
module matrixMult_N_M_1_N16_M32 ( clk, rst, x, y, o );
  input [511:0] x;
  input [8191:0] y;
  output [511:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N545, N546, N547, N548, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N673, N674, N675, N676, N677, N678, N679,
         N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690,
         N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701,
         N702, N703, N704, N737, N738, N739, N740, N741, N742, N743, N744,
         N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755,
         N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766,
         N767, N768, N801, N802, N803, N804, N805, N806, N807, N808, N809,
         N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885,
         N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N993,
         N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201,
         n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
         n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
         n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
         n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
         n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241,
         n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249,
         n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257,
         n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
         n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273,
         n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
         n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289,
         n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297,
         n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
         n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313,
         n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321,
         n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329,
         n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
         n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345,
         n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
         n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
         n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369,
         n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377,
         n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385,
         n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393,
         n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401,
         n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
         n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417,
         n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
         n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433,
         n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441,
         n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449,
         n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457,
         n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465,
         n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473,
         n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
         n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489,
         n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
         n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
         n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513,
         n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521,
         n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529,
         n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537,
         n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545,
         n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
         n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
         n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
         n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577,
         n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585,
         n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593,
         n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601,
         n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609,
         n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
         n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
         n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633,
         n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
         n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649,
         n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657,
         n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665,
         n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
         n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681,
         n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689,
         n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
         n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705,
         n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
         n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721,
         n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729,
         n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737,
         n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745,
         n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753,
         n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761,
         n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
         n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777,
         n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
         n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793,
         n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801,
         n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809,
         n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
         n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825,
         n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833,
         n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
         n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849,
         n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
         n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
         n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873,
         n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
         n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889,
         n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
         n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905,
         n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
         n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921,
         n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
         n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937,
         n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945,
         n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953,
         n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961,
         n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969,
         n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977,
         n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
         n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993,
         n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
         n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
         n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017,
         n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
         n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033,
         n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041,
         n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049,
         n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
         n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065,
         n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
         n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081,
         n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089,
         n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097,
         n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105,
         n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113,
         n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121,
         n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
         n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137,
         n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
         n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153,
         n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161,
         n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
         n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177,
         n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185,
         n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193,
         n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
         n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209,
         n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
         n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225,
         n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233,
         n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241,
         n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249,
         n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257,
         n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265,
         n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
         n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281,
         n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
         n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297,
         n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305,
         n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
         n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321,
         n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329,
         n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337,
         n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
         n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353,
         n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
         n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369,
         n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377,
         n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
         n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393,
         n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401,
         n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409,
         n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
         n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425,
         n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
         n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441,
         n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449,
         n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457,
         n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465,
         n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473,
         n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481,
         n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
         n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497,
         n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513,
         n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521,
         n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
         n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537,
         n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545,
         n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553,
         n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
         n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569,
         n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
         n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585,
         n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593,
         n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601,
         n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609,
         n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617,
         n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625,
         n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
         n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641,
         n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
         n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657,
         n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665,
         n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673,
         n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681,
         n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689,
         n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697,
         n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
         n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713,
         n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
         n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729,
         n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737,
         n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745,
         n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753,
         n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761,
         n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769,
         n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
         n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785,
         n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
         n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
         n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809,
         n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817,
         n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825,
         n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833,
         n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841,
         n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
         n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857,
         n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
         n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873,
         n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881,
         n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889,
         n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897,
         n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905,
         n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913,
         n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
         n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929,
         n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
         n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945,
         n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953,
         n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961,
         n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969,
         n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977,
         n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985,
         n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
         n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001,
         n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
         n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017,
         n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025,
         n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033,
         n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041,
         n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049,
         n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057,
         n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
         n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073,
         n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
         n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089,
         n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097,
         n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
         n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113,
         n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121,
         n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129,
         n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
         n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145,
         n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
         n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161,
         n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169,
         n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
         n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185,
         n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193,
         n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201,
         n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
         n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217,
         n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
         n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233,
         n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241,
         n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
         n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257,
         n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265,
         n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273,
         n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
         n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289,
         n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
         n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305,
         n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313,
         n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
         n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329,
         n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337,
         n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345,
         n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
         n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361,
         n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
         n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377,
         n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385,
         n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
         n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401,
         n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409,
         n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417,
         n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
         n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433,
         n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
         n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449,
         n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457,
         n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
         n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473,
         n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481,
         n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489,
         n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
         n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521,
         n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529,
         n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
         n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
         n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553,
         n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
         n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
         n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577,
         n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
         n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593,
         n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601,
         n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
         n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649,
         n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
         n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665,
         n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673,
         n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
         n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689,
         n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697,
         n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705,
         n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713,
         n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721,
         n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729,
         n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737,
         n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745,
         n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753,
         n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761,
         n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769,
         n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777,
         n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785,
         n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793,
         n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801,
         n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809,
         n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817,
         n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825,
         n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833,
         n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841,
         n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849,
         n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857,
         n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865,
         n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873,
         n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881,
         n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889,
         n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897,
         n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905,
         n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913,
         n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921,
         n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
         n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937,
         n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945,
         n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953,
         n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961,
         n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969,
         n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977,
         n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985,
         n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993,
         n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
         n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009,
         n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
         n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025,
         n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033,
         n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041,
         n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049,
         n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057,
         n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065,
         n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073,
         n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081,
         n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089,
         n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097,
         n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105,
         n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113,
         n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121,
         n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129,
         n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137,
         n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145,
         n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153,
         n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161,
         n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169,
         n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177,
         n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185,
         n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193,
         n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201,
         n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209,
         n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217,
         n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225,
         n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233,
         n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241,
         n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249,
         n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257,
         n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265,
         n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273,
         n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281,
         n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289,
         n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297,
         n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
         n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313,
         n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321,
         n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329,
         n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337,
         n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345,
         n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353,
         n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361,
         n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369,
         n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
         n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385,
         n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393,
         n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
         n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409,
         n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417,
         n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425,
         n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
         n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441,
         n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
         n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457,
         n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465,
         n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
         n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481,
         n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489,
         n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497,
         n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
         n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513,
         n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521,
         n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529,
         n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537,
         n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545,
         n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553,
         n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561,
         n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569,
         n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577,
         n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585,
         n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593,
         n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601,
         n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609,
         n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
         n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625,
         n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633,
         n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641,
         n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
         n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657,
         n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665,
         n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673,
         n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681,
         n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689,
         n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697,
         n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705,
         n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713,
         n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
         n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729,
         n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737,
         n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745,
         n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753,
         n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761,
         n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769,
         n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777,
         n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785,
         n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793,
         n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801,
         n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
         n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817,
         n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825,
         n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
         n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841,
         n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849,
         n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857,
         n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865,
         n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873,
         n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
         n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889,
         n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897,
         n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
         n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913,
         n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921,
         n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929,
         n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
         n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945,
         n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
         n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961,
         n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969,
         n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977,
         n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985,
         n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993,
         n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001,
         n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009,
         n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017,
         n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
         n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033,
         n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041,
         n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049,
         n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057,
         n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065,
         n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073,
         n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081,
         n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089,
         n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
         n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105,
         n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113,
         n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121,
         n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129,
         n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137,
         n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145,
         n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
         n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161,
         n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
         n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177,
         n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185,
         n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
         n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201,
         n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209,
         n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217,
         n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
         n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233,
         n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
         n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249,
         n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257,
         n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
         n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273,
         n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281,
         n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289,
         n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
         n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305,
         n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
         n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321,
         n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
         n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
         n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345,
         n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353,
         n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361,
         n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
         n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377,
         n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
         n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393,
         n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401,
         n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
         n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417,
         n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425,
         n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433,
         n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
         n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449,
         n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
         n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465,
         n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473,
         n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
         n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489,
         n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497,
         n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505,
         n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
         n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521,
         n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
         n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537,
         n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545,
         n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
         n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569,
         n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577,
         n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
         n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593,
         n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
         n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609,
         n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617,
         n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
         n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633,
         n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641,
         n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649,
         n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
         n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665,
         n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
         n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681,
         n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689,
         n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
         n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705,
         n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713,
         n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721,
         n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
         n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737,
         n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
         n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753,
         n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761,
         n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
         n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777,
         n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785,
         n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793,
         n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
         n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809,
         n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
         n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825,
         n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833,
         n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
         n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849,
         n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857,
         n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865,
         n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
         n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881,
         n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
         n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897,
         n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905,
         n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
         n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921,
         n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929,
         n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937,
         n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
         n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953,
         n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
         n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969,
         n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977,
         n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
         n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993,
         n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001,
         n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009,
         n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
         n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025,
         n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
         n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041,
         n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049,
         n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
         n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065,
         n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073,
         n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081,
         n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
         n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
         n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
         n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
         n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121,
         n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
         n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137,
         n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145,
         n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153,
         n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
         n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
         n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
         n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185,
         n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193,
         n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
         n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209,
         n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217,
         n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225,
         n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
         n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241,
         n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
         n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257,
         n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265,
         n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
         n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281,
         n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289,
         n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297,
         n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
         n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313,
         n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
         n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329,
         n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337,
         n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
         n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353,
         n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361,
         n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369,
         n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
         n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385,
         n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
         n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401,
         n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409,
         n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
         n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425,
         n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433,
         n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441,
         n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
         n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457,
         n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
         n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473,
         n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481,
         n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
         n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497,
         n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505,
         n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513,
         n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
         n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529,
         n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537,
         n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545,
         n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553,
         n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561,
         n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569,
         n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577,
         n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585,
         n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593,
         n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601,
         n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609,
         n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617,
         n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625,
         n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
         n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641,
         n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649,
         n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657,
         n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
         n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673,
         n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
         n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689,
         n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697,
         n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
         n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713,
         n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721,
         n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729,
         n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737,
         n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745,
         n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753,
         n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761,
         n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769,
         n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777,
         n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785,
         n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793,
         n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801,
         n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809,
         n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817,
         n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825,
         n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833,
         n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841,
         n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849,
         n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857,
         n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865,
         n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873,
         n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881,
         n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889,
         n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897,
         n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905,
         n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913,
         n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921,
         n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929,
         n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937,
         n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945,
         n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953,
         n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961,
         n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969,
         n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977,
         n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985,
         n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993,
         n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001,
         n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009,
         n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017,
         n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025,
         n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033,
         n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041,
         n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049,
         n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057,
         n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065,
         n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073,
         n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081,
         n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089,
         n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097,
         n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105,
         n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113,
         n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121,
         n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129,
         n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137,
         n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145,
         n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153,
         n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161,
         n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169,
         n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177,
         n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185,
         n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193,
         n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201,
         n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209,
         n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217,
         n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225,
         n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233,
         n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241,
         n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249,
         n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
         n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265,
         n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273,
         n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oi_reg[3][31]  ( .D(N256), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oi_reg[3][30]  ( .D(N255), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oi_reg[3][29]  ( .D(N254), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oi_reg[3][28]  ( .D(N253), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oi_reg[3][27]  ( .D(N252), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oi_reg[3][26]  ( .D(N251), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oi_reg[3][25]  ( .D(N250), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oi_reg[3][24]  ( .D(N249), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oi_reg[3][23]  ( .D(N248), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oi_reg[3][22]  ( .D(N247), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oi_reg[3][21]  ( .D(N246), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oi_reg[3][20]  ( .D(N245), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oi_reg[3][19]  ( .D(N244), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oi_reg[3][18]  ( .D(N243), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oi_reg[3][17]  ( .D(N242), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oi_reg[3][16]  ( .D(N241), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oi_reg[3][15]  ( .D(N240), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oi_reg[3][14]  ( .D(N239), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oi_reg[3][13]  ( .D(N238), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oi_reg[3][12]  ( .D(N237), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oi_reg[3][11]  ( .D(N236), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oi_reg[3][10]  ( .D(N235), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oi_reg[3][9]  ( .D(N234), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oi_reg[3][8]  ( .D(N233), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oi_reg[3][7]  ( .D(N232), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oi_reg[3][6]  ( .D(N231), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oi_reg[3][5]  ( .D(N230), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oi_reg[3][4]  ( .D(N229), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oi_reg[3][3]  ( .D(N228), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oi_reg[3][2]  ( .D(N227), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oi_reg[3][1]  ( .D(N226), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oi_reg[3][0]  ( .D(N225), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oi_reg[4][31]  ( .D(N320), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oi_reg[4][30]  ( .D(N319), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oi_reg[4][29]  ( .D(N318), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oi_reg[4][28]  ( .D(N317), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oi_reg[4][27]  ( .D(N316), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oi_reg[4][26]  ( .D(N315), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oi_reg[4][25]  ( .D(N314), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oi_reg[4][24]  ( .D(N313), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oi_reg[4][23]  ( .D(N312), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oi_reg[4][22]  ( .D(N311), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oi_reg[4][21]  ( .D(N310), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oi_reg[4][20]  ( .D(N309), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oi_reg[4][19]  ( .D(N308), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oi_reg[4][18]  ( .D(N307), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oi_reg[4][17]  ( .D(N306), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oi_reg[4][16]  ( .D(N305), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oi_reg[4][15]  ( .D(N304), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oi_reg[4][14]  ( .D(N303), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oi_reg[4][13]  ( .D(N302), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oi_reg[4][12]  ( .D(N301), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oi_reg[4][11]  ( .D(N300), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oi_reg[4][10]  ( .D(N299), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oi_reg[4][9]  ( .D(N298), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oi_reg[4][8]  ( .D(N297), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oi_reg[4][7]  ( .D(N296), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oi_reg[4][6]  ( .D(N295), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oi_reg[4][5]  ( .D(N294), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oi_reg[4][4]  ( .D(N293), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oi_reg[4][3]  ( .D(N292), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oi_reg[4][2]  ( .D(N291), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oi_reg[4][1]  ( .D(N290), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oi_reg[4][0]  ( .D(N289), .CLK(clk), .RST(rst), .Q(o[128]) );
  DFF \oi_reg[5][31]  ( .D(N384), .CLK(clk), .RST(rst), .Q(o[191]) );
  DFF \oi_reg[5][30]  ( .D(N383), .CLK(clk), .RST(rst), .Q(o[190]) );
  DFF \oi_reg[5][29]  ( .D(N382), .CLK(clk), .RST(rst), .Q(o[189]) );
  DFF \oi_reg[5][28]  ( .D(N381), .CLK(clk), .RST(rst), .Q(o[188]) );
  DFF \oi_reg[5][27]  ( .D(N380), .CLK(clk), .RST(rst), .Q(o[187]) );
  DFF \oi_reg[5][26]  ( .D(N379), .CLK(clk), .RST(rst), .Q(o[186]) );
  DFF \oi_reg[5][25]  ( .D(N378), .CLK(clk), .RST(rst), .Q(o[185]) );
  DFF \oi_reg[5][24]  ( .D(N377), .CLK(clk), .RST(rst), .Q(o[184]) );
  DFF \oi_reg[5][23]  ( .D(N376), .CLK(clk), .RST(rst), .Q(o[183]) );
  DFF \oi_reg[5][22]  ( .D(N375), .CLK(clk), .RST(rst), .Q(o[182]) );
  DFF \oi_reg[5][21]  ( .D(N374), .CLK(clk), .RST(rst), .Q(o[181]) );
  DFF \oi_reg[5][20]  ( .D(N373), .CLK(clk), .RST(rst), .Q(o[180]) );
  DFF \oi_reg[5][19]  ( .D(N372), .CLK(clk), .RST(rst), .Q(o[179]) );
  DFF \oi_reg[5][18]  ( .D(N371), .CLK(clk), .RST(rst), .Q(o[178]) );
  DFF \oi_reg[5][17]  ( .D(N370), .CLK(clk), .RST(rst), .Q(o[177]) );
  DFF \oi_reg[5][16]  ( .D(N369), .CLK(clk), .RST(rst), .Q(o[176]) );
  DFF \oi_reg[5][15]  ( .D(N368), .CLK(clk), .RST(rst), .Q(o[175]) );
  DFF \oi_reg[5][14]  ( .D(N367), .CLK(clk), .RST(rst), .Q(o[174]) );
  DFF \oi_reg[5][13]  ( .D(N366), .CLK(clk), .RST(rst), .Q(o[173]) );
  DFF \oi_reg[5][12]  ( .D(N365), .CLK(clk), .RST(rst), .Q(o[172]) );
  DFF \oi_reg[5][11]  ( .D(N364), .CLK(clk), .RST(rst), .Q(o[171]) );
  DFF \oi_reg[5][10]  ( .D(N363), .CLK(clk), .RST(rst), .Q(o[170]) );
  DFF \oi_reg[5][9]  ( .D(N362), .CLK(clk), .RST(rst), .Q(o[169]) );
  DFF \oi_reg[5][8]  ( .D(N361), .CLK(clk), .RST(rst), .Q(o[168]) );
  DFF \oi_reg[5][7]  ( .D(N360), .CLK(clk), .RST(rst), .Q(o[167]) );
  DFF \oi_reg[5][6]  ( .D(N359), .CLK(clk), .RST(rst), .Q(o[166]) );
  DFF \oi_reg[5][5]  ( .D(N358), .CLK(clk), .RST(rst), .Q(o[165]) );
  DFF \oi_reg[5][4]  ( .D(N357), .CLK(clk), .RST(rst), .Q(o[164]) );
  DFF \oi_reg[5][3]  ( .D(N356), .CLK(clk), .RST(rst), .Q(o[163]) );
  DFF \oi_reg[5][2]  ( .D(N355), .CLK(clk), .RST(rst), .Q(o[162]) );
  DFF \oi_reg[5][1]  ( .D(N354), .CLK(clk), .RST(rst), .Q(o[161]) );
  DFF \oi_reg[5][0]  ( .D(N353), .CLK(clk), .RST(rst), .Q(o[160]) );
  DFF \oi_reg[6][31]  ( .D(N448), .CLK(clk), .RST(rst), .Q(o[223]) );
  DFF \oi_reg[6][30]  ( .D(N447), .CLK(clk), .RST(rst), .Q(o[222]) );
  DFF \oi_reg[6][29]  ( .D(N446), .CLK(clk), .RST(rst), .Q(o[221]) );
  DFF \oi_reg[6][28]  ( .D(N445), .CLK(clk), .RST(rst), .Q(o[220]) );
  DFF \oi_reg[6][27]  ( .D(N444), .CLK(clk), .RST(rst), .Q(o[219]) );
  DFF \oi_reg[6][26]  ( .D(N443), .CLK(clk), .RST(rst), .Q(o[218]) );
  DFF \oi_reg[6][25]  ( .D(N442), .CLK(clk), .RST(rst), .Q(o[217]) );
  DFF \oi_reg[6][24]  ( .D(N441), .CLK(clk), .RST(rst), .Q(o[216]) );
  DFF \oi_reg[6][23]  ( .D(N440), .CLK(clk), .RST(rst), .Q(o[215]) );
  DFF \oi_reg[6][22]  ( .D(N439), .CLK(clk), .RST(rst), .Q(o[214]) );
  DFF \oi_reg[6][21]  ( .D(N438), .CLK(clk), .RST(rst), .Q(o[213]) );
  DFF \oi_reg[6][20]  ( .D(N437), .CLK(clk), .RST(rst), .Q(o[212]) );
  DFF \oi_reg[6][19]  ( .D(N436), .CLK(clk), .RST(rst), .Q(o[211]) );
  DFF \oi_reg[6][18]  ( .D(N435), .CLK(clk), .RST(rst), .Q(o[210]) );
  DFF \oi_reg[6][17]  ( .D(N434), .CLK(clk), .RST(rst), .Q(o[209]) );
  DFF \oi_reg[6][16]  ( .D(N433), .CLK(clk), .RST(rst), .Q(o[208]) );
  DFF \oi_reg[6][15]  ( .D(N432), .CLK(clk), .RST(rst), .Q(o[207]) );
  DFF \oi_reg[6][14]  ( .D(N431), .CLK(clk), .RST(rst), .Q(o[206]) );
  DFF \oi_reg[6][13]  ( .D(N430), .CLK(clk), .RST(rst), .Q(o[205]) );
  DFF \oi_reg[6][12]  ( .D(N429), .CLK(clk), .RST(rst), .Q(o[204]) );
  DFF \oi_reg[6][11]  ( .D(N428), .CLK(clk), .RST(rst), .Q(o[203]) );
  DFF \oi_reg[6][10]  ( .D(N427), .CLK(clk), .RST(rst), .Q(o[202]) );
  DFF \oi_reg[6][9]  ( .D(N426), .CLK(clk), .RST(rst), .Q(o[201]) );
  DFF \oi_reg[6][8]  ( .D(N425), .CLK(clk), .RST(rst), .Q(o[200]) );
  DFF \oi_reg[6][7]  ( .D(N424), .CLK(clk), .RST(rst), .Q(o[199]) );
  DFF \oi_reg[6][6]  ( .D(N423), .CLK(clk), .RST(rst), .Q(o[198]) );
  DFF \oi_reg[6][5]  ( .D(N422), .CLK(clk), .RST(rst), .Q(o[197]) );
  DFF \oi_reg[6][4]  ( .D(N421), .CLK(clk), .RST(rst), .Q(o[196]) );
  DFF \oi_reg[6][3]  ( .D(N420), .CLK(clk), .RST(rst), .Q(o[195]) );
  DFF \oi_reg[6][2]  ( .D(N419), .CLK(clk), .RST(rst), .Q(o[194]) );
  DFF \oi_reg[6][1]  ( .D(N418), .CLK(clk), .RST(rst), .Q(o[193]) );
  DFF \oi_reg[6][0]  ( .D(N417), .CLK(clk), .RST(rst), .Q(o[192]) );
  DFF \oi_reg[7][31]  ( .D(N512), .CLK(clk), .RST(rst), .Q(o[255]) );
  DFF \oi_reg[7][30]  ( .D(N511), .CLK(clk), .RST(rst), .Q(o[254]) );
  DFF \oi_reg[7][29]  ( .D(N510), .CLK(clk), .RST(rst), .Q(o[253]) );
  DFF \oi_reg[7][28]  ( .D(N509), .CLK(clk), .RST(rst), .Q(o[252]) );
  DFF \oi_reg[7][27]  ( .D(N508), .CLK(clk), .RST(rst), .Q(o[251]) );
  DFF \oi_reg[7][26]  ( .D(N507), .CLK(clk), .RST(rst), .Q(o[250]) );
  DFF \oi_reg[7][25]  ( .D(N506), .CLK(clk), .RST(rst), .Q(o[249]) );
  DFF \oi_reg[7][24]  ( .D(N505), .CLK(clk), .RST(rst), .Q(o[248]) );
  DFF \oi_reg[7][23]  ( .D(N504), .CLK(clk), .RST(rst), .Q(o[247]) );
  DFF \oi_reg[7][22]  ( .D(N503), .CLK(clk), .RST(rst), .Q(o[246]) );
  DFF \oi_reg[7][21]  ( .D(N502), .CLK(clk), .RST(rst), .Q(o[245]) );
  DFF \oi_reg[7][20]  ( .D(N501), .CLK(clk), .RST(rst), .Q(o[244]) );
  DFF \oi_reg[7][19]  ( .D(N500), .CLK(clk), .RST(rst), .Q(o[243]) );
  DFF \oi_reg[7][18]  ( .D(N499), .CLK(clk), .RST(rst), .Q(o[242]) );
  DFF \oi_reg[7][17]  ( .D(N498), .CLK(clk), .RST(rst), .Q(o[241]) );
  DFF \oi_reg[7][16]  ( .D(N497), .CLK(clk), .RST(rst), .Q(o[240]) );
  DFF \oi_reg[7][15]  ( .D(N496), .CLK(clk), .RST(rst), .Q(o[239]) );
  DFF \oi_reg[7][14]  ( .D(N495), .CLK(clk), .RST(rst), .Q(o[238]) );
  DFF \oi_reg[7][13]  ( .D(N494), .CLK(clk), .RST(rst), .Q(o[237]) );
  DFF \oi_reg[7][12]  ( .D(N493), .CLK(clk), .RST(rst), .Q(o[236]) );
  DFF \oi_reg[7][11]  ( .D(N492), .CLK(clk), .RST(rst), .Q(o[235]) );
  DFF \oi_reg[7][10]  ( .D(N491), .CLK(clk), .RST(rst), .Q(o[234]) );
  DFF \oi_reg[7][9]  ( .D(N490), .CLK(clk), .RST(rst), .Q(o[233]) );
  DFF \oi_reg[7][8]  ( .D(N489), .CLK(clk), .RST(rst), .Q(o[232]) );
  DFF \oi_reg[7][7]  ( .D(N488), .CLK(clk), .RST(rst), .Q(o[231]) );
  DFF \oi_reg[7][6]  ( .D(N487), .CLK(clk), .RST(rst), .Q(o[230]) );
  DFF \oi_reg[7][5]  ( .D(N486), .CLK(clk), .RST(rst), .Q(o[229]) );
  DFF \oi_reg[7][4]  ( .D(N485), .CLK(clk), .RST(rst), .Q(o[228]) );
  DFF \oi_reg[7][3]  ( .D(N484), .CLK(clk), .RST(rst), .Q(o[227]) );
  DFF \oi_reg[7][2]  ( .D(N483), .CLK(clk), .RST(rst), .Q(o[226]) );
  DFF \oi_reg[7][1]  ( .D(N482), .CLK(clk), .RST(rst), .Q(o[225]) );
  DFF \oi_reg[7][0]  ( .D(N481), .CLK(clk), .RST(rst), .Q(o[224]) );
  DFF \oi_reg[8][31]  ( .D(N576), .CLK(clk), .RST(rst), .Q(o[287]) );
  DFF \oi_reg[8][30]  ( .D(N575), .CLK(clk), .RST(rst), .Q(o[286]) );
  DFF \oi_reg[8][29]  ( .D(N574), .CLK(clk), .RST(rst), .Q(o[285]) );
  DFF \oi_reg[8][28]  ( .D(N573), .CLK(clk), .RST(rst), .Q(o[284]) );
  DFF \oi_reg[8][27]  ( .D(N572), .CLK(clk), .RST(rst), .Q(o[283]) );
  DFF \oi_reg[8][26]  ( .D(N571), .CLK(clk), .RST(rst), .Q(o[282]) );
  DFF \oi_reg[8][25]  ( .D(N570), .CLK(clk), .RST(rst), .Q(o[281]) );
  DFF \oi_reg[8][24]  ( .D(N569), .CLK(clk), .RST(rst), .Q(o[280]) );
  DFF \oi_reg[8][23]  ( .D(N568), .CLK(clk), .RST(rst), .Q(o[279]) );
  DFF \oi_reg[8][22]  ( .D(N567), .CLK(clk), .RST(rst), .Q(o[278]) );
  DFF \oi_reg[8][21]  ( .D(N566), .CLK(clk), .RST(rst), .Q(o[277]) );
  DFF \oi_reg[8][20]  ( .D(N565), .CLK(clk), .RST(rst), .Q(o[276]) );
  DFF \oi_reg[8][19]  ( .D(N564), .CLK(clk), .RST(rst), .Q(o[275]) );
  DFF \oi_reg[8][18]  ( .D(N563), .CLK(clk), .RST(rst), .Q(o[274]) );
  DFF \oi_reg[8][17]  ( .D(N562), .CLK(clk), .RST(rst), .Q(o[273]) );
  DFF \oi_reg[8][16]  ( .D(N561), .CLK(clk), .RST(rst), .Q(o[272]) );
  DFF \oi_reg[8][15]  ( .D(N560), .CLK(clk), .RST(rst), .Q(o[271]) );
  DFF \oi_reg[8][14]  ( .D(N559), .CLK(clk), .RST(rst), .Q(o[270]) );
  DFF \oi_reg[8][13]  ( .D(N558), .CLK(clk), .RST(rst), .Q(o[269]) );
  DFF \oi_reg[8][12]  ( .D(N557), .CLK(clk), .RST(rst), .Q(o[268]) );
  DFF \oi_reg[8][11]  ( .D(N556), .CLK(clk), .RST(rst), .Q(o[267]) );
  DFF \oi_reg[8][10]  ( .D(N555), .CLK(clk), .RST(rst), .Q(o[266]) );
  DFF \oi_reg[8][9]  ( .D(N554), .CLK(clk), .RST(rst), .Q(o[265]) );
  DFF \oi_reg[8][8]  ( .D(N553), .CLK(clk), .RST(rst), .Q(o[264]) );
  DFF \oi_reg[8][7]  ( .D(N552), .CLK(clk), .RST(rst), .Q(o[263]) );
  DFF \oi_reg[8][6]  ( .D(N551), .CLK(clk), .RST(rst), .Q(o[262]) );
  DFF \oi_reg[8][5]  ( .D(N550), .CLK(clk), .RST(rst), .Q(o[261]) );
  DFF \oi_reg[8][4]  ( .D(N549), .CLK(clk), .RST(rst), .Q(o[260]) );
  DFF \oi_reg[8][3]  ( .D(N548), .CLK(clk), .RST(rst), .Q(o[259]) );
  DFF \oi_reg[8][2]  ( .D(N547), .CLK(clk), .RST(rst), .Q(o[258]) );
  DFF \oi_reg[8][1]  ( .D(N546), .CLK(clk), .RST(rst), .Q(o[257]) );
  DFF \oi_reg[8][0]  ( .D(N545), .CLK(clk), .RST(rst), .Q(o[256]) );
  DFF \oi_reg[9][31]  ( .D(N640), .CLK(clk), .RST(rst), .Q(o[319]) );
  DFF \oi_reg[9][30]  ( .D(N639), .CLK(clk), .RST(rst), .Q(o[318]) );
  DFF \oi_reg[9][29]  ( .D(N638), .CLK(clk), .RST(rst), .Q(o[317]) );
  DFF \oi_reg[9][28]  ( .D(N637), .CLK(clk), .RST(rst), .Q(o[316]) );
  DFF \oi_reg[9][27]  ( .D(N636), .CLK(clk), .RST(rst), .Q(o[315]) );
  DFF \oi_reg[9][26]  ( .D(N635), .CLK(clk), .RST(rst), .Q(o[314]) );
  DFF \oi_reg[9][25]  ( .D(N634), .CLK(clk), .RST(rst), .Q(o[313]) );
  DFF \oi_reg[9][24]  ( .D(N633), .CLK(clk), .RST(rst), .Q(o[312]) );
  DFF \oi_reg[9][23]  ( .D(N632), .CLK(clk), .RST(rst), .Q(o[311]) );
  DFF \oi_reg[9][22]  ( .D(N631), .CLK(clk), .RST(rst), .Q(o[310]) );
  DFF \oi_reg[9][21]  ( .D(N630), .CLK(clk), .RST(rst), .Q(o[309]) );
  DFF \oi_reg[9][20]  ( .D(N629), .CLK(clk), .RST(rst), .Q(o[308]) );
  DFF \oi_reg[9][19]  ( .D(N628), .CLK(clk), .RST(rst), .Q(o[307]) );
  DFF \oi_reg[9][18]  ( .D(N627), .CLK(clk), .RST(rst), .Q(o[306]) );
  DFF \oi_reg[9][17]  ( .D(N626), .CLK(clk), .RST(rst), .Q(o[305]) );
  DFF \oi_reg[9][16]  ( .D(N625), .CLK(clk), .RST(rst), .Q(o[304]) );
  DFF \oi_reg[9][15]  ( .D(N624), .CLK(clk), .RST(rst), .Q(o[303]) );
  DFF \oi_reg[9][14]  ( .D(N623), .CLK(clk), .RST(rst), .Q(o[302]) );
  DFF \oi_reg[9][13]  ( .D(N622), .CLK(clk), .RST(rst), .Q(o[301]) );
  DFF \oi_reg[9][12]  ( .D(N621), .CLK(clk), .RST(rst), .Q(o[300]) );
  DFF \oi_reg[9][11]  ( .D(N620), .CLK(clk), .RST(rst), .Q(o[299]) );
  DFF \oi_reg[9][10]  ( .D(N619), .CLK(clk), .RST(rst), .Q(o[298]) );
  DFF \oi_reg[9][9]  ( .D(N618), .CLK(clk), .RST(rst), .Q(o[297]) );
  DFF \oi_reg[9][8]  ( .D(N617), .CLK(clk), .RST(rst), .Q(o[296]) );
  DFF \oi_reg[9][7]  ( .D(N616), .CLK(clk), .RST(rst), .Q(o[295]) );
  DFF \oi_reg[9][6]  ( .D(N615), .CLK(clk), .RST(rst), .Q(o[294]) );
  DFF \oi_reg[9][5]  ( .D(N614), .CLK(clk), .RST(rst), .Q(o[293]) );
  DFF \oi_reg[9][4]  ( .D(N613), .CLK(clk), .RST(rst), .Q(o[292]) );
  DFF \oi_reg[9][3]  ( .D(N612), .CLK(clk), .RST(rst), .Q(o[291]) );
  DFF \oi_reg[9][2]  ( .D(N611), .CLK(clk), .RST(rst), .Q(o[290]) );
  DFF \oi_reg[9][1]  ( .D(N610), .CLK(clk), .RST(rst), .Q(o[289]) );
  DFF \oi_reg[9][0]  ( .D(N609), .CLK(clk), .RST(rst), .Q(o[288]) );
  DFF \oi_reg[10][31]  ( .D(N704), .CLK(clk), .RST(rst), .Q(o[351]) );
  DFF \oi_reg[10][30]  ( .D(N703), .CLK(clk), .RST(rst), .Q(o[350]) );
  DFF \oi_reg[10][29]  ( .D(N702), .CLK(clk), .RST(rst), .Q(o[349]) );
  DFF \oi_reg[10][28]  ( .D(N701), .CLK(clk), .RST(rst), .Q(o[348]) );
  DFF \oi_reg[10][27]  ( .D(N700), .CLK(clk), .RST(rst), .Q(o[347]) );
  DFF \oi_reg[10][26]  ( .D(N699), .CLK(clk), .RST(rst), .Q(o[346]) );
  DFF \oi_reg[10][25]  ( .D(N698), .CLK(clk), .RST(rst), .Q(o[345]) );
  DFF \oi_reg[10][24]  ( .D(N697), .CLK(clk), .RST(rst), .Q(o[344]) );
  DFF \oi_reg[10][23]  ( .D(N696), .CLK(clk), .RST(rst), .Q(o[343]) );
  DFF \oi_reg[10][22]  ( .D(N695), .CLK(clk), .RST(rst), .Q(o[342]) );
  DFF \oi_reg[10][21]  ( .D(N694), .CLK(clk), .RST(rst), .Q(o[341]) );
  DFF \oi_reg[10][20]  ( .D(N693), .CLK(clk), .RST(rst), .Q(o[340]) );
  DFF \oi_reg[10][19]  ( .D(N692), .CLK(clk), .RST(rst), .Q(o[339]) );
  DFF \oi_reg[10][18]  ( .D(N691), .CLK(clk), .RST(rst), .Q(o[338]) );
  DFF \oi_reg[10][17]  ( .D(N690), .CLK(clk), .RST(rst), .Q(o[337]) );
  DFF \oi_reg[10][16]  ( .D(N689), .CLK(clk), .RST(rst), .Q(o[336]) );
  DFF \oi_reg[10][15]  ( .D(N688), .CLK(clk), .RST(rst), .Q(o[335]) );
  DFF \oi_reg[10][14]  ( .D(N687), .CLK(clk), .RST(rst), .Q(o[334]) );
  DFF \oi_reg[10][13]  ( .D(N686), .CLK(clk), .RST(rst), .Q(o[333]) );
  DFF \oi_reg[10][12]  ( .D(N685), .CLK(clk), .RST(rst), .Q(o[332]) );
  DFF \oi_reg[10][11]  ( .D(N684), .CLK(clk), .RST(rst), .Q(o[331]) );
  DFF \oi_reg[10][10]  ( .D(N683), .CLK(clk), .RST(rst), .Q(o[330]) );
  DFF \oi_reg[10][9]  ( .D(N682), .CLK(clk), .RST(rst), .Q(o[329]) );
  DFF \oi_reg[10][8]  ( .D(N681), .CLK(clk), .RST(rst), .Q(o[328]) );
  DFF \oi_reg[10][7]  ( .D(N680), .CLK(clk), .RST(rst), .Q(o[327]) );
  DFF \oi_reg[10][6]  ( .D(N679), .CLK(clk), .RST(rst), .Q(o[326]) );
  DFF \oi_reg[10][5]  ( .D(N678), .CLK(clk), .RST(rst), .Q(o[325]) );
  DFF \oi_reg[10][4]  ( .D(N677), .CLK(clk), .RST(rst), .Q(o[324]) );
  DFF \oi_reg[10][3]  ( .D(N676), .CLK(clk), .RST(rst), .Q(o[323]) );
  DFF \oi_reg[10][2]  ( .D(N675), .CLK(clk), .RST(rst), .Q(o[322]) );
  DFF \oi_reg[10][1]  ( .D(N674), .CLK(clk), .RST(rst), .Q(o[321]) );
  DFF \oi_reg[10][0]  ( .D(N673), .CLK(clk), .RST(rst), .Q(o[320]) );
  DFF \oi_reg[11][31]  ( .D(N768), .CLK(clk), .RST(rst), .Q(o[383]) );
  DFF \oi_reg[11][30]  ( .D(N767), .CLK(clk), .RST(rst), .Q(o[382]) );
  DFF \oi_reg[11][29]  ( .D(N766), .CLK(clk), .RST(rst), .Q(o[381]) );
  DFF \oi_reg[11][28]  ( .D(N765), .CLK(clk), .RST(rst), .Q(o[380]) );
  DFF \oi_reg[11][27]  ( .D(N764), .CLK(clk), .RST(rst), .Q(o[379]) );
  DFF \oi_reg[11][26]  ( .D(N763), .CLK(clk), .RST(rst), .Q(o[378]) );
  DFF \oi_reg[11][25]  ( .D(N762), .CLK(clk), .RST(rst), .Q(o[377]) );
  DFF \oi_reg[11][24]  ( .D(N761), .CLK(clk), .RST(rst), .Q(o[376]) );
  DFF \oi_reg[11][23]  ( .D(N760), .CLK(clk), .RST(rst), .Q(o[375]) );
  DFF \oi_reg[11][22]  ( .D(N759), .CLK(clk), .RST(rst), .Q(o[374]) );
  DFF \oi_reg[11][21]  ( .D(N758), .CLK(clk), .RST(rst), .Q(o[373]) );
  DFF \oi_reg[11][20]  ( .D(N757), .CLK(clk), .RST(rst), .Q(o[372]) );
  DFF \oi_reg[11][19]  ( .D(N756), .CLK(clk), .RST(rst), .Q(o[371]) );
  DFF \oi_reg[11][18]  ( .D(N755), .CLK(clk), .RST(rst), .Q(o[370]) );
  DFF \oi_reg[11][17]  ( .D(N754), .CLK(clk), .RST(rst), .Q(o[369]) );
  DFF \oi_reg[11][16]  ( .D(N753), .CLK(clk), .RST(rst), .Q(o[368]) );
  DFF \oi_reg[11][15]  ( .D(N752), .CLK(clk), .RST(rst), .Q(o[367]) );
  DFF \oi_reg[11][14]  ( .D(N751), .CLK(clk), .RST(rst), .Q(o[366]) );
  DFF \oi_reg[11][13]  ( .D(N750), .CLK(clk), .RST(rst), .Q(o[365]) );
  DFF \oi_reg[11][12]  ( .D(N749), .CLK(clk), .RST(rst), .Q(o[364]) );
  DFF \oi_reg[11][11]  ( .D(N748), .CLK(clk), .RST(rst), .Q(o[363]) );
  DFF \oi_reg[11][10]  ( .D(N747), .CLK(clk), .RST(rst), .Q(o[362]) );
  DFF \oi_reg[11][9]  ( .D(N746), .CLK(clk), .RST(rst), .Q(o[361]) );
  DFF \oi_reg[11][8]  ( .D(N745), .CLK(clk), .RST(rst), .Q(o[360]) );
  DFF \oi_reg[11][7]  ( .D(N744), .CLK(clk), .RST(rst), .Q(o[359]) );
  DFF \oi_reg[11][6]  ( .D(N743), .CLK(clk), .RST(rst), .Q(o[358]) );
  DFF \oi_reg[11][5]  ( .D(N742), .CLK(clk), .RST(rst), .Q(o[357]) );
  DFF \oi_reg[11][4]  ( .D(N741), .CLK(clk), .RST(rst), .Q(o[356]) );
  DFF \oi_reg[11][3]  ( .D(N740), .CLK(clk), .RST(rst), .Q(o[355]) );
  DFF \oi_reg[11][2]  ( .D(N739), .CLK(clk), .RST(rst), .Q(o[354]) );
  DFF \oi_reg[11][1]  ( .D(N738), .CLK(clk), .RST(rst), .Q(o[353]) );
  DFF \oi_reg[11][0]  ( .D(N737), .CLK(clk), .RST(rst), .Q(o[352]) );
  DFF \oi_reg[12][31]  ( .D(N832), .CLK(clk), .RST(rst), .Q(o[415]) );
  DFF \oi_reg[12][30]  ( .D(N831), .CLK(clk), .RST(rst), .Q(o[414]) );
  DFF \oi_reg[12][29]  ( .D(N830), .CLK(clk), .RST(rst), .Q(o[413]) );
  DFF \oi_reg[12][28]  ( .D(N829), .CLK(clk), .RST(rst), .Q(o[412]) );
  DFF \oi_reg[12][27]  ( .D(N828), .CLK(clk), .RST(rst), .Q(o[411]) );
  DFF \oi_reg[12][26]  ( .D(N827), .CLK(clk), .RST(rst), .Q(o[410]) );
  DFF \oi_reg[12][25]  ( .D(N826), .CLK(clk), .RST(rst), .Q(o[409]) );
  DFF \oi_reg[12][24]  ( .D(N825), .CLK(clk), .RST(rst), .Q(o[408]) );
  DFF \oi_reg[12][23]  ( .D(N824), .CLK(clk), .RST(rst), .Q(o[407]) );
  DFF \oi_reg[12][22]  ( .D(N823), .CLK(clk), .RST(rst), .Q(o[406]) );
  DFF \oi_reg[12][21]  ( .D(N822), .CLK(clk), .RST(rst), .Q(o[405]) );
  DFF \oi_reg[12][20]  ( .D(N821), .CLK(clk), .RST(rst), .Q(o[404]) );
  DFF \oi_reg[12][19]  ( .D(N820), .CLK(clk), .RST(rst), .Q(o[403]) );
  DFF \oi_reg[12][18]  ( .D(N819), .CLK(clk), .RST(rst), .Q(o[402]) );
  DFF \oi_reg[12][17]  ( .D(N818), .CLK(clk), .RST(rst), .Q(o[401]) );
  DFF \oi_reg[12][16]  ( .D(N817), .CLK(clk), .RST(rst), .Q(o[400]) );
  DFF \oi_reg[12][15]  ( .D(N816), .CLK(clk), .RST(rst), .Q(o[399]) );
  DFF \oi_reg[12][14]  ( .D(N815), .CLK(clk), .RST(rst), .Q(o[398]) );
  DFF \oi_reg[12][13]  ( .D(N814), .CLK(clk), .RST(rst), .Q(o[397]) );
  DFF \oi_reg[12][12]  ( .D(N813), .CLK(clk), .RST(rst), .Q(o[396]) );
  DFF \oi_reg[12][11]  ( .D(N812), .CLK(clk), .RST(rst), .Q(o[395]) );
  DFF \oi_reg[12][10]  ( .D(N811), .CLK(clk), .RST(rst), .Q(o[394]) );
  DFF \oi_reg[12][9]  ( .D(N810), .CLK(clk), .RST(rst), .Q(o[393]) );
  DFF \oi_reg[12][8]  ( .D(N809), .CLK(clk), .RST(rst), .Q(o[392]) );
  DFF \oi_reg[12][7]  ( .D(N808), .CLK(clk), .RST(rst), .Q(o[391]) );
  DFF \oi_reg[12][6]  ( .D(N807), .CLK(clk), .RST(rst), .Q(o[390]) );
  DFF \oi_reg[12][5]  ( .D(N806), .CLK(clk), .RST(rst), .Q(o[389]) );
  DFF \oi_reg[12][4]  ( .D(N805), .CLK(clk), .RST(rst), .Q(o[388]) );
  DFF \oi_reg[12][3]  ( .D(N804), .CLK(clk), .RST(rst), .Q(o[387]) );
  DFF \oi_reg[12][2]  ( .D(N803), .CLK(clk), .RST(rst), .Q(o[386]) );
  DFF \oi_reg[12][1]  ( .D(N802), .CLK(clk), .RST(rst), .Q(o[385]) );
  DFF \oi_reg[12][0]  ( .D(N801), .CLK(clk), .RST(rst), .Q(o[384]) );
  DFF \oi_reg[13][31]  ( .D(N896), .CLK(clk), .RST(rst), .Q(o[447]) );
  DFF \oi_reg[13][30]  ( .D(N895), .CLK(clk), .RST(rst), .Q(o[446]) );
  DFF \oi_reg[13][29]  ( .D(N894), .CLK(clk), .RST(rst), .Q(o[445]) );
  DFF \oi_reg[13][28]  ( .D(N893), .CLK(clk), .RST(rst), .Q(o[444]) );
  DFF \oi_reg[13][27]  ( .D(N892), .CLK(clk), .RST(rst), .Q(o[443]) );
  DFF \oi_reg[13][26]  ( .D(N891), .CLK(clk), .RST(rst), .Q(o[442]) );
  DFF \oi_reg[13][25]  ( .D(N890), .CLK(clk), .RST(rst), .Q(o[441]) );
  DFF \oi_reg[13][24]  ( .D(N889), .CLK(clk), .RST(rst), .Q(o[440]) );
  DFF \oi_reg[13][23]  ( .D(N888), .CLK(clk), .RST(rst), .Q(o[439]) );
  DFF \oi_reg[13][22]  ( .D(N887), .CLK(clk), .RST(rst), .Q(o[438]) );
  DFF \oi_reg[13][21]  ( .D(N886), .CLK(clk), .RST(rst), .Q(o[437]) );
  DFF \oi_reg[13][20]  ( .D(N885), .CLK(clk), .RST(rst), .Q(o[436]) );
  DFF \oi_reg[13][19]  ( .D(N884), .CLK(clk), .RST(rst), .Q(o[435]) );
  DFF \oi_reg[13][18]  ( .D(N883), .CLK(clk), .RST(rst), .Q(o[434]) );
  DFF \oi_reg[13][17]  ( .D(N882), .CLK(clk), .RST(rst), .Q(o[433]) );
  DFF \oi_reg[13][16]  ( .D(N881), .CLK(clk), .RST(rst), .Q(o[432]) );
  DFF \oi_reg[13][15]  ( .D(N880), .CLK(clk), .RST(rst), .Q(o[431]) );
  DFF \oi_reg[13][14]  ( .D(N879), .CLK(clk), .RST(rst), .Q(o[430]) );
  DFF \oi_reg[13][13]  ( .D(N878), .CLK(clk), .RST(rst), .Q(o[429]) );
  DFF \oi_reg[13][12]  ( .D(N877), .CLK(clk), .RST(rst), .Q(o[428]) );
  DFF \oi_reg[13][11]  ( .D(N876), .CLK(clk), .RST(rst), .Q(o[427]) );
  DFF \oi_reg[13][10]  ( .D(N875), .CLK(clk), .RST(rst), .Q(o[426]) );
  DFF \oi_reg[13][9]  ( .D(N874), .CLK(clk), .RST(rst), .Q(o[425]) );
  DFF \oi_reg[13][8]  ( .D(N873), .CLK(clk), .RST(rst), .Q(o[424]) );
  DFF \oi_reg[13][7]  ( .D(N872), .CLK(clk), .RST(rst), .Q(o[423]) );
  DFF \oi_reg[13][6]  ( .D(N871), .CLK(clk), .RST(rst), .Q(o[422]) );
  DFF \oi_reg[13][5]  ( .D(N870), .CLK(clk), .RST(rst), .Q(o[421]) );
  DFF \oi_reg[13][4]  ( .D(N869), .CLK(clk), .RST(rst), .Q(o[420]) );
  DFF \oi_reg[13][3]  ( .D(N868), .CLK(clk), .RST(rst), .Q(o[419]) );
  DFF \oi_reg[13][2]  ( .D(N867), .CLK(clk), .RST(rst), .Q(o[418]) );
  DFF \oi_reg[13][1]  ( .D(N866), .CLK(clk), .RST(rst), .Q(o[417]) );
  DFF \oi_reg[13][0]  ( .D(N865), .CLK(clk), .RST(rst), .Q(o[416]) );
  DFF \oi_reg[14][31]  ( .D(N960), .CLK(clk), .RST(rst), .Q(o[479]) );
  DFF \oi_reg[14][30]  ( .D(N959), .CLK(clk), .RST(rst), .Q(o[478]) );
  DFF \oi_reg[14][29]  ( .D(N958), .CLK(clk), .RST(rst), .Q(o[477]) );
  DFF \oi_reg[14][28]  ( .D(N957), .CLK(clk), .RST(rst), .Q(o[476]) );
  DFF \oi_reg[14][27]  ( .D(N956), .CLK(clk), .RST(rst), .Q(o[475]) );
  DFF \oi_reg[14][26]  ( .D(N955), .CLK(clk), .RST(rst), .Q(o[474]) );
  DFF \oi_reg[14][25]  ( .D(N954), .CLK(clk), .RST(rst), .Q(o[473]) );
  DFF \oi_reg[14][24]  ( .D(N953), .CLK(clk), .RST(rst), .Q(o[472]) );
  DFF \oi_reg[14][23]  ( .D(N952), .CLK(clk), .RST(rst), .Q(o[471]) );
  DFF \oi_reg[14][22]  ( .D(N951), .CLK(clk), .RST(rst), .Q(o[470]) );
  DFF \oi_reg[14][21]  ( .D(N950), .CLK(clk), .RST(rst), .Q(o[469]) );
  DFF \oi_reg[14][20]  ( .D(N949), .CLK(clk), .RST(rst), .Q(o[468]) );
  DFF \oi_reg[14][19]  ( .D(N948), .CLK(clk), .RST(rst), .Q(o[467]) );
  DFF \oi_reg[14][18]  ( .D(N947), .CLK(clk), .RST(rst), .Q(o[466]) );
  DFF \oi_reg[14][17]  ( .D(N946), .CLK(clk), .RST(rst), .Q(o[465]) );
  DFF \oi_reg[14][16]  ( .D(N945), .CLK(clk), .RST(rst), .Q(o[464]) );
  DFF \oi_reg[14][15]  ( .D(N944), .CLK(clk), .RST(rst), .Q(o[463]) );
  DFF \oi_reg[14][14]  ( .D(N943), .CLK(clk), .RST(rst), .Q(o[462]) );
  DFF \oi_reg[14][13]  ( .D(N942), .CLK(clk), .RST(rst), .Q(o[461]) );
  DFF \oi_reg[14][12]  ( .D(N941), .CLK(clk), .RST(rst), .Q(o[460]) );
  DFF \oi_reg[14][11]  ( .D(N940), .CLK(clk), .RST(rst), .Q(o[459]) );
  DFF \oi_reg[14][10]  ( .D(N939), .CLK(clk), .RST(rst), .Q(o[458]) );
  DFF \oi_reg[14][9]  ( .D(N938), .CLK(clk), .RST(rst), .Q(o[457]) );
  DFF \oi_reg[14][8]  ( .D(N937), .CLK(clk), .RST(rst), .Q(o[456]) );
  DFF \oi_reg[14][7]  ( .D(N936), .CLK(clk), .RST(rst), .Q(o[455]) );
  DFF \oi_reg[14][6]  ( .D(N935), .CLK(clk), .RST(rst), .Q(o[454]) );
  DFF \oi_reg[14][5]  ( .D(N934), .CLK(clk), .RST(rst), .Q(o[453]) );
  DFF \oi_reg[14][4]  ( .D(N933), .CLK(clk), .RST(rst), .Q(o[452]) );
  DFF \oi_reg[14][3]  ( .D(N932), .CLK(clk), .RST(rst), .Q(o[451]) );
  DFF \oi_reg[14][2]  ( .D(N931), .CLK(clk), .RST(rst), .Q(o[450]) );
  DFF \oi_reg[14][1]  ( .D(N930), .CLK(clk), .RST(rst), .Q(o[449]) );
  DFF \oi_reg[14][0]  ( .D(N929), .CLK(clk), .RST(rst), .Q(o[448]) );
  DFF \oi_reg[15][31]  ( .D(N1024), .CLK(clk), .RST(rst), .Q(o[511]) );
  DFF \oi_reg[15][30]  ( .D(N1023), .CLK(clk), .RST(rst), .Q(o[510]) );
  DFF \oi_reg[15][29]  ( .D(N1022), .CLK(clk), .RST(rst), .Q(o[509]) );
  DFF \oi_reg[15][28]  ( .D(N1021), .CLK(clk), .RST(rst), .Q(o[508]) );
  DFF \oi_reg[15][27]  ( .D(N1020), .CLK(clk), .RST(rst), .Q(o[507]) );
  DFF \oi_reg[15][26]  ( .D(N1019), .CLK(clk), .RST(rst), .Q(o[506]) );
  DFF \oi_reg[15][25]  ( .D(N1018), .CLK(clk), .RST(rst), .Q(o[505]) );
  DFF \oi_reg[15][24]  ( .D(N1017), .CLK(clk), .RST(rst), .Q(o[504]) );
  DFF \oi_reg[15][23]  ( .D(N1016), .CLK(clk), .RST(rst), .Q(o[503]) );
  DFF \oi_reg[15][22]  ( .D(N1015), .CLK(clk), .RST(rst), .Q(o[502]) );
  DFF \oi_reg[15][21]  ( .D(N1014), .CLK(clk), .RST(rst), .Q(o[501]) );
  DFF \oi_reg[15][20]  ( .D(N1013), .CLK(clk), .RST(rst), .Q(o[500]) );
  DFF \oi_reg[15][19]  ( .D(N1012), .CLK(clk), .RST(rst), .Q(o[499]) );
  DFF \oi_reg[15][18]  ( .D(N1011), .CLK(clk), .RST(rst), .Q(o[498]) );
  DFF \oi_reg[15][17]  ( .D(N1010), .CLK(clk), .RST(rst), .Q(o[497]) );
  DFF \oi_reg[15][16]  ( .D(N1009), .CLK(clk), .RST(rst), .Q(o[496]) );
  DFF \oi_reg[15][15]  ( .D(N1008), .CLK(clk), .RST(rst), .Q(o[495]) );
  DFF \oi_reg[15][14]  ( .D(N1007), .CLK(clk), .RST(rst), .Q(o[494]) );
  DFF \oi_reg[15][13]  ( .D(N1006), .CLK(clk), .RST(rst), .Q(o[493]) );
  DFF \oi_reg[15][12]  ( .D(N1005), .CLK(clk), .RST(rst), .Q(o[492]) );
  DFF \oi_reg[15][11]  ( .D(N1004), .CLK(clk), .RST(rst), .Q(o[491]) );
  DFF \oi_reg[15][10]  ( .D(N1003), .CLK(clk), .RST(rst), .Q(o[490]) );
  DFF \oi_reg[15][9]  ( .D(N1002), .CLK(clk), .RST(rst), .Q(o[489]) );
  DFF \oi_reg[15][8]  ( .D(N1001), .CLK(clk), .RST(rst), .Q(o[488]) );
  DFF \oi_reg[15][7]  ( .D(N1000), .CLK(clk), .RST(rst), .Q(o[487]) );
  DFF \oi_reg[15][6]  ( .D(N999), .CLK(clk), .RST(rst), .Q(o[486]) );
  DFF \oi_reg[15][5]  ( .D(N998), .CLK(clk), .RST(rst), .Q(o[485]) );
  DFF \oi_reg[15][4]  ( .D(N997), .CLK(clk), .RST(rst), .Q(o[484]) );
  DFF \oi_reg[15][3]  ( .D(N996), .CLK(clk), .RST(rst), .Q(o[483]) );
  DFF \oi_reg[15][2]  ( .D(N995), .CLK(clk), .RST(rst), .Q(o[482]) );
  DFF \oi_reg[15][1]  ( .D(N994), .CLK(clk), .RST(rst), .Q(o[481]) );
  DFF \oi_reg[15][0]  ( .D(N993), .CLK(clk), .RST(rst), .Q(o[480]) );
  XNOR U3 ( .A(n15367), .B(n15366), .Z(n15370) );
  NAND U4 ( .A(n47191), .B(n47192), .Z(n1) );
  NAND U5 ( .A(n47189), .B(n47190), .Z(n2) );
  NAND U6 ( .A(n1), .B(n2), .Z(n47334) );
  XNOR U7 ( .A(n40660), .B(n40659), .Z(n40641) );
  XNOR U8 ( .A(n24102), .B(n24101), .Z(n24141) );
  NAND U9 ( .A(n37516), .B(n37515), .Z(n3) );
  NANDN U10 ( .A(n38296), .B(n37709), .Z(n4) );
  NAND U11 ( .A(n3), .B(n4), .Z(n37622) );
  XNOR U12 ( .A(n38467), .B(n38466), .Z(n38468) );
  NAND U13 ( .A(n31425), .B(n31426), .Z(n5) );
  NAND U14 ( .A(n31603), .B(n32685), .Z(n6) );
  NAND U15 ( .A(n5), .B(n6), .Z(n31471) );
  AND U16 ( .A(n31849), .B(n31564), .Z(n7) );
  AND U17 ( .A(n31563), .B(y[8011]), .Z(n8) );
  NAND U18 ( .A(x[488]), .B(n8), .Z(n9) );
  NANDN U19 ( .A(n7), .B(n9), .Z(n31628) );
  NAND U20 ( .A(n19884), .B(n19885), .Z(n10) );
  NAND U21 ( .A(n19997), .B(n21407), .Z(n11) );
  NAND U22 ( .A(n10), .B(n11), .Z(n19930) );
  NAND U23 ( .A(n21216), .B(n21215), .Z(n12) );
  NAND U24 ( .A(n21214), .B(n21213), .Z(n13) );
  AND U25 ( .A(n12), .B(n13), .Z(n21365) );
  AND U26 ( .A(n17669), .B(n17668), .Z(n14) );
  ANDN U27 ( .B(x[481]), .A(n19135), .Z(n15) );
  NAND U28 ( .A(y[7849]), .B(n15), .Z(n16) );
  NANDN U29 ( .A(n14), .B(n16), .Z(n17839) );
  NAND U30 ( .A(n17845), .B(n17844), .Z(n17) );
  NAND U31 ( .A(n17842), .B(n17843), .Z(n18) );
  NAND U32 ( .A(n17), .B(n18), .Z(n17885) );
  XNOR U33 ( .A(n15655), .B(n15654), .Z(n15687) );
  NAND U34 ( .A(n15549), .B(n15550), .Z(n19) );
  NANDN U35 ( .A(n15552), .B(n15551), .Z(n20) );
  AND U36 ( .A(n19), .B(n20), .Z(n15620) );
  XNOR U37 ( .A(n15693), .B(n15692), .Z(n15694) );
  XNOR U38 ( .A(n2445), .B(n3319), .Z(n2438) );
  XNOR U39 ( .A(n3179), .B(n3178), .Z(n3133) );
  NAND U40 ( .A(n47712), .B(n47711), .Z(n21) );
  NAND U41 ( .A(n47709), .B(n47710), .Z(n22) );
  NAND U42 ( .A(n21), .B(n22), .Z(n47984) );
  XNOR U43 ( .A(n44442), .B(n44441), .Z(n44443) );
  XNOR U44 ( .A(n44836), .B(n44835), .Z(n44912) );
  NAND U45 ( .A(n37620), .B(n37619), .Z(n23) );
  NAND U46 ( .A(n37618), .B(n37617), .Z(n24) );
  AND U47 ( .A(n23), .B(n24), .Z(n37751) );
  XNOR U48 ( .A(n37698), .B(n37697), .Z(n37764) );
  NAND U49 ( .A(n39058), .B(n39059), .Z(n25) );
  NAND U50 ( .A(n39056), .B(n39057), .Z(n26) );
  NAND U51 ( .A(n25), .B(n26), .Z(n39307) );
  NAND U52 ( .A(n38946), .B(n38947), .Z(n27) );
  NAND U53 ( .A(n38944), .B(n38945), .Z(n28) );
  NAND U54 ( .A(n27), .B(n28), .Z(n39066) );
  NAND U55 ( .A(n36254), .B(n36253), .Z(n29) );
  NAND U56 ( .A(n36252), .B(n36403), .Z(n30) );
  NAND U57 ( .A(n29), .B(n30), .Z(n36454) );
  NAND U58 ( .A(n36222), .B(n36223), .Z(n31) );
  NAND U59 ( .A(n36220), .B(n36221), .Z(n32) );
  NAND U60 ( .A(n31), .B(n32), .Z(n36470) );
  NAND U61 ( .A(n36111), .B(n36112), .Z(n33) );
  NAND U62 ( .A(n36109), .B(n36110), .Z(n34) );
  NAND U63 ( .A(n33), .B(n34), .Z(n36213) );
  XNOR U64 ( .A(n22883), .B(n22882), .Z(n22884) );
  XNOR U65 ( .A(n24549), .B(n24550), .Z(n24631) );
  NAND U66 ( .A(n24430), .B(n24429), .Z(n35) );
  NAND U67 ( .A(n24428), .B(n24579), .Z(n36) );
  AND U68 ( .A(n35), .B(n36), .Z(n24540) );
  NAND U69 ( .A(n21371), .B(n21372), .Z(n37) );
  NAND U70 ( .A(n21369), .B(n21370), .Z(n38) );
  NAND U71 ( .A(n37), .B(n38), .Z(n21558) );
  NAND U72 ( .A(n21656), .B(n21655), .Z(n39) );
  NAND U73 ( .A(n21654), .B(n21813), .Z(n40) );
  NAND U74 ( .A(n39), .B(n40), .Z(n21861) );
  NAND U75 ( .A(n21629), .B(n21630), .Z(n41) );
  NAND U76 ( .A(n21627), .B(n21628), .Z(n42) );
  NAND U77 ( .A(n41), .B(n42), .Z(n21880) );
  NAND U78 ( .A(n21528), .B(n21529), .Z(n43) );
  NANDN U79 ( .A(n21531), .B(n21530), .Z(n44) );
  NAND U80 ( .A(n43), .B(n44), .Z(n21684) );
  NAND U81 ( .A(n21486), .B(n21487), .Z(n45) );
  NAND U82 ( .A(n21484), .B(n21485), .Z(n46) );
  NAND U83 ( .A(n45), .B(n46), .Z(n21693) );
  XNOR U84 ( .A(n18402), .B(n18401), .Z(n18405) );
  XNOR U85 ( .A(n15314), .B(n15313), .Z(n15315) );
  XNOR U86 ( .A(n15571), .B(n15570), .Z(n15593) );
  XNOR U87 ( .A(n15874), .B(n15873), .Z(n15876) );
  NAND U88 ( .A(n15627), .B(n15626), .Z(n47) );
  NAND U89 ( .A(n15624), .B(n15625), .Z(n48) );
  NAND U90 ( .A(n47), .B(n48), .Z(n15869) );
  XNOR U91 ( .A(n10942), .B(n10941), .Z(n10943) );
  NAND U92 ( .A(n11337), .B(n11336), .Z(n49) );
  NANDN U93 ( .A(n11335), .B(n11334), .Z(n50) );
  NAND U94 ( .A(n49), .B(n50), .Z(n11463) );
  XNOR U95 ( .A(n11457), .B(n11456), .Z(n11448) );
  XNOR U96 ( .A(n5578), .B(n5577), .Z(n5579) );
  XNOR U97 ( .A(n5644), .B(n5643), .Z(n5605) );
  XNOR U98 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U99 ( .A(n47684), .B(n47683), .Z(n47685) );
  XNOR U100 ( .A(n44830), .B(n44829), .Z(n44878) );
  XNOR U101 ( .A(n39114), .B(n39113), .Z(n39115) );
  NAND U102 ( .A(n39347), .B(n39348), .Z(n39351) );
  XNOR U103 ( .A(n27632), .B(n27631), .Z(n27600) );
  XNOR U104 ( .A(n24597), .B(n24596), .Z(n24616) );
  XNOR U105 ( .A(n24656), .B(n24655), .Z(n24647) );
  NAND U106 ( .A(n21713), .B(n21714), .Z(n51) );
  NAND U107 ( .A(n21711), .B(n21712), .Z(n52) );
  NAND U108 ( .A(n51), .B(n52), .Z(n21835) );
  XNOR U109 ( .A(n18943), .B(n18942), .Z(n18944) );
  XNOR U110 ( .A(n15310), .B(n15309), .Z(n15189) );
  NAND U111 ( .A(n15920), .B(n15919), .Z(n53) );
  NAND U112 ( .A(n15918), .B(n15917), .Z(n54) );
  AND U113 ( .A(n53), .B(n54), .Z(n16162) );
  XNOR U114 ( .A(n16435), .B(n16434), .Z(n16431) );
  XOR U115 ( .A(n16224), .B(n16223), .Z(n16222) );
  XNOR U116 ( .A(n9243), .B(n9242), .Z(n9138) );
  NAND U117 ( .A(n39141), .B(n39142), .Z(n55) );
  NAND U118 ( .A(n39139), .B(n39140), .Z(n56) );
  NAND U119 ( .A(n55), .B(n56), .Z(n39266) );
  NAND U120 ( .A(n39519), .B(n39518), .Z(n57) );
  NAND U121 ( .A(n39516), .B(n39517), .Z(n58) );
  NAND U122 ( .A(n57), .B(n58), .Z(n39520) );
  XOR U123 ( .A(n36512), .B(n36511), .Z(n36510) );
  NAND U124 ( .A(n28085), .B(n28086), .Z(n59) );
  NAND U125 ( .A(n28679), .B(n28883), .Z(n60) );
  NAND U126 ( .A(n59), .B(n60), .Z(n28098) );
  XNOR U127 ( .A(n24844), .B(n24843), .Z(n24841) );
  NAND U128 ( .A(n21797), .B(n21796), .Z(n61) );
  NAND U129 ( .A(n21795), .B(n22012), .Z(n62) );
  AND U130 ( .A(n61), .B(n62), .Z(n21908) );
  NAND U131 ( .A(n16543), .B(n16544), .Z(n63) );
  NAND U132 ( .A(n17340), .B(n17140), .Z(n64) );
  NAND U133 ( .A(n63), .B(n64), .Z(n16556) );
  XNOR U134 ( .A(n17634), .B(n17633), .Z(n17526) );
  NAND U135 ( .A(n16009), .B(n16010), .Z(n65) );
  NAND U136 ( .A(n16007), .B(n16008), .Z(n66) );
  NAND U137 ( .A(n65), .B(n66), .Z(n16149) );
  NAND U138 ( .A(n12878), .B(n12879), .Z(n67) );
  NANDN U139 ( .A(n12881), .B(n12880), .Z(n68) );
  AND U140 ( .A(n67), .B(n68), .Z(n13034) );
  XOR U141 ( .A(n48005), .B(n48004), .Z(n48003) );
  NAND U142 ( .A(n44952), .B(n44951), .Z(n69) );
  NANDN U143 ( .A(n44950), .B(n44949), .Z(n70) );
  AND U144 ( .A(n69), .B(n70), .Z(n45110) );
  XNOR U145 ( .A(n39314), .B(n39313), .Z(n39311) );
  XNOR U146 ( .A(n36728), .B(n36727), .Z(n36725) );
  XNOR U147 ( .A(n30941), .B(n30940), .Z(n30684) );
  NAND U148 ( .A(n21737), .B(n21736), .Z(n71) );
  NAND U149 ( .A(n21734), .B(n21735), .Z(n72) );
  NAND U150 ( .A(n71), .B(n72), .Z(n22139) );
  XNOR U151 ( .A(n16481), .B(n16480), .Z(n16478) );
  OR U152 ( .A(n3221), .B(n3222), .Z(n73) );
  NAND U153 ( .A(n3220), .B(n3219), .Z(n74) );
  AND U154 ( .A(n73), .B(n74), .Z(n3462) );
  XNOR U155 ( .A(n4570), .B(n4571), .Z(n4569) );
  XNOR U156 ( .A(n40579), .B(o[434]), .Z(n40559) );
  XNOR U157 ( .A(n32465), .B(n32464), .Z(n32428) );
  XNOR U158 ( .A(n24094), .B(n24093), .Z(n24095) );
  XNOR U159 ( .A(n5863), .B(o[50]), .Z(n5843) );
  XNOR U160 ( .A(n40545), .B(n40544), .Z(n40588) );
  XNOR U161 ( .A(n40693), .B(n40692), .Z(n40642) );
  XNOR U162 ( .A(n40655), .B(n40654), .Z(n40701) );
  XNOR U163 ( .A(n38378), .B(n38377), .Z(n38315) );
  XNOR U164 ( .A(n35822), .B(n35821), .Z(n35823) );
  XNOR U165 ( .A(n32153), .B(o[340]), .Z(n32144) );
  XNOR U166 ( .A(n32353), .B(n32586), .Z(n32300) );
  XNOR U167 ( .A(n32304), .B(n32303), .Z(n32315) );
  XNOR U168 ( .A(n26945), .B(n26944), .Z(n26950) );
  XNOR U169 ( .A(n23753), .B(n23752), .Z(n23790) );
  XOR U170 ( .A(n24120), .B(n24119), .Z(n24147) );
  XNOR U171 ( .A(n24064), .B(n24063), .Z(n24069) );
  XNOR U172 ( .A(n20149), .B(o[208]), .Z(n20163) );
  XNOR U173 ( .A(n20241), .B(n20240), .Z(n20255) );
  XNOR U174 ( .A(n20425), .B(o[211]), .Z(n20449) );
  XNOR U175 ( .A(n20659), .B(n20658), .Z(n20669) );
  XNOR U176 ( .A(n20678), .B(n20677), .Z(n20715) );
  XNOR U177 ( .A(n17473), .B(o[178]), .Z(n17453) );
  XNOR U178 ( .A(n17438), .B(n17437), .Z(n17482) );
  XNOR U179 ( .A(n18015), .B(n18014), .Z(n18052) );
  NAND U180 ( .A(n12529), .B(n12530), .Z(n75) );
  NAND U181 ( .A(n12527), .B(n12528), .Z(n76) );
  NAND U182 ( .A(n75), .B(n76), .Z(n12697) );
  XNOR U183 ( .A(n9727), .B(n9726), .Z(n9737) );
  XNOR U184 ( .A(n5948), .B(n5947), .Z(n5929) );
  XNOR U185 ( .A(n5943), .B(n5942), .Z(n5988) );
  NAND U186 ( .A(n47188), .B(n47187), .Z(n77) );
  NAND U187 ( .A(n47185), .B(n47186), .Z(n78) );
  NAND U188 ( .A(n77), .B(n78), .Z(n47336) );
  NAND U189 ( .A(n47146), .B(n47147), .Z(n79) );
  NANDN U190 ( .A(n47149), .B(n47148), .Z(n80) );
  NAND U191 ( .A(n79), .B(n80), .Z(n47280) );
  NAND U192 ( .A(n47345), .B(n47344), .Z(n81) );
  NAND U193 ( .A(n47342), .B(n47343), .Z(n82) );
  NAND U194 ( .A(n81), .B(n82), .Z(n47503) );
  XNOR U195 ( .A(n40836), .B(n40835), .Z(n40790) );
  XNOR U196 ( .A(n41366), .B(n41365), .Z(n41351) );
  NAND U197 ( .A(n41396), .B(n41397), .Z(n83) );
  NAND U198 ( .A(n41394), .B(n41395), .Z(n84) );
  NAND U199 ( .A(n83), .B(n84), .Z(n41469) );
  NAND U200 ( .A(n37514), .B(n37513), .Z(n85) );
  NANDN U201 ( .A(n37640), .B(n37512), .Z(n86) );
  NAND U202 ( .A(n85), .B(n86), .Z(n37621) );
  XNOR U203 ( .A(n36019), .B(n36018), .Z(n36020) );
  XNOR U204 ( .A(n31355), .B(n31354), .Z(n31318) );
  NAND U205 ( .A(n31476), .B(n32348), .Z(n87) );
  NAND U206 ( .A(n31475), .B(n31627), .Z(n88) );
  NAND U207 ( .A(n87), .B(n88), .Z(n31574) );
  NAND U208 ( .A(n31498), .B(n31499), .Z(n89) );
  NAND U209 ( .A(n31603), .B(n33069), .Z(n90) );
  NAND U210 ( .A(n89), .B(n90), .Z(n31535) );
  XNOR U211 ( .A(n32399), .B(n32398), .Z(n32474) );
  XOR U212 ( .A(n32411), .B(n32410), .Z(n32480) );
  XNOR U213 ( .A(n32669), .B(n32668), .Z(n32670) );
  NAND U214 ( .A(n26094), .B(n26095), .Z(n91) );
  NAND U215 ( .A(n26092), .B(n26093), .Z(n92) );
  NAND U216 ( .A(n91), .B(n92), .Z(n26203) );
  XNOR U217 ( .A(n22851), .B(n22850), .Z(n22852) );
  XNOR U218 ( .A(n24142), .B(n24141), .Z(n24143) );
  XNOR U219 ( .A(n24204), .B(n24203), .Z(n24205) );
  XNOR U220 ( .A(n24302), .B(n24301), .Z(n24303) );
  NAND U221 ( .A(n19862), .B(n20703), .Z(n93) );
  NAND U222 ( .A(n19861), .B(n20021), .Z(n94) );
  NAND U223 ( .A(n93), .B(n94), .Z(n19972) );
  NAND U224 ( .A(n19956), .B(n19957), .Z(n95) );
  NAND U225 ( .A(n19997), .B(n21647), .Z(n96) );
  NAND U226 ( .A(n95), .B(n96), .Z(n20023) );
  XNOR U227 ( .A(n20208), .B(o[209]), .Z(n20213) );
  XNOR U228 ( .A(n20541), .B(n20540), .Z(n20594) );
  XNOR U229 ( .A(n20411), .B(n20410), .Z(n20392) );
  XNOR U230 ( .A(n20420), .B(n20419), .Z(n20459) );
  XNOR U231 ( .A(n20603), .B(n20602), .Z(n20553) );
  XNOR U232 ( .A(n20772), .B(n20771), .Z(n20773) );
  NAND U233 ( .A(n21381), .B(n21380), .Z(n97) );
  NAND U234 ( .A(n21378), .B(n21379), .Z(n98) );
  NAND U235 ( .A(n97), .B(n98), .Z(n21477) );
  XNOR U236 ( .A(n16829), .B(n16828), .Z(n16847) );
  OR U237 ( .A(n17381), .B(n18294), .Z(n99) );
  NAND U238 ( .A(n17382), .B(n17383), .Z(n100) );
  AND U239 ( .A(n99), .B(n100), .Z(n17479) );
  XNOR U240 ( .A(n15135), .B(n15134), .Z(n15093) );
  OR U241 ( .A(n15489), .B(n15490), .Z(n101) );
  NAND U242 ( .A(n15488), .B(n15487), .Z(n102) );
  AND U243 ( .A(n101), .B(n102), .Z(n15664) );
  XNOR U244 ( .A(n15615), .B(n15614), .Z(n15616) );
  XNOR U245 ( .A(n15701), .B(n15700), .Z(n15695) );
  XNOR U246 ( .A(n11532), .B(n12246), .Z(n11494) );
  XNOR U247 ( .A(n11619), .B(n11618), .Z(n11624) );
  XNOR U248 ( .A(n11691), .B(n11690), .Z(n11692) );
  NAND U249 ( .A(n12486), .B(n12487), .Z(n103) );
  NANDN U250 ( .A(n12489), .B(n12488), .Z(n104) );
  NAND U251 ( .A(n103), .B(n104), .Z(n12644) );
  NAND U252 ( .A(n12708), .B(n12707), .Z(n105) );
  NANDN U253 ( .A(n12706), .B(n12705), .Z(n106) );
  NAND U254 ( .A(n105), .B(n106), .Z(n12865) );
  XNOR U255 ( .A(n8202), .B(n8201), .Z(n8165) );
  XNOR U256 ( .A(n5654), .B(n6366), .Z(n5617) );
  XNOR U257 ( .A(n5741), .B(n5740), .Z(n5746) );
  XNOR U258 ( .A(n5813), .B(n5812), .Z(n5814) );
  XNOR U259 ( .A(n5956), .B(n5955), .Z(n5994) );
  XNOR U260 ( .A(n6129), .B(n6128), .Z(n6079) );
  XNOR U261 ( .A(n3042), .B(n3159), .Z(n3013) );
  XNOR U262 ( .A(n3185), .B(n3184), .Z(n3135) );
  XNOR U263 ( .A(n46297), .B(n46296), .Z(n46319) );
  NAND U264 ( .A(n47707), .B(n47708), .Z(n107) );
  NAND U265 ( .A(n47705), .B(n47706), .Z(n108) );
  NAND U266 ( .A(n107), .B(n108), .Z(n47983) );
  XNOR U267 ( .A(n44444), .B(n44443), .Z(n44435) );
  XNOR U268 ( .A(n44859), .B(n44858), .Z(n44860) );
  XNOR U269 ( .A(n44867), .B(n44866), .Z(n44913) );
  XNOR U270 ( .A(n44843), .B(n44842), .Z(n44918) );
  NAND U271 ( .A(n44664), .B(n44663), .Z(n109) );
  NANDN U272 ( .A(n44662), .B(n44661), .Z(n110) );
  NAND U273 ( .A(n109), .B(n110), .Z(n44906) );
  XNOR U274 ( .A(n44788), .B(n44787), .Z(n44790) );
  XOR U275 ( .A(n40728), .B(n40727), .Z(n40732) );
  XOR U276 ( .A(n40848), .B(n40847), .Z(n40852) );
  XNOR U277 ( .A(n41022), .B(n41021), .Z(n41023) );
  XOR U278 ( .A(n42168), .B(n42167), .Z(n42170) );
  NAND U279 ( .A(n37616), .B(n37615), .Z(n111) );
  NAND U280 ( .A(n37614), .B(n37613), .Z(n112) );
  AND U281 ( .A(n111), .B(n112), .Z(n37752) );
  XOR U282 ( .A(n38568), .B(n38567), .Z(n38561) );
  NAND U283 ( .A(n39083), .B(n39082), .Z(n113) );
  NAND U284 ( .A(n39241), .B(n39081), .Z(n114) );
  AND U285 ( .A(n113), .B(n114), .Z(n39290) );
  NAND U286 ( .A(n39054), .B(n39055), .Z(n115) );
  NAND U287 ( .A(n39052), .B(n39053), .Z(n116) );
  NAND U288 ( .A(n115), .B(n116), .Z(n39306) );
  NAND U289 ( .A(n38943), .B(n38942), .Z(n117) );
  NAND U290 ( .A(n38940), .B(n38941), .Z(n118) );
  NAND U291 ( .A(n117), .B(n118), .Z(n39065) );
  NAND U292 ( .A(n35999), .B(n35998), .Z(n119) );
  NAND U293 ( .A(n35996), .B(n35997), .Z(n120) );
  NAND U294 ( .A(n119), .B(n120), .Z(n36152) );
  NAND U295 ( .A(n35973), .B(n35974), .Z(n121) );
  NAND U296 ( .A(n35971), .B(n35972), .Z(n122) );
  NAND U297 ( .A(n121), .B(n122), .Z(n36149) );
  NAND U298 ( .A(n36132), .B(n36131), .Z(n123) );
  NAND U299 ( .A(n36129), .B(n36130), .Z(n124) );
  NAND U300 ( .A(n123), .B(n124), .Z(n36305) );
  NAND U301 ( .A(n36146), .B(n36147), .Z(n125) );
  NAND U302 ( .A(n36144), .B(n36145), .Z(n126) );
  NAND U303 ( .A(n125), .B(n126), .Z(n36300) );
  NAND U304 ( .A(n36218), .B(n36219), .Z(n127) );
  NAND U305 ( .A(n36216), .B(n36217), .Z(n128) );
  NAND U306 ( .A(n127), .B(n128), .Z(n36469) );
  NAND U307 ( .A(n36107), .B(n36108), .Z(n129) );
  NAND U308 ( .A(n36105), .B(n36106), .Z(n130) );
  NAND U309 ( .A(n129), .B(n130), .Z(n36212) );
  XNOR U310 ( .A(n36294), .B(n36293), .Z(n36296) );
  NAND U311 ( .A(n31573), .B(n31572), .Z(n131) );
  NAND U312 ( .A(n31956), .B(n31571), .Z(n132) );
  AND U313 ( .A(n131), .B(n132), .Z(n31670) );
  XNOR U314 ( .A(n31667), .B(n31666), .Z(n31659) );
  XNOR U315 ( .A(n28523), .B(n28522), .Z(n28510) );
  XNOR U316 ( .A(n30412), .B(n30611), .Z(n30413) );
  XNOR U317 ( .A(n25837), .B(n25836), .Z(n25878) );
  NAND U318 ( .A(n25987), .B(n25986), .Z(n133) );
  NANDN U319 ( .A(n26937), .B(n26060), .Z(n134) );
  NAND U320 ( .A(n133), .B(n134), .Z(n26108) );
  NAND U321 ( .A(n26215), .B(n26214), .Z(n135) );
  NAND U322 ( .A(n26213), .B(n26212), .Z(n136) );
  AND U323 ( .A(n135), .B(n136), .Z(n26349) );
  XNOR U324 ( .A(n22917), .B(n22916), .Z(n22958) );
  XOR U325 ( .A(n24467), .B(n24466), .Z(n24484) );
  XNOR U326 ( .A(n24546), .B(n24545), .Z(n24630) );
  NAND U327 ( .A(n19971), .B(n19970), .Z(n137) );
  NAND U328 ( .A(n20346), .B(n19969), .Z(n138) );
  AND U329 ( .A(n137), .B(n138), .Z(n20064) );
  XNOR U330 ( .A(n20061), .B(n20060), .Z(n20053) );
  NAND U331 ( .A(n20012), .B(n20011), .Z(n139) );
  NAND U332 ( .A(n20152), .B(n20010), .Z(n140) );
  NAND U333 ( .A(n139), .B(n140), .Z(n20132) );
  XNOR U334 ( .A(n20456), .B(n20455), .Z(n20474) );
  XNOR U335 ( .A(n20520), .B(n20519), .Z(n20606) );
  XNOR U336 ( .A(n20870), .B(n20869), .Z(n20874) );
  NAND U337 ( .A(n21367), .B(n21368), .Z(n141) );
  NAND U338 ( .A(n21365), .B(n21366), .Z(n142) );
  NAND U339 ( .A(n141), .B(n142), .Z(n21559) );
  NAND U340 ( .A(n21540), .B(n21541), .Z(n143) );
  NAND U341 ( .A(n21538), .B(n21539), .Z(n144) );
  NAND U342 ( .A(n143), .B(n144), .Z(n21703) );
  NAND U343 ( .A(n21625), .B(n21626), .Z(n145) );
  NAND U344 ( .A(n21623), .B(n21624), .Z(n146) );
  NAND U345 ( .A(n145), .B(n146), .Z(n21879) );
  NAND U346 ( .A(n21510), .B(n21511), .Z(n147) );
  NAND U347 ( .A(n21508), .B(n21509), .Z(n148) );
  NAND U348 ( .A(n147), .B(n148), .Z(n21636) );
  NAND U349 ( .A(n21526), .B(n21527), .Z(n149) );
  NAND U350 ( .A(n21524), .B(n21525), .Z(n150) );
  NAND U351 ( .A(n149), .B(n150), .Z(n21683) );
  NAND U352 ( .A(n21480), .B(n21481), .Z(n151) );
  NANDN U353 ( .A(n21483), .B(n21482), .Z(n152) );
  NAND U354 ( .A(n151), .B(n152), .Z(n21695) );
  XNOR U355 ( .A(n17209), .B(n17208), .Z(n17200) );
  NAND U356 ( .A(n17290), .B(n17291), .Z(n153) );
  NAND U357 ( .A(n17288), .B(n17289), .Z(n154) );
  NAND U358 ( .A(n153), .B(n154), .Z(n17396) );
  NAND U359 ( .A(n17841), .B(n17840), .Z(n155) );
  NAND U360 ( .A(n17838), .B(n17839), .Z(n156) );
  NAND U361 ( .A(n155), .B(n156), .Z(n17887) );
  XNOR U362 ( .A(n15308), .B(n15307), .Z(n15309) );
  XNOR U363 ( .A(n15522), .B(n15521), .Z(n15483) );
  NAND U364 ( .A(n15671), .B(n15670), .Z(n157) );
  NAND U365 ( .A(n15668), .B(n15669), .Z(n158) );
  NAND U366 ( .A(n157), .B(n158), .Z(n15866) );
  XNOR U367 ( .A(n15888), .B(n15887), .Z(n15759) );
  NAND U368 ( .A(n15817), .B(n15818), .Z(n159) );
  NAND U369 ( .A(n15815), .B(n15816), .Z(n160) );
  NAND U370 ( .A(n159), .B(n160), .Z(n15918) );
  NAND U371 ( .A(n15943), .B(n15944), .Z(n161) );
  NAND U372 ( .A(n15945), .B(n15946), .Z(n162) );
  NAND U373 ( .A(n161), .B(n162), .Z(n16177) );
  NAND U374 ( .A(n15927), .B(n15928), .Z(n163) );
  NAND U375 ( .A(n15925), .B(n15926), .Z(n164) );
  NAND U376 ( .A(n163), .B(n164), .Z(n16181) );
  XNOR U377 ( .A(n11522), .B(n11521), .Z(n11482) );
  NAND U378 ( .A(n10026), .B(n10027), .Z(n165) );
  NAND U379 ( .A(n10024), .B(n10025), .Z(n166) );
  NAND U380 ( .A(n165), .B(n166), .Z(n10226) );
  XOR U381 ( .A(n10436), .B(n10435), .Z(n10437) );
  XNOR U382 ( .A(n7251), .B(n7250), .Z(n7281) );
  XOR U383 ( .A(n7490), .B(n7489), .Z(n7492) );
  XNOR U384 ( .A(n2484), .B(n2483), .Z(n2432) );
  XNOR U385 ( .A(n3257), .B(n3256), .Z(n3258) );
  XNOR U386 ( .A(n4201), .B(n4200), .Z(n4202) );
  XNOR U387 ( .A(n4158), .B(n4157), .Z(n4095) );
  XNOR U388 ( .A(n47974), .B(n47973), .Z(n47952) );
  NAND U389 ( .A(n47934), .B(n47933), .Z(n167) );
  NANDN U390 ( .A(n48159), .B(n47932), .Z(n168) );
  NAND U391 ( .A(n167), .B(n168), .Z(n48049) );
  NAND U392 ( .A(n43292), .B(n43293), .Z(n169) );
  NANDN U393 ( .A(n43295), .B(n43294), .Z(n170) );
  NAND U394 ( .A(n169), .B(n170), .Z(n43307) );
  XNOR U395 ( .A(n44881), .B(n44880), .Z(n44902) );
  NAND U396 ( .A(n37766), .B(n37765), .Z(n171) );
  NAND U397 ( .A(n37763), .B(n37764), .Z(n172) );
  NAND U398 ( .A(n171), .B(n172), .Z(n37873) );
  XOR U399 ( .A(n39033), .B(n39032), .Z(n39019) );
  NAND U400 ( .A(n39099), .B(n39100), .Z(n173) );
  NAND U401 ( .A(n39097), .B(n39098), .Z(n174) );
  NAND U402 ( .A(n173), .B(n174), .Z(n39219) );
  NAND U403 ( .A(n38978), .B(n38979), .Z(n175) );
  NAND U404 ( .A(n38976), .B(n38977), .Z(n176) );
  NAND U405 ( .A(n175), .B(n176), .Z(n39132) );
  NAND U406 ( .A(n39283), .B(n39284), .Z(n177) );
  NANDN U407 ( .A(n39286), .B(n39285), .Z(n178) );
  AND U408 ( .A(n177), .B(n178), .Z(n39518) );
  NAND U409 ( .A(n39051), .B(n39050), .Z(n179) );
  NAND U410 ( .A(n39049), .B(n39048), .Z(n180) );
  AND U411 ( .A(n179), .B(n180), .Z(n39274) );
  NAND U412 ( .A(n36309), .B(n36310), .Z(n181) );
  NAND U413 ( .A(n36307), .B(n36308), .Z(n182) );
  NAND U414 ( .A(n181), .B(n182), .Z(n36440) );
  XNOR U415 ( .A(n36466), .B(n36465), .Z(n36436) );
  NAND U416 ( .A(n36232), .B(n36231), .Z(n183) );
  NAND U417 ( .A(n36230), .B(n36229), .Z(n184) );
  AND U418 ( .A(n183), .B(n184), .Z(n36447) );
  XNOR U419 ( .A(n33566), .B(n33565), .Z(n33567) );
  XOR U420 ( .A(n33758), .B(n33595), .Z(n185) );
  NAND U421 ( .A(n185), .B(n33596), .Z(n186) );
  NAND U422 ( .A(n33758), .B(n33595), .Z(n187) );
  AND U423 ( .A(n186), .B(n187), .Z(n33845) );
  XNOR U424 ( .A(n30420), .B(n30419), .Z(n30480) );
  XNOR U425 ( .A(n30397), .B(n30396), .Z(n30486) );
  XNOR U426 ( .A(n30632), .B(n30631), .Z(n30633) );
  XNOR U427 ( .A(n27594), .B(n27593), .Z(n27595) );
  XOR U428 ( .A(n27600), .B(n27599), .Z(n27602) );
  XNOR U429 ( .A(n22891), .B(n22890), .Z(n22871) );
  XNOR U430 ( .A(n24490), .B(n24489), .Z(n24492) );
  XNOR U431 ( .A(n24540), .B(n24539), .Z(n24618) );
  NAND U432 ( .A(n24626), .B(n24627), .Z(n188) );
  NANDN U433 ( .A(n24629), .B(n24628), .Z(n189) );
  AND U434 ( .A(n188), .B(n189), .Z(n24757) );
  XNOR U435 ( .A(n19783), .B(n19782), .Z(n19784) );
  XNOR U436 ( .A(n20370), .B(n20369), .Z(n20295) );
  XNOR U437 ( .A(n20492), .B(n20491), .Z(n20495) );
  XNOR U438 ( .A(n21031), .B(n21030), .Z(n21032) );
  XNOR U439 ( .A(n21580), .B(n21579), .Z(n21465) );
  NAND U440 ( .A(n21709), .B(n21710), .Z(n190) );
  NAND U441 ( .A(n21707), .B(n21708), .Z(n191) );
  NAND U442 ( .A(n190), .B(n191), .Z(n21834) );
  XNOR U443 ( .A(n21855), .B(n21854), .Z(n21831) );
  NAND U444 ( .A(n21622), .B(n21621), .Z(n192) );
  NAND U445 ( .A(n21620), .B(n21619), .Z(n193) );
  AND U446 ( .A(n192), .B(n193), .Z(n21843) );
  XNOR U447 ( .A(n21594), .B(n21593), .Z(n21595) );
  NAND U448 ( .A(n17402), .B(n17403), .Z(n194) );
  NAND U449 ( .A(n17400), .B(n17401), .Z(n195) );
  NAND U450 ( .A(n194), .B(n195), .Z(n17415) );
  XNOR U451 ( .A(n18423), .B(n18422), .Z(n18424) );
  XOR U452 ( .A(n18949), .B(n18948), .Z(n18951) );
  NAND U453 ( .A(n14390), .B(n14389), .Z(n196) );
  NANDN U454 ( .A(n14388), .B(n14387), .Z(n197) );
  AND U455 ( .A(n196), .B(n197), .Z(n14393) );
  XNOR U456 ( .A(n15304), .B(n15303), .Z(n15191) );
  XNOR U457 ( .A(n15609), .B(n15608), .Z(n15610) );
  XNOR U458 ( .A(n15902), .B(n15901), .Z(n15903) );
  OR U459 ( .A(n15969), .B(n15970), .Z(n198) );
  NAND U460 ( .A(n15972), .B(n15971), .Z(n199) );
  NAND U461 ( .A(n198), .B(n199), .Z(n16081) );
  NAND U462 ( .A(n16141), .B(n16140), .Z(n200) );
  NAND U463 ( .A(n16139), .B(n16249), .Z(n201) );
  AND U464 ( .A(n200), .B(n201), .Z(n16221) );
  XNOR U465 ( .A(n10944), .B(n10943), .Z(n10957) );
  XNOR U466 ( .A(n11477), .B(n11476), .Z(n11478) );
  XNOR U467 ( .A(n13313), .B(n13312), .Z(n13233) );
  XNOR U468 ( .A(n9138), .B(n9137), .Z(n9139) );
  XNOR U469 ( .A(n10432), .B(n10431), .Z(n10408) );
  XNOR U470 ( .A(n10669), .B(n10668), .Z(n10666) );
  XNOR U471 ( .A(n10444), .B(n10443), .Z(n10418) );
  XNOR U472 ( .A(n5273), .B(n5272), .Z(n5274) );
  XNOR U473 ( .A(n5638), .B(n5637), .Z(n5607) );
  XNOR U474 ( .A(n5586), .B(n5585), .Z(n5566) );
  XNOR U475 ( .A(n7234), .B(n7233), .Z(n7323) );
  XNOR U476 ( .A(n7486), .B(n7485), .Z(n7377) );
  XNOR U477 ( .A(n7381), .B(n7380), .Z(n7382) );
  XNOR U478 ( .A(n2501), .B(n2500), .Z(n2502) );
  XNOR U479 ( .A(n4355), .B(n4354), .Z(n4249) );
  XNOR U480 ( .A(n47686), .B(n47685), .Z(n47678) );
  XNOR U481 ( .A(n48015), .B(n48014), .Z(n48231) );
  NAND U482 ( .A(n43313), .B(n43312), .Z(n202) );
  NANDN U483 ( .A(n43311), .B(n43310), .Z(n203) );
  AND U484 ( .A(n202), .B(n203), .Z(n43406) );
  XOR U485 ( .A(n45330), .B(n45329), .Z(n45328) );
  NAND U486 ( .A(n41719), .B(n41720), .Z(n204) );
  NAND U487 ( .A(n41717), .B(n41718), .Z(n205) );
  NAND U488 ( .A(n204), .B(n205), .Z(n41872) );
  XOR U489 ( .A(n42384), .B(n42385), .Z(n42233) );
  NAND U490 ( .A(n39137), .B(n39138), .Z(n206) );
  NAND U491 ( .A(n39135), .B(n39136), .Z(n207) );
  NAND U492 ( .A(n206), .B(n207), .Z(n39265) );
  NAND U493 ( .A(n39336), .B(n39335), .Z(n208) );
  NANDN U494 ( .A(n39338), .B(n39337), .Z(n209) );
  AND U495 ( .A(n208), .B(n209), .Z(n210) );
  NANDN U496 ( .A(n39342), .B(n39341), .Z(n211) );
  NANDN U497 ( .A(n39340), .B(n39339), .Z(n212) );
  AND U498 ( .A(n211), .B(n212), .Z(n213) );
  NAND U499 ( .A(n39344), .B(n39343), .Z(n214) );
  NAND U500 ( .A(n39345), .B(n39346), .Z(n215) );
  AND U501 ( .A(n214), .B(n215), .Z(n216) );
  XOR U502 ( .A(n39507), .B(n39506), .Z(n217) );
  XNOR U503 ( .A(n39477), .B(n39476), .Z(n218) );
  XNOR U504 ( .A(n217), .B(n218), .Z(n219) );
  AND U505 ( .A(n39351), .B(n39350), .Z(n220) );
  XNOR U506 ( .A(n39422), .B(n39421), .Z(n221) );
  XNOR U507 ( .A(n220), .B(n221), .Z(n222) );
  XOR U508 ( .A(n219), .B(n222), .Z(n223) );
  XNOR U509 ( .A(n213), .B(n216), .Z(n224) );
  XNOR U510 ( .A(n223), .B(n224), .Z(n225) );
  XNOR U511 ( .A(n210), .B(n225), .Z(n39508) );
  NAND U512 ( .A(n36677), .B(n36678), .Z(n36682) );
  XNOR U513 ( .A(n31182), .B(n31181), .Z(n31195) );
  XNOR U514 ( .A(n25654), .B(n25653), .Z(n25728) );
  XNOR U515 ( .A(n22911), .B(n22910), .Z(n22996) );
  XNOR U516 ( .A(n24648), .B(n24647), .Z(n24649) );
  XOR U517 ( .A(n25036), .B(n25035), .Z(n25034) );
  XOR U518 ( .A(n19838), .B(n19837), .Z(n19842) );
  XNOR U519 ( .A(n20762), .B(n20761), .Z(n20879) );
  NAND U520 ( .A(n22091), .B(n22092), .Z(n22096) );
  NAND U521 ( .A(n17421), .B(n17420), .Z(n226) );
  NANDN U522 ( .A(n17419), .B(n17418), .Z(n227) );
  AND U523 ( .A(n226), .B(n227), .Z(n17527) );
  NAND U524 ( .A(n16005), .B(n16006), .Z(n228) );
  NAND U525 ( .A(n16003), .B(n16004), .Z(n229) );
  NAND U526 ( .A(n228), .B(n229), .Z(n16148) );
  XNOR U527 ( .A(n16453), .B(n16452), .Z(n16450) );
  NAND U528 ( .A(n16115), .B(n16116), .Z(n230) );
  NAND U529 ( .A(n16113), .B(n16114), .Z(n231) );
  NAND U530 ( .A(n230), .B(n231), .Z(n16440) );
  NAND U531 ( .A(n11388), .B(n11389), .Z(n232) );
  XOR U532 ( .A(n11388), .B(n11389), .Z(n233) );
  NANDN U533 ( .A(n11387), .B(n233), .Z(n234) );
  NAND U534 ( .A(n232), .B(n234), .Z(n11565) );
  XNOR U535 ( .A(n13043), .B(n13042), .Z(n13035) );
  XNOR U536 ( .A(n13394), .B(n13393), .Z(n13391) );
  XNOR U537 ( .A(n8022), .B(n8021), .Z(n8035) );
  XNOR U538 ( .A(n8082), .B(n8081), .Z(n8084) );
  XNOR U539 ( .A(n9386), .B(n9385), .Z(n9514) );
  XOR U540 ( .A(n5332), .B(n5331), .Z(n5336) );
  XNOR U541 ( .A(n5602), .B(n5601), .Z(n5688) );
  XOR U542 ( .A(n7783), .B(n7782), .Z(n7781) );
  NAND U543 ( .A(n3201), .B(n3202), .Z(n235) );
  NANDN U544 ( .A(n3204), .B(n3203), .Z(n236) );
  AND U545 ( .A(n235), .B(n236), .Z(n3219) );
  XNOR U546 ( .A(n3474), .B(n3473), .Z(n3602) );
  XNOR U547 ( .A(n4439), .B(n4438), .Z(n4440) );
  XNOR U548 ( .A(n48263), .B(n48262), .Z(n48276) );
  XOR U549 ( .A(n42898), .B(n42897), .Z(n237) );
  NANDN U550 ( .A(n42896), .B(n237), .Z(n238) );
  NAND U551 ( .A(n42898), .B(n42897), .Z(n239) );
  AND U552 ( .A(n238), .B(n239), .Z(n43035) );
  XNOR U553 ( .A(n45111), .B(n45110), .Z(n45109) );
  XNOR U554 ( .A(n36837), .B(n36836), .Z(n36833) );
  XOR U555 ( .A(n39581), .B(n39582), .Z(n39580) );
  NAND U556 ( .A(n36334), .B(n36335), .Z(n240) );
  NANDN U557 ( .A(n36337), .B(n36336), .Z(n241) );
  AND U558 ( .A(n240), .B(n241), .Z(n36726) );
  XOR U559 ( .A(n33622), .B(n33621), .Z(n33620) );
  NAND U560 ( .A(n28100), .B(n28099), .Z(n242) );
  NAND U561 ( .A(n28098), .B(n28097), .Z(n243) );
  AND U562 ( .A(n242), .B(n243), .Z(n28152) );
  NAND U563 ( .A(n29086), .B(n29087), .Z(n244) );
  NANDN U564 ( .A(n29089), .B(n29088), .Z(n245) );
  NAND U565 ( .A(n244), .B(n245), .Z(n29311) );
  XNOR U566 ( .A(n30685), .B(n30684), .Z(n30682) );
  XNOR U567 ( .A(n19456), .B(n19455), .Z(n19461) );
  XNOR U568 ( .A(n20755), .B(n20754), .Z(n20751) );
  XOR U569 ( .A(n22142), .B(n22141), .Z(n22140) );
  NAND U570 ( .A(n16558), .B(n16557), .Z(n246) );
  NAND U571 ( .A(n16556), .B(n16555), .Z(n247) );
  AND U572 ( .A(n246), .B(n247), .Z(n16610) );
  XNOR U573 ( .A(n17647), .B(n17646), .Z(n17652) );
  NANDN U574 ( .A(n19359), .B(n19358), .Z(n19363) );
  XNOR U575 ( .A(n13740), .B(n13739), .Z(n13745) );
  NAND U576 ( .A(n16051), .B(n16050), .Z(n248) );
  NAND U577 ( .A(n16049), .B(n16048), .Z(n249) );
  AND U578 ( .A(n248), .B(n249), .Z(n16479) );
  NAND U579 ( .A(n10307), .B(n10306), .Z(n250) );
  NANDN U580 ( .A(n10305), .B(n10304), .Z(n251) );
  AND U581 ( .A(n250), .B(n251), .Z(n10464) );
  XNOR U582 ( .A(n3467), .B(n3466), .Z(n3463) );
  XNOR U583 ( .A(n4831), .B(n4830), .Z(n4850) );
  XNOR U584 ( .A(n11720), .B(n11719), .Z(n11722) );
  XNOR U585 ( .A(n44044), .B(n44043), .Z(n44081) );
  XNOR U586 ( .A(n44340), .B(n44339), .Z(n44345) );
  XNOR U587 ( .A(n40566), .B(n40565), .Z(n40583) );
  XNOR U588 ( .A(n40554), .B(n40553), .Z(n40589) );
  XNOR U589 ( .A(n40702), .B(n40701), .Z(n40703) );
  XNOR U590 ( .A(n41158), .B(n41157), .Z(n41195) );
  XNOR U591 ( .A(n38360), .B(n38359), .Z(n38317) );
  XNOR U592 ( .A(n38366), .B(n38365), .Z(n38371) );
  XNOR U593 ( .A(n35824), .B(n35823), .Z(n35833) );
  XNOR U594 ( .A(n35792), .B(n35791), .Z(n35797) );
  XNOR U595 ( .A(n35860), .B(n35859), .Z(n35876) );
  AND U596 ( .A(n31345), .B(o[331]), .Z(n31424) );
  XNOR U597 ( .A(n32317), .B(n32316), .Z(n32282) );
  XNOR U598 ( .A(n32350), .B(n32349), .Z(n32285) );
  XNOR U599 ( .A(n29920), .B(n29919), .Z(n29925) );
  XNOR U600 ( .A(n26949), .B(n26948), .Z(n26951) );
  XNOR U601 ( .A(n23746), .B(n23745), .Z(n23792) );
  XNOR U602 ( .A(n23742), .B(o[247]), .Z(n23764) );
  XNOR U603 ( .A(n24096), .B(n24095), .Z(n24106) );
  XNOR U604 ( .A(n24125), .B(n24124), .Z(n24126) );
  AND U605 ( .A(n19743), .B(o[203]), .Z(n19822) );
  XNOR U606 ( .A(n20544), .B(o[212]), .Z(n20535) );
  XNOR U607 ( .A(n20352), .B(o[210]), .Z(n20332) );
  XNOR U608 ( .A(n20431), .B(n20430), .Z(n20433) );
  XNOR U609 ( .A(n20693), .B(n20692), .Z(n20670) );
  XNOR U610 ( .A(n17452), .B(n17451), .Z(n17454) );
  XNOR U611 ( .A(n17460), .B(n17459), .Z(n17476) );
  XNOR U612 ( .A(n17448), .B(n17447), .Z(n17483) );
  XNOR U613 ( .A(n18053), .B(n18052), .Z(n18055) );
  XNOR U614 ( .A(n15008), .B(n15007), .Z(n14984) );
  XNOR U615 ( .A(n15154), .B(n15153), .Z(n15119) );
  XNOR U616 ( .A(n15342), .B(n15341), .Z(n15343) );
  XNOR U617 ( .A(n15348), .B(n15347), .Z(n15349) );
  XNOR U618 ( .A(n15498), .B(n15497), .Z(n15503) );
  XNOR U619 ( .A(n11419), .B(o[111]), .Z(n11391) );
  XNOR U620 ( .A(n11707), .B(n11706), .Z(n11750) );
  XNOR U621 ( .A(n12367), .B(n12366), .Z(n12368) );
  XOR U622 ( .A(n9758), .B(n9757), .Z(n9736) );
  XNOR U623 ( .A(n5455), .B(o[46]), .Z(n5447) );
  XNOR U624 ( .A(n5536), .B(o[47]), .Z(n5508) );
  XNOR U625 ( .A(n5829), .B(n5828), .Z(n5872) );
  XNOR U626 ( .A(n5980), .B(n5979), .Z(n5930) );
  XNOR U627 ( .A(n5989), .B(n5988), .Z(n5990) );
  XNOR U628 ( .A(n2833), .B(n2832), .Z(n2843) );
  XNOR U629 ( .A(n46303), .B(n46302), .Z(n46308) );
  XNOR U630 ( .A(n47049), .B(n47048), .Z(n47050) );
  NAND U631 ( .A(n47144), .B(n47145), .Z(n252) );
  NAND U632 ( .A(n47142), .B(n47143), .Z(n253) );
  NAND U633 ( .A(n252), .B(n253), .Z(n47279) );
  NAND U634 ( .A(n47131), .B(n47130), .Z(n254) );
  NAND U635 ( .A(n47129), .B(n47128), .Z(n255) );
  AND U636 ( .A(n254), .B(n255), .Z(n47271) );
  NAND U637 ( .A(n47336), .B(n47337), .Z(n256) );
  NAND U638 ( .A(n47334), .B(n47335), .Z(n257) );
  NAND U639 ( .A(n256), .B(n257), .Z(n47505) );
  XNOR U640 ( .A(n47401), .B(n47400), .Z(n47402) );
  XNOR U641 ( .A(n47452), .B(n47453), .Z(n47432) );
  XNOR U642 ( .A(n43609), .B(n43608), .Z(n43610) );
  XNOR U643 ( .A(n44561), .B(n44560), .Z(n44562) );
  XNOR U644 ( .A(n44671), .B(o[475]), .Z(n44663) );
  NAND U645 ( .A(n40456), .B(n40457), .Z(n258) );
  NANDN U646 ( .A(n40459), .B(n40458), .Z(n259) );
  AND U647 ( .A(n258), .B(n259), .Z(n40594) );
  XNOR U648 ( .A(n40828), .B(n40827), .Z(n40830) );
  XNOR U649 ( .A(n40842), .B(n40841), .Z(n40792) );
  XOR U650 ( .A(n40710), .B(n40709), .Z(n40720) );
  XNOR U651 ( .A(n40726), .B(n40725), .Z(n40727) );
  XOR U652 ( .A(n40781), .B(n40780), .Z(n40785) );
  NAND U653 ( .A(n41392), .B(n41393), .Z(n260) );
  NAND U654 ( .A(n41390), .B(n41391), .Z(n261) );
  NAND U655 ( .A(n260), .B(n261), .Z(n41468) );
  NAND U656 ( .A(n41389), .B(n41388), .Z(n262) );
  NAND U657 ( .A(n41387), .B(n41386), .Z(n263) );
  AND U658 ( .A(n262), .B(n263), .Z(n41460) );
  NAND U659 ( .A(n37519), .B(n37520), .Z(n264) );
  NAND U660 ( .A(n37517), .B(n37518), .Z(n265) );
  NAND U661 ( .A(n264), .B(n265), .Z(n37619) );
  OR U662 ( .A(n37634), .B(n38583), .Z(n266) );
  NAND U663 ( .A(n37635), .B(n37636), .Z(n267) );
  AND U664 ( .A(n266), .B(n267), .Z(n37742) );
  XNOR U665 ( .A(n37867), .B(n37866), .Z(n37868) );
  XNOR U666 ( .A(n37978), .B(n37977), .Z(n37932) );
  XNOR U667 ( .A(n38514), .B(n38513), .Z(n38516) );
  XNOR U668 ( .A(n34776), .B(n34775), .Z(n34789) );
  XNOR U669 ( .A(n35962), .B(n35961), .Z(n35986) );
  NAND U670 ( .A(n35983), .B(n35982), .Z(n268) );
  NAND U671 ( .A(n35980), .B(n35981), .Z(n269) );
  NAND U672 ( .A(n268), .B(n269), .Z(n36068) );
  NAND U673 ( .A(n31561), .B(n31562), .Z(n270) );
  NAND U674 ( .A(n31603), .B(n33338), .Z(n271) );
  NAND U675 ( .A(n270), .B(n271), .Z(n31629) );
  XNOR U676 ( .A(n32436), .B(n32435), .Z(n32408) );
  XNOR U677 ( .A(n32614), .B(n32613), .Z(n32616) );
  XNOR U678 ( .A(n29284), .B(n29283), .Z(n29238) );
  XNOR U679 ( .A(n30067), .B(n30066), .Z(n30071) );
  XNOR U680 ( .A(n30147), .B(n30146), .Z(n30148) );
  XNOR U681 ( .A(n30247), .B(n30246), .Z(n30248) );
  XNOR U682 ( .A(n30253), .B(n30252), .Z(n30255) );
  NAND U683 ( .A(n26050), .B(n26051), .Z(n272) );
  NAND U684 ( .A(n26423), .B(n26564), .Z(n273) );
  NAND U685 ( .A(n272), .B(n273), .Z(n26212) );
  XNOR U686 ( .A(n22592), .B(n22591), .Z(n22585) );
  XNOR U687 ( .A(n22836), .B(n22835), .Z(n22865) );
  XNOR U688 ( .A(n22845), .B(n22844), .Z(n22847) );
  XNOR U689 ( .A(n22915), .B(n22914), .Z(n22916) );
  XNOR U690 ( .A(n23205), .B(n23204), .Z(n23207) );
  XNOR U691 ( .A(n23973), .B(n23972), .Z(n23958) );
  XNOR U692 ( .A(n24150), .B(n24149), .Z(n24074) );
  XNOR U693 ( .A(n24292), .B(n24291), .Z(n24323) );
  XNOR U694 ( .A(n24477), .B(n24476), .Z(n24478) );
  XNOR U695 ( .A(n24461), .B(n24460), .Z(n24470) );
  NAND U696 ( .A(n19823), .B(n19824), .Z(n274) );
  NAND U697 ( .A(n19997), .B(n21100), .Z(n275) );
  NAND U698 ( .A(n274), .B(n275), .Z(n19857) );
  XNOR U699 ( .A(n20250), .B(n20249), .Z(n20227) );
  XNOR U700 ( .A(n20198), .B(n20197), .Z(n20221) );
  XNOR U701 ( .A(n20559), .B(n20558), .Z(n20595) );
  XNOR U702 ( .A(n20531), .B(n20530), .Z(n20523) );
  XNOR U703 ( .A(n20728), .B(n20727), .Z(n20646) );
  XNOR U704 ( .A(n20792), .B(n20791), .Z(n20779) );
  XNOR U705 ( .A(n21431), .B(n21430), .Z(n21432) );
  NAND U706 ( .A(n17386), .B(n17387), .Z(n276) );
  NANDN U707 ( .A(n17389), .B(n17388), .Z(n277) );
  AND U708 ( .A(n276), .B(n277), .Z(n17422) );
  XNOR U709 ( .A(n17626), .B(n17625), .Z(n17627) );
  XNOR U710 ( .A(n17939), .B(n17938), .Z(n17897) );
  XNOR U711 ( .A(n18137), .B(n18136), .Z(n18138) );
  AND U712 ( .A(n14843), .B(n14842), .Z(n278) );
  AND U713 ( .A(n16334), .B(y[7817]), .Z(n279) );
  NAND U714 ( .A(x[481]), .B(n279), .Z(n280) );
  NANDN U715 ( .A(n278), .B(n280), .Z(n15034) );
  XNOR U716 ( .A(n15520), .B(n15519), .Z(n15521) );
  XNOR U717 ( .A(n15661), .B(n15660), .Z(n15688) );
  XNOR U718 ( .A(n15739), .B(n15738), .Z(n15614) );
  XNOR U719 ( .A(n11367), .B(n11366), .Z(n11338) );
  XNOR U720 ( .A(n11423), .B(n11422), .Z(n11425) );
  XNOR U721 ( .A(n11623), .B(n11622), .Z(n11625) );
  NAND U722 ( .A(n12526), .B(n12525), .Z(n281) );
  NAND U723 ( .A(n12523), .B(n12524), .Z(n282) );
  NAND U724 ( .A(n281), .B(n282), .Z(n12699) );
  NAND U725 ( .A(n12471), .B(n12470), .Z(n283) );
  NAND U726 ( .A(n12469), .B(n12468), .Z(n284) );
  AND U727 ( .A(n283), .B(n284), .Z(n12635) );
  NAND U728 ( .A(n12484), .B(n12485), .Z(n285) );
  NAND U729 ( .A(n12482), .B(n12483), .Z(n286) );
  NAND U730 ( .A(n285), .B(n286), .Z(n12643) );
  NAND U731 ( .A(n12704), .B(n12703), .Z(n287) );
  NANDN U732 ( .A(n12702), .B(n12701), .Z(n288) );
  AND U733 ( .A(n287), .B(n288), .Z(n12866) );
  XNOR U734 ( .A(n8309), .B(n8308), .Z(n8310) );
  XNOR U735 ( .A(n8860), .B(n8859), .Z(n8862) );
  XNOR U736 ( .A(n8922), .B(n9076), .Z(n8894) );
  XNOR U737 ( .A(n9096), .B(n9095), .Z(n9050) );
  XNOR U738 ( .A(n9088), .B(n9087), .Z(n9090) );
  XNOR U739 ( .A(n9878), .B(n9877), .Z(n9913) );
  XOR U740 ( .A(n10112), .B(n10111), .Z(n10114) );
  XNOR U741 ( .A(n5540), .B(n5539), .Z(n5542) );
  XNOR U742 ( .A(n5745), .B(n5744), .Z(n5747) );
  XNOR U743 ( .A(n6123), .B(n6122), .Z(n6077) );
  XOR U744 ( .A(n6052), .B(n6051), .Z(n6044) );
  XNOR U745 ( .A(n6256), .B(n6255), .Z(n6257) );
  XNOR U746 ( .A(n6880), .B(n6879), .Z(n6911) );
  NAND U747 ( .A(n6739), .B(n6740), .Z(n289) );
  NANDN U748 ( .A(n6742), .B(n6741), .Z(n290) );
  AND U749 ( .A(n289), .B(n290), .Z(n6958) );
  XNOR U750 ( .A(n2464), .B(n3426), .Z(n2457) );
  XNOR U751 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U752 ( .A(n2840), .B(n2839), .Z(n291) );
  NANDN U753 ( .A(n3777), .B(n2838), .Z(n292) );
  NAND U754 ( .A(n291), .B(n292), .Z(n2937) );
  XNOR U755 ( .A(n3048), .B(n3047), .Z(n3014) );
  XOR U756 ( .A(n4185), .B(n4184), .Z(n4114) );
  XNOR U757 ( .A(n4040), .B(n4039), .Z(n4041) );
  XNOR U758 ( .A(n45870), .B(n45869), .Z(n45872) );
  XNOR U759 ( .A(n47079), .B(n47078), .Z(n47080) );
  NAND U760 ( .A(n47605), .B(n47604), .Z(n293) );
  NANDN U761 ( .A(n47603), .B(n47602), .Z(n294) );
  NAND U762 ( .A(n293), .B(n294), .Z(n47780) );
  XNOR U763 ( .A(n47937), .B(n47936), .Z(n47965) );
  NAND U764 ( .A(n43147), .B(n43146), .Z(n295) );
  NANDN U765 ( .A(n43240), .B(n43145), .Z(n296) );
  NAND U766 ( .A(n295), .B(n296), .Z(n43221) );
  NAND U767 ( .A(n43159), .B(n43160), .Z(n297) );
  NANDN U768 ( .A(n43162), .B(n43161), .Z(n298) );
  NAND U769 ( .A(n297), .B(n298), .Z(n43294) );
  NAND U770 ( .A(n43155), .B(n43156), .Z(n299) );
  NANDN U771 ( .A(n43158), .B(n43157), .Z(n300) );
  AND U772 ( .A(n299), .B(n300), .Z(n43263) );
  XNOR U773 ( .A(n44715), .B(n44714), .Z(n44716) );
  XNOR U774 ( .A(n44823), .B(n44822), .Z(n44824) );
  XNOR U775 ( .A(n45176), .B(n45087), .Z(n45089) );
  XNOR U776 ( .A(n40021), .B(n40020), .Z(n40014) );
  XNOR U777 ( .A(n40529), .B(n40528), .Z(n40530) );
  XOR U778 ( .A(n40740), .B(n40739), .Z(n40744) );
  XNOR U779 ( .A(n41260), .B(n41259), .Z(n41261) );
  XNOR U780 ( .A(n42156), .B(n42155), .Z(n42157) );
  XNOR U781 ( .A(n37185), .B(n37184), .Z(n37178) );
  XNOR U782 ( .A(n38125), .B(n38124), .Z(n38127) );
  XNOR U783 ( .A(n38560), .B(n38559), .Z(n38562) );
  XNOR U784 ( .A(n38566), .B(n38565), .Z(n38567) );
  XNOR U785 ( .A(n38951), .B(n38950), .Z(n39005) );
  NAND U786 ( .A(n38933), .B(n38934), .Z(n301) );
  NAND U787 ( .A(n38931), .B(n38932), .Z(n302) );
  NAND U788 ( .A(n301), .B(n302), .Z(n39105) );
  NAND U789 ( .A(n39213), .B(n39212), .Z(n303) );
  NAND U790 ( .A(n39210), .B(n39211), .Z(n304) );
  AND U791 ( .A(n303), .B(n304), .Z(n39469) );
  XNOR U792 ( .A(n34946), .B(n34945), .Z(n34948) );
  AND U793 ( .A(n36128), .B(n36127), .Z(n305) );
  AND U794 ( .A(n36556), .B(x[500]), .Z(n306) );
  NAND U795 ( .A(y[8035]), .B(n306), .Z(n307) );
  NANDN U796 ( .A(n305), .B(n307), .Z(n36309) );
  NAND U797 ( .A(n36142), .B(n36143), .Z(n308) );
  NAND U798 ( .A(n36140), .B(n36141), .Z(n309) );
  NAND U799 ( .A(n308), .B(n309), .Z(n36299) );
  NAND U800 ( .A(n36099), .B(n36098), .Z(n310) );
  NAND U801 ( .A(n36096), .B(n36097), .Z(n311) );
  NAND U802 ( .A(n310), .B(n311), .Z(n36273) );
  NAND U803 ( .A(n36237), .B(n36238), .Z(n312) );
  NAND U804 ( .A(n36239), .B(n36240), .Z(n313) );
  NAND U805 ( .A(n312), .B(n313), .Z(n36463) );
  NAND U806 ( .A(n36135), .B(n36136), .Z(n314) );
  NAND U807 ( .A(n36133), .B(n36134), .Z(n315) );
  NAND U808 ( .A(n314), .B(n315), .Z(n36231) );
  XNOR U809 ( .A(n36157), .B(n36156), .Z(n36159) );
  XNOR U810 ( .A(n31318), .B(n31317), .Z(n31348) );
  NAND U811 ( .A(n31618), .B(n31617), .Z(n316) );
  NAND U812 ( .A(n31726), .B(n31616), .Z(n317) );
  NAND U813 ( .A(n316), .B(n317), .Z(n31706) );
  XNOR U814 ( .A(n32789), .B(n32788), .Z(n32791) );
  XNOR U815 ( .A(n28509), .B(n28508), .Z(n28511) );
  XOR U816 ( .A(n30323), .B(n30322), .Z(n30325) );
  XNOR U817 ( .A(n30395), .B(n30394), .Z(n30396) );
  XNOR U818 ( .A(n30425), .B(n30424), .Z(n30426) );
  XNOR U819 ( .A(n30418), .B(n30417), .Z(n30419) );
  XNOR U820 ( .A(n25529), .B(n25528), .Z(n25522) );
  XNOR U821 ( .A(n25910), .B(n25909), .Z(n25880) );
  NAND U822 ( .A(n26205), .B(n26204), .Z(n318) );
  NAND U823 ( .A(n26203), .B(n26202), .Z(n319) );
  AND U824 ( .A(n318), .B(n319), .Z(n26352) );
  XNOR U825 ( .A(n22877), .B(n22876), .Z(n22878) );
  XNOR U826 ( .A(n23087), .B(n23086), .Z(n23088) );
  XNOR U827 ( .A(n23898), .B(n23897), .Z(n23899) );
  XNOR U828 ( .A(n24162), .B(n24161), .Z(n24166) );
  XNOR U829 ( .A(n24206), .B(n24205), .Z(n24193) );
  XNOR U830 ( .A(n24483), .B(n24482), .Z(n24485) );
  XNOR U831 ( .A(n24200), .B(n24199), .Z(n24241) );
  XNOR U832 ( .A(n24465), .B(n24464), .Z(n24466) );
  XNOR U833 ( .A(n24574), .B(n24573), .Z(n24575) );
  XNOR U834 ( .A(n24569), .B(n24568), .Z(n24626) );
  NAND U835 ( .A(n24382), .B(n24381), .Z(n320) );
  NANDN U836 ( .A(n24380), .B(n24379), .Z(n321) );
  NAND U837 ( .A(n320), .B(n321), .Z(n24620) );
  NAND U838 ( .A(n24440), .B(n24439), .Z(n322) );
  NANDN U839 ( .A(n24438), .B(n24437), .Z(n323) );
  NAND U840 ( .A(n322), .B(n323), .Z(n24537) );
  XNOR U841 ( .A(n24563), .B(n24562), .Z(n24594) );
  XNOR U842 ( .A(n19759), .B(n19758), .Z(n19762) );
  XNOR U843 ( .A(n20114), .B(n20113), .Z(n20169) );
  XNOR U844 ( .A(n20104), .B(n20103), .Z(n20134) );
  XNOR U845 ( .A(n20302), .B(n20301), .Z(n20304) );
  XNOR U846 ( .A(n20386), .B(n20385), .Z(n20388) );
  XOR U847 ( .A(n20474), .B(n20473), .Z(n20468) );
  XNOR U848 ( .A(n20732), .B(n20731), .Z(n20733) );
  XNOR U849 ( .A(n20512), .B(n20511), .Z(n20514) );
  XNOR U850 ( .A(n20607), .B(n20606), .Z(n20608) );
  XNOR U851 ( .A(n20874), .B(n20873), .Z(n20876) );
  XNOR U852 ( .A(n20774), .B(n20773), .Z(n20766) );
  XNOR U853 ( .A(n20997), .B(n20996), .Z(n20998) );
  XNOR U854 ( .A(n21009), .B(n21008), .Z(n21010) );
  XNOR U855 ( .A(n21015), .B(n21014), .Z(n21016) );
  NAND U856 ( .A(n21644), .B(n21645), .Z(n324) );
  NAND U857 ( .A(n21646), .B(n21647), .Z(n325) );
  NAND U858 ( .A(n324), .B(n325), .Z(n21852) );
  XNOR U859 ( .A(n21566), .B(n21565), .Z(n21568) );
  NAND U860 ( .A(n21479), .B(n21478), .Z(n326) );
  NAND U861 ( .A(n21476), .B(n21477), .Z(n327) );
  NAND U862 ( .A(n326), .B(n327), .Z(n21615) );
  XNOR U863 ( .A(n16640), .B(n16639), .Z(n16642) );
  XNOR U864 ( .A(n16847), .B(n16846), .Z(n16877) );
  XNOR U865 ( .A(n17201), .B(n17200), .Z(n17202) );
  NAND U866 ( .A(n17287), .B(n17286), .Z(n328) );
  NAND U867 ( .A(n17284), .B(n17285), .Z(n329) );
  NAND U868 ( .A(n328), .B(n329), .Z(n17398) );
  NAND U869 ( .A(n17367), .B(n17366), .Z(n330) );
  NAND U870 ( .A(n17365), .B(n17364), .Z(n331) );
  AND U871 ( .A(n330), .B(n331), .Z(n17488) );
  NAND U872 ( .A(n17781), .B(n17782), .Z(n332) );
  NAND U873 ( .A(n17779), .B(n17780), .Z(n333) );
  NAND U874 ( .A(n332), .B(n333), .Z(n17977) );
  XOR U875 ( .A(n17869), .B(n17868), .Z(n17861) );
  NAND U876 ( .A(n17974), .B(n17973), .Z(n334) );
  NANDN U877 ( .A(n17972), .B(n17971), .Z(n335) );
  AND U878 ( .A(n334), .B(n335), .Z(n18111) );
  NAND U879 ( .A(n17887), .B(n17888), .Z(n336) );
  NAND U880 ( .A(n17885), .B(n17886), .Z(n337) );
  NAND U881 ( .A(n336), .B(n337), .Z(n18108) );
  XNOR U882 ( .A(n14103), .B(n14102), .Z(n14096) );
  NAND U883 ( .A(n14275), .B(n14276), .Z(n338) );
  NAND U884 ( .A(n14274), .B(n14646), .Z(n339) );
  NAND U885 ( .A(n338), .B(n339), .Z(n14384) );
  XNOR U886 ( .A(n14687), .B(n14686), .Z(n14689) );
  XNOR U887 ( .A(n14786), .B(n14785), .Z(n14787) );
  XNOR U888 ( .A(n15298), .B(n15297), .Z(n15316) );
  XNOR U889 ( .A(n15593), .B(n15592), .Z(n15594) );
  NAND U890 ( .A(n15667), .B(n15666), .Z(n340) );
  NAND U891 ( .A(n15664), .B(n15665), .Z(n341) );
  NAND U892 ( .A(n340), .B(n341), .Z(n15867) );
  NAND U893 ( .A(n16103), .B(n16102), .Z(n342) );
  NAND U894 ( .A(n16100), .B(n16101), .Z(n343) );
  AND U895 ( .A(n342), .B(n343), .Z(n16365) );
  XNOR U896 ( .A(n11132), .B(n11131), .Z(n11135) );
  XNOR U897 ( .A(n11455), .B(n11454), .Z(n11456) );
  XNOR U898 ( .A(n11657), .B(n11656), .Z(n11658) );
  XNOR U899 ( .A(n11613), .B(n11612), .Z(n11663) );
  XOR U900 ( .A(n11893), .B(n11892), .Z(n11897) );
  XNOR U901 ( .A(n11693), .B(n11692), .Z(n11686) );
  XOR U902 ( .A(n11905), .B(n11904), .Z(n11909) );
  XOR U903 ( .A(n12013), .B(n12012), .Z(n12017) );
  XNOR U904 ( .A(n12023), .B(n12022), .Z(n12024) );
  XNOR U905 ( .A(n13132), .B(n13131), .Z(n13134) );
  XNOR U906 ( .A(n8165), .B(n8164), .Z(n8195) );
  XNOR U907 ( .A(n8378), .B(n8377), .Z(n8379) );
  XNOR U908 ( .A(n8354), .B(n8353), .Z(n8302) );
  XOR U909 ( .A(n8254), .B(n8253), .Z(n8275) );
  XNOR U910 ( .A(n8291), .B(n8290), .Z(n8293) );
  XOR U911 ( .A(n8969), .B(n8968), .Z(n8963) );
  XNOR U912 ( .A(n9041), .B(n9040), .Z(n9045) );
  XNOR U913 ( .A(n9235), .B(n9234), .Z(n9236) );
  XNOR U914 ( .A(n5253), .B(n5252), .Z(n5256) );
  XNOR U915 ( .A(n5572), .B(n5571), .Z(n5573) );
  XNOR U916 ( .A(n5779), .B(n5778), .Z(n5780) );
  XNOR U917 ( .A(n5735), .B(n5734), .Z(n5785) );
  XOR U918 ( .A(n6015), .B(n6014), .Z(n6019) );
  XNOR U919 ( .A(n5815), .B(n5814), .Z(n5808) );
  XOR U920 ( .A(n6027), .B(n6026), .Z(n6031) );
  XOR U921 ( .A(n6135), .B(n6134), .Z(n6139) );
  XNOR U922 ( .A(n6145), .B(n6144), .Z(n6146) );
  XOR U923 ( .A(n7157), .B(n7156), .Z(n7159) );
  XNOR U924 ( .A(n7203), .B(n7202), .Z(n7204) );
  XNOR U925 ( .A(n2215), .B(n2214), .Z(n2216) );
  XNOR U926 ( .A(n2392), .B(n3019), .Z(n2372) );
  XNOR U927 ( .A(n2362), .B(n2361), .Z(n2355) );
  XNOR U928 ( .A(n3128), .B(n3127), .Z(n3130) );
  XNOR U929 ( .A(n4321), .B(n4320), .Z(n4323) );
  XNOR U930 ( .A(n4084), .B(n4083), .Z(n4085) );
  NAND U931 ( .A(n45460), .B(n45461), .Z(n344) );
  XOR U932 ( .A(n45460), .B(n45461), .Z(n345) );
  NANDN U933 ( .A(n45530), .B(n345), .Z(n346) );
  NAND U934 ( .A(n344), .B(n346), .Z(n45482) );
  XNOR U935 ( .A(n46335), .B(n46334), .Z(n46336) );
  XNOR U936 ( .A(n47234), .B(n47233), .Z(n47235) );
  XOR U937 ( .A(n47657), .B(n47656), .Z(n47530) );
  XNOR U938 ( .A(n47829), .B(n47828), .Z(n47831) );
  XNOR U939 ( .A(n47958), .B(n47957), .Z(n47854) );
  XNOR U940 ( .A(n47950), .B(n47949), .Z(n47951) );
  XNOR U941 ( .A(n48191), .B(n48190), .Z(n48188) );
  XNOR U942 ( .A(n44458), .B(n44457), .Z(n44459) );
  XNOR U943 ( .A(n44808), .B(n44807), .Z(n44879) );
  NAND U944 ( .A(n44684), .B(n44685), .Z(n347) );
  NAND U945 ( .A(n44682), .B(n44683), .Z(n348) );
  NAND U946 ( .A(n347), .B(n348), .Z(n44884) );
  XOR U947 ( .A(n44861), .B(n44860), .Z(n44903) );
  XNOR U948 ( .A(n45054), .B(n45053), .Z(n44969) );
  NAND U949 ( .A(n45266), .B(n45265), .Z(n349) );
  NAND U950 ( .A(n45267), .B(n45268), .Z(n350) );
  AND U951 ( .A(n349), .B(n350), .Z(n45276) );
  XNOR U952 ( .A(n41024), .B(n41023), .Z(n41018) );
  XNOR U953 ( .A(n41286), .B(n41285), .Z(n41287) );
  XOR U954 ( .A(n42249), .B(n42248), .Z(n42247) );
  XOR U955 ( .A(n42237), .B(n42236), .Z(n42235) );
  XNOR U956 ( .A(n37680), .B(n37679), .Z(n37682) );
  NAND U957 ( .A(n39092), .B(n39091), .Z(n351) );
  NANDN U958 ( .A(n39090), .B(n39089), .Z(n352) );
  NAND U959 ( .A(n351), .B(n352), .Z(n39194) );
  NAND U960 ( .A(n39306), .B(n39307), .Z(n353) );
  NANDN U961 ( .A(n39309), .B(n39308), .Z(n354) );
  AND U962 ( .A(n353), .B(n354), .Z(n39511) );
  NAND U963 ( .A(n39254), .B(n39253), .Z(n355) );
  NAND U964 ( .A(n39252), .B(n39481), .Z(n356) );
  NAND U965 ( .A(n355), .B(n356), .Z(n39346) );
  NAND U966 ( .A(n39068), .B(n39067), .Z(n357) );
  NAND U967 ( .A(n39066), .B(n39065), .Z(n358) );
  AND U968 ( .A(n357), .B(n358), .Z(n39275) );
  NAND U969 ( .A(n36154), .B(n36155), .Z(n359) );
  NAND U970 ( .A(n36152), .B(n36153), .Z(n360) );
  NAND U971 ( .A(n359), .B(n360), .Z(n36197) );
  NAND U972 ( .A(n36305), .B(n36306), .Z(n361) );
  NAND U973 ( .A(n36303), .B(n36304), .Z(n362) );
  NAND U974 ( .A(n361), .B(n362), .Z(n36439) );
  XNOR U975 ( .A(n36434), .B(n36433), .Z(n36435) );
  NAND U976 ( .A(n36469), .B(n36470), .Z(n363) );
  NANDN U977 ( .A(n36472), .B(n36471), .Z(n364) );
  AND U978 ( .A(n363), .B(n364), .Z(n36671) );
  NAND U979 ( .A(n36215), .B(n36214), .Z(n365) );
  NAND U980 ( .A(n36213), .B(n36212), .Z(n366) );
  AND U981 ( .A(n365), .B(n366), .Z(n36449) );
  XNOR U982 ( .A(n31080), .B(n31079), .Z(n31082) );
  NAND U983 ( .A(n31067), .B(n31068), .Z(n367) );
  NAND U984 ( .A(n31066), .B(n31129), .Z(n368) );
  NAND U985 ( .A(n367), .B(n368), .Z(n31110) );
  NAND U986 ( .A(n31947), .B(n31161), .Z(n369) );
  NANDN U987 ( .A(n31163), .B(n31162), .Z(n370) );
  AND U988 ( .A(n369), .B(n370), .Z(n31201) );
  XOR U989 ( .A(n32628), .B(n32627), .Z(n32506) );
  XNOR U990 ( .A(n33360), .B(n33359), .Z(n33362) );
  XNOR U991 ( .A(n33610), .B(n33609), .Z(n33572) );
  XNOR U992 ( .A(n33392), .B(n33391), .Z(n33393) );
  XNOR U993 ( .A(n33560), .B(n33559), .Z(n33561) );
  XOR U994 ( .A(n33285), .B(n33284), .Z(n33271) );
  XNOR U995 ( .A(n30447), .B(n30446), .Z(n30468) );
  XNOR U996 ( .A(n30433), .B(n30432), .Z(n30481) );
  XNOR U997 ( .A(n30400), .B(n30401), .Z(n30487) );
  XNOR U998 ( .A(n30542), .B(n30541), .Z(n30548) );
  XNOR U999 ( .A(n30679), .B(n30678), .Z(n30638) );
  XNOR U1000 ( .A(n25652), .B(n25651), .Z(n25653) );
  XNOR U1001 ( .A(n26223), .B(n26222), .Z(n26226) );
  XNOR U1002 ( .A(n27511), .B(n27510), .Z(n27512) );
  XOR U1003 ( .A(n27404), .B(n27403), .Z(n27390) );
  XNOR U1004 ( .A(n27596), .B(n27595), .Z(n27601) );
  XNOR U1005 ( .A(n27731), .B(n27730), .Z(n27692) );
  XNOR U1006 ( .A(n22909), .B(n22908), .Z(n22910) );
  XNOR U1007 ( .A(n24765), .B(n24764), .Z(n24680) );
  NAND U1008 ( .A(n24630), .B(n24631), .Z(n371) );
  NANDN U1009 ( .A(n24633), .B(n24632), .Z(n372) );
  NAND U1010 ( .A(n371), .B(n372), .Z(n24756) );
  XNOR U1011 ( .A(n24813), .B(n24812), .Z(n24775) );
  XNOR U1012 ( .A(n19480), .B(n19479), .Z(n19482) );
  XOR U1013 ( .A(n20740), .B(n20739), .Z(n20635) );
  NAND U1014 ( .A(n21563), .B(n21564), .Z(n373) );
  NAND U1015 ( .A(n21561), .B(n21562), .Z(n374) );
  NAND U1016 ( .A(n373), .B(n374), .Z(n21606) );
  NAND U1017 ( .A(n21706), .B(n21705), .Z(n375) );
  NAND U1018 ( .A(n21703), .B(n21704), .Z(n376) );
  NAND U1019 ( .A(n375), .B(n376), .Z(n21836) );
  XNOR U1020 ( .A(n21829), .B(n21828), .Z(n21830) );
  NAND U1021 ( .A(n21681), .B(n21682), .Z(n377) );
  NAND U1022 ( .A(n21679), .B(n21680), .Z(n378) );
  NAND U1023 ( .A(n377), .B(n378), .Z(n21839) );
  NAND U1024 ( .A(n21879), .B(n21880), .Z(n379) );
  NANDN U1025 ( .A(n21882), .B(n21881), .Z(n380) );
  AND U1026 ( .A(n379), .B(n380), .Z(n22085) );
  NAND U1027 ( .A(n21639), .B(n21638), .Z(n381) );
  NAND U1028 ( .A(n21637), .B(n21636), .Z(n382) );
  AND U1029 ( .A(n381), .B(n382), .Z(n21844) );
  NAND U1030 ( .A(n21685), .B(n21686), .Z(n383) );
  NAND U1031 ( .A(n21683), .B(n21684), .Z(n384) );
  NAND U1032 ( .A(n383), .B(n384), .Z(n21742) );
  NAND U1033 ( .A(n21695), .B(n21696), .Z(n385) );
  NAND U1034 ( .A(n21693), .B(n21694), .Z(n386) );
  NAND U1035 ( .A(n385), .B(n386), .Z(n21740) );
  XNOR U1036 ( .A(n17233), .B(n17232), .Z(n17234) );
  XNOR U1037 ( .A(n18408), .B(n18407), .Z(n18271) );
  XNOR U1038 ( .A(n18567), .B(n18566), .Z(n18425) );
  XNOR U1039 ( .A(n18864), .B(n18863), .Z(n18865) );
  XOR U1040 ( .A(n18756), .B(n18755), .Z(n18742) );
  XNOR U1041 ( .A(n18945), .B(n18944), .Z(n18950) );
  XNOR U1042 ( .A(n19081), .B(n19080), .Z(n19040) );
  XNOR U1043 ( .A(n15745), .B(n15744), .Z(n15611) );
  NAND U1044 ( .A(n15871), .B(n15872), .Z(n387) );
  NAND U1045 ( .A(n15869), .B(n15870), .Z(n388) );
  NAND U1046 ( .A(n387), .B(n388), .Z(n16012) );
  NAND U1047 ( .A(n15975), .B(n15976), .Z(n389) );
  NAND U1048 ( .A(n15973), .B(n15974), .Z(n390) );
  NAND U1049 ( .A(n389), .B(n390), .Z(n16153) );
  NAND U1050 ( .A(n16176), .B(n16177), .Z(n391) );
  NANDN U1051 ( .A(n16179), .B(n16178), .Z(n392) );
  NAND U1052 ( .A(n391), .B(n392), .Z(n16422) );
  NAND U1053 ( .A(n16138), .B(n16137), .Z(n393) );
  NAND U1054 ( .A(n16135), .B(n16136), .Z(n394) );
  NAND U1055 ( .A(n393), .B(n394), .Z(n16235) );
  XNOR U1056 ( .A(n11156), .B(n11155), .Z(n11157) );
  XNOR U1057 ( .A(n11516), .B(n11515), .Z(n11484) );
  XOR U1058 ( .A(n12590), .B(n12589), .Z(n12583) );
  XNOR U1059 ( .A(n13355), .B(n13354), .Z(n13329) );
  XNOR U1060 ( .A(n13152), .B(n13151), .Z(n13191) );
  XNOR U1061 ( .A(n8764), .B(n8763), .Z(n8765) );
  XNOR U1062 ( .A(n9108), .B(n9107), .Z(n9112) );
  XNOR U1063 ( .A(n10120), .B(n10119), .Z(n9983) );
  NAND U1064 ( .A(n10061), .B(n10062), .Z(n395) );
  NAND U1065 ( .A(n10059), .B(n10060), .Z(n396) );
  NAND U1066 ( .A(n395), .B(n396), .Z(n10250) );
  XOR U1067 ( .A(n10321), .B(n10320), .Z(n10323) );
  XNOR U1068 ( .A(n10406), .B(n10405), .Z(n10407) );
  XNOR U1069 ( .A(n10700), .B(n10699), .Z(n10696) );
  XNOR U1070 ( .A(n10418), .B(n10417), .Z(n10420) );
  XNOR U1071 ( .A(n10663), .B(n10662), .Z(n10660) );
  NAND U1072 ( .A(n5848), .B(n5045), .Z(n397) );
  NANDN U1073 ( .A(n5047), .B(n5046), .Z(n398) );
  AND U1074 ( .A(n397), .B(n398), .Z(n5085) );
  XNOR U1075 ( .A(n5600), .B(n5599), .Z(n5601) );
  XNOR U1076 ( .A(n7268), .B(n7267), .Z(n7269) );
  XNOR U1077 ( .A(n7284), .B(n7283), .Z(n7305) );
  XNOR U1078 ( .A(n7257), .B(n7256), .Z(n7317) );
  XNOR U1079 ( .A(n7237), .B(n7238), .Z(n7324) );
  XNOR U1080 ( .A(n7377), .B(n7376), .Z(n7383) );
  XNOR U1081 ( .A(n7513), .B(n7512), .Z(n7472) );
  NAND U1082 ( .A(n2992), .B(n2991), .Z(n399) );
  NANDN U1083 ( .A(n2990), .B(n2989), .Z(n400) );
  AND U1084 ( .A(n399), .B(n400), .Z(n3197) );
  XNOR U1085 ( .A(n3259), .B(n3258), .Z(n3233) );
  XNOR U1086 ( .A(n3332), .B(n3331), .Z(n3227) );
  XNOR U1087 ( .A(n3452), .B(n3451), .Z(n3457) );
  XOR U1088 ( .A(n3762), .B(n3761), .Z(n3755) );
  XNOR U1089 ( .A(n4215), .B(n4214), .Z(n4078) );
  XNOR U1090 ( .A(n4441), .B(n4440), .Z(n4542) );
  XOR U1091 ( .A(n4412), .B(n4411), .Z(n4414) );
  XNOR U1092 ( .A(n4241), .B(n4240), .Z(n4234) );
  XNOR U1093 ( .A(n4249), .B(n4248), .Z(n4251) );
  XOR U1094 ( .A(n45614), .B(n45613), .Z(n45653) );
  XOR U1095 ( .A(n48225), .B(n48224), .Z(n48223) );
  XOR U1096 ( .A(n47836), .B(n47835), .Z(n401) );
  NANDN U1097 ( .A(n47837), .B(n401), .Z(n402) );
  NAND U1098 ( .A(n47836), .B(n47835), .Z(n403) );
  AND U1099 ( .A(n402), .B(n403), .Z(n48259) );
  XOR U1100 ( .A(n42720), .B(n42719), .Z(n42761) );
  XNOR U1101 ( .A(n43039), .B(n43038), .Z(n43041) );
  XNOR U1102 ( .A(n43623), .B(n43622), .Z(n43626) );
  XNOR U1103 ( .A(n45048), .B(n45047), .Z(n44961) );
  XNOR U1104 ( .A(n45136), .B(n45135), .Z(n45133) );
  XOR U1105 ( .A(n44934), .B(n44935), .Z(n404) );
  NANDN U1106 ( .A(n44936), .B(n404), .Z(n405) );
  NAND U1107 ( .A(n44934), .B(n44935), .Z(n406) );
  AND U1108 ( .A(n405), .B(n406), .Z(n45365) );
  XOR U1109 ( .A(n39622), .B(n39623), .Z(n407) );
  NANDN U1110 ( .A(n39624), .B(n407), .Z(n408) );
  NAND U1111 ( .A(n39622), .B(n39623), .Z(n409) );
  AND U1112 ( .A(n408), .B(n409), .Z(n39645) );
  NAND U1113 ( .A(n39715), .B(n39714), .Z(n410) );
  NAND U1114 ( .A(n39713), .B(n39712), .Z(n411) );
  AND U1115 ( .A(n410), .B(n411), .Z(n39725) );
  XNOR U1116 ( .A(n40854), .B(n40853), .Z(n40869) );
  XNOR U1117 ( .A(n42445), .B(n42444), .Z(n42442) );
  NAND U1118 ( .A(n36820), .B(n36819), .Z(n412) );
  XOR U1119 ( .A(n36820), .B(n36819), .Z(n413) );
  NANDN U1120 ( .A(n36889), .B(n413), .Z(n414) );
  NAND U1121 ( .A(n412), .B(n414), .Z(n36865) );
  XNOR U1122 ( .A(n37383), .B(n37382), .Z(n37385) );
  XOR U1123 ( .A(n37664), .B(n37663), .Z(n37666) );
  NAND U1124 ( .A(n37872), .B(n37873), .Z(n415) );
  NANDN U1125 ( .A(n37875), .B(n37874), .Z(n416) );
  AND U1126 ( .A(n415), .B(n416), .Z(n38009) );
  NAND U1127 ( .A(n39134), .B(n39133), .Z(n417) );
  NAND U1128 ( .A(n39131), .B(n39132), .Z(n418) );
  NAND U1129 ( .A(n417), .B(n418), .Z(n39267) );
  NAND U1130 ( .A(n39193), .B(n39192), .Z(n419) );
  NANDN U1131 ( .A(n39191), .B(n39190), .Z(n420) );
  AND U1132 ( .A(n419), .B(n420), .Z(n39563) );
  XOR U1133 ( .A(n39553), .B(n39552), .Z(n39551) );
  NAND U1134 ( .A(n39217), .B(n39216), .Z(n421) );
  NAND U1135 ( .A(n39214), .B(n39215), .Z(n422) );
  NAND U1136 ( .A(n421), .B(n422), .Z(n39323) );
  XOR U1137 ( .A(n34139), .B(n34138), .Z(n34180) );
  NAND U1138 ( .A(n36270), .B(n36269), .Z(n423) );
  NANDN U1139 ( .A(n36268), .B(n36267), .Z(n424) );
  NAND U1140 ( .A(n423), .B(n424), .Z(n36356) );
  NAND U1141 ( .A(n36533), .B(n36534), .Z(n425) );
  NANDN U1142 ( .A(n36535), .B(n36569), .Z(n426) );
  AND U1143 ( .A(n425), .B(n426), .Z(n427) );
  XOR U1144 ( .A(n36604), .B(n36603), .Z(n428) );
  XNOR U1145 ( .A(n36548), .B(n36547), .Z(n429) );
  XNOR U1146 ( .A(n428), .B(n429), .Z(n430) );
  XOR U1147 ( .A(n36638), .B(n36637), .Z(n431) );
  XNOR U1148 ( .A(n36624), .B(n36623), .Z(n432) );
  XNOR U1149 ( .A(n431), .B(n432), .Z(n433) );
  XOR U1150 ( .A(n36666), .B(n36665), .Z(n434) );
  XNOR U1151 ( .A(n36652), .B(n36651), .Z(n435) );
  XNOR U1152 ( .A(n434), .B(n435), .Z(n436) );
  XOR U1153 ( .A(n433), .B(n436), .Z(n437) );
  XNOR U1154 ( .A(n427), .B(n430), .Z(n438) );
  XNOR U1155 ( .A(n437), .B(n438), .Z(n439) );
  NAND U1156 ( .A(n36530), .B(n36529), .Z(n440) );
  NAND U1157 ( .A(n36531), .B(n36532), .Z(n441) );
  NAND U1158 ( .A(n440), .B(n441), .Z(n442) );
  XNOR U1159 ( .A(n439), .B(n442), .Z(n36667) );
  XNOR U1160 ( .A(n31244), .B(n31243), .Z(n31245) );
  NAND U1161 ( .A(n31657), .B(n31656), .Z(n443) );
  NANDN U1162 ( .A(n31655), .B(n31654), .Z(n444) );
  AND U1163 ( .A(n443), .B(n444), .Z(n31690) );
  XNOR U1164 ( .A(n32107), .B(n32106), .Z(n32110) );
  XNOR U1165 ( .A(n33507), .B(n33506), .Z(n33475) );
  XNOR U1166 ( .A(n33850), .B(n33849), .Z(n33864) );
  NAND U1167 ( .A(n28109), .B(n28108), .Z(n445) );
  XOR U1168 ( .A(n28109), .B(n28108), .Z(n446) );
  NANDN U1169 ( .A(n28169), .B(n446), .Z(n447) );
  NAND U1170 ( .A(n445), .B(n447), .Z(n28145) );
  XNOR U1171 ( .A(n25727), .B(n25726), .Z(n25729) );
  XNOR U1172 ( .A(n25936), .B(n25935), .Z(n26023) );
  XOR U1173 ( .A(n27979), .B(n27978), .Z(n27977) );
  XOR U1174 ( .A(n27755), .B(n27754), .Z(n27753) );
  XNOR U1175 ( .A(n22218), .B(n22217), .Z(n22222) );
  XNOR U1176 ( .A(n22995), .B(n22994), .Z(n22997) );
  XNOR U1177 ( .A(n24335), .B(n24334), .Z(n24337) );
  NAND U1178 ( .A(n24513), .B(n24512), .Z(n448) );
  NANDN U1179 ( .A(n24511), .B(n24510), .Z(n449) );
  AND U1180 ( .A(n448), .B(n449), .Z(n24672) );
  NAND U1181 ( .A(n25021), .B(n25022), .Z(n25026) );
  NAND U1182 ( .A(n24645), .B(n24644), .Z(n450) );
  XOR U1183 ( .A(n24645), .B(n24644), .Z(n451) );
  NANDN U1184 ( .A(n24646), .B(n451), .Z(n452) );
  NAND U1185 ( .A(n450), .B(n452), .Z(n25072) );
  XOR U1186 ( .A(n19528), .B(n19466), .Z(n453) );
  NANDN U1187 ( .A(n19467), .B(n453), .Z(n454) );
  NAND U1188 ( .A(n19528), .B(n19466), .Z(n455) );
  AND U1189 ( .A(n454), .B(n455), .Z(n19507) );
  XNOR U1190 ( .A(n19907), .B(n19906), .Z(n19908) );
  XOR U1191 ( .A(n19849), .B(n19848), .Z(n456) );
  NANDN U1192 ( .A(n19847), .B(n456), .Z(n457) );
  NAND U1193 ( .A(n19849), .B(n19848), .Z(n458) );
  AND U1194 ( .A(n457), .B(n458), .Z(n19914) );
  NAND U1195 ( .A(n20051), .B(n20050), .Z(n459) );
  NANDN U1196 ( .A(n20049), .B(n20048), .Z(n460) );
  AND U1197 ( .A(n459), .B(n460), .Z(n20080) );
  XNOR U1198 ( .A(n20505), .B(n20504), .Z(n20507) );
  XNOR U1199 ( .A(n20880), .B(n20879), .Z(n20881) );
  NAND U1200 ( .A(n21666), .B(n21665), .Z(n461) );
  NANDN U1201 ( .A(n21664), .B(n21663), .Z(n462) );
  NAND U1202 ( .A(n461), .B(n462), .Z(n21750) );
  NAND U1203 ( .A(n21932), .B(n21931), .Z(n463) );
  NAND U1204 ( .A(n21968), .B(n21933), .Z(n464) );
  AND U1205 ( .A(n463), .B(n464), .Z(n465) );
  XOR U1206 ( .A(n22002), .B(n22001), .Z(n466) );
  XNOR U1207 ( .A(n21946), .B(n21945), .Z(n467) );
  XNOR U1208 ( .A(n466), .B(n467), .Z(n468) );
  XOR U1209 ( .A(n22052), .B(n22051), .Z(n469) );
  XNOR U1210 ( .A(n22040), .B(n22039), .Z(n470) );
  XNOR U1211 ( .A(n469), .B(n470), .Z(n471) );
  XOR U1212 ( .A(n22080), .B(n22079), .Z(n472) );
  XNOR U1213 ( .A(n22066), .B(n22065), .Z(n473) );
  XNOR U1214 ( .A(n472), .B(n473), .Z(n474) );
  XOR U1215 ( .A(n471), .B(n474), .Z(n475) );
  XNOR U1216 ( .A(n465), .B(n468), .Z(n476) );
  XNOR U1217 ( .A(n475), .B(n476), .Z(n477) );
  NAND U1218 ( .A(n21928), .B(n21927), .Z(n478) );
  NAND U1219 ( .A(n21929), .B(n21930), .Z(n479) );
  NAND U1220 ( .A(n478), .B(n479), .Z(n480) );
  XNOR U1221 ( .A(n477), .B(n480), .Z(n22081) );
  NAND U1222 ( .A(n16567), .B(n16566), .Z(n481) );
  XOR U1223 ( .A(n16567), .B(n16566), .Z(n482) );
  NANDN U1224 ( .A(n16628), .B(n482), .Z(n483) );
  NAND U1225 ( .A(n481), .B(n483), .Z(n16603) );
  NAND U1226 ( .A(n13751), .B(n13750), .Z(n484) );
  XOR U1227 ( .A(n13751), .B(n13750), .Z(n485) );
  NANDN U1228 ( .A(n13811), .B(n485), .Z(n486) );
  NAND U1229 ( .A(n484), .B(n486), .Z(n13787) );
  XNOR U1230 ( .A(n14307), .B(n14306), .Z(n14309) );
  XNOR U1231 ( .A(n15191), .B(n15190), .Z(n15319) );
  NAND U1232 ( .A(n15963), .B(n15964), .Z(n487) );
  NAND U1233 ( .A(n15961), .B(n15962), .Z(n488) );
  NAND U1234 ( .A(n487), .B(n488), .Z(n16087) );
  NAND U1235 ( .A(n16160), .B(n16161), .Z(n489) );
  NANDN U1236 ( .A(n16163), .B(n16162), .Z(n490) );
  AND U1237 ( .A(n489), .B(n490), .Z(n16432) );
  XOR U1238 ( .A(n11213), .B(n11212), .Z(n11224) );
  XNOR U1239 ( .A(n11234), .B(n11233), .Z(n11235) );
  XNOR U1240 ( .A(n11479), .B(n11478), .Z(n11566) );
  XNOR U1241 ( .A(n13323), .B(n13322), .Z(n13324) );
  XNOR U1242 ( .A(n13610), .B(n13609), .Z(n13624) );
  XNOR U1243 ( .A(n7872), .B(n7871), .Z(n7876) );
  XOR U1244 ( .A(n8035), .B(n8034), .Z(n8037) );
  XNOR U1245 ( .A(n9140), .B(n9139), .Z(n9127) );
  XOR U1246 ( .A(n9377), .B(n9376), .Z(n9379) );
  XNOR U1247 ( .A(n10695), .B(n10694), .Z(n10692) );
  XNOR U1248 ( .A(n4917), .B(n4916), .Z(n4921) );
  XNOR U1249 ( .A(n5079), .B(n5078), .Z(n5080) );
  XNOR U1250 ( .A(n5413), .B(n5412), .Z(n5414) );
  XNOR U1251 ( .A(n5687), .B(n5686), .Z(n5689) );
  XOR U1252 ( .A(n2136), .B(n2135), .Z(n2149) );
  XOR U1253 ( .A(n2167), .B(n2166), .Z(n2157) );
  XNOR U1254 ( .A(n2503), .B(n2502), .Z(n2585) );
  XNOR U1255 ( .A(n2878), .B(n2877), .Z(n2970) );
  XNOR U1256 ( .A(n4557), .B(n4556), .Z(n4558) );
  NANDN U1257 ( .A(n45437), .B(n45439), .Z(n491) );
  OR U1258 ( .A(n45439), .B(n45440), .Z(n492) );
  NAND U1259 ( .A(n45438), .B(n492), .Z(n493) );
  NAND U1260 ( .A(n491), .B(n493), .Z(n45479) );
  NAND U1261 ( .A(n47520), .B(n47521), .Z(n494) );
  XOR U1262 ( .A(n47520), .B(n47521), .Z(n495) );
  NANDN U1263 ( .A(n47519), .B(n495), .Z(n496) );
  NAND U1264 ( .A(n494), .B(n496), .Z(n47666) );
  XNOR U1265 ( .A(n48277), .B(n48276), .Z(n48274) );
  NAND U1266 ( .A(n42902), .B(n42901), .Z(n497) );
  NAND U1267 ( .A(n42900), .B(n42899), .Z(n498) );
  AND U1268 ( .A(n497), .B(n498), .Z(n43036) );
  XOR U1269 ( .A(n43412), .B(n43413), .Z(n499) );
  NANDN U1270 ( .A(n43414), .B(n499), .Z(n500) );
  NAND U1271 ( .A(n43412), .B(n43413), .Z(n501) );
  AND U1272 ( .A(n500), .B(n501), .Z(n43632) );
  XNOR U1273 ( .A(n43755), .B(n43754), .Z(n43751) );
  NAND U1274 ( .A(n44298), .B(n44299), .Z(n502) );
  XOR U1275 ( .A(n44298), .B(n44299), .Z(n503) );
  NANDN U1276 ( .A(n44297), .B(n503), .Z(n504) );
  NAND U1277 ( .A(n502), .B(n504), .Z(n44448) );
  XNOR U1278 ( .A(n45384), .B(n45383), .Z(n45382) );
  XNOR U1279 ( .A(n39802), .B(n39801), .Z(n39798) );
  NAND U1280 ( .A(n40239), .B(n40240), .Z(n505) );
  XOR U1281 ( .A(n40239), .B(n40240), .Z(n506) );
  NANDN U1282 ( .A(n40238), .B(n506), .Z(n507) );
  NAND U1283 ( .A(n505), .B(n507), .Z(n40413) );
  XOR U1284 ( .A(n40638), .B(n40639), .Z(n508) );
  NANDN U1285 ( .A(n40640), .B(n508), .Z(n509) );
  NAND U1286 ( .A(n40638), .B(n40639), .Z(n510) );
  AND U1287 ( .A(n509), .B(n510), .Z(n40864) );
  NAND U1288 ( .A(n41863), .B(n41864), .Z(n511) );
  XOR U1289 ( .A(n41863), .B(n41864), .Z(n512) );
  NANDN U1290 ( .A(n41862), .B(n512), .Z(n513) );
  NAND U1291 ( .A(n511), .B(n513), .Z(n41877) );
  NAND U1292 ( .A(n41875), .B(n41874), .Z(n514) );
  NAND U1293 ( .A(n41873), .B(n41872), .Z(n515) );
  AND U1294 ( .A(n514), .B(n515), .Z(n42038) );
  XNOR U1295 ( .A(n42473), .B(n42472), .Z(n42470) );
  XOR U1296 ( .A(n36831), .B(n36832), .Z(n516) );
  NANDN U1297 ( .A(n36833), .B(n516), .Z(n517) );
  NAND U1298 ( .A(n36831), .B(n36832), .Z(n518) );
  AND U1299 ( .A(n517), .B(n518), .Z(n36872) );
  XOR U1300 ( .A(n37303), .B(n37304), .Z(n519) );
  NANDN U1301 ( .A(n37305), .B(n519), .Z(n520) );
  NAND U1302 ( .A(n37303), .B(n37304), .Z(n521) );
  AND U1303 ( .A(n520), .B(n521), .Z(n37389) );
  XOR U1304 ( .A(n37888), .B(n37889), .Z(n522) );
  NANDN U1305 ( .A(n37890), .B(n522), .Z(n523) );
  NAND U1306 ( .A(n37888), .B(n37889), .Z(n524) );
  AND U1307 ( .A(n523), .B(n524), .Z(n38005) );
  XOR U1308 ( .A(n39157), .B(n39158), .Z(n525) );
  NANDN U1309 ( .A(n39159), .B(n525), .Z(n526) );
  NAND U1310 ( .A(n39157), .B(n39158), .Z(n527) );
  AND U1311 ( .A(n526), .B(n527), .Z(n39573) );
  XOR U1312 ( .A(n34843), .B(n34842), .Z(n528) );
  NANDN U1313 ( .A(n34841), .B(n528), .Z(n529) );
  NAND U1314 ( .A(n34843), .B(n34842), .Z(n530) );
  AND U1315 ( .A(n529), .B(n530), .Z(n34958) );
  XNOR U1316 ( .A(n36494), .B(n36493), .Z(n36492) );
  NAND U1317 ( .A(n31192), .B(n31193), .Z(n531) );
  XOR U1318 ( .A(n31192), .B(n31193), .Z(n532) );
  NANDN U1319 ( .A(n31191), .B(n532), .Z(n533) );
  NAND U1320 ( .A(n531), .B(n533), .Z(n31250) );
  NAND U1321 ( .A(n31897), .B(n31898), .Z(n534) );
  XOR U1322 ( .A(n31897), .B(n31898), .Z(n535) );
  NANDN U1323 ( .A(n31896), .B(n535), .Z(n536) );
  NAND U1324 ( .A(n534), .B(n536), .Z(n32117) );
  XNOR U1325 ( .A(n32239), .B(n32238), .Z(n32235) );
  XOR U1326 ( .A(n33880), .B(n33879), .Z(n33900) );
  NAND U1327 ( .A(n28102), .B(n28103), .Z(n537) );
  XOR U1328 ( .A(n28102), .B(n28103), .Z(n538) );
  NANDN U1329 ( .A(n28101), .B(n538), .Z(n539) );
  NAND U1330 ( .A(n537), .B(n539), .Z(n28151) );
  XOR U1331 ( .A(n29079), .B(n29080), .Z(n540) );
  NANDN U1332 ( .A(n29081), .B(n540), .Z(n541) );
  NAND U1333 ( .A(n29079), .B(n29080), .Z(n542) );
  AND U1334 ( .A(n541), .B(n542), .Z(n29083) );
  XNOR U1335 ( .A(n29317), .B(n29316), .Z(n29313) );
  XNOR U1336 ( .A(n30691), .B(n30690), .Z(n30689) );
  XOR U1337 ( .A(n25647), .B(n25648), .Z(n543) );
  NANDN U1338 ( .A(n25649), .B(n543), .Z(n544) );
  NAND U1339 ( .A(n25647), .B(n25648), .Z(n545) );
  AND U1340 ( .A(n544), .B(n545), .Z(n25733) );
  XOR U1341 ( .A(n28020), .B(n28021), .Z(n28022) );
  XNOR U1342 ( .A(n25090), .B(n25089), .Z(n25087) );
  NAND U1343 ( .A(n19460), .B(n19461), .Z(n546) );
  XOR U1344 ( .A(n19460), .B(n19461), .Z(n547) );
  NANDN U1345 ( .A(n19459), .B(n547), .Z(n548) );
  NAND U1346 ( .A(n546), .B(n548), .Z(n19504) );
  NAND U1347 ( .A(n19596), .B(n19597), .Z(n549) );
  XOR U1348 ( .A(n19596), .B(n19597), .Z(n550) );
  NANDN U1349 ( .A(n19595), .B(n550), .Z(n551) );
  NAND U1350 ( .A(n549), .B(n551), .Z(n19648) );
  XOR U1351 ( .A(n20070), .B(n20071), .Z(n552) );
  NANDN U1352 ( .A(n20072), .B(n552), .Z(n553) );
  NAND U1353 ( .A(n20070), .B(n20071), .Z(n554) );
  AND U1354 ( .A(n553), .B(n554), .Z(n20087) );
  NAND U1355 ( .A(n20287), .B(n20288), .Z(n555) );
  XOR U1356 ( .A(n20287), .B(n20288), .Z(n556) );
  NANDN U1357 ( .A(n20286), .B(n556), .Z(n557) );
  NAND U1358 ( .A(n555), .B(n557), .Z(n20502) );
  NAND U1359 ( .A(n20750), .B(n20751), .Z(n558) );
  XOR U1360 ( .A(n20750), .B(n20751), .Z(n559) );
  NANDN U1361 ( .A(n20749), .B(n559), .Z(n560) );
  NAND U1362 ( .A(n558), .B(n560), .Z(n20886) );
  NAND U1363 ( .A(n21174), .B(n21175), .Z(n561) );
  XOR U1364 ( .A(n21174), .B(n21175), .Z(n562) );
  NANDN U1365 ( .A(n21176), .B(n562), .Z(n563) );
  NAND U1366 ( .A(n561), .B(n563), .Z(n21455) );
  XOR U1367 ( .A(n21723), .B(n21722), .Z(n564) );
  NANDN U1368 ( .A(n21721), .B(n564), .Z(n565) );
  NAND U1369 ( .A(n21723), .B(n21722), .Z(n566) );
  AND U1370 ( .A(n565), .B(n566), .Z(n21726) );
  XNOR U1371 ( .A(n21892), .B(n21891), .Z(n21890) );
  NAND U1372 ( .A(n16560), .B(n16561), .Z(n567) );
  XOR U1373 ( .A(n16560), .B(n16561), .Z(n568) );
  NANDN U1374 ( .A(n16559), .B(n568), .Z(n569) );
  NAND U1375 ( .A(n567), .B(n569), .Z(n16609) );
  NAND U1376 ( .A(n17533), .B(n17534), .Z(n570) );
  XOR U1377 ( .A(n17533), .B(n17534), .Z(n571) );
  NANDN U1378 ( .A(n17532), .B(n571), .Z(n572) );
  NAND U1379 ( .A(n570), .B(n572), .Z(n17650) );
  NAND U1380 ( .A(n18414), .B(n18411), .Z(n573) );
  NANDN U1381 ( .A(n18414), .B(n18413), .Z(n574) );
  NANDN U1382 ( .A(n18412), .B(n574), .Z(n575) );
  NAND U1383 ( .A(n573), .B(n575), .Z(n18571) );
  NAND U1384 ( .A(n18906), .B(n18907), .Z(n576) );
  XOR U1385 ( .A(n18906), .B(n18907), .Z(n577) );
  NANDN U1386 ( .A(n18905), .B(n577), .Z(n578) );
  NAND U1387 ( .A(n576), .B(n578), .Z(n18909) );
  XOR U1388 ( .A(n19372), .B(n19373), .Z(n19371) );
  NAND U1389 ( .A(n13744), .B(n13745), .Z(n579) );
  XOR U1390 ( .A(n13744), .B(n13745), .Z(n580) );
  NANDN U1391 ( .A(n13743), .B(n580), .Z(n581) );
  NAND U1392 ( .A(n579), .B(n581), .Z(n13794) );
  XNOR U1393 ( .A(n14226), .B(n14225), .Z(n14232) );
  XOR U1394 ( .A(n14580), .B(n14581), .Z(n582) );
  NANDN U1395 ( .A(n14582), .B(n582), .Z(n583) );
  NAND U1396 ( .A(n14580), .B(n14581), .Z(n584) );
  AND U1397 ( .A(n583), .B(n584), .Z(n14700) );
  XOR U1398 ( .A(n15066), .B(n15067), .Z(n585) );
  NANDN U1399 ( .A(n15068), .B(n585), .Z(n586) );
  NAND U1400 ( .A(n15066), .B(n15067), .Z(n587) );
  AND U1401 ( .A(n586), .B(n587), .Z(n15325) );
  NAND U1402 ( .A(n15605), .B(n15606), .Z(n588) );
  XOR U1403 ( .A(n15605), .B(n15606), .Z(n589) );
  NANDN U1404 ( .A(n15604), .B(n589), .Z(n590) );
  NAND U1405 ( .A(n588), .B(n590), .Z(n15755) );
  NAND U1406 ( .A(n16151), .B(n16150), .Z(n591) );
  NAND U1407 ( .A(n16149), .B(n16148), .Z(n592) );
  AND U1408 ( .A(n591), .B(n592), .Z(n16463) );
  XNOR U1409 ( .A(n10959), .B(n10958), .Z(n10955) );
  XOR U1410 ( .A(n11466), .B(n11467), .Z(n593) );
  NANDN U1411 ( .A(n11468), .B(n593), .Z(n594) );
  NAND U1412 ( .A(n11466), .B(n11467), .Z(n595) );
  AND U1413 ( .A(n594), .B(n595), .Z(n11571) );
  NAND U1414 ( .A(n13036), .B(n13035), .Z(n596) );
  NAND U1415 ( .A(n13034), .B(n13033), .Z(n597) );
  AND U1416 ( .A(n596), .B(n597), .Z(n13199) );
  XOR U1417 ( .A(n8098), .B(n8097), .Z(n598) );
  NANDN U1418 ( .A(n8099), .B(n598), .Z(n599) );
  NAND U1419 ( .A(n8098), .B(n8097), .Z(n600) );
  AND U1420 ( .A(n599), .B(n600), .Z(n8154) );
  NAND U1421 ( .A(n9531), .B(n9532), .Z(n601) );
  XOR U1422 ( .A(n9531), .B(n9532), .Z(n602) );
  NANDN U1423 ( .A(n9530), .B(n602), .Z(n603) );
  NAND U1424 ( .A(n601), .B(n603), .Z(n9809) );
  XNOR U1425 ( .A(n10465), .B(n10464), .Z(n10462) );
  NAND U1426 ( .A(n5342), .B(n5343), .Z(n604) );
  XOR U1427 ( .A(n5342), .B(n5343), .Z(n605) );
  NANDN U1428 ( .A(n5341), .B(n605), .Z(n606) );
  NAND U1429 ( .A(n604), .B(n606), .Z(n5419) );
  XOR U1430 ( .A(n5589), .B(n5590), .Z(n607) );
  NANDN U1431 ( .A(n5591), .B(n607), .Z(n608) );
  NAND U1432 ( .A(n5589), .B(n5590), .Z(n609) );
  AND U1433 ( .A(n608), .B(n609), .Z(n5693) );
  XOR U1434 ( .A(n7011), .B(n7012), .Z(n610) );
  NANDN U1435 ( .A(n7013), .B(n610), .Z(n611) );
  NAND U1436 ( .A(n7011), .B(n7012), .Z(n612) );
  AND U1437 ( .A(n611), .B(n612), .Z(n7168) );
  XNOR U1438 ( .A(n7775), .B(n7774), .Z(n7518) );
  XOR U1439 ( .A(n2865), .B(n2866), .Z(n613) );
  NANDN U1440 ( .A(n2867), .B(n613), .Z(n614) );
  NAND U1441 ( .A(n2865), .B(n2866), .Z(n615) );
  AND U1442 ( .A(n614), .B(n615), .Z(n2977) );
  NAND U1443 ( .A(n3224), .B(n3225), .Z(n616) );
  XOR U1444 ( .A(n3224), .B(n3225), .Z(n617) );
  NANDN U1445 ( .A(n3223), .B(n617), .Z(n618) );
  NAND U1446 ( .A(n616), .B(n618), .Z(n3461) );
  NAND U1447 ( .A(n3744), .B(n3745), .Z(n619) );
  XOR U1448 ( .A(n3744), .B(n3745), .Z(n620) );
  NANDN U1449 ( .A(n3743), .B(n620), .Z(n621) );
  NAND U1450 ( .A(n619), .B(n621), .Z(n3893) );
  XNOR U1451 ( .A(n4855), .B(n4854), .Z(n4851) );
  XNOR U1452 ( .A(n44208), .B(n44207), .Z(n44209) );
  XNOR U1453 ( .A(n40558), .B(n40557), .Z(n40560) );
  XNOR U1454 ( .A(n40679), .B(n40678), .Z(n40681) );
  XNOR U1455 ( .A(n35716), .B(n35715), .Z(n35717) );
  XNOR U1456 ( .A(n29821), .B(n29820), .Z(n29822) );
  XNOR U1457 ( .A(n26812), .B(n26811), .Z(n26813) );
  XNOR U1458 ( .A(n23644), .B(n23643), .Z(n23645) );
  XNOR U1459 ( .A(n23933), .B(o[248]), .Z(n23948) );
  XNOR U1460 ( .A(n24130), .B(n24227), .Z(n23990) );
  XNOR U1461 ( .A(n21112), .B(n21111), .Z(n21113) );
  XNOR U1462 ( .A(n15722), .B(n15558), .Z(n15366) );
  XNOR U1463 ( .A(n15361), .B(n15360), .Z(n15371) );
  XNOR U1464 ( .A(n5842), .B(n5841), .Z(n5844) );
  XNOR U1465 ( .A(n5967), .B(n5966), .Z(n5969) );
  XNOR U1466 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U1467 ( .A(n46504), .B(n46503), .Z(n46524) );
  XNOR U1468 ( .A(n46713), .B(n46712), .Z(n46714) );
  XNOR U1469 ( .A(n43543), .B(n43542), .Z(n43530) );
  XNOR U1470 ( .A(n44054), .B(n44053), .Z(n44056) );
  XNOR U1471 ( .A(n44344), .B(n44343), .Z(n44346) );
  XNOR U1472 ( .A(n44524), .B(n44523), .Z(n44525) );
  XNOR U1473 ( .A(n40892), .B(n40891), .Z(n40893) );
  XNOR U1474 ( .A(n40917), .B(n40916), .Z(n40954) );
  XNOR U1475 ( .A(n37802), .B(n37801), .Z(n37783) );
  XNOR U1476 ( .A(n38059), .B(n38058), .Z(n38065) );
  XNOR U1477 ( .A(n34980), .B(n34979), .Z(n34961) );
  XNOR U1478 ( .A(n35828), .B(n35827), .Z(n35829) );
  XNOR U1479 ( .A(n35796), .B(n35795), .Z(n35798) );
  XNOR U1480 ( .A(n35877), .B(n35876), .Z(n35878) );
  XNOR U1481 ( .A(n32391), .B(n32390), .Z(n32393) );
  XNOR U1482 ( .A(n32608), .B(n32607), .Z(n32610) );
  XNOR U1483 ( .A(n32545), .B(n32544), .Z(n32613) );
  XNOR U1484 ( .A(n29115), .B(n29114), .Z(n29096) );
  XNOR U1485 ( .A(n29809), .B(n29808), .Z(n29749) );
  XNOR U1486 ( .A(n29924), .B(n29923), .Z(n29926) );
  XNOR U1487 ( .A(n30004), .B(n30003), .Z(n30005) );
  XNOR U1488 ( .A(n26149), .B(n26148), .Z(n26130) );
  XNOR U1489 ( .A(n22760), .B(o[238]), .Z(n22752) );
  XNOR U1490 ( .A(n23256), .B(n23255), .Z(n23237) );
  XNOR U1491 ( .A(n23691), .B(o[246]), .Z(n23670) );
  XNOR U1492 ( .A(n24132), .B(n24131), .Z(n24148) );
  XOR U1493 ( .A(n24138), .B(n24137), .Z(n24154) );
  XOR U1494 ( .A(n24127), .B(n24126), .Z(n24105) );
  XNOR U1495 ( .A(n24050), .B(n24049), .Z(n24051) );
  XNOR U1496 ( .A(n24118), .B(n24117), .Z(n24119) );
  XNOR U1497 ( .A(n24112), .B(n24111), .Z(n24113) );
  XNOR U1498 ( .A(n24284), .B(n24283), .Z(n24285) );
  XNOR U1499 ( .A(n24278), .B(n24277), .Z(n24279) );
  XNOR U1500 ( .A(n20583), .B(n20582), .Z(n20585) );
  XNOR U1501 ( .A(n20331), .B(n20330), .Z(n20333) );
  XOR U1502 ( .A(n20655), .B(n20654), .Z(n20671) );
  XNOR U1503 ( .A(n20705), .B(n20704), .Z(n20725) );
  XNOR U1504 ( .A(n21105), .B(n21106), .Z(n21077) );
  AND U1505 ( .A(n21279), .B(o[217]), .Z(n21412) );
  XNOR U1506 ( .A(n18065), .B(n18064), .Z(n18066) );
  XNOR U1507 ( .A(n18071), .B(n18070), .Z(n18072) );
  XNOR U1508 ( .A(n14414), .B(o[144]), .Z(n14428) );
  XNOR U1509 ( .A(n15013), .B(n15012), .Z(n15015) );
  XNOR U1510 ( .A(n14968), .B(n14967), .Z(n14969) );
  XNOR U1511 ( .A(n14974), .B(n14973), .Z(n14985) );
  XNOR U1512 ( .A(n15020), .B(n15019), .Z(n15046) );
  XNOR U1513 ( .A(n15395), .B(n15394), .Z(n15389) );
  XNOR U1514 ( .A(n15540), .B(n15539), .Z(n15542) );
  AND U1515 ( .A(n11117), .B(o[107]), .Z(n11195) );
  XNOR U1516 ( .A(n11537), .B(o[112]), .Z(n11552) );
  XNOR U1517 ( .A(n11738), .B(n11737), .Z(n11698) );
  XNOR U1518 ( .A(n11728), .B(n11727), .Z(n11745) );
  XNOR U1519 ( .A(n11716), .B(n11715), .Z(n11751) );
  XNOR U1520 ( .A(n11847), .B(n11846), .Z(n11848) );
  XNOR U1521 ( .A(n8926), .B(n8925), .Z(n8927) );
  XNOR U1522 ( .A(n9550), .B(n9549), .Z(n9546) );
  XNOR U1523 ( .A(n5659), .B(o[48]), .Z(n5674) );
  XNOR U1524 ( .A(n5850), .B(n5849), .Z(n5866) );
  XNOR U1525 ( .A(n5838), .B(n5837), .Z(n5873) );
  XNOR U1526 ( .A(n6774), .B(n6773), .Z(n6775) );
  XNOR U1527 ( .A(n46307), .B(n46306), .Z(n46309) );
  XNOR U1528 ( .A(n46170), .B(n46169), .Z(n46144) );
  XNOR U1529 ( .A(n47043), .B(n47042), .Z(n47044) );
  XNOR U1530 ( .A(n47051), .B(n47050), .Z(n47038) );
  XNOR U1531 ( .A(n47057), .B(n47056), .Z(n46994) );
  NAND U1532 ( .A(n47340), .B(n47341), .Z(n622) );
  NAND U1533 ( .A(n47338), .B(n47339), .Z(n623) );
  NAND U1534 ( .A(n622), .B(n623), .Z(n47504) );
  AND U1535 ( .A(n47623), .B(o[507]), .Z(n47712) );
  XOR U1536 ( .A(n47639), .B(n47638), .Z(n47649) );
  XNOR U1537 ( .A(n42922), .B(n42921), .Z(n42915) );
  XNOR U1538 ( .A(n43597), .B(n43596), .Z(n43599) );
  XNOR U1539 ( .A(n44239), .B(n44238), .Z(n44240) );
  XNOR U1540 ( .A(n44599), .B(n44598), .Z(n44600) );
  XNOR U1541 ( .A(n44726), .B(n44725), .Z(n44727) );
  XNOR U1542 ( .A(n44732), .B(n44731), .Z(n44734) );
  XNOR U1543 ( .A(n44841), .B(n44840), .Z(n44842) );
  NAND U1544 ( .A(n40355), .B(n40354), .Z(n624) );
  NANDN U1545 ( .A(n41158), .B(n40552), .Z(n625) );
  NAND U1546 ( .A(n624), .B(n625), .Z(n40460) );
  XNOR U1547 ( .A(n40668), .B(n40667), .Z(n40707) );
  XNOR U1548 ( .A(n40714), .B(n40713), .Z(n40716) );
  XNOR U1549 ( .A(n40751), .B(n40750), .Z(n40753) );
  XNOR U1550 ( .A(n41198), .B(n41197), .Z(n41191) );
  XNOR U1551 ( .A(n41220), .B(n41219), .Z(n41183) );
  XNOR U1552 ( .A(n41352), .B(n41351), .Z(n41353) );
  NAND U1553 ( .A(n41448), .B(n41449), .Z(n626) );
  NANDN U1554 ( .A(n41451), .B(n41450), .Z(n627) );
  AND U1555 ( .A(n626), .B(n627), .Z(n41668) );
  XNOR U1556 ( .A(n37855), .B(n37854), .Z(n37857) );
  XNOR U1557 ( .A(n37984), .B(n37983), .Z(n37934) );
  XNOR U1558 ( .A(n38469), .B(n38468), .Z(n38419) );
  XNOR U1559 ( .A(n38780), .B(n38779), .Z(n38773) );
  XNOR U1560 ( .A(n34351), .B(n34350), .Z(n34344) );
  NAND U1561 ( .A(n34426), .B(n34425), .Z(n628) );
  NANDN U1562 ( .A(n34988), .B(n34424), .Z(n629) );
  NAND U1563 ( .A(n628), .B(n629), .Z(n34530) );
  XNOR U1564 ( .A(n34609), .B(n34608), .Z(n34611) );
  NAND U1565 ( .A(n34889), .B(n34888), .Z(n630) );
  NANDN U1566 ( .A(n36093), .B(n34887), .Z(n631) );
  NAND U1567 ( .A(n630), .B(n631), .Z(n35003) );
  XNOR U1568 ( .A(n35544), .B(n35543), .Z(n35545) );
  XNOR U1569 ( .A(n35564), .B(n35563), .Z(n35501) );
  XNOR U1570 ( .A(n35704), .B(n35703), .Z(n35706) );
  XNOR U1571 ( .A(n35836), .B(n35835), .Z(n35807) );
  XNOR U1572 ( .A(n35985), .B(n35984), .Z(n35987) );
  XNOR U1573 ( .A(n35914), .B(n35913), .Z(n35915) );
  NAND U1574 ( .A(n35928), .B(n35927), .Z(n632) );
  NAND U1575 ( .A(n35925), .B(n35926), .Z(n633) );
  NAND U1576 ( .A(n632), .B(n633), .Z(n36113) );
  NAND U1577 ( .A(n35936), .B(n35937), .Z(n634) );
  NAND U1578 ( .A(n36139), .B(n35935), .Z(n635) );
  NAND U1579 ( .A(n634), .B(n635), .Z(n36082) );
  NAND U1580 ( .A(n31424), .B(n31423), .Z(n636) );
  NANDN U1581 ( .A(n31851), .B(n31477), .Z(n637) );
  NAND U1582 ( .A(n636), .B(n637), .Z(n31473) );
  XOR U1583 ( .A(n31651), .B(n31650), .Z(n31631) );
  XNOR U1584 ( .A(n32036), .B(n32035), .Z(n32074) );
  XNOR U1585 ( .A(n32459), .B(n32458), .Z(n32409) );
  XNOR U1586 ( .A(n32431), .B(n32430), .Z(n32475) );
  XNOR U1587 ( .A(n32469), .B(n32468), .Z(n32471) );
  XNOR U1588 ( .A(n28326), .B(o[298]), .Z(n28337) );
  XNOR U1589 ( .A(n28478), .B(n28477), .Z(n28479) );
  XNOR U1590 ( .A(n28494), .B(n29108), .Z(n28473) );
  NAND U1591 ( .A(n28924), .B(n28925), .Z(n638) );
  NAND U1592 ( .A(n29007), .B(n29912), .Z(n639) );
  NAND U1593 ( .A(n638), .B(n639), .Z(n29061) );
  XNOR U1594 ( .A(n29290), .B(n29289), .Z(n29240) );
  XNOR U1595 ( .A(n29664), .B(n29663), .Z(n29665) );
  XNOR U1596 ( .A(n29684), .B(n29683), .Z(n29621) );
  XNOR U1597 ( .A(n29827), .B(n29826), .Z(n29829) );
  XNOR U1598 ( .A(n30054), .B(n30055), .Z(n30034) );
  XNOR U1599 ( .A(n30071), .B(n30070), .Z(n30073) );
  XNOR U1600 ( .A(n30777), .B(n30592), .Z(n30593) );
  NAND U1601 ( .A(n25993), .B(n25994), .Z(n640) );
  NANDN U1602 ( .A(n25996), .B(n25995), .Z(n641) );
  AND U1603 ( .A(n640), .B(n641), .Z(n26041) );
  AND U1604 ( .A(n26049), .B(n26048), .Z(n642) );
  AND U1605 ( .A(n26047), .B(x[486]), .Z(n643) );
  NAND U1606 ( .A(y[7949]), .B(n643), .Z(n644) );
  NANDN U1607 ( .A(n642), .B(n644), .Z(n26214) );
  NAND U1608 ( .A(n26090), .B(n26091), .Z(n645) );
  NAND U1609 ( .A(n26088), .B(n26089), .Z(n646) );
  NAND U1610 ( .A(n645), .B(n646), .Z(n26202) );
  XNOR U1611 ( .A(n27192), .B(n27191), .Z(n27194) );
  XNOR U1612 ( .A(n27206), .B(n27205), .Z(n27207) );
  XNOR U1613 ( .A(n27202), .B(n27201), .Z(n27124) );
  XNOR U1614 ( .A(n27180), .B(n27179), .Z(n27181) );
  XNOR U1615 ( .A(n27218), .B(n27217), .Z(n27219) );
  XOR U1616 ( .A(n22602), .B(n22603), .Z(n22587) );
  XNOR U1617 ( .A(n22965), .B(n22964), .Z(n22967) );
  XNOR U1618 ( .A(n23959), .B(n23958), .Z(n23960) );
  XNOR U1619 ( .A(n23942), .B(n23943), .Z(n23935) );
  XNOR U1620 ( .A(n24304), .B(n24303), .Z(n24249) );
  XNOR U1621 ( .A(n24544), .B(n24543), .Z(n24545) );
  XNOR U1622 ( .A(n19698), .B(n19697), .Z(n19672) );
  NAND U1623 ( .A(n19822), .B(n19821), .Z(n647) );
  NANDN U1624 ( .A(n20241), .B(n19863), .Z(n648) );
  NAND U1625 ( .A(n647), .B(n648), .Z(n19859) );
  XOR U1626 ( .A(n20045), .B(n20044), .Z(n20025) );
  XNOR U1627 ( .A(n20154), .B(n20153), .Z(n20137) );
  XNOR U1628 ( .A(n20230), .B(n20229), .Z(n20235) );
  XNOR U1629 ( .A(n20589), .B(n20588), .Z(n20591) );
  XNOR U1630 ( .A(n20406), .B(n20405), .Z(n20453) );
  XNOR U1631 ( .A(n20552), .B(n20551), .Z(n20554) );
  XNOR U1632 ( .A(n20778), .B(n20777), .Z(n20780) );
  XNOR U1633 ( .A(n20985), .B(n20984), .Z(n20986) );
  XNOR U1634 ( .A(n20993), .B(n20992), .Z(n20930) );
  NAND U1635 ( .A(n21277), .B(n21278), .Z(n649) );
  NAND U1636 ( .A(n21275), .B(n21276), .Z(n650) );
  NAND U1637 ( .A(n649), .B(n650), .Z(n21320) );
  NAND U1638 ( .A(n21419), .B(n21420), .Z(n651) );
  NAND U1639 ( .A(n21556), .B(n21418), .Z(n652) );
  NAND U1640 ( .A(n651), .B(n652), .Z(n21487) );
  XNOR U1641 ( .A(n17086), .B(n17085), .Z(n17058) );
  NAND U1642 ( .A(n17268), .B(n17269), .Z(n653) );
  NAND U1643 ( .A(n17266), .B(n17267), .Z(n654) );
  NAND U1644 ( .A(n653), .B(n654), .Z(n17366) );
  NAND U1645 ( .A(n17265), .B(n17264), .Z(n655) );
  NANDN U1646 ( .A(n18015), .B(n17446), .Z(n656) );
  NAND U1647 ( .A(n655), .B(n656), .Z(n17369) );
  XOR U1648 ( .A(n17604), .B(n17603), .Z(n17621) );
  XNOR U1649 ( .A(n17614), .B(n17613), .Z(n17616) );
  NAND U1650 ( .A(n17925), .B(n17926), .Z(n657) );
  NAND U1651 ( .A(n17923), .B(n17924), .Z(n658) );
  NAND U1652 ( .A(n657), .B(n658), .Z(n18040) );
  NAND U1653 ( .A(n14278), .B(n14277), .Z(n659) );
  NAND U1654 ( .A(n14320), .B(n15946), .Z(n660) );
  AND U1655 ( .A(n659), .B(n660), .Z(n14348) );
  XNOR U1656 ( .A(n15164), .B(n15163), .Z(n15166) );
  XNOR U1657 ( .A(n15286), .B(n15285), .Z(n15273) );
  XNOR U1658 ( .A(n15292), .B(n15291), .Z(n15229) );
  XNOR U1659 ( .A(n15379), .B(n15378), .Z(n15436) );
  XNOR U1660 ( .A(n15705), .B(n15704), .Z(n15706) );
  XNOR U1661 ( .A(n15699), .B(n15698), .Z(n15700) );
  XNOR U1662 ( .A(n15642), .B(n15643), .Z(n15625) );
  NAND U1663 ( .A(n11198), .B(n11199), .Z(n661) );
  NAND U1664 ( .A(n11395), .B(n12507), .Z(n662) );
  NAND U1665 ( .A(n661), .B(n662), .Z(n11257) );
  XNOR U1666 ( .A(n11414), .B(n11413), .Z(n11443) );
  XNOR U1667 ( .A(n11506), .B(n11505), .Z(n11495) );
  XNOR U1668 ( .A(n11489), .B(n11488), .Z(n11491) );
  XNOR U1669 ( .A(n11651), .B(n11650), .Z(n11653) );
  XNOR U1670 ( .A(n11520), .B(n11519), .Z(n11521) );
  XOR U1671 ( .A(n11843), .B(n11842), .Z(n11885) );
  XNOR U1672 ( .A(n11810), .B(n11809), .Z(n11890) );
  XNOR U1673 ( .A(n11916), .B(n11915), .Z(n11918) );
  XNOR U1674 ( .A(n12491), .B(n12490), .Z(n12492) );
  NAND U1675 ( .A(n12620), .B(n12619), .Z(n663) );
  NAND U1676 ( .A(n12618), .B(n12617), .Z(n664) );
  AND U1677 ( .A(n663), .B(n664), .Z(n12794) );
  NAND U1678 ( .A(n12699), .B(n12700), .Z(n665) );
  NAND U1679 ( .A(n12697), .B(n12698), .Z(n666) );
  NAND U1680 ( .A(n665), .B(n666), .Z(n12867) );
  XNOR U1681 ( .A(n8193), .B(o[75]), .Z(n8173) );
  XNOR U1682 ( .A(n8267), .B(n8900), .Z(n8247) );
  XNOR U1683 ( .A(n8237), .B(n8236), .Z(n8230) );
  XNOR U1684 ( .A(n9051), .B(n9050), .Z(n9053) );
  XNOR U1685 ( .A(n9150), .B(n9149), .Z(n9152) );
  XNOR U1686 ( .A(n9739), .B(n9738), .Z(n9710) );
  XNOR U1687 ( .A(n5020), .B(o[39]), .Z(n5015) );
  XNOR U1688 ( .A(n5179), .B(n5178), .Z(n5153) );
  XNOR U1689 ( .A(n5531), .B(n5530), .Z(n5560) );
  XNOR U1690 ( .A(n5546), .B(n5545), .Z(n5547) );
  XNOR U1691 ( .A(n5628), .B(n5627), .Z(n5618) );
  XNOR U1692 ( .A(n5612), .B(n5611), .Z(n5614) );
  XNOR U1693 ( .A(n5773), .B(n5772), .Z(n5775) );
  XNOR U1694 ( .A(n5642), .B(n5641), .Z(n5643) );
  XOR U1695 ( .A(n5997), .B(n5996), .Z(n6007) );
  XNOR U1696 ( .A(n5932), .B(n5931), .Z(n6012) );
  XNOR U1697 ( .A(n6038), .B(n6037), .Z(n6040) );
  XNOR U1698 ( .A(n6946), .B(n6945), .Z(n6947) );
  XNOR U1699 ( .A(n6910), .B(n6909), .Z(n6912) );
  NAND U1700 ( .A(n6743), .B(n6744), .Z(n667) );
  NANDN U1701 ( .A(n6746), .B(n6745), .Z(n668) );
  AND U1702 ( .A(n667), .B(n668), .Z(n6959) );
  XNOR U1703 ( .A(n7075), .B(n7074), .Z(n7076) );
  XNOR U1704 ( .A(n7081), .B(n7080), .Z(n7083) );
  XNOR U1705 ( .A(n2116), .B(o[8]), .Z(n2111) );
  XNOR U1706 ( .A(n2367), .B(o[12]), .Z(n2386) );
  NAND U1707 ( .A(n2843), .B(n2844), .Z(n669) );
  NANDN U1708 ( .A(n2846), .B(n2845), .Z(n670) );
  AND U1709 ( .A(n669), .B(n670), .Z(n2887) );
  NAND U1710 ( .A(n2929), .B(n2930), .Z(n671) );
  NAND U1711 ( .A(n2927), .B(n2928), .Z(n672) );
  NAND U1712 ( .A(n671), .B(n672), .Z(n3015) );
  XNOR U1713 ( .A(n3060), .B(n3059), .Z(n3008) );
  XNOR U1714 ( .A(n3122), .B(n3121), .Z(n3123) );
  XNOR U1715 ( .A(n3134), .B(n3133), .Z(n3136) );
  XNOR U1716 ( .A(n3171), .B(n3170), .Z(n3173) );
  XNOR U1717 ( .A(n3660), .B(n3659), .Z(n3661) );
  XNOR U1718 ( .A(n3942), .B(n3941), .Z(n3923) );
  XNOR U1719 ( .A(n47353), .B(n47352), .Z(n47354) );
  XNOR U1720 ( .A(n47645), .B(n47644), .Z(n47657) );
  NAND U1721 ( .A(n47279), .B(n47280), .Z(n673) );
  NANDN U1722 ( .A(n47282), .B(n47281), .Z(n674) );
  NAND U1723 ( .A(n673), .B(n674), .Z(n47386) );
  NAND U1724 ( .A(n47278), .B(n47277), .Z(n675) );
  NAND U1725 ( .A(n47276), .B(n47275), .Z(n676) );
  AND U1726 ( .A(n675), .B(n676), .Z(n47509) );
  NAND U1727 ( .A(n47598), .B(n47599), .Z(n677) );
  NANDN U1728 ( .A(n47601), .B(n47600), .Z(n678) );
  AND U1729 ( .A(n677), .B(n678), .Z(n47781) );
  XNOR U1730 ( .A(n47727), .B(n47726), .Z(n47816) );
  XOR U1731 ( .A(n47978), .B(n47977), .Z(n47979) );
  NAND U1732 ( .A(n43148), .B(n43149), .Z(n679) );
  NAND U1733 ( .A(n43961), .B(n43541), .Z(n680) );
  NAND U1734 ( .A(n679), .B(n680), .Z(n43259) );
  XNOR U1735 ( .A(n43428), .B(n43427), .Z(n43429) );
  XOR U1736 ( .A(n43611), .B(n43610), .Z(n43519) );
  XOR U1737 ( .A(n43617), .B(n43616), .Z(n43621) );
  XNOR U1738 ( .A(n43744), .B(n43743), .Z(n43745) );
  XNOR U1739 ( .A(n44320), .B(n44319), .Z(n44322) );
  XNOR U1740 ( .A(n44436), .B(n44435), .Z(n44437) );
  XNOR U1741 ( .A(n44846), .B(n44847), .Z(n44919) );
  XNOR U1742 ( .A(n44802), .B(n44801), .Z(n44908) );
  XNOR U1743 ( .A(n40031), .B(n40032), .Z(n40017) );
  XNOR U1744 ( .A(n40787), .B(n40786), .Z(n40845) );
  XNOR U1745 ( .A(n40858), .B(n40857), .Z(n40859) );
  XNOR U1746 ( .A(n40880), .B(n40879), .Z(n40881) );
  XNOR U1747 ( .A(n41358), .B(n41357), .Z(n41360) );
  XNOR U1748 ( .A(n41292), .B(n41291), .Z(n41293) );
  OR U1749 ( .A(n41470), .B(n41471), .Z(n681) );
  NAND U1750 ( .A(n41468), .B(n41469), .Z(n682) );
  NAND U1751 ( .A(n681), .B(n682), .Z(n41589) );
  NAND U1752 ( .A(n41467), .B(n41466), .Z(n683) );
  NAND U1753 ( .A(n41465), .B(n41464), .Z(n684) );
  AND U1754 ( .A(n683), .B(n684), .Z(n41712) );
  NAND U1755 ( .A(n41787), .B(n41786), .Z(n685) );
  NANDN U1756 ( .A(n41785), .B(n41784), .Z(n686) );
  AND U1757 ( .A(n685), .B(n686), .Z(n41984) );
  XOR U1758 ( .A(n37195), .B(n37196), .Z(n37180) );
  NAND U1759 ( .A(n37607), .B(n37608), .Z(n687) );
  NAND U1760 ( .A(n37605), .B(n37606), .Z(n688) );
  NAND U1761 ( .A(n687), .B(n688), .Z(n37763) );
  XNOR U1762 ( .A(n37748), .B(n37747), .Z(n37756) );
  XOR U1763 ( .A(n37869), .B(n37868), .Z(n37778) );
  XNOR U1764 ( .A(n38532), .B(n38531), .Z(n38533) );
  XNOR U1765 ( .A(n38963), .B(n38962), .Z(n38905) );
  XNOR U1766 ( .A(n39006), .B(n39005), .Z(n39008) );
  NAND U1767 ( .A(n39073), .B(n39074), .Z(n689) );
  NAND U1768 ( .A(n39075), .B(n39076), .Z(n690) );
  NAND U1769 ( .A(n689), .B(n690), .Z(n39284) );
  XNOR U1770 ( .A(n39501), .B(n39500), .Z(n39499) );
  NAND U1771 ( .A(n39300), .B(n39301), .Z(n691) );
  NAND U1772 ( .A(n39298), .B(n39299), .Z(n692) );
  NAND U1773 ( .A(n691), .B(n692), .Z(n39461) );
  NAND U1774 ( .A(n38982), .B(n38983), .Z(n693) );
  NAND U1775 ( .A(n38980), .B(n38981), .Z(n694) );
  NAND U1776 ( .A(n693), .B(n694), .Z(n39050) );
  XNOR U1777 ( .A(n36634), .B(n36633), .Z(n36631) );
  NAND U1778 ( .A(n36119), .B(n36120), .Z(n695) );
  NAND U1779 ( .A(n36117), .B(n36118), .Z(n696) );
  NAND U1780 ( .A(n695), .B(n696), .Z(n36276) );
  XNOR U1781 ( .A(n31075), .B(o[325]), .Z(n31062) );
  XNOR U1782 ( .A(n31309), .B(n31308), .Z(n31310) );
  XNOR U1783 ( .A(n31454), .B(n31453), .Z(n31456) );
  NAND U1784 ( .A(n31497), .B(n31496), .Z(n697) );
  NANDN U1785 ( .A(n31616), .B(n32034), .Z(n698) );
  NAND U1786 ( .A(n697), .B(n698), .Z(n31536) );
  NAND U1787 ( .A(n31486), .B(n31485), .Z(n699) );
  NAND U1788 ( .A(n31484), .B(n31483), .Z(n700) );
  AND U1789 ( .A(n699), .B(n700), .Z(n31528) );
  NAND U1790 ( .A(n31577), .B(n31576), .Z(n701) );
  NAND U1791 ( .A(n31575), .B(n31574), .Z(n702) );
  AND U1792 ( .A(n701), .B(n702), .Z(n31672) );
  NAND U1793 ( .A(n31540), .B(n31541), .Z(n703) );
  NAND U1794 ( .A(n31538), .B(n31539), .Z(n704) );
  NAND U1795 ( .A(n703), .B(n704), .Z(n31658) );
  XOR U1796 ( .A(n31780), .B(n31779), .Z(n31782) );
  XNOR U1797 ( .A(n32127), .B(n32126), .Z(n32129) );
  XOR U1798 ( .A(n32483), .B(n32482), .Z(n32486) );
  XNOR U1799 ( .A(n32795), .B(n32794), .Z(n32797) );
  XNOR U1800 ( .A(n33704), .B(n33545), .Z(n33546) );
  XNOR U1801 ( .A(n33499), .B(n33498), .Z(n33500) );
  XOR U1802 ( .A(n33242), .B(n33241), .Z(n33252) );
  XOR U1803 ( .A(n28200), .B(n29019), .Z(n28202) );
  XNOR U1804 ( .A(n29401), .B(n29400), .Z(n29403) );
  XNOR U1805 ( .A(n30200), .B(n30199), .Z(n30202) );
  XNOR U1806 ( .A(n30414), .B(n30413), .Z(n30444) );
  XNOR U1807 ( .A(n30366), .B(n30365), .Z(n30367) );
  XOR U1808 ( .A(n25539), .B(n25540), .Z(n25524) );
  XNOR U1809 ( .A(n25835), .B(n25834), .Z(n25836) );
  XNOR U1810 ( .A(n26097), .B(n26096), .Z(n26098) );
  XNOR U1811 ( .A(n26109), .B(n26108), .Z(n26111) );
  XNOR U1812 ( .A(n26115), .B(n26114), .Z(n26117) );
  XNOR U1813 ( .A(n26784), .B(n26783), .Z(n26785) );
  XNOR U1814 ( .A(n27043), .B(n27042), .Z(n27046) );
  XOR U1815 ( .A(n27361), .B(n27360), .Z(n27371) );
  XNOR U1816 ( .A(n27479), .B(n27478), .Z(n27481) );
  XNOR U1817 ( .A(n27790), .B(n27646), .Z(n27647) );
  XNOR U1818 ( .A(n27264), .B(n27263), .Z(n27365) );
  XNOR U1819 ( .A(n22889), .B(n22888), .Z(n22890) );
  XNOR U1820 ( .A(n23115), .B(n23114), .Z(n23117) );
  XNOR U1821 ( .A(n23335), .B(n23334), .Z(n23338) );
  XNOR U1822 ( .A(n23965), .B(n23964), .Z(n23967) );
  XOR U1823 ( .A(n24088), .B(n24087), .Z(n24046) );
  XNOR U1824 ( .A(n24144), .B(n24143), .Z(n24160) );
  XNOR U1825 ( .A(n24242), .B(n24241), .Z(n24244) );
  XNOR U1826 ( .A(n24538), .B(n24537), .Z(n24539) );
  XNOR U1827 ( .A(n24726), .B(n24725), .Z(n24780) );
  XNOR U1828 ( .A(n19763), .B(n19762), .Z(n19764) );
  NAND U1829 ( .A(n19883), .B(n19882), .Z(n705) );
  NANDN U1830 ( .A(n20010), .B(n20418), .Z(n706) );
  NAND U1831 ( .A(n705), .B(n706), .Z(n19931) );
  NAND U1832 ( .A(n19872), .B(n19871), .Z(n707) );
  NAND U1833 ( .A(n19870), .B(n19869), .Z(n708) );
  AND U1834 ( .A(n707), .B(n708), .Z(n19923) );
  NAND U1835 ( .A(n19975), .B(n19974), .Z(n709) );
  NAND U1836 ( .A(n19973), .B(n19972), .Z(n710) );
  AND U1837 ( .A(n709), .B(n710), .Z(n20066) );
  NAND U1838 ( .A(n19935), .B(n19936), .Z(n711) );
  NAND U1839 ( .A(n19933), .B(n19934), .Z(n712) );
  NAND U1840 ( .A(n711), .B(n712), .Z(n20052) );
  XNOR U1841 ( .A(n20158), .B(n20157), .Z(n20170) );
  XOR U1842 ( .A(n20126), .B(n20125), .Z(n20128) );
  XNOR U1843 ( .A(n20224), .B(n20223), .Z(n20274) );
  XNOR U1844 ( .A(n20380), .B(n20379), .Z(n20382) );
  XNOR U1845 ( .A(n20395), .B(n20394), .Z(n20478) );
  XNOR U1846 ( .A(n20472), .B(n20471), .Z(n20473) );
  XOR U1847 ( .A(n20526), .B(n20525), .Z(n20518) );
  NAND U1848 ( .A(n21643), .B(n21642), .Z(n713) );
  NAND U1849 ( .A(n21640), .B(n21641), .Z(n714) );
  NAND U1850 ( .A(n713), .B(n714), .Z(n21853) );
  NAND U1851 ( .A(n21552), .B(n21553), .Z(n715) );
  NAND U1852 ( .A(n21550), .B(n21551), .Z(n716) );
  NAND U1853 ( .A(n715), .B(n716), .Z(n21621) );
  XNOR U1854 ( .A(n16808), .B(n16807), .Z(n16809) );
  XNOR U1855 ( .A(n17021), .B(n17020), .Z(n17023) );
  XNOR U1856 ( .A(n17207), .B(n17206), .Z(n17208) );
  XNOR U1857 ( .A(n17423), .B(n17422), .Z(n17425) );
  NAND U1858 ( .A(n17363), .B(n17362), .Z(n717) );
  NAND U1859 ( .A(n17361), .B(n17360), .Z(n718) );
  AND U1860 ( .A(n717), .B(n718), .Z(n17489) );
  XOR U1861 ( .A(n17628), .B(n17627), .Z(n17536) );
  XNOR U1862 ( .A(n17683), .B(n17682), .Z(n17685) );
  NAND U1863 ( .A(n17889), .B(n17890), .Z(n719) );
  NANDN U1864 ( .A(n17892), .B(n17891), .Z(n720) );
  NAND U1865 ( .A(n719), .B(n720), .Z(n18102) );
  XOR U1866 ( .A(n18239), .B(n18238), .Z(n18133) );
  XNOR U1867 ( .A(n18654), .B(n18653), .Z(n18720) );
  XOR U1868 ( .A(n18704), .B(n18703), .Z(n18714) );
  XNOR U1869 ( .A(n18832), .B(n18831), .Z(n18834) );
  XNOR U1870 ( .A(n19139), .B(n18995), .Z(n18996) );
  XNOR U1871 ( .A(n14113), .B(n14114), .Z(n14099) );
  XOR U1872 ( .A(n14788), .B(n14787), .Z(n14782) );
  NAND U1873 ( .A(n14903), .B(n14904), .Z(n721) );
  NANDN U1874 ( .A(n14906), .B(n14905), .Z(n722) );
  NAND U1875 ( .A(n721), .B(n722), .Z(n14955) );
  XNOR U1876 ( .A(n15296), .B(n15295), .Z(n15297) );
  XNOR U1877 ( .A(n15482), .B(n15481), .Z(n15484) );
  XNOR U1878 ( .A(n15595), .B(n15594), .Z(n15586) );
  XNOR U1879 ( .A(n15617), .B(n15616), .Z(n15742) );
  NAND U1880 ( .A(n15622), .B(n15623), .Z(n723) );
  NAND U1881 ( .A(n15620), .B(n15621), .Z(n724) );
  NAND U1882 ( .A(n723), .B(n724), .Z(n15871) );
  XOR U1883 ( .A(n15759), .B(n15758), .Z(n15761) );
  XNOR U1884 ( .A(n15765), .B(n15764), .Z(n15767) );
  NAND U1885 ( .A(n15804), .B(n15805), .Z(n725) );
  NAND U1886 ( .A(n15802), .B(n15803), .Z(n726) );
  NAND U1887 ( .A(n725), .B(n726), .Z(n15975) );
  NAND U1888 ( .A(n15801), .B(n15800), .Z(n727) );
  NANDN U1889 ( .A(n15799), .B(n15798), .Z(n728) );
  NAND U1890 ( .A(n727), .B(n728), .Z(n15972) );
  NAND U1891 ( .A(n15813), .B(n15814), .Z(n729) );
  NAND U1892 ( .A(n15811), .B(n15812), .Z(n730) );
  NAND U1893 ( .A(n729), .B(n730), .Z(n15917) );
  NAND U1894 ( .A(n15941), .B(n15942), .Z(n731) );
  NAND U1895 ( .A(n15939), .B(n15940), .Z(n732) );
  NAND U1896 ( .A(n731), .B(n732), .Z(n16176) );
  NAND U1897 ( .A(n15923), .B(n15924), .Z(n733) );
  NAND U1898 ( .A(n15921), .B(n15922), .Z(n734) );
  NAND U1899 ( .A(n733), .B(n734), .Z(n16180) );
  NAND U1900 ( .A(n16187), .B(n16186), .Z(n735) );
  NAND U1901 ( .A(n16184), .B(n16185), .Z(n736) );
  AND U1902 ( .A(n735), .B(n736), .Z(n16358) );
  XNOR U1903 ( .A(n10863), .B(o[102]), .Z(n10855) );
  XNOR U1904 ( .A(n11136), .B(n11135), .Z(n11137) );
  NAND U1905 ( .A(n11276), .B(n11275), .Z(n737) );
  NAND U1906 ( .A(n11274), .B(n11273), .Z(n738) );
  AND U1907 ( .A(n737), .B(n738), .Z(n11307) );
  XNOR U1908 ( .A(n11461), .B(n11460), .Z(n11462) );
  XNOR U1909 ( .A(n11685), .B(n11684), .Z(n11687) );
  XNOR U1910 ( .A(n11899), .B(n11898), .Z(n11911) );
  XOR U1911 ( .A(n12301), .B(n12300), .Z(n12192) );
  NAND U1912 ( .A(n12642), .B(n12641), .Z(n739) );
  NAND U1913 ( .A(n12640), .B(n12639), .Z(n740) );
  AND U1914 ( .A(n739), .B(n740), .Z(n12823) );
  NAND U1915 ( .A(n12643), .B(n12644), .Z(n741) );
  NANDN U1916 ( .A(n12646), .B(n12645), .Z(n742) );
  NAND U1917 ( .A(n741), .B(n742), .Z(n12743) );
  NAND U1918 ( .A(n12914), .B(n12915), .Z(n743) );
  NAND U1919 ( .A(n12912), .B(n12913), .Z(n744) );
  NAND U1920 ( .A(n743), .B(n744), .Z(n13133) );
  XOR U1921 ( .A(n13335), .B(n13334), .Z(n13337) );
  XNOR U1922 ( .A(n7935), .B(o[70]), .Z(n7927) );
  XNOR U1923 ( .A(n8147), .B(n8146), .Z(n8148) );
  XNOR U1924 ( .A(n8305), .B(n8304), .Z(n8292) );
  XNOR U1925 ( .A(n8329), .B(n8328), .Z(n8297) );
  XNOR U1926 ( .A(n8967), .B(n8966), .Z(n8968) );
  XNOR U1927 ( .A(n8987), .B(n8986), .Z(n8990) );
  XNOR U1928 ( .A(n9045), .B(n9044), .Z(n9047) );
  XNOR U1929 ( .A(n9834), .B(n9833), .Z(n9836) );
  XOR U1930 ( .A(n10225), .B(n10224), .Z(n10227) );
  NAND U1931 ( .A(n10083), .B(n10082), .Z(n745) );
  NANDN U1932 ( .A(n10081), .B(n10080), .Z(n746) );
  NAND U1933 ( .A(n745), .B(n746), .Z(n10270) );
  XNOR U1934 ( .A(n5109), .B(o[41]), .Z(n5099) );
  XNOR U1935 ( .A(n5257), .B(n5256), .Z(n5258) );
  XNOR U1936 ( .A(n5291), .B(n5290), .Z(n5284) );
  XNOR U1937 ( .A(n5584), .B(n5583), .Z(n5585) );
  XNOR U1938 ( .A(n5807), .B(n5806), .Z(n5809) );
  XNOR U1939 ( .A(n6046), .B(n6045), .Z(n6132) );
  XNOR U1940 ( .A(n6021), .B(n6020), .Z(n6033) );
  XNOR U1941 ( .A(n6258), .B(n6257), .Z(n6170) );
  XNOR U1942 ( .A(n7232), .B(n7231), .Z(n7233) );
  XNOR U1943 ( .A(n7453), .B(n7452), .Z(n7477) );
  XNOR U1944 ( .A(n2076), .B(o[7]), .Z(n2071) );
  XOR U1945 ( .A(n2124), .B(n2918), .Z(n2126) );
  XOR U1946 ( .A(n2204), .B(n2203), .Z(n2192) );
  XOR U1947 ( .A(n2320), .B(n2319), .Z(n2322) );
  XNOR U1948 ( .A(n2372), .B(n2373), .Z(n2358) );
  XNOR U1949 ( .A(n2667), .B(n2666), .Z(n2669) );
  XNOR U1950 ( .A(n2663), .B(n2662), .Z(n2655) );
  NAND U1951 ( .A(n2836), .B(n2837), .Z(n747) );
  NAND U1952 ( .A(n2906), .B(n3778), .Z(n748) );
  NAND U1953 ( .A(n747), .B(n748), .Z(n2958) );
  AND U1954 ( .A(n2897), .B(n2896), .Z(n749) );
  AND U1955 ( .A(n3268), .B(y[7687]), .Z(n750) );
  NAND U1956 ( .A(x[496]), .B(n750), .Z(n751) );
  NANDN U1957 ( .A(n749), .B(n751), .Z(n2993) );
  XNOR U1958 ( .A(n3883), .B(n3882), .Z(n3886) );
  NAND U1959 ( .A(n4176), .B(n4175), .Z(n752) );
  NANDN U1960 ( .A(n4174), .B(n4173), .Z(n753) );
  NAND U1961 ( .A(n752), .B(n753), .Z(n4322) );
  XOR U1962 ( .A(n4263), .B(n4262), .Z(n4367) );
  XNOR U1963 ( .A(n4213), .B(n4212), .Z(n4214) );
  XNOR U1964 ( .A(n45542), .B(n45541), .Z(n45543) );
  XNOR U1965 ( .A(n47105), .B(n47104), .Z(n47106) );
  XNOR U1966 ( .A(n47101), .B(n47100), .Z(n47220) );
  XOR U1967 ( .A(n47236), .B(n47235), .Z(n47229) );
  XOR U1968 ( .A(n47825), .B(n47824), .Z(n47830) );
  NAND U1969 ( .A(n48095), .B(n48096), .Z(n754) );
  NAND U1970 ( .A(n48107), .B(n48097), .Z(n755) );
  AND U1971 ( .A(n754), .B(n755), .Z(n756) );
  NAND U1972 ( .A(n48098), .B(n48099), .Z(n757) );
  NAND U1973 ( .A(n48100), .B(n48101), .Z(n758) );
  AND U1974 ( .A(n757), .B(n758), .Z(n759) );
  NAND U1975 ( .A(n48102), .B(n48103), .Z(n760) );
  NAND U1976 ( .A(n48127), .B(n48104), .Z(n761) );
  AND U1977 ( .A(n760), .B(n761), .Z(n762) );
  XOR U1978 ( .A(n48147), .B(n48146), .Z(n763) );
  XNOR U1979 ( .A(n48141), .B(n48140), .Z(n764) );
  XNOR U1980 ( .A(n763), .B(n764), .Z(n765) );
  AND U1981 ( .A(x[484]), .B(y[8187]), .Z(n766) );
  XNOR U1982 ( .A(n48112), .B(n48111), .Z(n767) );
  XNOR U1983 ( .A(n766), .B(n767), .Z(n768) );
  XOR U1984 ( .A(n765), .B(n768), .Z(n769) );
  XNOR U1985 ( .A(n759), .B(n762), .Z(n770) );
  XNOR U1986 ( .A(n769), .B(n770), .Z(n771) );
  XNOR U1987 ( .A(n756), .B(n771), .Z(n48148) );
  XNOR U1988 ( .A(n48039), .B(n48038), .Z(n48040) );
  XNOR U1989 ( .A(n47956), .B(n47955), .Z(n47957) );
  XNOR U1990 ( .A(n42654), .B(n42653), .Z(n42661) );
  NAND U1991 ( .A(n43263), .B(n43264), .Z(n772) );
  NANDN U1992 ( .A(n43266), .B(n43265), .Z(n773) );
  NAND U1993 ( .A(n772), .B(n773), .Z(n43308) );
  XNOR U1994 ( .A(n44023), .B(n44022), .Z(n44024) );
  XNOR U1995 ( .A(n44464), .B(n44463), .Z(n44465) );
  XOR U1996 ( .A(n44778), .B(n44777), .Z(n44772) );
  XOR U1997 ( .A(n44915), .B(n44914), .Z(n44891) );
  NAND U1998 ( .A(n44678), .B(n44679), .Z(n774) );
  NANDN U1999 ( .A(n44681), .B(n44680), .Z(n775) );
  AND U2000 ( .A(n774), .B(n775), .Z(n44885) );
  XNOR U2001 ( .A(n45052), .B(n45051), .Z(n45053) );
  NAND U2002 ( .A(n45174), .B(n45175), .Z(n776) );
  NANDN U2003 ( .A(n45176), .B(n45200), .Z(n777) );
  AND U2004 ( .A(n776), .B(n777), .Z(n45226) );
  XOR U2005 ( .A(n45269), .B(n45270), .Z(n45271) );
  XNOR U2006 ( .A(n45148), .B(n45147), .Z(n45145) );
  NAND U2007 ( .A(n39966), .B(n39965), .Z(n778) );
  NAND U2008 ( .A(n40930), .B(n39964), .Z(n779) );
  NAND U2009 ( .A(n778), .B(n779), .Z(n40003) );
  XNOR U2010 ( .A(n40226), .B(n40225), .Z(n40228) );
  XOR U2011 ( .A(n40979), .B(n40978), .Z(n40874) );
  XNOR U2012 ( .A(n41018), .B(n41017), .Z(n41002) );
  XNOR U2013 ( .A(n41280), .B(n41279), .Z(n41281) );
  XNOR U2014 ( .A(n42132), .B(n42131), .Z(n42133) );
  XNOR U2015 ( .A(n42378), .B(n42379), .Z(n42376) );
  NAND U2016 ( .A(n37754), .B(n37753), .Z(n780) );
  NAND U2017 ( .A(n37752), .B(n37751), .Z(n781) );
  AND U2018 ( .A(n780), .B(n781), .Z(n37876) );
  NAND U2019 ( .A(n37762), .B(n37761), .Z(n782) );
  NAND U2020 ( .A(n37759), .B(n37760), .Z(n783) );
  NAND U2021 ( .A(n782), .B(n783), .Z(n37872) );
  XNOR U2022 ( .A(n38149), .B(n38148), .Z(n38142) );
  XNOR U2023 ( .A(n39014), .B(n39013), .Z(n38892) );
  XNOR U2024 ( .A(n39126), .B(n39125), .Z(n39128) );
  NAND U2025 ( .A(n39095), .B(n39096), .Z(n784) );
  NAND U2026 ( .A(n39093), .B(n39094), .Z(n785) );
  NAND U2027 ( .A(n784), .B(n785), .Z(n39218) );
  XNOR U2028 ( .A(n39116), .B(n39115), .Z(n39036) );
  NAND U2029 ( .A(n39251), .B(n39250), .Z(n786) );
  NAND U2030 ( .A(n39248), .B(n39249), .Z(n787) );
  NAND U2031 ( .A(n786), .B(n787), .Z(n39343) );
  NAND U2032 ( .A(n39080), .B(n39079), .Z(n788) );
  NAND U2033 ( .A(n39077), .B(n39078), .Z(n789) );
  NAND U2034 ( .A(n788), .B(n789), .Z(n39203) );
  XNOR U2035 ( .A(n34073), .B(n34072), .Z(n34080) );
  XNOR U2036 ( .A(n35059), .B(n35058), .Z(n35062) );
  XNOR U2037 ( .A(n36171), .B(n36170), .Z(n36050) );
  XNOR U2038 ( .A(n36284), .B(n36283), .Z(n36200) );
  NAND U2039 ( .A(n36148), .B(n36149), .Z(n790) );
  NANDN U2040 ( .A(n36151), .B(n36150), .Z(n791) );
  NAND U2041 ( .A(n790), .B(n791), .Z(n36196) );
  NAND U2042 ( .A(n36302), .B(n36301), .Z(n792) );
  NAND U2043 ( .A(n36299), .B(n36300), .Z(n793) );
  NAND U2044 ( .A(n792), .B(n793), .Z(n36441) );
  NAND U2045 ( .A(n36273), .B(n36274), .Z(n794) );
  NAND U2046 ( .A(n36271), .B(n36272), .Z(n795) );
  NAND U2047 ( .A(n794), .B(n795), .Z(n36444) );
  NAND U2048 ( .A(n36535), .B(n36474), .Z(n796) );
  XOR U2049 ( .A(n36535), .B(n36474), .Z(n797) );
  NANDN U2050 ( .A(n36473), .B(n797), .Z(n798) );
  NAND U2051 ( .A(n796), .B(n798), .Z(n36674) );
  NAND U2052 ( .A(n36611), .B(n36612), .Z(n799) );
  NAND U2053 ( .A(n36614), .B(n36613), .Z(n800) );
  AND U2054 ( .A(n799), .B(n800), .Z(n801) );
  NAND U2055 ( .A(n36615), .B(n36616), .Z(n802) );
  NAND U2056 ( .A(n36617), .B(n36618), .Z(n803) );
  AND U2057 ( .A(n802), .B(n803), .Z(n804) );
  AND U2058 ( .A(y[8033]), .B(x[510]), .Z(n805) );
  NAND U2059 ( .A(y[8034]), .B(x[509]), .Z(n806) );
  XNOR U2060 ( .A(n805), .B(n806), .Z(n807) );
  AND U2061 ( .A(y[8054]), .B(x[489]), .Z(n808) );
  NAND U2062 ( .A(x[494]), .B(y[8049]), .Z(n809) );
  XNOR U2063 ( .A(n808), .B(n809), .Z(n810) );
  XOR U2064 ( .A(n36622), .B(n36621), .Z(n811) );
  XNOR U2065 ( .A(n36620), .B(n36619), .Z(n812) );
  XNOR U2066 ( .A(n811), .B(n812), .Z(n813) );
  XOR U2067 ( .A(n810), .B(n813), .Z(n814) );
  XNOR U2068 ( .A(n804), .B(n807), .Z(n815) );
  XNOR U2069 ( .A(n814), .B(n815), .Z(n816) );
  XNOR U2070 ( .A(n801), .B(n816), .Z(n36623) );
  XNOR U2071 ( .A(n36524), .B(n36523), .Z(n36521) );
  XOR U2072 ( .A(n32244), .B(n32243), .Z(n32246) );
  XNOR U2073 ( .A(n32387), .B(n32386), .Z(n32378) );
  XOR U2074 ( .A(n32622), .B(n32621), .Z(n32508) );
  XNOR U2075 ( .A(n33266), .B(n33265), .Z(n33125) );
  XNOR U2076 ( .A(n33572), .B(n33571), .Z(n33574) );
  XNOR U2077 ( .A(n33394), .B(n33393), .Z(n33288) );
  XNOR U2078 ( .A(n33586), .B(n33585), .Z(n33562) );
  XOR U2079 ( .A(n33590), .B(n33589), .Z(n33591) );
  XNOR U2080 ( .A(n33846), .B(n33845), .Z(n33844) );
  XNOR U2081 ( .A(n33660), .B(n33659), .Z(n33657) );
  NAND U2082 ( .A(n28294), .B(n28293), .Z(n817) );
  NANDN U2083 ( .A(n28926), .B(n28633), .Z(n818) );
  AND U2084 ( .A(n817), .B(n818), .Z(n28297) );
  XOR U2085 ( .A(n30483), .B(n30482), .Z(n30457) );
  NAND U2086 ( .A(n30262), .B(n30263), .Z(n819) );
  NANDN U2087 ( .A(n30265), .B(n30264), .Z(n820) );
  AND U2088 ( .A(n819), .B(n820), .Z(n30451) );
  XOR U2089 ( .A(n30427), .B(n30426), .Z(n30469) );
  XOR U2090 ( .A(n30656), .B(n30655), .Z(n30658) );
  XNOR U2091 ( .A(n30638), .B(n30637), .Z(n30639) );
  XNOR U2092 ( .A(n30907), .B(n30906), .Z(n30905) );
  XNOR U2093 ( .A(n25589), .B(n25588), .Z(n25576) );
  XNOR U2094 ( .A(n27686), .B(n27685), .Z(n27687) );
  XNOR U2095 ( .A(n27692), .B(n27691), .Z(n27694) );
  XOR U2096 ( .A(n27761), .B(n27760), .Z(n27759) );
  XNOR U2097 ( .A(n27767), .B(n27766), .Z(n27764) );
  XNOR U2098 ( .A(n27513), .B(n27512), .Z(n27407) );
  NAND U2099 ( .A(n23156), .B(n22366), .Z(n821) );
  NANDN U2100 ( .A(n22368), .B(n22367), .Z(n822) );
  NAND U2101 ( .A(n821), .B(n822), .Z(n22387) );
  XNOR U2102 ( .A(n22991), .B(n22990), .Z(n22960) );
  XOR U2103 ( .A(n22879), .B(n22878), .Z(n22870) );
  XNOR U2104 ( .A(n23109), .B(n23108), .Z(n23110) );
  XOR U2105 ( .A(n23013), .B(n23012), .Z(n23102) );
  XNOR U2106 ( .A(n24194), .B(n24193), .Z(n24328) );
  XNOR U2107 ( .A(n24473), .B(n24472), .Z(n24344) );
  XNOR U2108 ( .A(n24498), .B(n24497), .Z(n24491) );
  XOR U2109 ( .A(n24576), .B(n24575), .Z(n24617) );
  XNOR U2110 ( .A(n24502), .B(n24501), .Z(n24503) );
  XNOR U2111 ( .A(n24775), .B(n24774), .Z(n24777) );
  XNOR U2112 ( .A(n25018), .B(n25017), .Z(n25015) );
  XOR U2113 ( .A(n24854), .B(n24853), .Z(n24852) );
  XNOR U2114 ( .A(n24769), .B(n24768), .Z(n24770) );
  XNOR U2115 ( .A(n19487), .B(n19486), .Z(n19479) );
  NAND U2116 ( .A(n20337), .B(n19570), .Z(n823) );
  NANDN U2117 ( .A(n19572), .B(n19571), .Z(n824) );
  NAND U2118 ( .A(n823), .B(n824), .Z(n19600) );
  XOR U2119 ( .A(n19716), .B(n19715), .Z(n19746) );
  XNOR U2120 ( .A(n20296), .B(n20295), .Z(n20298) );
  XNOR U2121 ( .A(n20613), .B(n20612), .Z(n20615) );
  XNOR U2122 ( .A(n20734), .B(n20733), .Z(n20640) );
  XNOR U2123 ( .A(n20768), .B(n20767), .Z(n20762) );
  XNOR U2124 ( .A(n21011), .B(n21010), .Z(n20890) );
  XNOR U2125 ( .A(n21155), .B(n21154), .Z(n21156) );
  XNOR U2126 ( .A(n21459), .B(n21458), .Z(n21460) );
  XNOR U2127 ( .A(n21465), .B(n21464), .Z(n21467) );
  NAND U2128 ( .A(n21557), .B(n21558), .Z(n825) );
  NANDN U2129 ( .A(n21560), .B(n21559), .Z(n826) );
  NAND U2130 ( .A(n825), .B(n826), .Z(n21605) );
  NAND U2131 ( .A(n22044), .B(n22043), .Z(n827) );
  NAND U2132 ( .A(n22042), .B(n22041), .Z(n828) );
  AND U2133 ( .A(n827), .B(n828), .Z(n22052) );
  XNOR U2134 ( .A(n21922), .B(n21921), .Z(n21919) );
  NAND U2135 ( .A(n21617), .B(n21618), .Z(n829) );
  NAND U2136 ( .A(n21615), .B(n21616), .Z(n830) );
  NAND U2137 ( .A(n829), .B(n830), .Z(n21746) );
  XNOR U2138 ( .A(n17215), .B(n17214), .Z(n17195) );
  NAND U2139 ( .A(n17398), .B(n17399), .Z(n831) );
  NAND U2140 ( .A(n17396), .B(n17397), .Z(n832) );
  NAND U2141 ( .A(n831), .B(n832), .Z(n17414) );
  XOR U2142 ( .A(n17640), .B(n17639), .Z(n17632) );
  XOR U2143 ( .A(n17768), .B(n17767), .Z(n17770) );
  NAND U2144 ( .A(n17978), .B(n17977), .Z(n833) );
  NANDN U2145 ( .A(n17976), .B(n17975), .Z(n834) );
  AND U2146 ( .A(n833), .B(n834), .Z(n17993) );
  XNOR U2147 ( .A(n17880), .B(n17879), .Z(n17881) );
  NAND U2148 ( .A(n18112), .B(n18113), .Z(n835) );
  NAND U2149 ( .A(n18110), .B(n18111), .Z(n836) );
  NAND U2150 ( .A(n835), .B(n836), .Z(n18255) );
  XNOR U2151 ( .A(n18277), .B(n18276), .Z(n18279) );
  XNOR U2152 ( .A(n18271), .B(n18270), .Z(n18272) );
  XNOR U2153 ( .A(n18728), .B(n18727), .Z(n18587) );
  XNOR U2154 ( .A(n19034), .B(n19033), .Z(n19035) );
  XOR U2155 ( .A(n19040), .B(n19039), .Z(n19042) );
  XNOR U2156 ( .A(n19131), .B(n19130), .Z(n19128) );
  XOR U2157 ( .A(n19117), .B(n19116), .Z(n19115) );
  XNOR U2158 ( .A(n18866), .B(n18865), .Z(n18759) );
  XNOR U2159 ( .A(n14237), .B(n14236), .Z(n14239) );
  XNOR U2160 ( .A(n14800), .B(n14799), .Z(n14803) );
  XNOR U2161 ( .A(n15189), .B(n15188), .Z(n15190) );
  NAND U2162 ( .A(n15822), .B(n15821), .Z(n837) );
  NANDN U2163 ( .A(n15820), .B(n15819), .Z(n838) );
  AND U2164 ( .A(n837), .B(n838), .Z(n15980) );
  NAND U2165 ( .A(n15865), .B(n15866), .Z(n839) );
  NANDN U2166 ( .A(n15868), .B(n15867), .Z(n840) );
  NAND U2167 ( .A(n839), .B(n840), .Z(n16011) );
  NAND U2168 ( .A(n16147), .B(n16146), .Z(n841) );
  NAND U2169 ( .A(n16145), .B(n16331), .Z(n842) );
  NAND U2170 ( .A(n841), .B(n842), .Z(n16237) );
  NAND U2171 ( .A(n15949), .B(n15950), .Z(n843) );
  NAND U2172 ( .A(n15947), .B(n15948), .Z(n844) );
  NAND U2173 ( .A(n843), .B(n844), .Z(n16111) );
  XNOR U2174 ( .A(n10948), .B(n10947), .Z(n10949) );
  XNOR U2175 ( .A(n11451), .B(n11450), .Z(n11387) );
  XNOR U2176 ( .A(n11679), .B(n11678), .Z(n11680) );
  XOR U2177 ( .A(n11577), .B(n11576), .Z(n11672) );
  XNOR U2178 ( .A(n12319), .B(n12318), .Z(n12320) );
  XOR U2179 ( .A(n13016), .B(n13015), .Z(n12873) );
  XOR U2180 ( .A(n13329), .B(n13328), .Z(n13331) );
  XNOR U2181 ( .A(n13150), .B(n13149), .Z(n13151) );
  XNOR U2182 ( .A(n13264), .B(n13263), .Z(n13232) );
  XNOR U2183 ( .A(n13349), .B(n13348), .Z(n13313) );
  XNOR U2184 ( .A(n13612), .B(n13611), .Z(n13609) );
  XOR U2185 ( .A(n13420), .B(n13419), .Z(n13418) );
  XOR U2186 ( .A(n13188), .B(n13187), .Z(n13041) );
  XNOR U2187 ( .A(n7920), .B(n7919), .Z(n7912) );
  XNOR U2188 ( .A(n7958), .B(n7957), .Z(n7976) );
  XNOR U2189 ( .A(n9112), .B(n9111), .Z(n9114) );
  XNOR U2190 ( .A(n9237), .B(n9236), .Z(n9144) );
  XNOR U2191 ( .A(n9254), .B(n9253), .Z(n9256) );
  XNOR U2192 ( .A(n9983), .B(n9982), .Z(n9985) );
  XOR U2193 ( .A(n10152), .B(n10151), .Z(n10138) );
  NAND U2194 ( .A(n10055), .B(n10056), .Z(n845) );
  NANDN U2195 ( .A(n10058), .B(n10057), .Z(n846) );
  AND U2196 ( .A(n845), .B(n846), .Z(n10251) );
  XNOR U2197 ( .A(n10412), .B(n10411), .Z(n10413) );
  XNOR U2198 ( .A(n5114), .B(n5113), .Z(n5087) );
  XOR U2199 ( .A(n5210), .B(n5209), .Z(n5240) );
  XOR U2200 ( .A(n5574), .B(n5573), .Z(n5565) );
  XNOR U2201 ( .A(n5801), .B(n5800), .Z(n5802) );
  XOR U2202 ( .A(n5699), .B(n5698), .Z(n5794) );
  XOR U2203 ( .A(n6179), .B(n6178), .Z(n6165) );
  XOR U2204 ( .A(n7320), .B(n7319), .Z(n7294) );
  NAND U2205 ( .A(n7090), .B(n7091), .Z(n847) );
  NANDN U2206 ( .A(n7093), .B(n7092), .Z(n848) );
  AND U2207 ( .A(n847), .B(n848), .Z(n7288) );
  XOR U2208 ( .A(n7264), .B(n7263), .Z(n7306) );
  XNOR U2209 ( .A(n7312), .B(n7311), .Z(n7314) );
  XNOR U2210 ( .A(n7375), .B(n7374), .Z(n7376) );
  XNOR U2211 ( .A(n7741), .B(n7740), .Z(n7739) );
  XNOR U2212 ( .A(n2030), .B(n2029), .Z(n2032) );
  XOR U2213 ( .A(n2078), .B(n2007), .Z(n849) );
  NANDN U2214 ( .A(n2008), .B(n849), .Z(n850) );
  NAND U2215 ( .A(n2078), .B(n2007), .Z(n851) );
  AND U2216 ( .A(n850), .B(n851), .Z(n2056) );
  XNOR U2217 ( .A(n2209), .B(n2208), .Z(n2210) );
  XNOR U2218 ( .A(n2217), .B(n2216), .Z(n2269) );
  XNOR U2219 ( .A(n2460), .B(n2459), .Z(n2494) );
  XNOR U2220 ( .A(n2435), .B(n2434), .Z(n2489) );
  XOR U2221 ( .A(n2862), .B(n2861), .Z(n2783) );
  XNOR U2222 ( .A(n2876), .B(n2875), .Z(n2877) );
  OR U2223 ( .A(n3005), .B(n3006), .Z(n852) );
  NAND U2224 ( .A(n3004), .B(n3003), .Z(n853) );
  AND U2225 ( .A(n852), .B(n853), .Z(n3201) );
  XNOR U2226 ( .A(n3233), .B(n3232), .Z(n3235) );
  XNOR U2227 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U2228 ( .A(n4203), .B(n4202), .Z(n4077) );
  XNOR U2229 ( .A(n4086), .B(n4085), .Z(n4072) );
  XNOR U2230 ( .A(n4435), .B(n4434), .Z(n4394) );
  XOR U2231 ( .A(n4589), .B(n4588), .Z(n4587) );
  XNOR U2232 ( .A(n4609), .B(n4608), .Z(n4606) );
  XNOR U2233 ( .A(n45483), .B(n45482), .Z(n45485) );
  XNOR U2234 ( .A(n45717), .B(n45716), .Z(n45719) );
  XNOR U2235 ( .A(n45940), .B(n45939), .Z(n45942) );
  XNOR U2236 ( .A(n46337), .B(n46336), .Z(n46436) );
  NAND U2237 ( .A(n47964), .B(n47963), .Z(n854) );
  NAND U2238 ( .A(n47962), .B(n47961), .Z(n855) );
  AND U2239 ( .A(n854), .B(n855), .Z(n48222) );
  NAND U2240 ( .A(n42568), .B(n42567), .Z(n856) );
  XOR U2241 ( .A(n42568), .B(n42567), .Z(n857) );
  NANDN U2242 ( .A(n42640), .B(n857), .Z(n858) );
  NAND U2243 ( .A(n856), .B(n858), .Z(n42613) );
  XNOR U2244 ( .A(n42823), .B(n42822), .Z(n42825) );
  XNOR U2245 ( .A(n45060), .B(n45059), .Z(n44953) );
  NAND U2246 ( .A(n44904), .B(n44905), .Z(n859) );
  NAND U2247 ( .A(n44902), .B(n44903), .Z(n860) );
  NAND U2248 ( .A(n859), .B(n860), .Z(n44960) );
  XOR U2249 ( .A(n45354), .B(n45353), .Z(n45352) );
  NAND U2250 ( .A(n45315), .B(n45316), .Z(n45320) );
  XNOR U2251 ( .A(n39800), .B(n39799), .Z(n39801) );
  XOR U2252 ( .A(n40746), .B(n40745), .Z(n40633) );
  XNOR U2253 ( .A(n41553), .B(n41552), .Z(n41554) );
  XNOR U2254 ( .A(n42096), .B(n42095), .Z(n42058) );
  XOR U2255 ( .A(n37078), .B(n37077), .Z(n37080) );
  XNOR U2256 ( .A(n37676), .B(n37675), .Z(n37770) );
  XNOR U2257 ( .A(n38134), .B(n38133), .Z(n38136) );
  XNOR U2258 ( .A(n38704), .B(n38703), .Z(n38706) );
  NAND U2259 ( .A(n39269), .B(n39270), .Z(n861) );
  NANDN U2260 ( .A(n39272), .B(n39271), .Z(n862) );
  NAND U2261 ( .A(n861), .B(n862), .Z(n39546) );
  XOR U2262 ( .A(n39529), .B(n39528), .Z(n39527) );
  NAND U2263 ( .A(n33986), .B(n33985), .Z(n863) );
  XOR U2264 ( .A(n33986), .B(n33985), .Z(n864) );
  NANDN U2265 ( .A(n34059), .B(n864), .Z(n865) );
  NAND U2266 ( .A(n863), .B(n865), .Z(n34031) );
  XNOR U2267 ( .A(n34244), .B(n34243), .Z(n34246) );
  XNOR U2268 ( .A(n34465), .B(n34464), .Z(n34467) );
  XOR U2269 ( .A(n34756), .B(n34755), .Z(n34845) );
  XNOR U2270 ( .A(n35606), .B(n35605), .Z(n35607) );
  XNOR U2271 ( .A(n36436), .B(n36435), .Z(n36358) );
  NAND U2272 ( .A(n36447), .B(n36448), .Z(n866) );
  NANDN U2273 ( .A(n36450), .B(n36449), .Z(n867) );
  AND U2274 ( .A(n866), .B(n867), .Z(n36689) );
  NAND U2275 ( .A(n36265), .B(n36266), .Z(n868) );
  NAND U2276 ( .A(n36263), .B(n36264), .Z(n869) );
  NAND U2277 ( .A(n868), .B(n869), .Z(n36386) );
  NAND U2278 ( .A(n30986), .B(n30985), .Z(n870) );
  NAND U2279 ( .A(n30984), .B(n30993), .Z(n871) );
  AND U2280 ( .A(n870), .B(n871), .Z(n30999) );
  XOR U2281 ( .A(n31195), .B(n31194), .Z(n31197) );
  XNOR U2282 ( .A(n31447), .B(n31446), .Z(n31449) );
  XNOR U2283 ( .A(n31787), .B(n31786), .Z(n31789) );
  XNOR U2284 ( .A(n32648), .B(n32647), .Z(n32649) );
  XOR U2285 ( .A(n33475), .B(n33474), .Z(n33477) );
  XNOR U2286 ( .A(n33870), .B(n33869), .Z(n33868) );
  NAND U2287 ( .A(n28084), .B(n28083), .Z(n872) );
  NANDN U2288 ( .A(n28169), .B(n28161), .Z(n873) );
  NAND U2289 ( .A(n872), .B(n873), .Z(n28097) );
  XOR U2290 ( .A(n28223), .B(n28222), .Z(n28240) );
  XNOR U2291 ( .A(n28247), .B(n28246), .Z(n28248) );
  XNOR U2292 ( .A(n28579), .B(n28578), .Z(n28581) );
  XNOR U2293 ( .A(n28588), .B(n28587), .Z(n28669) );
  XNOR U2294 ( .A(n29712), .B(n29711), .Z(n29713) );
  XNOR U2295 ( .A(n30627), .B(n30626), .Z(n30534) );
  XNOR U2296 ( .A(n30652), .B(n30651), .Z(n30542) );
  XNOR U2297 ( .A(n30695), .B(n30694), .Z(n30931) );
  XNOR U2298 ( .A(n26023), .B(n26022), .Z(n26025) );
  XNOR U2299 ( .A(n26356), .B(n26355), .Z(n26357) );
  NAND U2300 ( .A(n26484), .B(n26485), .Z(n874) );
  NANDN U2301 ( .A(n26487), .B(n26486), .Z(n875) );
  AND U2302 ( .A(n874), .B(n875), .Z(n26615) );
  XNOR U2303 ( .A(n27067), .B(n27066), .Z(n27069) );
  XOR U2304 ( .A(n28003), .B(n28002), .Z(n28001) );
  XOR U2305 ( .A(n27717), .B(n27715), .Z(n876) );
  NANDN U2306 ( .A(n27716), .B(n876), .Z(n877) );
  NAND U2307 ( .A(n27717), .B(n27715), .Z(n878) );
  AND U2308 ( .A(n877), .B(n878), .Z(n27748) );
  XNOR U2309 ( .A(n22252), .B(n22251), .Z(n22253) );
  XNOR U2310 ( .A(n22806), .B(n22805), .Z(n22807) );
  XNOR U2311 ( .A(n23877), .B(n23876), .Z(n23878) );
  XNOR U2312 ( .A(n24759), .B(n24758), .Z(n24659) );
  NAND U2313 ( .A(n24509), .B(n24508), .Z(n879) );
  XOR U2314 ( .A(n24509), .B(n24508), .Z(n880) );
  NANDN U2315 ( .A(n24507), .B(n880), .Z(n881) );
  NAND U2316 ( .A(n879), .B(n881), .Z(n24653) );
  XOR U2317 ( .A(n25060), .B(n25059), .Z(n25058) );
  XOR U2318 ( .A(n24982), .B(n24981), .Z(n882) );
  XNOR U2319 ( .A(n24968), .B(n24967), .Z(n883) );
  XNOR U2320 ( .A(n882), .B(n883), .Z(n884) );
  XOR U2321 ( .A(n25010), .B(n25009), .Z(n885) );
  XNOR U2322 ( .A(n24996), .B(n24995), .Z(n886) );
  XNOR U2323 ( .A(n885), .B(n886), .Z(n887) );
  XOR U2324 ( .A(n884), .B(n887), .Z(n888) );
  NAND U2325 ( .A(n24860), .B(n24859), .Z(n889) );
  NAND U2326 ( .A(n24861), .B(n24862), .Z(n890) );
  AND U2327 ( .A(n889), .B(n890), .Z(n891) );
  XOR U2328 ( .A(n24930), .B(n24929), .Z(n892) );
  XNOR U2329 ( .A(n24874), .B(n24873), .Z(n893) );
  XNOR U2330 ( .A(n892), .B(n893), .Z(n894) );
  XNOR U2331 ( .A(n891), .B(n894), .Z(n895) );
  XNOR U2332 ( .A(n888), .B(n895), .Z(n896) );
  NAND U2333 ( .A(n24855), .B(n24856), .Z(n897) );
  NAND U2334 ( .A(n24857), .B(n24858), .Z(n898) );
  NAND U2335 ( .A(n897), .B(n898), .Z(n899) );
  XNOR U2336 ( .A(n896), .B(n899), .Z(n25011) );
  XNOR U2337 ( .A(n19542), .B(n19541), .Z(n19546) );
  XNOR U2338 ( .A(n20177), .B(n20176), .Z(n20179) );
  XNOR U2339 ( .A(n20625), .B(n20624), .Z(n20626) );
  XNOR U2340 ( .A(n21033), .B(n21032), .Z(n21160) );
  NAND U2341 ( .A(n21837), .B(n21836), .Z(n900) );
  NAND U2342 ( .A(n21835), .B(n21834), .Z(n901) );
  AND U2343 ( .A(n900), .B(n901), .Z(n22130) );
  NAND U2344 ( .A(n21838), .B(n21839), .Z(n902) );
  NANDN U2345 ( .A(n21841), .B(n21840), .Z(n903) );
  NAND U2346 ( .A(n902), .B(n903), .Z(n22123) );
  XNOR U2347 ( .A(n22106), .B(n22105), .Z(n22103) );
  NAND U2348 ( .A(n21745), .B(n21744), .Z(n904) );
  NAND U2349 ( .A(n21743), .B(n21742), .Z(n905) );
  AND U2350 ( .A(n904), .B(n905), .Z(n22148) );
  XOR U2351 ( .A(n16959), .B(n16958), .Z(n16961) );
  XNOR U2352 ( .A(n17235), .B(n17234), .Z(n17312) );
  XNOR U2353 ( .A(n17759), .B(n17758), .Z(n17761) );
  XNOR U2354 ( .A(n18732), .B(n18731), .Z(n18733) );
  XOR U2355 ( .A(n19353), .B(n19352), .Z(n19351) );
  XOR U2356 ( .A(n19329), .B(n19328), .Z(n19327) );
  XOR U2357 ( .A(n19105), .B(n19104), .Z(n19103) );
  NAND U2358 ( .A(n13901), .B(n13902), .Z(n906) );
  NANDN U2359 ( .A(n13904), .B(n13903), .Z(n907) );
  AND U2360 ( .A(n906), .B(n907), .Z(n14002) );
  NAND U2361 ( .A(n14394), .B(n14395), .Z(n908) );
  NAND U2362 ( .A(n14392), .B(n14393), .Z(n909) );
  NAND U2363 ( .A(n908), .B(n909), .Z(n14585) );
  XOR U2364 ( .A(n15332), .B(n15331), .Z(n15463) );
  NAND U2365 ( .A(n15916), .B(n15915), .Z(n910) );
  NANDN U2366 ( .A(n15914), .B(n15913), .Z(n911) );
  AND U2367 ( .A(n910), .B(n911), .Z(n16068) );
  NAND U2368 ( .A(n16002), .B(n16001), .Z(n912) );
  NAND U2369 ( .A(n15999), .B(n16000), .Z(n913) );
  NAND U2370 ( .A(n912), .B(n913), .Z(n16150) );
  XNOR U2371 ( .A(n16206), .B(n16205), .Z(n16203) );
  XNOR U2372 ( .A(n10957), .B(n10956), .Z(n10958) );
  XOR U2373 ( .A(n10979), .B(n10978), .Z(n10965) );
  XNOR U2374 ( .A(n12019), .B(n12018), .Z(n12038) );
  XNOR U2375 ( .A(n12720), .B(n12719), .Z(n12722) );
  XNOR U2376 ( .A(n13630), .B(n13629), .Z(n13628) );
  XNOR U2377 ( .A(n13210), .B(n13209), .Z(n13202) );
  XNOR U2378 ( .A(n7906), .B(n7905), .Z(n7907) );
  XOR U2379 ( .A(n8044), .B(n8043), .Z(n8083) );
  XNOR U2380 ( .A(n8284), .B(n8283), .Z(n8286) );
  XNOR U2381 ( .A(n8374), .B(n8373), .Z(n8455) );
  XNOR U2382 ( .A(n8766), .B(n8765), .Z(n8865) );
  XNOR U2383 ( .A(n9515), .B(n9514), .Z(n9516) );
  XNOR U2384 ( .A(n9813), .B(n9812), .Z(n9815) );
  NAND U2385 ( .A(n10164), .B(n10163), .Z(n914) );
  NANDN U2386 ( .A(n10162), .B(n10161), .Z(n915) );
  AND U2387 ( .A(n914), .B(n915), .Z(n10309) );
  XNOR U2388 ( .A(n4951), .B(n4950), .Z(n4952) );
  XNOR U2389 ( .A(n6141), .B(n6140), .Z(n6160) );
  XNOR U2390 ( .A(n7175), .B(n7174), .Z(n7334) );
  XNOR U2391 ( .A(n7468), .B(n7467), .Z(n7362) );
  XNOR U2392 ( .A(n7460), .B(n7459), .Z(n7461) );
  XNOR U2393 ( .A(n7529), .B(n7528), .Z(n7765) );
  NAND U2394 ( .A(n1943), .B(n1942), .Z(n916) );
  NAND U2395 ( .A(n1941), .B(n1950), .Z(n917) );
  AND U2396 ( .A(n916), .B(n917), .Z(n1956) );
  XNOR U2397 ( .A(n2156), .B(n2155), .Z(n2158) );
  XNOR U2398 ( .A(n2768), .B(n2767), .Z(n2770) );
  XNOR U2399 ( .A(n3603), .B(n3602), .Z(n3604) );
  XNOR U2400 ( .A(n3903), .B(n3902), .Z(n3905) );
  XNOR U2401 ( .A(n4408), .B(n4407), .Z(n4532) );
  XNOR U2402 ( .A(n4839), .B(n4838), .Z(n4836) );
  XNOR U2403 ( .A(n4810), .B(n4811), .Z(n4812) );
  NAND U2404 ( .A(n4247), .B(n4246), .Z(n918) );
  NANDN U2405 ( .A(n4245), .B(n4244), .Z(n919) );
  NAND U2406 ( .A(n918), .B(n919), .Z(n4389) );
  NAND U2407 ( .A(n45479), .B(n45480), .Z(n920) );
  XOR U2408 ( .A(n45479), .B(n45480), .Z(n921) );
  NANDN U2409 ( .A(n45478), .B(n921), .Z(n922) );
  NAND U2410 ( .A(n920), .B(n922), .Z(n45489) );
  NAND U2411 ( .A(n45658), .B(n45659), .Z(n923) );
  XOR U2412 ( .A(n45658), .B(n45659), .Z(n924) );
  NANDN U2413 ( .A(n45657), .B(n924), .Z(n925) );
  NAND U2414 ( .A(n923), .B(n925), .Z(n45713) );
  XOR U2415 ( .A(n46324), .B(n46325), .Z(n926) );
  NANDN U2416 ( .A(n46326), .B(n926), .Z(n927) );
  NAND U2417 ( .A(n46324), .B(n46325), .Z(n928) );
  AND U2418 ( .A(n927), .B(n928), .Z(n46443) );
  NAND U2419 ( .A(n46944), .B(n46945), .Z(n929) );
  XOR U2420 ( .A(n46944), .B(n46945), .Z(n930) );
  NAND U2421 ( .A(n930), .B(n46943), .Z(n931) );
  NAND U2422 ( .A(n929), .B(n931), .Z(n47085) );
  XOR U2423 ( .A(n47666), .B(n47667), .Z(n932) );
  NANDN U2424 ( .A(n47668), .B(n932), .Z(n933) );
  NAND U2425 ( .A(n47666), .B(n47667), .Z(n934) );
  AND U2426 ( .A(n933), .B(n934), .Z(n47681) );
  NAND U2427 ( .A(n47679), .B(n47678), .Z(n935) );
  NAND U2428 ( .A(n47677), .B(n47676), .Z(n936) );
  AND U2429 ( .A(n935), .B(n936), .Z(n47836) );
  NAND U2430 ( .A(n48243), .B(n48242), .Z(n937) );
  NAND U2431 ( .A(n48241), .B(n48240), .Z(n938) );
  AND U2432 ( .A(n937), .B(n938), .Z(n48251) );
  XOR U2433 ( .A(n42579), .B(n42580), .Z(n939) );
  NANDN U2434 ( .A(n42581), .B(n939), .Z(n940) );
  NAND U2435 ( .A(n42579), .B(n42580), .Z(n941) );
  AND U2436 ( .A(n940), .B(n941), .Z(n42620) );
  NAND U2437 ( .A(n42766), .B(n42767), .Z(n942) );
  XOR U2438 ( .A(n42766), .B(n42767), .Z(n943) );
  NANDN U2439 ( .A(n42765), .B(n943), .Z(n944) );
  NAND U2440 ( .A(n942), .B(n944), .Z(n42819) );
  NAND U2441 ( .A(n43036), .B(n43035), .Z(n945) );
  XOR U2442 ( .A(n43036), .B(n43035), .Z(n946) );
  NANDN U2443 ( .A(n43037), .B(n946), .Z(n947) );
  NAND U2444 ( .A(n945), .B(n947), .Z(n43116) );
  XOR U2445 ( .A(n43302), .B(n43303), .Z(n948) );
  NANDN U2446 ( .A(n43304), .B(n948), .Z(n949) );
  NAND U2447 ( .A(n43302), .B(n43303), .Z(n950) );
  AND U2448 ( .A(n949), .B(n950), .Z(n43396) );
  XOR U2449 ( .A(n43633), .B(n43632), .Z(n951) );
  NANDN U2450 ( .A(n43634), .B(n951), .Z(n952) );
  NAND U2451 ( .A(n43633), .B(n43632), .Z(n953) );
  AND U2452 ( .A(n952), .B(n953), .Z(n43749) );
  XOR U2453 ( .A(n44604), .B(n44605), .Z(n954) );
  NANDN U2454 ( .A(n44606), .B(n954), .Z(n955) );
  NAND U2455 ( .A(n44604), .B(n44605), .Z(n956) );
  AND U2456 ( .A(n955), .B(n956), .Z(n44762) );
  XNOR U2457 ( .A(n45366), .B(n45365), .Z(n45364) );
  NAND U2458 ( .A(n39600), .B(n39599), .Z(n957) );
  NAND U2459 ( .A(n39605), .B(n39598), .Z(n958) );
  NAND U2460 ( .A(n957), .B(n958), .Z(n39610) );
  NAND U2461 ( .A(n39726), .B(n39723), .Z(n959) );
  NANDN U2462 ( .A(n39726), .B(n39725), .Z(n960) );
  NANDN U2463 ( .A(n39724), .B(n960), .Z(n961) );
  NAND U2464 ( .A(n959), .B(n961), .Z(n39796) );
  XOR U2465 ( .A(n39979), .B(n39980), .Z(n962) );
  NANDN U2466 ( .A(n39981), .B(n962), .Z(n963) );
  NAND U2467 ( .A(n39979), .B(n39980), .Z(n964) );
  AND U2468 ( .A(n963), .B(n964), .Z(n39996) );
  NAND U2469 ( .A(n40413), .B(n40414), .Z(n965) );
  XOR U2470 ( .A(n40413), .B(n40414), .Z(n966) );
  NANDN U2471 ( .A(n40412), .B(n966), .Z(n967) );
  NAND U2472 ( .A(n965), .B(n967), .Z(n40506) );
  XNOR U2473 ( .A(n40869), .B(n40868), .Z(n40863) );
  XOR U2474 ( .A(n41877), .B(n41876), .Z(n968) );
  NANDN U2475 ( .A(n41878), .B(n968), .Z(n969) );
  NAND U2476 ( .A(n41877), .B(n41876), .Z(n970) );
  AND U2477 ( .A(n969), .B(n970), .Z(n42037) );
  NAND U2478 ( .A(n42231), .B(n42230), .Z(n971) );
  NANDN U2479 ( .A(n42233), .B(n42232), .Z(n972) );
  AND U2480 ( .A(n971), .B(n972), .Z(n973) );
  AND U2481 ( .A(n42441), .B(n42440), .Z(n974) );
  NAND U2482 ( .A(n42435), .B(n42434), .Z(n975) );
  XNOR U2483 ( .A(n974), .B(n975), .Z(n976) );
  AND U2484 ( .A(n42239), .B(n42238), .Z(n977) );
  XNOR U2485 ( .A(n42429), .B(n42428), .Z(n978) );
  XNOR U2486 ( .A(n977), .B(n978), .Z(n979) );
  NAND U2487 ( .A(n42443), .B(n42442), .Z(n980) );
  NANDN U2488 ( .A(n42445), .B(n42444), .Z(n981) );
  AND U2489 ( .A(n980), .B(n981), .Z(n982) );
  NAND U2490 ( .A(n42449), .B(n42448), .Z(n983) );
  NANDN U2491 ( .A(n42447), .B(n42446), .Z(n984) );
  AND U2492 ( .A(n983), .B(n984), .Z(n985) );
  XOR U2493 ( .A(n982), .B(n985), .Z(n986) );
  XNOR U2494 ( .A(n976), .B(n979), .Z(n987) );
  XNOR U2495 ( .A(n986), .B(n987), .Z(n988) );
  XNOR U2496 ( .A(n973), .B(n988), .Z(n42450) );
  NAND U2497 ( .A(n36782), .B(n36783), .Z(n989) );
  NAND U2498 ( .A(n36781), .B(n36881), .Z(n990) );
  NAND U2499 ( .A(n989), .B(n990), .Z(n36811) );
  NAND U2500 ( .A(n36872), .B(n36873), .Z(n991) );
  XOR U2501 ( .A(n36872), .B(n36873), .Z(n992) );
  NANDN U2502 ( .A(n36871), .B(n992), .Z(n993) );
  NAND U2503 ( .A(n991), .B(n993), .Z(n36906) );
  XOR U2504 ( .A(n37390), .B(n37389), .Z(n994) );
  NANDN U2505 ( .A(n37388), .B(n994), .Z(n995) );
  NAND U2506 ( .A(n37390), .B(n37389), .Z(n996) );
  AND U2507 ( .A(n995), .B(n996), .Z(n37476) );
  XOR U2508 ( .A(n37669), .B(n37670), .Z(n997) );
  NANDN U2509 ( .A(n37671), .B(n997), .Z(n998) );
  NAND U2510 ( .A(n37669), .B(n37670), .Z(n999) );
  AND U2511 ( .A(n998), .B(n999), .Z(n37767) );
  XOR U2512 ( .A(n38005), .B(n38006), .Z(n1000) );
  NANDN U2513 ( .A(n38007), .B(n1000), .Z(n1001) );
  NAND U2514 ( .A(n38005), .B(n38006), .Z(n1002) );
  AND U2515 ( .A(n1001), .B(n1002), .Z(n38130) );
  NAND U2516 ( .A(n38556), .B(n38557), .Z(n1003) );
  XOR U2517 ( .A(n38556), .B(n38557), .Z(n1004) );
  NANDN U2518 ( .A(n38555), .B(n1004), .Z(n1005) );
  NAND U2519 ( .A(n1003), .B(n1005), .Z(n38700) );
  NAND U2520 ( .A(n39268), .B(n39267), .Z(n1006) );
  NAND U2521 ( .A(n39266), .B(n39265), .Z(n1007) );
  AND U2522 ( .A(n1006), .B(n1007), .Z(n39564) );
  XOR U2523 ( .A(n33998), .B(n33997), .Z(n1008) );
  NANDN U2524 ( .A(n33999), .B(n1008), .Z(n1009) );
  NAND U2525 ( .A(n33998), .B(n33997), .Z(n1010) );
  AND U2526 ( .A(n1009), .B(n1010), .Z(n34038) );
  NAND U2527 ( .A(n34185), .B(n34186), .Z(n1011) );
  XOR U2528 ( .A(n34185), .B(n34186), .Z(n1012) );
  NANDN U2529 ( .A(n34184), .B(n1012), .Z(n1013) );
  NAND U2530 ( .A(n1011), .B(n1013), .Z(n34240) );
  XOR U2531 ( .A(n34737), .B(n34738), .Z(n1014) );
  NANDN U2532 ( .A(n34739), .B(n1014), .Z(n1015) );
  NAND U2533 ( .A(n34737), .B(n34738), .Z(n1016) );
  AND U2534 ( .A(n1015), .B(n1016), .Z(n34842) );
  XOR U2535 ( .A(n35069), .B(n35068), .Z(n1017) );
  NANDN U2536 ( .A(n35070), .B(n1017), .Z(n1018) );
  NAND U2537 ( .A(n35069), .B(n35068), .Z(n1019) );
  AND U2538 ( .A(n1018), .B(n1019), .Z(n35192) );
  NAND U2539 ( .A(n35451), .B(n35452), .Z(n1020) );
  XOR U2540 ( .A(n35451), .B(n35452), .Z(n1021) );
  NAND U2541 ( .A(n1021), .B(n35450), .Z(n1022) );
  NAND U2542 ( .A(n1020), .B(n1022), .Z(n35592) );
  XOR U2543 ( .A(n36325), .B(n36326), .Z(n1023) );
  NANDN U2544 ( .A(n36327), .B(n1023), .Z(n1024) );
  NAND U2545 ( .A(n36325), .B(n36326), .Z(n1025) );
  AND U2546 ( .A(n1024), .B(n1025), .Z(n36745) );
  NAND U2547 ( .A(n31155), .B(n31152), .Z(n1026) );
  NANDN U2548 ( .A(n31155), .B(n31154), .Z(n1027) );
  NANDN U2549 ( .A(n31153), .B(n1027), .Z(n1028) );
  NAND U2550 ( .A(n1026), .B(n1028), .Z(n31192) );
  XOR U2551 ( .A(n31260), .B(n31259), .Z(n1029) );
  NANDN U2552 ( .A(n31261), .B(n1029), .Z(n1030) );
  NAND U2553 ( .A(n31260), .B(n31259), .Z(n1031) );
  AND U2554 ( .A(n1030), .B(n1031), .Z(n31377) );
  NAND U2555 ( .A(n31697), .B(n31698), .Z(n1032) );
  XOR U2556 ( .A(n31697), .B(n31698), .Z(n1033) );
  NANDN U2557 ( .A(n31696), .B(n1033), .Z(n1034) );
  NAND U2558 ( .A(n1032), .B(n1034), .Z(n31792) );
  NAND U2559 ( .A(n32117), .B(n32118), .Z(n1035) );
  XOR U2560 ( .A(n32117), .B(n32118), .Z(n1036) );
  NANDN U2561 ( .A(n32116), .B(n1036), .Z(n1037) );
  NAND U2562 ( .A(n1035), .B(n1037), .Z(n32233) );
  NAND U2563 ( .A(n32638), .B(n32639), .Z(n1038) );
  XOR U2564 ( .A(n32638), .B(n32639), .Z(n1039) );
  NANDN U2565 ( .A(n32637), .B(n1039), .Z(n1040) );
  NAND U2566 ( .A(n1038), .B(n1040), .Z(n32653) );
  XNOR U2567 ( .A(n32939), .B(n32938), .Z(n32932) );
  XOR U2568 ( .A(n33441), .B(n33442), .Z(n1041) );
  NANDN U2569 ( .A(n33443), .B(n1041), .Z(n1042) );
  NAND U2570 ( .A(n33441), .B(n33442), .Z(n1043) );
  AND U2571 ( .A(n1042), .B(n1043), .Z(n33615) );
  XOR U2572 ( .A(n28087), .B(n28088), .Z(n1044) );
  NANDN U2573 ( .A(n28089), .B(n1044), .Z(n1045) );
  NAND U2574 ( .A(n28087), .B(n28088), .Z(n1046) );
  AND U2575 ( .A(n1045), .B(n1046), .Z(n28102) );
  XOR U2576 ( .A(n28186), .B(n28187), .Z(n1047) );
  NANDN U2577 ( .A(n28188), .B(n1047), .Z(n1048) );
  NAND U2578 ( .A(n28186), .B(n28187), .Z(n1049) );
  AND U2579 ( .A(n1048), .B(n1049), .Z(n28233) );
  XOR U2580 ( .A(n29083), .B(n29084), .Z(n1050) );
  NANDN U2581 ( .A(n29085), .B(n1050), .Z(n1051) );
  NAND U2582 ( .A(n29083), .B(n29084), .Z(n1052) );
  AND U2583 ( .A(n1051), .B(n1052), .Z(n29312) );
  NAND U2584 ( .A(n29571), .B(n29572), .Z(n1053) );
  XOR U2585 ( .A(n29571), .B(n29572), .Z(n1054) );
  NAND U2586 ( .A(n1054), .B(n29570), .Z(n1055) );
  NAND U2587 ( .A(n1053), .B(n1055), .Z(n29718) );
  XOR U2588 ( .A(n29872), .B(n29873), .Z(n1056) );
  NANDN U2589 ( .A(n29874), .B(n1056), .Z(n1057) );
  NAND U2590 ( .A(n29872), .B(n29873), .Z(n1058) );
  AND U2591 ( .A(n1057), .B(n1058), .Z(n30171) );
  XOR U2592 ( .A(n30506), .B(n30507), .Z(n1059) );
  NANDN U2593 ( .A(n30508), .B(n1059), .Z(n1060) );
  NAND U2594 ( .A(n30506), .B(n30507), .Z(n1061) );
  AND U2595 ( .A(n1060), .B(n1061), .Z(n30968) );
  NANDN U2596 ( .A(n25157), .B(n25159), .Z(n1062) );
  OR U2597 ( .A(n25159), .B(n25160), .Z(n1063) );
  NAND U2598 ( .A(n25158), .B(n1063), .Z(n1064) );
  NAND U2599 ( .A(n1062), .B(n1064), .Z(n25178) );
  NAND U2600 ( .A(n25233), .B(n25234), .Z(n1065) );
  XOR U2601 ( .A(n25233), .B(n25234), .Z(n1066) );
  NANDN U2602 ( .A(n25232), .B(n1066), .Z(n1067) );
  NAND U2603 ( .A(n1065), .B(n1067), .Z(n25274) );
  XOR U2604 ( .A(n25376), .B(n25377), .Z(n1068) );
  NANDN U2605 ( .A(n25378), .B(n1068), .Z(n1069) );
  NAND U2606 ( .A(n25376), .B(n25377), .Z(n1070) );
  AND U2607 ( .A(n1069), .B(n1070), .Z(n25488) );
  XOR U2608 ( .A(n25734), .B(n25733), .Z(n1071) );
  NANDN U2609 ( .A(n25732), .B(n1071), .Z(n1072) );
  NAND U2610 ( .A(n25734), .B(n25733), .Z(n1073) );
  AND U2611 ( .A(n1072), .B(n1073), .Z(n25819) );
  XOR U2612 ( .A(n26233), .B(n26232), .Z(n1074) );
  NANDN U2613 ( .A(n26234), .B(n1074), .Z(n1075) );
  NAND U2614 ( .A(n26233), .B(n26232), .Z(n1076) );
  AND U2615 ( .A(n1075), .B(n1076), .Z(n26362) );
  XOR U2616 ( .A(n26902), .B(n26903), .Z(n1077) );
  NANDN U2617 ( .A(n26904), .B(n1077), .Z(n1078) );
  NAND U2618 ( .A(n26902), .B(n26903), .Z(n1079) );
  AND U2619 ( .A(n1078), .B(n1079), .Z(n27053) );
  XOR U2620 ( .A(n27560), .B(n27561), .Z(n1080) );
  NANDN U2621 ( .A(n27562), .B(n1080), .Z(n1081) );
  NAND U2622 ( .A(n27560), .B(n27561), .Z(n1082) );
  AND U2623 ( .A(n1081), .B(n1082), .Z(n27736) );
  NANDN U2624 ( .A(n22227), .B(n22229), .Z(n1083) );
  OR U2625 ( .A(n22229), .B(n22230), .Z(n1084) );
  NAND U2626 ( .A(n22228), .B(n1084), .Z(n1085) );
  NAND U2627 ( .A(n1083), .B(n1085), .Z(n22248) );
  XOR U2628 ( .A(n22348), .B(n22349), .Z(n1086) );
  NANDN U2629 ( .A(n22350), .B(n1086), .Z(n1087) );
  NAND U2630 ( .A(n22348), .B(n22349), .Z(n1088) );
  AND U2631 ( .A(n1087), .B(n1088), .Z(n22435) );
  XOR U2632 ( .A(n22636), .B(n22637), .Z(n1089) );
  NANDN U2633 ( .A(n22638), .B(n1089), .Z(n1090) );
  NAND U2634 ( .A(n22636), .B(n22637), .Z(n1091) );
  AND U2635 ( .A(n1090), .B(n1091), .Z(n22714) );
  XOR U2636 ( .A(n23002), .B(n23001), .Z(n1092) );
  NANDN U2637 ( .A(n23000), .B(n1092), .Z(n1093) );
  NAND U2638 ( .A(n23002), .B(n23001), .Z(n1094) );
  AND U2639 ( .A(n1093), .B(n1094), .Z(n23099) );
  XOR U2640 ( .A(n23721), .B(n23722), .Z(n1095) );
  NANDN U2641 ( .A(n23723), .B(n1095), .Z(n1096) );
  NAND U2642 ( .A(n23721), .B(n23722), .Z(n1097) );
  AND U2643 ( .A(n1096), .B(n1097), .Z(n23863) );
  NAND U2644 ( .A(n24341), .B(n24342), .Z(n1098) );
  XOR U2645 ( .A(n24341), .B(n24342), .Z(n1099) );
  NANDN U2646 ( .A(n24340), .B(n1099), .Z(n1100) );
  NAND U2647 ( .A(n1098), .B(n1100), .Z(n24635) );
  XNOR U2648 ( .A(n25072), .B(n25071), .Z(n25070) );
  NAND U2649 ( .A(n19504), .B(n19505), .Z(n1101) );
  XOR U2650 ( .A(n19504), .B(n19505), .Z(n1102) );
  NANDN U2651 ( .A(n19503), .B(n1102), .Z(n1103) );
  NAND U2652 ( .A(n1101), .B(n1103), .Z(n19552) );
  NAND U2653 ( .A(n19648), .B(n19649), .Z(n1104) );
  XOR U2654 ( .A(n19648), .B(n19649), .Z(n1105) );
  NANDN U2655 ( .A(n19647), .B(n1105), .Z(n1106) );
  NAND U2656 ( .A(n1104), .B(n1106), .Z(n19657) );
  NAND U2657 ( .A(n19915), .B(n19912), .Z(n1107) );
  NANDN U2658 ( .A(n19915), .B(n19914), .Z(n1108) );
  NANDN U2659 ( .A(n19913), .B(n1108), .Z(n1109) );
  NAND U2660 ( .A(n1107), .B(n1109), .Z(n19989) );
  NAND U2661 ( .A(n20087), .B(n20088), .Z(n1110) );
  XOR U2662 ( .A(n20087), .B(n20088), .Z(n1111) );
  NANDN U2663 ( .A(n20086), .B(n1111), .Z(n1112) );
  NAND U2664 ( .A(n1110), .B(n1112), .Z(n20182) );
  NAND U2665 ( .A(n20502), .B(n20503), .Z(n1113) );
  XOR U2666 ( .A(n20502), .B(n20503), .Z(n1114) );
  NANDN U2667 ( .A(n20501), .B(n1114), .Z(n1115) );
  NAND U2668 ( .A(n1113), .B(n1115), .Z(n20631) );
  NAND U2669 ( .A(n20886), .B(n20885), .Z(n1116) );
  XOR U2670 ( .A(n20886), .B(n20885), .Z(n1117) );
  NANDN U2671 ( .A(n20887), .B(n1117), .Z(n1118) );
  NAND U2672 ( .A(n1116), .B(n1118), .Z(n21021) );
  XOR U2673 ( .A(n21455), .B(n21454), .Z(n1119) );
  NANDN U2674 ( .A(n21456), .B(n1119), .Z(n1120) );
  NAND U2675 ( .A(n21455), .B(n21454), .Z(n1121) );
  AND U2676 ( .A(n1120), .B(n1121), .Z(n21589) );
  XOR U2677 ( .A(n21726), .B(n21725), .Z(n1122) );
  NANDN U2678 ( .A(n21727), .B(n1122), .Z(n1123) );
  NAND U2679 ( .A(n21726), .B(n21725), .Z(n1124) );
  AND U2680 ( .A(n1123), .B(n1124), .Z(n22159) );
  NAND U2681 ( .A(n16526), .B(n16527), .Z(n1125) );
  NAND U2682 ( .A(n16525), .B(n16619), .Z(n1126) );
  NAND U2683 ( .A(n1125), .B(n1126), .Z(n16545) );
  XOR U2684 ( .A(n16610), .B(n16609), .Z(n1127) );
  NANDN U2685 ( .A(n16611), .B(n1127), .Z(n1128) );
  NAND U2686 ( .A(n16610), .B(n16609), .Z(n1129) );
  AND U2687 ( .A(n1128), .B(n1129), .Z(n16645) );
  XNOR U2688 ( .A(n16701), .B(n16700), .Z(n16694) );
  NAND U2689 ( .A(n16889), .B(n16890), .Z(n1130) );
  XOR U2690 ( .A(n16889), .B(n16890), .Z(n1131) );
  NANDN U2691 ( .A(n16888), .B(n1131), .Z(n1132) );
  NAND U2692 ( .A(n1130), .B(n1132), .Z(n16955) );
  XOR U2693 ( .A(n17651), .B(n17650), .Z(n1133) );
  NANDN U2694 ( .A(n17652), .B(n1133), .Z(n1134) );
  NAND U2695 ( .A(n17651), .B(n17650), .Z(n1135) );
  AND U2696 ( .A(n1134), .B(n1135), .Z(n17765) );
  NAND U2697 ( .A(n18121), .B(n18122), .Z(n1136) );
  XOR U2698 ( .A(n18121), .B(n18122), .Z(n1137) );
  NANDN U2699 ( .A(n18120), .B(n1137), .Z(n1138) );
  NAND U2700 ( .A(n1136), .B(n1138), .Z(n18261) );
  NAND U2701 ( .A(n18571), .B(n18572), .Z(n1139) );
  XOR U2702 ( .A(n18571), .B(n18572), .Z(n1140) );
  NANDN U2703 ( .A(n18570), .B(n1140), .Z(n1141) );
  NAND U2704 ( .A(n1139), .B(n1141), .Z(n18738) );
  XOR U2705 ( .A(n18909), .B(n18910), .Z(n1142) );
  NANDN U2706 ( .A(n18911), .B(n1142), .Z(n1143) );
  NAND U2707 ( .A(n18909), .B(n18910), .Z(n1144) );
  AND U2708 ( .A(n1143), .B(n1144), .Z(n19086) );
  XOR U2709 ( .A(n13710), .B(n13709), .Z(n1145) );
  NANDN U2710 ( .A(n13711), .B(n1145), .Z(n1146) );
  NAND U2711 ( .A(n13710), .B(n13709), .Z(n1147) );
  AND U2712 ( .A(n1146), .B(n1147), .Z(n13727) );
  NAND U2713 ( .A(n13794), .B(n13795), .Z(n1148) );
  XOR U2714 ( .A(n13794), .B(n13795), .Z(n1149) );
  NANDN U2715 ( .A(n13793), .B(n1149), .Z(n1150) );
  NAND U2716 ( .A(n1148), .B(n1150), .Z(n13828) );
  XOR U2717 ( .A(n14154), .B(n14155), .Z(n1151) );
  NANDN U2718 ( .A(n14156), .B(n1151), .Z(n1152) );
  NAND U2719 ( .A(n14154), .B(n14155), .Z(n1153) );
  AND U2720 ( .A(n1152), .B(n1153), .Z(n14230) );
  NAND U2721 ( .A(n14483), .B(n14484), .Z(n1154) );
  XOR U2722 ( .A(n14483), .B(n14484), .Z(n1155) );
  NANDN U2723 ( .A(n14482), .B(n1155), .Z(n1156) );
  NAND U2724 ( .A(n1154), .B(n1156), .Z(n14580) );
  XOR U2725 ( .A(n14809), .B(n14810), .Z(n1157) );
  NANDN U2726 ( .A(n14811), .B(n1157), .Z(n1158) );
  NAND U2727 ( .A(n14809), .B(n14810), .Z(n1159) );
  AND U2728 ( .A(n1158), .B(n1159), .Z(n14926) );
  XOR U2729 ( .A(n15325), .B(n15326), .Z(n1160) );
  NANDN U2730 ( .A(n15327), .B(n1160), .Z(n1161) );
  NAND U2731 ( .A(n15325), .B(n15326), .Z(n1162) );
  AND U2732 ( .A(n1161), .B(n1162), .Z(n15459) );
  NAND U2733 ( .A(n15755), .B(n15756), .Z(n1163) );
  XOR U2734 ( .A(n15755), .B(n15756), .Z(n1164) );
  NANDN U2735 ( .A(n15754), .B(n1164), .Z(n1165) );
  NAND U2736 ( .A(n1163), .B(n1165), .Z(n15891) );
  NAND U2737 ( .A(n16451), .B(n16450), .Z(n1166) );
  NANDN U2738 ( .A(n16453), .B(n16452), .Z(n1167) );
  AND U2739 ( .A(n1166), .B(n1167), .Z(n1168) );
  NAND U2740 ( .A(n16455), .B(n16454), .Z(n1169) );
  NAND U2741 ( .A(n16457), .B(n16456), .Z(n1170) );
  NAND U2742 ( .A(n1169), .B(n1170), .Z(n1171) );
  XNOR U2743 ( .A(n1168), .B(n1171), .Z(n16458) );
  NANDN U2744 ( .A(n10809), .B(n10811), .Z(n1172) );
  OR U2745 ( .A(n10811), .B(n10812), .Z(n1173) );
  NAND U2746 ( .A(n10810), .B(n1173), .Z(n1174) );
  NAND U2747 ( .A(n1172), .B(n1174), .Z(n10830) );
  NAND U2748 ( .A(n10885), .B(n10886), .Z(n1175) );
  XOR U2749 ( .A(n10885), .B(n10886), .Z(n1176) );
  NANDN U2750 ( .A(n10884), .B(n1176), .Z(n1177) );
  NAND U2751 ( .A(n1175), .B(n1177), .Z(n10953) );
  XOR U2752 ( .A(n11232), .B(n11231), .Z(n1178) );
  NANDN U2753 ( .A(n11230), .B(n1178), .Z(n1179) );
  NAND U2754 ( .A(n11232), .B(n11231), .Z(n1180) );
  AND U2755 ( .A(n1179), .B(n1180), .Z(n11384) );
  NAND U2756 ( .A(n11571), .B(n11572), .Z(n1181) );
  XOR U2757 ( .A(n11571), .B(n11572), .Z(n1182) );
  NANDN U2758 ( .A(n11570), .B(n1182), .Z(n1183) );
  NAND U2759 ( .A(n1181), .B(n1183), .Z(n11668) );
  NAND U2760 ( .A(n12710), .B(n12711), .Z(n1184) );
  XOR U2761 ( .A(n12710), .B(n12711), .Z(n1185) );
  NANDN U2762 ( .A(n12709), .B(n1185), .Z(n1186) );
  NAND U2763 ( .A(n1184), .B(n1186), .Z(n12725) );
  NAND U2764 ( .A(n13038), .B(n13039), .Z(n1187) );
  XOR U2765 ( .A(n13038), .B(n13039), .Z(n1188) );
  NANDN U2766 ( .A(n13037), .B(n1188), .Z(n1189) );
  NAND U2767 ( .A(n1187), .B(n1189), .Z(n13198) );
  XOR U2768 ( .A(n13380), .B(n13379), .Z(n13660) );
  NANDN U2769 ( .A(n7881), .B(n7883), .Z(n1190) );
  OR U2770 ( .A(n7883), .B(n7884), .Z(n1191) );
  NAND U2771 ( .A(n7882), .B(n1191), .Z(n1192) );
  NAND U2772 ( .A(n1190), .B(n1192), .Z(n7902) );
  NAND U2773 ( .A(n8032), .B(n8033), .Z(n1193) );
  XOR U2774 ( .A(n8032), .B(n8033), .Z(n1194) );
  NANDN U2775 ( .A(n8031), .B(n1194), .Z(n1195) );
  NAND U2776 ( .A(n1193), .B(n1195), .Z(n8088) );
  XOR U2777 ( .A(n8154), .B(n8153), .Z(n1196) );
  NANDN U2778 ( .A(n8155), .B(n1196), .Z(n1197) );
  NAND U2779 ( .A(n8154), .B(n8153), .Z(n1198) );
  AND U2780 ( .A(n1197), .B(n1198), .Z(n8281) );
  NAND U2781 ( .A(n9374), .B(n9375), .Z(n1199) );
  XOR U2782 ( .A(n9374), .B(n9375), .Z(n1200) );
  NANDN U2783 ( .A(n9373), .B(n1200), .Z(n1201) );
  NAND U2784 ( .A(n1199), .B(n1201), .Z(n9521) );
  NAND U2785 ( .A(n9809), .B(n9810), .Z(n1202) );
  XOR U2786 ( .A(n9809), .B(n9810), .Z(n1203) );
  NANDN U2787 ( .A(n9808), .B(n1203), .Z(n1204) );
  NAND U2788 ( .A(n1202), .B(n1204), .Z(n9818) );
  NAND U2789 ( .A(n10481), .B(n10480), .Z(n1205) );
  NAND U2790 ( .A(n10482), .B(n10483), .Z(n1206) );
  AND U2791 ( .A(n1205), .B(n1206), .Z(n1207) );
  AND U2792 ( .A(n10691), .B(n10690), .Z(n1208) );
  NAND U2793 ( .A(n10685), .B(n10684), .Z(n1209) );
  XNOR U2794 ( .A(n1208), .B(n1209), .Z(n1210) );
  AND U2795 ( .A(n10489), .B(n10488), .Z(n1211) );
  XNOR U2796 ( .A(n10679), .B(n10678), .Z(n1212) );
  XNOR U2797 ( .A(n1211), .B(n1212), .Z(n1213) );
  NAND U2798 ( .A(n10693), .B(n10692), .Z(n1214) );
  NANDN U2799 ( .A(n10695), .B(n10694), .Z(n1215) );
  AND U2800 ( .A(n1214), .B(n1215), .Z(n1216) );
  NANDN U2801 ( .A(n10698), .B(n10697), .Z(n1217) );
  NANDN U2802 ( .A(n10700), .B(n10699), .Z(n1218) );
  AND U2803 ( .A(n1217), .B(n1218), .Z(n1219) );
  XOR U2804 ( .A(n1216), .B(n1219), .Z(n1220) );
  XNOR U2805 ( .A(n1210), .B(n1213), .Z(n1221) );
  XNOR U2806 ( .A(n1220), .B(n1221), .Z(n1222) );
  XNOR U2807 ( .A(n1207), .B(n1222), .Z(n10701) );
  NANDN U2808 ( .A(n4926), .B(n4928), .Z(n1223) );
  OR U2809 ( .A(n4928), .B(n4929), .Z(n1224) );
  NAND U2810 ( .A(n4927), .B(n1224), .Z(n1225) );
  NAND U2811 ( .A(n1223), .B(n1225), .Z(n4947) );
  XNOR U2812 ( .A(n5081), .B(n5080), .Z(n5077) );
  NAND U2813 ( .A(n5419), .B(n5420), .Z(n1226) );
  XOR U2814 ( .A(n5419), .B(n5420), .Z(n1227) );
  NANDN U2815 ( .A(n5418), .B(n1227), .Z(n1228) );
  NAND U2816 ( .A(n1226), .B(n1228), .Z(n5504) );
  XOR U2817 ( .A(n5694), .B(n5693), .Z(n1229) );
  NANDN U2818 ( .A(n5692), .B(n1229), .Z(n1230) );
  NAND U2819 ( .A(n5694), .B(n5693), .Z(n1231) );
  AND U2820 ( .A(n1230), .B(n1231), .Z(n5791) );
  XOR U2821 ( .A(n7168), .B(n7169), .Z(n1232) );
  NANDN U2822 ( .A(n7170), .B(n1232), .Z(n1233) );
  NAND U2823 ( .A(n7168), .B(n7169), .Z(n1234) );
  AND U2824 ( .A(n1233), .B(n1234), .Z(n7330) );
  XNOR U2825 ( .A(n7519), .B(n7518), .Z(n7516) );
  XOR U2826 ( .A(n2026), .B(n2025), .Z(n1235) );
  NANDN U2827 ( .A(n2027), .B(n1235), .Z(n1236) );
  NAND U2828 ( .A(n2026), .B(n2025), .Z(n1237) );
  AND U2829 ( .A(n1236), .B(n1237), .Z(n2053) );
  NAND U2830 ( .A(n2146), .B(n2147), .Z(n1238) );
  XOR U2831 ( .A(n2146), .B(n2147), .Z(n1239) );
  NANDN U2832 ( .A(n2145), .B(n1239), .Z(n1240) );
  NAND U2833 ( .A(n1238), .B(n1240), .Z(n2161) );
  NAND U2834 ( .A(n2679), .B(n2678), .Z(n1241) );
  XOR U2835 ( .A(n2679), .B(n2678), .Z(n1242) );
  NANDN U2836 ( .A(n2680), .B(n1242), .Z(n1243) );
  NAND U2837 ( .A(n1241), .B(n1243), .Z(n2774) );
  NAND U2838 ( .A(n2977), .B(n2978), .Z(n1244) );
  XOR U2839 ( .A(n2977), .B(n2978), .Z(n1245) );
  NANDN U2840 ( .A(n2976), .B(n1245), .Z(n1246) );
  NAND U2841 ( .A(n1244), .B(n1246), .Z(n2986) );
  XOR U2842 ( .A(n3462), .B(n3461), .Z(n1247) );
  NANDN U2843 ( .A(n3463), .B(n1247), .Z(n1248) );
  NAND U2844 ( .A(n3462), .B(n3461), .Z(n1249) );
  AND U2845 ( .A(n1248), .B(n1249), .Z(n3609) );
  NAND U2846 ( .A(n3893), .B(n3894), .Z(n1250) );
  XOR U2847 ( .A(n3893), .B(n3894), .Z(n1251) );
  NANDN U2848 ( .A(n3892), .B(n1251), .Z(n1252) );
  NAND U2849 ( .A(n1250), .B(n1252), .Z(n3908) );
  NAND U2850 ( .A(n4554), .B(n4555), .Z(n1253) );
  XOR U2851 ( .A(n4554), .B(n4555), .Z(n1254) );
  NANDN U2852 ( .A(n4553), .B(n1254), .Z(n1255) );
  NAND U2853 ( .A(n1253), .B(n1255), .Z(n4564) );
  XNOR U2854 ( .A(n32343), .B(n32342), .Z(n32345) );
  XNOR U2855 ( .A(n32440), .B(n32439), .Z(n32442) );
  XNOR U2856 ( .A(n32453), .B(n32452), .Z(n32429) );
  XNOR U2857 ( .A(n29807), .B(n29806), .Z(n29808) );
  XNOR U2858 ( .A(n29986), .B(n30140), .Z(n29762) );
  XNOR U2859 ( .A(n23926), .B(n23925), .Z(n23928) );
  XNOR U2860 ( .A(n23947), .B(n23946), .Z(n23949) );
  XNOR U2861 ( .A(n23744), .B(n23743), .Z(n23745) );
  XNOR U2862 ( .A(n24100), .B(n24099), .Z(n24101) );
  XNOR U2863 ( .A(n9725), .B(n9724), .Z(n9726) );
  XNOR U2864 ( .A(n6804), .B(n6987), .Z(n6599) );
  XNOR U2865 ( .A(n46168), .B(n46167), .Z(n46169) );
  XNOR U2866 ( .A(n46301), .B(n46300), .Z(n46302) );
  XNOR U2867 ( .A(n46489), .B(n46488), .Z(n46525) );
  XOR U2868 ( .A(n46715), .B(n46714), .Z(n46731) );
  XNOR U2869 ( .A(n46916), .B(n46915), .Z(n46879) );
  XNOR U2870 ( .A(n46975), .B(n46974), .Z(n47013) );
  NAND U2871 ( .A(n47133), .B(n47134), .Z(n1256) );
  NAND U2872 ( .A(n47132), .B(n48097), .Z(n1257) );
  NAND U2873 ( .A(n1256), .B(n1257), .Z(n47340) );
  XNOR U2874 ( .A(n43367), .B(n43366), .Z(n43344) );
  XNOR U2875 ( .A(n43588), .B(n43587), .Z(n43531) );
  XNOR U2876 ( .A(n44082), .B(n44081), .Z(n44084) );
  XNOR U2877 ( .A(n44210), .B(n44209), .Z(n44262) );
  XNOR U2878 ( .A(n44197), .B(n44198), .Z(n44286) );
  XNOR U2879 ( .A(n44567), .B(n44566), .Z(n44568) );
  XNOR U2880 ( .A(n40477), .B(n40476), .Z(n40456) );
  XNOR U2881 ( .A(n40576), .B(n40575), .Z(n40536) );
  XNOR U2882 ( .A(n40675), .B(n40816), .Z(n40647) );
  XNOR U2883 ( .A(n40779), .B(n40778), .Z(n40780) );
  XOR U2884 ( .A(n40894), .B(n40893), .Z(n40910) );
  XNOR U2885 ( .A(n41108), .B(n41107), .Z(n41071) );
  XNOR U2886 ( .A(n41196), .B(n41195), .Z(n41197) );
  NAND U2887 ( .A(n41204), .B(n41203), .Z(n1258) );
  NAND U2888 ( .A(n41201), .B(n41202), .Z(n1259) );
  NAND U2889 ( .A(n1258), .B(n1259), .Z(n41388) );
  XNOR U2890 ( .A(n37797), .B(n37796), .Z(n37842) );
  XNOR U2891 ( .A(n37834), .B(n37833), .Z(n37784) );
  XNOR U2892 ( .A(n38233), .B(n38232), .Z(n38196) );
  XNOR U2893 ( .A(n38065), .B(n38064), .Z(n38115) );
  XNOR U2894 ( .A(n38296), .B(n38295), .Z(n38333) );
  XNOR U2895 ( .A(n38370), .B(n38369), .Z(n38372) );
  XNOR U2896 ( .A(n38479), .B(n38478), .Z(n38473) );
  XNOR U2897 ( .A(n38634), .B(n38633), .Z(n38636) );
  XNOR U2898 ( .A(n35024), .B(n35023), .Z(n34962) );
  XNOR U2899 ( .A(n35423), .B(n35422), .Z(n35386) );
  XNOR U2900 ( .A(n35482), .B(n35481), .Z(n35519) );
  XNOR U2901 ( .A(n35393), .B(n35392), .Z(n35360) );
  XNOR U2902 ( .A(n35680), .B(n35679), .Z(n35674) );
  XNOR U2903 ( .A(n35718), .B(n35717), .Z(n35639) );
  XNOR U2904 ( .A(n35834), .B(n35833), .Z(n35835) );
  XNOR U2905 ( .A(n35883), .B(n35882), .Z(n35884) );
  XNOR U2906 ( .A(n35830), .B(n35829), .Z(n35870) );
  XNOR U2907 ( .A(n32457), .B(n32456), .Z(n32458) );
  XNOR U2908 ( .A(n32300), .B(n32299), .Z(n32317) );
  XNOR U2909 ( .A(n32588), .B(n32587), .Z(n32518) );
  XNOR U2910 ( .A(n32681), .B(n32680), .Z(n32675) );
  XNOR U2911 ( .A(n32863), .B(n32862), .Z(n32865) );
  XNOR U2912 ( .A(n28934), .B(n28933), .Z(n28935) );
  XNOR U2913 ( .A(n29110), .B(n29109), .Z(n29155) );
  XNOR U2914 ( .A(n29147), .B(n29146), .Z(n29097) );
  XNOR U2915 ( .A(n29543), .B(n29542), .Z(n29506) );
  XNOR U2916 ( .A(n29513), .B(n29512), .Z(n29480) );
  XNOR U2917 ( .A(n29791), .B(n29790), .Z(n29785) );
  XNOR U2918 ( .A(n29823), .B(n29822), .Z(n29750) );
  XNOR U2919 ( .A(n30010), .B(n30009), .Z(n30011) );
  XNOR U2920 ( .A(n25983), .B(n25982), .Z(n25993) );
  NAND U2921 ( .A(n26062), .B(n26061), .Z(n1260) );
  NANDN U2922 ( .A(n27153), .B(n26060), .Z(n1261) );
  NAND U2923 ( .A(n1260), .B(n1261), .Z(n26173) );
  XNOR U2924 ( .A(n26194), .B(n26193), .Z(n26131) );
  XNOR U2925 ( .A(n26554), .B(n26553), .Z(n26556) );
  XNOR U2926 ( .A(n26579), .B(n26578), .Z(n26542) );
  XNOR U2927 ( .A(n26708), .B(n26707), .Z(n26638) );
  XNOR U2928 ( .A(n26814), .B(n26813), .Z(n26866) );
  XNOR U2929 ( .A(n26801), .B(n26802), .Z(n26891) );
  XNOR U2930 ( .A(n23017), .B(n23016), .Z(n23040) );
  XNOR U2931 ( .A(n23031), .B(n23030), .Z(n23033) );
  XNOR U2932 ( .A(n23288), .B(n23287), .Z(n23238) );
  XNOR U2933 ( .A(n23669), .B(n23668), .Z(n23671) );
  XNOR U2934 ( .A(n23694), .B(n23693), .Z(n23657) );
  XNOR U2935 ( .A(n23675), .B(n23674), .Z(n23631) );
  XNOR U2936 ( .A(n23646), .B(n23645), .Z(n23625) );
  XNOR U2937 ( .A(n23791), .B(n23790), .Z(n23793) );
  XNOR U2938 ( .A(n23763), .B(n23762), .Z(n23765) );
  XOR U2939 ( .A(n24058), .B(n24057), .Z(n24062) );
  XNOR U2940 ( .A(n23910), .B(n23909), .Z(n23904) );
  XNOR U2941 ( .A(n24068), .B(n24067), .Z(n24070) );
  XNOR U2942 ( .A(n23915), .B(n23916), .Z(n24006) );
  XNOR U2943 ( .A(n23984), .B(n23983), .Z(n24000) );
  XNOR U2944 ( .A(n24136), .B(n24135), .Z(n24137) );
  XOR U2945 ( .A(n24280), .B(n24279), .Z(n24290) );
  XNOR U2946 ( .A(n20162), .B(n20161), .Z(n20164) );
  XNOR U2947 ( .A(n20203), .B(n20202), .Z(n20257) );
  XNOR U2948 ( .A(n20698), .B(n20697), .Z(n20700) );
  XNOR U2949 ( .A(n20653), .B(n20652), .Z(n20654) );
  XNOR U2950 ( .A(n20720), .B(n20719), .Z(n20721) );
  XNOR U2951 ( .A(n20714), .B(n20713), .Z(n20716) );
  XNOR U2952 ( .A(n20852), .B(n20851), .Z(n20815) );
  XNOR U2953 ( .A(n21114), .B(n21113), .Z(n21065) );
  XNOR U2954 ( .A(n21102), .B(n21101), .Z(n21078) );
  NAND U2955 ( .A(n17720), .B(n17719), .Z(n1262) );
  NAND U2956 ( .A(n17717), .B(n17718), .Z(n1263) );
  NAND U2957 ( .A(n1262), .B(n1263), .Z(n17843) );
  XNOR U2958 ( .A(n18019), .B(n18018), .Z(n18021) );
  XNOR U2959 ( .A(n18025), .B(n18024), .Z(n18027) );
  XNOR U2960 ( .A(n18190), .B(n18189), .Z(n18184) );
  XNOR U2961 ( .A(n18345), .B(n18344), .Z(n18347) );
  XNOR U2962 ( .A(n14542), .B(n14541), .Z(n14556) );
  XNOR U2963 ( .A(n14849), .B(o[148]), .Z(n14842) );
  XOR U2964 ( .A(n14970), .B(n14969), .Z(n14986) );
  NAND U2965 ( .A(n14890), .B(n14889), .Z(n1264) );
  NANDN U2966 ( .A(n14888), .B(n14887), .Z(n1265) );
  NAND U2967 ( .A(n1264), .B(n1265), .Z(n15040) );
  XNOR U2968 ( .A(n15210), .B(n15209), .Z(n15247) );
  XNOR U2969 ( .A(n15356), .B(n15355), .Z(n15344) );
  XNOR U2970 ( .A(n15373), .B(n15372), .Z(n15350) );
  XNOR U2971 ( .A(n15502), .B(n15501), .Z(n15504) );
  XOR U2972 ( .A(n15577), .B(n15576), .Z(n15508) );
  XNOR U2973 ( .A(n11360), .B(o[110]), .Z(n11352) );
  XNOR U2974 ( .A(n11551), .B(n11550), .Z(n11553) );
  XNOR U2975 ( .A(n11592), .B(n11591), .Z(n11646) );
  XNOR U2976 ( .A(n11639), .B(n11638), .Z(n11616) );
  XNOR U2977 ( .A(n12277), .B(n12276), .Z(n12240) );
  XNOR U2978 ( .A(n12369), .B(n12368), .Z(n12356) );
  XNOR U2979 ( .A(n12400), .B(n12399), .Z(n12331) );
  NAND U2980 ( .A(n12502), .B(n12503), .Z(n1266) );
  NAND U2981 ( .A(n12501), .B(n13505), .Z(n1267) );
  NAND U2982 ( .A(n1266), .B(n1267), .Z(n12663) );
  NAND U2983 ( .A(n12473), .B(n12474), .Z(n1268) );
  NAND U2984 ( .A(n12472), .B(n13429), .Z(n1269) );
  NAND U2985 ( .A(n1268), .B(n1269), .Z(n12703) );
  XNOR U2986 ( .A(n8580), .B(o[80]), .Z(n8594) );
  XNOR U2987 ( .A(n8711), .B(n8710), .Z(n8725) );
  XNOR U2988 ( .A(n8720), .B(n8719), .Z(n8697) );
  XNOR U2989 ( .A(n8668), .B(n8667), .Z(n8691) );
  XNOR U2990 ( .A(n8682), .B(n8681), .Z(n8684) );
  XNOR U2991 ( .A(n9346), .B(n9345), .Z(n9309) );
  XNOR U2992 ( .A(n9465), .B(n9464), .Z(n9395) );
  XOR U2993 ( .A(n9785), .B(n9784), .Z(n9787) );
  XNOR U2994 ( .A(n9779), .B(n9778), .Z(n9781) );
  XOR U2995 ( .A(n9882), .B(n9881), .Z(n9884) );
  XNOR U2996 ( .A(n5673), .B(n5672), .Z(n5675) );
  XNOR U2997 ( .A(n5714), .B(n5713), .Z(n5768) );
  XNOR U2998 ( .A(n5761), .B(n5760), .Z(n5738) );
  XNOR U2999 ( .A(n5860), .B(n5859), .Z(n5820) );
  XNOR U3000 ( .A(n5963), .B(n6103), .Z(n5935) );
  XOR U3001 ( .A(n6072), .B(n6071), .Z(n6074) );
  XNOR U3002 ( .A(n6050), .B(n6049), .Z(n6051) );
  XNOR U3003 ( .A(n6397), .B(n6396), .Z(n6360) );
  XNOR U3004 ( .A(n6447), .B(n6446), .Z(n6482) );
  NAND U3005 ( .A(n6354), .B(n6355), .Z(n1270) );
  NAND U3006 ( .A(n6356), .B(n6357), .Z(n1271) );
  NAND U3007 ( .A(n1270), .B(n1271), .Z(n6476) );
  XNOR U3008 ( .A(n6806), .B(n6805), .Z(n6821) );
  XNOR U3009 ( .A(n6776), .B(n6775), .Z(n6815) );
  NAND U3010 ( .A(n6603), .B(n6604), .Z(n1272) );
  NANDN U3011 ( .A(n6606), .B(n6605), .Z(n1273) );
  AND U3012 ( .A(n1272), .B(n1273), .Z(n6749) );
  XNOR U3013 ( .A(n3046), .B(n3045), .Z(n3047) );
  XNOR U3014 ( .A(n3428), .B(n3427), .Z(n3392) );
  XNOR U3015 ( .A(n3493), .B(n3492), .Z(n3530) );
  XNOR U3016 ( .A(n3675), .B(n3676), .Z(n3654) );
  XNOR U3017 ( .A(n3690), .B(n3689), .Z(n3630) );
  XNOR U3018 ( .A(n45812), .B(n45811), .Z(n45814) );
  XOR U3019 ( .A(n45834), .B(n45835), .Z(n45819) );
  XNOR U3020 ( .A(n46188), .B(n46187), .Z(n46190) );
  XNOR U3021 ( .A(n46512), .B(n46511), .Z(n46459) );
  XNOR U3022 ( .A(n46738), .B(n46737), .Z(n46782) );
  XNOR U3023 ( .A(n46897), .B(n46896), .Z(n46853) );
  XNOR U3024 ( .A(n47037), .B(n47036), .Z(n47039) );
  XNOR U3025 ( .A(n47045), .B(n47044), .Z(n46996) );
  XOR U3026 ( .A(n47403), .B(n47402), .Z(n47429) );
  XNOR U3027 ( .A(n47548), .B(n47547), .Z(n47549) );
  NAND U3028 ( .A(n47476), .B(n47475), .Z(n1274) );
  XOR U3029 ( .A(n47476), .B(n47475), .Z(n1275) );
  NANDN U3030 ( .A(n47474), .B(n1275), .Z(n1276) );
  NAND U3031 ( .A(n1274), .B(n1276), .Z(n47663) );
  XOR U3032 ( .A(n42932), .B(n42933), .Z(n42917) );
  NAND U3033 ( .A(n42853), .B(n42854), .Z(n1277) );
  NAND U3034 ( .A(n42852), .B(n43143), .Z(n1278) );
  NAND U3035 ( .A(n1277), .B(n1278), .Z(n42909) );
  NAND U3036 ( .A(n43071), .B(n43070), .Z(n1279) );
  NANDN U3037 ( .A(n43543), .B(n43069), .Z(n1280) );
  AND U3038 ( .A(n1279), .B(n1280), .Z(n43161) );
  NAND U3039 ( .A(n43086), .B(n43087), .Z(n1281) );
  NAND U3040 ( .A(n43131), .B(n44849), .Z(n1282) );
  NAND U3041 ( .A(n1281), .B(n1282), .Z(n43155) );
  XNOR U3042 ( .A(n43552), .B(n43551), .Z(n43558) );
  XNOR U3043 ( .A(n43440), .B(n43439), .Z(n43512) );
  XNOR U3044 ( .A(n43484), .B(n43483), .Z(n43507) );
  XNOR U3045 ( .A(n43490), .B(n43489), .Z(n43500) );
  XNOR U3046 ( .A(n44227), .B(n44226), .Z(n44229) );
  XNOR U3047 ( .A(n44526), .B(n44525), .Z(n44519) );
  XOR U3048 ( .A(n44635), .B(n44634), .Z(n44738) );
  OR U3049 ( .A(n40351), .B(n40483), .Z(n1283) );
  NAND U3050 ( .A(n40352), .B(n40353), .Z(n1284) );
  AND U3051 ( .A(n1283), .B(n1284), .Z(n40461) );
  NAND U3052 ( .A(n40452), .B(n40453), .Z(n1285) );
  NANDN U3053 ( .A(n40455), .B(n40454), .Z(n1286) );
  AND U3054 ( .A(n1285), .B(n1286), .Z(n40595) );
  XNOR U3055 ( .A(n40541), .B(n40540), .Z(n40613) );
  XNOR U3056 ( .A(n40585), .B(n40584), .Z(n40608) );
  XNOR U3057 ( .A(n40591), .B(n40590), .Z(n40601) );
  XOR U3058 ( .A(n40759), .B(n40758), .Z(n40829) );
  XNOR U3059 ( .A(n40791), .B(n40790), .Z(n40793) );
  XOR U3060 ( .A(n40704), .B(n40703), .Z(n40721) );
  XNOR U3061 ( .A(n40644), .B(n40643), .Z(n40725) );
  XNOR U3062 ( .A(n40971), .B(n40970), .Z(n40973) );
  XNOR U3063 ( .A(n41089), .B(n41088), .Z(n41045) );
  XNOR U3064 ( .A(n37810), .B(n37809), .Z(n37848) );
  XNOR U3065 ( .A(n37933), .B(n37932), .Z(n37935) );
  XNOR U3066 ( .A(n37970), .B(n37969), .Z(n37972) );
  XNOR U3067 ( .A(n38420), .B(n38419), .Z(n38422) );
  XNOR U3068 ( .A(n38778), .B(n38777), .Z(n38779) );
  XOR U3069 ( .A(n34361), .B(n34362), .Z(n34346) );
  NAND U3070 ( .A(n34515), .B(n34514), .Z(n1287) );
  NAND U3071 ( .A(n34561), .B(n36240), .Z(n1288) );
  AND U3072 ( .A(n1287), .B(n1288), .Z(n34589) );
  XNOR U3073 ( .A(n34760), .B(n34759), .Z(n34783) );
  XNOR U3074 ( .A(n34774), .B(n34773), .Z(n34775) );
  XNOR U3075 ( .A(n34988), .B(n34987), .Z(n34994) );
  XNOR U3076 ( .A(n35558), .B(n35557), .Z(n35546) );
  XNOR U3077 ( .A(n35552), .B(n35551), .Z(n35503) );
  XOR U3078 ( .A(n35879), .B(n35878), .Z(n35802) );
  AND U3079 ( .A(n35938), .B(o[378]), .Z(n36112) );
  XNOR U3080 ( .A(n36025), .B(n36024), .Z(n36026) );
  XOR U3081 ( .A(n36021), .B(n36020), .Z(n35960) );
  NAND U3082 ( .A(n35979), .B(n35978), .Z(n1289) );
  NAND U3083 ( .A(n35977), .B(n36100), .Z(n1290) );
  NAND U3084 ( .A(n1289), .B(n1290), .Z(n36069) );
  XNOR U3085 ( .A(n31391), .B(n31390), .Z(n31393) );
  XOR U3086 ( .A(n31413), .B(n31414), .Z(n31398) );
  NAND U3087 ( .A(n31479), .B(n31478), .Z(n1291) );
  NANDN U3088 ( .A(n32036), .B(n31477), .Z(n1292) );
  NAND U3089 ( .A(n1291), .B(n1292), .Z(n31575) );
  XNOR U3090 ( .A(n32274), .B(n32273), .Z(n32276) );
  XNOR U3091 ( .A(n32735), .B(n32734), .Z(n32737) );
  XNOR U3092 ( .A(n28451), .B(n28450), .Z(n28453) );
  XOR U3093 ( .A(n28473), .B(n28474), .Z(n28458) );
  XNOR U3094 ( .A(n28729), .B(n28728), .Z(n28708) );
  NAND U3095 ( .A(n28802), .B(n28803), .Z(n1293) );
  NAND U3096 ( .A(n29007), .B(n29601), .Z(n1294) );
  NAND U3097 ( .A(n1293), .B(n1294), .Z(n28913) );
  NAND U3098 ( .A(n28903), .B(n28904), .Z(n1295) );
  NANDN U3099 ( .A(n28906), .B(n28905), .Z(n1296) );
  AND U3100 ( .A(n1295), .B(n1296), .Z(n29050) );
  XNOR U3101 ( .A(n29123), .B(n29122), .Z(n29161) );
  XNOR U3102 ( .A(n29239), .B(n29238), .Z(n29241) );
  XNOR U3103 ( .A(n29276), .B(n29275), .Z(n29278) );
  XNOR U3104 ( .A(n29678), .B(n29677), .Z(n29666) );
  XNOR U3105 ( .A(n29672), .B(n29671), .Z(n29623) );
  XOR U3106 ( .A(n30006), .B(n30005), .Z(n29930) );
  XNOR U3107 ( .A(n30077), .B(n30076), .Z(n30079) );
  OR U3108 ( .A(n25988), .B(n26936), .Z(n1297) );
  NANDN U3109 ( .A(n25990), .B(n25989), .Z(n1298) );
  NAND U3110 ( .A(n1297), .B(n1298), .Z(n26090) );
  XNOR U3111 ( .A(n26158), .B(n26157), .Z(n26164) );
  XNOR U3112 ( .A(n26560), .B(n26559), .Z(n26516) );
  XNOR U3113 ( .A(n26831), .B(n26830), .Z(n26833) );
  XNOR U3114 ( .A(n27216), .B(o[282]), .Z(n27162) );
  XNOR U3115 ( .A(n27208), .B(n27207), .Z(n27148) );
  XNOR U3116 ( .A(n22692), .B(o[237]), .Z(n22680) );
  XNOR U3117 ( .A(n22776), .B(n23058), .Z(n22785) );
  XNOR U3118 ( .A(n22687), .B(n23692), .Z(n22670) );
  XNOR U3119 ( .A(n22791), .B(n22790), .Z(n22793) );
  XNOR U3120 ( .A(n22767), .B(n22766), .Z(n22739) );
  XOR U3121 ( .A(n22832), .B(n22831), .Z(n22866) );
  XNOR U3122 ( .A(n23264), .B(n23263), .Z(n23302) );
  XNOR U3123 ( .A(n23739), .B(n23738), .Z(n23820) );
  XNOR U3124 ( .A(n24108), .B(n24107), .Z(n24080) );
  XNOR U3125 ( .A(n24074), .B(n24073), .Z(n24076) );
  XNOR U3126 ( .A(n24322), .B(n24321), .Z(n24324) );
  XNOR U3127 ( .A(n24198), .B(n24197), .Z(n24199) );
  XNOR U3128 ( .A(n24296), .B(n24295), .Z(n24298) );
  XNOR U3129 ( .A(n24254), .B(n24253), .Z(n24256) );
  XNOR U3130 ( .A(n24248), .B(n24247), .Z(n24250) );
  XNOR U3131 ( .A(n24561), .B(n24743), .Z(n24562) );
  NAND U3132 ( .A(n19865), .B(n19864), .Z(n1299) );
  NANDN U3133 ( .A(n20420), .B(n19863), .Z(n1300) );
  NAND U3134 ( .A(n1299), .B(n1300), .Z(n19973) );
  XNOR U3135 ( .A(n20262), .B(n20261), .Z(n20264) );
  XNOR U3136 ( .A(n20119), .B(n20118), .Z(n20108) );
  XNOR U3137 ( .A(n20234), .B(n20233), .Z(n20236) );
  XNOR U3138 ( .A(n20212), .B(n20211), .Z(n20214) );
  XNOR U3139 ( .A(n20339), .B(n20338), .Z(n20356) );
  XOR U3140 ( .A(n20548), .B(n20547), .Z(n20590) );
  XNOR U3141 ( .A(n20524), .B(n20523), .Z(n20525) );
  XNOR U3142 ( .A(n20454), .B(n20453), .Z(n20455) );
  XNOR U3143 ( .A(n20445), .B(n20444), .Z(n20393) );
  XNOR U3144 ( .A(n20427), .B(n20577), .Z(n20398) );
  XNOR U3145 ( .A(n20597), .B(n20596), .Z(n20551) );
  XNOR U3146 ( .A(n20647), .B(n20646), .Z(n20649) );
  XNOR U3147 ( .A(n20786), .B(n20785), .Z(n20861) );
  XNOR U3148 ( .A(n20856), .B(n20855), .Z(n20858) );
  XNOR U3149 ( .A(n20981), .B(n20980), .Z(n20987) );
  XNOR U3150 ( .A(n20975), .B(n20974), .Z(n20932) );
  NAND U3151 ( .A(n21293), .B(n21292), .Z(n1301) );
  NAND U3152 ( .A(n21291), .B(n21290), .Z(n1302) );
  AND U3153 ( .A(n1301), .B(n1302), .Z(n21327) );
  NAND U3154 ( .A(n21274), .B(n21273), .Z(n1303) );
  NAND U3155 ( .A(n21272), .B(n21271), .Z(n1304) );
  AND U3156 ( .A(n1303), .B(n1304), .Z(n21319) );
  NAND U3157 ( .A(n21283), .B(n21282), .Z(n1305) );
  NAND U3158 ( .A(n21281), .B(n21280), .Z(n1306) );
  AND U3159 ( .A(n1305), .B(n1306), .Z(n21371) );
  NAND U3160 ( .A(n21220), .B(n21219), .Z(n1307) );
  NAND U3161 ( .A(n21218), .B(n21217), .Z(n1308) );
  AND U3162 ( .A(n1307), .B(n1308), .Z(n21367) );
  XNOR U3163 ( .A(n21401), .B(n21400), .Z(n21403) );
  NAND U3164 ( .A(n21377), .B(n21376), .Z(n1309) );
  NAND U3165 ( .A(n21375), .B(n21503), .Z(n1310) );
  NAND U3166 ( .A(n1309), .B(n1310), .Z(n21476) );
  NAND U3167 ( .A(n21334), .B(n21333), .Z(n1311) );
  NAND U3168 ( .A(n21331), .B(n21332), .Z(n1312) );
  NAND U3169 ( .A(n1311), .B(n1312), .Z(n21480) );
  XNOR U3170 ( .A(n16899), .B(n16898), .Z(n16901) );
  XOR U3171 ( .A(n16921), .B(n16922), .Z(n16906) );
  XNOR U3172 ( .A(n17378), .B(n17377), .Z(n17361) );
  NAND U3173 ( .A(n17666), .B(n17667), .Z(n1313) );
  NAND U3174 ( .A(n17665), .B(n18453), .Z(n1314) );
  NAND U3175 ( .A(n1313), .B(n1314), .Z(n17838) );
  NAND U3176 ( .A(n17695), .B(n17696), .Z(n1315) );
  NAND U3177 ( .A(n17694), .B(n18446), .Z(n1316) );
  NAND U3178 ( .A(n1315), .B(n1316), .Z(n17779) );
  NAND U3179 ( .A(n17835), .B(n18013), .Z(n1317) );
  NAND U3180 ( .A(n17956), .B(n18985), .Z(n1318) );
  NAND U3181 ( .A(n1317), .B(n1318), .Z(n17899) );
  NAND U3182 ( .A(n17828), .B(n17829), .Z(n1319) );
  NAND U3183 ( .A(n17826), .B(n17827), .Z(n1320) );
  NAND U3184 ( .A(n1319), .B(n1320), .Z(n17889) );
  NAND U3185 ( .A(n17790), .B(n17789), .Z(n1321) );
  NANDN U3186 ( .A(n18455), .B(n17927), .Z(n1322) );
  AND U3187 ( .A(n1321), .B(n1322), .Z(n17906) );
  XNOR U3188 ( .A(n18067), .B(n18066), .Z(n18083) );
  XNOR U3189 ( .A(n18073), .B(n18072), .Z(n18095) );
  XNOR U3190 ( .A(n18237), .B(n18236), .Z(n18238) );
  NAND U3191 ( .A(n14174), .B(n14175), .Z(n1323) );
  NAND U3192 ( .A(n14173), .B(n14734), .Z(n1324) );
  NAND U3193 ( .A(n1323), .B(n1324), .Z(n14293) );
  XNOR U3194 ( .A(n14551), .B(n14550), .Z(n14528) );
  XNOR U3195 ( .A(n14499), .B(n14498), .Z(n14522) );
  XNOR U3196 ( .A(n14513), .B(n14512), .Z(n14515) );
  XOR U3197 ( .A(n14993), .B(n14992), .Z(n15037) );
  XOR U3198 ( .A(n15096), .B(n15095), .Z(n15084) );
  NAND U3199 ( .A(n15046), .B(n15047), .Z(n1325) );
  NANDN U3200 ( .A(n15049), .B(n15048), .Z(n1326) );
  NAND U3201 ( .A(n1325), .B(n1326), .Z(n15075) );
  XNOR U3202 ( .A(n15272), .B(n15271), .Z(n15274) );
  XNOR U3203 ( .A(n15280), .B(n15279), .Z(n15231) );
  NAND U3204 ( .A(n15119), .B(n15120), .Z(n1327) );
  NANDN U3205 ( .A(n15122), .B(n15121), .Z(n1328) );
  NAND U3206 ( .A(n1327), .B(n1328), .Z(n15236) );
  XNOR U3207 ( .A(n15569), .B(n15568), .Z(n15570) );
  XNOR U3208 ( .A(n15514), .B(n15513), .Z(n15516) );
  XNOR U3209 ( .A(n15687), .B(n15686), .Z(n15689) );
  XNOR U3210 ( .A(n15737), .B(n15736), .Z(n15738) );
  NAND U3211 ( .A(n15563), .B(n15564), .Z(n1329) );
  NANDN U3212 ( .A(n15566), .B(n15565), .Z(n1330) );
  AND U3213 ( .A(n1329), .B(n1330), .Z(n15626) );
  NAND U3214 ( .A(n15545), .B(n15546), .Z(n1331) );
  NANDN U3215 ( .A(n15548), .B(n15547), .Z(n1332) );
  AND U3216 ( .A(n1331), .B(n1332), .Z(n15621) );
  NAND U3217 ( .A(n15557), .B(n15556), .Z(n1333) );
  NAND U3218 ( .A(n15555), .B(n15554), .Z(n1334) );
  AND U3219 ( .A(n1333), .B(n1334), .Z(n15670) );
  NAND U3220 ( .A(n15491), .B(n15492), .Z(n1335) );
  NANDN U3221 ( .A(n15494), .B(n15493), .Z(n1336) );
  AND U3222 ( .A(n1335), .B(n1336), .Z(n15666) );
  NAND U3223 ( .A(n11282), .B(n11281), .Z(n1337) );
  NAND U3224 ( .A(n11395), .B(n12847), .Z(n1338) );
  AND U3225 ( .A(n1337), .B(n1338), .Z(n11339) );
  XOR U3226 ( .A(n11410), .B(n11409), .Z(n11444) );
  XNOR U3227 ( .A(n11429), .B(n11428), .Z(n11430) );
  XNOR U3228 ( .A(n11501), .B(n11500), .Z(n11558) );
  XNOR U3229 ( .A(n11703), .B(n11702), .Z(n11775) );
  XNOR U3230 ( .A(n11747), .B(n11746), .Z(n11770) );
  XNOR U3231 ( .A(n11753), .B(n11752), .Z(n11763) );
  XOR U3232 ( .A(n11849), .B(n11848), .Z(n11886) );
  XNOR U3233 ( .A(n11891), .B(n11890), .Z(n11892) );
  XNOR U3234 ( .A(n11879), .B(n11878), .Z(n11881) );
  XNOR U3235 ( .A(n12258), .B(n12257), .Z(n12214) );
  AND U3236 ( .A(n12679), .B(o[121]), .Z(n12853) );
  XNOR U3237 ( .A(n8252), .B(n8251), .Z(n8253) );
  XNOR U3238 ( .A(n8225), .B(n8224), .Z(n8227) );
  XOR U3239 ( .A(n8247), .B(n8248), .Z(n8232) );
  XNOR U3240 ( .A(n8613), .B(n8612), .Z(n8615) );
  XNOR U3241 ( .A(n8902), .B(n8901), .Z(n8949) );
  XNOR U3242 ( .A(n8928), .B(n8927), .Z(n8895) );
  XNOR U3243 ( .A(n8940), .B(n8939), .Z(n8889) );
  XNOR U3244 ( .A(n9039), .B(n9038), .Z(n9040) );
  XNOR U3245 ( .A(n9102), .B(n9101), .Z(n9052) );
  XNOR U3246 ( .A(n9058), .B(n9057), .Z(n9094) );
  XOR U3247 ( .A(n9019), .B(n9018), .Z(n9089) );
  XNOR U3248 ( .A(n9327), .B(n9326), .Z(n9283) );
  XNOR U3249 ( .A(n9434), .B(n9433), .Z(n9490) );
  NAND U3250 ( .A(n9547), .B(n9546), .Z(n1339) );
  NAND U3251 ( .A(n9687), .B(n9545), .Z(n1340) );
  NAND U3252 ( .A(n1339), .B(n1340), .Z(n9711) );
  XNOR U3253 ( .A(n9913), .B(n9912), .Z(n9914) );
  XNOR U3254 ( .A(n9925), .B(n9924), .Z(n9927) );
  XOR U3255 ( .A(n10096), .B(n10095), .Z(n10106) );
  XNOR U3256 ( .A(n5055), .B(o[40]), .Z(n5049) );
  XNOR U3257 ( .A(n5391), .B(o[45]), .Z(n5379) );
  XNOR U3258 ( .A(n5471), .B(n5750), .Z(n5480) );
  XNOR U3259 ( .A(n5386), .B(n6395), .Z(n5369) );
  XNOR U3260 ( .A(n5486), .B(n5485), .Z(n5488) );
  XNOR U3261 ( .A(n5462), .B(n5461), .Z(n5434) );
  XOR U3262 ( .A(n5527), .B(n5526), .Z(n5561) );
  XNOR U3263 ( .A(n5624), .B(n5623), .Z(n5680) );
  XNOR U3264 ( .A(n5825), .B(n5824), .Z(n5897) );
  XNOR U3265 ( .A(n5869), .B(n5868), .Z(n5892) );
  XNOR U3266 ( .A(n5875), .B(n5874), .Z(n5885) );
  XNOR U3267 ( .A(n6115), .B(n6114), .Z(n6117) );
  XNOR U3268 ( .A(n6078), .B(n6077), .Z(n6080) );
  XOR U3269 ( .A(n5991), .B(n5990), .Z(n6008) );
  XNOR U3270 ( .A(n6013), .B(n6012), .Z(n6014) );
  XNOR U3271 ( .A(n6001), .B(n6000), .Z(n6003) );
  XNOR U3272 ( .A(n6378), .B(n6377), .Z(n6336) );
  NAND U3273 ( .A(n6613), .B(n6614), .Z(n1341) );
  NANDN U3274 ( .A(n6616), .B(n6615), .Z(n1342) );
  NAND U3275 ( .A(n1341), .B(n1342), .Z(n6759) );
  NAND U3276 ( .A(n6453), .B(n6452), .Z(n1343) );
  NANDN U3277 ( .A(n6451), .B(n6450), .Z(n1344) );
  NAND U3278 ( .A(n1343), .B(n1344), .Z(n6586) );
  XNOR U3279 ( .A(n6941), .B(n6942), .Z(n6921) );
  XNOR U3280 ( .A(n6952), .B(n6951), .Z(n6953) );
  XOR U3281 ( .A(n6948), .B(n6947), .Z(n6878) );
  XNOR U3282 ( .A(n7249), .B(n7427), .Z(n7250) );
  XNOR U3283 ( .A(n2256), .B(n2255), .Z(n2257) );
  XNOR U3284 ( .A(n2318), .B(o[11]), .Z(n2299) );
  XNOR U3285 ( .A(n2695), .B(n2694), .Z(n2697) );
  XNOR U3286 ( .A(n3021), .B(n3020), .Z(n3069) );
  XNOR U3287 ( .A(n3141), .B(n3140), .Z(n3177) );
  XOR U3288 ( .A(n3118), .B(n3117), .Z(n3172) );
  XNOR U3289 ( .A(n3263), .B(n3262), .Z(n3265) );
  XNOR U3290 ( .A(n3410), .B(n3409), .Z(n3366) );
  XNOR U3291 ( .A(n3708), .B(n3707), .Z(n3710) );
  XNOR U3292 ( .A(n3662), .B(n3661), .Z(n3612) );
  XNOR U3293 ( .A(n3796), .B(n3795), .Z(n3797) );
  XNOR U3294 ( .A(n4008), .B(n4007), .Z(n4009) );
  XOR U3295 ( .A(n45576), .B(n46382), .Z(n45578) );
  XOR U3296 ( .A(n45773), .B(n45772), .Z(n45775) );
  XNOR U3297 ( .A(n46341), .B(n46340), .Z(n46342) );
  XOR U3298 ( .A(n46557), .B(n46556), .Z(n46561) );
  XNOR U3299 ( .A(n47151), .B(n47150), .Z(n47152) );
  XNOR U3300 ( .A(n47355), .B(n47354), .Z(n47347) );
  XNOR U3301 ( .A(n47637), .B(n47636), .Z(n47638) );
  XNOR U3302 ( .A(n47643), .B(n47642), .Z(n47644) );
  NAND U3303 ( .A(n47635), .B(n47634), .Z(n1345) );
  NANDN U3304 ( .A(n47633), .B(n47632), .Z(n1346) );
  NAND U3305 ( .A(n1345), .B(n1346), .Z(n47798) );
  NAND U3306 ( .A(n47555), .B(n47554), .Z(n1347) );
  NAND U3307 ( .A(n47760), .B(n47553), .Z(n1348) );
  AND U3308 ( .A(n1347), .B(n1348), .Z(n47721) );
  XNOR U3309 ( .A(n48159), .B(n47932), .Z(n47933) );
  XNOR U3310 ( .A(n47750), .B(n47749), .Z(n47724) );
  NAND U3311 ( .A(n42812), .B(n42811), .Z(n1349) );
  NAND U3312 ( .A(n42810), .B(n42991), .Z(n1350) );
  NAND U3313 ( .A(n1349), .B(n1350), .Z(n42842) );
  XOR U3314 ( .A(n42890), .B(n42889), .Z(n42892) );
  XOR U3315 ( .A(n44241), .B(n44240), .Z(n44246) );
  XNOR U3316 ( .A(n44438), .B(n44437), .Z(n44307) );
  XNOR U3317 ( .A(n44563), .B(n44562), .Z(n44557) );
  XNOR U3318 ( .A(n44601), .B(n44600), .Z(n44469) );
  XNOR U3319 ( .A(n44828), .B(n45032), .Z(n44829) );
  XNOR U3320 ( .A(n44806), .B(n44805), .Z(n44807) );
  XNOR U3321 ( .A(n44728), .B(n44727), .Z(n44682) );
  XNOR U3322 ( .A(n44717), .B(n44716), .Z(n44678) );
  NAND U3323 ( .A(n44710), .B(n44711), .Z(n1351) );
  NANDN U3324 ( .A(n44713), .B(n44712), .Z(n1352) );
  AND U3325 ( .A(n1351), .B(n1352), .Z(n44861) );
  XNOR U3326 ( .A(n44907), .B(n44906), .Z(n44909) );
  XNOR U3327 ( .A(n44834), .B(n44833), .Z(n44835) );
  XNOR U3328 ( .A(n45076), .B(n45075), .Z(n45078) );
  XNOR U3329 ( .A(n45082), .B(n45081), .Z(n45083) );
  XNOR U3330 ( .A(n44839), .B(o[476]), .Z(n44871) );
  XNOR U3331 ( .A(n44865), .B(n44864), .Z(n44866) );
  XOR U3332 ( .A(n40017), .B(n40016), .Z(n40011) );
  XNOR U3333 ( .A(n40088), .B(n40087), .Z(n40090) );
  XNOR U3334 ( .A(n40846), .B(n40845), .Z(n40847) );
  XOR U3335 ( .A(n41354), .B(n41353), .Z(n41359) );
  XNOR U3336 ( .A(n41549), .B(n41548), .Z(n41541) );
  NAND U3337 ( .A(n41637), .B(n41636), .Z(n1353) );
  NAND U3338 ( .A(n41635), .B(n41634), .Z(n1354) );
  AND U3339 ( .A(n1353), .B(n1354), .Z(n41839) );
  XNOR U3340 ( .A(n42158), .B(n42157), .Z(n42175) );
  XNOR U3341 ( .A(n42101), .B(n42100), .Z(n42189) );
  NAND U3342 ( .A(n41748), .B(n41747), .Z(n1355) );
  NAND U3343 ( .A(n41746), .B(n41745), .Z(n1356) );
  AND U3344 ( .A(n1355), .B(n1356), .Z(n41995) );
  XOR U3345 ( .A(n36933), .B(n37721), .Z(n36935) );
  XNOR U3346 ( .A(n37470), .B(n37469), .Z(n37472) );
  XOR U3347 ( .A(n37466), .B(n37465), .Z(n37458) );
  XOR U3348 ( .A(n37538), .B(n37537), .Z(n37494) );
  NAND U3349 ( .A(n37624), .B(n37623), .Z(n1357) );
  NAND U3350 ( .A(n37622), .B(n37621), .Z(n1358) );
  AND U3351 ( .A(n1357), .B(n1358), .Z(n37753) );
  XNOR U3352 ( .A(n37742), .B(n37741), .Z(n37761) );
  XNOR U3353 ( .A(n38000), .B(n37999), .Z(n38001) );
  XNOR U3354 ( .A(n38402), .B(n38401), .Z(n38388) );
  XNOR U3355 ( .A(n38691), .B(n38690), .Z(n38694) );
  XNOR U3356 ( .A(n38898), .B(n38897), .Z(n38900) );
  XNOR U3357 ( .A(n38912), .B(n38911), .Z(n38994) );
  XNOR U3358 ( .A(n38906), .B(n38905), .Z(n38988) );
  NAND U3359 ( .A(n38930), .B(n38929), .Z(n1359) );
  NANDN U3360 ( .A(n38928), .B(n38927), .Z(n1360) );
  NAND U3361 ( .A(n1359), .B(n1360), .Z(n39091) );
  NAND U3362 ( .A(n39072), .B(n39071), .Z(n1361) );
  NAND U3363 ( .A(n39069), .B(n39070), .Z(n1362) );
  NAND U3364 ( .A(n1361), .B(n1362), .Z(n39283) );
  XNOR U3365 ( .A(n39258), .B(n39257), .Z(n39277) );
  AND U3366 ( .A(n39263), .B(o[413]), .Z(n39436) );
  XOR U3367 ( .A(n34101), .B(n34897), .Z(n34103) );
  XOR U3368 ( .A(n34300), .B(n34299), .Z(n34302) );
  NAND U3369 ( .A(n34529), .B(n34528), .Z(n1363) );
  NANDN U3370 ( .A(n34527), .B(n34906), .Z(n1364) );
  AND U3371 ( .A(n1363), .B(n1364), .Z(n34632) );
  XNOR U3372 ( .A(n34697), .B(n34696), .Z(n34698) );
  XNOR U3373 ( .A(n35445), .B(n35444), .Z(n35446) );
  XNOR U3374 ( .A(n35891), .B(n35890), .Z(n35894) );
  XNOR U3375 ( .A(n35916), .B(n35915), .Z(n35910) );
  NAND U3376 ( .A(n36236), .B(n36235), .Z(n1365) );
  NAND U3377 ( .A(n36233), .B(n36234), .Z(n1366) );
  NAND U3378 ( .A(n1365), .B(n1366), .Z(n36464) );
  XNOR U3379 ( .A(n36628), .B(n36627), .Z(n36626) );
  NAND U3380 ( .A(n36428), .B(n36427), .Z(n1367) );
  NAND U3381 ( .A(n36426), .B(n36656), .Z(n1368) );
  AND U3382 ( .A(n1367), .B(n1368), .Z(n36632) );
  XNOR U3383 ( .A(n36282), .B(n36281), .Z(n36283) );
  NAND U3384 ( .A(n36113), .B(n36114), .Z(n1369) );
  NANDN U3385 ( .A(n36116), .B(n36115), .Z(n1370) );
  NAND U3386 ( .A(n1369), .B(n1370), .Z(n36277) );
  XNOR U3387 ( .A(n31102), .B(o[326]), .Z(n31094) );
  XNOR U3388 ( .A(n31223), .B(o[329]), .Z(n31215) );
  NAND U3389 ( .A(n31474), .B(n31473), .Z(n1371) );
  NAND U3390 ( .A(n31472), .B(n31471), .Z(n1372) );
  AND U3391 ( .A(n1371), .B(n1372), .Z(n31530) );
  XNOR U3392 ( .A(n31671), .B(n31670), .Z(n31673) );
  NAND U3393 ( .A(n31534), .B(n31535), .Z(n1373) );
  NANDN U3394 ( .A(n31537), .B(n31536), .Z(n1374) );
  NAND U3395 ( .A(n1373), .B(n1374), .Z(n31660) );
  XNOR U3396 ( .A(n31708), .B(n31707), .Z(n31750) );
  XOR U3397 ( .A(n32101), .B(n32100), .Z(n32105) );
  XNOR U3398 ( .A(n32228), .B(n32227), .Z(n32229) );
  XOR U3399 ( .A(n32218), .B(n32217), .Z(n32222) );
  XNOR U3400 ( .A(n32385), .B(n32384), .Z(n32386) );
  XNOR U3401 ( .A(n32626), .B(n32625), .Z(n32627) );
  XNOR U3402 ( .A(n32634), .B(n32633), .Z(n32620) );
  XNOR U3403 ( .A(n32671), .B(n32670), .Z(n32664) );
  XOR U3404 ( .A(n33174), .B(n33173), .Z(n33204) );
  XNOR U3405 ( .A(n33145), .B(n33144), .Z(n33246) );
  XOR U3406 ( .A(n33258), .B(n33257), .Z(n33260) );
  XOR U3407 ( .A(n28412), .B(n28411), .Z(n28414) );
  XNOR U3408 ( .A(n28572), .B(n28571), .Z(n28520) );
  XNOR U3409 ( .A(n28480), .B(n28479), .Z(n28501) );
  XOR U3410 ( .A(n29188), .B(n29187), .Z(n29192) );
  XNOR U3411 ( .A(n29890), .B(n29889), .Z(n29893) );
  XNOR U3412 ( .A(n30149), .B(n30148), .Z(n30155) );
  XOR U3413 ( .A(n30249), .B(n30248), .Z(n30267) );
  XNOR U3414 ( .A(n30594), .B(n30593), .Z(n30643) );
  XNOR U3415 ( .A(n30891), .B(n30890), .Z(n30888) );
  XNOR U3416 ( .A(n25347), .B(n25346), .Z(n25348) );
  XNOR U3417 ( .A(n25560), .B(n26142), .Z(n25539) );
  XNOR U3418 ( .A(n25638), .B(n25637), .Z(n25586) );
  XNOR U3419 ( .A(n25813), .B(n25812), .Z(n25815) );
  XOR U3420 ( .A(n25809), .B(n25808), .Z(n25801) );
  XNOR U3421 ( .A(n25873), .B(n25872), .Z(n25874) );
  XNOR U3422 ( .A(n25879), .B(n25878), .Z(n25881) );
  XNOR U3423 ( .A(n26103), .B(n26102), .Z(n26105) );
  XNOR U3424 ( .A(n26099), .B(n26098), .Z(n26035) );
  XNOR U3425 ( .A(n26849), .B(n26848), .Z(n26851) );
  XNOR U3426 ( .A(n26919), .B(n26918), .Z(n26921) );
  XNOR U3427 ( .A(n27182), .B(n27181), .Z(n27176) );
  XNOR U3428 ( .A(n27220), .B(n27219), .Z(n27087) );
  XOR U3429 ( .A(n27293), .B(n27292), .Z(n27323) );
  XOR U3430 ( .A(n27377), .B(n27376), .Z(n27379) );
  XNOR U3431 ( .A(n22885), .B(n22884), .Z(n22876) );
  XOR U3432 ( .A(n22973), .B(n22972), .Z(n22988) );
  XOR U3433 ( .A(n23095), .B(n23094), .Z(n23010) );
  XNOR U3434 ( .A(n23333), .B(n23332), .Z(n23334) );
  XOR U3435 ( .A(n23961), .B(n23960), .Z(n23966) );
  XNOR U3436 ( .A(n23900), .B(n23899), .Z(n23894) );
  XNOR U3437 ( .A(n24160), .B(n24159), .Z(n24161) );
  XNOR U3438 ( .A(n24479), .B(n24478), .Z(n24355) );
  XNOR U3439 ( .A(n24459), .B(n24458), .Z(n24460) );
  XNOR U3440 ( .A(n24567), .B(n24566), .Z(n24568) );
  XNOR U3441 ( .A(n24580), .B(n24579), .Z(n24581) );
  XNOR U3442 ( .A(n24496), .B(n24495), .Z(n24497) );
  XNOR U3443 ( .A(n19707), .B(n19706), .Z(n19708) );
  XNOR U3444 ( .A(n19714), .B(n19713), .Z(n19715) );
  XOR U3445 ( .A(n19811), .B(n19812), .Z(n19796) );
  NAND U3446 ( .A(n19860), .B(n19859), .Z(n1375) );
  NAND U3447 ( .A(n19858), .B(n19857), .Z(n1376) );
  AND U3448 ( .A(n1375), .B(n1376), .Z(n19925) );
  XNOR U3449 ( .A(n20065), .B(n20064), .Z(n20067) );
  NAND U3450 ( .A(n19929), .B(n19930), .Z(n1377) );
  NANDN U3451 ( .A(n19932), .B(n19931), .Z(n1378) );
  NAND U3452 ( .A(n1377), .B(n1378), .Z(n20054) );
  XNOR U3453 ( .A(n20134), .B(n20133), .Z(n20096) );
  XNOR U3454 ( .A(n20368), .B(n20367), .Z(n20369) );
  XNOR U3455 ( .A(n20374), .B(n20373), .Z(n20376) );
  XNOR U3456 ( .A(n20462), .B(n20461), .Z(n20472) );
  XOR U3457 ( .A(n20484), .B(n20483), .Z(n20486) );
  XNOR U3458 ( .A(n20766), .B(n20765), .Z(n20767) );
  XNOR U3459 ( .A(n20999), .B(n20998), .Z(n21017) );
  XNOR U3460 ( .A(n21433), .B(n21432), .Z(n21388) );
  AND U3461 ( .A(n21533), .B(n21532), .Z(n1379) );
  AND U3462 ( .A(n21954), .B(y[7875]), .Z(n1380) );
  NAND U3463 ( .A(x[500]), .B(n1380), .Z(n1381) );
  NANDN U3464 ( .A(n1379), .B(n1381), .Z(n21713) );
  NAND U3465 ( .A(n21537), .B(n21536), .Z(n1382) );
  NAND U3466 ( .A(n21534), .B(n21535), .Z(n1383) );
  NAND U3467 ( .A(n1382), .B(n1383), .Z(n21709) );
  NAND U3468 ( .A(n21502), .B(n21501), .Z(n1384) );
  NAND U3469 ( .A(n21499), .B(n21500), .Z(n1385) );
  NAND U3470 ( .A(n1384), .B(n1385), .Z(n21681) );
  NAND U3471 ( .A(n21520), .B(n21521), .Z(n1386) );
  NANDN U3472 ( .A(n21523), .B(n21522), .Z(n1387) );
  NAND U3473 ( .A(n1386), .B(n1387), .Z(n21685) );
  XNOR U3474 ( .A(n16727), .B(o[169]), .Z(n16719) );
  XNOR U3475 ( .A(n17213), .B(n17212), .Z(n17214) );
  XNOR U3476 ( .A(n17434), .B(n17433), .Z(n17507) );
  XNOR U3477 ( .A(n17479), .B(n17478), .Z(n17502) );
  XNOR U3478 ( .A(n17485), .B(n17484), .Z(n17495) );
  NAND U3479 ( .A(n17371), .B(n17370), .Z(n1388) );
  NAND U3480 ( .A(n17369), .B(n17368), .Z(n1389) );
  AND U3481 ( .A(n1388), .B(n1389), .Z(n17490) );
  XOR U3482 ( .A(n17742), .B(n17741), .Z(n17746) );
  XNOR U3483 ( .A(n17752), .B(n17751), .Z(n17753) );
  NAND U3484 ( .A(n17895), .B(n17896), .Z(n1390) );
  NAND U3485 ( .A(n17893), .B(n17894), .Z(n1391) );
  NAND U3486 ( .A(n1390), .B(n1391), .Z(n18101) );
  NAND U3487 ( .A(n17963), .B(n17964), .Z(n1392) );
  NAND U3488 ( .A(n17961), .B(n17962), .Z(n1393) );
  NAND U3489 ( .A(n1392), .B(n1393), .Z(n18112) );
  XNOR U3490 ( .A(n18283), .B(n18282), .Z(n18285) );
  XNOR U3491 ( .A(n18406), .B(n18405), .Z(n18407) );
  XOR U3492 ( .A(n18636), .B(n18635), .Z(n18666) );
  XNOR U3493 ( .A(n19135), .B(n19136), .Z(n19202) );
  XNOR U3494 ( .A(n19209), .B(n19208), .Z(n19207) );
  XNOR U3495 ( .A(n18607), .B(n18606), .Z(n18708) );
  XOR U3496 ( .A(n14099), .B(n14098), .Z(n14093) );
  XNOR U3497 ( .A(n14158), .B(n14157), .Z(n14160) );
  NAND U3498 ( .A(n14292), .B(n14291), .Z(n1394) );
  NANDN U3499 ( .A(n14290), .B(n14647), .Z(n1395) );
  AND U3500 ( .A(n1394), .B(n1395), .Z(n14387) );
  NAND U3501 ( .A(n14350), .B(n14349), .Z(n1396) );
  NANDN U3502 ( .A(n14348), .B(n14347), .Z(n1397) );
  NAND U3503 ( .A(n1396), .B(n1397), .Z(n14441) );
  XOR U3504 ( .A(n14703), .B(n14702), .Z(n14705) );
  XNOR U3505 ( .A(n15587), .B(n15586), .Z(n15589) );
  XNOR U3506 ( .A(n15743), .B(n15742), .Z(n15744) );
  XNOR U3507 ( .A(n16390), .B(n16389), .Z(n16387) );
  AND U3508 ( .A(n16144), .B(o[157]), .Z(n16374) );
  XOR U3509 ( .A(n11039), .B(n11038), .Z(n11066) );
  XOR U3510 ( .A(n11184), .B(n11185), .Z(n11169) );
  NAND U3511 ( .A(n11260), .B(n11259), .Z(n1398) );
  NAND U3512 ( .A(n11258), .B(n11257), .Z(n1399) );
  AND U3513 ( .A(n1398), .B(n1399), .Z(n11309) );
  XNOR U3514 ( .A(n11449), .B(n11448), .Z(n11450) );
  XOR U3515 ( .A(n11497), .B(n11496), .Z(n11513) );
  XOR U3516 ( .A(n11665), .B(n11664), .Z(n11580) );
  XNOR U3517 ( .A(n12588), .B(n12587), .Z(n12589) );
  XOR U3518 ( .A(n12924), .B(n12923), .Z(n12954) );
  XNOR U3519 ( .A(n12897), .B(n12896), .Z(n12996) );
  XOR U3520 ( .A(n13008), .B(n13007), .Z(n13010) );
  XOR U3521 ( .A(n12992), .B(n12991), .Z(n13002) );
  XNOR U3522 ( .A(n8183), .B(n8182), .Z(n8206) );
  XNOR U3523 ( .A(n8188), .B(n8187), .Z(n8202) );
  XNOR U3524 ( .A(n8311), .B(n8310), .Z(n8303) );
  XNOR U3525 ( .A(n8770), .B(n8769), .Z(n8772) );
  XOR U3526 ( .A(n8979), .B(n8978), .Z(n8981) );
  XNOR U3527 ( .A(n8985), .B(n8984), .Z(n8986) );
  XNOR U3528 ( .A(n9669), .B(n9668), .Z(n9671) );
  XNOR U3529 ( .A(n5118), .B(n5117), .Z(n5119) );
  XNOR U3530 ( .A(n5188), .B(n5187), .Z(n5189) );
  XNOR U3531 ( .A(n5208), .B(n5207), .Z(n5209) );
  XOR U3532 ( .A(n5301), .B(n5302), .Z(n5286) );
  XNOR U3533 ( .A(n5580), .B(n5579), .Z(n5571) );
  XOR U3534 ( .A(n5620), .B(n5619), .Z(n5635) );
  XOR U3535 ( .A(n5787), .B(n5786), .Z(n5702) );
  XNOR U3536 ( .A(n6133), .B(n6132), .Z(n6134) );
  XOR U3537 ( .A(n7077), .B(n7076), .Z(n7095) );
  NAND U3538 ( .A(n6959), .B(n6960), .Z(n1400) );
  NAND U3539 ( .A(n6957), .B(n6958), .Z(n1401) );
  NAND U3540 ( .A(n1400), .B(n1401), .Z(n7027) );
  XNOR U3541 ( .A(n7022), .B(n7021), .Z(n7023) );
  XNOR U3542 ( .A(n7262), .B(n7261), .Z(n7263) );
  XNOR U3543 ( .A(n7255), .B(n7254), .Z(n7256) );
  XNOR U3544 ( .A(n7689), .B(n7451), .Z(n7452) );
  XNOR U3545 ( .A(n2198), .B(n2197), .Z(n2199) );
  XOR U3546 ( .A(n2358), .B(n2357), .Z(n2352) );
  XNOR U3547 ( .A(n2472), .B(n2471), .Z(n2481) );
  XNOR U3548 ( .A(n2441), .B(n2440), .Z(n2433) );
  XNOR U3549 ( .A(n2507), .B(n2506), .Z(n2508) );
  XNOR U3550 ( .A(n2882), .B(n2881), .Z(n2884) );
  NAND U3551 ( .A(n2890), .B(n2889), .Z(n1402) );
  NANDN U3552 ( .A(n2888), .B(n2887), .Z(n1403) );
  NAND U3553 ( .A(n1402), .B(n1403), .Z(n2991) );
  NAND U3554 ( .A(n2936), .B(n2937), .Z(n1404) );
  NAND U3555 ( .A(n2934), .B(n2935), .Z(n1405) );
  NAND U3556 ( .A(n1404), .B(n1405), .Z(n3003) );
  XNOR U3557 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U3558 ( .A(n3124), .B(n3123), .Z(n3128) );
  XNOR U3559 ( .A(n3760), .B(n3759), .Z(n3761) );
  XNOR U3560 ( .A(n4042), .B(n4041), .Z(n3995) );
  NAND U3561 ( .A(n4107), .B(n4108), .Z(n1406) );
  NANDN U3562 ( .A(n4110), .B(n4109), .Z(n1407) );
  NAND U3563 ( .A(n1406), .B(n1407), .Z(n4347) );
  XNOR U3564 ( .A(n4365), .B(n4364), .Z(n4366) );
  XNOR U3565 ( .A(n4353), .B(n4352), .Z(n4354) );
  NAND U3566 ( .A(n3926), .B(n3925), .Z(n1408) );
  NAND U3567 ( .A(n3924), .B(n3923), .Z(n1409) );
  AND U3568 ( .A(n1408), .B(n1409), .Z(n4096) );
  XNOR U3569 ( .A(n4152), .B(n4151), .Z(n4089) );
  XNOR U3570 ( .A(n45544), .B(n45543), .Z(n45555) );
  NAND U3571 ( .A(n45650), .B(n45649), .Z(n1410) );
  NANDN U3572 ( .A(n46251), .B(n45994), .Z(n1411) );
  AND U3573 ( .A(n1410), .B(n1411), .Z(n45662) );
  XOR U3574 ( .A(n46321), .B(n46320), .Z(n46236) );
  XNOR U3575 ( .A(n47099), .B(n47098), .Z(n47100) );
  NAND U3576 ( .A(n47387), .B(n47386), .Z(n1412) );
  NANDN U3577 ( .A(n47385), .B(n47384), .Z(n1413) );
  AND U3578 ( .A(n1412), .B(n1413), .Z(n47531) );
  NAND U3579 ( .A(n47509), .B(n47510), .Z(n1414) );
  NANDN U3580 ( .A(n47512), .B(n47511), .Z(n1415) );
  AND U3581 ( .A(n1414), .B(n1415), .Z(n47523) );
  NAND U3582 ( .A(n47704), .B(n47703), .Z(n1416) );
  NAND U3583 ( .A(n47702), .B(n47701), .Z(n1417) );
  AND U3584 ( .A(n1416), .B(n1417), .Z(n47962) );
  NAND U3585 ( .A(n47983), .B(n47984), .Z(n1418) );
  NANDN U3586 ( .A(n47986), .B(n47985), .Z(n1419) );
  AND U3587 ( .A(n1418), .B(n1419), .Z(n48204) );
  NAND U3588 ( .A(n48169), .B(n48168), .Z(n1420) );
  NAND U3589 ( .A(n48167), .B(n48166), .Z(n1421) );
  AND U3590 ( .A(n1420), .B(n1421), .Z(n48177) );
  XOR U3591 ( .A(n48026), .B(n48027), .Z(n48028) );
  XOR U3592 ( .A(n48033), .B(n48032), .Z(n48034) );
  XNOR U3593 ( .A(n42652), .B(n42651), .Z(n42653) );
  XOR U3594 ( .A(n43178), .B(n43177), .Z(n43180) );
  NAND U3595 ( .A(n43221), .B(n43222), .Z(n1422) );
  NANDN U3596 ( .A(n43224), .B(n43223), .Z(n1423) );
  NAND U3597 ( .A(n1422), .B(n1423), .Z(n43312) );
  XNOR U3598 ( .A(n43521), .B(n43520), .Z(n43623) );
  XNOR U3599 ( .A(n43430), .B(n43429), .Z(n43423) );
  XNOR U3600 ( .A(n44466), .B(n44465), .Z(n44460) );
  XOR U3601 ( .A(n44752), .B(n44751), .Z(n44615) );
  XOR U3602 ( .A(n44921), .B(n44920), .Z(n44893) );
  NAND U3603 ( .A(n44677), .B(n44676), .Z(n1424) );
  NANDN U3604 ( .A(n44675), .B(n44674), .Z(n1425) );
  AND U3605 ( .A(n1424), .B(n1425), .Z(n44887) );
  XNOR U3606 ( .A(n44825), .B(n44824), .Z(n44904) );
  XNOR U3607 ( .A(n45046), .B(n45045), .Z(n45047) );
  XNOR U3608 ( .A(n45064), .B(n45063), .Z(n45066) );
  XNOR U3609 ( .A(n45312), .B(n45311), .Z(n45309) );
  XOR U3610 ( .A(n45142), .B(n45141), .Z(n45140) );
  XNOR U3611 ( .A(n44853), .B(n44852), .Z(n44855) );
  XNOR U3612 ( .A(n39754), .B(n39753), .Z(n39756) );
  NAND U3613 ( .A(n39671), .B(n39670), .Z(n1426) );
  XOR U3614 ( .A(n39671), .B(n39670), .Z(n1427) );
  NANDN U3615 ( .A(n39742), .B(n1427), .Z(n1428) );
  NAND U3616 ( .A(n1426), .B(n1428), .Z(n39713) );
  NAND U3617 ( .A(n39845), .B(n39844), .Z(n1429) );
  NANDN U3618 ( .A(n40475), .B(n40204), .Z(n1430) );
  AND U3619 ( .A(n1429), .B(n1430), .Z(n39861) );
  XOR U3620 ( .A(n40157), .B(n40156), .Z(n40159) );
  XNOR U3621 ( .A(n40734), .B(n40733), .Z(n40746) );
  XNOR U3622 ( .A(n40531), .B(n40530), .Z(n40524) );
  XOR U3623 ( .A(n40882), .B(n40881), .Z(n40875) );
  XNOR U3624 ( .A(n41294), .B(n41293), .Z(n41288) );
  XNOR U3625 ( .A(n41282), .B(n41281), .Z(n41411) );
  XOR U3626 ( .A(n41425), .B(n41424), .Z(n41427) );
  NAND U3627 ( .A(n41590), .B(n41589), .Z(n1431) );
  NAND U3628 ( .A(n41588), .B(n41587), .Z(n1432) );
  AND U3629 ( .A(n1431), .B(n1432), .Z(n41723) );
  NAND U3630 ( .A(n41712), .B(n41713), .Z(n1433) );
  NANDN U3631 ( .A(n41715), .B(n41714), .Z(n1434) );
  AND U3632 ( .A(n1433), .B(n1434), .Z(n41718) );
  XOR U3633 ( .A(n42257), .B(n42256), .Z(n42255) );
  XNOR U3634 ( .A(n42439), .B(n42438), .Z(n42437) );
  XNOR U3635 ( .A(n42094), .B(n42093), .Z(n42095) );
  XNOR U3636 ( .A(n37231), .B(n37230), .Z(n37233) );
  XNOR U3637 ( .A(n37780), .B(n37779), .Z(n37879) );
  NAND U3638 ( .A(n37757), .B(n37758), .Z(n1435) );
  NAND U3639 ( .A(n37755), .B(n37756), .Z(n1436) );
  NAND U3640 ( .A(n1435), .B(n1436), .Z(n37874) );
  XNOR U3641 ( .A(n38147), .B(n38146), .Z(n38148) );
  XNOR U3642 ( .A(n38141), .B(n38140), .Z(n38143) );
  XNOR U3643 ( .A(n38534), .B(n38533), .Z(n38540) );
  XNOR U3644 ( .A(n38892), .B(n38891), .Z(n38894) );
  XOR U3645 ( .A(n39027), .B(n39026), .Z(n39021) );
  XNOR U3646 ( .A(n39037), .B(n39036), .Z(n39038) );
  AND U3647 ( .A(n38967), .B(n38966), .Z(n1437) );
  AND U3648 ( .A(n39373), .B(y[8067]), .Z(n1438) );
  NAND U3649 ( .A(x[500]), .B(n1438), .Z(n1439) );
  NANDN U3650 ( .A(n1437), .B(n1439), .Z(n39141) );
  NAND U3651 ( .A(n38970), .B(n38971), .Z(n1440) );
  NAND U3652 ( .A(n38968), .B(n38969), .Z(n1441) );
  NAND U3653 ( .A(n1440), .B(n1441), .Z(n39137) );
  NAND U3654 ( .A(n38974), .B(n38975), .Z(n1442) );
  NAND U3655 ( .A(n38972), .B(n38973), .Z(n1443) );
  NAND U3656 ( .A(n1442), .B(n1443), .Z(n39131) );
  NAND U3657 ( .A(n39105), .B(n39106), .Z(n1444) );
  NAND U3658 ( .A(n39103), .B(n39104), .Z(n1445) );
  NAND U3659 ( .A(n1444), .B(n1445), .Z(n39270) );
  XNOR U3660 ( .A(n39332), .B(n39331), .Z(n39329) );
  XOR U3661 ( .A(n39468), .B(n39469), .Z(n39470) );
  NAND U3662 ( .A(n39087), .B(n39086), .Z(n1446) );
  NAND U3663 ( .A(n39084), .B(n39085), .Z(n1447) );
  NAND U3664 ( .A(n1446), .B(n1447), .Z(n39225) );
  XNOR U3665 ( .A(n39513), .B(n39512), .Z(n39510) );
  XOR U3666 ( .A(n39342), .B(n39341), .Z(n39340) );
  XNOR U3667 ( .A(n34071), .B(n34070), .Z(n34072) );
  XOR U3668 ( .A(n34734), .B(n34733), .Z(n34705) );
  XNOR U3669 ( .A(n35057), .B(n35056), .Z(n35058) );
  XNOR U3670 ( .A(n35766), .B(n35765), .Z(n35768) );
  XNOR U3671 ( .A(n36051), .B(n36050), .Z(n36052) );
  NAND U3672 ( .A(n36094), .B(n36095), .Z(n1448) );
  NAND U3673 ( .A(n36092), .B(n36093), .Z(n1449) );
  NAND U3674 ( .A(n1448), .B(n1449), .Z(n36269) );
  NAND U3675 ( .A(n36250), .B(n36249), .Z(n1450) );
  NAND U3676 ( .A(n36247), .B(n36248), .Z(n1451) );
  NAND U3677 ( .A(n1450), .B(n1451), .Z(n36413) );
  NAND U3678 ( .A(n36425), .B(n36424), .Z(n1452) );
  NAND U3679 ( .A(n36423), .B(n36613), .Z(n1453) );
  NAND U3680 ( .A(n1452), .B(n1453), .Z(n36532) );
  XOR U3681 ( .A(n36518), .B(n36517), .Z(n36516) );
  XOR U3682 ( .A(n36193), .B(n36192), .Z(n36187) );
  XNOR U3683 ( .A(n31115), .B(n31114), .Z(n31116) );
  XNOR U3684 ( .A(n31141), .B(n31140), .Z(n31143) );
  XNOR U3685 ( .A(n31180), .B(n31179), .Z(n31181) );
  XNOR U3686 ( .A(n31186), .B(n31185), .Z(n31187) );
  XOR U3687 ( .A(n31348), .B(n31347), .Z(n31350) );
  XNOR U3688 ( .A(n31802), .B(n31801), .Z(n31804) );
  XOR U3689 ( .A(n31796), .B(n31795), .Z(n31798) );
  XNOR U3690 ( .A(n32489), .B(n32488), .Z(n32380) );
  XNOR U3691 ( .A(n33125), .B(n33124), .Z(n33127) );
  XNOR U3692 ( .A(n33404), .B(n33403), .Z(n33406) );
  XNOR U3693 ( .A(n33289), .B(n33288), .Z(n33290) );
  XNOR U3694 ( .A(n33547), .B(n33546), .Z(n33577) );
  XOR U3695 ( .A(n33758), .B(n33595), .Z(n1454) );
  XNOR U3696 ( .A(n33596), .B(n1454), .Z(n33507) );
  XOR U3697 ( .A(n33663), .B(n33664), .Z(n33665) );
  XNOR U3698 ( .A(n33652), .B(n33651), .Z(n33649) );
  XNOR U3699 ( .A(n28221), .B(n28220), .Z(n28222) );
  XNOR U3700 ( .A(n28227), .B(n28226), .Z(n28228) );
  XNOR U3701 ( .A(n28586), .B(n28585), .Z(n28587) );
  XNOR U3702 ( .A(n29457), .B(n29456), .Z(n29459) );
  XNOR U3703 ( .A(n29451), .B(n29450), .Z(n29453) );
  XNOR U3704 ( .A(n29882), .B(n29881), .Z(n29884) );
  XNOR U3705 ( .A(n30194), .B(n30193), .Z(n30196) );
  XNOR U3706 ( .A(n30431), .B(n30430), .Z(n30432) );
  XOR U3707 ( .A(n30489), .B(n30488), .Z(n30459) );
  NAND U3708 ( .A(n30261), .B(n30260), .Z(n1455) );
  NANDN U3709 ( .A(n30259), .B(n30258), .Z(n1456) );
  AND U3710 ( .A(n1455), .B(n1456), .Z(n30452) );
  XOR U3711 ( .A(n30368), .B(n30367), .Z(n30471) );
  XNOR U3712 ( .A(n30475), .B(n30474), .Z(n30477) );
  XNOR U3713 ( .A(n30546), .B(n30545), .Z(n30547) );
  XNOR U3714 ( .A(n30885), .B(n30884), .Z(n30882) );
  XOR U3715 ( .A(n30709), .B(n30708), .Z(n30707) );
  XOR U3716 ( .A(n30721), .B(n30720), .Z(n30719) );
  XNOR U3717 ( .A(n25575), .B(n25574), .Z(n25577) );
  XNOR U3718 ( .A(n26221), .B(n26220), .Z(n26222) );
  OR U3719 ( .A(n26217), .B(n26216), .Z(n1457) );
  NAND U3720 ( .A(n26218), .B(n26219), .Z(n1458) );
  AND U3721 ( .A(n1457), .B(n1458), .Z(n26345) );
  XNOR U3722 ( .A(n26913), .B(n26912), .Z(n26915) );
  XNOR U3723 ( .A(n26786), .B(n26785), .Z(n26779) );
  XOR U3724 ( .A(n27385), .B(n27384), .Z(n27238) );
  XNOR U3725 ( .A(n27523), .B(n27522), .Z(n27525) );
  XNOR U3726 ( .A(n27706), .B(n27705), .Z(n27596) );
  XNOR U3727 ( .A(n27715), .B(n27716), .Z(n1459) );
  XNOR U3728 ( .A(n27717), .B(n1459), .Z(n27632) );
  XNOR U3729 ( .A(n27624), .B(n27623), .Z(n27625) );
  XNOR U3730 ( .A(n27648), .B(n27647), .Z(n27697) );
  XOR U3731 ( .A(n27710), .B(n27709), .Z(n27711) );
  XNOR U3732 ( .A(n27775), .B(n27774), .Z(n27772) );
  XNOR U3733 ( .A(n27408), .B(n27407), .Z(n27409) );
  XOR U3734 ( .A(n22324), .B(n22236), .Z(n1460) );
  NANDN U3735 ( .A(n22237), .B(n1460), .Z(n1461) );
  NAND U3736 ( .A(n22324), .B(n22236), .Z(n1462) );
  AND U3737 ( .A(n1461), .B(n1462), .Z(n22289) );
  XNOR U3738 ( .A(n22702), .B(n22701), .Z(n22704) );
  XNOR U3739 ( .A(n22959), .B(n22958), .Z(n22961) );
  XOR U3740 ( .A(n23089), .B(n23088), .Z(n23005) );
  XNOR U3741 ( .A(n23111), .B(n23110), .Z(n23217) );
  XNOR U3742 ( .A(n23466), .B(n23465), .Z(n23467) );
  XOR U3743 ( .A(n23718), .B(n23717), .Z(n23609) );
  XOR U3744 ( .A(n24038), .B(n24037), .Z(n24040) );
  XNOR U3745 ( .A(n24328), .B(n24327), .Z(n24330) );
  XNOR U3746 ( .A(n24344), .B(n24343), .Z(n24345) );
  NAND U3747 ( .A(n24456), .B(n24455), .Z(n1463) );
  NANDN U3748 ( .A(n24454), .B(n24453), .Z(n1464) );
  NAND U3749 ( .A(n1463), .B(n1464), .Z(n24600) );
  XNOR U3750 ( .A(n24678), .B(n24677), .Z(n24679) );
  XNOR U3751 ( .A(n24789), .B(n24788), .Z(n24765) );
  XNOR U3752 ( .A(n24757), .B(n24756), .Z(n24758) );
  XNOR U3753 ( .A(n24870), .B(n24724), .Z(n24725) );
  NAND U3754 ( .A(n24877), .B(n24799), .Z(n1465) );
  XOR U3755 ( .A(n24877), .B(n24799), .Z(n1466) );
  NANDN U3756 ( .A(n24798), .B(n1466), .Z(n1467) );
  NAND U3757 ( .A(n1465), .B(n1467), .Z(n25017) );
  XOR U3758 ( .A(n24975), .B(n24976), .Z(n24977) );
  XNOR U3759 ( .A(n24972), .B(n24971), .Z(n24969) );
  XNOR U3760 ( .A(n19442), .B(o[196]), .Z(n19444) );
  XNOR U3761 ( .A(n19540), .B(n19539), .Z(n19541) );
  XOR U3762 ( .A(n19675), .B(n19674), .Z(n19667) );
  XOR U3763 ( .A(n19765), .B(n19764), .Z(n19747) );
  XOR U3764 ( .A(n20192), .B(n20191), .Z(n20194) );
  XNOR U3765 ( .A(n20186), .B(n20185), .Z(n20188) );
  XNOR U3766 ( .A(n20490), .B(n20489), .Z(n20491) );
  XNOR U3767 ( .A(n20609), .B(n20608), .Z(n20613) );
  XOR U3768 ( .A(n20643), .B(n20642), .Z(n20636) );
  XOR U3769 ( .A(n20890), .B(n20889), .Z(n20892) );
  XNOR U3770 ( .A(n21190), .B(n21189), .Z(n21192) );
  NAND U3771 ( .A(n21497), .B(n21498), .Z(n1468) );
  NAND U3772 ( .A(n21495), .B(n21496), .Z(n1469) );
  NAND U3773 ( .A(n1468), .B(n1469), .Z(n21665) );
  NAND U3774 ( .A(n21661), .B(n21660), .Z(n1470) );
  NAND U3775 ( .A(n21658), .B(n21659), .Z(n1471) );
  NAND U3776 ( .A(n1470), .B(n1471), .Z(n21823) );
  XNOR U3777 ( .A(n22088), .B(n22087), .Z(n22086) );
  NAND U3778 ( .A(n21794), .B(n21793), .Z(n1472) );
  NAND U3779 ( .A(n21792), .B(n21942), .Z(n1473) );
  NAND U3780 ( .A(n1472), .B(n1473), .Z(n21930) );
  XOR U3781 ( .A(n22048), .B(n22047), .Z(n22046) );
  XOR U3782 ( .A(n21916), .B(n21915), .Z(n21914) );
  XOR U3783 ( .A(n21602), .B(n21601), .Z(n21596) );
  XNOR U3784 ( .A(n16706), .B(n16705), .Z(n16708) );
  XOR U3785 ( .A(n16877), .B(n16876), .Z(n16879) );
  XOR U3786 ( .A(n17203), .B(n17202), .Z(n17194) );
  XNOR U3787 ( .A(n17538), .B(n17537), .Z(n17634) );
  XNOR U3788 ( .A(n17774), .B(n17773), .Z(n17776) );
  NAND U3789 ( .A(n18108), .B(n18109), .Z(n1474) );
  NAND U3790 ( .A(n18106), .B(n18107), .Z(n1475) );
  NAND U3791 ( .A(n1474), .B(n1475), .Z(n18256) );
  XNOR U3792 ( .A(n18565), .B(n18564), .Z(n18566) );
  XNOR U3793 ( .A(n18587), .B(n18586), .Z(n18589) );
  XNOR U3794 ( .A(n18876), .B(n18875), .Z(n18878) );
  XOR U3795 ( .A(n18750), .B(n18749), .Z(n18744) );
  XNOR U3796 ( .A(n18973), .B(n18972), .Z(n18974) );
  XNOR U3797 ( .A(n18997), .B(n18996), .Z(n19045) );
  XOR U3798 ( .A(n19058), .B(n19057), .Z(n19060) );
  XNOR U3799 ( .A(n19125), .B(n19124), .Z(n19122) );
  XNOR U3800 ( .A(n18760), .B(n18759), .Z(n18761) );
  NAND U3801 ( .A(n14383), .B(n14384), .Z(n1476) );
  NANDN U3802 ( .A(n14386), .B(n14385), .Z(n1477) );
  NAND U3803 ( .A(n1476), .B(n1477), .Z(n14392) );
  XNOR U3804 ( .A(n14798), .B(n14797), .Z(n14799) );
  XNOR U3805 ( .A(n14914), .B(n14913), .Z(n14915) );
  NAND U3806 ( .A(n14951), .B(n14952), .Z(n1478) );
  NANDN U3807 ( .A(n14954), .B(n14953), .Z(n1479) );
  AND U3808 ( .A(n1478), .B(n1479), .Z(n15070) );
  XNOR U3809 ( .A(n15454), .B(n15453), .Z(n15455) );
  XNOR U3810 ( .A(n15330), .B(n15329), .Z(n15331) );
  XNOR U3811 ( .A(n15476), .B(n15475), .Z(n15478) );
  NAND U3812 ( .A(n15823), .B(n15824), .Z(n1480) );
  NANDN U3813 ( .A(n15826), .B(n15825), .Z(n1481) );
  AND U3814 ( .A(n1480), .B(n1481), .Z(n15978) );
  NAND U3815 ( .A(n15791), .B(n15790), .Z(n1482) );
  NAND U3816 ( .A(n15789), .B(n15788), .Z(n1483) );
  AND U3817 ( .A(n1482), .B(n1483), .Z(n15990) );
  XOR U3818 ( .A(n15910), .B(n15909), .Z(n15904) );
  NAND U3819 ( .A(n15958), .B(n15957), .Z(n1484) );
  NAND U3820 ( .A(n16117), .B(n15956), .Z(n1485) );
  AND U3821 ( .A(n1484), .B(n1485), .Z(n16167) );
  XOR U3822 ( .A(n16218), .B(n16217), .Z(n16216) );
  XOR U3823 ( .A(n16366), .B(n16365), .Z(n16364) );
  NAND U3824 ( .A(n15953), .B(n15954), .Z(n1486) );
  NAND U3825 ( .A(n15951), .B(n15952), .Z(n1487) );
  NAND U3826 ( .A(n1486), .B(n1487), .Z(n16115) );
  NAND U3827 ( .A(n15938), .B(n15937), .Z(n1488) );
  NAND U3828 ( .A(n15936), .B(n15935), .Z(n1489) );
  AND U3829 ( .A(n1488), .B(n1489), .Z(n16160) );
  XNOR U3830 ( .A(n16422), .B(n16421), .Z(n16419) );
  NAND U3831 ( .A(n16180), .B(n16181), .Z(n1490) );
  NANDN U3832 ( .A(n16183), .B(n16182), .Z(n1491) );
  AND U3833 ( .A(n1490), .B(n1491), .Z(n16414) );
  XOR U3834 ( .A(n16230), .B(n16229), .Z(n16228) );
  XNOR U3835 ( .A(n10888), .B(n10887), .Z(n10889) );
  XNOR U3836 ( .A(n10913), .B(n10912), .Z(n10915) );
  NAND U3837 ( .A(n11726), .B(n10934), .Z(n1492) );
  NANDN U3838 ( .A(n10936), .B(n10935), .Z(n1493) );
  NAND U3839 ( .A(n1492), .B(n1493), .Z(n10976) );
  XNOR U3840 ( .A(n11483), .B(n11482), .Z(n11485) );
  XNOR U3841 ( .A(n11463), .B(n11462), .Z(n11388) );
  XOR U3842 ( .A(n11659), .B(n11658), .Z(n11575) );
  XNOR U3843 ( .A(n11681), .B(n11680), .Z(n11787) );
  XNOR U3844 ( .A(n11911), .B(n11910), .Z(n11794) );
  XOR U3845 ( .A(n12051), .B(n12050), .Z(n12044) );
  XNOR U3846 ( .A(n12321), .B(n12320), .Z(n12305) );
  XNOR U3847 ( .A(n12582), .B(n12581), .Z(n12584) );
  NAND U3848 ( .A(n12823), .B(n12824), .Z(n1494) );
  NANDN U3849 ( .A(n12826), .B(n12825), .Z(n1495) );
  NAND U3850 ( .A(n1494), .B(n1495), .Z(n12878) );
  OR U3851 ( .A(n12740), .B(n12741), .Z(n1496) );
  NAND U3852 ( .A(n12743), .B(n12742), .Z(n1497) );
  NAND U3853 ( .A(n1496), .B(n1497), .Z(n12874) );
  XNOR U3854 ( .A(n13162), .B(n13161), .Z(n13164) );
  XNOR U3855 ( .A(n13192), .B(n13191), .Z(n13193) );
  XOR U3856 ( .A(n13232), .B(n13231), .Z(n13234) );
  XNOR U3857 ( .A(n13311), .B(n13310), .Z(n13312) );
  XOR U3858 ( .A(n13426), .B(n13425), .Z(n13424) );
  XOR U3859 ( .A(n13412), .B(n13411), .Z(n13410) );
  XNOR U3860 ( .A(n7951), .B(n7950), .Z(n7952) );
  XNOR U3861 ( .A(n7913), .B(n7912), .Z(n7915) );
  XOR U3862 ( .A(n7964), .B(n7890), .Z(n1498) );
  NANDN U3863 ( .A(n7891), .B(n1498), .Z(n1499) );
  NAND U3864 ( .A(n7964), .B(n7890), .Z(n1500) );
  AND U3865 ( .A(n1499), .B(n1500), .Z(n7943) );
  XNOR U3866 ( .A(n7976), .B(n7975), .Z(n7978) );
  XNOR U3867 ( .A(n8020), .B(n8019), .Z(n8021) );
  XNOR U3868 ( .A(n8026), .B(n8025), .Z(n8027) );
  XOR U3869 ( .A(n8195), .B(n8194), .Z(n8197) );
  NAND U3870 ( .A(n8067), .B(n8068), .Z(n1501) );
  NANDN U3871 ( .A(n8070), .B(n8069), .Z(n1502) );
  AND U3872 ( .A(n1501), .B(n1502), .Z(n8102) );
  XNOR U3873 ( .A(n8372), .B(n8371), .Z(n8373) );
  XOR U3874 ( .A(n8521), .B(n8520), .Z(n8549) );
  XOR U3875 ( .A(n8746), .B(n8745), .Z(n8661) );
  XNOR U3876 ( .A(n9144), .B(n9143), .Z(n9146) );
  XOR U3877 ( .A(n9370), .B(n9369), .Z(n9261) );
  XNOR U3878 ( .A(n9384), .B(n9383), .Z(n9385) );
  XNOR U3879 ( .A(n9663), .B(n9662), .Z(n9665) );
  XNOR U3880 ( .A(n9991), .B(n9990), .Z(n9969) );
  NAND U3881 ( .A(n10054), .B(n10053), .Z(n1503) );
  NANDN U3882 ( .A(n10052), .B(n10051), .Z(n1504) );
  AND U3883 ( .A(n1503), .B(n1504), .Z(n10253) );
  XNOR U3884 ( .A(n10408), .B(n10407), .Z(n10322) );
  XOR U3885 ( .A(n10487), .B(n10486), .Z(n10485) );
  XNOR U3886 ( .A(n10507), .B(n10506), .Z(n10504) );
  XNOR U3887 ( .A(n10689), .B(n10688), .Z(n10687) );
  XNOR U3888 ( .A(n10499), .B(n10498), .Z(n10496) );
  XNOR U3889 ( .A(n5035), .B(n5034), .Z(n5037) );
  XOR U3890 ( .A(n5023), .B(n4935), .Z(n1505) );
  NANDN U3891 ( .A(n4936), .B(n1505), .Z(n1506) );
  NAND U3892 ( .A(n5023), .B(n4935), .Z(n1507) );
  AND U3893 ( .A(n1506), .B(n1507), .Z(n4988) );
  XNOR U3894 ( .A(n5086), .B(n5085), .Z(n5088) );
  XOR U3895 ( .A(n5156), .B(n5155), .Z(n5148) );
  XOR U3896 ( .A(n5259), .B(n5258), .Z(n5241) );
  XNOR U3897 ( .A(n5606), .B(n5605), .Z(n5608) );
  XOR U3898 ( .A(n5781), .B(n5780), .Z(n5697) );
  XNOR U3899 ( .A(n5803), .B(n5802), .Z(n5909) );
  XNOR U3900 ( .A(n6033), .B(n6032), .Z(n5916) );
  XOR U3901 ( .A(n6173), .B(n6172), .Z(n6166) );
  XOR U3902 ( .A(n7326), .B(n7325), .Z(n7296) );
  NAND U3903 ( .A(n7089), .B(n7088), .Z(n1508) );
  NANDN U3904 ( .A(n7087), .B(n7086), .Z(n1509) );
  AND U3905 ( .A(n1508), .B(n1509), .Z(n7289) );
  XOR U3906 ( .A(n7205), .B(n7204), .Z(n7308) );
  XNOR U3907 ( .A(n7270), .B(n7269), .Z(n7318) );
  XNOR U3908 ( .A(n7466), .B(n7465), .Z(n7467) );
  XNOR U3909 ( .A(n7725), .B(n7724), .Z(n7722) );
  XOR U3910 ( .A(n7719), .B(n7718), .Z(n7717) );
  XOR U3911 ( .A(n7543), .B(n7542), .Z(n7541) );
  XNOR U3912 ( .A(n7472), .B(n7471), .Z(n7473) );
  XNOR U3913 ( .A(n7555), .B(n7554), .Z(n7552) );
  XNOR U3914 ( .A(n2134), .B(n2133), .Z(n2135) );
  XNOR U3915 ( .A(n2140), .B(n2139), .Z(n2141) );
  XOR U3916 ( .A(n2649), .B(n2648), .Z(n2651) );
  XNOR U3917 ( .A(n3191), .B(n3190), .Z(n3196) );
  NAND U3918 ( .A(n2996), .B(n2995), .Z(n1510) );
  NAND U3919 ( .A(n2994), .B(n2993), .Z(n1511) );
  AND U3920 ( .A(n1510), .B(n1511), .Z(n3203) );
  XNOR U3921 ( .A(n3456), .B(n3455), .Z(n3458) );
  XNOR U3922 ( .A(n3472), .B(n3471), .Z(n3473) );
  XNOR U3923 ( .A(n3754), .B(n3753), .Z(n3756) );
  XNOR U3924 ( .A(n4078), .B(n4077), .Z(n4080) );
  XNOR U3925 ( .A(n4072), .B(n4071), .Z(n4073) );
  XOR U3926 ( .A(n4445), .B(n4444), .Z(n4447) );
  XOR U3927 ( .A(n4526), .B(n4525), .Z(n4548) );
  XOR U3928 ( .A(n4394), .B(n4393), .Z(n4396) );
  XOR U3929 ( .A(n4603), .B(n4602), .Z(n4601) );
  XNOR U3930 ( .A(n4595), .B(n4594), .Z(n4592) );
  XNOR U3931 ( .A(n4239), .B(n4238), .Z(n4240) );
  XNOR U3932 ( .A(n46029), .B(n46028), .Z(n46031) );
  XNOR U3933 ( .A(n47359), .B(n47358), .Z(n47360) );
  XNOR U3934 ( .A(n47952), .B(n47951), .Z(n47869) );
  XNOR U3935 ( .A(n47845), .B(n47844), .Z(n47846) );
  NAND U3936 ( .A(n47853), .B(n47852), .Z(n1512) );
  NANDN U3937 ( .A(n47851), .B(n47850), .Z(n1513) );
  AND U3938 ( .A(n1512), .B(n1513), .Z(n48247) );
  NAND U3939 ( .A(n48210), .B(n48211), .Z(n48215) );
  NAND U3940 ( .A(n43306), .B(n43307), .Z(n1514) );
  NANDN U3941 ( .A(n43309), .B(n43308), .Z(n1515) );
  AND U3942 ( .A(n1514), .B(n1515), .Z(n43409) );
  XNOR U3943 ( .A(n43882), .B(n43881), .Z(n43884) );
  XNOR U3944 ( .A(n44025), .B(n44024), .Z(n44161) );
  XNOR U3945 ( .A(n45058), .B(n45057), .Z(n45059) );
  NAND U3946 ( .A(n45158), .B(n45157), .Z(n1516) );
  NAND U3947 ( .A(n45159), .B(n45160), .Z(n1517) );
  AND U3948 ( .A(n1516), .B(n1517), .Z(n1518) );
  XOR U3949 ( .A(n45226), .B(n45225), .Z(n1519) );
  XNOR U3950 ( .A(n45173), .B(n45172), .Z(n1520) );
  XNOR U3951 ( .A(n1519), .B(n1520), .Z(n1521) );
  XOR U3952 ( .A(n45276), .B(n45275), .Z(n1522) );
  XNOR U3953 ( .A(n45264), .B(n45263), .Z(n1523) );
  XNOR U3954 ( .A(n1522), .B(n1523), .Z(n1524) );
  XOR U3955 ( .A(n45304), .B(n45303), .Z(n1525) );
  XNOR U3956 ( .A(n45290), .B(n45289), .Z(n1526) );
  XNOR U3957 ( .A(n1525), .B(n1526), .Z(n1527) );
  XOR U3958 ( .A(n1524), .B(n1527), .Z(n1528) );
  XNOR U3959 ( .A(n1518), .B(n1521), .Z(n1529) );
  XNOR U3960 ( .A(n1528), .B(n1529), .Z(n1530) );
  NAND U3961 ( .A(n45153), .B(n45154), .Z(n1531) );
  NAND U3962 ( .A(n45155), .B(n45156), .Z(n1532) );
  NAND U3963 ( .A(n1531), .B(n1532), .Z(n1533) );
  XNOR U3964 ( .A(n1530), .B(n1533), .Z(n45305) );
  XOR U3965 ( .A(n45372), .B(n45371), .Z(n45370) );
  XOR U3966 ( .A(n39657), .B(n39658), .Z(n1534) );
  NANDN U3967 ( .A(n39659), .B(n1534), .Z(n1535) );
  NAND U3968 ( .A(n39657), .B(n39658), .Z(n1536) );
  AND U3969 ( .A(n1535), .B(n1536), .Z(n39706) );
  XNOR U3970 ( .A(n40233), .B(n40232), .Z(n40235) );
  XNOR U3971 ( .A(n40996), .B(n40995), .Z(n40998) );
  XNOR U3972 ( .A(n41003), .B(n41002), .Z(n41004) );
  XOR U3973 ( .A(n41273), .B(n41272), .Z(n41275) );
  XNOR U3974 ( .A(n42134), .B(n42133), .Z(n42055) );
  XOR U3975 ( .A(n42461), .B(n42460), .Z(n42459) );
  XNOR U3976 ( .A(n42455), .B(n42454), .Z(n42452) );
  XNOR U3977 ( .A(n42225), .B(n42224), .Z(n42449) );
  XNOR U3978 ( .A(n42090), .B(n42089), .Z(n42059) );
  XNOR U3979 ( .A(n42479), .B(n42478), .Z(n42476) );
  XNOR U3980 ( .A(n38711), .B(n38710), .Z(n38713) );
  NAND U3981 ( .A(n39221), .B(n39220), .Z(n1537) );
  NAND U3982 ( .A(n39219), .B(n39218), .Z(n1538) );
  AND U3983 ( .A(n1537), .B(n1538), .Z(n39310) );
  XOR U3984 ( .A(n39564), .B(n39563), .Z(n1539) );
  XNOR U3985 ( .A(n39565), .B(n1539), .Z(n39545) );
  NAND U3986 ( .A(n39276), .B(n39275), .Z(n1540) );
  NAND U3987 ( .A(n39274), .B(n39273), .Z(n1541) );
  AND U3988 ( .A(n1540), .B(n1541), .Z(n39526) );
  NAND U3989 ( .A(n39203), .B(n39202), .Z(n1542) );
  NAND U3990 ( .A(n39200), .B(n39201), .Z(n1543) );
  AND U3991 ( .A(n1542), .B(n1543), .Z(n39313) );
  OR U3992 ( .A(n36198), .B(n36199), .Z(n1544) );
  NAND U3993 ( .A(n36197), .B(n36196), .Z(n1545) );
  AND U3994 ( .A(n1544), .B(n1545), .Z(n36335) );
  NAND U3995 ( .A(n36442), .B(n36441), .Z(n1546) );
  NAND U3996 ( .A(n36440), .B(n36439), .Z(n1547) );
  AND U3997 ( .A(n1546), .B(n1547), .Z(n36716) );
  NAND U3998 ( .A(n36445), .B(n36446), .Z(n1548) );
  NAND U3999 ( .A(n36443), .B(n36444), .Z(n1549) );
  NAND U4000 ( .A(n1548), .B(n1549), .Z(n36709) );
  XOR U4001 ( .A(n36692), .B(n36691), .Z(n36690) );
  NAND U4002 ( .A(n36262), .B(n36261), .Z(n1550) );
  NAND U4003 ( .A(n36259), .B(n36260), .Z(n1551) );
  NAND U4004 ( .A(n1550), .B(n1551), .Z(n36387) );
  NAND U4005 ( .A(n31112), .B(n31111), .Z(n1552) );
  NAND U4006 ( .A(n31110), .B(n31109), .Z(n1553) );
  AND U4007 ( .A(n1552), .B(n1553), .Z(n31154) );
  XNOR U4008 ( .A(n31516), .B(n31515), .Z(n31518) );
  XNOR U4009 ( .A(n31592), .B(n31591), .Z(n31594) );
  XNOR U4010 ( .A(n32944), .B(n32943), .Z(n32946) );
  XNOR U4011 ( .A(n33273), .B(n33272), .Z(n33429) );
  XNOR U4012 ( .A(n33562), .B(n33561), .Z(n33476) );
  XNOR U4013 ( .A(n33628), .B(n33627), .Z(n33625) );
  XNOR U4014 ( .A(n33568), .B(n33567), .Z(n33463) );
  XOR U4015 ( .A(n33640), .B(n33639), .Z(n33638) );
  XOR U4016 ( .A(n28356), .B(n28355), .Z(n28358) );
  XNOR U4017 ( .A(n28668), .B(n28667), .Z(n28670) );
  XOR U4018 ( .A(n28876), .B(n28875), .Z(n28958) );
  XNOR U4019 ( .A(n30338), .B(n30337), .Z(n30494) );
  XNOR U4020 ( .A(n30634), .B(n30633), .Z(n30527) );
  XNOR U4021 ( .A(n30540), .B(n30539), .Z(n30541) );
  XNOR U4022 ( .A(n30625), .B(n30624), .Z(n30626) );
  XOR U4023 ( .A(n30949), .B(n30948), .Z(n30947) );
  XNOR U4024 ( .A(n30925), .B(n30924), .Z(n30922) );
  NAND U4025 ( .A(n25167), .B(n25250), .Z(n1554) );
  XOR U4026 ( .A(n25167), .B(n25250), .Z(n1555) );
  NANDN U4027 ( .A(n25166), .B(n1555), .Z(n1556) );
  NAND U4028 ( .A(n1554), .B(n1556), .Z(n25220) );
  XNOR U4029 ( .A(n27392), .B(n27391), .Z(n27548) );
  XNOR U4030 ( .A(n27688), .B(n27687), .Z(n27588) );
  XNOR U4031 ( .A(n27985), .B(n27984), .Z(n27983) );
  XNOR U4032 ( .A(n27749), .B(n27748), .Z(n27747) );
  XNOR U4033 ( .A(n27965), .B(n27964), .Z(n27743) );
  XOR U4034 ( .A(n22873), .B(n22872), .Z(n22902) );
  XNOR U4035 ( .A(n24771), .B(n24770), .Z(n24671) );
  NAND U4036 ( .A(n24609), .B(n24608), .Z(n1557) );
  NAND U4037 ( .A(n24607), .B(n24606), .Z(n1558) );
  AND U4038 ( .A(n1557), .B(n1558), .Z(n24665) );
  NAND U4039 ( .A(n24619), .B(n24618), .Z(n1559) );
  NAND U4040 ( .A(n24616), .B(n24617), .Z(n1560) );
  AND U4041 ( .A(n1559), .B(n1560), .Z(n24660) );
  XNOR U4042 ( .A(n24654), .B(n24653), .Z(n24655) );
  NAND U4043 ( .A(n24848), .B(n24847), .Z(n1561) );
  NAND U4044 ( .A(n24849), .B(n24850), .Z(n1562) );
  AND U4045 ( .A(n1561), .B(n1562), .Z(n1563) );
  NANDN U4046 ( .A(n24854), .B(n24853), .Z(n1564) );
  NANDN U4047 ( .A(n24852), .B(n24851), .Z(n1565) );
  NAND U4048 ( .A(n1564), .B(n1565), .Z(n1566) );
  XNOR U4049 ( .A(n1563), .B(n1566), .Z(n25012) );
  XNOR U4050 ( .A(n19785), .B(n19784), .Z(n19843) );
  XNOR U4051 ( .A(n20292), .B(n20291), .Z(n20280) );
  XNOR U4052 ( .A(n21161), .B(n21160), .Z(n21162) );
  XNOR U4053 ( .A(n21716), .B(n21715), .Z(n21718) );
  XNOR U4054 ( .A(n21831), .B(n21830), .Z(n21752) );
  NAND U4055 ( .A(n21605), .B(n21606), .Z(n1567) );
  NANDN U4056 ( .A(n21608), .B(n21607), .Z(n1568) );
  NAND U4057 ( .A(n1567), .B(n1568), .Z(n21734) );
  NAND U4058 ( .A(n21845), .B(n21844), .Z(n1569) );
  NAND U4059 ( .A(n21843), .B(n21842), .Z(n1570) );
  AND U4060 ( .A(n1569), .B(n1570), .Z(n22104) );
  NAND U4061 ( .A(n21669), .B(n21670), .Z(n1571) );
  NAND U4062 ( .A(n21667), .B(n21668), .Z(n1572) );
  NAND U4063 ( .A(n1571), .B(n1572), .Z(n21781) );
  NAND U4064 ( .A(n21749), .B(n21748), .Z(n1573) );
  NAND U4065 ( .A(n21747), .B(n21746), .Z(n1574) );
  AND U4066 ( .A(n1573), .B(n1574), .Z(n22147) );
  NAND U4067 ( .A(n21741), .B(n21740), .Z(n1575) );
  NAND U4068 ( .A(n21739), .B(n21738), .Z(n1576) );
  AND U4069 ( .A(n1575), .B(n1576), .Z(n22146) );
  NAND U4070 ( .A(n16542), .B(n16541), .Z(n1577) );
  NANDN U4071 ( .A(n16628), .B(n16619), .Z(n1578) );
  NAND U4072 ( .A(n1577), .B(n1578), .Z(n16555) );
  XNOR U4073 ( .A(n16699), .B(n16698), .Z(n16700) );
  XNOR U4074 ( .A(n17040), .B(n17039), .Z(n17042) );
  XNOR U4075 ( .A(n17129), .B(n17128), .Z(n17130) );
  OR U4076 ( .A(n17416), .B(n17417), .Z(n1579) );
  NAND U4077 ( .A(n17414), .B(n17415), .Z(n1580) );
  NAND U4078 ( .A(n1579), .B(n1580), .Z(n17528) );
  XOR U4079 ( .A(n17876), .B(n17875), .Z(n17987) );
  XOR U4080 ( .A(n18273), .B(n18272), .Z(n18416) );
  XNOR U4081 ( .A(n19036), .B(n19035), .Z(n18931) );
  XOR U4082 ( .A(n19359), .B(n19358), .Z(n1581) );
  XNOR U4083 ( .A(n19360), .B(n1581), .Z(n19345) );
  XNOR U4084 ( .A(n19335), .B(n19334), .Z(n19333) );
  XNOR U4085 ( .A(n19099), .B(n19098), .Z(n19097) );
  XNOR U4086 ( .A(n19315), .B(n19314), .Z(n19093) );
  NAND U4087 ( .A(n13677), .B(n13676), .Z(n1582) );
  NAND U4088 ( .A(n13675), .B(n13684), .Z(n1583) );
  AND U4089 ( .A(n1582), .B(n1583), .Z(n13690) );
  XNOR U4090 ( .A(n16029), .B(n16028), .Z(n16031) );
  NAND U4091 ( .A(n15997), .B(n15998), .Z(n1584) );
  NAND U4092 ( .A(n15995), .B(n15996), .Z(n1585) );
  NAND U4093 ( .A(n1584), .B(n1585), .Z(n16052) );
  NAND U4094 ( .A(n15967), .B(n15968), .Z(n1586) );
  NAND U4095 ( .A(n15965), .B(n15966), .Z(n1587) );
  NAND U4096 ( .A(n1586), .B(n1587), .Z(n16088) );
  NAND U4097 ( .A(n16011), .B(n16012), .Z(n1588) );
  NANDN U4098 ( .A(n16014), .B(n16013), .Z(n1589) );
  NAND U4099 ( .A(n1588), .B(n1589), .Z(n16048) );
  XOR U4100 ( .A(n16463), .B(n16462), .Z(n1590) );
  XNOR U4101 ( .A(n16464), .B(n1590), .Z(n16451) );
  NAND U4102 ( .A(n16107), .B(n16106), .Z(n1591) );
  NAND U4103 ( .A(n16104), .B(n16105), .Z(n1592) );
  NAND U4104 ( .A(n1591), .B(n1592), .Z(n16209) );
  NAND U4105 ( .A(n16111), .B(n16110), .Z(n1593) );
  NAND U4106 ( .A(n16108), .B(n16109), .Z(n1594) );
  AND U4107 ( .A(n1593), .B(n1594), .Z(n16199) );
  XOR U4108 ( .A(n10901), .B(n10818), .Z(n1595) );
  NANDN U4109 ( .A(n10819), .B(n1595), .Z(n1596) );
  NAND U4110 ( .A(n10901), .B(n10818), .Z(n1597) );
  AND U4111 ( .A(n1596), .B(n1597), .Z(n10872) );
  XNOR U4112 ( .A(n10964), .B(n10963), .Z(n10966) );
  XNOR U4113 ( .A(n11079), .B(n11078), .Z(n11081) );
  XNOR U4114 ( .A(n11158), .B(n11157), .Z(n11225) );
  XNOR U4115 ( .A(n12165), .B(n12164), .Z(n12167) );
  XNOR U4116 ( .A(n12172), .B(n12171), .Z(n12173) );
  XNOR U4117 ( .A(n13388), .B(n13387), .Z(n13385) );
  XNOR U4118 ( .A(n13325), .B(n13324), .Z(n13226) );
  XOR U4119 ( .A(n13648), .B(n13647), .Z(n13646) );
  XNOR U4120 ( .A(n13400), .B(n13399), .Z(n13397) );
  XNOR U4121 ( .A(n8365), .B(n8364), .Z(n8367) );
  XNOR U4122 ( .A(n8454), .B(n8453), .Z(n8456) );
  XNOR U4123 ( .A(n8649), .B(n8648), .Z(n8651) );
  XNOR U4124 ( .A(n10414), .B(n10413), .Z(n10308) );
  NAND U4125 ( .A(n10259), .B(n10258), .Z(n1598) );
  NAND U4126 ( .A(n10257), .B(n10256), .Z(n1599) );
  AND U4127 ( .A(n1598), .B(n1599), .Z(n10304) );
  NAND U4128 ( .A(n10268), .B(n10269), .Z(n1600) );
  NAND U4129 ( .A(n10266), .B(n10267), .Z(n1601) );
  NAND U4130 ( .A(n1600), .B(n1601), .Z(n10314) );
  XNOR U4131 ( .A(n10706), .B(n10705), .Z(n10703) );
  XNOR U4132 ( .A(n10477), .B(n10476), .Z(n10474) );
  XOR U4133 ( .A(n10730), .B(n10729), .Z(n10728) );
  NAND U4134 ( .A(n10290), .B(n10291), .Z(n1602) );
  XOR U4135 ( .A(n10290), .B(n10291), .Z(n1603) );
  NANDN U4136 ( .A(n10289), .B(n1603), .Z(n1604) );
  NAND U4137 ( .A(n1602), .B(n1604), .Z(n10724) );
  XNOR U4138 ( .A(n5275), .B(n5274), .Z(n5337) );
  XOR U4139 ( .A(n5568), .B(n5567), .Z(n5593) );
  XNOR U4140 ( .A(n6287), .B(n6286), .Z(n6289) );
  XNOR U4141 ( .A(n6294), .B(n6293), .Z(n6295) );
  XOR U4142 ( .A(n6712), .B(n6711), .Z(n6853) );
  XNOR U4143 ( .A(n7462), .B(n7461), .Z(n7369) );
  XOR U4144 ( .A(n7794), .B(n7793), .Z(n1605) );
  XNOR U4145 ( .A(n7795), .B(n1605), .Z(n7774) );
  XNOR U4146 ( .A(n7759), .B(n7758), .Z(n7756) );
  NAND U4147 ( .A(n1970), .B(n1971), .Z(n1606) );
  NAND U4148 ( .A(n2017), .B(n2595), .Z(n1607) );
  NAND U4149 ( .A(n1606), .B(n1607), .Z(n1978) );
  XOR U4150 ( .A(n1963), .B(n1962), .Z(n1608) );
  NANDN U4151 ( .A(n1964), .B(n1608), .Z(n1609) );
  NAND U4152 ( .A(n1963), .B(n1962), .Z(n1610) );
  AND U4153 ( .A(n1609), .B(n1610), .Z(n1982) );
  XNOR U4154 ( .A(n2269), .B(n2268), .Z(n2271) );
  XNOR U4155 ( .A(n2276), .B(n2275), .Z(n2277) );
  XNOR U4156 ( .A(n2413), .B(n2412), .Z(n2415) );
  XNOR U4157 ( .A(n2869), .B(n2868), .Z(n2871) );
  XNOR U4158 ( .A(n3229), .B(n3228), .Z(n3221) );
  XNOR U4159 ( .A(n4530), .B(n4529), .Z(n4531) );
  XNOR U4160 ( .A(n4833), .B(n4832), .Z(n4830) );
  XNOR U4161 ( .A(n4787), .B(n4786), .Z(n4821) );
  XNOR U4162 ( .A(n4795), .B(n4794), .Z(n4793) );
  XOR U4163 ( .A(n45488), .B(n45489), .Z(n1611) );
  NANDN U4164 ( .A(n45490), .B(n1611), .Z(n1612) );
  NAND U4165 ( .A(n45488), .B(n45489), .Z(n1613) );
  AND U4166 ( .A(n1612), .B(n1613), .Z(n45549) );
  XOR U4167 ( .A(n45713), .B(n45714), .Z(n1614) );
  NANDN U4168 ( .A(n45715), .B(n1614), .Z(n1615) );
  NAND U4169 ( .A(n45713), .B(n45714), .Z(n1616) );
  AND U4170 ( .A(n1615), .B(n1616), .Z(n45780) );
  XOR U4171 ( .A(n45936), .B(n45937), .Z(n1617) );
  NANDN U4172 ( .A(n45938), .B(n1617), .Z(n1618) );
  NAND U4173 ( .A(n45936), .B(n45937), .Z(n1619) );
  AND U4174 ( .A(n1618), .B(n1619), .Z(n46023) );
  XOR U4175 ( .A(n46456), .B(n46457), .Z(n1620) );
  NANDN U4176 ( .A(n46458), .B(n1620), .Z(n1621) );
  NAND U4177 ( .A(n46456), .B(n46457), .Z(n1622) );
  AND U4178 ( .A(n1621), .B(n1622), .Z(n46682) );
  XOR U4179 ( .A(n47217), .B(n47218), .Z(n1623) );
  NANDN U4180 ( .A(n47219), .B(n1623), .Z(n1624) );
  NAND U4181 ( .A(n47217), .B(n47218), .Z(n1625) );
  AND U4182 ( .A(n1624), .B(n1625), .Z(n47365) );
  NAND U4183 ( .A(n47681), .B(n47682), .Z(n1626) );
  XOR U4184 ( .A(n47681), .B(n47682), .Z(n1627) );
  NANDN U4185 ( .A(n47680), .B(n1627), .Z(n1628) );
  NAND U4186 ( .A(n1626), .B(n1628), .Z(n47835) );
  XNOR U4187 ( .A(n48011), .B(n48010), .Z(n48009) );
  NANDN U4188 ( .A(n42558), .B(n42560), .Z(n1629) );
  OR U4189 ( .A(n42560), .B(n42561), .Z(n1630) );
  NAND U4190 ( .A(n42559), .B(n1630), .Z(n1631) );
  NAND U4191 ( .A(n1629), .B(n1631), .Z(n42579) );
  XOR U4192 ( .A(n42657), .B(n42658), .Z(n1632) );
  NANDN U4193 ( .A(n42659), .B(n1632), .Z(n1633) );
  NAND U4194 ( .A(n42657), .B(n42658), .Z(n1634) );
  AND U4195 ( .A(n1633), .B(n1634), .Z(n42710) );
  XOR U4196 ( .A(n42819), .B(n42820), .Z(n1635) );
  NANDN U4197 ( .A(n42821), .B(n1635), .Z(n1636) );
  NAND U4198 ( .A(n42819), .B(n42820), .Z(n1637) );
  AND U4199 ( .A(n1636), .B(n1637), .Z(n42837) );
  XOR U4200 ( .A(n43116), .B(n43117), .Z(n1638) );
  NANDN U4201 ( .A(n43118), .B(n1638), .Z(n1639) );
  NAND U4202 ( .A(n43116), .B(n43117), .Z(n1640) );
  AND U4203 ( .A(n1639), .B(n1640), .Z(n43208) );
  XOR U4204 ( .A(n43396), .B(n43397), .Z(n1641) );
  NANDN U4205 ( .A(n43398), .B(n1641), .Z(n1642) );
  NAND U4206 ( .A(n43396), .B(n43397), .Z(n1643) );
  AND U4207 ( .A(n1642), .B(n1643), .Z(n43412) );
  XOR U4208 ( .A(n43749), .B(n43750), .Z(n1644) );
  NANDN U4209 ( .A(n43751), .B(n1644), .Z(n1645) );
  NAND U4210 ( .A(n43749), .B(n43750), .Z(n1646) );
  AND U4211 ( .A(n1645), .B(n1646), .Z(n43876) );
  NAND U4212 ( .A(n44448), .B(n44449), .Z(n1647) );
  XOR U4213 ( .A(n44448), .B(n44449), .Z(n1648) );
  NANDN U4214 ( .A(n44447), .B(n1648), .Z(n1649) );
  NAND U4215 ( .A(n1647), .B(n1649), .Z(n44604) );
  NAND U4216 ( .A(n44931), .B(n44932), .Z(n1650) );
  XOR U4217 ( .A(n44931), .B(n44932), .Z(n1651) );
  NANDN U4218 ( .A(n44930), .B(n1651), .Z(n1652) );
  NAND U4219 ( .A(n1650), .B(n1652), .Z(n44934) );
  XNOR U4220 ( .A(n45118), .B(n45117), .Z(n45115) );
  NAND U4221 ( .A(n39611), .B(n39612), .Z(n1653) );
  XOR U4222 ( .A(n39611), .B(n39612), .Z(n1654) );
  NANDN U4223 ( .A(n39610), .B(n1654), .Z(n1655) );
  NAND U4224 ( .A(n1653), .B(n1655), .Z(n39622) );
  XOR U4225 ( .A(n39796), .B(n39797), .Z(n1656) );
  NANDN U4226 ( .A(n39798), .B(n1656), .Z(n1657) );
  NAND U4227 ( .A(n39796), .B(n39797), .Z(n1658) );
  AND U4228 ( .A(n1657), .B(n1658), .Z(n39848) );
  XOR U4229 ( .A(n40072), .B(n40073), .Z(n1659) );
  NANDN U4230 ( .A(n40074), .B(n1659), .Z(n1660) );
  NAND U4231 ( .A(n40072), .B(n40073), .Z(n1661) );
  AND U4232 ( .A(n1660), .B(n1661), .Z(n40150) );
  XOR U4233 ( .A(n40506), .B(n40507), .Z(n1662) );
  NANDN U4234 ( .A(n40508), .B(n1662), .Z(n1663) );
  NAND U4235 ( .A(n40506), .B(n40507), .Z(n1664) );
  AND U4236 ( .A(n1663), .B(n1664), .Z(n40625) );
  NAND U4237 ( .A(n40864), .B(n40865), .Z(n1665) );
  XOR U4238 ( .A(n40864), .B(n40865), .Z(n1666) );
  NAND U4239 ( .A(n1666), .B(n40863), .Z(n1667) );
  NAND U4240 ( .A(n1665), .B(n1667), .Z(n40990) );
  NAND U4241 ( .A(n41573), .B(n41574), .Z(n1668) );
  XOR U4242 ( .A(n41573), .B(n41574), .Z(n1669) );
  NANDN U4243 ( .A(n41572), .B(n1669), .Z(n1670) );
  NAND U4244 ( .A(n1668), .B(n1670), .Z(n41863) );
  XOR U4245 ( .A(n42038), .B(n42037), .Z(n1671) );
  NANDN U4246 ( .A(n42039), .B(n1671), .Z(n1672) );
  NAND U4247 ( .A(n42038), .B(n42037), .Z(n1673) );
  AND U4248 ( .A(n1672), .B(n1673), .Z(n42488) );
  XOR U4249 ( .A(n36811), .B(n36812), .Z(n1674) );
  NANDN U4250 ( .A(n36813), .B(n1674), .Z(n1675) );
  NAND U4251 ( .A(n36811), .B(n36812), .Z(n1676) );
  AND U4252 ( .A(n1675), .B(n1676), .Z(n36831) );
  XOR U4253 ( .A(n36906), .B(n36907), .Z(n1677) );
  NANDN U4254 ( .A(n36908), .B(n1677), .Z(n1678) );
  NAND U4255 ( .A(n36906), .B(n36907), .Z(n1679) );
  AND U4256 ( .A(n1678), .B(n1679), .Z(n36924) );
  XOR U4257 ( .A(n37074), .B(n37075), .Z(n1680) );
  NANDN U4258 ( .A(n37076), .B(n1680), .Z(n1681) );
  NAND U4259 ( .A(n37074), .B(n37075), .Z(n1682) );
  AND U4260 ( .A(n1681), .B(n1682), .Z(n37141) );
  XOR U4261 ( .A(n37476), .B(n37475), .Z(n1683) );
  NANDN U4262 ( .A(n37477), .B(n1683), .Z(n1684) );
  NAND U4263 ( .A(n37476), .B(n37475), .Z(n1685) );
  AND U4264 ( .A(n1684), .B(n1685), .Z(n37572) );
  XOR U4265 ( .A(n37767), .B(n37768), .Z(n1686) );
  NANDN U4266 ( .A(n37769), .B(n1686), .Z(n1687) );
  NAND U4267 ( .A(n37767), .B(n37768), .Z(n1688) );
  AND U4268 ( .A(n1687), .B(n1688), .Z(n37888) );
  XOR U4269 ( .A(n38131), .B(n38130), .Z(n1689) );
  NANDN U4270 ( .A(n38132), .B(n1689), .Z(n1690) );
  NAND U4271 ( .A(n38131), .B(n38130), .Z(n1691) );
  AND U4272 ( .A(n1690), .B(n1691), .Z(n38262) );
  XOR U4273 ( .A(n38700), .B(n38701), .Z(n1692) );
  NANDN U4274 ( .A(n38702), .B(n1692), .Z(n1693) );
  NAND U4275 ( .A(n38700), .B(n38701), .Z(n1694) );
  AND U4276 ( .A(n1693), .B(n1694), .Z(n38718) );
  XNOR U4277 ( .A(n39574), .B(n39573), .Z(n39572) );
  NAND U4278 ( .A(n33978), .B(n33977), .Z(n1695) );
  XOR U4279 ( .A(n33978), .B(n33977), .Z(n1696) );
  NANDN U4280 ( .A(n33979), .B(n1696), .Z(n1697) );
  NAND U4281 ( .A(n1695), .B(n1697), .Z(n33998) );
  XOR U4282 ( .A(n34076), .B(n34077), .Z(n1698) );
  NANDN U4283 ( .A(n34078), .B(n1698), .Z(n1699) );
  NAND U4284 ( .A(n34076), .B(n34077), .Z(n1700) );
  AND U4285 ( .A(n1699), .B(n1700), .Z(n34129) );
  XOR U4286 ( .A(n34240), .B(n34241), .Z(n1701) );
  NANDN U4287 ( .A(n34242), .B(n1701), .Z(n1702) );
  NAND U4288 ( .A(n34240), .B(n34241), .Z(n1703) );
  AND U4289 ( .A(n1702), .B(n1703), .Z(n34307) );
  XOR U4290 ( .A(n34461), .B(n34462), .Z(n1704) );
  NANDN U4291 ( .A(n34463), .B(n1704), .Z(n1705) );
  NAND U4292 ( .A(n34461), .B(n34462), .Z(n1706) );
  AND U4293 ( .A(n1705), .B(n1706), .Z(n34544) );
  NAND U4294 ( .A(n34958), .B(n34957), .Z(n1707) );
  XOR U4295 ( .A(n34958), .B(n34957), .Z(n1708) );
  NANDN U4296 ( .A(n34959), .B(n1708), .Z(n1709) );
  NAND U4297 ( .A(n1707), .B(n1709), .Z(n35069) );
  XOR U4298 ( .A(n35320), .B(n35321), .Z(n1710) );
  NANDN U4299 ( .A(n35322), .B(n1710), .Z(n1711) );
  NAND U4300 ( .A(n35320), .B(n35321), .Z(n1712) );
  AND U4301 ( .A(n1711), .B(n1712), .Z(n35451) );
  XOR U4302 ( .A(n35611), .B(n35612), .Z(n1713) );
  NANDN U4303 ( .A(n35613), .B(n1713), .Z(n1714) );
  NAND U4304 ( .A(n35611), .B(n35612), .Z(n1715) );
  AND U4305 ( .A(n1714), .B(n1715), .Z(n35754) );
  XOR U4306 ( .A(n36174), .B(n36175), .Z(n1716) );
  NANDN U4307 ( .A(n36176), .B(n1716), .Z(n1717) );
  NAND U4308 ( .A(n36174), .B(n36175), .Z(n1718) );
  AND U4309 ( .A(n1717), .B(n1718), .Z(n36318) );
  XNOR U4310 ( .A(n36746), .B(n36745), .Z(n36744) );
  XOR U4311 ( .A(n31014), .B(n31013), .Z(n1719) );
  NANDN U4312 ( .A(n31015), .B(n1719), .Z(n1720) );
  NAND U4313 ( .A(n31014), .B(n31013), .Z(n1721) );
  AND U4314 ( .A(n1720), .B(n1721), .Z(n31037) );
  XNOR U4315 ( .A(n31059), .B(n31058), .Z(n31052) );
  NAND U4316 ( .A(n31250), .B(n31249), .Z(n1722) );
  XOR U4317 ( .A(n31250), .B(n31249), .Z(n1723) );
  NANDN U4318 ( .A(n31251), .B(n1723), .Z(n1724) );
  NAND U4319 ( .A(n1722), .B(n1724), .Z(n31260) );
  XOR U4320 ( .A(n31443), .B(n31444), .Z(n1725) );
  NANDN U4321 ( .A(n31445), .B(n1725), .Z(n1726) );
  NAND U4322 ( .A(n31443), .B(n31444), .Z(n1727) );
  AND U4323 ( .A(n1726), .B(n1727), .Z(n31510) );
  XOR U4324 ( .A(n31793), .B(n31792), .Z(n1728) );
  NANDN U4325 ( .A(n31794), .B(n1728), .Z(n1729) );
  NAND U4326 ( .A(n31793), .B(n31792), .Z(n1730) );
  AND U4327 ( .A(n1729), .B(n1730), .Z(n31897) );
  XOR U4328 ( .A(n32233), .B(n32234), .Z(n1731) );
  NANDN U4329 ( .A(n32235), .B(n1731), .Z(n1732) );
  NAND U4330 ( .A(n32233), .B(n32234), .Z(n1733) );
  AND U4331 ( .A(n1732), .B(n1733), .Z(n32360) );
  XNOR U4332 ( .A(n32502), .B(n32501), .Z(n32495) );
  XOR U4333 ( .A(n32653), .B(n32654), .Z(n1734) );
  NANDN U4334 ( .A(n32655), .B(n1734), .Z(n1735) );
  NAND U4335 ( .A(n32653), .B(n32654), .Z(n1736) );
  AND U4336 ( .A(n1735), .B(n1736), .Z(n32931) );
  XNOR U4337 ( .A(n33616), .B(n33615), .Z(n33614) );
  NAND U4338 ( .A(n28068), .B(n28069), .Z(n1737) );
  NAND U4339 ( .A(n28067), .B(n28161), .Z(n1738) );
  NAND U4340 ( .A(n1737), .B(n1738), .Z(n28087) );
  XOR U4341 ( .A(n28152), .B(n28151), .Z(n1739) );
  NANDN U4342 ( .A(n28153), .B(n1739), .Z(n1740) );
  NAND U4343 ( .A(n28152), .B(n28151), .Z(n1741) );
  AND U4344 ( .A(n1740), .B(n1741), .Z(n28186) );
  XOR U4345 ( .A(n28252), .B(n28253), .Z(n1742) );
  NANDN U4346 ( .A(n28254), .B(n1742), .Z(n1743) );
  NAND U4347 ( .A(n28252), .B(n28253), .Z(n1744) );
  AND U4348 ( .A(n1743), .B(n1744), .Z(n28350) );
  XOR U4349 ( .A(n28575), .B(n28576), .Z(n1745) );
  NANDN U4350 ( .A(n28577), .B(n1745), .Z(n1746) );
  NAND U4351 ( .A(n28575), .B(n28576), .Z(n1747) );
  AND U4352 ( .A(n1746), .B(n1747), .Z(n28662) );
  XOR U4353 ( .A(n29311), .B(n29312), .Z(n1748) );
  NANDN U4354 ( .A(n29313), .B(n1748), .Z(n1749) );
  NAND U4355 ( .A(n29311), .B(n29312), .Z(n1750) );
  AND U4356 ( .A(n1749), .B(n1750), .Z(n29438) );
  NAND U4357 ( .A(n29863), .B(n29864), .Z(n1751) );
  XOR U4358 ( .A(n29863), .B(n29864), .Z(n1752) );
  NANDN U4359 ( .A(n29862), .B(n1752), .Z(n1753) );
  NAND U4360 ( .A(n1751), .B(n1753), .Z(n29872) );
  XOR U4361 ( .A(n30184), .B(n30185), .Z(n1754) );
  NANDN U4362 ( .A(n30186), .B(n1754), .Z(n1755) );
  NAND U4363 ( .A(n30184), .B(n30185), .Z(n1756) );
  AND U4364 ( .A(n1755), .B(n1756), .Z(n30499) );
  XNOR U4365 ( .A(n30969), .B(n30968), .Z(n30967) );
  XOR U4366 ( .A(n25178), .B(n25179), .Z(n1757) );
  NANDN U4367 ( .A(n25180), .B(n1757), .Z(n1758) );
  NAND U4368 ( .A(n25178), .B(n25179), .Z(n1759) );
  AND U4369 ( .A(n1758), .B(n1759), .Z(n25213) );
  XOR U4370 ( .A(n25274), .B(n25275), .Z(n1760) );
  NANDN U4371 ( .A(n25276), .B(n1760), .Z(n1761) );
  NAND U4372 ( .A(n25274), .B(n25275), .Z(n1762) );
  AND U4373 ( .A(n1761), .B(n1762), .Z(n25363) );
  NAND U4374 ( .A(n25508), .B(n25509), .Z(n1763) );
  XOR U4375 ( .A(n25508), .B(n25509), .Z(n1764) );
  NANDN U4376 ( .A(n25507), .B(n1764), .Z(n1765) );
  NAND U4377 ( .A(n1763), .B(n1765), .Z(n25647) );
  XOR U4378 ( .A(n25819), .B(n25818), .Z(n1766) );
  NANDN U4379 ( .A(n25820), .B(n1766), .Z(n1767) );
  NAND U4380 ( .A(n25819), .B(n25818), .Z(n1768) );
  AND U4381 ( .A(n1767), .B(n1768), .Z(n25915) );
  NAND U4382 ( .A(n26127), .B(n26126), .Z(n1769) );
  XOR U4383 ( .A(n26127), .B(n26126), .Z(n1770) );
  NANDN U4384 ( .A(n26128), .B(n1770), .Z(n1771) );
  NAND U4385 ( .A(n1769), .B(n1771), .Z(n26233) );
  NAND U4386 ( .A(n26489), .B(n26490), .Z(n1772) );
  XOR U4387 ( .A(n26489), .B(n26490), .Z(n1773) );
  NANDN U4388 ( .A(n26488), .B(n1773), .Z(n1774) );
  NAND U4389 ( .A(n1772), .B(n1774), .Z(n26616) );
  XOR U4390 ( .A(n27072), .B(n27073), .Z(n1775) );
  NANDN U4391 ( .A(n27074), .B(n1775), .Z(n1776) );
  NAND U4392 ( .A(n27072), .B(n27073), .Z(n1777) );
  AND U4393 ( .A(n1776), .B(n1777), .Z(n27232) );
  XNOR U4394 ( .A(n27737), .B(n27736), .Z(n27735) );
  XOR U4395 ( .A(n22248), .B(n22249), .Z(n1778) );
  NANDN U4396 ( .A(n22250), .B(n1778), .Z(n1779) );
  NAND U4397 ( .A(n22248), .B(n22249), .Z(n1780) );
  AND U4398 ( .A(n1779), .B(n1780), .Z(n22284) );
  XOR U4399 ( .A(n22448), .B(n22449), .Z(n1781) );
  NANDN U4400 ( .A(n22450), .B(n1781), .Z(n1782) );
  NAND U4401 ( .A(n22448), .B(n22449), .Z(n1783) );
  AND U4402 ( .A(n1782), .B(n1783), .Z(n22566) );
  XOR U4403 ( .A(n22802), .B(n22803), .Z(n1784) );
  NANDN U4404 ( .A(n22804), .B(n1784), .Z(n1785) );
  NAND U4405 ( .A(n22802), .B(n22803), .Z(n1786) );
  AND U4406 ( .A(n1785), .B(n1786), .Z(n22896) );
  XOR U4407 ( .A(n23099), .B(n23098), .Z(n1787) );
  NANDN U4408 ( .A(n23100), .B(n1787), .Z(n1788) );
  NAND U4409 ( .A(n23099), .B(n23098), .Z(n1789) );
  AND U4410 ( .A(n1788), .B(n1789), .Z(n23212) );
  XOR U4411 ( .A(n23882), .B(n23883), .Z(n1790) );
  NANDN U4412 ( .A(n23884), .B(n1790), .Z(n1791) );
  NAND U4413 ( .A(n23882), .B(n23883), .Z(n1792) );
  AND U4414 ( .A(n1791), .B(n1792), .Z(n24026) );
  NAND U4415 ( .A(n24635), .B(n24636), .Z(n1793) );
  XOR U4416 ( .A(n24635), .B(n24636), .Z(n1794) );
  NANDN U4417 ( .A(n24634), .B(n1794), .Z(n1795) );
  NAND U4418 ( .A(n1793), .B(n1795), .Z(n24645) );
  XNOR U4419 ( .A(n24826), .B(n24825), .Z(n24823) );
  NANDN U4420 ( .A(n19434), .B(n19436), .Z(n1796) );
  OR U4421 ( .A(n19436), .B(n19437), .Z(n1797) );
  NAND U4422 ( .A(n19435), .B(n1797), .Z(n1798) );
  NAND U4423 ( .A(n1796), .B(n1798), .Z(n19460) );
  NAND U4424 ( .A(n19552), .B(n19553), .Z(n1799) );
  XOR U4425 ( .A(n19552), .B(n19553), .Z(n1800) );
  NANDN U4426 ( .A(n19551), .B(n1800), .Z(n1801) );
  NAND U4427 ( .A(n1799), .B(n1801), .Z(n19596) );
  XOR U4428 ( .A(n19657), .B(n19658), .Z(n1802) );
  NANDN U4429 ( .A(n19659), .B(n1802), .Z(n1803) );
  NAND U4430 ( .A(n19657), .B(n19658), .Z(n1804) );
  AND U4431 ( .A(n1803), .B(n1804), .Z(n19769) );
  NAND U4432 ( .A(n19989), .B(n19990), .Z(n1805) );
  XOR U4433 ( .A(n19989), .B(n19990), .Z(n1806) );
  NANDN U4434 ( .A(n19988), .B(n1806), .Z(n1807) );
  NAND U4435 ( .A(n1805), .B(n1807), .Z(n20070) );
  XOR U4436 ( .A(n20183), .B(n20182), .Z(n1808) );
  NANDN U4437 ( .A(n20184), .B(n1808), .Z(n1809) );
  NAND U4438 ( .A(n20183), .B(n20182), .Z(n1810) );
  AND U4439 ( .A(n1809), .B(n1810), .Z(n20287) );
  NAND U4440 ( .A(n20631), .B(n20632), .Z(n1811) );
  XOR U4441 ( .A(n20631), .B(n20632), .Z(n1812) );
  NANDN U4442 ( .A(n20630), .B(n1812), .Z(n1813) );
  NAND U4443 ( .A(n1811), .B(n1813), .Z(n20750) );
  XOR U4444 ( .A(n21021), .B(n21020), .Z(n1814) );
  NANDN U4445 ( .A(n21022), .B(n1814), .Z(n1815) );
  NAND U4446 ( .A(n21021), .B(n21020), .Z(n1816) );
  AND U4447 ( .A(n1815), .B(n1816), .Z(n21168) );
  XOR U4448 ( .A(n21589), .B(n21590), .Z(n1817) );
  NANDN U4449 ( .A(n21591), .B(n1817), .Z(n1818) );
  NAND U4450 ( .A(n21589), .B(n21590), .Z(n1819) );
  AND U4451 ( .A(n1818), .B(n1819), .Z(n21722) );
  XNOR U4452 ( .A(n22160), .B(n22159), .Z(n22158) );
  XOR U4453 ( .A(n16545), .B(n16546), .Z(n1820) );
  NANDN U4454 ( .A(n16547), .B(n1820), .Z(n1821) );
  NAND U4455 ( .A(n16545), .B(n16546), .Z(n1822) );
  AND U4456 ( .A(n1821), .B(n1822), .Z(n16560) );
  XOR U4457 ( .A(n16645), .B(n16646), .Z(n1823) );
  NANDN U4458 ( .A(n16647), .B(n1823), .Z(n1824) );
  NAND U4459 ( .A(n16645), .B(n16646), .Z(n1825) );
  AND U4460 ( .A(n1824), .B(n1825), .Z(n16693) );
  XOR U4461 ( .A(n16955), .B(n16956), .Z(n1826) );
  NANDN U4462 ( .A(n16957), .B(n1826), .Z(n1827) );
  NAND U4463 ( .A(n16955), .B(n16956), .Z(n1828) );
  AND U4464 ( .A(n1827), .B(n1828), .Z(n17034) );
  XOR U4465 ( .A(n17404), .B(n17405), .Z(n1829) );
  NANDN U4466 ( .A(n17406), .B(n1829), .Z(n1830) );
  NAND U4467 ( .A(n17404), .B(n17405), .Z(n1831) );
  AND U4468 ( .A(n1830), .B(n1831), .Z(n17514) );
  NAND U4469 ( .A(n17765), .B(n17766), .Z(n1832) );
  XOR U4470 ( .A(n17765), .B(n17766), .Z(n1833) );
  NANDN U4471 ( .A(n17764), .B(n1833), .Z(n1834) );
  NAND U4472 ( .A(n1832), .B(n1834), .Z(n17982) );
  XOR U4473 ( .A(n18261), .B(n18260), .Z(n1835) );
  NANDN U4474 ( .A(n18262), .B(n1835), .Z(n1836) );
  NAND U4475 ( .A(n18261), .B(n18260), .Z(n1837) );
  AND U4476 ( .A(n1836), .B(n1837), .Z(n18412) );
  NAND U4477 ( .A(n18738), .B(n18739), .Z(n1838) );
  XOR U4478 ( .A(n18738), .B(n18739), .Z(n1839) );
  NANDN U4479 ( .A(n18737), .B(n1839), .Z(n1840) );
  NAND U4480 ( .A(n1838), .B(n1840), .Z(n18906) );
  XNOR U4481 ( .A(n19087), .B(n19086), .Z(n19085) );
  XOR U4482 ( .A(n13727), .B(n13728), .Z(n1841) );
  NANDN U4483 ( .A(n13729), .B(n1841), .Z(n1842) );
  NAND U4484 ( .A(n13727), .B(n13728), .Z(n1843) );
  AND U4485 ( .A(n1842), .B(n1843), .Z(n13744) );
  XOR U4486 ( .A(n13828), .B(n13829), .Z(n1844) );
  NANDN U4487 ( .A(n13830), .B(n1844), .Z(n1845) );
  NAND U4488 ( .A(n13828), .B(n13829), .Z(n1846) );
  AND U4489 ( .A(n1845), .B(n1846), .Z(n13846) );
  XOR U4490 ( .A(n14062), .B(n14061), .Z(n1847) );
  NANDN U4491 ( .A(n14063), .B(n1847), .Z(n1848) );
  NAND U4492 ( .A(n14062), .B(n14061), .Z(n1849) );
  AND U4493 ( .A(n1848), .B(n1849), .Z(n14078) );
  NAND U4494 ( .A(n14313), .B(n14314), .Z(n1850) );
  XOR U4495 ( .A(n14313), .B(n14314), .Z(n1851) );
  NANDN U4496 ( .A(n14312), .B(n1851), .Z(n1852) );
  NAND U4497 ( .A(n1850), .B(n1852), .Z(n14483) );
  NAND U4498 ( .A(n14698), .B(n14699), .Z(n1853) );
  XOR U4499 ( .A(n14698), .B(n14699), .Z(n1854) );
  NANDN U4500 ( .A(n14700), .B(n1854), .Z(n1855) );
  NAND U4501 ( .A(n1853), .B(n1855), .Z(n14809) );
  XOR U4502 ( .A(n15056), .B(n15057), .Z(n1856) );
  NANDN U4503 ( .A(n15058), .B(n1856), .Z(n1857) );
  NAND U4504 ( .A(n15056), .B(n15057), .Z(n1858) );
  AND U4505 ( .A(n1857), .B(n1858), .Z(n15066) );
  NAND U4506 ( .A(n15460), .B(n15461), .Z(n1859) );
  XOR U4507 ( .A(n15460), .B(n15461), .Z(n1860) );
  NANDN U4508 ( .A(n15459), .B(n1860), .Z(n1861) );
  NAND U4509 ( .A(n1859), .B(n1861), .Z(n15605) );
  XOR U4510 ( .A(n15891), .B(n15892), .Z(n1862) );
  NANDN U4511 ( .A(n15893), .B(n1862), .Z(n1863) );
  NAND U4512 ( .A(n15891), .B(n15892), .Z(n1864) );
  AND U4513 ( .A(n1863), .B(n1864), .Z(n16023) );
  XNOR U4514 ( .A(n16487), .B(n16486), .Z(n16485) );
  XOR U4515 ( .A(n10830), .B(n10831), .Z(n1865) );
  NANDN U4516 ( .A(n10832), .B(n1865), .Z(n1866) );
  NAND U4517 ( .A(n10830), .B(n10831), .Z(n1867) );
  AND U4518 ( .A(n1866), .B(n1867), .Z(n10865) );
  XOR U4519 ( .A(n10953), .B(n10954), .Z(n1868) );
  NANDN U4520 ( .A(n10955), .B(n1868), .Z(n1869) );
  NAND U4521 ( .A(n10953), .B(n10954), .Z(n1870) );
  AND U4522 ( .A(n1869), .B(n1870), .Z(n10971) );
  XOR U4523 ( .A(n11384), .B(n11383), .Z(n1871) );
  NANDN U4524 ( .A(n11385), .B(n1871), .Z(n1872) );
  NAND U4525 ( .A(n11384), .B(n11383), .Z(n1873) );
  AND U4526 ( .A(n1872), .B(n1873), .Z(n11466) );
  NAND U4527 ( .A(n11670), .B(n11668), .Z(n1874) );
  XOR U4528 ( .A(n11670), .B(n11668), .Z(n1875) );
  NAND U4529 ( .A(n1875), .B(n11669), .Z(n1876) );
  NAND U4530 ( .A(n1874), .B(n1876), .Z(n11782) );
  XNOR U4531 ( .A(n12038), .B(n12037), .Z(n12031) );
  XOR U4532 ( .A(n12725), .B(n12726), .Z(n1877) );
  NANDN U4533 ( .A(n12727), .B(n1877), .Z(n1878) );
  NAND U4534 ( .A(n12725), .B(n12726), .Z(n1879) );
  AND U4535 ( .A(n1878), .B(n1879), .Z(n13027) );
  XOR U4536 ( .A(n13199), .B(n13198), .Z(n1880) );
  NANDN U4537 ( .A(n13200), .B(n1880), .Z(n1881) );
  NAND U4538 ( .A(n13199), .B(n13198), .Z(n1882) );
  AND U4539 ( .A(n1881), .B(n1882), .Z(n13376) );
  XOR U4540 ( .A(n7902), .B(n7903), .Z(n1883) );
  NANDN U4541 ( .A(n7904), .B(n1883), .Z(n1884) );
  NAND U4542 ( .A(n7902), .B(n7903), .Z(n1885) );
  AND U4543 ( .A(n1884), .B(n1885), .Z(n7938) );
  NAND U4544 ( .A(n8088), .B(n8087), .Z(n1886) );
  XOR U4545 ( .A(n8088), .B(n8087), .Z(n1887) );
  NANDN U4546 ( .A(n8089), .B(n1887), .Z(n1888) );
  NAND U4547 ( .A(n1886), .B(n1888), .Z(n8098) );
  XOR U4548 ( .A(n8280), .B(n8281), .Z(n1889) );
  NANDN U4549 ( .A(n8282), .B(n1889), .Z(n1890) );
  NAND U4550 ( .A(n8280), .B(n8281), .Z(n1891) );
  AND U4551 ( .A(n1890), .B(n1891), .Z(n8359) );
  XOR U4552 ( .A(n8885), .B(n8886), .Z(n1892) );
  NANDN U4553 ( .A(n8887), .B(n1892), .Z(n1893) );
  NAND U4554 ( .A(n8885), .B(n8886), .Z(n1894) );
  AND U4555 ( .A(n1893), .B(n1894), .Z(n9005) );
  XNOR U4556 ( .A(n9127), .B(n9126), .Z(n9133) );
  NAND U4557 ( .A(n9521), .B(n9522), .Z(n1895) );
  XOR U4558 ( .A(n9521), .B(n9522), .Z(n1896) );
  NANDN U4559 ( .A(n9520), .B(n1896), .Z(n1897) );
  NAND U4560 ( .A(n1895), .B(n1897), .Z(n9531) );
  XOR U4561 ( .A(n9818), .B(n9819), .Z(n1898) );
  NANDN U4562 ( .A(n9820), .B(n1898), .Z(n1899) );
  NAND U4563 ( .A(n9818), .B(n9819), .Z(n1900) );
  AND U4564 ( .A(n1899), .B(n1900), .Z(n9977) );
  XNOR U4565 ( .A(n10471), .B(n10470), .Z(n10468) );
  XOR U4566 ( .A(n4947), .B(n4948), .Z(n1901) );
  NANDN U4567 ( .A(n4949), .B(n1901), .Z(n1902) );
  NAND U4568 ( .A(n4947), .B(n4948), .Z(n1903) );
  AND U4569 ( .A(n1902), .B(n1903), .Z(n4983) );
  XOR U4570 ( .A(n5075), .B(n5076), .Z(n1904) );
  NANDN U4571 ( .A(n5077), .B(n1904), .Z(n1905) );
  NAND U4572 ( .A(n5075), .B(n5076), .Z(n1906) );
  AND U4573 ( .A(n1905), .B(n1906), .Z(n5129) );
  NAND U4574 ( .A(n5263), .B(n5264), .Z(n1907) );
  XOR U4575 ( .A(n5263), .B(n5264), .Z(n1908) );
  NANDN U4576 ( .A(n5262), .B(n1908), .Z(n1909) );
  NAND U4577 ( .A(n1907), .B(n1909), .Z(n5342) );
  NAND U4578 ( .A(n5504), .B(n5505), .Z(n1910) );
  XOR U4579 ( .A(n5504), .B(n5505), .Z(n1911) );
  NANDN U4580 ( .A(n5503), .B(n1911), .Z(n1912) );
  NAND U4581 ( .A(n1910), .B(n1912), .Z(n5589) );
  XOR U4582 ( .A(n5791), .B(n5790), .Z(n1913) );
  NANDN U4583 ( .A(n5792), .B(n1913), .Z(n1914) );
  NAND U4584 ( .A(n5791), .B(n5790), .Z(n1915) );
  AND U4585 ( .A(n1914), .B(n1915), .Z(n5904) );
  XNOR U4586 ( .A(n6160), .B(n6159), .Z(n6153) );
  XOR U4587 ( .A(n7329), .B(n7330), .Z(n1916) );
  NANDN U4588 ( .A(n7331), .B(n1916), .Z(n1917) );
  NAND U4589 ( .A(n7329), .B(n7330), .Z(n1918) );
  AND U4590 ( .A(n1917), .B(n1918), .Z(n7340) );
  NAND U4591 ( .A(n7355), .B(n7354), .Z(n1919) );
  NANDN U4592 ( .A(n7353), .B(n7352), .Z(n1920) );
  AND U4593 ( .A(n1919), .B(n1920), .Z(n7517) );
  XOR U4594 ( .A(n2053), .B(n2054), .Z(n1921) );
  NANDN U4595 ( .A(n2055), .B(n1921), .Z(n1922) );
  NAND U4596 ( .A(n2053), .B(n2054), .Z(n1923) );
  AND U4597 ( .A(n1922), .B(n1923), .Z(n2103) );
  XOR U4598 ( .A(n2161), .B(n2162), .Z(n1924) );
  NANDN U4599 ( .A(n2163), .B(n1924), .Z(n1925) );
  NAND U4600 ( .A(n2161), .B(n2162), .Z(n1926) );
  AND U4601 ( .A(n1925), .B(n1926), .Z(n2263) );
  XNOR U4602 ( .A(n2586), .B(n2585), .Z(n2579) );
  XOR U4603 ( .A(n2774), .B(n2773), .Z(n1927) );
  NANDN U4604 ( .A(n2775), .B(n1927), .Z(n1928) );
  NAND U4605 ( .A(n2774), .B(n2773), .Z(n1929) );
  AND U4606 ( .A(n1928), .B(n1929), .Z(n2865) );
  XOR U4607 ( .A(n2986), .B(n2987), .Z(n1930) );
  NANDN U4608 ( .A(n2988), .B(n1930), .Z(n1931) );
  NAND U4609 ( .A(n2986), .B(n2987), .Z(n1932) );
  AND U4610 ( .A(n1931), .B(n1932), .Z(n3213) );
  NAND U4611 ( .A(n3609), .B(n3610), .Z(n1933) );
  XOR U4612 ( .A(n3609), .B(n3610), .Z(n1934) );
  NANDN U4613 ( .A(n3608), .B(n1934), .Z(n1935) );
  NAND U4614 ( .A(n1933), .B(n1935), .Z(n3744) );
  XOR U4615 ( .A(n3908), .B(n3909), .Z(n1936) );
  NANDN U4616 ( .A(n3910), .B(n1936), .Z(n1937) );
  NAND U4617 ( .A(n3908), .B(n3909), .Z(n1938) );
  AND U4618 ( .A(n1937), .B(n1938), .Z(n4066) );
  XNOR U4619 ( .A(n4559), .B(n4558), .Z(n4555) );
  NAND U4620 ( .A(n4392), .B(n4391), .Z(n1939) );
  NAND U4621 ( .A(n4390), .B(n4389), .Z(n1940) );
  AND U4622 ( .A(n1939), .B(n1940), .Z(n4849) );
  AND U4623 ( .A(x[480]), .B(y[7680]), .Z(n2595) );
  XOR U4624 ( .A(n2595), .B(o[0]), .Z(N33) );
  NAND U4625 ( .A(y[7680]), .B(x[481]), .Z(n1950) );
  AND U4626 ( .A(x[480]), .B(y[7681]), .Z(n1946) );
  XNOR U4627 ( .A(n1946), .B(o[1]), .Z(n1941) );
  XOR U4628 ( .A(n1950), .B(n1941), .Z(n1943) );
  NAND U4629 ( .A(n2595), .B(o[0]), .Z(n1942) );
  XNOR U4630 ( .A(n1943), .B(n1942), .Z(N34) );
  AND U4631 ( .A(x[480]), .B(y[7682]), .Z(n1947) );
  XNOR U4632 ( .A(n1947), .B(o[2]), .Z(n1955) );
  XNOR U4633 ( .A(n1956), .B(n1955), .Z(n1958) );
  AND U4634 ( .A(x[481]), .B(y[7681]), .Z(n1945) );
  NAND U4635 ( .A(x[482]), .B(y[7680]), .Z(n1944) );
  XNOR U4636 ( .A(n1945), .B(n1944), .Z(n1952) );
  AND U4637 ( .A(n1946), .B(o[1]), .Z(n1951) );
  XNOR U4638 ( .A(n1952), .B(n1951), .Z(n1957) );
  XNOR U4639 ( .A(n1958), .B(n1957), .Z(N35) );
  AND U4640 ( .A(x[481]), .B(y[7682]), .Z(n2069) );
  AND U4641 ( .A(y[7681]), .B(x[482]), .Z(n1974) );
  XOR U4642 ( .A(n1974), .B(o[3]), .Z(n1965) );
  XOR U4643 ( .A(n2069), .B(n1965), .Z(n1967) );
  AND U4644 ( .A(n1947), .B(o[2]), .Z(n1971) );
  AND U4645 ( .A(y[7680]), .B(x[483]), .Z(n1949) );
  AND U4646 ( .A(y[7683]), .B(x[480]), .Z(n1948) );
  XOR U4647 ( .A(n1949), .B(n1948), .Z(n1970) );
  XOR U4648 ( .A(n1971), .B(n1970), .Z(n1966) );
  XNOR U4649 ( .A(n1967), .B(n1966), .Z(n1964) );
  NANDN U4650 ( .A(n1950), .B(n1974), .Z(n1954) );
  NAND U4651 ( .A(n1952), .B(n1951), .Z(n1953) );
  NAND U4652 ( .A(n1954), .B(n1953), .Z(n1962) );
  NANDN U4653 ( .A(n1956), .B(n1955), .Z(n1960) );
  NAND U4654 ( .A(n1958), .B(n1957), .Z(n1959) );
  AND U4655 ( .A(n1960), .B(n1959), .Z(n1963) );
  XOR U4656 ( .A(n1962), .B(n1963), .Z(n1961) );
  XNOR U4657 ( .A(n1964), .B(n1961), .Z(N36) );
  NAND U4658 ( .A(n2069), .B(n1965), .Z(n1969) );
  NAND U4659 ( .A(n1967), .B(n1966), .Z(n1968) );
  NAND U4660 ( .A(n1969), .B(n1968), .Z(n1983) );
  XNOR U4661 ( .A(n1982), .B(n1983), .Z(n1985) );
  AND U4662 ( .A(x[483]), .B(y[7683]), .Z(n2017) );
  AND U4663 ( .A(y[7684]), .B(x[480]), .Z(n1973) );
  NAND U4664 ( .A(y[7680]), .B(x[484]), .Z(n1972) );
  XNOR U4665 ( .A(n1973), .B(n1972), .Z(n1998) );
  AND U4666 ( .A(n1974), .B(o[3]), .Z(n1999) );
  XOR U4667 ( .A(n1998), .B(n1999), .Z(n1977) );
  AND U4668 ( .A(x[482]), .B(y[7682]), .Z(n2129) );
  NAND U4669 ( .A(y[7683]), .B(x[481]), .Z(n1975) );
  XNOR U4670 ( .A(n2129), .B(n1975), .Z(n1995) );
  AND U4671 ( .A(y[7681]), .B(x[483]), .Z(n1992) );
  XOR U4672 ( .A(o[4]), .B(n1992), .Z(n1994) );
  XOR U4673 ( .A(n1995), .B(n1994), .Z(n1976) );
  XNOR U4674 ( .A(n1977), .B(n1976), .Z(n1979) );
  XOR U4675 ( .A(n1978), .B(n1979), .Z(n1984) );
  XNOR U4676 ( .A(n1985), .B(n1984), .Z(N37) );
  NAND U4677 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U4678 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U4679 ( .A(n1981), .B(n1980), .Z(n2026) );
  NANDN U4680 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U4681 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U4682 ( .A(n1987), .B(n1986), .Z(n2025) );
  AND U4683 ( .A(y[7682]), .B(x[483]), .Z(n1989) );
  NAND U4684 ( .A(y[7684]), .B(x[481]), .Z(n1988) );
  XNOR U4685 ( .A(n1989), .B(n1988), .Z(n2004) );
  AND U4686 ( .A(x[484]), .B(y[7681]), .Z(n2015) );
  XOR U4687 ( .A(n2015), .B(o[5]), .Z(n2003) );
  XNOR U4688 ( .A(n2004), .B(n2003), .Z(n2007) );
  NAND U4689 ( .A(x[482]), .B(y[7683]), .Z(n2078) );
  AND U4690 ( .A(x[485]), .B(y[7680]), .Z(n1991) );
  NAND U4691 ( .A(y[7685]), .B(x[480]), .Z(n1990) );
  XNOR U4692 ( .A(n1991), .B(n1990), .Z(n2010) );
  AND U4693 ( .A(o[4]), .B(n1992), .Z(n2009) );
  XOR U4694 ( .A(n2010), .B(n2009), .Z(n2008) );
  XOR U4695 ( .A(n2078), .B(n2008), .Z(n1993) );
  XOR U4696 ( .A(n2007), .B(n1993), .Z(n2022) );
  NANDN U4697 ( .A(n2078), .B(n2069), .Z(n1997) );
  NAND U4698 ( .A(n1995), .B(n1994), .Z(n1996) );
  NAND U4699 ( .A(n1997), .B(n1996), .Z(n2020) );
  AND U4700 ( .A(x[484]), .B(y[7684]), .Z(n2793) );
  NAND U4701 ( .A(n2793), .B(n2595), .Z(n2001) );
  NAND U4702 ( .A(n1999), .B(n1998), .Z(n2000) );
  NAND U4703 ( .A(n2001), .B(n2000), .Z(n2019) );
  XOR U4704 ( .A(n2020), .B(n2019), .Z(n2021) );
  XOR U4705 ( .A(n2022), .B(n2021), .Z(n2027) );
  XOR U4706 ( .A(n2025), .B(n2027), .Z(n2002) );
  XOR U4707 ( .A(n2026), .B(n2002), .Z(N38) );
  AND U4708 ( .A(x[483]), .B(y[7684]), .Z(n2079) );
  NAND U4709 ( .A(n2079), .B(n2069), .Z(n2006) );
  NAND U4710 ( .A(n2004), .B(n2003), .Z(n2005) );
  NAND U4711 ( .A(n2006), .B(n2005), .Z(n2057) );
  XOR U4712 ( .A(n2057), .B(n2056), .Z(n2059) );
  AND U4713 ( .A(y[7685]), .B(x[485]), .Z(n2251) );
  NAND U4714 ( .A(n2595), .B(n2251), .Z(n2012) );
  NAND U4715 ( .A(n2010), .B(n2009), .Z(n2011) );
  AND U4716 ( .A(n2012), .B(n2011), .Z(n2030) );
  AND U4717 ( .A(x[486]), .B(y[7680]), .Z(n2014) );
  NAND U4718 ( .A(x[480]), .B(y[7686]), .Z(n2013) );
  XNOR U4719 ( .A(n2014), .B(n2013), .Z(n2036) );
  AND U4720 ( .A(n2015), .B(o[5]), .Z(n2037) );
  XOR U4721 ( .A(n2036), .B(n2037), .Z(n2029) );
  NAND U4722 ( .A(y[7684]), .B(x[482]), .Z(n2016) );
  XNOR U4723 ( .A(n2017), .B(n2016), .Z(n2041) );
  AND U4724 ( .A(y[7685]), .B(x[481]), .Z(n2298) );
  NAND U4725 ( .A(y[7682]), .B(x[484]), .Z(n2018) );
  XNOR U4726 ( .A(n2298), .B(n2018), .Z(n2045) );
  AND U4727 ( .A(y[7681]), .B(x[485]), .Z(n2052) );
  XOR U4728 ( .A(o[6]), .B(n2052), .Z(n2044) );
  XOR U4729 ( .A(n2045), .B(n2044), .Z(n2040) );
  XOR U4730 ( .A(n2041), .B(n2040), .Z(n2031) );
  XOR U4731 ( .A(n2032), .B(n2031), .Z(n2058) );
  XNOR U4732 ( .A(n2059), .B(n2058), .Z(n2055) );
  NAND U4733 ( .A(n2020), .B(n2019), .Z(n2024) );
  NAND U4734 ( .A(n2022), .B(n2021), .Z(n2023) );
  NAND U4735 ( .A(n2024), .B(n2023), .Z(n2054) );
  XOR U4736 ( .A(n2054), .B(n2053), .Z(n2028) );
  XNOR U4737 ( .A(n2055), .B(n2028), .Z(N39) );
  NANDN U4738 ( .A(n2030), .B(n2029), .Z(n2034) );
  NAND U4739 ( .A(n2032), .B(n2031), .Z(n2033) );
  AND U4740 ( .A(n2034), .B(n2033), .Z(n2099) );
  AND U4741 ( .A(x[485]), .B(y[7682]), .Z(n2170) );
  NAND U4742 ( .A(x[481]), .B(y[7686]), .Z(n2035) );
  XNOR U4743 ( .A(n2170), .B(n2035), .Z(n2072) );
  NAND U4744 ( .A(y[7681]), .B(x[486]), .Z(n2076) );
  XNOR U4745 ( .A(n2072), .B(n2071), .Z(n2091) );
  AND U4746 ( .A(y[7686]), .B(x[486]), .Z(n2317) );
  NAND U4747 ( .A(n2595), .B(n2317), .Z(n2039) );
  NAND U4748 ( .A(n2037), .B(n2036), .Z(n2038) );
  AND U4749 ( .A(n2039), .B(n2038), .Z(n2090) );
  XOR U4750 ( .A(n2091), .B(n2090), .Z(n2092) );
  NANDN U4751 ( .A(n2078), .B(n2079), .Z(n2043) );
  NAND U4752 ( .A(n2041), .B(n2040), .Z(n2042) );
  AND U4753 ( .A(n2043), .B(n2042), .Z(n2093) );
  XOR U4754 ( .A(n2092), .B(n2093), .Z(n2097) );
  AND U4755 ( .A(x[484]), .B(y[7685]), .Z(n2600) );
  NAND U4756 ( .A(n2600), .B(n2069), .Z(n2047) );
  NAND U4757 ( .A(n2045), .B(n2044), .Z(n2046) );
  AND U4758 ( .A(n2047), .B(n2046), .Z(n2066) );
  AND U4759 ( .A(y[7685]), .B(x[482]), .Z(n2049) );
  NAND U4760 ( .A(y[7683]), .B(x[484]), .Z(n2048) );
  XNOR U4761 ( .A(n2049), .B(n2048), .Z(n2080) );
  XNOR U4762 ( .A(n2080), .B(n2079), .Z(n2064) );
  AND U4763 ( .A(x[487]), .B(y[7680]), .Z(n2051) );
  NAND U4764 ( .A(y[7687]), .B(x[480]), .Z(n2050) );
  XNOR U4765 ( .A(n2051), .B(n2050), .Z(n2085) );
  AND U4766 ( .A(o[6]), .B(n2052), .Z(n2084) );
  XNOR U4767 ( .A(n2085), .B(n2084), .Z(n2063) );
  XOR U4768 ( .A(n2064), .B(n2063), .Z(n2065) );
  XOR U4769 ( .A(n2066), .B(n2065), .Z(n2096) );
  XOR U4770 ( .A(n2097), .B(n2096), .Z(n2098) );
  XNOR U4771 ( .A(n2099), .B(n2098), .Z(n2105) );
  NAND U4772 ( .A(n2057), .B(n2056), .Z(n2061) );
  NAND U4773 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U4774 ( .A(n2061), .B(n2060), .Z(n2104) );
  IV U4775 ( .A(n2104), .Z(n2102) );
  XOR U4776 ( .A(n2103), .B(n2102), .Z(n2062) );
  XNOR U4777 ( .A(n2105), .B(n2062), .Z(N40) );
  NAND U4778 ( .A(n2064), .B(n2063), .Z(n2068) );
  NAND U4779 ( .A(n2066), .B(n2065), .Z(n2067) );
  AND U4780 ( .A(n2068), .B(n2067), .Z(n2142) );
  AND U4781 ( .A(y[7686]), .B(x[485]), .Z(n2070) );
  NAND U4782 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U4783 ( .A(n2072), .B(n2071), .Z(n2073) );
  AND U4784 ( .A(n2074), .B(n2073), .Z(n2140) );
  AND U4785 ( .A(x[485]), .B(y[7683]), .Z(n2735) );
  NAND U4786 ( .A(x[481]), .B(y[7687]), .Z(n2075) );
  XNOR U4787 ( .A(n2735), .B(n2075), .Z(n2121) );
  ANDN U4788 ( .B(o[7]), .A(n2076), .Z(n2120) );
  XNOR U4789 ( .A(n2121), .B(n2120), .Z(n2125) );
  NAND U4790 ( .A(x[483]), .B(y[7685]), .Z(n2918) );
  AND U4791 ( .A(y[7682]), .B(x[486]), .Z(n2077) );
  AND U4792 ( .A(x[482]), .B(y[7686]), .Z(n3024) );
  XOR U4793 ( .A(n2077), .B(n3024), .Z(n2130) );
  XOR U4794 ( .A(n2793), .B(n2130), .Z(n2124) );
  XOR U4795 ( .A(n2125), .B(n2126), .Z(n2139) );
  XOR U4796 ( .A(n2142), .B(n2141), .Z(n2151) );
  NANDN U4797 ( .A(n2078), .B(n2600), .Z(n2082) );
  NAND U4798 ( .A(n2080), .B(n2079), .Z(n2081) );
  AND U4799 ( .A(n2082), .B(n2081), .Z(n2136) );
  AND U4800 ( .A(y[7687]), .B(x[487]), .Z(n2083) );
  NAND U4801 ( .A(n2595), .B(n2083), .Z(n2087) );
  NAND U4802 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U4803 ( .A(n2087), .B(n2086), .Z(n2134) );
  AND U4804 ( .A(x[488]), .B(y[7680]), .Z(n2089) );
  NAND U4805 ( .A(y[7688]), .B(x[480]), .Z(n2088) );
  XNOR U4806 ( .A(n2089), .B(n2088), .Z(n2112) );
  NAND U4807 ( .A(y[7681]), .B(x[487]), .Z(n2116) );
  XOR U4808 ( .A(n2112), .B(n2111), .Z(n2133) );
  NAND U4809 ( .A(n2091), .B(n2090), .Z(n2095) );
  NAND U4810 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U4811 ( .A(n2095), .B(n2094), .Z(n2148) );
  XOR U4812 ( .A(n2149), .B(n2148), .Z(n2150) );
  XOR U4813 ( .A(n2151), .B(n2150), .Z(n2147) );
  NAND U4814 ( .A(n2097), .B(n2096), .Z(n2101) );
  NAND U4815 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U4816 ( .A(n2101), .B(n2100), .Z(n2145) );
  NANDN U4817 ( .A(n2102), .B(n2103), .Z(n2108) );
  NOR U4818 ( .A(n2104), .B(n2103), .Z(n2106) );
  OR U4819 ( .A(n2106), .B(n2105), .Z(n2107) );
  AND U4820 ( .A(n2108), .B(n2107), .Z(n2146) );
  XOR U4821 ( .A(n2145), .B(n2146), .Z(n2109) );
  XNOR U4822 ( .A(n2147), .B(n2109), .Z(N41) );
  AND U4823 ( .A(x[488]), .B(y[7688]), .Z(n2110) );
  NAND U4824 ( .A(n2110), .B(n2595), .Z(n2114) );
  NAND U4825 ( .A(n2112), .B(n2111), .Z(n2113) );
  AND U4826 ( .A(n2114), .B(n2113), .Z(n2200) );
  AND U4827 ( .A(y[7682]), .B(x[487]), .Z(n2524) );
  NAND U4828 ( .A(x[485]), .B(y[7684]), .Z(n2115) );
  XNOR U4829 ( .A(n2524), .B(n2115), .Z(n2172) );
  ANDN U4830 ( .B(o[8]), .A(n2116), .Z(n2171) );
  XOR U4831 ( .A(n2172), .B(n2171), .Z(n2198) );
  AND U4832 ( .A(x[489]), .B(y[7680]), .Z(n2118) );
  NAND U4833 ( .A(y[7689]), .B(x[480]), .Z(n2117) );
  XNOR U4834 ( .A(n2118), .B(n2117), .Z(n2179) );
  AND U4835 ( .A(y[7681]), .B(x[488]), .Z(n2189) );
  XOR U4836 ( .A(o[9]), .B(n2189), .Z(n2178) );
  XNOR U4837 ( .A(n2179), .B(n2178), .Z(n2197) );
  XNOR U4838 ( .A(n2200), .B(n2199), .Z(n2194) );
  AND U4839 ( .A(y[7683]), .B(x[486]), .Z(n2538) );
  NAND U4840 ( .A(y[7688]), .B(x[481]), .Z(n2119) );
  XNOR U4841 ( .A(n2538), .B(n2119), .Z(n2184) );
  XOR U4842 ( .A(n2600), .B(n2184), .Z(n2204) );
  AND U4843 ( .A(y[7687]), .B(x[482]), .Z(n2838) );
  AND U4844 ( .A(y[7686]), .B(x[483]), .Z(n2549) );
  XOR U4845 ( .A(n2838), .B(n2549), .Z(n2203) );
  NAND U4846 ( .A(y[7687]), .B(x[485]), .Z(n2371) );
  AND U4847 ( .A(x[481]), .B(y[7683]), .Z(n2182) );
  NANDN U4848 ( .A(n2371), .B(n2182), .Z(n2123) );
  NAND U4849 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U4850 ( .A(n2123), .B(n2122), .Z(n2191) );
  XOR U4851 ( .A(n2192), .B(n2191), .Z(n2193) );
  XNOR U4852 ( .A(n2194), .B(n2193), .Z(n2166) );
  NANDN U4853 ( .A(n2124), .B(n2918), .Z(n2128) );
  NANDN U4854 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U4855 ( .A(n2128), .B(n2127), .Z(n2164) );
  NAND U4856 ( .A(n2317), .B(n2129), .Z(n2132) );
  NAND U4857 ( .A(n2793), .B(n2130), .Z(n2131) );
  AND U4858 ( .A(n2132), .B(n2131), .Z(n2165) );
  XNOR U4859 ( .A(n2164), .B(n2165), .Z(n2167) );
  NANDN U4860 ( .A(n2134), .B(n2133), .Z(n2138) );
  NANDN U4861 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U4862 ( .A(n2138), .B(n2137), .Z(n2156) );
  NANDN U4863 ( .A(n2140), .B(n2139), .Z(n2144) );
  NAND U4864 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U4865 ( .A(n2144), .B(n2143), .Z(n2155) );
  XNOR U4866 ( .A(n2157), .B(n2158), .Z(n2163) );
  NAND U4867 ( .A(n2149), .B(n2148), .Z(n2153) );
  NANDN U4868 ( .A(n2151), .B(n2150), .Z(n2152) );
  AND U4869 ( .A(n2153), .B(n2152), .Z(n2162) );
  XOR U4870 ( .A(n2161), .B(n2162), .Z(n2154) );
  XNOR U4871 ( .A(n2163), .B(n2154), .Z(N42) );
  NANDN U4872 ( .A(n2156), .B(n2155), .Z(n2160) );
  NAND U4873 ( .A(n2158), .B(n2157), .Z(n2159) );
  NAND U4874 ( .A(n2160), .B(n2159), .Z(n2262) );
  IV U4875 ( .A(n2262), .Z(n2261) );
  NAND U4876 ( .A(n2165), .B(n2164), .Z(n2169) );
  NANDN U4877 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U4878 ( .A(n2169), .B(n2168), .Z(n2270) );
  AND U4879 ( .A(y[7684]), .B(x[487]), .Z(n2245) );
  NAND U4880 ( .A(n2245), .B(n2170), .Z(n2174) );
  NAND U4881 ( .A(n2172), .B(n2171), .Z(n2173) );
  AND U4882 ( .A(n2174), .B(n2173), .Z(n2258) );
  AND U4883 ( .A(x[487]), .B(y[7683]), .Z(n2176) );
  NAND U4884 ( .A(x[484]), .B(y[7686]), .Z(n2175) );
  XNOR U4885 ( .A(n2176), .B(n2175), .Z(n2228) );
  AND U4886 ( .A(y[7684]), .B(x[486]), .Z(n2229) );
  XOR U4887 ( .A(n2228), .B(n2229), .Z(n2256) );
  AND U4888 ( .A(x[488]), .B(y[7682]), .Z(n2444) );
  AND U4889 ( .A(y[7681]), .B(x[489]), .Z(n2239) );
  XOR U4890 ( .A(o[10]), .B(n2239), .Z(n2250) );
  XOR U4891 ( .A(n2444), .B(n2250), .Z(n2252) );
  XNOR U4892 ( .A(n2252), .B(n2251), .Z(n2255) );
  XOR U4893 ( .A(n2258), .B(n2257), .Z(n2217) );
  AND U4894 ( .A(x[489]), .B(y[7689]), .Z(n2177) );
  NAND U4895 ( .A(n2177), .B(n2595), .Z(n2181) );
  NAND U4896 ( .A(n2179), .B(n2178), .Z(n2180) );
  AND U4897 ( .A(n2181), .B(n2180), .Z(n2215) );
  AND U4898 ( .A(y[7688]), .B(x[486]), .Z(n2183) );
  NAND U4899 ( .A(n2183), .B(n2182), .Z(n2186) );
  NAND U4900 ( .A(n2600), .B(n2184), .Z(n2185) );
  NAND U4901 ( .A(n2186), .B(n2185), .Z(n2223) );
  AND U4902 ( .A(x[490]), .B(y[7680]), .Z(n2188) );
  NAND U4903 ( .A(y[7690]), .B(x[480]), .Z(n2187) );
  XNOR U4904 ( .A(n2188), .B(n2187), .Z(n2234) );
  AND U4905 ( .A(o[9]), .B(n2189), .Z(n2233) );
  XOR U4906 ( .A(n2234), .B(n2233), .Z(n2221) );
  AND U4907 ( .A(y[7689]), .B(x[481]), .Z(n3104) );
  NAND U4908 ( .A(x[483]), .B(y[7687]), .Z(n2190) );
  XNOR U4909 ( .A(n3104), .B(n2190), .Z(n2246) );
  AND U4910 ( .A(y[7688]), .B(x[482]), .Z(n2247) );
  XOR U4911 ( .A(n2246), .B(n2247), .Z(n2220) );
  XOR U4912 ( .A(n2221), .B(n2220), .Z(n2222) );
  XOR U4913 ( .A(n2223), .B(n2222), .Z(n2214) );
  NAND U4914 ( .A(n2192), .B(n2191), .Z(n2196) );
  NAND U4915 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U4916 ( .A(n2196), .B(n2195), .Z(n2211) );
  NANDN U4917 ( .A(n2198), .B(n2197), .Z(n2202) );
  NAND U4918 ( .A(n2200), .B(n2199), .Z(n2201) );
  AND U4919 ( .A(n2202), .B(n2201), .Z(n2208) );
  NOR U4920 ( .A(n2549), .B(n2838), .Z(n2206) );
  NANDN U4921 ( .A(n2204), .B(n2203), .Z(n2205) );
  NANDN U4922 ( .A(n2206), .B(n2205), .Z(n2209) );
  XOR U4923 ( .A(n2211), .B(n2210), .Z(n2268) );
  XOR U4924 ( .A(n2270), .B(n2271), .Z(n2264) );
  XNOR U4925 ( .A(n2263), .B(n2264), .Z(n2207) );
  XOR U4926 ( .A(n2261), .B(n2207), .Z(N43) );
  NANDN U4927 ( .A(n2209), .B(n2208), .Z(n2213) );
  NANDN U4928 ( .A(n2211), .B(n2210), .Z(n2212) );
  AND U4929 ( .A(n2213), .B(n2212), .Z(n2278) );
  NANDN U4930 ( .A(n2215), .B(n2214), .Z(n2219) );
  NANDN U4931 ( .A(n2217), .B(n2216), .Z(n2218) );
  AND U4932 ( .A(n2219), .B(n2218), .Z(n2276) );
  NAND U4933 ( .A(n2221), .B(n2220), .Z(n2225) );
  NAND U4934 ( .A(n2223), .B(n2222), .Z(n2224) );
  NAND U4935 ( .A(n2225), .B(n2224), .Z(n2339) );
  AND U4936 ( .A(y[7686]), .B(x[487]), .Z(n2227) );
  AND U4937 ( .A(x[484]), .B(y[7683]), .Z(n2226) );
  NAND U4938 ( .A(n2227), .B(n2226), .Z(n2231) );
  NAND U4939 ( .A(n2229), .B(n2228), .Z(n2230) );
  NAND U4940 ( .A(n2231), .B(n2230), .Z(n2337) );
  AND U4941 ( .A(x[490]), .B(y[7690]), .Z(n2232) );
  NAND U4942 ( .A(n2232), .B(n2595), .Z(n2236) );
  NAND U4943 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U4944 ( .A(n2236), .B(n2235), .Z(n2333) );
  AND U4945 ( .A(x[491]), .B(y[7680]), .Z(n2238) );
  NAND U4946 ( .A(x[480]), .B(y[7691]), .Z(n2237) );
  XNOR U4947 ( .A(n2238), .B(n2237), .Z(n2309) );
  AND U4948 ( .A(o[10]), .B(n2239), .Z(n2308) );
  XOR U4949 ( .A(n2309), .B(n2308), .Z(n2331) );
  AND U4950 ( .A(x[486]), .B(y[7685]), .Z(n2241) );
  NAND U4951 ( .A(y[7690]), .B(x[481]), .Z(n2240) );
  XNOR U4952 ( .A(n2241), .B(n2240), .Z(n2300) );
  NAND U4953 ( .A(y[7681]), .B(x[490]), .Z(n2318) );
  XOR U4954 ( .A(n2300), .B(n2299), .Z(n2330) );
  XOR U4955 ( .A(n2331), .B(n2330), .Z(n2332) );
  XOR U4956 ( .A(n2333), .B(n2332), .Z(n2336) );
  XOR U4957 ( .A(n2337), .B(n2336), .Z(n2338) );
  XNOR U4958 ( .A(n2339), .B(n2338), .Z(n2321) );
  NAND U4959 ( .A(y[7688]), .B(x[483]), .Z(n3307) );
  AND U4960 ( .A(x[482]), .B(y[7689]), .Z(n2243) );
  NAND U4961 ( .A(x[485]), .B(y[7686]), .Z(n2242) );
  XNOR U4962 ( .A(n2243), .B(n2242), .Z(n2295) );
  AND U4963 ( .A(x[484]), .B(y[7687]), .Z(n2294) );
  XNOR U4964 ( .A(n2295), .B(n2294), .Z(n2325) );
  XOR U4965 ( .A(n3307), .B(n2325), .Z(n2327) );
  NAND U4966 ( .A(y[7682]), .B(x[489]), .Z(n2244) );
  XNOR U4967 ( .A(n2245), .B(n2244), .Z(n2313) );
  AND U4968 ( .A(x[488]), .B(y[7683]), .Z(n2312) );
  XNOR U4969 ( .A(n2313), .B(n2312), .Z(n2326) );
  XNOR U4970 ( .A(n2327), .B(n2326), .Z(n2291) );
  NAND U4971 ( .A(y[7689]), .B(x[483]), .Z(n2362) );
  AND U4972 ( .A(y[7687]), .B(x[481]), .Z(n2590) );
  NANDN U4973 ( .A(n2362), .B(n2590), .Z(n2249) );
  NAND U4974 ( .A(n2247), .B(n2246), .Z(n2248) );
  NAND U4975 ( .A(n2249), .B(n2248), .Z(n2289) );
  NAND U4976 ( .A(n2444), .B(n2250), .Z(n2254) );
  NAND U4977 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U4978 ( .A(n2254), .B(n2253), .Z(n2288) );
  XOR U4979 ( .A(n2289), .B(n2288), .Z(n2290) );
  XOR U4980 ( .A(n2291), .B(n2290), .Z(n2320) );
  NANDN U4981 ( .A(n2256), .B(n2255), .Z(n2260) );
  NAND U4982 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U4983 ( .A(n2260), .B(n2259), .Z(n2319) );
  XOR U4984 ( .A(n2321), .B(n2322), .Z(n2275) );
  XOR U4985 ( .A(n2278), .B(n2277), .Z(n2284) );
  OR U4986 ( .A(n2263), .B(n2261), .Z(n2267) );
  ANDN U4987 ( .B(n2263), .A(n2262), .Z(n2265) );
  OR U4988 ( .A(n2265), .B(n2264), .Z(n2266) );
  AND U4989 ( .A(n2267), .B(n2266), .Z(n2283) );
  NANDN U4990 ( .A(n2269), .B(n2268), .Z(n2273) );
  NAND U4991 ( .A(n2271), .B(n2270), .Z(n2272) );
  AND U4992 ( .A(n2273), .B(n2272), .Z(n2282) );
  IV U4993 ( .A(n2282), .Z(n2281) );
  XOR U4994 ( .A(n2283), .B(n2281), .Z(n2274) );
  XNOR U4995 ( .A(n2284), .B(n2274), .Z(N44) );
  NANDN U4996 ( .A(n2276), .B(n2275), .Z(n2280) );
  NANDN U4997 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U4998 ( .A(n2280), .B(n2279), .Z(n2406) );
  IV U4999 ( .A(n2406), .Z(n2405) );
  OR U5000 ( .A(n2283), .B(n2281), .Z(n2287) );
  ANDN U5001 ( .B(n2283), .A(n2282), .Z(n2285) );
  OR U5002 ( .A(n2285), .B(n2284), .Z(n2286) );
  AND U5003 ( .A(n2287), .B(n2286), .Z(n2407) );
  NAND U5004 ( .A(n2289), .B(n2288), .Z(n2293) );
  NAND U5005 ( .A(n2291), .B(n2290), .Z(n2292) );
  NAND U5006 ( .A(n2293), .B(n2292), .Z(n2402) );
  AND U5007 ( .A(y[7689]), .B(x[485]), .Z(n2831) );
  NAND U5008 ( .A(n3024), .B(n2831), .Z(n2297) );
  NAND U5009 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U5010 ( .A(n2297), .B(n2296), .Z(n2350) );
  AND U5011 ( .A(x[486]), .B(y[7690]), .Z(n2607) );
  NAND U5012 ( .A(n2607), .B(n2298), .Z(n2302) );
  NAND U5013 ( .A(n2300), .B(n2299), .Z(n2301) );
  NAND U5014 ( .A(n2302), .B(n2301), .Z(n2349) );
  XOR U5015 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U5016 ( .A(x[489]), .B(y[7683]), .Z(n3019) );
  AND U5017 ( .A(y[7682]), .B(x[490]), .Z(n3063) );
  NAND U5018 ( .A(y[7688]), .B(x[484]), .Z(n2303) );
  XOR U5019 ( .A(n3063), .B(n2303), .Z(n2392) );
  NAND U5020 ( .A(x[487]), .B(y[7685]), .Z(n2370) );
  XOR U5021 ( .A(n2371), .B(n2370), .Z(n2373) );
  AND U5022 ( .A(x[492]), .B(y[7680]), .Z(n2305) );
  NAND U5023 ( .A(y[7692]), .B(x[480]), .Z(n2304) );
  XNOR U5024 ( .A(n2305), .B(n2304), .Z(n2387) );
  NAND U5025 ( .A(y[7681]), .B(x[491]), .Z(n2367) );
  XOR U5026 ( .A(n2387), .B(n2386), .Z(n2356) );
  AND U5027 ( .A(y[7690]), .B(x[482]), .Z(n2307) );
  NAND U5028 ( .A(y[7684]), .B(x[488]), .Z(n2306) );
  XNOR U5029 ( .A(n2307), .B(n2306), .Z(n2361) );
  XOR U5030 ( .A(n2356), .B(n2355), .Z(n2357) );
  XNOR U5031 ( .A(n2351), .B(n2352), .Z(n2400) );
  AND U5032 ( .A(y[7691]), .B(x[491]), .Z(n3387) );
  NAND U5033 ( .A(n3387), .B(n2595), .Z(n2311) );
  NAND U5034 ( .A(n2309), .B(n2308), .Z(n2310) );
  NAND U5035 ( .A(n2311), .B(n2310), .Z(n2379) );
  AND U5036 ( .A(x[489]), .B(y[7684]), .Z(n2369) );
  NAND U5037 ( .A(n2524), .B(n2369), .Z(n2315) );
  NAND U5038 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U5039 ( .A(n2315), .B(n2314), .Z(n2377) );
  NAND U5040 ( .A(x[481]), .B(y[7691]), .Z(n2316) );
  XNOR U5041 ( .A(n2317), .B(n2316), .Z(n2383) );
  ANDN U5042 ( .B(o[11]), .A(n2318), .Z(n2382) );
  XOR U5043 ( .A(n2383), .B(n2382), .Z(n2376) );
  XOR U5044 ( .A(n2377), .B(n2376), .Z(n2378) );
  XOR U5045 ( .A(n2379), .B(n2378), .Z(n2399) );
  XOR U5046 ( .A(n2400), .B(n2399), .Z(n2401) );
  XOR U5047 ( .A(n2402), .B(n2401), .Z(n2413) );
  NANDN U5048 ( .A(n2320), .B(n2319), .Z(n2324) );
  NANDN U5049 ( .A(n2322), .B(n2321), .Z(n2323) );
  NAND U5050 ( .A(n2324), .B(n2323), .Z(n2412) );
  IV U5051 ( .A(n3307), .Z(n3033) );
  NANDN U5052 ( .A(n3033), .B(n2325), .Z(n2329) );
  NAND U5053 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U5054 ( .A(n2329), .B(n2328), .Z(n2344) );
  NAND U5055 ( .A(n2331), .B(n2330), .Z(n2335) );
  NAND U5056 ( .A(n2333), .B(n2332), .Z(n2334) );
  AND U5057 ( .A(n2335), .B(n2334), .Z(n2343) );
  XOR U5058 ( .A(n2344), .B(n2343), .Z(n2346) );
  NAND U5059 ( .A(n2337), .B(n2336), .Z(n2341) );
  NAND U5060 ( .A(n2339), .B(n2338), .Z(n2340) );
  AND U5061 ( .A(n2341), .B(n2340), .Z(n2345) );
  XOR U5062 ( .A(n2346), .B(n2345), .Z(n2414) );
  XOR U5063 ( .A(n2415), .B(n2414), .Z(n2408) );
  XNOR U5064 ( .A(n2407), .B(n2408), .Z(n2342) );
  XOR U5065 ( .A(n2405), .B(n2342), .Z(N45) );
  NAND U5066 ( .A(n2344), .B(n2343), .Z(n2348) );
  NAND U5067 ( .A(n2346), .B(n2345), .Z(n2347) );
  NAND U5068 ( .A(n2348), .B(n2347), .Z(n2422) );
  NAND U5069 ( .A(n2350), .B(n2349), .Z(n2354) );
  NANDN U5070 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND U5071 ( .A(n2354), .B(n2353), .Z(n2487) );
  NAND U5072 ( .A(n2356), .B(n2355), .Z(n2360) );
  NANDN U5073 ( .A(n2358), .B(n2357), .Z(n2359) );
  NAND U5074 ( .A(n2360), .B(n2359), .Z(n2495) );
  AND U5075 ( .A(y[7690]), .B(x[488]), .Z(n3670) );
  AND U5076 ( .A(x[482]), .B(y[7684]), .Z(n2534) );
  NAND U5077 ( .A(n3670), .B(n2534), .Z(n2364) );
  NANDN U5078 ( .A(n2362), .B(n2361), .Z(n2363) );
  AND U5079 ( .A(n2364), .B(n2363), .Z(n2460) );
  AND U5080 ( .A(y[7692]), .B(x[481]), .Z(n2366) );
  NAND U5081 ( .A(x[487]), .B(y[7686]), .Z(n2365) );
  XNOR U5082 ( .A(n2366), .B(n2365), .Z(n2450) );
  ANDN U5083 ( .B(o[12]), .A(n2367), .Z(n2449) );
  XOR U5084 ( .A(n2450), .B(n2449), .Z(n2458) );
  AND U5085 ( .A(y[7687]), .B(x[486]), .Z(n3426) );
  NAND U5086 ( .A(x[482]), .B(y[7691]), .Z(n2368) );
  XOR U5087 ( .A(n2369), .B(n2368), .Z(n2464) );
  XOR U5088 ( .A(n2458), .B(n2457), .Z(n2459) );
  NAND U5089 ( .A(n2371), .B(n2370), .Z(n2375) );
  ANDN U5090 ( .B(n2373), .A(n2372), .Z(n2374) );
  ANDN U5091 ( .B(n2375), .A(n2374), .Z(n2493) );
  XOR U5092 ( .A(n2494), .B(n2493), .Z(n2496) );
  XOR U5093 ( .A(n2495), .B(n2496), .Z(n2488) );
  XOR U5094 ( .A(n2487), .B(n2488), .Z(n2490) );
  NAND U5095 ( .A(n2377), .B(n2376), .Z(n2381) );
  NAND U5096 ( .A(n2379), .B(n2378), .Z(n2380) );
  AND U5097 ( .A(n2381), .B(n2380), .Z(n2435) );
  NAND U5098 ( .A(y[7691]), .B(x[486]), .Z(n2833) );
  AND U5099 ( .A(y[7686]), .B(x[481]), .Z(n2448) );
  NANDN U5100 ( .A(n2833), .B(n2448), .Z(n2385) );
  NAND U5101 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U5102 ( .A(n2385), .B(n2384), .Z(n2441) );
  AND U5103 ( .A(x[492]), .B(y[7692]), .Z(n3678) );
  NAND U5104 ( .A(n3678), .B(n2595), .Z(n2389) );
  NAND U5105 ( .A(n2387), .B(n2386), .Z(n2388) );
  AND U5106 ( .A(n2389), .B(n2388), .Z(n2439) );
  AND U5107 ( .A(x[490]), .B(y[7683]), .Z(n3319) );
  AND U5108 ( .A(y[7682]), .B(x[491]), .Z(n3268) );
  NAND U5109 ( .A(y[7685]), .B(x[488]), .Z(n2390) );
  XOR U5110 ( .A(n3268), .B(n2390), .Z(n2445) );
  AND U5111 ( .A(x[490]), .B(y[7688]), .Z(n2799) );
  AND U5112 ( .A(x[484]), .B(y[7682]), .Z(n2391) );
  NAND U5113 ( .A(n2799), .B(n2391), .Z(n2394) );
  NANDN U5114 ( .A(n2392), .B(n3019), .Z(n2393) );
  AND U5115 ( .A(n2394), .B(n2393), .Z(n2484) );
  AND U5116 ( .A(x[493]), .B(y[7680]), .Z(n2396) );
  NAND U5117 ( .A(y[7693]), .B(x[480]), .Z(n2395) );
  XNOR U5118 ( .A(n2396), .B(n2395), .Z(n2476) );
  AND U5119 ( .A(y[7681]), .B(x[492]), .Z(n2469) );
  XOR U5120 ( .A(o[13]), .B(n2469), .Z(n2475) );
  XOR U5121 ( .A(n2476), .B(n2475), .Z(n2482) );
  AND U5122 ( .A(y[7690]), .B(x[483]), .Z(n2398) );
  NAND U5123 ( .A(x[485]), .B(y[7688]), .Z(n2397) );
  XNOR U5124 ( .A(n2398), .B(n2397), .Z(n2471) );
  NAND U5125 ( .A(x[484]), .B(y[7689]), .Z(n2472) );
  XOR U5126 ( .A(n2482), .B(n2481), .Z(n2483) );
  XOR U5127 ( .A(n2433), .B(n2432), .Z(n2434) );
  XNOR U5128 ( .A(n2490), .B(n2489), .Z(n2420) );
  NAND U5129 ( .A(n2400), .B(n2399), .Z(n2404) );
  NAND U5130 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U5131 ( .A(n2404), .B(n2403), .Z(n2419) );
  XOR U5132 ( .A(n2420), .B(n2419), .Z(n2421) );
  XOR U5133 ( .A(n2422), .B(n2421), .Z(n2428) );
  OR U5134 ( .A(n2407), .B(n2405), .Z(n2411) );
  ANDN U5135 ( .B(n2407), .A(n2406), .Z(n2409) );
  OR U5136 ( .A(n2409), .B(n2408), .Z(n2410) );
  AND U5137 ( .A(n2411), .B(n2410), .Z(n2427) );
  NANDN U5138 ( .A(n2413), .B(n2412), .Z(n2417) );
  NAND U5139 ( .A(n2415), .B(n2414), .Z(n2416) );
  AND U5140 ( .A(n2417), .B(n2416), .Z(n2426) );
  IV U5141 ( .A(n2426), .Z(n2425) );
  XOR U5142 ( .A(n2427), .B(n2425), .Z(n2418) );
  XNOR U5143 ( .A(n2428), .B(n2418), .Z(N46) );
  NAND U5144 ( .A(n2420), .B(n2419), .Z(n2424) );
  NAND U5145 ( .A(n2422), .B(n2421), .Z(n2423) );
  NAND U5146 ( .A(n2424), .B(n2423), .Z(n2578) );
  IV U5147 ( .A(n2578), .Z(n2576) );
  OR U5148 ( .A(n2427), .B(n2425), .Z(n2431) );
  ANDN U5149 ( .B(n2427), .A(n2426), .Z(n2429) );
  OR U5150 ( .A(n2429), .B(n2428), .Z(n2430) );
  AND U5151 ( .A(n2431), .B(n2430), .Z(n2577) );
  NAND U5152 ( .A(n2433), .B(n2432), .Z(n2437) );
  NANDN U5153 ( .A(n2435), .B(n2434), .Z(n2436) );
  AND U5154 ( .A(n2437), .B(n2436), .Z(n2503) );
  NANDN U5155 ( .A(n2439), .B(n2438), .Z(n2443) );
  NANDN U5156 ( .A(n2441), .B(n2440), .Z(n2442) );
  AND U5157 ( .A(n2443), .B(n2442), .Z(n2509) );
  AND U5158 ( .A(x[491]), .B(y[7685]), .Z(n2621) );
  NAND U5159 ( .A(n2621), .B(n2444), .Z(n2447) );
  NANDN U5160 ( .A(n2445), .B(n3319), .Z(n2446) );
  NAND U5161 ( .A(n2447), .B(n2446), .Z(n2565) );
  AND U5162 ( .A(y[7692]), .B(x[487]), .Z(n3034) );
  NAND U5163 ( .A(n3034), .B(n2448), .Z(n2452) );
  NAND U5164 ( .A(n2450), .B(n2449), .Z(n2451) );
  NAND U5165 ( .A(n2452), .B(n2451), .Z(n2564) );
  XOR U5166 ( .A(n2565), .B(n2564), .Z(n2567) );
  AND U5167 ( .A(x[484]), .B(y[7690]), .Z(n2927) );
  AND U5168 ( .A(x[488]), .B(y[7686]), .Z(n2454) );
  NAND U5169 ( .A(x[483]), .B(y[7691]), .Z(n2453) );
  XNOR U5170 ( .A(n2454), .B(n2453), .Z(n2550) );
  XOR U5171 ( .A(n2831), .B(n2550), .Z(n2559) );
  XOR U5172 ( .A(n2927), .B(n2559), .Z(n2561) );
  AND U5173 ( .A(x[489]), .B(y[7685]), .Z(n3109) );
  AND U5174 ( .A(x[482]), .B(y[7692]), .Z(n2456) );
  NAND U5175 ( .A(y[7684]), .B(x[490]), .Z(n2455) );
  XNOR U5176 ( .A(n2456), .B(n2455), .Z(n2535) );
  XOR U5177 ( .A(n3109), .B(n2535), .Z(n2560) );
  XOR U5178 ( .A(n2561), .B(n2560), .Z(n2566) );
  XOR U5179 ( .A(n2567), .B(n2566), .Z(n2507) );
  NAND U5180 ( .A(n2458), .B(n2457), .Z(n2462) );
  NANDN U5181 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U5182 ( .A(n2462), .B(n2461), .Z(n2506) );
  XOR U5183 ( .A(n2509), .B(n2508), .Z(n2501) );
  AND U5184 ( .A(y[7691]), .B(x[489]), .Z(n2463) );
  NAND U5185 ( .A(n2463), .B(n2534), .Z(n2466) );
  NANDN U5186 ( .A(n2464), .B(n3426), .Z(n2465) );
  NAND U5187 ( .A(n2466), .B(n2465), .Z(n2520) );
  AND U5188 ( .A(x[494]), .B(y[7680]), .Z(n2468) );
  NAND U5189 ( .A(y[7694]), .B(x[480]), .Z(n2467) );
  XNOR U5190 ( .A(n2468), .B(n2467), .Z(n2545) );
  AND U5191 ( .A(o[13]), .B(n2469), .Z(n2544) );
  XOR U5192 ( .A(n2545), .B(n2544), .Z(n2519) );
  AND U5193 ( .A(y[7682]), .B(x[492]), .Z(n3099) );
  NAND U5194 ( .A(x[487]), .B(y[7687]), .Z(n2470) );
  XNOR U5195 ( .A(n3099), .B(n2470), .Z(n2526) );
  AND U5196 ( .A(y[7681]), .B(x[493]), .Z(n2533) );
  XOR U5197 ( .A(o[14]), .B(n2533), .Z(n2525) );
  XOR U5198 ( .A(n2526), .B(n2525), .Z(n2518) );
  XOR U5199 ( .A(n2519), .B(n2518), .Z(n2521) );
  XNOR U5200 ( .A(n2520), .B(n2521), .Z(n2571) );
  AND U5201 ( .A(y[7690]), .B(x[485]), .Z(n2608) );
  NANDN U5202 ( .A(n3307), .B(n2608), .Z(n2474) );
  NANDN U5203 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U5204 ( .A(n2474), .B(n2473), .Z(n2514) );
  AND U5205 ( .A(y[7693]), .B(x[493]), .Z(n4022) );
  NAND U5206 ( .A(n4022), .B(n2595), .Z(n2478) );
  NAND U5207 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U5208 ( .A(n2478), .B(n2477), .Z(n2512) );
  AND U5209 ( .A(y[7683]), .B(x[491]), .Z(n2480) );
  NAND U5210 ( .A(x[486]), .B(y[7688]), .Z(n2479) );
  XNOR U5211 ( .A(n2480), .B(n2479), .Z(n2541) );
  AND U5212 ( .A(x[481]), .B(y[7693]), .Z(n2540) );
  XOR U5213 ( .A(n2541), .B(n2540), .Z(n2513) );
  XNOR U5214 ( .A(n2512), .B(n2513), .Z(n2515) );
  XOR U5215 ( .A(n2514), .B(n2515), .Z(n2570) );
  XOR U5216 ( .A(n2571), .B(n2570), .Z(n2573) );
  NAND U5217 ( .A(n2482), .B(n2481), .Z(n2486) );
  NANDN U5218 ( .A(n2484), .B(n2483), .Z(n2485) );
  AND U5219 ( .A(n2486), .B(n2485), .Z(n2572) );
  XNOR U5220 ( .A(n2573), .B(n2572), .Z(n2500) );
  NAND U5221 ( .A(n2488), .B(n2487), .Z(n2492) );
  NAND U5222 ( .A(n2490), .B(n2489), .Z(n2491) );
  NAND U5223 ( .A(n2492), .B(n2491), .Z(n2584) );
  NAND U5224 ( .A(n2494), .B(n2493), .Z(n2498) );
  NAND U5225 ( .A(n2496), .B(n2495), .Z(n2497) );
  NAND U5226 ( .A(n2498), .B(n2497), .Z(n2583) );
  XNOR U5227 ( .A(n2584), .B(n2583), .Z(n2586) );
  XNOR U5228 ( .A(n2577), .B(n2579), .Z(n2499) );
  XOR U5229 ( .A(n2576), .B(n2499), .Z(N47) );
  NANDN U5230 ( .A(n2501), .B(n2500), .Z(n2505) );
  NANDN U5231 ( .A(n2503), .B(n2502), .Z(n2504) );
  AND U5232 ( .A(n2505), .B(n2504), .Z(n2675) );
  NANDN U5233 ( .A(n2507), .B(n2506), .Z(n2511) );
  NAND U5234 ( .A(n2509), .B(n2508), .Z(n2510) );
  NAND U5235 ( .A(n2511), .B(n2510), .Z(n2650) );
  NAND U5236 ( .A(n2513), .B(n2512), .Z(n2517) );
  NANDN U5237 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U5238 ( .A(n2517), .B(n2516), .Z(n2656) );
  NAND U5239 ( .A(n2519), .B(n2518), .Z(n2523) );
  NAND U5240 ( .A(n2521), .B(n2520), .Z(n2522) );
  NAND U5241 ( .A(n2523), .B(n2522), .Z(n2654) );
  AND U5242 ( .A(y[7687]), .B(x[492]), .Z(n3025) );
  NAND U5243 ( .A(n3025), .B(n2524), .Z(n2528) );
  NAND U5244 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U5245 ( .A(n2528), .B(n2527), .Z(n2631) );
  AND U5246 ( .A(y[7684]), .B(x[491]), .Z(n2530) );
  NAND U5247 ( .A(y[7682]), .B(x[493]), .Z(n2529) );
  XNOR U5248 ( .A(n2530), .B(n2529), .Z(n2635) );
  AND U5249 ( .A(x[492]), .B(y[7683]), .Z(n2634) );
  XNOR U5250 ( .A(n2635), .B(n2634), .Z(n2629) );
  AND U5251 ( .A(x[495]), .B(y[7680]), .Z(n2532) );
  NAND U5252 ( .A(y[7695]), .B(x[480]), .Z(n2531) );
  XNOR U5253 ( .A(n2532), .B(n2531), .Z(n2597) );
  AND U5254 ( .A(o[14]), .B(n2533), .Z(n2596) );
  XNOR U5255 ( .A(n2597), .B(n2596), .Z(n2628) );
  XOR U5256 ( .A(n2629), .B(n2628), .Z(n2630) );
  XOR U5257 ( .A(n2631), .B(n2630), .Z(n2663) );
  NAND U5258 ( .A(x[490]), .B(y[7692]), .Z(n3428) );
  NANDN U5259 ( .A(n3428), .B(n2534), .Z(n2537) );
  NAND U5260 ( .A(n3109), .B(n2535), .Z(n2536) );
  NAND U5261 ( .A(n2537), .B(n2536), .Z(n2661) );
  AND U5262 ( .A(y[7688]), .B(x[491]), .Z(n2539) );
  NAND U5263 ( .A(n2539), .B(n2538), .Z(n2543) );
  NAND U5264 ( .A(n2541), .B(n2540), .Z(n2542) );
  NAND U5265 ( .A(n2543), .B(n2542), .Z(n2660) );
  XOR U5266 ( .A(n2661), .B(n2660), .Z(n2662) );
  XOR U5267 ( .A(n2654), .B(n2655), .Z(n2657) );
  XOR U5268 ( .A(n2656), .B(n2657), .Z(n2649) );
  AND U5269 ( .A(y[7694]), .B(x[494]), .Z(n4298) );
  NAND U5270 ( .A(n4298), .B(n2595), .Z(n2547) );
  NAND U5271 ( .A(n2545), .B(n2544), .Z(n2546) );
  NAND U5272 ( .A(n2547), .B(n2546), .Z(n2623) );
  AND U5273 ( .A(y[7691]), .B(x[488]), .Z(n2548) );
  NAND U5274 ( .A(n2549), .B(n2548), .Z(n2552) );
  NAND U5275 ( .A(n2831), .B(n2550), .Z(n2551) );
  NAND U5276 ( .A(n2552), .B(n2551), .Z(n2622) );
  XOR U5277 ( .A(n2623), .B(n2622), .Z(n2625) );
  AND U5278 ( .A(y[7685]), .B(x[490]), .Z(n2554) );
  NAND U5279 ( .A(x[484]), .B(y[7691]), .Z(n2553) );
  XNOR U5280 ( .A(n2554), .B(n2553), .Z(n2603) );
  AND U5281 ( .A(y[7688]), .B(x[487]), .Z(n2602) );
  XNOR U5282 ( .A(n2603), .B(n2602), .Z(n2610) );
  NAND U5283 ( .A(y[7689]), .B(x[486]), .Z(n2744) );
  XNOR U5284 ( .A(n2744), .B(n2608), .Z(n2609) );
  XNOR U5285 ( .A(n2610), .B(n2609), .Z(n2644) );
  AND U5286 ( .A(y[7693]), .B(x[482]), .Z(n2556) );
  NAND U5287 ( .A(x[489]), .B(y[7686]), .Z(n2555) );
  XNOR U5288 ( .A(n2556), .B(n2555), .Z(n2613) );
  AND U5289 ( .A(y[7692]), .B(x[483]), .Z(n2614) );
  XOR U5290 ( .A(n2613), .B(n2614), .Z(n2643) );
  AND U5291 ( .A(y[7694]), .B(x[481]), .Z(n2558) );
  NAND U5292 ( .A(y[7687]), .B(x[488]), .Z(n2557) );
  XNOR U5293 ( .A(n2558), .B(n2557), .Z(n2592) );
  AND U5294 ( .A(y[7681]), .B(x[494]), .Z(n2619) );
  XOR U5295 ( .A(o[15]), .B(n2619), .Z(n2591) );
  XOR U5296 ( .A(n2592), .B(n2591), .Z(n2642) );
  XOR U5297 ( .A(n2643), .B(n2642), .Z(n2645) );
  XOR U5298 ( .A(n2644), .B(n2645), .Z(n2624) );
  XOR U5299 ( .A(n2625), .B(n2624), .Z(n2667) );
  NAND U5300 ( .A(n2927), .B(n2559), .Z(n2563) );
  NAND U5301 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U5302 ( .A(n2563), .B(n2562), .Z(n2666) );
  NAND U5303 ( .A(n2565), .B(n2564), .Z(n2569) );
  NAND U5304 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U5305 ( .A(n2569), .B(n2568), .Z(n2668) );
  XOR U5306 ( .A(n2669), .B(n2668), .Z(n2648) );
  XOR U5307 ( .A(n2650), .B(n2651), .Z(n2672) );
  NAND U5308 ( .A(n2571), .B(n2570), .Z(n2575) );
  NAND U5309 ( .A(n2573), .B(n2572), .Z(n2574) );
  AND U5310 ( .A(n2575), .B(n2574), .Z(n2673) );
  XOR U5311 ( .A(n2672), .B(n2673), .Z(n2674) );
  XOR U5312 ( .A(n2675), .B(n2674), .Z(n2680) );
  NANDN U5313 ( .A(n2576), .B(n2577), .Z(n2582) );
  NOR U5314 ( .A(n2578), .B(n2577), .Z(n2580) );
  OR U5315 ( .A(n2580), .B(n2579), .Z(n2581) );
  AND U5316 ( .A(n2582), .B(n2581), .Z(n2679) );
  NAND U5317 ( .A(n2584), .B(n2583), .Z(n2588) );
  NANDN U5318 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U5319 ( .A(n2588), .B(n2587), .Z(n2678) );
  XOR U5320 ( .A(n2679), .B(n2678), .Z(n2589) );
  XNOR U5321 ( .A(n2680), .B(n2589), .Z(N48) );
  AND U5322 ( .A(x[488]), .B(y[7694]), .Z(n2928) );
  NAND U5323 ( .A(n2928), .B(n2590), .Z(n2594) );
  NAND U5324 ( .A(n2592), .B(n2591), .Z(n2593) );
  AND U5325 ( .A(n2594), .B(n2593), .Z(n2695) );
  AND U5326 ( .A(x[495]), .B(y[7695]), .Z(n4670) );
  NAND U5327 ( .A(n4670), .B(n2595), .Z(n2599) );
  NAND U5328 ( .A(n2597), .B(n2596), .Z(n2598) );
  NAND U5329 ( .A(n2599), .B(n2598), .Z(n2694) );
  AND U5330 ( .A(y[7691]), .B(x[490]), .Z(n2601) );
  NAND U5331 ( .A(n2601), .B(n2600), .Z(n2605) );
  NAND U5332 ( .A(n2603), .B(n2602), .Z(n2604) );
  NAND U5333 ( .A(n2605), .B(n2604), .Z(n2731) );
  AND U5334 ( .A(x[480]), .B(y[7696]), .Z(n2753) );
  AND U5335 ( .A(y[7680]), .B(x[496]), .Z(n2754) );
  XOR U5336 ( .A(n2753), .B(n2754), .Z(n2755) );
  NAND U5337 ( .A(y[7681]), .B(x[495]), .Z(n2741) );
  XNOR U5338 ( .A(o[16]), .B(n2741), .Z(n2756) );
  XOR U5339 ( .A(n2755), .B(n2756), .Z(n2730) );
  NAND U5340 ( .A(x[487]), .B(y[7689]), .Z(n2606) );
  XNOR U5341 ( .A(n2607), .B(n2606), .Z(n2746) );
  AND U5342 ( .A(y[7686]), .B(x[490]), .Z(n2745) );
  XOR U5343 ( .A(n2746), .B(n2745), .Z(n2729) );
  XOR U5344 ( .A(n2730), .B(n2729), .Z(n2732) );
  XOR U5345 ( .A(n2731), .B(n2732), .Z(n2696) );
  XNOR U5346 ( .A(n2697), .B(n2696), .Z(n2726) );
  NANDN U5347 ( .A(n2608), .B(n2744), .Z(n2612) );
  NAND U5348 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U5349 ( .A(n2612), .B(n2611), .Z(n2724) );
  NAND U5350 ( .A(x[489]), .B(y[7693]), .Z(n3410) );
  NANDN U5351 ( .A(n3410), .B(n3024), .Z(n2616) );
  NAND U5352 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U5353 ( .A(n2616), .B(n2615), .Z(n2764) );
  AND U5354 ( .A(y[7695]), .B(x[481]), .Z(n2618) );
  NAND U5355 ( .A(y[7688]), .B(x[488]), .Z(n2617) );
  XNOR U5356 ( .A(n2618), .B(n2617), .Z(n2750) );
  AND U5357 ( .A(o[15]), .B(n2619), .Z(n2749) );
  XOR U5358 ( .A(n2750), .B(n2749), .Z(n2761) );
  NAND U5359 ( .A(y[7682]), .B(x[494]), .Z(n2620) );
  XNOR U5360 ( .A(n2621), .B(n2620), .Z(n2706) );
  NAND U5361 ( .A(x[484]), .B(y[7692]), .Z(n2707) );
  XNOR U5362 ( .A(n2706), .B(n2707), .Z(n2762) );
  XOR U5363 ( .A(n2761), .B(n2762), .Z(n2763) );
  XOR U5364 ( .A(n2764), .B(n2763), .Z(n2723) );
  XOR U5365 ( .A(n2724), .B(n2723), .Z(n2725) );
  XOR U5366 ( .A(n2726), .B(n2725), .Z(n2688) );
  NAND U5367 ( .A(n2623), .B(n2622), .Z(n2627) );
  NAND U5368 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U5369 ( .A(n2627), .B(n2626), .Z(n2689) );
  XOR U5370 ( .A(n2688), .B(n2689), .Z(n2691) );
  NAND U5371 ( .A(n2629), .B(n2628), .Z(n2633) );
  NAND U5372 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U5373 ( .A(n2633), .B(n2632), .Z(n2720) );
  AND U5374 ( .A(x[493]), .B(y[7684]), .Z(n2716) );
  NAND U5375 ( .A(n3268), .B(n2716), .Z(n2637) );
  NAND U5376 ( .A(n2635), .B(n2634), .Z(n2636) );
  NAND U5377 ( .A(n2637), .B(n2636), .Z(n2703) );
  AND U5378 ( .A(x[482]), .B(y[7694]), .Z(n2639) );
  NAND U5379 ( .A(y[7687]), .B(x[489]), .Z(n2638) );
  XNOR U5380 ( .A(n2639), .B(n2638), .Z(n2710) );
  NAND U5381 ( .A(x[483]), .B(y[7693]), .Z(n2711) );
  XNOR U5382 ( .A(n2710), .B(n2711), .Z(n2701) );
  AND U5383 ( .A(x[492]), .B(y[7684]), .Z(n3398) );
  AND U5384 ( .A(y[7683]), .B(x[493]), .Z(n2641) );
  NAND U5385 ( .A(x[485]), .B(y[7691]), .Z(n2640) );
  XNOR U5386 ( .A(n2641), .B(n2640), .Z(n2736) );
  XOR U5387 ( .A(n3398), .B(n2736), .Z(n2700) );
  XOR U5388 ( .A(n2701), .B(n2700), .Z(n2702) );
  XNOR U5389 ( .A(n2703), .B(n2702), .Z(n2717) );
  NAND U5390 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U5391 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U5392 ( .A(n2647), .B(n2646), .Z(n2718) );
  XOR U5393 ( .A(n2717), .B(n2718), .Z(n2719) );
  XOR U5394 ( .A(n2720), .B(n2719), .Z(n2690) );
  XOR U5395 ( .A(n2691), .B(n2690), .Z(n2768) );
  NANDN U5396 ( .A(n2649), .B(n2648), .Z(n2653) );
  NANDN U5397 ( .A(n2651), .B(n2650), .Z(n2652) );
  AND U5398 ( .A(n2653), .B(n2652), .Z(n2767) );
  NAND U5399 ( .A(n2655), .B(n2654), .Z(n2659) );
  NAND U5400 ( .A(n2657), .B(n2656), .Z(n2658) );
  NAND U5401 ( .A(n2659), .B(n2658), .Z(n2684) );
  NAND U5402 ( .A(n2661), .B(n2660), .Z(n2665) );
  NANDN U5403 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U5404 ( .A(n2665), .B(n2664), .Z(n2682) );
  NANDN U5405 ( .A(n2667), .B(n2666), .Z(n2671) );
  NAND U5406 ( .A(n2669), .B(n2668), .Z(n2670) );
  AND U5407 ( .A(n2671), .B(n2670), .Z(n2683) );
  XOR U5408 ( .A(n2682), .B(n2683), .Z(n2685) );
  XOR U5409 ( .A(n2684), .B(n2685), .Z(n2769) );
  XNOR U5410 ( .A(n2770), .B(n2769), .Z(n2775) );
  NAND U5411 ( .A(n2673), .B(n2672), .Z(n2677) );
  NANDN U5412 ( .A(n2675), .B(n2674), .Z(n2676) );
  NAND U5413 ( .A(n2677), .B(n2676), .Z(n2773) );
  XOR U5414 ( .A(n2773), .B(n2774), .Z(n2681) );
  XNOR U5415 ( .A(n2775), .B(n2681), .Z(N49) );
  NAND U5416 ( .A(n2683), .B(n2682), .Z(n2687) );
  NAND U5417 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U5418 ( .A(n2687), .B(n2686), .Z(n2870) );
  NAND U5419 ( .A(n2689), .B(n2688), .Z(n2693) );
  NAND U5420 ( .A(n2691), .B(n2690), .Z(n2692) );
  NAND U5421 ( .A(n2693), .B(n2692), .Z(n2780) );
  NANDN U5422 ( .A(n2695), .B(n2694), .Z(n2699) );
  NAND U5423 ( .A(n2697), .B(n2696), .Z(n2698) );
  NAND U5424 ( .A(n2699), .B(n2698), .Z(n2856) );
  NAND U5425 ( .A(n2701), .B(n2700), .Z(n2705) );
  NAND U5426 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U5427 ( .A(n2705), .B(n2704), .Z(n2854) );
  NAND U5428 ( .A(x[494]), .B(y[7685]), .Z(n3060) );
  NANDN U5429 ( .A(n3060), .B(n3268), .Z(n2709) );
  NANDN U5430 ( .A(n2707), .B(n2706), .Z(n2708) );
  AND U5431 ( .A(n2709), .B(n2708), .Z(n2848) );
  AND U5432 ( .A(x[489]), .B(y[7694]), .Z(n3665) );
  NAND U5433 ( .A(n2838), .B(n3665), .Z(n2713) );
  NANDN U5434 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U5435 ( .A(n2713), .B(n2712), .Z(n2847) );
  XNOR U5436 ( .A(n2848), .B(n2847), .Z(n2849) );
  AND U5437 ( .A(x[487]), .B(y[7690]), .Z(n2844) );
  AND U5438 ( .A(x[485]), .B(y[7692]), .Z(n2891) );
  NAND U5439 ( .A(y[7689]), .B(x[488]), .Z(n2714) );
  XNOR U5440 ( .A(n2891), .B(n2714), .Z(n2832) );
  XOR U5441 ( .A(n2844), .B(n2843), .Z(n2845) );
  NAND U5442 ( .A(y[7693]), .B(x[484]), .Z(n2715) );
  XNOR U5443 ( .A(n2716), .B(n2715), .Z(n2794) );
  NAND U5444 ( .A(y[7686]), .B(x[491]), .Z(n2795) );
  XOR U5445 ( .A(n2794), .B(n2795), .Z(n2846) );
  XOR U5446 ( .A(n2845), .B(n2846), .Z(n2850) );
  XNOR U5447 ( .A(n2849), .B(n2850), .Z(n2853) );
  XOR U5448 ( .A(n2854), .B(n2853), .Z(n2855) );
  XNOR U5449 ( .A(n2856), .B(n2855), .Z(n2778) );
  NAND U5450 ( .A(n2718), .B(n2717), .Z(n2722) );
  NAND U5451 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U5452 ( .A(n2722), .B(n2721), .Z(n2777) );
  XOR U5453 ( .A(n2778), .B(n2777), .Z(n2779) );
  XOR U5454 ( .A(n2780), .B(n2779), .Z(n2869) );
  NAND U5455 ( .A(n2724), .B(n2723), .Z(n2728) );
  NAND U5456 ( .A(n2726), .B(n2725), .Z(n2727) );
  AND U5457 ( .A(n2728), .B(n2727), .Z(n2786) );
  NAND U5458 ( .A(n2730), .B(n2729), .Z(n2734) );
  NAND U5459 ( .A(n2732), .B(n2731), .Z(n2733) );
  AND U5460 ( .A(n2734), .B(n2733), .Z(n2862) );
  AND U5461 ( .A(y[7691]), .B(x[493]), .Z(n3684) );
  NAND U5462 ( .A(n3684), .B(n2735), .Z(n2738) );
  NAND U5463 ( .A(n2736), .B(n3398), .Z(n2737) );
  NAND U5464 ( .A(n2738), .B(n2737), .Z(n2816) );
  AND U5465 ( .A(y[7696]), .B(x[481]), .Z(n2740) );
  NAND U5466 ( .A(y[7688]), .B(x[489]), .Z(n2739) );
  XNOR U5467 ( .A(n2740), .B(n2739), .Z(n2837) );
  ANDN U5468 ( .B(o[16]), .A(n2741), .Z(n2836) );
  XOR U5469 ( .A(n2837), .B(n2836), .Z(n2814) );
  AND U5470 ( .A(y[7682]), .B(x[495]), .Z(n2743) );
  NAND U5471 ( .A(y[7685]), .B(x[492]), .Z(n2742) );
  XNOR U5472 ( .A(n2743), .B(n2742), .Z(n2790) );
  AND U5473 ( .A(x[494]), .B(y[7683]), .Z(n2789) );
  XOR U5474 ( .A(n2790), .B(n2789), .Z(n2813) );
  XOR U5475 ( .A(n2814), .B(n2813), .Z(n2815) );
  XOR U5476 ( .A(n2816), .B(n2815), .Z(n2860) );
  NANDN U5477 ( .A(n2744), .B(n2844), .Z(n2748) );
  NAND U5478 ( .A(n2746), .B(n2745), .Z(n2747) );
  NAND U5479 ( .A(n2748), .B(n2747), .Z(n2826) );
  NAND U5480 ( .A(x[488]), .B(y[7695]), .Z(n3493) );
  AND U5481 ( .A(x[481]), .B(y[7688]), .Z(n2906) );
  NANDN U5482 ( .A(n3493), .B(n2906), .Z(n2752) );
  NAND U5483 ( .A(n2750), .B(n2749), .Z(n2751) );
  NAND U5484 ( .A(n2752), .B(n2751), .Z(n2825) );
  XOR U5485 ( .A(n2826), .B(n2825), .Z(n2828) );
  NAND U5486 ( .A(n2754), .B(n2753), .Z(n2758) );
  NAND U5487 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U5488 ( .A(n2758), .B(n2757), .Z(n2822) );
  AND U5489 ( .A(x[480]), .B(y[7697]), .Z(n2804) );
  AND U5490 ( .A(x[497]), .B(y[7680]), .Z(n2803) );
  XOR U5491 ( .A(n2804), .B(n2803), .Z(n2806) );
  AND U5492 ( .A(y[7681]), .B(x[496]), .Z(n2798) );
  XOR U5493 ( .A(n2798), .B(o[17]), .Z(n2805) );
  XOR U5494 ( .A(n2806), .B(n2805), .Z(n2820) );
  AND U5495 ( .A(y[7695]), .B(x[482]), .Z(n2760) );
  NAND U5496 ( .A(y[7687]), .B(x[490]), .Z(n2759) );
  XNOR U5497 ( .A(n2760), .B(n2759), .Z(n2840) );
  AND U5498 ( .A(y[7694]), .B(x[483]), .Z(n2839) );
  XOR U5499 ( .A(n2840), .B(n2839), .Z(n2819) );
  XOR U5500 ( .A(n2820), .B(n2819), .Z(n2821) );
  XOR U5501 ( .A(n2822), .B(n2821), .Z(n2827) );
  XOR U5502 ( .A(n2828), .B(n2827), .Z(n2859) );
  XOR U5503 ( .A(n2860), .B(n2859), .Z(n2861) );
  NAND U5504 ( .A(n2762), .B(n2761), .Z(n2766) );
  NANDN U5505 ( .A(n2764), .B(n2763), .Z(n2765) );
  AND U5506 ( .A(n2766), .B(n2765), .Z(n2784) );
  XOR U5507 ( .A(n2783), .B(n2784), .Z(n2785) );
  XOR U5508 ( .A(n2786), .B(n2785), .Z(n2868) );
  XOR U5509 ( .A(n2870), .B(n2871), .Z(n2867) );
  NANDN U5510 ( .A(n2768), .B(n2767), .Z(n2772) );
  NAND U5511 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U5512 ( .A(n2772), .B(n2771), .Z(n2866) );
  XNOR U5513 ( .A(n2866), .B(n2865), .Z(n2776) );
  XNOR U5514 ( .A(n2867), .B(n2776), .Z(N50) );
  NAND U5515 ( .A(n2778), .B(n2777), .Z(n2782) );
  NAND U5516 ( .A(n2780), .B(n2779), .Z(n2781) );
  AND U5517 ( .A(n2782), .B(n2781), .Z(n2973) );
  NAND U5518 ( .A(n2784), .B(n2783), .Z(n2788) );
  NANDN U5519 ( .A(n2786), .B(n2785), .Z(n2787) );
  AND U5520 ( .A(n2788), .B(n2787), .Z(n2971) );
  AND U5521 ( .A(x[495]), .B(y[7685]), .Z(n3032) );
  NAND U5522 ( .A(n3099), .B(n3032), .Z(n2792) );
  NAND U5523 ( .A(n2790), .B(n2789), .Z(n2791) );
  NAND U5524 ( .A(n2792), .B(n2791), .Z(n2952) );
  NAND U5525 ( .A(n4022), .B(n2793), .Z(n2797) );
  NANDN U5526 ( .A(n2795), .B(n2794), .Z(n2796) );
  NAND U5527 ( .A(n2797), .B(n2796), .Z(n2941) );
  AND U5528 ( .A(n2798), .B(o[17]), .Z(n2908) );
  AND U5529 ( .A(y[7697]), .B(x[481]), .Z(n2800) );
  XOR U5530 ( .A(n2800), .B(n2799), .Z(n2907) );
  XOR U5531 ( .A(n2908), .B(n2907), .Z(n2939) );
  AND U5532 ( .A(y[7683]), .B(x[495]), .Z(n2802) );
  NAND U5533 ( .A(y[7689]), .B(x[489]), .Z(n2801) );
  XNOR U5534 ( .A(n2802), .B(n2801), .Z(n2899) );
  AND U5535 ( .A(x[494]), .B(y[7684]), .Z(n2898) );
  XOR U5536 ( .A(n2899), .B(n2898), .Z(n2938) );
  XOR U5537 ( .A(n2939), .B(n2938), .Z(n2942) );
  XOR U5538 ( .A(n2941), .B(n2942), .Z(n2953) );
  XOR U5539 ( .A(n2952), .B(n2953), .Z(n2955) );
  NAND U5540 ( .A(n2804), .B(n2803), .Z(n2808) );
  NAND U5541 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U5542 ( .A(n2808), .B(n2807), .Z(n2964) );
  AND U5543 ( .A(y[7682]), .B(x[496]), .Z(n2810) );
  NAND U5544 ( .A(x[491]), .B(y[7687]), .Z(n2809) );
  XNOR U5545 ( .A(n2810), .B(n2809), .Z(n2897) );
  AND U5546 ( .A(x[482]), .B(y[7696]), .Z(n2896) );
  XOR U5547 ( .A(n2897), .B(n2896), .Z(n2965) );
  XOR U5548 ( .A(n2964), .B(n2965), .Z(n2967) );
  AND U5549 ( .A(y[7693]), .B(x[485]), .Z(n3041) );
  NAND U5550 ( .A(x[486]), .B(y[7692]), .Z(n2811) );
  XNOR U5551 ( .A(n3041), .B(n2811), .Z(n2893) );
  NAND U5552 ( .A(y[7694]), .B(x[484]), .Z(n2812) );
  XNOR U5553 ( .A(n3670), .B(n2812), .Z(n2930) );
  AND U5554 ( .A(y[7691]), .B(x[487]), .Z(n2929) );
  XOR U5555 ( .A(n2930), .B(n2929), .Z(n2892) );
  XOR U5556 ( .A(n2893), .B(n2892), .Z(n2966) );
  XOR U5557 ( .A(n2967), .B(n2966), .Z(n2954) );
  XOR U5558 ( .A(n2955), .B(n2954), .Z(n2882) );
  NAND U5559 ( .A(n2814), .B(n2813), .Z(n2818) );
  NAND U5560 ( .A(n2816), .B(n2815), .Z(n2817) );
  AND U5561 ( .A(n2818), .B(n2817), .Z(n2947) );
  NAND U5562 ( .A(n2820), .B(n2819), .Z(n2824) );
  NAND U5563 ( .A(n2822), .B(n2821), .Z(n2823) );
  AND U5564 ( .A(n2824), .B(n2823), .Z(n2946) );
  XOR U5565 ( .A(n2947), .B(n2946), .Z(n2949) );
  NAND U5566 ( .A(n2826), .B(n2825), .Z(n2830) );
  NAND U5567 ( .A(n2828), .B(n2827), .Z(n2829) );
  AND U5568 ( .A(n2830), .B(n2829), .Z(n2948) );
  XOR U5569 ( .A(n2949), .B(n2948), .Z(n2881) );
  AND U5570 ( .A(x[488]), .B(y[7692]), .Z(n3145) );
  NAND U5571 ( .A(n3145), .B(n2831), .Z(n2835) );
  NANDN U5572 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U5573 ( .A(n2835), .B(n2834), .Z(n2959) );
  AND U5574 ( .A(x[489]), .B(y[7696]), .Z(n3778) );
  XOR U5575 ( .A(n2959), .B(n2958), .Z(n2960) );
  AND U5576 ( .A(x[490]), .B(y[7695]), .Z(n3693) );
  IV U5577 ( .A(n3693), .Z(n3777) );
  AND U5578 ( .A(x[480]), .B(y[7698]), .Z(n2912) );
  AND U5579 ( .A(y[7680]), .B(x[498]), .Z(n2911) );
  XOR U5580 ( .A(n2912), .B(n2911), .Z(n2914) );
  AND U5581 ( .A(x[497]), .B(y[7681]), .Z(n2931) );
  XOR U5582 ( .A(n2931), .B(o[18]), .Z(n2913) );
  XOR U5583 ( .A(n2914), .B(n2913), .Z(n2935) );
  AND U5584 ( .A(y[7685]), .B(x[493]), .Z(n2842) );
  NAND U5585 ( .A(y[7695]), .B(x[483]), .Z(n2841) );
  XNOR U5586 ( .A(n2842), .B(n2841), .Z(n2920) );
  AND U5587 ( .A(y[7686]), .B(x[492]), .Z(n2919) );
  XOR U5588 ( .A(n2920), .B(n2919), .Z(n2934) );
  XOR U5589 ( .A(n2935), .B(n2934), .Z(n2936) );
  XNOR U5590 ( .A(n2937), .B(n2936), .Z(n2961) );
  XNOR U5591 ( .A(n2960), .B(n2961), .Z(n2888) );
  XNOR U5592 ( .A(n2888), .B(n2887), .Z(n2890) );
  NANDN U5593 ( .A(n2848), .B(n2847), .Z(n2852) );
  NANDN U5594 ( .A(n2850), .B(n2849), .Z(n2851) );
  AND U5595 ( .A(n2852), .B(n2851), .Z(n2889) );
  XOR U5596 ( .A(n2890), .B(n2889), .Z(n2883) );
  XOR U5597 ( .A(n2884), .B(n2883), .Z(n2878) );
  NAND U5598 ( .A(n2854), .B(n2853), .Z(n2858) );
  NAND U5599 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U5600 ( .A(n2858), .B(n2857), .Z(n2876) );
  NAND U5601 ( .A(n2860), .B(n2859), .Z(n2864) );
  NANDN U5602 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U5603 ( .A(n2864), .B(n2863), .Z(n2875) );
  XOR U5604 ( .A(n2971), .B(n2970), .Z(n2972) );
  XOR U5605 ( .A(n2973), .B(n2972), .Z(n2978) );
  NANDN U5606 ( .A(n2869), .B(n2868), .Z(n2873) );
  NAND U5607 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U5608 ( .A(n2873), .B(n2872), .Z(n2976) );
  XOR U5609 ( .A(n2977), .B(n2976), .Z(n2874) );
  XNOR U5610 ( .A(n2978), .B(n2874), .Z(N51) );
  NANDN U5611 ( .A(n2876), .B(n2875), .Z(n2880) );
  NANDN U5612 ( .A(n2878), .B(n2877), .Z(n2879) );
  AND U5613 ( .A(n2880), .B(n2879), .Z(n2983) );
  NANDN U5614 ( .A(n2882), .B(n2881), .Z(n2886) );
  NAND U5615 ( .A(n2884), .B(n2883), .Z(n2885) );
  AND U5616 ( .A(n2886), .B(n2885), .Z(n2981) );
  AND U5617 ( .A(y[7693]), .B(x[486]), .Z(n2933) );
  NAND U5618 ( .A(n2933), .B(n2891), .Z(n2895) );
  NAND U5619 ( .A(n2893), .B(n2892), .Z(n2894) );
  NAND U5620 ( .A(n2895), .B(n2894), .Z(n2995) );
  AND U5621 ( .A(x[495]), .B(y[7689]), .Z(n3698) );
  NAND U5622 ( .A(n3698), .B(n3019), .Z(n2901) );
  NAND U5623 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U5624 ( .A(n2901), .B(n2900), .Z(n3009) );
  AND U5625 ( .A(x[481]), .B(y[7698]), .Z(n2903) );
  NAND U5626 ( .A(x[488]), .B(y[7691]), .Z(n2902) );
  XNOR U5627 ( .A(n2903), .B(n2902), .Z(n3059) );
  AND U5628 ( .A(x[482]), .B(y[7697]), .Z(n2905) );
  NAND U5629 ( .A(x[493]), .B(y[7686]), .Z(n2904) );
  XNOR U5630 ( .A(n2905), .B(n2904), .Z(n3026) );
  XOR U5631 ( .A(n3026), .B(n3025), .Z(n3007) );
  XOR U5632 ( .A(n3008), .B(n3007), .Z(n3010) );
  XOR U5633 ( .A(n3009), .B(n3010), .Z(n2994) );
  XOR U5634 ( .A(n2993), .B(n2994), .Z(n2996) );
  XOR U5635 ( .A(n2995), .B(n2996), .Z(n2990) );
  AND U5636 ( .A(x[490]), .B(y[7697]), .Z(n4174) );
  IV U5637 ( .A(n4174), .Z(n3975) );
  NANDN U5638 ( .A(n3975), .B(n2906), .Z(n2910) );
  NAND U5639 ( .A(n2908), .B(n2907), .Z(n2909) );
  NAND U5640 ( .A(n2910), .B(n2909), .Z(n3070) );
  NAND U5641 ( .A(n2912), .B(n2911), .Z(n2916) );
  NAND U5642 ( .A(n2914), .B(n2913), .Z(n2915) );
  NAND U5643 ( .A(n2916), .B(n2915), .Z(n3068) );
  AND U5644 ( .A(y[7683]), .B(x[496]), .Z(n3636) );
  NAND U5645 ( .A(y[7690]), .B(x[489]), .Z(n2917) );
  XNOR U5646 ( .A(n3636), .B(n2917), .Z(n3020) );
  NAND U5647 ( .A(x[495]), .B(y[7684]), .Z(n3021) );
  XOR U5648 ( .A(n3068), .B(n3069), .Z(n3071) );
  XOR U5649 ( .A(n3070), .B(n3071), .Z(n3000) );
  AND U5650 ( .A(x[493]), .B(y[7695]), .Z(n4327) );
  NANDN U5651 ( .A(n2918), .B(n4327), .Z(n2922) );
  NAND U5652 ( .A(n2920), .B(n2919), .Z(n2921) );
  NAND U5653 ( .A(n2922), .B(n2921), .Z(n3076) );
  AND U5654 ( .A(y[7689]), .B(x[490]), .Z(n2924) );
  NAND U5655 ( .A(y[7682]), .B(x[497]), .Z(n2923) );
  XNOR U5656 ( .A(n2924), .B(n2923), .Z(n3065) );
  AND U5657 ( .A(y[7681]), .B(x[498]), .Z(n3040) );
  XOR U5658 ( .A(o[19]), .B(n3040), .Z(n3064) );
  XOR U5659 ( .A(n3065), .B(n3064), .Z(n3075) );
  AND U5660 ( .A(y[7696]), .B(x[483]), .Z(n2926) );
  NAND U5661 ( .A(x[491]), .B(y[7688]), .Z(n2925) );
  XNOR U5662 ( .A(n2926), .B(n2925), .Z(n3035) );
  XOR U5663 ( .A(n3035), .B(n3034), .Z(n3074) );
  XOR U5664 ( .A(n3075), .B(n3074), .Z(n3077) );
  XOR U5665 ( .A(n3076), .B(n3077), .Z(n2998) );
  AND U5666 ( .A(x[480]), .B(y[7699]), .Z(n3045) );
  NAND U5667 ( .A(y[7680]), .B(x[499]), .Z(n3046) );
  NAND U5668 ( .A(n2931), .B(o[18]), .Z(n3048) );
  AND U5669 ( .A(x[484]), .B(y[7695]), .Z(n3159) );
  NAND U5670 ( .A(x[485]), .B(y[7694]), .Z(n2932) );
  XOR U5671 ( .A(n2933), .B(n2932), .Z(n3042) );
  XOR U5672 ( .A(n3014), .B(n3013), .Z(n3016) );
  XNOR U5673 ( .A(n3015), .B(n3016), .Z(n2997) );
  IV U5674 ( .A(n2938), .Z(n2940) );
  NANDN U5675 ( .A(n2940), .B(n2939), .Z(n2945) );
  IV U5676 ( .A(n2941), .Z(n2943) );
  NANDN U5677 ( .A(n2943), .B(n2942), .Z(n2944) );
  NAND U5678 ( .A(n2945), .B(n2944), .Z(n3004) );
  XNOR U5679 ( .A(n3003), .B(n3004), .Z(n3006) );
  XNOR U5680 ( .A(n3005), .B(n3006), .Z(n2989) );
  XNOR U5681 ( .A(n2990), .B(n2989), .Z(n2992) );
  XNOR U5682 ( .A(n2991), .B(n2992), .Z(n3089) );
  NAND U5683 ( .A(n2947), .B(n2946), .Z(n2951) );
  NAND U5684 ( .A(n2949), .B(n2948), .Z(n2950) );
  AND U5685 ( .A(n2951), .B(n2950), .Z(n3086) );
  NAND U5686 ( .A(n2953), .B(n2952), .Z(n2957) );
  NAND U5687 ( .A(n2955), .B(n2954), .Z(n2956) );
  NAND U5688 ( .A(n2957), .B(n2956), .Z(n3082) );
  NAND U5689 ( .A(n2959), .B(n2958), .Z(n2963) );
  NANDN U5690 ( .A(n2961), .B(n2960), .Z(n2962) );
  NAND U5691 ( .A(n2963), .B(n2962), .Z(n3081) );
  NAND U5692 ( .A(n2965), .B(n2964), .Z(n2969) );
  NAND U5693 ( .A(n2967), .B(n2966), .Z(n2968) );
  NAND U5694 ( .A(n2969), .B(n2968), .Z(n3080) );
  XOR U5695 ( .A(n3081), .B(n3080), .Z(n3083) );
  XNOR U5696 ( .A(n3082), .B(n3083), .Z(n3087) );
  XNOR U5697 ( .A(n3086), .B(n3087), .Z(n3088) );
  XOR U5698 ( .A(n3089), .B(n3088), .Z(n2980) );
  XOR U5699 ( .A(n2981), .B(n2980), .Z(n2982) );
  XOR U5700 ( .A(n2983), .B(n2982), .Z(n2988) );
  NAND U5701 ( .A(n2971), .B(n2970), .Z(n2975) );
  NAND U5702 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U5703 ( .A(n2975), .B(n2974), .Z(n2987) );
  XOR U5704 ( .A(n2987), .B(n2986), .Z(n2979) );
  XNOR U5705 ( .A(n2988), .B(n2979), .Z(N52) );
  NAND U5706 ( .A(n2981), .B(n2980), .Z(n2985) );
  NANDN U5707 ( .A(n2983), .B(n2982), .Z(n2984) );
  NAND U5708 ( .A(n2985), .B(n2984), .Z(n3212) );
  IV U5709 ( .A(n3212), .Z(n3211) );
  NANDN U5710 ( .A(n2998), .B(n2997), .Z(n3002) );
  NANDN U5711 ( .A(n3000), .B(n2999), .Z(n3001) );
  NAND U5712 ( .A(n3002), .B(n3001), .Z(n3202) );
  XNOR U5713 ( .A(n3202), .B(n3201), .Z(n3204) );
  XOR U5714 ( .A(n3203), .B(n3204), .Z(n3195) );
  NAND U5715 ( .A(n3008), .B(n3007), .Z(n3012) );
  NAND U5716 ( .A(n3010), .B(n3009), .Z(n3011) );
  NAND U5717 ( .A(n3012), .B(n3011), .Z(n3094) );
  NAND U5718 ( .A(n3014), .B(n3013), .Z(n3018) );
  NAND U5719 ( .A(n3016), .B(n3015), .Z(n3017) );
  NAND U5720 ( .A(n3018), .B(n3017), .Z(n3093) );
  XOR U5721 ( .A(n3094), .B(n3093), .Z(n3096) );
  AND U5722 ( .A(x[496]), .B(y[7690]), .Z(n3933) );
  NAND U5723 ( .A(n3933), .B(n3019), .Z(n3023) );
  NANDN U5724 ( .A(n3021), .B(n3020), .Z(n3022) );
  AND U5725 ( .A(n3023), .B(n3022), .Z(n3134) );
  AND U5726 ( .A(y[7697]), .B(x[493]), .Z(n4429) );
  NAND U5727 ( .A(n4429), .B(n3024), .Z(n3028) );
  NAND U5728 ( .A(n3026), .B(n3025), .Z(n3027) );
  AND U5729 ( .A(n3028), .B(n3027), .Z(n3179) );
  AND U5730 ( .A(y[7684]), .B(x[496]), .Z(n3030) );
  NAND U5731 ( .A(y[7690]), .B(x[490]), .Z(n3029) );
  XNOR U5732 ( .A(n3030), .B(n3029), .Z(n3140) );
  NAND U5733 ( .A(y[7698]), .B(x[482]), .Z(n3141) );
  NAND U5734 ( .A(x[489]), .B(y[7691]), .Z(n3031) );
  XNOR U5735 ( .A(n3032), .B(n3031), .Z(n3110) );
  AND U5736 ( .A(y[7686]), .B(x[494]), .Z(n3111) );
  XOR U5737 ( .A(n3110), .B(n3111), .Z(n3176) );
  XOR U5738 ( .A(n3177), .B(n3176), .Z(n3178) );
  NAND U5739 ( .A(x[491]), .B(y[7696]), .Z(n4175) );
  NANDN U5740 ( .A(n4175), .B(n3033), .Z(n3037) );
  NAND U5741 ( .A(n3035), .B(n3034), .Z(n3036) );
  AND U5742 ( .A(n3037), .B(n3036), .Z(n3185) );
  AND U5743 ( .A(x[491]), .B(y[7689]), .Z(n3039) );
  NAND U5744 ( .A(x[481]), .B(y[7699]), .Z(n3038) );
  XNOR U5745 ( .A(n3039), .B(n3038), .Z(n3106) );
  AND U5746 ( .A(y[7681]), .B(x[499]), .Z(n3114) );
  XOR U5747 ( .A(o[20]), .B(n3114), .Z(n3105) );
  XOR U5748 ( .A(n3106), .B(n3105), .Z(n3183) );
  AND U5749 ( .A(x[480]), .B(y[7700]), .Z(n3164) );
  AND U5750 ( .A(y[7680]), .B(x[500]), .Z(n3165) );
  XOR U5751 ( .A(n3164), .B(n3165), .Z(n3167) );
  AND U5752 ( .A(o[19]), .B(n3040), .Z(n3166) );
  XOR U5753 ( .A(n3167), .B(n3166), .Z(n3182) );
  XOR U5754 ( .A(n3183), .B(n3182), .Z(n3184) );
  XOR U5755 ( .A(n3136), .B(n3135), .Z(n3095) );
  XOR U5756 ( .A(n3096), .B(n3095), .Z(n3191) );
  AND U5757 ( .A(y[7694]), .B(x[486]), .Z(n3116) );
  IV U5758 ( .A(n3116), .Z(n3057) );
  NANDN U5759 ( .A(n3057), .B(n3041), .Z(n3044) );
  NANDN U5760 ( .A(n3042), .B(n3159), .Z(n3043) );
  AND U5761 ( .A(n3044), .B(n3043), .Z(n3124) );
  NANDN U5762 ( .A(n3046), .B(n3045), .Z(n3050) );
  NANDN U5763 ( .A(n3048), .B(n3047), .Z(n3049) );
  AND U5764 ( .A(n3050), .B(n3049), .Z(n3122) );
  AND U5765 ( .A(y[7682]), .B(x[498]), .Z(n3052) );
  NAND U5766 ( .A(y[7688]), .B(x[492]), .Z(n3051) );
  XNOR U5767 ( .A(n3052), .B(n3051), .Z(n3100) );
  AND U5768 ( .A(x[497]), .B(y[7683]), .Z(n3101) );
  XOR U5769 ( .A(n3100), .B(n3101), .Z(n3121) );
  AND U5770 ( .A(x[483]), .B(y[7697]), .Z(n3054) );
  NAND U5771 ( .A(x[493]), .B(y[7687]), .Z(n3053) );
  XNOR U5772 ( .A(n3054), .B(n3053), .Z(n3146) );
  XOR U5773 ( .A(n3146), .B(n3145), .Z(n3118) );
  AND U5774 ( .A(x[485]), .B(y[7695]), .Z(n3056) );
  NAND U5775 ( .A(y[7696]), .B(x[484]), .Z(n3055) );
  XNOR U5776 ( .A(n3056), .B(n3055), .Z(n3161) );
  AND U5777 ( .A(y[7693]), .B(x[487]), .Z(n3160) );
  XNOR U5778 ( .A(n3161), .B(n3160), .Z(n3115) );
  XOR U5779 ( .A(n3057), .B(n3115), .Z(n3117) );
  AND U5780 ( .A(x[488]), .B(y[7698]), .Z(n4278) );
  AND U5781 ( .A(y[7691]), .B(x[481]), .Z(n3058) );
  NAND U5782 ( .A(n4278), .B(n3058), .Z(n3062) );
  NANDN U5783 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U5784 ( .A(n3062), .B(n3061), .Z(n3171) );
  NAND U5785 ( .A(x[497]), .B(y[7689]), .Z(n3942) );
  NANDN U5786 ( .A(n3942), .B(n3063), .Z(n3067) );
  NAND U5787 ( .A(n3065), .B(n3064), .Z(n3066) );
  NAND U5788 ( .A(n3067), .B(n3066), .Z(n3170) );
  XNOR U5789 ( .A(n3172), .B(n3173), .Z(n3127) );
  NAND U5790 ( .A(n3069), .B(n3068), .Z(n3073) );
  NAND U5791 ( .A(n3071), .B(n3070), .Z(n3072) );
  AND U5792 ( .A(n3073), .B(n3072), .Z(n3129) );
  XOR U5793 ( .A(n3130), .B(n3129), .Z(n3189) );
  NAND U5794 ( .A(n3075), .B(n3074), .Z(n3079) );
  NAND U5795 ( .A(n3077), .B(n3076), .Z(n3078) );
  AND U5796 ( .A(n3079), .B(n3078), .Z(n3188) );
  XOR U5797 ( .A(n3189), .B(n3188), .Z(n3190) );
  XOR U5798 ( .A(n3195), .B(n3196), .Z(n3198) );
  XOR U5799 ( .A(n3197), .B(n3198), .Z(n3207) );
  NAND U5800 ( .A(n3081), .B(n3080), .Z(n3085) );
  NAND U5801 ( .A(n3083), .B(n3082), .Z(n3084) );
  AND U5802 ( .A(n3085), .B(n3084), .Z(n3206) );
  NANDN U5803 ( .A(n3087), .B(n3086), .Z(n3091) );
  NAND U5804 ( .A(n3089), .B(n3088), .Z(n3090) );
  AND U5805 ( .A(n3091), .B(n3090), .Z(n3205) );
  XOR U5806 ( .A(n3206), .B(n3205), .Z(n3208) );
  XOR U5807 ( .A(n3207), .B(n3208), .Z(n3214) );
  XNOR U5808 ( .A(n3213), .B(n3214), .Z(n3092) );
  XOR U5809 ( .A(n3211), .B(n3092), .Z(N53) );
  NAND U5810 ( .A(n3094), .B(n3093), .Z(n3098) );
  NAND U5811 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U5812 ( .A(n3098), .B(n3097), .Z(n3234) );
  AND U5813 ( .A(y[7688]), .B(x[498]), .Z(n3940) );
  NAND U5814 ( .A(n3940), .B(n3099), .Z(n3103) );
  NAND U5815 ( .A(n3101), .B(n3100), .Z(n3102) );
  NAND U5816 ( .A(n3103), .B(n3102), .Z(n3239) );
  AND U5817 ( .A(y[7699]), .B(x[491]), .Z(n4619) );
  NAND U5818 ( .A(n4619), .B(n3104), .Z(n3108) );
  NAND U5819 ( .A(n3106), .B(n3105), .Z(n3107) );
  NAND U5820 ( .A(n3108), .B(n3107), .Z(n3238) );
  XOR U5821 ( .A(n3239), .B(n3238), .Z(n3241) );
  AND U5822 ( .A(y[7691]), .B(x[495]), .Z(n3928) );
  NAND U5823 ( .A(n3928), .B(n3109), .Z(n3113) );
  NAND U5824 ( .A(n3111), .B(n3110), .Z(n3112) );
  NAND U5825 ( .A(n3113), .B(n3112), .Z(n3294) );
  AND U5826 ( .A(o[20]), .B(n3114), .Z(n3316) );
  AND U5827 ( .A(x[480]), .B(y[7701]), .Z(n3313) );
  AND U5828 ( .A(y[7680]), .B(x[501]), .Z(n3314) );
  XOR U5829 ( .A(n3313), .B(n3314), .Z(n3315) );
  XOR U5830 ( .A(n3316), .B(n3315), .Z(n3292) );
  AND U5831 ( .A(y[7696]), .B(x[485]), .Z(n3300) );
  AND U5832 ( .A(x[496]), .B(y[7685]), .Z(n3299) );
  XOR U5833 ( .A(n3300), .B(n3299), .Z(n3298) );
  AND U5834 ( .A(y[7686]), .B(x[495]), .Z(n3297) );
  XOR U5835 ( .A(n3298), .B(n3297), .Z(n3291) );
  XOR U5836 ( .A(n3292), .B(n3291), .Z(n3293) );
  XOR U5837 ( .A(n3294), .B(n3293), .Z(n3240) );
  XOR U5838 ( .A(n3241), .B(n3240), .Z(n3257) );
  NANDN U5839 ( .A(n3116), .B(n3115), .Z(n3120) );
  NANDN U5840 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U5841 ( .A(n3120), .B(n3119), .Z(n3256) );
  NANDN U5842 ( .A(n3122), .B(n3121), .Z(n3126) );
  NANDN U5843 ( .A(n3124), .B(n3123), .Z(n3125) );
  NAND U5844 ( .A(n3126), .B(n3125), .Z(n3259) );
  NANDN U5845 ( .A(n3128), .B(n3127), .Z(n3132) );
  NAND U5846 ( .A(n3130), .B(n3129), .Z(n3131) );
  AND U5847 ( .A(n3132), .B(n3131), .Z(n3232) );
  XOR U5848 ( .A(n3234), .B(n3235), .Z(n3229) );
  NANDN U5849 ( .A(n3134), .B(n3133), .Z(n3138) );
  NAND U5850 ( .A(n3136), .B(n3135), .Z(n3137) );
  AND U5851 ( .A(n3138), .B(n3137), .Z(n3332) );
  AND U5852 ( .A(x[490]), .B(y[7684]), .Z(n3139) );
  NAND U5853 ( .A(n3933), .B(n3139), .Z(n3143) );
  NANDN U5854 ( .A(n3141), .B(n3140), .Z(n3142) );
  AND U5855 ( .A(n3143), .B(n3142), .Z(n3263) );
  AND U5856 ( .A(y[7687]), .B(x[483]), .Z(n3144) );
  NAND U5857 ( .A(n4429), .B(n3144), .Z(n3148) );
  NAND U5858 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U5859 ( .A(n3148), .B(n3147), .Z(n3253) );
  AND U5860 ( .A(y[7682]), .B(x[499]), .Z(n3150) );
  NAND U5861 ( .A(y[7690]), .B(x[491]), .Z(n3149) );
  XNOR U5862 ( .A(n3150), .B(n3149), .Z(n3270) );
  AND U5863 ( .A(y[7681]), .B(x[500]), .Z(n3312) );
  XOR U5864 ( .A(o[21]), .B(n3312), .Z(n3269) );
  XOR U5865 ( .A(n3270), .B(n3269), .Z(n3251) );
  AND U5866 ( .A(y[7683]), .B(x[498]), .Z(n3152) );
  NAND U5867 ( .A(x[490]), .B(y[7691]), .Z(n3151) );
  XNOR U5868 ( .A(n3152), .B(n3151), .Z(n3320) );
  AND U5869 ( .A(y[7700]), .B(x[481]), .Z(n3321) );
  XOR U5870 ( .A(n3320), .B(n3321), .Z(n3250) );
  XOR U5871 ( .A(n3251), .B(n3250), .Z(n3252) );
  XOR U5872 ( .A(n3253), .B(n3252), .Z(n3262) );
  AND U5873 ( .A(y[7694]), .B(x[487]), .Z(n3491) );
  AND U5874 ( .A(x[486]), .B(y[7695]), .Z(n3154) );
  NAND U5875 ( .A(x[494]), .B(y[7687]), .Z(n3153) );
  XNOR U5876 ( .A(n3154), .B(n3153), .Z(n3324) );
  XNOR U5877 ( .A(n3491), .B(n3324), .Z(n3282) );
  NAND U5878 ( .A(x[489]), .B(y[7692]), .Z(n3280) );
  NAND U5879 ( .A(x[488]), .B(y[7693]), .Z(n3279) );
  XOR U5880 ( .A(n3280), .B(n3279), .Z(n3281) );
  XNOR U5881 ( .A(n3282), .B(n3281), .Z(n3287) );
  AND U5882 ( .A(y[7689]), .B(x[492]), .Z(n3156) );
  NAND U5883 ( .A(y[7684]), .B(x[497]), .Z(n3155) );
  XNOR U5884 ( .A(n3156), .B(n3155), .Z(n3273) );
  AND U5885 ( .A(y[7699]), .B(x[482]), .Z(n3274) );
  XOR U5886 ( .A(n3273), .B(n3274), .Z(n3286) );
  AND U5887 ( .A(x[493]), .B(y[7688]), .Z(n3158) );
  NAND U5888 ( .A(x[483]), .B(y[7698]), .Z(n3157) );
  XNOR U5889 ( .A(n3158), .B(n3157), .Z(n3308) );
  AND U5890 ( .A(x[484]), .B(y[7697]), .Z(n3309) );
  XOR U5891 ( .A(n3308), .B(n3309), .Z(n3285) );
  XOR U5892 ( .A(n3286), .B(n3285), .Z(n3288) );
  XOR U5893 ( .A(n3287), .B(n3288), .Z(n3247) );
  NAND U5894 ( .A(n3300), .B(n3159), .Z(n3163) );
  NAND U5895 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U5896 ( .A(n3163), .B(n3162), .Z(n3245) );
  NAND U5897 ( .A(n3165), .B(n3164), .Z(n3169) );
  NAND U5898 ( .A(n3167), .B(n3166), .Z(n3168) );
  NAND U5899 ( .A(n3169), .B(n3168), .Z(n3244) );
  XOR U5900 ( .A(n3245), .B(n3244), .Z(n3246) );
  XOR U5901 ( .A(n3247), .B(n3246), .Z(n3264) );
  XOR U5902 ( .A(n3265), .B(n3264), .Z(n3330) );
  NANDN U5903 ( .A(n3171), .B(n3170), .Z(n3175) );
  NAND U5904 ( .A(n3173), .B(n3172), .Z(n3174) );
  NAND U5905 ( .A(n3175), .B(n3174), .Z(n3337) );
  NAND U5906 ( .A(n3177), .B(n3176), .Z(n3181) );
  NANDN U5907 ( .A(n3179), .B(n3178), .Z(n3180) );
  NAND U5908 ( .A(n3181), .B(n3180), .Z(n3336) );
  NAND U5909 ( .A(n3183), .B(n3182), .Z(n3187) );
  NANDN U5910 ( .A(n3185), .B(n3184), .Z(n3186) );
  NAND U5911 ( .A(n3187), .B(n3186), .Z(n3335) );
  XOR U5912 ( .A(n3336), .B(n3335), .Z(n3338) );
  XOR U5913 ( .A(n3337), .B(n3338), .Z(n3329) );
  XOR U5914 ( .A(n3330), .B(n3329), .Z(n3331) );
  IV U5915 ( .A(n3227), .Z(n3194) );
  NAND U5916 ( .A(n3189), .B(n3188), .Z(n3193) );
  NANDN U5917 ( .A(n3191), .B(n3190), .Z(n3192) );
  NAND U5918 ( .A(n3193), .B(n3192), .Z(n3226) );
  XOR U5919 ( .A(n3194), .B(n3226), .Z(n3228) );
  NANDN U5920 ( .A(n3196), .B(n3195), .Z(n3200) );
  NANDN U5921 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U5922 ( .A(n3200), .B(n3199), .Z(n3220) );
  XNOR U5923 ( .A(n3220), .B(n3219), .Z(n3222) );
  XNOR U5924 ( .A(n3221), .B(n3222), .Z(n3225) );
  NAND U5925 ( .A(n3206), .B(n3205), .Z(n3210) );
  NAND U5926 ( .A(n3208), .B(n3207), .Z(n3209) );
  AND U5927 ( .A(n3210), .B(n3209), .Z(n3223) );
  OR U5928 ( .A(n3213), .B(n3211), .Z(n3217) );
  ANDN U5929 ( .B(n3213), .A(n3212), .Z(n3215) );
  OR U5930 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U5931 ( .A(n3217), .B(n3216), .Z(n3224) );
  XNOR U5932 ( .A(n3223), .B(n3224), .Z(n3218) );
  XNOR U5933 ( .A(n3225), .B(n3218), .Z(N54) );
  NANDN U5934 ( .A(n3227), .B(n3226), .Z(n3231) );
  NANDN U5935 ( .A(n3229), .B(n3228), .Z(n3230) );
  AND U5936 ( .A(n3231), .B(n3230), .Z(n3466) );
  NANDN U5937 ( .A(n3233), .B(n3232), .Z(n3237) );
  NAND U5938 ( .A(n3235), .B(n3234), .Z(n3236) );
  NAND U5939 ( .A(n3237), .B(n3236), .Z(n3464) );
  NAND U5940 ( .A(n3239), .B(n3238), .Z(n3243) );
  NAND U5941 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U5942 ( .A(n3243), .B(n3242), .Z(n3351) );
  NAND U5943 ( .A(n3245), .B(n3244), .Z(n3249) );
  NAND U5944 ( .A(n3247), .B(n3246), .Z(n3248) );
  NAND U5945 ( .A(n3249), .B(n3248), .Z(n3349) );
  NAND U5946 ( .A(n3251), .B(n3250), .Z(n3255) );
  NAND U5947 ( .A(n3253), .B(n3252), .Z(n3254) );
  NAND U5948 ( .A(n3255), .B(n3254), .Z(n3348) );
  XOR U5949 ( .A(n3349), .B(n3348), .Z(n3350) );
  XOR U5950 ( .A(n3351), .B(n3350), .Z(n3455) );
  NANDN U5951 ( .A(n3257), .B(n3256), .Z(n3261) );
  NANDN U5952 ( .A(n3259), .B(n3258), .Z(n3260) );
  NAND U5953 ( .A(n3261), .B(n3260), .Z(n3456) );
  NANDN U5954 ( .A(n3263), .B(n3262), .Z(n3267) );
  NAND U5955 ( .A(n3265), .B(n3264), .Z(n3266) );
  AND U5956 ( .A(n3267), .B(n3266), .Z(n3452) );
  AND U5957 ( .A(x[499]), .B(y[7690]), .Z(n4462) );
  NAND U5958 ( .A(n4462), .B(n3268), .Z(n3272) );
  NAND U5959 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U5960 ( .A(n3272), .B(n3271), .Z(n3444) );
  NANDN U5961 ( .A(n3942), .B(n3398), .Z(n3276) );
  NAND U5962 ( .A(n3274), .B(n3273), .Z(n3275) );
  NAND U5963 ( .A(n3276), .B(n3275), .Z(n3374) );
  AND U5964 ( .A(y[7697]), .B(x[485]), .Z(n3419) );
  AND U5965 ( .A(x[497]), .B(y[7685]), .Z(n3420) );
  XOR U5966 ( .A(n3419), .B(n3420), .Z(n3421) );
  AND U5967 ( .A(y[7686]), .B(x[496]), .Z(n3422) );
  XOR U5968 ( .A(n3421), .B(n3422), .Z(n3373) );
  AND U5969 ( .A(y[7684]), .B(x[498]), .Z(n3278) );
  NAND U5970 ( .A(y[7690]), .B(x[492]), .Z(n3277) );
  XNOR U5971 ( .A(n3278), .B(n3277), .Z(n3400) );
  AND U5972 ( .A(x[484]), .B(y[7698]), .Z(n3399) );
  XOR U5973 ( .A(n3400), .B(n3399), .Z(n3372) );
  XOR U5974 ( .A(n3373), .B(n3372), .Z(n3375) );
  XOR U5975 ( .A(n3374), .B(n3375), .Z(n3443) );
  XOR U5976 ( .A(n3444), .B(n3443), .Z(n3445) );
  NAND U5977 ( .A(n3280), .B(n3279), .Z(n3284) );
  NAND U5978 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U5979 ( .A(n3284), .B(n3283), .Z(n3446) );
  XOR U5980 ( .A(n3445), .B(n3446), .Z(n3450) );
  NAND U5981 ( .A(n3286), .B(n3285), .Z(n3290) );
  NAND U5982 ( .A(n3288), .B(n3287), .Z(n3289) );
  NAND U5983 ( .A(n3290), .B(n3289), .Z(n3432) );
  NAND U5984 ( .A(n3292), .B(n3291), .Z(n3296) );
  NAND U5985 ( .A(n3294), .B(n3293), .Z(n3295) );
  NAND U5986 ( .A(n3296), .B(n3295), .Z(n3431) );
  XOR U5987 ( .A(n3432), .B(n3431), .Z(n3434) );
  AND U5988 ( .A(n3298), .B(n3297), .Z(n3302) );
  NAND U5989 ( .A(n3300), .B(n3299), .Z(n3301) );
  NANDN U5990 ( .A(n3302), .B(n3301), .Z(n3395) );
  AND U5991 ( .A(x[493]), .B(y[7689]), .Z(n3304) );
  NAND U5992 ( .A(y[7682]), .B(x[500]), .Z(n3303) );
  XNOR U5993 ( .A(n3304), .B(n3303), .Z(n3415) );
  AND U5994 ( .A(y[7700]), .B(x[482]), .Z(n3416) );
  XOR U5995 ( .A(n3415), .B(n3416), .Z(n3393) );
  AND U5996 ( .A(x[486]), .B(y[7696]), .Z(n3306) );
  NAND U5997 ( .A(x[495]), .B(y[7687]), .Z(n3305) );
  XNOR U5998 ( .A(n3306), .B(n3305), .Z(n3427) );
  XOR U5999 ( .A(n3393), .B(n3392), .Z(n3394) );
  XOR U6000 ( .A(n3395), .B(n3394), .Z(n3438) );
  AND U6001 ( .A(y[7698]), .B(x[493]), .Z(n4707) );
  NANDN U6002 ( .A(n3307), .B(n4707), .Z(n3311) );
  NAND U6003 ( .A(n3309), .B(n3308), .Z(n3310) );
  NAND U6004 ( .A(n3311), .B(n3310), .Z(n3363) );
  AND U6005 ( .A(x[481]), .B(y[7701]), .Z(n3386) );
  XOR U6006 ( .A(n3387), .B(n3386), .Z(n3385) );
  AND U6007 ( .A(o[21]), .B(n3312), .Z(n3384) );
  XOR U6008 ( .A(n3385), .B(n3384), .Z(n3361) );
  AND U6009 ( .A(y[7688]), .B(x[494]), .Z(n3378) );
  AND U6010 ( .A(y[7699]), .B(x[483]), .Z(n3379) );
  XOR U6011 ( .A(n3378), .B(n3379), .Z(n3380) );
  AND U6012 ( .A(y[7683]), .B(x[499]), .Z(n3381) );
  XOR U6013 ( .A(n3380), .B(n3381), .Z(n3360) );
  XOR U6014 ( .A(n3361), .B(n3360), .Z(n3362) );
  XOR U6015 ( .A(n3363), .B(n3362), .Z(n3437) );
  XOR U6016 ( .A(n3438), .B(n3437), .Z(n3440) );
  NAND U6017 ( .A(n3314), .B(n3313), .Z(n3318) );
  NAND U6018 ( .A(n3316), .B(n3315), .Z(n3317) );
  NAND U6019 ( .A(n3318), .B(n3317), .Z(n3355) );
  AND U6020 ( .A(y[7691]), .B(x[498]), .Z(n4465) );
  NAND U6021 ( .A(n4465), .B(n3319), .Z(n3323) );
  NAND U6022 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U6023 ( .A(n3323), .B(n3322), .Z(n3354) );
  XOR U6024 ( .A(n3355), .B(n3354), .Z(n3357) );
  AND U6025 ( .A(x[494]), .B(y[7695]), .Z(n4481) );
  NAND U6026 ( .A(n4481), .B(n3426), .Z(n3326) );
  NAND U6027 ( .A(n3491), .B(n3324), .Z(n3325) );
  NAND U6028 ( .A(n3326), .B(n3325), .Z(n3369) );
  AND U6029 ( .A(x[480]), .B(y[7702]), .Z(n3403) );
  AND U6030 ( .A(x[502]), .B(y[7680]), .Z(n3404) );
  XOR U6031 ( .A(n3403), .B(n3404), .Z(n3406) );
  AND U6032 ( .A(y[7681]), .B(x[501]), .Z(n3425) );
  XOR U6033 ( .A(o[22]), .B(n3425), .Z(n3405) );
  XOR U6034 ( .A(n3406), .B(n3405), .Z(n3367) );
  AND U6035 ( .A(x[487]), .B(y[7695]), .Z(n3328) );
  NAND U6036 ( .A(y[7694]), .B(x[488]), .Z(n3327) );
  XNOR U6037 ( .A(n3328), .B(n3327), .Z(n3409) );
  XOR U6038 ( .A(n3367), .B(n3366), .Z(n3368) );
  XOR U6039 ( .A(n3369), .B(n3368), .Z(n3356) );
  XOR U6040 ( .A(n3357), .B(n3356), .Z(n3439) );
  XOR U6041 ( .A(n3440), .B(n3439), .Z(n3433) );
  XOR U6042 ( .A(n3434), .B(n3433), .Z(n3449) );
  XOR U6043 ( .A(n3450), .B(n3449), .Z(n3451) );
  XOR U6044 ( .A(n3458), .B(n3457), .Z(n3345) );
  NAND U6045 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U6046 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U6047 ( .A(n3334), .B(n3333), .Z(n3343) );
  NAND U6048 ( .A(n3336), .B(n3335), .Z(n3340) );
  NAND U6049 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U6050 ( .A(n3340), .B(n3339), .Z(n3342) );
  XOR U6051 ( .A(n3345), .B(n3344), .Z(n3465) );
  XNOR U6052 ( .A(n3464), .B(n3465), .Z(n3467) );
  XOR U6053 ( .A(n3461), .B(n3463), .Z(n3341) );
  XOR U6054 ( .A(n3462), .B(n3341), .Z(N55) );
  NANDN U6055 ( .A(n3343), .B(n3342), .Z(n3347) );
  NAND U6056 ( .A(n3345), .B(n3344), .Z(n3346) );
  AND U6057 ( .A(n3347), .B(n3346), .Z(n3605) );
  NAND U6058 ( .A(n3349), .B(n3348), .Z(n3353) );
  NAND U6059 ( .A(n3351), .B(n3350), .Z(n3352) );
  NAND U6060 ( .A(n3353), .B(n3352), .Z(n3587) );
  NAND U6061 ( .A(n3355), .B(n3354), .Z(n3359) );
  NAND U6062 ( .A(n3357), .B(n3356), .Z(n3358) );
  NAND U6063 ( .A(n3359), .B(n3358), .Z(n3581) );
  NAND U6064 ( .A(n3361), .B(n3360), .Z(n3365) );
  NAND U6065 ( .A(n3363), .B(n3362), .Z(n3364) );
  NAND U6066 ( .A(n3365), .B(n3364), .Z(n3579) );
  NAND U6067 ( .A(n3367), .B(n3366), .Z(n3371) );
  NAND U6068 ( .A(n3369), .B(n3368), .Z(n3370) );
  NAND U6069 ( .A(n3371), .B(n3370), .Z(n3578) );
  XOR U6070 ( .A(n3579), .B(n3578), .Z(n3580) );
  XOR U6071 ( .A(n3581), .B(n3580), .Z(n3599) );
  NAND U6072 ( .A(n3373), .B(n3372), .Z(n3377) );
  NAND U6073 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND U6074 ( .A(n3377), .B(n3376), .Z(n3597) );
  NAND U6075 ( .A(n3379), .B(n3378), .Z(n3383) );
  NAND U6076 ( .A(n3381), .B(n3380), .Z(n3382) );
  NAND U6077 ( .A(n3383), .B(n3382), .Z(n3525) );
  AND U6078 ( .A(n3385), .B(n3384), .Z(n3389) );
  NAND U6079 ( .A(n3387), .B(n3386), .Z(n3388) );
  NANDN U6080 ( .A(n3389), .B(n3388), .Z(n3524) );
  XOR U6081 ( .A(n3525), .B(n3524), .Z(n3527) );
  AND U6082 ( .A(x[487]), .B(y[7696]), .Z(n3391) );
  NAND U6083 ( .A(y[7694]), .B(x[489]), .Z(n3390) );
  XNOR U6084 ( .A(n3391), .B(n3390), .Z(n3492) );
  AND U6085 ( .A(x[490]), .B(y[7693]), .Z(n3531) );
  XOR U6086 ( .A(n3530), .B(n3531), .Z(n3533) );
  AND U6087 ( .A(y[7697]), .B(x[486]), .Z(n3483) );
  AND U6088 ( .A(x[495]), .B(y[7688]), .Z(n3484) );
  XOR U6089 ( .A(n3483), .B(n3484), .Z(n3485) );
  AND U6090 ( .A(y[7692]), .B(x[491]), .Z(n3486) );
  XOR U6091 ( .A(n3485), .B(n3486), .Z(n3532) );
  XOR U6092 ( .A(n3533), .B(n3532), .Z(n3526) );
  XOR U6093 ( .A(n3527), .B(n3526), .Z(n3596) );
  XOR U6094 ( .A(n3597), .B(n3596), .Z(n3598) );
  XOR U6095 ( .A(n3599), .B(n3598), .Z(n3585) );
  NAND U6096 ( .A(n3393), .B(n3392), .Z(n3397) );
  NAND U6097 ( .A(n3395), .B(n3394), .Z(n3396) );
  NAND U6098 ( .A(n3397), .B(n3396), .Z(n3519) );
  AND U6099 ( .A(x[498]), .B(y[7690]), .Z(n4308) );
  NAND U6100 ( .A(n4308), .B(n3398), .Z(n3402) );
  NAND U6101 ( .A(n3400), .B(n3399), .Z(n3401) );
  NAND U6102 ( .A(n3402), .B(n3401), .Z(n3567) );
  NAND U6103 ( .A(n3404), .B(n3403), .Z(n3408) );
  NAND U6104 ( .A(n3406), .B(n3405), .Z(n3407) );
  NAND U6105 ( .A(n3408), .B(n3407), .Z(n3566) );
  XOR U6106 ( .A(n3567), .B(n3566), .Z(n3569) );
  NANDN U6107 ( .A(n3493), .B(n3491), .Z(n3412) );
  NANDN U6108 ( .A(n3410), .B(n3409), .Z(n3411) );
  NAND U6109 ( .A(n3412), .B(n3411), .Z(n3563) );
  AND U6110 ( .A(x[480]), .B(y[7703]), .Z(n3502) );
  AND U6111 ( .A(y[7680]), .B(x[503]), .Z(n3503) );
  XOR U6112 ( .A(n3502), .B(n3503), .Z(n3505) );
  AND U6113 ( .A(x[502]), .B(y[7681]), .Z(n3482) );
  XOR U6114 ( .A(o[23]), .B(n3482), .Z(n3504) );
  XOR U6115 ( .A(n3505), .B(n3504), .Z(n3561) );
  AND U6116 ( .A(y[7683]), .B(x[500]), .Z(n4117) );
  NAND U6117 ( .A(x[496]), .B(y[7687]), .Z(n3413) );
  XNOR U6118 ( .A(n4117), .B(n3413), .Z(n3478) );
  AND U6119 ( .A(y[7684]), .B(x[499]), .Z(n3479) );
  XOR U6120 ( .A(n3478), .B(n3479), .Z(n3560) );
  XOR U6121 ( .A(n3561), .B(n3560), .Z(n3562) );
  XOR U6122 ( .A(n3563), .B(n3562), .Z(n3568) );
  XOR U6123 ( .A(n3569), .B(n3568), .Z(n3518) );
  XOR U6124 ( .A(n3519), .B(n3518), .Z(n3521) );
  AND U6125 ( .A(x[500]), .B(y[7689]), .Z(n4492) );
  AND U6126 ( .A(x[493]), .B(y[7682]), .Z(n3414) );
  NAND U6127 ( .A(n4492), .B(n3414), .Z(n3418) );
  NAND U6128 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U6129 ( .A(n3418), .B(n3417), .Z(n3513) );
  NAND U6130 ( .A(n3420), .B(n3419), .Z(n3424) );
  NAND U6131 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U6132 ( .A(n3424), .B(n3423), .Z(n3575) );
  AND U6133 ( .A(x[493]), .B(y[7690]), .Z(n3548) );
  AND U6134 ( .A(x[482]), .B(y[7701]), .Z(n3549) );
  XOR U6135 ( .A(n3548), .B(n3549), .Z(n3550) );
  AND U6136 ( .A(x[501]), .B(y[7682]), .Z(n3551) );
  XOR U6137 ( .A(n3550), .B(n3551), .Z(n3573) );
  AND U6138 ( .A(y[7691]), .B(x[492]), .Z(n3496) );
  AND U6139 ( .A(x[481]), .B(y[7702]), .Z(n3497) );
  XOR U6140 ( .A(n3496), .B(n3497), .Z(n3499) );
  AND U6141 ( .A(o[22]), .B(n3425), .Z(n3498) );
  XOR U6142 ( .A(n3499), .B(n3498), .Z(n3572) );
  XOR U6143 ( .A(n3573), .B(n3572), .Z(n3574) );
  XOR U6144 ( .A(n3575), .B(n3574), .Z(n3512) );
  XOR U6145 ( .A(n3513), .B(n3512), .Z(n3515) );
  AND U6146 ( .A(x[495]), .B(y[7696]), .Z(n4717) );
  NAND U6147 ( .A(n4717), .B(n3426), .Z(n3430) );
  NANDN U6148 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U6149 ( .A(n3430), .B(n3429), .Z(n3557) );
  AND U6150 ( .A(y[7689]), .B(x[494]), .Z(n3542) );
  AND U6151 ( .A(y[7700]), .B(x[483]), .Z(n3543) );
  XOR U6152 ( .A(n3542), .B(n3543), .Z(n3544) );
  AND U6153 ( .A(x[484]), .B(y[7699]), .Z(n3545) );
  XOR U6154 ( .A(n3544), .B(n3545), .Z(n3555) );
  AND U6155 ( .A(y[7698]), .B(x[485]), .Z(n3536) );
  AND U6156 ( .A(x[498]), .B(y[7685]), .Z(n3537) );
  XOR U6157 ( .A(n3536), .B(n3537), .Z(n3538) );
  AND U6158 ( .A(x[497]), .B(y[7686]), .Z(n3539) );
  XOR U6159 ( .A(n3538), .B(n3539), .Z(n3554) );
  XOR U6160 ( .A(n3555), .B(n3554), .Z(n3556) );
  XOR U6161 ( .A(n3557), .B(n3556), .Z(n3514) );
  XOR U6162 ( .A(n3515), .B(n3514), .Z(n3520) );
  XOR U6163 ( .A(n3521), .B(n3520), .Z(n3584) );
  XOR U6164 ( .A(n3585), .B(n3584), .Z(n3586) );
  XOR U6165 ( .A(n3587), .B(n3586), .Z(n3474) );
  NAND U6166 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U6167 ( .A(n3434), .B(n3433), .Z(n3435) );
  NAND U6168 ( .A(n3436), .B(n3435), .Z(n3593) );
  NAND U6169 ( .A(n3438), .B(n3437), .Z(n3442) );
  NAND U6170 ( .A(n3440), .B(n3439), .Z(n3441) );
  NAND U6171 ( .A(n3442), .B(n3441), .Z(n3591) );
  NAND U6172 ( .A(n3444), .B(n3443), .Z(n3448) );
  NAND U6173 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U6174 ( .A(n3448), .B(n3447), .Z(n3590) );
  XOR U6175 ( .A(n3591), .B(n3590), .Z(n3592) );
  XOR U6176 ( .A(n3593), .B(n3592), .Z(n3472) );
  NAND U6177 ( .A(n3450), .B(n3449), .Z(n3454) );
  NANDN U6178 ( .A(n3452), .B(n3451), .Z(n3453) );
  AND U6179 ( .A(n3454), .B(n3453), .Z(n3471) );
  NANDN U6180 ( .A(n3456), .B(n3455), .Z(n3460) );
  NAND U6181 ( .A(n3458), .B(n3457), .Z(n3459) );
  NAND U6182 ( .A(n3460), .B(n3459), .Z(n3603) );
  XNOR U6183 ( .A(n3605), .B(n3604), .Z(n3610) );
  NAND U6184 ( .A(n3465), .B(n3464), .Z(n3469) );
  NANDN U6185 ( .A(n3467), .B(n3466), .Z(n3468) );
  AND U6186 ( .A(n3469), .B(n3468), .Z(n3608) );
  XOR U6187 ( .A(n3609), .B(n3608), .Z(n3470) );
  XNOR U6188 ( .A(n3610), .B(n3470), .Z(N56) );
  NANDN U6189 ( .A(n3472), .B(n3471), .Z(n3476) );
  NANDN U6190 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U6191 ( .A(n3476), .B(n3475), .Z(n3748) );
  AND U6192 ( .A(y[7687]), .B(x[500]), .Z(n3477) );
  NAND U6193 ( .A(n3477), .B(n3636), .Z(n3481) );
  NAND U6194 ( .A(n3479), .B(n3478), .Z(n3480) );
  NAND U6195 ( .A(n3481), .B(n3480), .Z(n3656) );
  AND U6196 ( .A(x[502]), .B(y[7682]), .Z(n3677) );
  XOR U6197 ( .A(n3678), .B(n3677), .Z(n3676) );
  NAND U6198 ( .A(x[482]), .B(y[7702]), .Z(n3675) );
  AND U6199 ( .A(x[481]), .B(y[7703]), .Z(n3683) );
  XOR U6200 ( .A(n3684), .B(n3683), .Z(n3682) );
  AND U6201 ( .A(o[23]), .B(n3482), .Z(n3681) );
  XOR U6202 ( .A(n3682), .B(n3681), .Z(n3653) );
  XOR U6203 ( .A(n3654), .B(n3653), .Z(n3655) );
  XOR U6204 ( .A(n3656), .B(n3655), .Z(n3714) );
  NAND U6205 ( .A(n3484), .B(n3483), .Z(n3488) );
  NAND U6206 ( .A(n3486), .B(n3485), .Z(n3487) );
  NAND U6207 ( .A(n3488), .B(n3487), .Z(n3650) );
  AND U6208 ( .A(x[496]), .B(y[7688]), .Z(n3490) );
  NAND U6209 ( .A(y[7683]), .B(x[501]), .Z(n3489) );
  XNOR U6210 ( .A(n3490), .B(n3489), .Z(n3637) );
  AND U6211 ( .A(y[7699]), .B(x[485]), .Z(n3638) );
  XOR U6212 ( .A(n3637), .B(n3638), .Z(n3648) );
  AND U6213 ( .A(y[7698]), .B(x[486]), .Z(n4033) );
  AND U6214 ( .A(x[500]), .B(y[7684]), .Z(n3851) );
  XOR U6215 ( .A(n4033), .B(n3851), .Z(n3643) );
  AND U6216 ( .A(y[7685]), .B(x[499]), .Z(n3644) );
  XOR U6217 ( .A(n3643), .B(n3644), .Z(n3647) );
  XOR U6218 ( .A(n3648), .B(n3647), .Z(n3649) );
  XOR U6219 ( .A(n3650), .B(n3649), .Z(n3627) );
  NAND U6220 ( .A(n3778), .B(n3491), .Z(n3495) );
  NANDN U6221 ( .A(n3493), .B(n3492), .Z(n3494) );
  NAND U6222 ( .A(n3495), .B(n3494), .Z(n3625) );
  NAND U6223 ( .A(n3497), .B(n3496), .Z(n3501) );
  NAND U6224 ( .A(n3499), .B(n3498), .Z(n3500) );
  NAND U6225 ( .A(n3501), .B(n3500), .Z(n3624) );
  XOR U6226 ( .A(n3625), .B(n3624), .Z(n3626) );
  XOR U6227 ( .A(n3627), .B(n3626), .Z(n3713) );
  XOR U6228 ( .A(n3714), .B(n3713), .Z(n3716) );
  NAND U6229 ( .A(n3503), .B(n3502), .Z(n3507) );
  NAND U6230 ( .A(n3505), .B(n3504), .Z(n3506) );
  AND U6231 ( .A(n3507), .B(n3506), .Z(n3708) );
  AND U6232 ( .A(x[483]), .B(y[7701]), .Z(n3697) );
  XOR U6233 ( .A(n3698), .B(n3697), .Z(n3696) );
  AND U6234 ( .A(x[484]), .B(y[7700]), .Z(n3695) );
  XOR U6235 ( .A(n3696), .B(n3695), .Z(n3707) );
  AND U6236 ( .A(y[7695]), .B(x[489]), .Z(n3509) );
  NAND U6237 ( .A(y[7694]), .B(x[490]), .Z(n3508) );
  XNOR U6238 ( .A(n3509), .B(n3508), .Z(n3667) );
  AND U6239 ( .A(y[7690]), .B(x[494]), .Z(n3511) );
  NAND U6240 ( .A(y[7696]), .B(x[488]), .Z(n3510) );
  XNOR U6241 ( .A(n3511), .B(n3510), .Z(n3671) );
  AND U6242 ( .A(y[7693]), .B(x[491]), .Z(n3672) );
  XOR U6243 ( .A(n3671), .B(n3672), .Z(n3666) );
  XOR U6244 ( .A(n3667), .B(n3666), .Z(n3709) );
  XOR U6245 ( .A(n3710), .B(n3709), .Z(n3715) );
  XNOR U6246 ( .A(n3716), .B(n3715), .Z(n3726) );
  NAND U6247 ( .A(n3513), .B(n3512), .Z(n3517) );
  NAND U6248 ( .A(n3515), .B(n3514), .Z(n3516) );
  AND U6249 ( .A(n3517), .B(n3516), .Z(n3725) );
  XOR U6250 ( .A(n3726), .B(n3725), .Z(n3727) );
  NAND U6251 ( .A(n3519), .B(n3518), .Z(n3523) );
  NAND U6252 ( .A(n3521), .B(n3520), .Z(n3522) );
  AND U6253 ( .A(n3523), .B(n3522), .Z(n3728) );
  XOR U6254 ( .A(n3727), .B(n3728), .Z(n3734) );
  NAND U6255 ( .A(n3525), .B(n3524), .Z(n3529) );
  NAND U6256 ( .A(n3527), .B(n3526), .Z(n3528) );
  NAND U6257 ( .A(n3529), .B(n3528), .Z(n3722) );
  NAND U6258 ( .A(n3531), .B(n3530), .Z(n3535) );
  NAND U6259 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U6260 ( .A(n3535), .B(n3534), .Z(n3720) );
  NAND U6261 ( .A(n3537), .B(n3536), .Z(n3541) );
  NAND U6262 ( .A(n3539), .B(n3538), .Z(n3540) );
  NAND U6263 ( .A(n3541), .B(n3540), .Z(n3633) );
  AND U6264 ( .A(y[7704]), .B(x[480]), .Z(n3701) );
  AND U6265 ( .A(y[7680]), .B(x[504]), .Z(n3702) );
  XOR U6266 ( .A(n3701), .B(n3702), .Z(n3703) );
  NAND U6267 ( .A(y[7681]), .B(x[503]), .Z(n3694) );
  XNOR U6268 ( .A(o[24]), .B(n3694), .Z(n3704) );
  XOR U6269 ( .A(n3703), .B(n3704), .Z(n3631) );
  AND U6270 ( .A(y[7697]), .B(x[487]), .Z(n3687) );
  NAND U6271 ( .A(y[7686]), .B(x[498]), .Z(n3688) );
  NAND U6272 ( .A(x[497]), .B(y[7687]), .Z(n3690) );
  XOR U6273 ( .A(n3631), .B(n3630), .Z(n3632) );
  XOR U6274 ( .A(n3633), .B(n3632), .Z(n3621) );
  NAND U6275 ( .A(n3543), .B(n3542), .Z(n3547) );
  NAND U6276 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U6277 ( .A(n3547), .B(n3546), .Z(n3619) );
  NAND U6278 ( .A(n3549), .B(n3548), .Z(n3553) );
  NAND U6279 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U6280 ( .A(n3553), .B(n3552), .Z(n3618) );
  XOR U6281 ( .A(n3619), .B(n3618), .Z(n3620) );
  XOR U6282 ( .A(n3621), .B(n3620), .Z(n3719) );
  XOR U6283 ( .A(n3720), .B(n3719), .Z(n3721) );
  XNOR U6284 ( .A(n3722), .B(n3721), .Z(n3614) );
  NAND U6285 ( .A(n3555), .B(n3554), .Z(n3559) );
  NAND U6286 ( .A(n3557), .B(n3556), .Z(n3558) );
  AND U6287 ( .A(n3559), .B(n3558), .Z(n3659) );
  NAND U6288 ( .A(n3561), .B(n3560), .Z(n3565) );
  NAND U6289 ( .A(n3563), .B(n3562), .Z(n3564) );
  NAND U6290 ( .A(n3565), .B(n3564), .Z(n3660) );
  NAND U6291 ( .A(n3567), .B(n3566), .Z(n3571) );
  NAND U6292 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U6293 ( .A(n3571), .B(n3570), .Z(n3662) );
  NAND U6294 ( .A(n3573), .B(n3572), .Z(n3577) );
  NAND U6295 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U6296 ( .A(n3577), .B(n3576), .Z(n3613) );
  XOR U6297 ( .A(n3612), .B(n3613), .Z(n3615) );
  XOR U6298 ( .A(n3614), .B(n3615), .Z(n3731) );
  NAND U6299 ( .A(n3579), .B(n3578), .Z(n3583) );
  NAND U6300 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U6301 ( .A(n3583), .B(n3582), .Z(n3732) );
  XOR U6302 ( .A(n3731), .B(n3732), .Z(n3733) );
  XNOR U6303 ( .A(n3734), .B(n3733), .Z(n3746) );
  NAND U6304 ( .A(n3585), .B(n3584), .Z(n3589) );
  NAND U6305 ( .A(n3587), .B(n3586), .Z(n3588) );
  NAND U6306 ( .A(n3589), .B(n3588), .Z(n3740) );
  NAND U6307 ( .A(n3591), .B(n3590), .Z(n3595) );
  NAND U6308 ( .A(n3593), .B(n3592), .Z(n3594) );
  NAND U6309 ( .A(n3595), .B(n3594), .Z(n3738) );
  NAND U6310 ( .A(n3597), .B(n3596), .Z(n3601) );
  NAND U6311 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND U6312 ( .A(n3601), .B(n3600), .Z(n3737) );
  XOR U6313 ( .A(n3738), .B(n3737), .Z(n3739) );
  XNOR U6314 ( .A(n3740), .B(n3739), .Z(n3747) );
  XOR U6315 ( .A(n3746), .B(n3747), .Z(n3749) );
  XNOR U6316 ( .A(n3748), .B(n3749), .Z(n3745) );
  NANDN U6317 ( .A(n3603), .B(n3602), .Z(n3607) );
  NAND U6318 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U6319 ( .A(n3607), .B(n3606), .Z(n3743) );
  XOR U6320 ( .A(n3743), .B(n3744), .Z(n3611) );
  XNOR U6321 ( .A(n3745), .B(n3611), .Z(N57) );
  NAND U6322 ( .A(n3613), .B(n3612), .Z(n3617) );
  NAND U6323 ( .A(n3615), .B(n3614), .Z(n3616) );
  AND U6324 ( .A(n3617), .B(n3616), .Z(n3762) );
  NAND U6325 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U6326 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U6327 ( .A(n3623), .B(n3622), .Z(n3766) );
  NAND U6328 ( .A(n3625), .B(n3624), .Z(n3629) );
  NAND U6329 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U6330 ( .A(n3629), .B(n3628), .Z(n3765) );
  XOR U6331 ( .A(n3766), .B(n3765), .Z(n3768) );
  NAND U6332 ( .A(n3631), .B(n3630), .Z(n3635) );
  NAND U6333 ( .A(n3633), .B(n3632), .Z(n3634) );
  AND U6334 ( .A(n3635), .B(n3634), .Z(n3798) );
  AND U6335 ( .A(x[501]), .B(y[7688]), .Z(n4612) );
  NAND U6336 ( .A(n4612), .B(n3636), .Z(n3640) );
  NAND U6337 ( .A(n3638), .B(n3637), .Z(n3639) );
  NAND U6338 ( .A(n3640), .B(n3639), .Z(n3871) );
  AND U6339 ( .A(x[502]), .B(y[7683]), .Z(n3840) );
  AND U6340 ( .A(y[7700]), .B(x[485]), .Z(n3839) );
  NAND U6341 ( .A(x[497]), .B(y[7688]), .Z(n3838) );
  XOR U6342 ( .A(n3839), .B(n3838), .Z(n3841) );
  XNOR U6343 ( .A(n3840), .B(n3841), .Z(n3869) );
  AND U6344 ( .A(y[7685]), .B(x[500]), .Z(n3642) );
  NAND U6345 ( .A(y[7684]), .B(x[501]), .Z(n3641) );
  XNOR U6346 ( .A(n3642), .B(n3641), .Z(n3852) );
  AND U6347 ( .A(y[7686]), .B(x[499]), .Z(n3853) );
  XOR U6348 ( .A(n3852), .B(n3853), .Z(n3868) );
  XOR U6349 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U6350 ( .A(n3871), .B(n3870), .Z(n3796) );
  NAND U6351 ( .A(n3851), .B(n4033), .Z(n3646) );
  NAND U6352 ( .A(n3644), .B(n3643), .Z(n3645) );
  AND U6353 ( .A(n3646), .B(n3645), .Z(n3877) );
  AND U6354 ( .A(x[495]), .B(y[7690]), .Z(n3858) );
  AND U6355 ( .A(y[7687]), .B(x[498]), .Z(n3857) );
  NAND U6356 ( .A(y[7699]), .B(x[486]), .Z(n3856) );
  XOR U6357 ( .A(n3857), .B(n3856), .Z(n3859) );
  XNOR U6358 ( .A(n3858), .B(n3859), .Z(n3875) );
  AND U6359 ( .A(x[503]), .B(y[7682]), .Z(n3834) );
  AND U6360 ( .A(x[484]), .B(y[7701]), .Z(n3833) );
  NAND U6361 ( .A(y[7689]), .B(x[496]), .Z(n3832) );
  XOR U6362 ( .A(n3833), .B(n3832), .Z(n3835) );
  XNOR U6363 ( .A(n3834), .B(n3835), .Z(n3874) );
  XOR U6364 ( .A(n3875), .B(n3874), .Z(n3876) );
  XOR U6365 ( .A(n3877), .B(n3876), .Z(n3795) );
  XNOR U6366 ( .A(n3798), .B(n3797), .Z(n3810) );
  NAND U6367 ( .A(n3648), .B(n3647), .Z(n3652) );
  NAND U6368 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND U6369 ( .A(n3652), .B(n3651), .Z(n3808) );
  NAND U6370 ( .A(n3654), .B(n3653), .Z(n3658) );
  NAND U6371 ( .A(n3656), .B(n3655), .Z(n3657) );
  NAND U6372 ( .A(n3658), .B(n3657), .Z(n3807) );
  XOR U6373 ( .A(n3808), .B(n3807), .Z(n3809) );
  XOR U6374 ( .A(n3810), .B(n3809), .Z(n3767) );
  XOR U6375 ( .A(n3768), .B(n3767), .Z(n3760) );
  NANDN U6376 ( .A(n3660), .B(n3659), .Z(n3664) );
  NANDN U6377 ( .A(n3662), .B(n3661), .Z(n3663) );
  NAND U6378 ( .A(n3664), .B(n3663), .Z(n3759) );
  NANDN U6379 ( .A(n3777), .B(n3665), .Z(n3669) );
  NAND U6380 ( .A(n3667), .B(n3666), .Z(n3668) );
  NAND U6381 ( .A(n3669), .B(n3668), .Z(n3802) );
  AND U6382 ( .A(x[494]), .B(y[7696]), .Z(n4632) );
  NAND U6383 ( .A(n4632), .B(n3670), .Z(n3674) );
  NAND U6384 ( .A(n3672), .B(n3671), .Z(n3673) );
  NAND U6385 ( .A(n3674), .B(n3673), .Z(n3829) );
  AND U6386 ( .A(y[7694]), .B(x[491]), .Z(n3847) );
  AND U6387 ( .A(x[492]), .B(y[7693]), .Z(n3846) );
  NAND U6388 ( .A(y[7698]), .B(x[487]), .Z(n3845) );
  XOR U6389 ( .A(n3846), .B(n3845), .Z(n3848) );
  XNOR U6390 ( .A(n3847), .B(n3848), .Z(n3827) );
  NAND U6391 ( .A(y[7681]), .B(x[504]), .Z(n3844) );
  XNOR U6392 ( .A(o[25]), .B(n3844), .Z(n3814) );
  AND U6393 ( .A(y[7704]), .B(x[481]), .Z(n3815) );
  XOR U6394 ( .A(n3814), .B(n3815), .Z(n3816) );
  AND U6395 ( .A(y[7692]), .B(x[493]), .Z(n3817) );
  XOR U6396 ( .A(n3816), .B(n3817), .Z(n3826) );
  XOR U6397 ( .A(n3827), .B(n3826), .Z(n3828) );
  XOR U6398 ( .A(n3829), .B(n3828), .Z(n3801) );
  XOR U6399 ( .A(n3802), .B(n3801), .Z(n3804) );
  ANDN U6400 ( .B(n3676), .A(n3675), .Z(n3680) );
  NAND U6401 ( .A(n3678), .B(n3677), .Z(n3679) );
  NANDN U6402 ( .A(n3680), .B(n3679), .Z(n3790) );
  AND U6403 ( .A(n3682), .B(n3681), .Z(n3686) );
  NAND U6404 ( .A(n3684), .B(n3683), .Z(n3685) );
  NANDN U6405 ( .A(n3686), .B(n3685), .Z(n3789) );
  XOR U6406 ( .A(n3790), .B(n3789), .Z(n3792) );
  NANDN U6407 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U6408 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U6409 ( .A(n3692), .B(n3691), .Z(n3786) );
  AND U6410 ( .A(x[488]), .B(y[7697]), .Z(n3780) );
  XOR U6411 ( .A(n3778), .B(n3693), .Z(n3779) );
  XOR U6412 ( .A(n3780), .B(n3779), .Z(n3784) );
  ANDN U6413 ( .B(o[24]), .A(n3694), .Z(n3773) );
  AND U6414 ( .A(y[7680]), .B(x[505]), .Z(n3772) );
  NAND U6415 ( .A(x[480]), .B(y[7705]), .Z(n3771) );
  XOR U6416 ( .A(n3772), .B(n3771), .Z(n3774) );
  XNOR U6417 ( .A(n3773), .B(n3774), .Z(n3783) );
  XOR U6418 ( .A(n3784), .B(n3783), .Z(n3785) );
  XOR U6419 ( .A(n3786), .B(n3785), .Z(n3791) );
  XOR U6420 ( .A(n3792), .B(n3791), .Z(n3803) );
  XOR U6421 ( .A(n3804), .B(n3803), .Z(n3883) );
  AND U6422 ( .A(n3696), .B(n3695), .Z(n3700) );
  NAND U6423 ( .A(n3698), .B(n3697), .Z(n3699) );
  NANDN U6424 ( .A(n3700), .B(n3699), .Z(n3865) );
  NAND U6425 ( .A(n3702), .B(n3701), .Z(n3706) );
  NAND U6426 ( .A(n3704), .B(n3703), .Z(n3705) );
  NAND U6427 ( .A(n3706), .B(n3705), .Z(n3863) );
  AND U6428 ( .A(y[7691]), .B(x[494]), .Z(n3820) );
  AND U6429 ( .A(x[482]), .B(y[7703]), .Z(n3821) );
  XOR U6430 ( .A(n3820), .B(n3821), .Z(n3822) );
  AND U6431 ( .A(x[483]), .B(y[7702]), .Z(n3823) );
  XOR U6432 ( .A(n3822), .B(n3823), .Z(n3862) );
  XOR U6433 ( .A(n3863), .B(n3862), .Z(n3864) );
  XNOR U6434 ( .A(n3865), .B(n3864), .Z(n3880) );
  NANDN U6435 ( .A(n3708), .B(n3707), .Z(n3712) );
  NAND U6436 ( .A(n3710), .B(n3709), .Z(n3711) );
  AND U6437 ( .A(n3712), .B(n3711), .Z(n3881) );
  XOR U6438 ( .A(n3880), .B(n3881), .Z(n3882) );
  NAND U6439 ( .A(n3714), .B(n3713), .Z(n3718) );
  NAND U6440 ( .A(n3716), .B(n3715), .Z(n3717) );
  AND U6441 ( .A(n3718), .B(n3717), .Z(n3887) );
  XOR U6442 ( .A(n3886), .B(n3887), .Z(n3889) );
  NAND U6443 ( .A(n3720), .B(n3719), .Z(n3724) );
  NAND U6444 ( .A(n3722), .B(n3721), .Z(n3723) );
  AND U6445 ( .A(n3724), .B(n3723), .Z(n3888) );
  XOR U6446 ( .A(n3889), .B(n3888), .Z(n3754) );
  NAND U6447 ( .A(n3726), .B(n3725), .Z(n3730) );
  NAND U6448 ( .A(n3728), .B(n3727), .Z(n3729) );
  AND U6449 ( .A(n3730), .B(n3729), .Z(n3753) );
  XNOR U6450 ( .A(n3755), .B(n3756), .Z(n3896) );
  NAND U6451 ( .A(n3732), .B(n3731), .Z(n3736) );
  NAND U6452 ( .A(n3734), .B(n3733), .Z(n3735) );
  NAND U6453 ( .A(n3736), .B(n3735), .Z(n3895) );
  XOR U6454 ( .A(n3896), .B(n3895), .Z(n3898) );
  NAND U6455 ( .A(n3738), .B(n3737), .Z(n3742) );
  NAND U6456 ( .A(n3740), .B(n3739), .Z(n3741) );
  AND U6457 ( .A(n3742), .B(n3741), .Z(n3897) );
  XNOR U6458 ( .A(n3898), .B(n3897), .Z(n3894) );
  NANDN U6459 ( .A(n3747), .B(n3746), .Z(n3751) );
  NANDN U6460 ( .A(n3749), .B(n3748), .Z(n3750) );
  AND U6461 ( .A(n3751), .B(n3750), .Z(n3892) );
  XOR U6462 ( .A(n3893), .B(n3892), .Z(n3752) );
  XNOR U6463 ( .A(n3894), .B(n3752), .Z(N58) );
  NANDN U6464 ( .A(n3754), .B(n3753), .Z(n3758) );
  NAND U6465 ( .A(n3756), .B(n3755), .Z(n3757) );
  AND U6466 ( .A(n3758), .B(n3757), .Z(n3903) );
  NANDN U6467 ( .A(n3760), .B(n3759), .Z(n3764) );
  NANDN U6468 ( .A(n3762), .B(n3761), .Z(n3763) );
  AND U6469 ( .A(n3764), .B(n3763), .Z(n3902) );
  NAND U6470 ( .A(n3766), .B(n3765), .Z(n3770) );
  NAND U6471 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U6472 ( .A(n3770), .B(n3769), .Z(n4054) );
  AND U6473 ( .A(y[7704]), .B(x[482]), .Z(n3927) );
  XOR U6474 ( .A(n3928), .B(n3927), .Z(n3930) );
  AND U6475 ( .A(x[504]), .B(y[7682]), .Z(n3929) );
  XOR U6476 ( .A(n3930), .B(n3929), .Z(n3963) );
  NANDN U6477 ( .A(n3772), .B(n3771), .Z(n3776) );
  OR U6478 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U6479 ( .A(n3776), .B(n3775), .Z(n3964) );
  XNOR U6480 ( .A(n3963), .B(n3964), .Z(n3966) );
  NANDN U6481 ( .A(n3778), .B(n3777), .Z(n3782) );
  NANDN U6482 ( .A(n3780), .B(n3779), .Z(n3781) );
  AND U6483 ( .A(n3782), .B(n3781), .Z(n3965) );
  XNOR U6484 ( .A(n3966), .B(n3965), .Z(n4002) );
  NAND U6485 ( .A(n3784), .B(n3783), .Z(n3788) );
  NAND U6486 ( .A(n3786), .B(n3785), .Z(n3787) );
  AND U6487 ( .A(n3788), .B(n3787), .Z(n4001) );
  XOR U6488 ( .A(n4002), .B(n4001), .Z(n4003) );
  NAND U6489 ( .A(n3790), .B(n3789), .Z(n3794) );
  NAND U6490 ( .A(n3792), .B(n3791), .Z(n3793) );
  AND U6491 ( .A(n3794), .B(n3793), .Z(n4004) );
  XOR U6492 ( .A(n4003), .B(n4004), .Z(n4048) );
  NANDN U6493 ( .A(n3796), .B(n3795), .Z(n3800) );
  NAND U6494 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U6495 ( .A(n3800), .B(n3799), .Z(n4045) );
  NAND U6496 ( .A(n3802), .B(n3801), .Z(n3806) );
  NAND U6497 ( .A(n3804), .B(n3803), .Z(n3805) );
  AND U6498 ( .A(n3806), .B(n3805), .Z(n4046) );
  XOR U6499 ( .A(n4045), .B(n4046), .Z(n4047) );
  XNOR U6500 ( .A(n4048), .B(n4047), .Z(n4052) );
  NAND U6501 ( .A(n3808), .B(n3807), .Z(n3812) );
  NAND U6502 ( .A(n3810), .B(n3809), .Z(n3811) );
  NAND U6503 ( .A(n3812), .B(n3811), .Z(n3997) );
  AND U6504 ( .A(x[492]), .B(y[7694]), .Z(n4183) );
  AND U6505 ( .A(y[7701]), .B(x[485]), .Z(n3978) );
  XOR U6506 ( .A(n4183), .B(n3978), .Z(n3979) );
  NAND U6507 ( .A(x[490]), .B(y[7696]), .Z(n3980) );
  XNOR U6508 ( .A(n3979), .B(n3980), .Z(n4010) );
  NAND U6509 ( .A(x[486]), .B(y[7700]), .Z(n3813) );
  XNOR U6510 ( .A(n4278), .B(n3813), .Z(n4034) );
  NAND U6511 ( .A(x[489]), .B(y[7697]), .Z(n4035) );
  XNOR U6512 ( .A(n4034), .B(n4035), .Z(n4007) );
  NAND U6513 ( .A(y[7699]), .B(x[487]), .Z(n4008) );
  XOR U6514 ( .A(n4010), .B(n4009), .Z(n3954) );
  NAND U6515 ( .A(n3815), .B(n3814), .Z(n3819) );
  NAND U6516 ( .A(n3817), .B(n3816), .Z(n3818) );
  NAND U6517 ( .A(n3819), .B(n3818), .Z(n3952) );
  NAND U6518 ( .A(n3821), .B(n3820), .Z(n3825) );
  NAND U6519 ( .A(n3823), .B(n3822), .Z(n3824) );
  NAND U6520 ( .A(n3825), .B(n3824), .Z(n3951) );
  XOR U6521 ( .A(n3952), .B(n3951), .Z(n3953) );
  XNOR U6522 ( .A(n3954), .B(n3953), .Z(n3990) );
  NAND U6523 ( .A(n3827), .B(n3826), .Z(n3831) );
  NAND U6524 ( .A(n3829), .B(n3828), .Z(n3830) );
  AND U6525 ( .A(n3831), .B(n3830), .Z(n3989) );
  XOR U6526 ( .A(n3990), .B(n3989), .Z(n3992) );
  NANDN U6527 ( .A(n3833), .B(n3832), .Z(n3837) );
  OR U6528 ( .A(n3835), .B(n3834), .Z(n3836) );
  AND U6529 ( .A(n3837), .B(n3836), .Z(n3917) );
  NANDN U6530 ( .A(n3839), .B(n3838), .Z(n3843) );
  OR U6531 ( .A(n3841), .B(n3840), .Z(n3842) );
  NAND U6532 ( .A(n3843), .B(n3842), .Z(n3918) );
  XNOR U6533 ( .A(n3917), .B(n3918), .Z(n3920) );
  ANDN U6534 ( .B(o[25]), .A(n3844), .Z(n4028) );
  AND U6535 ( .A(y[7692]), .B(x[494]), .Z(n4027) );
  XOR U6536 ( .A(n4028), .B(n4027), .Z(n4030) );
  AND U6537 ( .A(x[481]), .B(y[7705]), .Z(n4029) );
  XOR U6538 ( .A(n4030), .B(n4029), .Z(n3969) );
  AND U6539 ( .A(y[7681]), .B(x[505]), .Z(n4038) );
  XOR U6540 ( .A(o[26]), .B(n4038), .Z(n3983) );
  NAND U6541 ( .A(y[7680]), .B(x[506]), .Z(n3984) );
  XNOR U6542 ( .A(n3983), .B(n3984), .Z(n3985) );
  NAND U6543 ( .A(x[480]), .B(y[7706]), .Z(n3986) );
  XOR U6544 ( .A(n3985), .B(n3986), .Z(n3970) );
  XNOR U6545 ( .A(n3969), .B(n3970), .Z(n3971) );
  NANDN U6546 ( .A(n3846), .B(n3845), .Z(n3850) );
  OR U6547 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U6548 ( .A(n3850), .B(n3849), .Z(n3972) );
  XNOR U6549 ( .A(n3971), .B(n3972), .Z(n3919) );
  XNOR U6550 ( .A(n3920), .B(n3919), .Z(n3960) );
  AND U6551 ( .A(x[501]), .B(y[7685]), .Z(n4021) );
  NAND U6552 ( .A(n3851), .B(n4021), .Z(n3855) );
  NAND U6553 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U6554 ( .A(n3855), .B(n3854), .Z(n3948) );
  XOR U6555 ( .A(n4022), .B(n4021), .Z(n4024) );
  NAND U6556 ( .A(y[7686]), .B(x[500]), .Z(n4023) );
  XNOR U6557 ( .A(n4024), .B(n4023), .Z(n3945) );
  NAND U6558 ( .A(y[7683]), .B(x[503]), .Z(n3934) );
  XNOR U6559 ( .A(n3933), .B(n3934), .Z(n3935) );
  NAND U6560 ( .A(x[502]), .B(y[7684]), .Z(n3936) );
  XNOR U6561 ( .A(n3935), .B(n3936), .Z(n3946) );
  XOR U6562 ( .A(n3945), .B(n3946), .Z(n3947) );
  XNOR U6563 ( .A(n3948), .B(n3947), .Z(n3958) );
  AND U6564 ( .A(x[483]), .B(y[7703]), .Z(n4014) );
  AND U6565 ( .A(y[7687]), .B(x[499]), .Z(n4013) );
  XOR U6566 ( .A(n4014), .B(n4013), .Z(n4016) );
  AND U6567 ( .A(y[7695]), .B(x[491]), .Z(n4015) );
  XOR U6568 ( .A(n4016), .B(n4015), .Z(n3924) );
  AND U6569 ( .A(x[484]), .B(y[7702]), .Z(n3939) );
  XOR U6570 ( .A(n3940), .B(n3939), .Z(n3941) );
  XOR U6571 ( .A(n3924), .B(n3923), .Z(n3926) );
  NANDN U6572 ( .A(n3857), .B(n3856), .Z(n3861) );
  OR U6573 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U6574 ( .A(n3861), .B(n3860), .Z(n3925) );
  XNOR U6575 ( .A(n3926), .B(n3925), .Z(n3957) );
  XOR U6576 ( .A(n3958), .B(n3957), .Z(n3959) );
  XOR U6577 ( .A(n3960), .B(n3959), .Z(n3991) );
  XNOR U6578 ( .A(n3992), .B(n3991), .Z(n3996) );
  NAND U6579 ( .A(n3863), .B(n3862), .Z(n3867) );
  NAND U6580 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U6581 ( .A(n3867), .B(n3866), .Z(n4042) );
  NAND U6582 ( .A(n3869), .B(n3868), .Z(n3873) );
  NAND U6583 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U6584 ( .A(n3873), .B(n3872), .Z(n4040) );
  NAND U6585 ( .A(n3875), .B(n3874), .Z(n3879) );
  NANDN U6586 ( .A(n3877), .B(n3876), .Z(n3878) );
  NAND U6587 ( .A(n3879), .B(n3878), .Z(n4039) );
  XOR U6588 ( .A(n3996), .B(n3995), .Z(n3998) );
  XOR U6589 ( .A(n3997), .B(n3998), .Z(n4051) );
  XOR U6590 ( .A(n4052), .B(n4051), .Z(n4053) );
  XOR U6591 ( .A(n4054), .B(n4053), .Z(n3914) );
  NAND U6592 ( .A(n3881), .B(n3880), .Z(n3885) );
  NANDN U6593 ( .A(n3883), .B(n3882), .Z(n3884) );
  AND U6594 ( .A(n3885), .B(n3884), .Z(n3911) );
  NAND U6595 ( .A(n3887), .B(n3886), .Z(n3891) );
  NAND U6596 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U6597 ( .A(n3891), .B(n3890), .Z(n3912) );
  XOR U6598 ( .A(n3911), .B(n3912), .Z(n3913) );
  XOR U6599 ( .A(n3914), .B(n3913), .Z(n3904) );
  XNOR U6600 ( .A(n3905), .B(n3904), .Z(n3910) );
  NAND U6601 ( .A(n3896), .B(n3895), .Z(n3900) );
  NAND U6602 ( .A(n3898), .B(n3897), .Z(n3899) );
  AND U6603 ( .A(n3900), .B(n3899), .Z(n3909) );
  XOR U6604 ( .A(n3908), .B(n3909), .Z(n3901) );
  XNOR U6605 ( .A(n3910), .B(n3901), .Z(N59) );
  NANDN U6606 ( .A(n3903), .B(n3902), .Z(n3907) );
  NAND U6607 ( .A(n3905), .B(n3904), .Z(n3906) );
  NAND U6608 ( .A(n3907), .B(n3906), .Z(n4065) );
  IV U6609 ( .A(n4065), .Z(n4064) );
  NAND U6610 ( .A(n3912), .B(n3911), .Z(n3916) );
  NAND U6611 ( .A(n3914), .B(n3913), .Z(n3915) );
  AND U6612 ( .A(n3916), .B(n3915), .Z(n4061) );
  NANDN U6613 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U6614 ( .A(n3920), .B(n3919), .Z(n3921) );
  AND U6615 ( .A(n3922), .B(n3921), .Z(n4097) );
  AND U6616 ( .A(n3928), .B(n3927), .Z(n3932) );
  NAND U6617 ( .A(n3930), .B(n3929), .Z(n3931) );
  NANDN U6618 ( .A(n3932), .B(n3931), .Z(n4156) );
  NANDN U6619 ( .A(n3934), .B(n3933), .Z(n3938) );
  NANDN U6620 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U6621 ( .A(n3938), .B(n3937), .Z(n4155) );
  XOR U6622 ( .A(n4156), .B(n4155), .Z(n4157) );
  AND U6623 ( .A(n3940), .B(n3939), .Z(n3944) );
  NANDN U6624 ( .A(n3942), .B(n3941), .Z(n3943) );
  NANDN U6625 ( .A(n3944), .B(n3943), .Z(n4169) );
  AND U6626 ( .A(x[480]), .B(y[7707]), .Z(n4135) );
  AND U6627 ( .A(y[7680]), .B(x[507]), .Z(n4134) );
  XOR U6628 ( .A(n4135), .B(n4134), .Z(n4137) );
  AND U6629 ( .A(x[506]), .B(y[7681]), .Z(n4146) );
  XOR U6630 ( .A(n4146), .B(o[27]), .Z(n4136) );
  XOR U6631 ( .A(n4137), .B(n4136), .Z(n4168) );
  AND U6632 ( .A(y[7698]), .B(x[489]), .Z(n4141) );
  AND U6633 ( .A(y[7686]), .B(x[501]), .Z(n4140) );
  XOR U6634 ( .A(n4141), .B(n4140), .Z(n4143) );
  AND U6635 ( .A(y[7689]), .B(x[498]), .Z(n4142) );
  XOR U6636 ( .A(n4143), .B(n4142), .Z(n4167) );
  XOR U6637 ( .A(n4168), .B(n4167), .Z(n4170) );
  XNOR U6638 ( .A(n4169), .B(n4170), .Z(n4158) );
  XOR U6639 ( .A(n4096), .B(n4095), .Z(n4098) );
  XOR U6640 ( .A(n4097), .B(n4098), .Z(n4215) );
  NAND U6641 ( .A(n3946), .B(n3945), .Z(n3950) );
  NAND U6642 ( .A(n3948), .B(n3947), .Z(n3949) );
  AND U6643 ( .A(n3950), .B(n3949), .Z(n4212) );
  NAND U6644 ( .A(n3952), .B(n3951), .Z(n3956) );
  NAND U6645 ( .A(n3954), .B(n3953), .Z(n3955) );
  NAND U6646 ( .A(n3956), .B(n3955), .Z(n4213) );
  NAND U6647 ( .A(n3958), .B(n3957), .Z(n3962) );
  NAND U6648 ( .A(n3960), .B(n3959), .Z(n3961) );
  AND U6649 ( .A(n3962), .B(n3961), .Z(n4200) );
  NANDN U6650 ( .A(n3964), .B(n3963), .Z(n3968) );
  NAND U6651 ( .A(n3966), .B(n3965), .Z(n3967) );
  AND U6652 ( .A(n3968), .B(n3967), .Z(n4092) );
  NANDN U6653 ( .A(n3970), .B(n3969), .Z(n3974) );
  NANDN U6654 ( .A(n3972), .B(n3971), .Z(n3973) );
  AND U6655 ( .A(n3974), .B(n3973), .Z(n4090) );
  AND U6656 ( .A(y[7688]), .B(x[499]), .Z(n4123) );
  AND U6657 ( .A(x[505]), .B(y[7682]), .Z(n4122) );
  XOR U6658 ( .A(n4123), .B(n4122), .Z(n4125) );
  AND U6659 ( .A(y[7701]), .B(x[486]), .Z(n4124) );
  XOR U6660 ( .A(n4125), .B(n4124), .Z(n4112) );
  AND U6661 ( .A(x[495]), .B(y[7692]), .Z(n4189) );
  AND U6662 ( .A(x[482]), .B(y[7705]), .Z(n4188) );
  XOR U6663 ( .A(n4189), .B(n4188), .Z(n4191) );
  AND U6664 ( .A(y[7704]), .B(x[483]), .Z(n4190) );
  XOR U6665 ( .A(n4191), .B(n4190), .Z(n4111) );
  XOR U6666 ( .A(n4112), .B(n4111), .Z(n4113) );
  NAND U6667 ( .A(y[7691]), .B(x[496]), .Z(n4173) );
  XOR U6668 ( .A(n4173), .B(n3975), .Z(n4176) );
  XOR U6669 ( .A(n4175), .B(n4176), .Z(n4185) );
  AND U6670 ( .A(y[7694]), .B(x[493]), .Z(n3977) );
  AND U6671 ( .A(y[7695]), .B(x[492]), .Z(n3976) );
  XOR U6672 ( .A(n3977), .B(n3976), .Z(n4184) );
  XNOR U6673 ( .A(n4113), .B(n4114), .Z(n4151) );
  AND U6674 ( .A(n4183), .B(n3978), .Z(n3982) );
  NANDN U6675 ( .A(n3980), .B(n3979), .Z(n3981) );
  NANDN U6676 ( .A(n3982), .B(n3981), .Z(n4150) );
  NANDN U6677 ( .A(n3984), .B(n3983), .Z(n3988) );
  NANDN U6678 ( .A(n3986), .B(n3985), .Z(n3987) );
  NAND U6679 ( .A(n3988), .B(n3987), .Z(n4149) );
  XNOR U6680 ( .A(n4150), .B(n4149), .Z(n4152) );
  XNOR U6681 ( .A(n4090), .B(n4089), .Z(n4091) );
  XOR U6682 ( .A(n4092), .B(n4091), .Z(n4201) );
  NAND U6683 ( .A(n3990), .B(n3989), .Z(n3994) );
  NAND U6684 ( .A(n3992), .B(n3991), .Z(n3993) );
  NAND U6685 ( .A(n3994), .B(n3993), .Z(n4203) );
  NAND U6686 ( .A(n3996), .B(n3995), .Z(n4000) );
  NAND U6687 ( .A(n3998), .B(n3997), .Z(n3999) );
  NAND U6688 ( .A(n4000), .B(n3999), .Z(n4079) );
  XOR U6689 ( .A(n4080), .B(n4079), .Z(n4074) );
  NAND U6690 ( .A(n4002), .B(n4001), .Z(n4006) );
  NAND U6691 ( .A(n4004), .B(n4003), .Z(n4005) );
  AND U6692 ( .A(n4006), .B(n4005), .Z(n4084) );
  NANDN U6693 ( .A(n4008), .B(n4007), .Z(n4012) );
  NAND U6694 ( .A(n4010), .B(n4009), .Z(n4011) );
  AND U6695 ( .A(n4012), .B(n4011), .Z(n4209) );
  NAND U6696 ( .A(n4014), .B(n4013), .Z(n4018) );
  NAND U6697 ( .A(n4016), .B(n4015), .Z(n4017) );
  AND U6698 ( .A(n4018), .B(n4017), .Z(n4110) );
  AND U6699 ( .A(y[7683]), .B(x[504]), .Z(n4020) );
  NAND U6700 ( .A(x[500]), .B(y[7687]), .Z(n4019) );
  XNOR U6701 ( .A(n4020), .B(n4019), .Z(n4119) );
  AND U6702 ( .A(y[7700]), .B(x[487]), .Z(n4118) );
  XOR U6703 ( .A(n4119), .B(n4118), .Z(n4108) );
  AND U6704 ( .A(x[488]), .B(y[7699]), .Z(n4178) );
  AND U6705 ( .A(y[7684]), .B(x[503]), .Z(n4177) );
  XOR U6706 ( .A(n4178), .B(n4177), .Z(n4180) );
  AND U6707 ( .A(x[502]), .B(y[7685]), .Z(n4179) );
  XOR U6708 ( .A(n4180), .B(n4179), .Z(n4107) );
  XOR U6709 ( .A(n4108), .B(n4107), .Z(n4109) );
  XOR U6710 ( .A(n4110), .B(n4109), .Z(n4207) );
  NAND U6711 ( .A(n4022), .B(n4021), .Z(n4026) );
  ANDN U6712 ( .B(n4024), .A(n4023), .Z(n4025) );
  ANDN U6713 ( .B(n4026), .A(n4025), .Z(n4102) );
  NAND U6714 ( .A(n4028), .B(n4027), .Z(n4032) );
  NAND U6715 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U6716 ( .A(n4032), .B(n4031), .Z(n4101) );
  XNOR U6717 ( .A(n4102), .B(n4101), .Z(n4104) );
  AND U6718 ( .A(x[488]), .B(y[7700]), .Z(n4148) );
  NAND U6719 ( .A(n4148), .B(n4033), .Z(n4037) );
  NANDN U6720 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U6721 ( .A(n4037), .B(n4036), .Z(n4163) );
  AND U6722 ( .A(x[494]), .B(y[7693]), .Z(n4195) );
  AND U6723 ( .A(x[481]), .B(y[7706]), .Z(n4194) );
  XOR U6724 ( .A(n4195), .B(n4194), .Z(n4197) );
  AND U6725 ( .A(n4038), .B(o[26]), .Z(n4196) );
  XOR U6726 ( .A(n4197), .B(n4196), .Z(n4162) );
  AND U6727 ( .A(x[497]), .B(y[7690]), .Z(n4129) );
  AND U6728 ( .A(x[484]), .B(y[7703]), .Z(n4128) );
  XOR U6729 ( .A(n4129), .B(n4128), .Z(n4131) );
  AND U6730 ( .A(y[7702]), .B(x[485]), .Z(n4130) );
  XOR U6731 ( .A(n4131), .B(n4130), .Z(n4161) );
  XOR U6732 ( .A(n4162), .B(n4161), .Z(n4164) );
  XOR U6733 ( .A(n4163), .B(n4164), .Z(n4103) );
  XNOR U6734 ( .A(n4104), .B(n4103), .Z(n4206) );
  XOR U6735 ( .A(n4207), .B(n4206), .Z(n4208) );
  XOR U6736 ( .A(n4209), .B(n4208), .Z(n4083) );
  NANDN U6737 ( .A(n4040), .B(n4039), .Z(n4044) );
  NANDN U6738 ( .A(n4042), .B(n4041), .Z(n4043) );
  NAND U6739 ( .A(n4044), .B(n4043), .Z(n4086) );
  NAND U6740 ( .A(n4046), .B(n4045), .Z(n4050) );
  NAND U6741 ( .A(n4048), .B(n4047), .Z(n4049) );
  AND U6742 ( .A(n4050), .B(n4049), .Z(n4071) );
  XNOR U6743 ( .A(n4074), .B(n4073), .Z(n4059) );
  NAND U6744 ( .A(n4052), .B(n4051), .Z(n4056) );
  NAND U6745 ( .A(n4054), .B(n4053), .Z(n4055) );
  AND U6746 ( .A(n4056), .B(n4055), .Z(n4058) );
  XOR U6747 ( .A(n4059), .B(n4058), .Z(n4060) );
  XOR U6748 ( .A(n4061), .B(n4060), .Z(n4067) );
  XNOR U6749 ( .A(n4066), .B(n4067), .Z(n4057) );
  XOR U6750 ( .A(n4064), .B(n4057), .Z(N60) );
  NAND U6751 ( .A(n4059), .B(n4058), .Z(n4063) );
  NAND U6752 ( .A(n4061), .B(n4060), .Z(n4062) );
  NAND U6753 ( .A(n4063), .B(n4062), .Z(n4227) );
  IV U6754 ( .A(n4227), .Z(n4225) );
  OR U6755 ( .A(n4066), .B(n4064), .Z(n4070) );
  ANDN U6756 ( .B(n4066), .A(n4065), .Z(n4068) );
  OR U6757 ( .A(n4068), .B(n4067), .Z(n4069) );
  AND U6758 ( .A(n4070), .B(n4069), .Z(n4226) );
  NANDN U6759 ( .A(n4072), .B(n4071), .Z(n4076) );
  NAND U6760 ( .A(n4074), .B(n4073), .Z(n4075) );
  NAND U6761 ( .A(n4076), .B(n4075), .Z(n4220) );
  NANDN U6762 ( .A(n4078), .B(n4077), .Z(n4082) );
  NAND U6763 ( .A(n4080), .B(n4079), .Z(n4081) );
  NAND U6764 ( .A(n4082), .B(n4081), .Z(n4219) );
  XOR U6765 ( .A(n4220), .B(n4219), .Z(n4222) );
  NANDN U6766 ( .A(n4084), .B(n4083), .Z(n4088) );
  NANDN U6767 ( .A(n4086), .B(n4085), .Z(n4087) );
  AND U6768 ( .A(n4088), .B(n4087), .Z(n4233) );
  NANDN U6769 ( .A(n4090), .B(n4089), .Z(n4094) );
  NANDN U6770 ( .A(n4092), .B(n4091), .Z(n4093) );
  AND U6771 ( .A(n4094), .B(n4093), .Z(n4245) );
  NANDN U6772 ( .A(n4096), .B(n4095), .Z(n4100) );
  OR U6773 ( .A(n4098), .B(n4097), .Z(n4099) );
  NAND U6774 ( .A(n4100), .B(n4099), .Z(n4244) );
  XNOR U6775 ( .A(n4245), .B(n4244), .Z(n4247) );
  NANDN U6776 ( .A(n4102), .B(n4101), .Z(n4106) );
  NAND U6777 ( .A(n4104), .B(n4103), .Z(n4105) );
  NAND U6778 ( .A(n4106), .B(n4105), .Z(n4348) );
  NAND U6779 ( .A(n4112), .B(n4111), .Z(n4116) );
  NANDN U6780 ( .A(n4114), .B(n4113), .Z(n4115) );
  NAND U6781 ( .A(n4116), .B(n4115), .Z(n4346) );
  XOR U6782 ( .A(n4347), .B(n4346), .Z(n4349) );
  XOR U6783 ( .A(n4348), .B(n4349), .Z(n4248) );
  AND U6784 ( .A(y[7687]), .B(x[504]), .Z(n4728) );
  NAND U6785 ( .A(n4728), .B(n4117), .Z(n4121) );
  NAND U6786 ( .A(n4119), .B(n4118), .Z(n4120) );
  NAND U6787 ( .A(n4121), .B(n4120), .Z(n4384) );
  AND U6788 ( .A(x[505]), .B(y[7683]), .Z(n4297) );
  XOR U6789 ( .A(n4298), .B(n4297), .Z(n4296) );
  AND U6790 ( .A(x[481]), .B(y[7707]), .Z(n4295) );
  XOR U6791 ( .A(n4296), .B(n4295), .Z(n4383) );
  AND U6792 ( .A(y[7692]), .B(x[496]), .Z(n4290) );
  AND U6793 ( .A(x[504]), .B(y[7684]), .Z(n4289) );
  XOR U6794 ( .A(n4290), .B(n4289), .Z(n4292) );
  AND U6795 ( .A(x[482]), .B(y[7706]), .Z(n4291) );
  XOR U6796 ( .A(n4292), .B(n4291), .Z(n4382) );
  XOR U6797 ( .A(n4383), .B(n4382), .Z(n4385) );
  XOR U6798 ( .A(n4384), .B(n4385), .Z(n4355) );
  NAND U6799 ( .A(n4123), .B(n4122), .Z(n4127) );
  NAND U6800 ( .A(n4125), .B(n4124), .Z(n4126) );
  NAND U6801 ( .A(n4127), .B(n4126), .Z(n4378) );
  AND U6802 ( .A(y[7705]), .B(x[483]), .Z(n4326) );
  XOR U6803 ( .A(n4327), .B(n4326), .Z(n4329) );
  AND U6804 ( .A(x[503]), .B(y[7685]), .Z(n4328) );
  XOR U6805 ( .A(n4329), .B(n4328), .Z(n4377) );
  AND U6806 ( .A(y[7703]), .B(x[485]), .Z(n4313) );
  AND U6807 ( .A(y[7687]), .B(x[501]), .Z(n4312) );
  XOR U6808 ( .A(n4313), .B(n4312), .Z(n4315) );
  AND U6809 ( .A(y[7688]), .B(x[500]), .Z(n4314) );
  XOR U6810 ( .A(n4315), .B(n4314), .Z(n4376) );
  XOR U6811 ( .A(n4377), .B(n4376), .Z(n4379) );
  XOR U6812 ( .A(n4378), .B(n4379), .Z(n4353) );
  NAND U6813 ( .A(n4129), .B(n4128), .Z(n4133) );
  NAND U6814 ( .A(n4131), .B(n4130), .Z(n4132) );
  NAND U6815 ( .A(n4133), .B(n4132), .Z(n4371) );
  NAND U6816 ( .A(n4135), .B(n4134), .Z(n4139) );
  NAND U6817 ( .A(n4137), .B(n4136), .Z(n4138) );
  NAND U6818 ( .A(n4139), .B(n4138), .Z(n4370) );
  XOR U6819 ( .A(n4371), .B(n4370), .Z(n4373) );
  NAND U6820 ( .A(n4141), .B(n4140), .Z(n4145) );
  NAND U6821 ( .A(n4143), .B(n4142), .Z(n4144) );
  NAND U6822 ( .A(n4145), .B(n4144), .Z(n4285) );
  AND U6823 ( .A(x[480]), .B(y[7708]), .Z(n4273) );
  AND U6824 ( .A(x[508]), .B(y[7680]), .Z(n4272) );
  XOR U6825 ( .A(n4273), .B(n4272), .Z(n4275) );
  AND U6826 ( .A(n4146), .B(o[27]), .Z(n4274) );
  XOR U6827 ( .A(n4275), .B(n4274), .Z(n4284) );
  NAND U6828 ( .A(y[7698]), .B(x[490]), .Z(n4147) );
  XNOR U6829 ( .A(n4148), .B(n4147), .Z(n4280) );
  AND U6830 ( .A(x[489]), .B(y[7699]), .Z(n4279) );
  XOR U6831 ( .A(n4280), .B(n4279), .Z(n4283) );
  XOR U6832 ( .A(n4284), .B(n4283), .Z(n4286) );
  XOR U6833 ( .A(n4285), .B(n4286), .Z(n4372) );
  XNOR U6834 ( .A(n4373), .B(n4372), .Z(n4352) );
  NAND U6835 ( .A(n4150), .B(n4149), .Z(n4154) );
  NANDN U6836 ( .A(n4152), .B(n4151), .Z(n4153) );
  NAND U6837 ( .A(n4154), .B(n4153), .Z(n4254) );
  NAND U6838 ( .A(n4156), .B(n4155), .Z(n4160) );
  NANDN U6839 ( .A(n4158), .B(n4157), .Z(n4159) );
  NAND U6840 ( .A(n4160), .B(n4159), .Z(n4360) );
  NAND U6841 ( .A(n4162), .B(n4161), .Z(n4166) );
  NAND U6842 ( .A(n4164), .B(n4163), .Z(n4165) );
  NAND U6843 ( .A(n4166), .B(n4165), .Z(n4359) );
  NAND U6844 ( .A(n4168), .B(n4167), .Z(n4172) );
  NAND U6845 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U6846 ( .A(n4172), .B(n4171), .Z(n4358) );
  XOR U6847 ( .A(n4359), .B(n4358), .Z(n4361) );
  XOR U6848 ( .A(n4360), .B(n4361), .Z(n4255) );
  XOR U6849 ( .A(n4254), .B(n4255), .Z(n4257) );
  AND U6850 ( .A(x[487]), .B(y[7701]), .Z(n4302) );
  AND U6851 ( .A(x[492]), .B(y[7696]), .Z(n4301) );
  XOR U6852 ( .A(n4302), .B(n4301), .Z(n4304) );
  AND U6853 ( .A(y[7697]), .B(x[491]), .Z(n4303) );
  XOR U6854 ( .A(n4304), .B(n4303), .Z(n4321) );
  AND U6855 ( .A(x[495]), .B(y[7693]), .Z(n4335) );
  AND U6856 ( .A(y[7681]), .B(x[507]), .Z(n4318) );
  XOR U6857 ( .A(o[28]), .B(n4318), .Z(n4333) );
  AND U6858 ( .A(x[506]), .B(y[7682]), .Z(n4332) );
  XOR U6859 ( .A(n4333), .B(n4332), .Z(n4334) );
  XNOR U6860 ( .A(n4335), .B(n4334), .Z(n4320) );
  XOR U6861 ( .A(n4322), .B(n4323), .Z(n4365) );
  NAND U6862 ( .A(n4178), .B(n4177), .Z(n4182) );
  NAND U6863 ( .A(n4180), .B(n4179), .Z(n4181) );
  NAND U6864 ( .A(n4182), .B(n4181), .Z(n4342) );
  AND U6865 ( .A(x[497]), .B(y[7691]), .Z(n4267) );
  AND U6866 ( .A(x[502]), .B(y[7686]), .Z(n4266) );
  XOR U6867 ( .A(n4267), .B(n4266), .Z(n4269) );
  AND U6868 ( .A(x[484]), .B(y[7704]), .Z(n4268) );
  XOR U6869 ( .A(n4269), .B(n4268), .Z(n4341) );
  AND U6870 ( .A(x[486]), .B(y[7702]), .Z(n4510) );
  AND U6871 ( .A(y[7689]), .B(x[499]), .Z(n4307) );
  XOR U6872 ( .A(n4510), .B(n4307), .Z(n4309) );
  XOR U6873 ( .A(n4309), .B(n4308), .Z(n4340) );
  XOR U6874 ( .A(n4341), .B(n4340), .Z(n4343) );
  XOR U6875 ( .A(n4342), .B(n4343), .Z(n4364) );
  NAND U6876 ( .A(n4327), .B(n4183), .Z(n4187) );
  NANDN U6877 ( .A(n4185), .B(n4184), .Z(n4186) );
  NAND U6878 ( .A(n4187), .B(n4186), .Z(n4262) );
  NAND U6879 ( .A(n4189), .B(n4188), .Z(n4193) );
  NAND U6880 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U6881 ( .A(n4193), .B(n4192), .Z(n4261) );
  NAND U6882 ( .A(n4195), .B(n4194), .Z(n4199) );
  NAND U6883 ( .A(n4197), .B(n4196), .Z(n4198) );
  NAND U6884 ( .A(n4199), .B(n4198), .Z(n4260) );
  XNOR U6885 ( .A(n4261), .B(n4260), .Z(n4263) );
  XNOR U6886 ( .A(n4366), .B(n4367), .Z(n4256) );
  XOR U6887 ( .A(n4257), .B(n4256), .Z(n4250) );
  XOR U6888 ( .A(n4251), .B(n4250), .Z(n4246) );
  XOR U6889 ( .A(n4247), .B(n4246), .Z(n4232) );
  XOR U6890 ( .A(n4233), .B(n4232), .Z(n4235) );
  NANDN U6891 ( .A(n4201), .B(n4200), .Z(n4205) );
  NANDN U6892 ( .A(n4203), .B(n4202), .Z(n4204) );
  AND U6893 ( .A(n4205), .B(n4204), .Z(n4241) );
  NAND U6894 ( .A(n4207), .B(n4206), .Z(n4211) );
  NAND U6895 ( .A(n4209), .B(n4208), .Z(n4210) );
  AND U6896 ( .A(n4211), .B(n4210), .Z(n4238) );
  NANDN U6897 ( .A(n4213), .B(n4212), .Z(n4217) );
  NANDN U6898 ( .A(n4215), .B(n4214), .Z(n4216) );
  NAND U6899 ( .A(n4217), .B(n4216), .Z(n4239) );
  XOR U6900 ( .A(n4235), .B(n4234), .Z(n4221) );
  XOR U6901 ( .A(n4222), .B(n4221), .Z(n4228) );
  XNOR U6902 ( .A(n4226), .B(n4228), .Z(n4218) );
  XOR U6903 ( .A(n4225), .B(n4218), .Z(N61) );
  NAND U6904 ( .A(n4220), .B(n4219), .Z(n4224) );
  NAND U6905 ( .A(n4222), .B(n4221), .Z(n4223) );
  AND U6906 ( .A(n4224), .B(n4223), .Z(n4553) );
  NANDN U6907 ( .A(n4225), .B(n4226), .Z(n4231) );
  NOR U6908 ( .A(n4227), .B(n4226), .Z(n4229) );
  OR U6909 ( .A(n4229), .B(n4228), .Z(n4230) );
  AND U6910 ( .A(n4231), .B(n4230), .Z(n4554) );
  NAND U6911 ( .A(n4233), .B(n4232), .Z(n4237) );
  NAND U6912 ( .A(n4235), .B(n4234), .Z(n4236) );
  AND U6913 ( .A(n4237), .B(n4236), .Z(n4559) );
  NANDN U6914 ( .A(n4239), .B(n4238), .Z(n4243) );
  NANDN U6915 ( .A(n4241), .B(n4240), .Z(n4242) );
  AND U6916 ( .A(n4243), .B(n4242), .Z(n4557) );
  NANDN U6917 ( .A(n4249), .B(n4248), .Z(n4253) );
  NAND U6918 ( .A(n4251), .B(n4250), .Z(n4252) );
  NAND U6919 ( .A(n4253), .B(n4252), .Z(n4390) );
  XOR U6920 ( .A(n4389), .B(n4390), .Z(n4392) );
  NAND U6921 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U6922 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U6923 ( .A(n4259), .B(n4258), .Z(n4541) );
  NAND U6924 ( .A(n4261), .B(n4260), .Z(n4265) );
  NANDN U6925 ( .A(n4263), .B(n4262), .Z(n4264) );
  AND U6926 ( .A(n4265), .B(n4264), .Z(n4395) );
  NAND U6927 ( .A(n4267), .B(n4266), .Z(n4271) );
  NAND U6928 ( .A(n4269), .B(n4268), .Z(n4270) );
  NAND U6929 ( .A(n4271), .B(n4270), .Z(n4433) );
  NAND U6930 ( .A(n4273), .B(n4272), .Z(n4277) );
  NAND U6931 ( .A(n4275), .B(n4274), .Z(n4276) );
  NAND U6932 ( .A(n4277), .B(n4276), .Z(n4432) );
  XOR U6933 ( .A(n4433), .B(n4432), .Z(n4434) );
  AND U6934 ( .A(y[7700]), .B(x[490]), .Z(n4430) );
  NAND U6935 ( .A(n4430), .B(n4278), .Z(n4282) );
  NAND U6936 ( .A(n4280), .B(n4279), .Z(n4281) );
  NAND U6937 ( .A(n4282), .B(n4281), .Z(n4401) );
  AND U6938 ( .A(x[502]), .B(y[7687]), .Z(n4488) );
  AND U6939 ( .A(x[492]), .B(y[7697]), .Z(n4617) );
  AND U6940 ( .A(y[7708]), .B(x[481]), .Z(n4486) );
  XOR U6941 ( .A(n4617), .B(n4486), .Z(n4487) );
  XOR U6942 ( .A(n4488), .B(n4487), .Z(n4400) );
  AND U6943 ( .A(x[495]), .B(y[7694]), .Z(n4491) );
  XOR U6944 ( .A(n4491), .B(n4612), .Z(n4493) );
  XOR U6945 ( .A(n4493), .B(n4492), .Z(n4399) );
  XOR U6946 ( .A(n4400), .B(n4399), .Z(n4402) );
  XNOR U6947 ( .A(n4401), .B(n4402), .Z(n4435) );
  NAND U6948 ( .A(n4284), .B(n4283), .Z(n4288) );
  NAND U6949 ( .A(n4286), .B(n4285), .Z(n4287) );
  AND U6950 ( .A(n4288), .B(n4287), .Z(n4393) );
  XNOR U6951 ( .A(n4395), .B(n4396), .Z(n4441) );
  NAND U6952 ( .A(n4290), .B(n4289), .Z(n4294) );
  NAND U6953 ( .A(n4292), .B(n4291), .Z(n4293) );
  NAND U6954 ( .A(n4294), .B(n4293), .Z(n4406) );
  AND U6955 ( .A(n4296), .B(n4295), .Z(n4300) );
  NAND U6956 ( .A(n4298), .B(n4297), .Z(n4299) );
  NANDN U6957 ( .A(n4300), .B(n4299), .Z(n4405) );
  XOR U6958 ( .A(n4406), .B(n4405), .Z(n4407) );
  NAND U6959 ( .A(n4302), .B(n4301), .Z(n4306) );
  NAND U6960 ( .A(n4304), .B(n4303), .Z(n4305) );
  NAND U6961 ( .A(n4306), .B(n4305), .Z(n4452) );
  AND U6962 ( .A(y[7698]), .B(x[491]), .Z(n4507) );
  AND U6963 ( .A(x[483]), .B(y[7706]), .Z(n4505) );
  AND U6964 ( .A(x[497]), .B(y[7692]), .Z(n4504) );
  XOR U6965 ( .A(n4505), .B(n4504), .Z(n4506) );
  XOR U6966 ( .A(n4507), .B(n4506), .Z(n4451) );
  AND U6967 ( .A(y[7686]), .B(x[503]), .Z(n4501) );
  AND U6968 ( .A(x[493]), .B(y[7696]), .Z(n4499) );
  AND U6969 ( .A(x[504]), .B(y[7685]), .Z(n4626) );
  XOR U6970 ( .A(n4499), .B(n4626), .Z(n4500) );
  XOR U6971 ( .A(n4501), .B(n4500), .Z(n4450) );
  XOR U6972 ( .A(n4451), .B(n4450), .Z(n4453) );
  XNOR U6973 ( .A(n4452), .B(n4453), .Z(n4408) );
  IV U6974 ( .A(n4532), .Z(n4319) );
  NAND U6975 ( .A(n4510), .B(n4307), .Z(n4311) );
  NAND U6976 ( .A(n4309), .B(n4308), .Z(n4310) );
  AND U6977 ( .A(n4311), .B(n4310), .Z(n4413) );
  AND U6978 ( .A(x[505]), .B(y[7684]), .Z(n4483) );
  AND U6979 ( .A(x[506]), .B(y[7683]), .Z(n4480) );
  XOR U6980 ( .A(n4481), .B(n4480), .Z(n4482) );
  XOR U6981 ( .A(n4483), .B(n4482), .Z(n4412) );
  AND U6982 ( .A(x[508]), .B(y[7681]), .Z(n4498) );
  XOR U6983 ( .A(o[29]), .B(n4498), .Z(n4425) );
  AND U6984 ( .A(x[480]), .B(y[7709]), .Z(n4423) );
  AND U6985 ( .A(y[7680]), .B(x[509]), .Z(n4422) );
  XOR U6986 ( .A(n4423), .B(n4422), .Z(n4424) );
  XNOR U6987 ( .A(n4425), .B(n4424), .Z(n4411) );
  XNOR U6988 ( .A(n4413), .B(n4414), .Z(n4529) );
  NAND U6989 ( .A(n4313), .B(n4312), .Z(n4317) );
  NAND U6990 ( .A(n4315), .B(n4314), .Z(n4316) );
  NAND U6991 ( .A(n4317), .B(n4316), .Z(n4519) );
  AND U6992 ( .A(n4318), .B(o[28]), .Z(n4471) );
  AND U6993 ( .A(y[7693]), .B(x[496]), .Z(n4469) );
  AND U6994 ( .A(x[507]), .B(y[7682]), .Z(n4468) );
  XOR U6995 ( .A(n4469), .B(n4468), .Z(n4470) );
  XOR U6996 ( .A(n4471), .B(n4470), .Z(n4518) );
  AND U6997 ( .A(x[482]), .B(y[7707]), .Z(n4463) );
  XOR U6998 ( .A(n4463), .B(n4462), .Z(n4464) );
  XOR U6999 ( .A(n4465), .B(n4464), .Z(n4517) );
  XOR U7000 ( .A(n4518), .B(n4517), .Z(n4520) );
  XOR U7001 ( .A(n4519), .B(n4520), .Z(n4530) );
  XOR U7002 ( .A(n4319), .B(n4531), .Z(n4446) );
  NANDN U7003 ( .A(n4321), .B(n4320), .Z(n4325) );
  NAND U7004 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U7005 ( .A(n4325), .B(n4324), .Z(n4444) );
  NAND U7006 ( .A(n4327), .B(n4326), .Z(n4331) );
  NAND U7007 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U7008 ( .A(n4331), .B(n4330), .Z(n4475) );
  NAND U7009 ( .A(n4333), .B(n4332), .Z(n4337) );
  NAND U7010 ( .A(n4335), .B(n4334), .Z(n4336) );
  NAND U7011 ( .A(n4337), .B(n4336), .Z(n4474) );
  XOR U7012 ( .A(n4475), .B(n4474), .Z(n4477) );
  AND U7013 ( .A(y[7704]), .B(x[485]), .Z(n4459) );
  AND U7014 ( .A(x[484]), .B(y[7705]), .Z(n4457) );
  AND U7015 ( .A(x[490]), .B(y[7699]), .Z(n4456) );
  XOR U7016 ( .A(n4457), .B(n4456), .Z(n4458) );
  XOR U7017 ( .A(n4459), .B(n4458), .Z(n4419) );
  AND U7018 ( .A(x[488]), .B(y[7701]), .Z(n4512) );
  AND U7019 ( .A(y[7703]), .B(x[486]), .Z(n4339) );
  AND U7020 ( .A(y[7702]), .B(x[487]), .Z(n4338) );
  XOR U7021 ( .A(n4339), .B(n4338), .Z(n4511) );
  XOR U7022 ( .A(n4512), .B(n4511), .Z(n4417) );
  AND U7023 ( .A(y[7700]), .B(x[489]), .Z(n4701) );
  XOR U7024 ( .A(n4417), .B(n4701), .Z(n4418) );
  XOR U7025 ( .A(n4419), .B(n4418), .Z(n4476) );
  XOR U7026 ( .A(n4477), .B(n4476), .Z(n4445) );
  XNOR U7027 ( .A(n4446), .B(n4447), .Z(n4439) );
  NAND U7028 ( .A(n4341), .B(n4340), .Z(n4345) );
  NAND U7029 ( .A(n4343), .B(n4342), .Z(n4344) );
  NAND U7030 ( .A(n4345), .B(n4344), .Z(n4438) );
  XOR U7031 ( .A(n4541), .B(n4542), .Z(n4544) );
  NAND U7032 ( .A(n4347), .B(n4346), .Z(n4351) );
  NAND U7033 ( .A(n4349), .B(n4348), .Z(n4350) );
  NAND U7034 ( .A(n4351), .B(n4350), .Z(n4535) );
  NANDN U7035 ( .A(n4353), .B(n4352), .Z(n4357) );
  NANDN U7036 ( .A(n4355), .B(n4354), .Z(n4356) );
  AND U7037 ( .A(n4357), .B(n4356), .Z(n4536) );
  XOR U7038 ( .A(n4535), .B(n4536), .Z(n4537) );
  NAND U7039 ( .A(n4359), .B(n4358), .Z(n4363) );
  NAND U7040 ( .A(n4361), .B(n4360), .Z(n4362) );
  NAND U7041 ( .A(n4363), .B(n4362), .Z(n4549) );
  NANDN U7042 ( .A(n4365), .B(n4364), .Z(n4369) );
  NANDN U7043 ( .A(n4367), .B(n4366), .Z(n4368) );
  NAND U7044 ( .A(n4369), .B(n4368), .Z(n4547) );
  NAND U7045 ( .A(n4371), .B(n4370), .Z(n4375) );
  NAND U7046 ( .A(n4373), .B(n4372), .Z(n4374) );
  NAND U7047 ( .A(n4375), .B(n4374), .Z(n4525) );
  NAND U7048 ( .A(n4377), .B(n4376), .Z(n4381) );
  NAND U7049 ( .A(n4379), .B(n4378), .Z(n4380) );
  NAND U7050 ( .A(n4381), .B(n4380), .Z(n4524) );
  NAND U7051 ( .A(n4383), .B(n4382), .Z(n4387) );
  NAND U7052 ( .A(n4385), .B(n4384), .Z(n4386) );
  NAND U7053 ( .A(n4387), .B(n4386), .Z(n4523) );
  XNOR U7054 ( .A(n4524), .B(n4523), .Z(n4526) );
  XOR U7055 ( .A(n4547), .B(n4548), .Z(n4550) );
  XOR U7056 ( .A(n4549), .B(n4550), .Z(n4538) );
  XNOR U7057 ( .A(n4537), .B(n4538), .Z(n4543) );
  XOR U7058 ( .A(n4544), .B(n4543), .Z(n4391) );
  XOR U7059 ( .A(n4392), .B(n4391), .Z(n4556) );
  XNOR U7060 ( .A(n4554), .B(n4555), .Z(n4388) );
  XOR U7061 ( .A(n4553), .B(n4388), .Z(N62) );
  NANDN U7062 ( .A(n4394), .B(n4393), .Z(n4398) );
  NANDN U7063 ( .A(n4396), .B(n4395), .Z(n4397) );
  AND U7064 ( .A(n4398), .B(n4397), .Z(n4813) );
  NAND U7065 ( .A(n4400), .B(n4399), .Z(n4404) );
  NAND U7066 ( .A(n4402), .B(n4401), .Z(n4403) );
  AND U7067 ( .A(n4404), .B(n4403), .Z(n4794) );
  NAND U7068 ( .A(n4406), .B(n4405), .Z(n4410) );
  NANDN U7069 ( .A(n4408), .B(n4407), .Z(n4409) );
  NAND U7070 ( .A(n4410), .B(n4409), .Z(n4795) );
  NANDN U7071 ( .A(n4412), .B(n4411), .Z(n4416) );
  NANDN U7072 ( .A(n4414), .B(n4413), .Z(n4415) );
  NAND U7073 ( .A(n4416), .B(n4415), .Z(n4792) );
  XOR U7074 ( .A(n4793), .B(n4792), .Z(n4810) );
  NAND U7075 ( .A(n4417), .B(n4701), .Z(n4421) );
  NAND U7076 ( .A(n4419), .B(n4418), .Z(n4420) );
  AND U7077 ( .A(n4421), .B(n4420), .Z(n4577) );
  NAND U7078 ( .A(n4423), .B(n4422), .Z(n4427) );
  NAND U7079 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U7080 ( .A(n4427), .B(n4426), .Z(n4580) );
  AND U7081 ( .A(x[492]), .B(y[7698]), .Z(n4428) );
  XOR U7082 ( .A(n4429), .B(n4428), .Z(n4618) );
  XOR U7083 ( .A(n4619), .B(n4618), .Z(n4700) );
  AND U7084 ( .A(y[7701]), .B(x[489]), .Z(n4431) );
  XOR U7085 ( .A(n4431), .B(n4430), .Z(n4699) );
  XOR U7086 ( .A(n4700), .B(n4699), .Z(n4583) );
  AND U7087 ( .A(y[7683]), .B(x[507]), .Z(n4668) );
  AND U7088 ( .A(x[481]), .B(y[7709]), .Z(n4667) );
  XOR U7089 ( .A(n4668), .B(n4667), .Z(n4669) );
  XOR U7090 ( .A(n4670), .B(n4669), .Z(n4582) );
  XOR U7091 ( .A(n4583), .B(n4582), .Z(n4581) );
  XNOR U7092 ( .A(n4580), .B(n4581), .Z(n4576) );
  XOR U7093 ( .A(n4577), .B(n4576), .Z(n4575) );
  NAND U7094 ( .A(n4433), .B(n4432), .Z(n4437) );
  NANDN U7095 ( .A(n4435), .B(n4434), .Z(n4436) );
  AND U7096 ( .A(n4437), .B(n4436), .Z(n4574) );
  XNOR U7097 ( .A(n4575), .B(n4574), .Z(n4811) );
  XOR U7098 ( .A(n4813), .B(n4812), .Z(n4855) );
  NANDN U7099 ( .A(n4439), .B(n4438), .Z(n4443) );
  NANDN U7100 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U7101 ( .A(n4443), .B(n4442), .Z(n4857) );
  NANDN U7102 ( .A(n4445), .B(n4444), .Z(n4449) );
  NANDN U7103 ( .A(n4447), .B(n4446), .Z(n4448) );
  AND U7104 ( .A(n4449), .B(n4448), .Z(n4837) );
  NAND U7105 ( .A(n4451), .B(n4450), .Z(n4455) );
  NAND U7106 ( .A(n4453), .B(n4452), .Z(n4454) );
  AND U7107 ( .A(n4455), .B(n4454), .Z(n4807) );
  NAND U7108 ( .A(n4457), .B(n4456), .Z(n4461) );
  NAND U7109 ( .A(n4459), .B(n4458), .Z(n4460) );
  AND U7110 ( .A(n4461), .B(n4460), .Z(n4772) );
  AND U7111 ( .A(y[7704]), .B(x[486]), .Z(n4664) );
  AND U7112 ( .A(y[7705]), .B(x[485]), .Z(n4662) );
  AND U7113 ( .A(y[7691]), .B(x[499]), .Z(n4661) );
  XOR U7114 ( .A(n4662), .B(n4661), .Z(n4663) );
  XNOR U7115 ( .A(n4664), .B(n4663), .Z(n4600) );
  AND U7116 ( .A(x[484]), .B(y[7706]), .Z(n4636) );
  AND U7117 ( .A(x[483]), .B(y[7707]), .Z(n4638) );
  AND U7118 ( .A(x[498]), .B(y[7692]), .Z(n4637) );
  XOR U7119 ( .A(n4638), .B(n4637), .Z(n4635) );
  XOR U7120 ( .A(n4636), .B(n4635), .Z(n4603) );
  NAND U7121 ( .A(n4463), .B(n4462), .Z(n4467) );
  NAND U7122 ( .A(n4465), .B(n4464), .Z(n4466) );
  AND U7123 ( .A(n4467), .B(n4466), .Z(n4602) );
  XOR U7124 ( .A(n4600), .B(n4601), .Z(n4773) );
  XNOR U7125 ( .A(n4772), .B(n4773), .Z(n4771) );
  NAND U7126 ( .A(n4469), .B(n4468), .Z(n4473) );
  NAND U7127 ( .A(n4471), .B(n4470), .Z(n4472) );
  AND U7128 ( .A(n4473), .B(n4472), .Z(n4770) );
  XOR U7129 ( .A(n4771), .B(n4770), .Z(n4806) );
  XOR U7130 ( .A(n4807), .B(n4806), .Z(n4805) );
  NAND U7131 ( .A(n4475), .B(n4474), .Z(n4479) );
  NAND U7132 ( .A(n4477), .B(n4476), .Z(n4478) );
  AND U7133 ( .A(n4479), .B(n4478), .Z(n4804) );
  XOR U7134 ( .A(n4805), .B(n4804), .Z(n4839) );
  AND U7135 ( .A(n4481), .B(n4480), .Z(n4485) );
  NAND U7136 ( .A(n4483), .B(n4482), .Z(n4484) );
  NANDN U7137 ( .A(n4485), .B(n4484), .Z(n4764) );
  AND U7138 ( .A(n4617), .B(n4486), .Z(n4490) );
  NAND U7139 ( .A(n4488), .B(n4487), .Z(n4489) );
  NANDN U7140 ( .A(n4490), .B(n4489), .Z(n4767) );
  NAND U7141 ( .A(n4491), .B(n4612), .Z(n4495) );
  NAND U7142 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U7143 ( .A(n4495), .B(n4494), .Z(n4593) );
  AND U7144 ( .A(y[7687]), .B(x[503]), .Z(n4625) );
  AND U7145 ( .A(y[7685]), .B(x[505]), .Z(n4497) );
  AND U7146 ( .A(x[504]), .B(y[7686]), .Z(n4496) );
  XOR U7147 ( .A(n4497), .B(n4496), .Z(n4624) );
  XOR U7148 ( .A(n4625), .B(n4624), .Z(n4595) );
  AND U7149 ( .A(n4498), .B(o[29]), .Z(n4692) );
  AND U7150 ( .A(x[508]), .B(y[7682]), .Z(n4694) );
  AND U7151 ( .A(y[7694]), .B(x[496]), .Z(n4693) );
  XOR U7152 ( .A(n4694), .B(n4693), .Z(n4691) );
  XNOR U7153 ( .A(n4692), .B(n4691), .Z(n4594) );
  XNOR U7154 ( .A(n4593), .B(n4592), .Z(n4766) );
  XOR U7155 ( .A(n4767), .B(n4766), .Z(n4765) );
  XOR U7156 ( .A(n4764), .B(n4765), .Z(n4819) );
  NAND U7157 ( .A(n4499), .B(n4626), .Z(n4503) );
  NAND U7158 ( .A(n4501), .B(n4500), .Z(n4502) );
  NAND U7159 ( .A(n4503), .B(n4502), .Z(n4789) );
  NAND U7160 ( .A(n4505), .B(n4504), .Z(n4509) );
  NAND U7161 ( .A(n4507), .B(n4506), .Z(n4508) );
  AND U7162 ( .A(n4509), .B(n4508), .Z(n4607) );
  AND U7163 ( .A(x[480]), .B(y[7710]), .Z(n4680) );
  AND U7164 ( .A(y[7681]), .B(x[509]), .Z(n4704) );
  XOR U7165 ( .A(o[30]), .B(n4704), .Z(n4682) );
  AND U7166 ( .A(y[7680]), .B(x[510]), .Z(n4681) );
  XOR U7167 ( .A(n4682), .B(n4681), .Z(n4679) );
  XOR U7168 ( .A(n4680), .B(n4679), .Z(n4609) );
  AND U7169 ( .A(x[500]), .B(y[7690]), .Z(n4631) );
  XOR U7170 ( .A(n4632), .B(n4631), .Z(n4630) );
  AND U7171 ( .A(x[488]), .B(y[7702]), .Z(n4629) );
  XNOR U7172 ( .A(n4630), .B(n4629), .Z(n4608) );
  XNOR U7173 ( .A(n4607), .B(n4606), .Z(n4788) );
  XOR U7174 ( .A(n4789), .B(n4788), .Z(n4786) );
  AND U7175 ( .A(x[487]), .B(y[7703]), .Z(n4614) );
  NAND U7176 ( .A(n4510), .B(n4614), .Z(n4514) );
  NAND U7177 ( .A(n4512), .B(n4511), .Z(n4513) );
  AND U7178 ( .A(n4514), .B(n4513), .Z(n4586) );
  AND U7179 ( .A(y[7689]), .B(x[501]), .Z(n4516) );
  AND U7180 ( .A(y[7688]), .B(x[502]), .Z(n4515) );
  XOR U7181 ( .A(n4516), .B(n4515), .Z(n4613) );
  XOR U7182 ( .A(n4614), .B(n4613), .Z(n4589) );
  AND U7183 ( .A(x[497]), .B(y[7693]), .Z(n4686) );
  AND U7184 ( .A(y[7708]), .B(x[482]), .Z(n4688) );
  AND U7185 ( .A(x[506]), .B(y[7684]), .Z(n4687) );
  XOR U7186 ( .A(n4688), .B(n4687), .Z(n4685) );
  XNOR U7187 ( .A(n4686), .B(n4685), .Z(n4588) );
  XNOR U7188 ( .A(n4586), .B(n4587), .Z(n4787) );
  NAND U7189 ( .A(n4518), .B(n4517), .Z(n4522) );
  NAND U7190 ( .A(n4520), .B(n4519), .Z(n4521) );
  NAND U7191 ( .A(n4522), .B(n4521), .Z(n4820) );
  XOR U7192 ( .A(n4821), .B(n4820), .Z(n4818) );
  XOR U7193 ( .A(n4819), .B(n4818), .Z(n4838) );
  XOR U7194 ( .A(n4837), .B(n4836), .Z(n4570) );
  NAND U7195 ( .A(n4524), .B(n4523), .Z(n4528) );
  NANDN U7196 ( .A(n4526), .B(n4525), .Z(n4527) );
  AND U7197 ( .A(n4528), .B(n4527), .Z(n4571) );
  NANDN U7198 ( .A(n4530), .B(n4529), .Z(n4534) );
  NANDN U7199 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U7200 ( .A(n4534), .B(n4533), .Z(n4568) );
  XOR U7201 ( .A(n4569), .B(n4568), .Z(n4856) );
  XOR U7202 ( .A(n4857), .B(n4856), .Z(n4854) );
  NAND U7203 ( .A(n4536), .B(n4535), .Z(n4540) );
  NANDN U7204 ( .A(n4538), .B(n4537), .Z(n4539) );
  AND U7205 ( .A(n4540), .B(n4539), .Z(n4832) );
  NAND U7206 ( .A(n4542), .B(n4541), .Z(n4546) );
  NAND U7207 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U7208 ( .A(n4546), .B(n4545), .Z(n4833) );
  NANDN U7209 ( .A(n4548), .B(n4547), .Z(n4552) );
  NANDN U7210 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U7211 ( .A(n4552), .B(n4551), .Z(n4831) );
  XOR U7212 ( .A(n4851), .B(n4850), .Z(n4848) );
  XOR U7213 ( .A(n4849), .B(n4848), .Z(n4563) );
  NANDN U7214 ( .A(n4557), .B(n4556), .Z(n4561) );
  NANDN U7215 ( .A(n4559), .B(n4558), .Z(n4560) );
  AND U7216 ( .A(n4561), .B(n4560), .Z(n4565) );
  XNOR U7217 ( .A(n4564), .B(n4565), .Z(n4562) );
  XNOR U7218 ( .A(n4563), .B(n4562), .Z(N63) );
  NAND U7219 ( .A(n4563), .B(n4562), .Z(n4567) );
  ANDN U7220 ( .B(n4565), .A(n4564), .Z(n4566) );
  ANDN U7221 ( .B(n4567), .A(n4566), .Z(n4847) );
  NAND U7222 ( .A(n4569), .B(n4568), .Z(n4573) );
  ANDN U7223 ( .B(n4571), .A(n4570), .Z(n4572) );
  ANDN U7224 ( .B(n4573), .A(n4572), .Z(n4829) );
  NAND U7225 ( .A(n4575), .B(n4574), .Z(n4579) );
  NAND U7226 ( .A(n4577), .B(n4576), .Z(n4578) );
  AND U7227 ( .A(n4579), .B(n4578), .Z(n4803) );
  NAND U7228 ( .A(n4581), .B(n4580), .Z(n4585) );
  NAND U7229 ( .A(n4583), .B(n4582), .Z(n4584) );
  AND U7230 ( .A(n4585), .B(n4584), .Z(n4785) );
  NANDN U7231 ( .A(n4587), .B(n4586), .Z(n4591) );
  NANDN U7232 ( .A(n4589), .B(n4588), .Z(n4590) );
  AND U7233 ( .A(n4591), .B(n4590), .Z(n4599) );
  NAND U7234 ( .A(n4593), .B(n4592), .Z(n4597) );
  NANDN U7235 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U7236 ( .A(n4597), .B(n4596), .Z(n4598) );
  XNOR U7237 ( .A(n4599), .B(n4598), .Z(n4783) );
  NANDN U7238 ( .A(n4601), .B(n4600), .Z(n4605) );
  NANDN U7239 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U7240 ( .A(n4605), .B(n4604), .Z(n4781) );
  NAND U7241 ( .A(n4607), .B(n4606), .Z(n4611) );
  NANDN U7242 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U7243 ( .A(n4611), .B(n4610), .Z(n4763) );
  AND U7244 ( .A(x[502]), .B(y[7689]), .Z(n4729) );
  AND U7245 ( .A(n4612), .B(n4729), .Z(n4616) );
  AND U7246 ( .A(n4614), .B(n4613), .Z(n4615) );
  NOR U7247 ( .A(n4616), .B(n4615), .Z(n4623) );
  NAND U7248 ( .A(n4617), .B(n4707), .Z(n4621) );
  NAND U7249 ( .A(n4619), .B(n4618), .Z(n4620) );
  AND U7250 ( .A(n4621), .B(n4620), .Z(n4622) );
  XNOR U7251 ( .A(n4623), .B(n4622), .Z(n4678) );
  NAND U7252 ( .A(n4625), .B(n4624), .Z(n4628) );
  AND U7253 ( .A(y[7686]), .B(x[505]), .Z(n4705) );
  NAND U7254 ( .A(n4626), .B(n4705), .Z(n4627) );
  AND U7255 ( .A(n4628), .B(n4627), .Z(n4660) );
  NAND U7256 ( .A(n4630), .B(n4629), .Z(n4634) );
  NAND U7257 ( .A(n4632), .B(n4631), .Z(n4633) );
  AND U7258 ( .A(n4634), .B(n4633), .Z(n4642) );
  NAND U7259 ( .A(n4636), .B(n4635), .Z(n4640) );
  NAND U7260 ( .A(n4638), .B(n4637), .Z(n4639) );
  NAND U7261 ( .A(n4640), .B(n4639), .Z(n4641) );
  XNOR U7262 ( .A(n4642), .B(n4641), .Z(n4658) );
  AND U7263 ( .A(y[7685]), .B(x[506]), .Z(n4644) );
  NAND U7264 ( .A(y[7683]), .B(x[508]), .Z(n4643) );
  XNOR U7265 ( .A(n4644), .B(n4643), .Z(n4648) );
  AND U7266 ( .A(y[7709]), .B(x[482]), .Z(n4646) );
  NAND U7267 ( .A(x[503]), .B(y[7688]), .Z(n4645) );
  XNOR U7268 ( .A(n4646), .B(n4645), .Z(n4647) );
  XOR U7269 ( .A(n4648), .B(n4647), .Z(n4656) );
  AND U7270 ( .A(x[507]), .B(y[7684]), .Z(n4650) );
  NAND U7271 ( .A(y[7710]), .B(x[481]), .Z(n4649) );
  XNOR U7272 ( .A(n4650), .B(n4649), .Z(n4654) );
  AND U7273 ( .A(x[486]), .B(y[7705]), .Z(n4652) );
  NAND U7274 ( .A(x[487]), .B(y[7704]), .Z(n4651) );
  XNOR U7275 ( .A(n4652), .B(n4651), .Z(n4653) );
  XNOR U7276 ( .A(n4654), .B(n4653), .Z(n4655) );
  XNOR U7277 ( .A(n4656), .B(n4655), .Z(n4657) );
  XNOR U7278 ( .A(n4658), .B(n4657), .Z(n4659) );
  XNOR U7279 ( .A(n4660), .B(n4659), .Z(n4676) );
  AND U7280 ( .A(n4662), .B(n4661), .Z(n4666) );
  AND U7281 ( .A(n4664), .B(n4663), .Z(n4665) );
  NOR U7282 ( .A(n4666), .B(n4665), .Z(n4674) );
  NAND U7283 ( .A(n4668), .B(n4667), .Z(n4672) );
  NAND U7284 ( .A(n4670), .B(n4669), .Z(n4671) );
  AND U7285 ( .A(n4672), .B(n4671), .Z(n4673) );
  XNOR U7286 ( .A(n4674), .B(n4673), .Z(n4675) );
  XNOR U7287 ( .A(n4676), .B(n4675), .Z(n4677) );
  XNOR U7288 ( .A(n4678), .B(n4677), .Z(n4761) );
  NAND U7289 ( .A(n4680), .B(n4679), .Z(n4684) );
  NAND U7290 ( .A(n4682), .B(n4681), .Z(n4683) );
  AND U7291 ( .A(n4684), .B(n4683), .Z(n4759) );
  NAND U7292 ( .A(n4686), .B(n4685), .Z(n4690) );
  NAND U7293 ( .A(n4688), .B(n4687), .Z(n4689) );
  AND U7294 ( .A(n4690), .B(n4689), .Z(n4698) );
  NAND U7295 ( .A(n4692), .B(n4691), .Z(n4696) );
  NAND U7296 ( .A(n4694), .B(n4693), .Z(n4695) );
  NAND U7297 ( .A(n4696), .B(n4695), .Z(n4697) );
  XNOR U7298 ( .A(n4698), .B(n4697), .Z(n4757) );
  NAND U7299 ( .A(n4700), .B(n4699), .Z(n4703) );
  AND U7300 ( .A(x[490]), .B(y[7701]), .Z(n4706) );
  NAND U7301 ( .A(n4701), .B(n4706), .Z(n4702) );
  AND U7302 ( .A(n4703), .B(n4702), .Z(n4755) );
  AND U7303 ( .A(x[483]), .B(y[7708]), .Z(n4713) );
  AND U7304 ( .A(n4704), .B(o[30]), .Z(n4711) );
  XOR U7305 ( .A(n4705), .B(o[31]), .Z(n4709) );
  XNOR U7306 ( .A(n4707), .B(n4706), .Z(n4708) );
  XNOR U7307 ( .A(n4709), .B(n4708), .Z(n4710) );
  XNOR U7308 ( .A(n4711), .B(n4710), .Z(n4712) );
  XNOR U7309 ( .A(n4713), .B(n4712), .Z(n4753) );
  AND U7310 ( .A(x[492]), .B(y[7699]), .Z(n4719) );
  AND U7311 ( .A(x[491]), .B(y[7700]), .Z(n4715) );
  NAND U7312 ( .A(y[7694]), .B(x[497]), .Z(n4714) );
  XNOR U7313 ( .A(n4715), .B(n4714), .Z(n4716) );
  XNOR U7314 ( .A(n4717), .B(n4716), .Z(n4718) );
  XNOR U7315 ( .A(n4719), .B(n4718), .Z(n4743) );
  AND U7316 ( .A(x[499]), .B(y[7692]), .Z(n4721) );
  NAND U7317 ( .A(y[7690]), .B(x[501]), .Z(n4720) );
  XNOR U7318 ( .A(n4721), .B(n4720), .Z(n4733) );
  AND U7319 ( .A(y[7702]), .B(x[489]), .Z(n4723) );
  NAND U7320 ( .A(y[7703]), .B(x[488]), .Z(n4722) );
  XNOR U7321 ( .A(n4723), .B(n4722), .Z(n4727) );
  AND U7322 ( .A(y[7682]), .B(x[509]), .Z(n4725) );
  NAND U7323 ( .A(x[494]), .B(y[7697]), .Z(n4724) );
  XNOR U7324 ( .A(n4725), .B(n4724), .Z(n4726) );
  XOR U7325 ( .A(n4727), .B(n4726), .Z(n4731) );
  XNOR U7326 ( .A(n4729), .B(n4728), .Z(n4730) );
  XNOR U7327 ( .A(n4731), .B(n4730), .Z(n4732) );
  XOR U7328 ( .A(n4733), .B(n4732), .Z(n4741) );
  AND U7329 ( .A(y[7693]), .B(x[498]), .Z(n4735) );
  NAND U7330 ( .A(x[511]), .B(y[7680]), .Z(n4734) );
  XNOR U7331 ( .A(n4735), .B(n4734), .Z(n4739) );
  AND U7332 ( .A(x[485]), .B(y[7706]), .Z(n4737) );
  NAND U7333 ( .A(y[7707]), .B(x[484]), .Z(n4736) );
  XNOR U7334 ( .A(n4737), .B(n4736), .Z(n4738) );
  XNOR U7335 ( .A(n4739), .B(n4738), .Z(n4740) );
  XNOR U7336 ( .A(n4741), .B(n4740), .Z(n4742) );
  XOR U7337 ( .A(n4743), .B(n4742), .Z(n4751) );
  AND U7338 ( .A(x[496]), .B(y[7695]), .Z(n4745) );
  NAND U7339 ( .A(x[510]), .B(y[7681]), .Z(n4744) );
  XNOR U7340 ( .A(n4745), .B(n4744), .Z(n4749) );
  AND U7341 ( .A(y[7711]), .B(x[480]), .Z(n4747) );
  NAND U7342 ( .A(x[500]), .B(y[7691]), .Z(n4746) );
  XNOR U7343 ( .A(n4747), .B(n4746), .Z(n4748) );
  XNOR U7344 ( .A(n4749), .B(n4748), .Z(n4750) );
  XNOR U7345 ( .A(n4751), .B(n4750), .Z(n4752) );
  XNOR U7346 ( .A(n4753), .B(n4752), .Z(n4754) );
  XNOR U7347 ( .A(n4755), .B(n4754), .Z(n4756) );
  XNOR U7348 ( .A(n4757), .B(n4756), .Z(n4758) );
  XNOR U7349 ( .A(n4759), .B(n4758), .Z(n4760) );
  XNOR U7350 ( .A(n4761), .B(n4760), .Z(n4762) );
  XNOR U7351 ( .A(n4763), .B(n4762), .Z(n4779) );
  NAND U7352 ( .A(n4765), .B(n4764), .Z(n4769) );
  NAND U7353 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U7354 ( .A(n4769), .B(n4768), .Z(n4777) );
  NAND U7355 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U7356 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U7357 ( .A(n4775), .B(n4774), .Z(n4776) );
  XNOR U7358 ( .A(n4777), .B(n4776), .Z(n4778) );
  XNOR U7359 ( .A(n4779), .B(n4778), .Z(n4780) );
  XNOR U7360 ( .A(n4781), .B(n4780), .Z(n4782) );
  XNOR U7361 ( .A(n4783), .B(n4782), .Z(n4784) );
  XNOR U7362 ( .A(n4785), .B(n4784), .Z(n4801) );
  NANDN U7363 ( .A(n4787), .B(n4786), .Z(n4791) );
  NAND U7364 ( .A(n4789), .B(n4788), .Z(n4790) );
  AND U7365 ( .A(n4791), .B(n4790), .Z(n4799) );
  NAND U7366 ( .A(n4793), .B(n4792), .Z(n4797) );
  NANDN U7367 ( .A(n4795), .B(n4794), .Z(n4796) );
  NAND U7368 ( .A(n4797), .B(n4796), .Z(n4798) );
  XNOR U7369 ( .A(n4799), .B(n4798), .Z(n4800) );
  XNOR U7370 ( .A(n4801), .B(n4800), .Z(n4802) );
  XNOR U7371 ( .A(n4803), .B(n4802), .Z(n4827) );
  NAND U7372 ( .A(n4805), .B(n4804), .Z(n4809) );
  NAND U7373 ( .A(n4807), .B(n4806), .Z(n4808) );
  AND U7374 ( .A(n4809), .B(n4808), .Z(n4817) );
  ANDN U7375 ( .B(n4811), .A(n4810), .Z(n4815) );
  AND U7376 ( .A(n4813), .B(n4812), .Z(n4814) );
  OR U7377 ( .A(n4815), .B(n4814), .Z(n4816) );
  XNOR U7378 ( .A(n4817), .B(n4816), .Z(n4825) );
  NAND U7379 ( .A(n4819), .B(n4818), .Z(n4823) );
  NAND U7380 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U7381 ( .A(n4823), .B(n4822), .Z(n4824) );
  XNOR U7382 ( .A(n4825), .B(n4824), .Z(n4826) );
  XNOR U7383 ( .A(n4827), .B(n4826), .Z(n4828) );
  XNOR U7384 ( .A(n4829), .B(n4828), .Z(n4845) );
  NANDN U7385 ( .A(n4831), .B(n4830), .Z(n4835) );
  NANDN U7386 ( .A(n4833), .B(n4832), .Z(n4834) );
  AND U7387 ( .A(n4835), .B(n4834), .Z(n4843) );
  NAND U7388 ( .A(n4837), .B(n4836), .Z(n4841) );
  NANDN U7389 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U7390 ( .A(n4841), .B(n4840), .Z(n4842) );
  XNOR U7391 ( .A(n4843), .B(n4842), .Z(n4844) );
  XNOR U7392 ( .A(n4845), .B(n4844), .Z(n4846) );
  XNOR U7393 ( .A(n4847), .B(n4846), .Z(n4863) );
  NAND U7394 ( .A(n4849), .B(n4848), .Z(n4853) );
  NAND U7395 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U7396 ( .A(n4853), .B(n4852), .Z(n4861) );
  NANDN U7397 ( .A(n4855), .B(n4854), .Z(n4859) );
  NAND U7398 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U7399 ( .A(n4859), .B(n4858), .Z(n4860) );
  XNOR U7400 ( .A(n4861), .B(n4860), .Z(n4862) );
  XNOR U7401 ( .A(n4863), .B(n4862), .Z(N64) );
  AND U7402 ( .A(x[480]), .B(y[7712]), .Z(n5512) );
  XOR U7403 ( .A(n5512), .B(o[32]), .Z(N97) );
  AND U7404 ( .A(x[481]), .B(y[7712]), .Z(n4872) );
  AND U7405 ( .A(x[480]), .B(y[7713]), .Z(n4871) );
  XNOR U7406 ( .A(n4871), .B(o[33]), .Z(n4864) );
  XNOR U7407 ( .A(n4872), .B(n4864), .Z(n4866) );
  NAND U7408 ( .A(n5512), .B(o[32]), .Z(n4865) );
  XNOR U7409 ( .A(n4866), .B(n4865), .Z(N98) );
  NANDN U7410 ( .A(n4872), .B(n4864), .Z(n4868) );
  NAND U7411 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U7412 ( .A(n4868), .B(n4867), .Z(n4878) );
  AND U7413 ( .A(x[480]), .B(y[7714]), .Z(n4885) );
  XNOR U7414 ( .A(n4885), .B(o[34]), .Z(n4877) );
  XNOR U7415 ( .A(n4878), .B(n4877), .Z(n4880) );
  AND U7416 ( .A(y[7712]), .B(x[482]), .Z(n4870) );
  NAND U7417 ( .A(y[7713]), .B(x[481]), .Z(n4869) );
  XNOR U7418 ( .A(n4870), .B(n4869), .Z(n4874) );
  AND U7419 ( .A(n4871), .B(o[33]), .Z(n4873) );
  XNOR U7420 ( .A(n4874), .B(n4873), .Z(n4879) );
  XNOR U7421 ( .A(n4880), .B(n4879), .Z(N99) );
  AND U7422 ( .A(x[482]), .B(y[7713]), .Z(n4892) );
  NAND U7423 ( .A(n4892), .B(n4872), .Z(n4876) );
  NAND U7424 ( .A(n4874), .B(n4873), .Z(n4875) );
  AND U7425 ( .A(n4876), .B(n4875), .Z(n4895) );
  NANDN U7426 ( .A(n4878), .B(n4877), .Z(n4882) );
  NAND U7427 ( .A(n4880), .B(n4879), .Z(n4881) );
  AND U7428 ( .A(n4882), .B(n4881), .Z(n4894) );
  XNOR U7429 ( .A(n4895), .B(n4894), .Z(n4897) );
  AND U7430 ( .A(x[481]), .B(y[7714]), .Z(n5014) );
  XOR U7431 ( .A(n4892), .B(o[35]), .Z(n4900) );
  XOR U7432 ( .A(n5014), .B(n4900), .Z(n4902) );
  AND U7433 ( .A(y[7712]), .B(x[483]), .Z(n4884) );
  NAND U7434 ( .A(y[7715]), .B(x[480]), .Z(n4883) );
  XNOR U7435 ( .A(n4884), .B(n4883), .Z(n4887) );
  AND U7436 ( .A(n4885), .B(o[34]), .Z(n4886) );
  XOR U7437 ( .A(n4887), .B(n4886), .Z(n4901) );
  XOR U7438 ( .A(n4902), .B(n4901), .Z(n4896) );
  XOR U7439 ( .A(n4897), .B(n4896), .Z(N100) );
  AND U7440 ( .A(x[483]), .B(y[7715]), .Z(n4945) );
  NAND U7441 ( .A(n5512), .B(n4945), .Z(n4889) );
  NAND U7442 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U7443 ( .A(n4889), .B(n4888), .Z(n4923) );
  AND U7444 ( .A(y[7716]), .B(x[480]), .Z(n4891) );
  NAND U7445 ( .A(y[7712]), .B(x[484]), .Z(n4890) );
  XNOR U7446 ( .A(n4891), .B(n4890), .Z(n4916) );
  NAND U7447 ( .A(n4892), .B(o[35]), .Z(n4917) );
  AND U7448 ( .A(y[7714]), .B(x[482]), .Z(n5041) );
  NAND U7449 ( .A(y[7715]), .B(x[481]), .Z(n4893) );
  XNOR U7450 ( .A(n5041), .B(n4893), .Z(n4913) );
  AND U7451 ( .A(x[483]), .B(y[7713]), .Z(n4908) );
  XOR U7452 ( .A(o[36]), .B(n4908), .Z(n4912) );
  XOR U7453 ( .A(n4913), .B(n4912), .Z(n4920) );
  XOR U7454 ( .A(n4921), .B(n4920), .Z(n4922) );
  XOR U7455 ( .A(n4923), .B(n4922), .Z(n4927) );
  NANDN U7456 ( .A(n4895), .B(n4894), .Z(n4899) );
  NAND U7457 ( .A(n4897), .B(n4896), .Z(n4898) );
  NAND U7458 ( .A(n4899), .B(n4898), .Z(n4928) );
  NAND U7459 ( .A(n5014), .B(n4900), .Z(n4904) );
  NAND U7460 ( .A(n4902), .B(n4901), .Z(n4903) );
  NAND U7461 ( .A(n4904), .B(n4903), .Z(n4929) );
  IV U7462 ( .A(n4929), .Z(n4926) );
  XOR U7463 ( .A(n4928), .B(n4926), .Z(n4905) );
  XNOR U7464 ( .A(n4927), .B(n4905), .Z(N101) );
  AND U7465 ( .A(y[7714]), .B(x[483]), .Z(n4907) );
  NAND U7466 ( .A(y[7716]), .B(x[481]), .Z(n4906) );
  XNOR U7467 ( .A(n4907), .B(n4906), .Z(n4932) );
  AND U7468 ( .A(x[484]), .B(y[7713]), .Z(n4941) );
  XOR U7469 ( .A(n4941), .B(o[37]), .Z(n4931) );
  XNOR U7470 ( .A(n4932), .B(n4931), .Z(n4935) );
  NAND U7471 ( .A(x[482]), .B(y[7715]), .Z(n5023) );
  AND U7472 ( .A(o[36]), .B(n4908), .Z(n4937) );
  AND U7473 ( .A(y[7712]), .B(x[485]), .Z(n4910) );
  NAND U7474 ( .A(y[7717]), .B(x[480]), .Z(n4909) );
  XNOR U7475 ( .A(n4910), .B(n4909), .Z(n4938) );
  XOR U7476 ( .A(n4937), .B(n4938), .Z(n4936) );
  XOR U7477 ( .A(n5023), .B(n4936), .Z(n4911) );
  XOR U7478 ( .A(n4935), .B(n4911), .Z(n4953) );
  NANDN U7479 ( .A(n5023), .B(n5014), .Z(n4915) );
  NAND U7480 ( .A(n4913), .B(n4912), .Z(n4914) );
  AND U7481 ( .A(n4915), .B(n4914), .Z(n4951) );
  AND U7482 ( .A(x[484]), .B(y[7716]), .Z(n5712) );
  NAND U7483 ( .A(n5712), .B(n5512), .Z(n4919) );
  NANDN U7484 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U7485 ( .A(n4919), .B(n4918), .Z(n4950) );
  XNOR U7486 ( .A(n4953), .B(n4952), .Z(n4949) );
  NAND U7487 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U7488 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U7489 ( .A(n4925), .B(n4924), .Z(n4948) );
  XOR U7490 ( .A(n4948), .B(n4947), .Z(n4930) );
  XNOR U7491 ( .A(n4949), .B(n4930), .Z(N102) );
  AND U7492 ( .A(x[483]), .B(y[7716]), .Z(n5025) );
  NAND U7493 ( .A(n5014), .B(n5025), .Z(n4934) );
  NAND U7494 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U7495 ( .A(n4934), .B(n4933), .Z(n4989) );
  XOR U7496 ( .A(n4989), .B(n4988), .Z(n4991) );
  AND U7497 ( .A(x[485]), .B(y[7717]), .Z(n5183) );
  NAND U7498 ( .A(n5512), .B(n5183), .Z(n4940) );
  NAND U7499 ( .A(n4938), .B(n4937), .Z(n4939) );
  NAND U7500 ( .A(n4940), .B(n4939), .Z(n4958) );
  AND U7501 ( .A(n4941), .B(o[37]), .Z(n4964) );
  AND U7502 ( .A(y[7712]), .B(x[486]), .Z(n4943) );
  NAND U7503 ( .A(y[7718]), .B(x[480]), .Z(n4942) );
  XNOR U7504 ( .A(n4943), .B(n4942), .Z(n4965) );
  XOR U7505 ( .A(n4964), .B(n4965), .Z(n4957) );
  XOR U7506 ( .A(n4958), .B(n4957), .Z(n4960) );
  NAND U7507 ( .A(y[7716]), .B(x[482]), .Z(n4944) );
  XNOR U7508 ( .A(n4945), .B(n4944), .Z(n4969) );
  AND U7509 ( .A(y[7717]), .B(x[481]), .Z(n5217) );
  NAND U7510 ( .A(y[7714]), .B(x[484]), .Z(n4946) );
  XNOR U7511 ( .A(n5217), .B(n4946), .Z(n4973) );
  AND U7512 ( .A(x[485]), .B(y[7713]), .Z(n4978) );
  XOR U7513 ( .A(o[38]), .B(n4978), .Z(n4972) );
  XOR U7514 ( .A(n4973), .B(n4972), .Z(n4968) );
  XOR U7515 ( .A(n4969), .B(n4968), .Z(n4959) );
  XOR U7516 ( .A(n4960), .B(n4959), .Z(n4990) );
  XNOR U7517 ( .A(n4991), .B(n4990), .Z(n4984) );
  NANDN U7518 ( .A(n4951), .B(n4950), .Z(n4955) );
  NAND U7519 ( .A(n4953), .B(n4952), .Z(n4954) );
  NAND U7520 ( .A(n4955), .B(n4954), .Z(n4982) );
  IV U7521 ( .A(n4982), .Z(n4981) );
  XOR U7522 ( .A(n4983), .B(n4981), .Z(n4956) );
  XNOR U7523 ( .A(n4984), .B(n4956), .Z(N103) );
  NAND U7524 ( .A(n4958), .B(n4957), .Z(n4962) );
  NAND U7525 ( .A(n4960), .B(n4959), .Z(n4961) );
  AND U7526 ( .A(n4962), .B(n4961), .Z(n4998) );
  AND U7527 ( .A(x[485]), .B(y[7714]), .Z(n5091) );
  NAND U7528 ( .A(y[7718]), .B(x[481]), .Z(n4963) );
  XNOR U7529 ( .A(n5091), .B(n4963), .Z(n5016) );
  NAND U7530 ( .A(x[486]), .B(y[7713]), .Z(n5020) );
  XOR U7531 ( .A(n5016), .B(n5015), .Z(n5035) );
  AND U7532 ( .A(x[486]), .B(y[7718]), .Z(n5237) );
  NAND U7533 ( .A(n5512), .B(n5237), .Z(n4967) );
  NAND U7534 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U7535 ( .A(n4967), .B(n4966), .Z(n5034) );
  NANDN U7536 ( .A(n5023), .B(n5025), .Z(n4971) );
  NAND U7537 ( .A(n4969), .B(n4968), .Z(n4970) );
  AND U7538 ( .A(n4971), .B(n4970), .Z(n5036) );
  XOR U7539 ( .A(n5037), .B(n5036), .Z(n4996) );
  AND U7540 ( .A(x[484]), .B(y[7717]), .Z(n5517) );
  NAND U7541 ( .A(n5517), .B(n5014), .Z(n4975) );
  NAND U7542 ( .A(n4973), .B(n4972), .Z(n4974) );
  AND U7543 ( .A(n4975), .B(n4974), .Z(n5011) );
  AND U7544 ( .A(y[7717]), .B(x[482]), .Z(n4977) );
  NAND U7545 ( .A(y[7715]), .B(x[484]), .Z(n4976) );
  XNOR U7546 ( .A(n4977), .B(n4976), .Z(n5024) );
  XNOR U7547 ( .A(n5025), .B(n5024), .Z(n5009) );
  AND U7548 ( .A(o[38]), .B(n4978), .Z(n5029) );
  AND U7549 ( .A(y[7712]), .B(x[487]), .Z(n4980) );
  NAND U7550 ( .A(y[7719]), .B(x[480]), .Z(n4979) );
  XNOR U7551 ( .A(n4980), .B(n4979), .Z(n5028) );
  XNOR U7552 ( .A(n5029), .B(n5028), .Z(n5008) );
  XOR U7553 ( .A(n5009), .B(n5008), .Z(n5010) );
  XOR U7554 ( .A(n5011), .B(n5010), .Z(n4995) );
  XOR U7555 ( .A(n4996), .B(n4995), .Z(n4997) );
  XNOR U7556 ( .A(n4998), .B(n4997), .Z(n5004) );
  OR U7557 ( .A(n4983), .B(n4981), .Z(n4987) );
  ANDN U7558 ( .B(n4983), .A(n4982), .Z(n4985) );
  OR U7559 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U7560 ( .A(n4987), .B(n4986), .Z(n5002) );
  NAND U7561 ( .A(n4989), .B(n4988), .Z(n4993) );
  NAND U7562 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U7563 ( .A(n4993), .B(n4992), .Z(n5003) );
  IV U7564 ( .A(n5003), .Z(n5001) );
  XOR U7565 ( .A(n5002), .B(n5001), .Z(n4994) );
  XNOR U7566 ( .A(n5004), .B(n4994), .Z(N104) );
  NAND U7567 ( .A(n4996), .B(n4995), .Z(n5000) );
  NAND U7568 ( .A(n4998), .B(n4997), .Z(n4999) );
  AND U7569 ( .A(n5000), .B(n4999), .Z(n5076) );
  NANDN U7570 ( .A(n5001), .B(n5002), .Z(n5007) );
  NOR U7571 ( .A(n5003), .B(n5002), .Z(n5005) );
  OR U7572 ( .A(n5005), .B(n5004), .Z(n5006) );
  AND U7573 ( .A(n5007), .B(n5006), .Z(n5075) );
  NAND U7574 ( .A(n5009), .B(n5008), .Z(n5013) );
  NAND U7575 ( .A(n5011), .B(n5010), .Z(n5012) );
  AND U7576 ( .A(n5013), .B(n5012), .Z(n5072) );
  AND U7577 ( .A(x[485]), .B(y[7718]), .Z(n5175) );
  NAND U7578 ( .A(n5175), .B(n5014), .Z(n5018) );
  NAND U7579 ( .A(n5016), .B(n5015), .Z(n5017) );
  NAND U7580 ( .A(n5018), .B(n5017), .Z(n5070) );
  AND U7581 ( .A(x[485]), .B(y[7715]), .Z(n5653) );
  NAND U7582 ( .A(y[7719]), .B(x[481]), .Z(n5019) );
  XNOR U7583 ( .A(n5653), .B(n5019), .Z(n5060) );
  ANDN U7584 ( .B(o[39]), .A(n5020), .Z(n5059) );
  XOR U7585 ( .A(n5060), .B(n5059), .Z(n5047) );
  NAND U7586 ( .A(x[483]), .B(y[7717]), .Z(n5848) );
  AND U7587 ( .A(y[7714]), .B(x[486]), .Z(n5022) );
  NAND U7588 ( .A(y[7718]), .B(x[482]), .Z(n5021) );
  XNOR U7589 ( .A(n5022), .B(n5021), .Z(n5042) );
  XNOR U7590 ( .A(n5712), .B(n5042), .Z(n5045) );
  XOR U7591 ( .A(n5848), .B(n5045), .Z(n5046) );
  XOR U7592 ( .A(n5047), .B(n5046), .Z(n5069) );
  XOR U7593 ( .A(n5070), .B(n5069), .Z(n5071) );
  XOR U7594 ( .A(n5072), .B(n5071), .Z(n5081) );
  NANDN U7595 ( .A(n5023), .B(n5517), .Z(n5027) );
  NAND U7596 ( .A(n5025), .B(n5024), .Z(n5026) );
  NAND U7597 ( .A(n5027), .B(n5026), .Z(n5066) );
  AND U7598 ( .A(x[487]), .B(y[7719]), .Z(n5393) );
  NAND U7599 ( .A(n5512), .B(n5393), .Z(n5031) );
  NAND U7600 ( .A(n5029), .B(n5028), .Z(n5030) );
  NAND U7601 ( .A(n5031), .B(n5030), .Z(n5064) );
  AND U7602 ( .A(y[7712]), .B(x[488]), .Z(n5033) );
  NAND U7603 ( .A(y[7720]), .B(x[480]), .Z(n5032) );
  XNOR U7604 ( .A(n5033), .B(n5032), .Z(n5050) );
  NAND U7605 ( .A(x[487]), .B(y[7713]), .Z(n5055) );
  XOR U7606 ( .A(n5050), .B(n5049), .Z(n5063) );
  XOR U7607 ( .A(n5064), .B(n5063), .Z(n5065) );
  XOR U7608 ( .A(n5066), .B(n5065), .Z(n5079) );
  NANDN U7609 ( .A(n5035), .B(n5034), .Z(n5039) );
  NAND U7610 ( .A(n5037), .B(n5036), .Z(n5038) );
  NAND U7611 ( .A(n5039), .B(n5038), .Z(n5078) );
  XNOR U7612 ( .A(n5075), .B(n5077), .Z(n5040) );
  XOR U7613 ( .A(n5076), .B(n5040), .Z(N105) );
  NAND U7614 ( .A(n5237), .B(n5041), .Z(n5044) );
  NAND U7615 ( .A(n5712), .B(n5042), .Z(n5043) );
  AND U7616 ( .A(n5044), .B(n5043), .Z(n5086) );
  AND U7617 ( .A(x[488]), .B(y[7720]), .Z(n5048) );
  NAND U7618 ( .A(n5048), .B(n5512), .Z(n5052) );
  NAND U7619 ( .A(n5050), .B(n5049), .Z(n5051) );
  AND U7620 ( .A(n5052), .B(n5051), .Z(n5120) );
  AND U7621 ( .A(y[7716]), .B(x[485]), .Z(n5054) );
  NAND U7622 ( .A(y[7714]), .B(x[487]), .Z(n5053) );
  XNOR U7623 ( .A(n5054), .B(n5053), .Z(n5093) );
  ANDN U7624 ( .B(o[40]), .A(n5055), .Z(n5092) );
  XOR U7625 ( .A(n5093), .B(n5092), .Z(n5118) );
  AND U7626 ( .A(y[7712]), .B(x[489]), .Z(n5057) );
  NAND U7627 ( .A(y[7721]), .B(x[480]), .Z(n5056) );
  XNOR U7628 ( .A(n5057), .B(n5056), .Z(n5100) );
  NAND U7629 ( .A(x[488]), .B(y[7713]), .Z(n5109) );
  XNOR U7630 ( .A(n5100), .B(n5099), .Z(n5117) );
  XOR U7631 ( .A(n5120), .B(n5119), .Z(n5114) );
  AND U7632 ( .A(y[7715]), .B(x[486]), .Z(n5460) );
  NAND U7633 ( .A(y[7720]), .B(x[481]), .Z(n5058) );
  XNOR U7634 ( .A(n5460), .B(n5058), .Z(n5104) );
  XNOR U7635 ( .A(n5517), .B(n5104), .Z(n5123) );
  NAND U7636 ( .A(x[482]), .B(y[7719]), .Z(n5759) );
  AND U7637 ( .A(x[483]), .B(y[7718]), .Z(n5470) );
  XOR U7638 ( .A(n5759), .B(n5470), .Z(n5124) );
  XOR U7639 ( .A(n5123), .B(n5124), .Z(n5112) );
  NAND U7640 ( .A(x[485]), .B(y[7719]), .Z(n5300) );
  AND U7641 ( .A(x[481]), .B(y[7715]), .Z(n5103) );
  NANDN U7642 ( .A(n5300), .B(n5103), .Z(n5062) );
  NAND U7643 ( .A(n5060), .B(n5059), .Z(n5061) );
  NAND U7644 ( .A(n5062), .B(n5061), .Z(n5111) );
  XOR U7645 ( .A(n5112), .B(n5111), .Z(n5113) );
  XOR U7646 ( .A(n5088), .B(n5087), .Z(n5137) );
  NAND U7647 ( .A(n5064), .B(n5063), .Z(n5068) );
  NAND U7648 ( .A(n5066), .B(n5065), .Z(n5067) );
  NAND U7649 ( .A(n5068), .B(n5067), .Z(n5135) );
  NAND U7650 ( .A(n5070), .B(n5069), .Z(n5074) );
  NAND U7651 ( .A(n5072), .B(n5071), .Z(n5073) );
  NAND U7652 ( .A(n5074), .B(n5073), .Z(n5134) );
  XOR U7653 ( .A(n5135), .B(n5134), .Z(n5136) );
  XNOR U7654 ( .A(n5137), .B(n5136), .Z(n5130) );
  NANDN U7655 ( .A(n5079), .B(n5078), .Z(n5083) );
  NANDN U7656 ( .A(n5081), .B(n5080), .Z(n5082) );
  AND U7657 ( .A(n5083), .B(n5082), .Z(n5128) );
  IV U7658 ( .A(n5128), .Z(n5127) );
  XOR U7659 ( .A(n5129), .B(n5127), .Z(n5084) );
  XNOR U7660 ( .A(n5130), .B(n5084), .Z(N106) );
  NANDN U7661 ( .A(n5086), .B(n5085), .Z(n5090) );
  NAND U7662 ( .A(n5088), .B(n5087), .Z(n5089) );
  AND U7663 ( .A(n5090), .B(n5089), .Z(n5196) );
  AND U7664 ( .A(x[487]), .B(y[7716]), .Z(n5177) );
  NAND U7665 ( .A(n5177), .B(n5091), .Z(n5095) );
  NAND U7666 ( .A(n5093), .B(n5092), .Z(n5094) );
  AND U7667 ( .A(n5095), .B(n5094), .Z(n5190) );
  AND U7668 ( .A(y[7715]), .B(x[487]), .Z(n5097) );
  NAND U7669 ( .A(y[7718]), .B(x[484]), .Z(n5096) );
  XNOR U7670 ( .A(n5097), .B(n5096), .Z(n5161) );
  AND U7671 ( .A(x[486]), .B(y[7716]), .Z(n5160) );
  XOR U7672 ( .A(n5161), .B(n5160), .Z(n5188) );
  AND U7673 ( .A(x[488]), .B(y[7714]), .Z(n5357) );
  AND U7674 ( .A(x[489]), .B(y[7713]), .Z(n5171) );
  XOR U7675 ( .A(o[42]), .B(n5171), .Z(n5182) );
  XOR U7676 ( .A(n5357), .B(n5182), .Z(n5184) );
  XNOR U7677 ( .A(n5184), .B(n5183), .Z(n5187) );
  XNOR U7678 ( .A(n5190), .B(n5189), .Z(n5149) );
  AND U7679 ( .A(x[489]), .B(y[7721]), .Z(n5098) );
  NAND U7680 ( .A(n5098), .B(n5512), .Z(n5102) );
  NAND U7681 ( .A(n5100), .B(n5099), .Z(n5101) );
  NAND U7682 ( .A(n5102), .B(n5101), .Z(n5147) );
  AND U7683 ( .A(x[486]), .B(y[7720]), .Z(n5384) );
  NAND U7684 ( .A(n5384), .B(n5103), .Z(n5106) );
  NAND U7685 ( .A(n5104), .B(n5517), .Z(n5105) );
  AND U7686 ( .A(n5106), .B(n5105), .Z(n5156) );
  AND U7687 ( .A(y[7712]), .B(x[490]), .Z(n5108) );
  NAND U7688 ( .A(y[7722]), .B(x[480]), .Z(n5107) );
  XNOR U7689 ( .A(n5108), .B(n5107), .Z(n5166) );
  ANDN U7690 ( .B(o[41]), .A(n5109), .Z(n5165) );
  XOR U7691 ( .A(n5166), .B(n5165), .Z(n5154) );
  AND U7692 ( .A(y[7719]), .B(x[483]), .Z(n6088) );
  NAND U7693 ( .A(y[7721]), .B(x[481]), .Z(n5110) );
  XNOR U7694 ( .A(n6088), .B(n5110), .Z(n5178) );
  NAND U7695 ( .A(x[482]), .B(y[7720]), .Z(n5179) );
  XOR U7696 ( .A(n5154), .B(n5153), .Z(n5155) );
  XOR U7697 ( .A(n5147), .B(n5148), .Z(n5150) );
  XOR U7698 ( .A(n5149), .B(n5150), .Z(n5194) );
  NAND U7699 ( .A(n5112), .B(n5111), .Z(n5116) );
  NANDN U7700 ( .A(n5114), .B(n5113), .Z(n5115) );
  NAND U7701 ( .A(n5116), .B(n5115), .Z(n5143) );
  NANDN U7702 ( .A(n5118), .B(n5117), .Z(n5122) );
  NAND U7703 ( .A(n5120), .B(n5119), .Z(n5121) );
  AND U7704 ( .A(n5122), .B(n5121), .Z(n5142) );
  NANDN U7705 ( .A(n5124), .B(n5123), .Z(n5126) );
  ANDN U7706 ( .B(n5759), .A(n5470), .Z(n5125) );
  ANDN U7707 ( .B(n5126), .A(n5125), .Z(n5141) );
  XOR U7708 ( .A(n5142), .B(n5141), .Z(n5144) );
  XNOR U7709 ( .A(n5143), .B(n5144), .Z(n5193) );
  XOR U7710 ( .A(n5194), .B(n5193), .Z(n5195) );
  XNOR U7711 ( .A(n5196), .B(n5195), .Z(n5202) );
  OR U7712 ( .A(n5129), .B(n5127), .Z(n5133) );
  ANDN U7713 ( .B(n5129), .A(n5128), .Z(n5131) );
  OR U7714 ( .A(n5131), .B(n5130), .Z(n5132) );
  AND U7715 ( .A(n5133), .B(n5132), .Z(n5200) );
  NAND U7716 ( .A(n5135), .B(n5134), .Z(n5139) );
  NAND U7717 ( .A(n5137), .B(n5136), .Z(n5138) );
  AND U7718 ( .A(n5139), .B(n5138), .Z(n5201) );
  IV U7719 ( .A(n5201), .Z(n5199) );
  XOR U7720 ( .A(n5200), .B(n5199), .Z(n5140) );
  XNOR U7721 ( .A(n5202), .B(n5140), .Z(N107) );
  NAND U7722 ( .A(n5142), .B(n5141), .Z(n5146) );
  NAND U7723 ( .A(n5144), .B(n5143), .Z(n5145) );
  NAND U7724 ( .A(n5146), .B(n5145), .Z(n5267) );
  NANDN U7725 ( .A(n5148), .B(n5147), .Z(n5152) );
  NANDN U7726 ( .A(n5150), .B(n5149), .Z(n5151) );
  NAND U7727 ( .A(n5152), .B(n5151), .Z(n5266) );
  NAND U7728 ( .A(n5154), .B(n5153), .Z(n5158) );
  NANDN U7729 ( .A(n5156), .B(n5155), .Z(n5157) );
  AND U7730 ( .A(n5158), .B(n5157), .Z(n5259) );
  AND U7731 ( .A(x[487]), .B(y[7718]), .Z(n5295) );
  AND U7732 ( .A(x[484]), .B(y[7715]), .Z(n5159) );
  NAND U7733 ( .A(n5295), .B(n5159), .Z(n5163) );
  NAND U7734 ( .A(n5161), .B(n5160), .Z(n5162) );
  AND U7735 ( .A(n5163), .B(n5162), .Z(n5257) );
  AND U7736 ( .A(x[490]), .B(y[7722]), .Z(n5164) );
  NAND U7737 ( .A(n5164), .B(n5512), .Z(n5168) );
  NAND U7738 ( .A(n5166), .B(n5165), .Z(n5167) );
  AND U7739 ( .A(n5168), .B(n5167), .Z(n5253) );
  AND U7740 ( .A(y[7712]), .B(x[491]), .Z(n5170) );
  NAND U7741 ( .A(y[7723]), .B(x[480]), .Z(n5169) );
  XNOR U7742 ( .A(n5170), .B(n5169), .Z(n5228) );
  AND U7743 ( .A(o[42]), .B(n5171), .Z(n5227) );
  XOR U7744 ( .A(n5228), .B(n5227), .Z(n5251) );
  AND U7745 ( .A(y[7717]), .B(x[486]), .Z(n5173) );
  NAND U7746 ( .A(y[7722]), .B(x[481]), .Z(n5172) );
  XNOR U7747 ( .A(n5173), .B(n5172), .Z(n5219) );
  AND U7748 ( .A(x[490]), .B(y[7713]), .Z(n5238) );
  XOR U7749 ( .A(o[43]), .B(n5238), .Z(n5218) );
  XOR U7750 ( .A(n5219), .B(n5218), .Z(n5250) );
  XOR U7751 ( .A(n5251), .B(n5250), .Z(n5252) );
  AND U7752 ( .A(x[483]), .B(y[7720]), .Z(n6233) );
  NAND U7753 ( .A(y[7721]), .B(x[482]), .Z(n5174) );
  XNOR U7754 ( .A(n5175), .B(n5174), .Z(n5214) );
  AND U7755 ( .A(x[484]), .B(y[7719]), .Z(n5213) );
  XNOR U7756 ( .A(n5214), .B(n5213), .Z(n5245) );
  XNOR U7757 ( .A(n6233), .B(n5245), .Z(n5247) );
  NAND U7758 ( .A(y[7714]), .B(x[489]), .Z(n5176) );
  XNOR U7759 ( .A(n5177), .B(n5176), .Z(n5233) );
  AND U7760 ( .A(x[488]), .B(y[7715]), .Z(n5232) );
  XNOR U7761 ( .A(n5233), .B(n5232), .Z(n5246) );
  XOR U7762 ( .A(n5247), .B(n5246), .Z(n5210) );
  NAND U7763 ( .A(x[483]), .B(y[7721]), .Z(n5291) );
  AND U7764 ( .A(x[481]), .B(y[7719]), .Z(n5507) );
  NANDN U7765 ( .A(n5291), .B(n5507), .Z(n5181) );
  NANDN U7766 ( .A(n5179), .B(n5178), .Z(n5180) );
  AND U7767 ( .A(n5181), .B(n5180), .Z(n5208) );
  NAND U7768 ( .A(n5357), .B(n5182), .Z(n5186) );
  NAND U7769 ( .A(n5184), .B(n5183), .Z(n5185) );
  NAND U7770 ( .A(n5186), .B(n5185), .Z(n5207) );
  NANDN U7771 ( .A(n5188), .B(n5187), .Z(n5192) );
  NAND U7772 ( .A(n5190), .B(n5189), .Z(n5191) );
  NAND U7773 ( .A(n5192), .B(n5191), .Z(n5239) );
  XOR U7774 ( .A(n5240), .B(n5239), .Z(n5242) );
  XNOR U7775 ( .A(n5241), .B(n5242), .Z(n5265) );
  XOR U7776 ( .A(n5266), .B(n5265), .Z(n5268) );
  XOR U7777 ( .A(n5267), .B(n5268), .Z(n5264) );
  NAND U7778 ( .A(n5194), .B(n5193), .Z(n5198) );
  NAND U7779 ( .A(n5196), .B(n5195), .Z(n5197) );
  NAND U7780 ( .A(n5198), .B(n5197), .Z(n5262) );
  NANDN U7781 ( .A(n5199), .B(n5200), .Z(n5205) );
  NOR U7782 ( .A(n5201), .B(n5200), .Z(n5203) );
  OR U7783 ( .A(n5203), .B(n5202), .Z(n5204) );
  AND U7784 ( .A(n5205), .B(n5204), .Z(n5263) );
  XOR U7785 ( .A(n5262), .B(n5263), .Z(n5206) );
  XNOR U7786 ( .A(n5264), .B(n5206), .Z(N108) );
  NANDN U7787 ( .A(n5208), .B(n5207), .Z(n5212) );
  NANDN U7788 ( .A(n5210), .B(n5209), .Z(n5211) );
  AND U7789 ( .A(n5212), .B(n5211), .Z(n5332) );
  AND U7790 ( .A(x[482]), .B(y[7718]), .Z(n5946) );
  AND U7791 ( .A(x[485]), .B(y[7721]), .Z(n5750) );
  NAND U7792 ( .A(n5946), .B(n5750), .Z(n5216) );
  NAND U7793 ( .A(n5214), .B(n5213), .Z(n5215) );
  NAND U7794 ( .A(n5216), .B(n5215), .Z(n5279) );
  AND U7795 ( .A(y[7722]), .B(x[486]), .Z(n5524) );
  NAND U7796 ( .A(n5524), .B(n5217), .Z(n5221) );
  NAND U7797 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U7798 ( .A(n5221), .B(n5220), .Z(n5278) );
  XOR U7799 ( .A(n5279), .B(n5278), .Z(n5281) );
  AND U7800 ( .A(x[489]), .B(y[7715]), .Z(n5941) );
  AND U7801 ( .A(x[490]), .B(y[7714]), .Z(n5983) );
  AND U7802 ( .A(y[7720]), .B(x[484]), .Z(n5222) );
  XOR U7803 ( .A(n5983), .B(n5222), .Z(n5322) );
  XOR U7804 ( .A(n5941), .B(n5322), .Z(n5301) );
  NAND U7805 ( .A(x[487]), .B(y[7717]), .Z(n5299) );
  XOR U7806 ( .A(n5300), .B(n5299), .Z(n5302) );
  AND U7807 ( .A(y[7712]), .B(x[492]), .Z(n5224) );
  NAND U7808 ( .A(y[7724]), .B(x[480]), .Z(n5223) );
  XNOR U7809 ( .A(n5224), .B(n5223), .Z(n5316) );
  AND U7810 ( .A(x[491]), .B(y[7713]), .Z(n5296) );
  XOR U7811 ( .A(o[44]), .B(n5296), .Z(n5315) );
  XOR U7812 ( .A(n5316), .B(n5315), .Z(n5285) );
  AND U7813 ( .A(y[7722]), .B(x[482]), .Z(n5226) );
  NAND U7814 ( .A(y[7716]), .B(x[488]), .Z(n5225) );
  XNOR U7815 ( .A(n5226), .B(n5225), .Z(n5290) );
  XOR U7816 ( .A(n5285), .B(n5284), .Z(n5287) );
  XOR U7817 ( .A(n5286), .B(n5287), .Z(n5280) );
  XOR U7818 ( .A(n5281), .B(n5280), .Z(n5330) );
  AND U7819 ( .A(x[491]), .B(y[7723]), .Z(n6357) );
  NAND U7820 ( .A(n6357), .B(n5512), .Z(n5230) );
  NAND U7821 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U7822 ( .A(n5230), .B(n5229), .Z(n5308) );
  AND U7823 ( .A(x[487]), .B(y[7714]), .Z(n5446) );
  AND U7824 ( .A(x[489]), .B(y[7716]), .Z(n5231) );
  NAND U7825 ( .A(n5446), .B(n5231), .Z(n5235) );
  NAND U7826 ( .A(n5233), .B(n5232), .Z(n5234) );
  NAND U7827 ( .A(n5235), .B(n5234), .Z(n5306) );
  NAND U7828 ( .A(y[7723]), .B(x[481]), .Z(n5236) );
  XNOR U7829 ( .A(n5237), .B(n5236), .Z(n5312) );
  AND U7830 ( .A(o[43]), .B(n5238), .Z(n5311) );
  XOR U7831 ( .A(n5312), .B(n5311), .Z(n5305) );
  XOR U7832 ( .A(n5306), .B(n5305), .Z(n5307) );
  XOR U7833 ( .A(n5308), .B(n5307), .Z(n5329) );
  XOR U7834 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U7835 ( .A(n5240), .B(n5239), .Z(n5244) );
  NAND U7836 ( .A(n5242), .B(n5241), .Z(n5243) );
  NAND U7837 ( .A(n5244), .B(n5243), .Z(n5335) );
  XOR U7838 ( .A(n5336), .B(n5335), .Z(n5338) );
  NANDN U7839 ( .A(n6233), .B(n5245), .Z(n5249) );
  NAND U7840 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U7841 ( .A(n5249), .B(n5248), .Z(n5273) );
  NAND U7842 ( .A(n5251), .B(n5250), .Z(n5255) );
  NANDN U7843 ( .A(n5253), .B(n5252), .Z(n5254) );
  AND U7844 ( .A(n5255), .B(n5254), .Z(n5272) );
  NANDN U7845 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U7846 ( .A(n5259), .B(n5258), .Z(n5260) );
  NAND U7847 ( .A(n5261), .B(n5260), .Z(n5275) );
  XNOR U7848 ( .A(n5338), .B(n5337), .Z(n5343) );
  NAND U7849 ( .A(n5266), .B(n5265), .Z(n5270) );
  NAND U7850 ( .A(n5268), .B(n5267), .Z(n5269) );
  AND U7851 ( .A(n5270), .B(n5269), .Z(n5341) );
  XOR U7852 ( .A(n5342), .B(n5341), .Z(n5271) );
  XNOR U7853 ( .A(n5343), .B(n5271), .Z(N109) );
  NANDN U7854 ( .A(n5273), .B(n5272), .Z(n5277) );
  NANDN U7855 ( .A(n5275), .B(n5274), .Z(n5276) );
  AND U7856 ( .A(n5277), .B(n5276), .Z(n5415) );
  NAND U7857 ( .A(n5279), .B(n5278), .Z(n5283) );
  NAND U7858 ( .A(n5281), .B(n5280), .Z(n5282) );
  NAND U7859 ( .A(n5283), .B(n5282), .Z(n5401) );
  NAND U7860 ( .A(n5285), .B(n5284), .Z(n5289) );
  NAND U7861 ( .A(n5287), .B(n5286), .Z(n5288) );
  NAND U7862 ( .A(n5289), .B(n5288), .Z(n5408) );
  AND U7863 ( .A(y[7722]), .B(x[488]), .Z(n6628) );
  AND U7864 ( .A(x[482]), .B(y[7716]), .Z(n5456) );
  NAND U7865 ( .A(n6628), .B(n5456), .Z(n5293) );
  NANDN U7866 ( .A(n5291), .B(n5290), .Z(n5292) );
  NAND U7867 ( .A(n5293), .B(n5292), .Z(n5372) );
  NAND U7868 ( .A(y[7724]), .B(x[481]), .Z(n5294) );
  XNOR U7869 ( .A(n5295), .B(n5294), .Z(n5363) );
  AND U7870 ( .A(o[44]), .B(n5296), .Z(n5362) );
  XOR U7871 ( .A(n5363), .B(n5362), .Z(n5370) );
  AND U7872 ( .A(x[486]), .B(y[7719]), .Z(n6395) );
  AND U7873 ( .A(y[7723]), .B(x[482]), .Z(n5298) );
  NAND U7874 ( .A(y[7716]), .B(x[489]), .Z(n5297) );
  XOR U7875 ( .A(n5298), .B(n5297), .Z(n5386) );
  XOR U7876 ( .A(n5370), .B(n5369), .Z(n5371) );
  XOR U7877 ( .A(n5372), .B(n5371), .Z(n5407) );
  NAND U7878 ( .A(n5300), .B(n5299), .Z(n5304) );
  ANDN U7879 ( .B(n5302), .A(n5301), .Z(n5303) );
  ANDN U7880 ( .B(n5304), .A(n5303), .Z(n5406) );
  XOR U7881 ( .A(n5407), .B(n5406), .Z(n5409) );
  XOR U7882 ( .A(n5408), .B(n5409), .Z(n5400) );
  XOR U7883 ( .A(n5401), .B(n5400), .Z(n5403) );
  NAND U7884 ( .A(n5306), .B(n5305), .Z(n5310) );
  NAND U7885 ( .A(n5308), .B(n5307), .Z(n5309) );
  NAND U7886 ( .A(n5310), .B(n5309), .Z(n5347) );
  AND U7887 ( .A(x[486]), .B(y[7723]), .Z(n5632) );
  IV U7888 ( .A(n5632), .Z(n5752) );
  AND U7889 ( .A(x[481]), .B(y[7718]), .Z(n5361) );
  NANDN U7890 ( .A(n5752), .B(n5361), .Z(n5314) );
  NAND U7891 ( .A(n5312), .B(n5311), .Z(n5313) );
  NAND U7892 ( .A(n5314), .B(n5313), .Z(n5354) );
  AND U7893 ( .A(x[492]), .B(y[7724]), .Z(n6634) );
  NAND U7894 ( .A(n6634), .B(n5512), .Z(n5318) );
  NAND U7895 ( .A(n5316), .B(n5315), .Z(n5317) );
  NAND U7896 ( .A(n5318), .B(n5317), .Z(n5352) );
  AND U7897 ( .A(x[490]), .B(y[7715]), .Z(n6245) );
  AND U7898 ( .A(y[7714]), .B(x[491]), .Z(n6206) );
  NAND U7899 ( .A(y[7717]), .B(x[488]), .Z(n5319) );
  XNOR U7900 ( .A(n6206), .B(n5319), .Z(n5358) );
  XOR U7901 ( .A(n6245), .B(n5358), .Z(n5351) );
  XOR U7902 ( .A(n5352), .B(n5351), .Z(n5353) );
  XOR U7903 ( .A(n5354), .B(n5353), .Z(n5345) );
  AND U7904 ( .A(x[490]), .B(y[7720]), .Z(n5321) );
  AND U7905 ( .A(x[484]), .B(y[7714]), .Z(n5320) );
  NAND U7906 ( .A(n5321), .B(n5320), .Z(n5324) );
  NAND U7907 ( .A(n5941), .B(n5322), .Z(n5323) );
  NAND U7908 ( .A(n5324), .B(n5323), .Z(n5396) );
  AND U7909 ( .A(y[7712]), .B(x[493]), .Z(n5326) );
  NAND U7910 ( .A(y[7725]), .B(x[480]), .Z(n5325) );
  XNOR U7911 ( .A(n5326), .B(n5325), .Z(n5380) );
  NAND U7912 ( .A(x[492]), .B(y[7713]), .Z(n5391) );
  XOR U7913 ( .A(n5380), .B(n5379), .Z(n5395) );
  AND U7914 ( .A(y[7720]), .B(x[485]), .Z(n5328) );
  NAND U7915 ( .A(y[7722]), .B(x[483]), .Z(n5327) );
  XNOR U7916 ( .A(n5328), .B(n5327), .Z(n5375) );
  AND U7917 ( .A(x[484]), .B(y[7721]), .Z(n5376) );
  XOR U7918 ( .A(n5375), .B(n5376), .Z(n5394) );
  XOR U7919 ( .A(n5395), .B(n5394), .Z(n5397) );
  XOR U7920 ( .A(n5396), .B(n5397), .Z(n5346) );
  XOR U7921 ( .A(n5345), .B(n5346), .Z(n5348) );
  XOR U7922 ( .A(n5347), .B(n5348), .Z(n5402) );
  XOR U7923 ( .A(n5403), .B(n5402), .Z(n5413) );
  NAND U7924 ( .A(n5330), .B(n5329), .Z(n5334) );
  NANDN U7925 ( .A(n5332), .B(n5331), .Z(n5333) );
  AND U7926 ( .A(n5334), .B(n5333), .Z(n5412) );
  XOR U7927 ( .A(n5415), .B(n5414), .Z(n5420) );
  NAND U7928 ( .A(n5336), .B(n5335), .Z(n5340) );
  NAND U7929 ( .A(n5338), .B(n5337), .Z(n5339) );
  NAND U7930 ( .A(n5340), .B(n5339), .Z(n5418) );
  XOR U7931 ( .A(n5418), .B(n5419), .Z(n5344) );
  XNOR U7932 ( .A(n5420), .B(n5344), .Z(N110) );
  NAND U7933 ( .A(n5346), .B(n5345), .Z(n5350) );
  NAND U7934 ( .A(n5348), .B(n5347), .Z(n5349) );
  NAND U7935 ( .A(n5350), .B(n5349), .Z(n5424) );
  NAND U7936 ( .A(n5352), .B(n5351), .Z(n5356) );
  NAND U7937 ( .A(n5354), .B(n5353), .Z(n5355) );
  AND U7938 ( .A(n5356), .B(n5355), .Z(n5431) );
  AND U7939 ( .A(y[7717]), .B(x[491]), .Z(n5538) );
  NAND U7940 ( .A(n5538), .B(n5357), .Z(n5360) );
  NAND U7941 ( .A(n5358), .B(n6245), .Z(n5359) );
  AND U7942 ( .A(n5360), .B(n5359), .Z(n5486) );
  NAND U7943 ( .A(x[487]), .B(y[7724]), .Z(n5956) );
  NANDN U7944 ( .A(n5956), .B(n5361), .Z(n5365) );
  NAND U7945 ( .A(n5363), .B(n5362), .Z(n5364) );
  NAND U7946 ( .A(n5365), .B(n5364), .Z(n5485) );
  AND U7947 ( .A(x[484]), .B(y[7722]), .Z(n5857) );
  AND U7948 ( .A(y[7723]), .B(x[483]), .Z(n5367) );
  NAND U7949 ( .A(y[7718]), .B(x[488]), .Z(n5366) );
  XOR U7950 ( .A(n5367), .B(n5366), .Z(n5471) );
  XOR U7951 ( .A(n5857), .B(n5480), .Z(n5482) );
  AND U7952 ( .A(x[489]), .B(y[7717]), .Z(n6065) );
  AND U7953 ( .A(y[7724]), .B(x[482]), .Z(n5368) );
  AND U7954 ( .A(y[7716]), .B(x[490]), .Z(n6083) );
  XOR U7955 ( .A(n5368), .B(n6083), .Z(n5457) );
  XOR U7956 ( .A(n6065), .B(n5457), .Z(n5481) );
  XOR U7957 ( .A(n5482), .B(n5481), .Z(n5487) );
  XNOR U7958 ( .A(n5488), .B(n5487), .Z(n5429) );
  NAND U7959 ( .A(n5370), .B(n5369), .Z(n5374) );
  NAND U7960 ( .A(n5372), .B(n5371), .Z(n5373) );
  AND U7961 ( .A(n5374), .B(n5373), .Z(n5428) );
  XOR U7962 ( .A(n5429), .B(n5428), .Z(n5430) );
  XNOR U7963 ( .A(n5431), .B(n5430), .Z(n5423) );
  AND U7964 ( .A(x[485]), .B(y[7722]), .Z(n5525) );
  NAND U7965 ( .A(n6233), .B(n5525), .Z(n5378) );
  NAND U7966 ( .A(n5376), .B(n5375), .Z(n5377) );
  NAND U7967 ( .A(n5378), .B(n5377), .Z(n5437) );
  AND U7968 ( .A(x[493]), .B(y[7725]), .Z(n6976) );
  NAND U7969 ( .A(n6976), .B(n5512), .Z(n5382) );
  NAND U7970 ( .A(n5380), .B(n5379), .Z(n5381) );
  NAND U7971 ( .A(n5382), .B(n5381), .Z(n5435) );
  NAND U7972 ( .A(y[7715]), .B(x[491]), .Z(n5383) );
  XNOR U7973 ( .A(n5384), .B(n5383), .Z(n5461) );
  NAND U7974 ( .A(x[481]), .B(y[7725]), .Z(n5462) );
  XOR U7975 ( .A(n5435), .B(n5434), .Z(n5436) );
  XNOR U7976 ( .A(n5437), .B(n5436), .Z(n5492) );
  AND U7977 ( .A(x[489]), .B(y[7723]), .Z(n5385) );
  NAND U7978 ( .A(n5385), .B(n5456), .Z(n5388) );
  NANDN U7979 ( .A(n5386), .B(n6395), .Z(n5387) );
  AND U7980 ( .A(n5388), .B(n5387), .Z(n5443) );
  AND U7981 ( .A(y[7712]), .B(x[494]), .Z(n5390) );
  NAND U7982 ( .A(y[7726]), .B(x[480]), .Z(n5389) );
  XNOR U7983 ( .A(n5390), .B(n5389), .Z(n5466) );
  ANDN U7984 ( .B(o[45]), .A(n5391), .Z(n5465) );
  XOR U7985 ( .A(n5466), .B(n5465), .Z(n5441) );
  NAND U7986 ( .A(y[7714]), .B(x[492]), .Z(n5392) );
  XNOR U7987 ( .A(n5393), .B(n5392), .Z(n5448) );
  NAND U7988 ( .A(x[493]), .B(y[7713]), .Z(n5455) );
  XOR U7989 ( .A(n5448), .B(n5447), .Z(n5440) );
  XOR U7990 ( .A(n5441), .B(n5440), .Z(n5442) );
  XOR U7991 ( .A(n5443), .B(n5442), .Z(n5491) );
  XOR U7992 ( .A(n5492), .B(n5491), .Z(n5494) );
  NAND U7993 ( .A(n5395), .B(n5394), .Z(n5399) );
  NAND U7994 ( .A(n5397), .B(n5396), .Z(n5398) );
  AND U7995 ( .A(n5399), .B(n5398), .Z(n5493) );
  XNOR U7996 ( .A(n5494), .B(n5493), .Z(n5422) );
  XOR U7997 ( .A(n5423), .B(n5422), .Z(n5425) );
  XOR U7998 ( .A(n5424), .B(n5425), .Z(n5500) );
  NAND U7999 ( .A(n5401), .B(n5400), .Z(n5405) );
  NAND U8000 ( .A(n5403), .B(n5402), .Z(n5404) );
  NAND U8001 ( .A(n5405), .B(n5404), .Z(n5498) );
  NAND U8002 ( .A(n5407), .B(n5406), .Z(n5411) );
  NAND U8003 ( .A(n5409), .B(n5408), .Z(n5410) );
  NAND U8004 ( .A(n5411), .B(n5410), .Z(n5497) );
  XOR U8005 ( .A(n5498), .B(n5497), .Z(n5499) );
  XOR U8006 ( .A(n5500), .B(n5499), .Z(n5505) );
  NANDN U8007 ( .A(n5413), .B(n5412), .Z(n5417) );
  NANDN U8008 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U8009 ( .A(n5417), .B(n5416), .Z(n5503) );
  XOR U8010 ( .A(n5503), .B(n5504), .Z(n5421) );
  XNOR U8011 ( .A(n5505), .B(n5421), .Z(N111) );
  NAND U8012 ( .A(n5423), .B(n5422), .Z(n5427) );
  NAND U8013 ( .A(n5425), .B(n5424), .Z(n5426) );
  NAND U8014 ( .A(n5427), .B(n5426), .Z(n5594) );
  NAND U8015 ( .A(n5429), .B(n5428), .Z(n5433) );
  NAND U8016 ( .A(n5431), .B(n5430), .Z(n5432) );
  AND U8017 ( .A(n5433), .B(n5432), .Z(n5568) );
  NAND U8018 ( .A(n5435), .B(n5434), .Z(n5439) );
  NAND U8019 ( .A(n5437), .B(n5436), .Z(n5438) );
  AND U8020 ( .A(n5439), .B(n5438), .Z(n5574) );
  NAND U8021 ( .A(n5441), .B(n5440), .Z(n5445) );
  NANDN U8022 ( .A(n5443), .B(n5442), .Z(n5444) );
  AND U8023 ( .A(n5445), .B(n5444), .Z(n5572) );
  NAND U8024 ( .A(x[492]), .B(y[7719]), .Z(n5948) );
  NANDN U8025 ( .A(n5948), .B(n5446), .Z(n5450) );
  NAND U8026 ( .A(n5448), .B(n5447), .Z(n5449) );
  AND U8027 ( .A(n5450), .B(n5449), .Z(n5548) );
  AND U8028 ( .A(y[7716]), .B(x[491]), .Z(n5452) );
  NAND U8029 ( .A(y[7714]), .B(x[493]), .Z(n5451) );
  XNOR U8030 ( .A(n5452), .B(n5451), .Z(n5552) );
  AND U8031 ( .A(x[492]), .B(y[7715]), .Z(n5551) );
  XOR U8032 ( .A(n5552), .B(n5551), .Z(n5546) );
  AND U8033 ( .A(y[7712]), .B(x[495]), .Z(n5454) );
  NAND U8034 ( .A(y[7727]), .B(x[480]), .Z(n5453) );
  XNOR U8035 ( .A(n5454), .B(n5453), .Z(n5514) );
  ANDN U8036 ( .B(o[46]), .A(n5455), .Z(n5513) );
  XNOR U8037 ( .A(n5514), .B(n5513), .Z(n5545) );
  XOR U8038 ( .A(n5548), .B(n5547), .Z(n5580) );
  NAND U8039 ( .A(x[490]), .B(y[7724]), .Z(n6397) );
  NANDN U8040 ( .A(n6397), .B(n5456), .Z(n5459) );
  NAND U8041 ( .A(n6065), .B(n5457), .Z(n5458) );
  AND U8042 ( .A(n5459), .B(n5458), .Z(n5578) );
  AND U8043 ( .A(y[7720]), .B(x[491]), .Z(n5856) );
  NAND U8044 ( .A(n5856), .B(n5460), .Z(n5464) );
  NANDN U8045 ( .A(n5462), .B(n5461), .Z(n5463) );
  NAND U8046 ( .A(n5464), .B(n5463), .Z(n5577) );
  AND U8047 ( .A(x[494]), .B(y[7726]), .Z(n7240) );
  NAND U8048 ( .A(n7240), .B(n5512), .Z(n5468) );
  NAND U8049 ( .A(n5466), .B(n5465), .Z(n5467) );
  AND U8050 ( .A(n5468), .B(n5467), .Z(n5540) );
  AND U8051 ( .A(x[488]), .B(y[7723]), .Z(n5469) );
  NAND U8052 ( .A(n5470), .B(n5469), .Z(n5473) );
  NANDN U8053 ( .A(n5471), .B(n5750), .Z(n5472) );
  NAND U8054 ( .A(n5473), .B(n5472), .Z(n5539) );
  AND U8055 ( .A(y[7717]), .B(x[490]), .Z(n5475) );
  NAND U8056 ( .A(y[7723]), .B(x[484]), .Z(n5474) );
  XNOR U8057 ( .A(n5475), .B(n5474), .Z(n5520) );
  AND U8058 ( .A(x[487]), .B(y[7720]), .Z(n5519) );
  XOR U8059 ( .A(n5520), .B(n5519), .Z(n5527) );
  NAND U8060 ( .A(x[486]), .B(y[7721]), .Z(n5663) );
  XNOR U8061 ( .A(n5663), .B(n5525), .Z(n5526) );
  AND U8062 ( .A(y[7725]), .B(x[482]), .Z(n5477) );
  NAND U8063 ( .A(y[7718]), .B(x[489]), .Z(n5476) );
  XNOR U8064 ( .A(n5477), .B(n5476), .Z(n5530) );
  NAND U8065 ( .A(x[483]), .B(y[7724]), .Z(n5531) );
  AND U8066 ( .A(y[7726]), .B(x[481]), .Z(n5479) );
  NAND U8067 ( .A(y[7719]), .B(x[488]), .Z(n5478) );
  XNOR U8068 ( .A(n5479), .B(n5478), .Z(n5509) );
  NAND U8069 ( .A(x[494]), .B(y[7713]), .Z(n5536) );
  XOR U8070 ( .A(n5509), .B(n5508), .Z(n5559) );
  XOR U8071 ( .A(n5560), .B(n5559), .Z(n5562) );
  XOR U8072 ( .A(n5561), .B(n5562), .Z(n5541) );
  XOR U8073 ( .A(n5542), .B(n5541), .Z(n5584) );
  NAND U8074 ( .A(n5857), .B(n5480), .Z(n5484) );
  NAND U8075 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U8076 ( .A(n5484), .B(n5483), .Z(n5583) );
  NANDN U8077 ( .A(n5486), .B(n5485), .Z(n5490) );
  NAND U8078 ( .A(n5488), .B(n5487), .Z(n5489) );
  NAND U8079 ( .A(n5490), .B(n5489), .Z(n5586) );
  XOR U8080 ( .A(n5565), .B(n5566), .Z(n5567) );
  NAND U8081 ( .A(n5492), .B(n5491), .Z(n5496) );
  NAND U8082 ( .A(n5494), .B(n5493), .Z(n5495) );
  AND U8083 ( .A(n5496), .B(n5495), .Z(n5592) );
  XNOR U8084 ( .A(n5593), .B(n5592), .Z(n5595) );
  XOR U8085 ( .A(n5594), .B(n5595), .Z(n5591) );
  NAND U8086 ( .A(n5498), .B(n5497), .Z(n5502) );
  NAND U8087 ( .A(n5500), .B(n5499), .Z(n5501) );
  NAND U8088 ( .A(n5502), .B(n5501), .Z(n5590) );
  XOR U8089 ( .A(n5590), .B(n5589), .Z(n5506) );
  XNOR U8090 ( .A(n5591), .B(n5506), .Z(N112) );
  AND U8091 ( .A(x[488]), .B(y[7726]), .Z(n5858) );
  NAND U8092 ( .A(n5858), .B(n5507), .Z(n5511) );
  NAND U8093 ( .A(n5509), .B(n5508), .Z(n5510) );
  AND U8094 ( .A(n5511), .B(n5510), .Z(n5612) );
  AND U8095 ( .A(x[495]), .B(y[7727]), .Z(n7566) );
  NAND U8096 ( .A(n7566), .B(n5512), .Z(n5516) );
  NAND U8097 ( .A(n5514), .B(n5513), .Z(n5515) );
  NAND U8098 ( .A(n5516), .B(n5515), .Z(n5611) );
  AND U8099 ( .A(x[490]), .B(y[7723]), .Z(n5518) );
  NAND U8100 ( .A(n5518), .B(n5517), .Z(n5522) );
  NAND U8101 ( .A(n5520), .B(n5519), .Z(n5521) );
  NAND U8102 ( .A(n5522), .B(n5521), .Z(n5649) );
  AND U8103 ( .A(x[480]), .B(y[7728]), .Z(n5672) );
  NAND U8104 ( .A(x[496]), .B(y[7712]), .Z(n5673) );
  NAND U8105 ( .A(x[495]), .B(y[7713]), .Z(n5659) );
  XOR U8106 ( .A(n5675), .B(n5674), .Z(n5648) );
  NAND U8107 ( .A(y[7721]), .B(x[487]), .Z(n5523) );
  XNOR U8108 ( .A(n5524), .B(n5523), .Z(n5665) );
  AND U8109 ( .A(x[490]), .B(y[7718]), .Z(n5664) );
  XOR U8110 ( .A(n5665), .B(n5664), .Z(n5647) );
  XOR U8111 ( .A(n5648), .B(n5647), .Z(n5650) );
  XOR U8112 ( .A(n5649), .B(n5650), .Z(n5613) );
  XOR U8113 ( .A(n5614), .B(n5613), .Z(n5644) );
  NANDN U8114 ( .A(n5525), .B(n5663), .Z(n5529) );
  NANDN U8115 ( .A(n5527), .B(n5526), .Z(n5528) );
  AND U8116 ( .A(n5529), .B(n5528), .Z(n5642) );
  NAND U8117 ( .A(x[489]), .B(y[7725]), .Z(n6378) );
  NANDN U8118 ( .A(n6378), .B(n5946), .Z(n5533) );
  NANDN U8119 ( .A(n5531), .B(n5530), .Z(n5532) );
  AND U8120 ( .A(n5533), .B(n5532), .Z(n5683) );
  AND U8121 ( .A(y[7727]), .B(x[481]), .Z(n5535) );
  NAND U8122 ( .A(y[7720]), .B(x[488]), .Z(n5534) );
  XNOR U8123 ( .A(n5535), .B(n5534), .Z(n5669) );
  ANDN U8124 ( .B(o[47]), .A(n5536), .Z(n5668) );
  XOR U8125 ( .A(n5669), .B(n5668), .Z(n5681) );
  NAND U8126 ( .A(y[7714]), .B(x[494]), .Z(n5537) );
  XNOR U8127 ( .A(n5538), .B(n5537), .Z(n5623) );
  NAND U8128 ( .A(x[484]), .B(y[7724]), .Z(n5624) );
  XOR U8129 ( .A(n5681), .B(n5680), .Z(n5682) );
  XOR U8130 ( .A(n5683), .B(n5682), .Z(n5641) );
  NANDN U8131 ( .A(n5540), .B(n5539), .Z(n5544) );
  NAND U8132 ( .A(n5542), .B(n5541), .Z(n5543) );
  NAND U8133 ( .A(n5544), .B(n5543), .Z(n5606) );
  NANDN U8134 ( .A(n5546), .B(n5545), .Z(n5550) );
  NAND U8135 ( .A(n5548), .B(n5547), .Z(n5549) );
  AND U8136 ( .A(n5550), .B(n5549), .Z(n5638) );
  AND U8137 ( .A(y[7716]), .B(x[493]), .Z(n5634) );
  NAND U8138 ( .A(n6206), .B(n5634), .Z(n5554) );
  NAND U8139 ( .A(n5552), .B(n5551), .Z(n5553) );
  AND U8140 ( .A(n5554), .B(n5553), .Z(n5620) );
  AND U8141 ( .A(y[7726]), .B(x[482]), .Z(n5556) );
  NAND U8142 ( .A(y[7719]), .B(x[489]), .Z(n5555) );
  XNOR U8143 ( .A(n5556), .B(n5555), .Z(n5627) );
  NAND U8144 ( .A(x[483]), .B(y[7725]), .Z(n5628) );
  AND U8145 ( .A(x[492]), .B(y[7716]), .Z(n6366) );
  AND U8146 ( .A(y[7723]), .B(x[485]), .Z(n5558) );
  NAND U8147 ( .A(y[7715]), .B(x[493]), .Z(n5557) );
  XOR U8148 ( .A(n5558), .B(n5557), .Z(n5654) );
  XOR U8149 ( .A(n5618), .B(n5617), .Z(n5619) );
  NAND U8150 ( .A(n5560), .B(n5559), .Z(n5564) );
  NAND U8151 ( .A(n5562), .B(n5561), .Z(n5563) );
  AND U8152 ( .A(n5564), .B(n5563), .Z(n5636) );
  XOR U8153 ( .A(n5635), .B(n5636), .Z(n5637) );
  XOR U8154 ( .A(n5608), .B(n5607), .Z(n5687) );
  NAND U8155 ( .A(n5566), .B(n5565), .Z(n5570) );
  NANDN U8156 ( .A(n5568), .B(n5567), .Z(n5569) );
  AND U8157 ( .A(n5570), .B(n5569), .Z(n5686) );
  NANDN U8158 ( .A(n5572), .B(n5571), .Z(n5576) );
  NANDN U8159 ( .A(n5574), .B(n5573), .Z(n5575) );
  AND U8160 ( .A(n5576), .B(n5575), .Z(n5602) );
  NANDN U8161 ( .A(n5578), .B(n5577), .Z(n5582) );
  NANDN U8162 ( .A(n5580), .B(n5579), .Z(n5581) );
  AND U8163 ( .A(n5582), .B(n5581), .Z(n5600) );
  NANDN U8164 ( .A(n5584), .B(n5583), .Z(n5588) );
  NANDN U8165 ( .A(n5586), .B(n5585), .Z(n5587) );
  AND U8166 ( .A(n5588), .B(n5587), .Z(n5599) );
  XNOR U8167 ( .A(n5689), .B(n5688), .Z(n5694) );
  NAND U8168 ( .A(n5593), .B(n5592), .Z(n5597) );
  NANDN U8169 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U8170 ( .A(n5597), .B(n5596), .Z(n5692) );
  XNOR U8171 ( .A(n5693), .B(n5692), .Z(n5598) );
  XNOR U8172 ( .A(n5694), .B(n5598), .Z(N113) );
  NANDN U8173 ( .A(n5600), .B(n5599), .Z(n5604) );
  NANDN U8174 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U8175 ( .A(n5604), .B(n5603), .Z(n5796) );
  NANDN U8176 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U8177 ( .A(n5608), .B(n5607), .Z(n5609) );
  AND U8178 ( .A(n5610), .B(n5609), .Z(n5699) );
  NANDN U8179 ( .A(n5612), .B(n5611), .Z(n5616) );
  NAND U8180 ( .A(n5614), .B(n5613), .Z(n5615) );
  AND U8181 ( .A(n5616), .B(n5615), .Z(n5781) );
  NAND U8182 ( .A(n5618), .B(n5617), .Z(n5622) );
  NANDN U8183 ( .A(n5620), .B(n5619), .Z(n5621) );
  AND U8184 ( .A(n5622), .B(n5621), .Z(n5779) );
  NAND U8185 ( .A(x[494]), .B(y[7717]), .Z(n5980) );
  NANDN U8186 ( .A(n5980), .B(n6206), .Z(n5626) );
  NANDN U8187 ( .A(n5624), .B(n5623), .Z(n5625) );
  AND U8188 ( .A(n5626), .B(n5625), .Z(n5773) );
  AND U8189 ( .A(x[489]), .B(y[7726]), .Z(n6623) );
  NANDN U8190 ( .A(n5759), .B(n6623), .Z(n5630) );
  NANDN U8191 ( .A(n5628), .B(n5627), .Z(n5629) );
  NAND U8192 ( .A(n5630), .B(n5629), .Z(n5772) );
  AND U8193 ( .A(x[485]), .B(y[7724]), .Z(n5818) );
  NAND U8194 ( .A(y[7721]), .B(x[488]), .Z(n5631) );
  XNOR U8195 ( .A(n5818), .B(n5631), .Z(n5751) );
  XOR U8196 ( .A(n5751), .B(n5632), .Z(n5766) );
  NAND U8197 ( .A(x[487]), .B(y[7722]), .Z(n5767) );
  IV U8198 ( .A(n5767), .Z(n5662) );
  XOR U8199 ( .A(n5766), .B(n5662), .Z(n5769) );
  NAND U8200 ( .A(y[7725]), .B(x[484]), .Z(n5633) );
  XNOR U8201 ( .A(n5634), .B(n5633), .Z(n5713) );
  NAND U8202 ( .A(x[491]), .B(y[7718]), .Z(n5714) );
  XOR U8203 ( .A(n5769), .B(n5768), .Z(n5774) );
  XOR U8204 ( .A(n5775), .B(n5774), .Z(n5778) );
  NAND U8205 ( .A(n5636), .B(n5635), .Z(n5640) );
  NANDN U8206 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U8207 ( .A(n5640), .B(n5639), .Z(n5696) );
  XOR U8208 ( .A(n5697), .B(n5696), .Z(n5698) );
  NANDN U8209 ( .A(n5642), .B(n5641), .Z(n5646) );
  NANDN U8210 ( .A(n5644), .B(n5643), .Z(n5645) );
  AND U8211 ( .A(n5646), .B(n5645), .Z(n5705) );
  NAND U8212 ( .A(n5648), .B(n5647), .Z(n5652) );
  NAND U8213 ( .A(n5650), .B(n5649), .Z(n5651) );
  AND U8214 ( .A(n5652), .B(n5651), .Z(n5787) );
  AND U8215 ( .A(x[493]), .B(y[7723]), .Z(n6642) );
  NAND U8216 ( .A(n6642), .B(n5653), .Z(n5656) );
  NANDN U8217 ( .A(n5654), .B(n6366), .Z(n5655) );
  AND U8218 ( .A(n5656), .B(n5655), .Z(n5735) );
  AND U8219 ( .A(y[7728]), .B(x[481]), .Z(n5658) );
  NAND U8220 ( .A(y[7720]), .B(x[489]), .Z(n5657) );
  XNOR U8221 ( .A(n5658), .B(n5657), .Z(n5756) );
  ANDN U8222 ( .B(o[48]), .A(n5659), .Z(n5755) );
  XOR U8223 ( .A(n5756), .B(n5755), .Z(n5733) );
  AND U8224 ( .A(y[7714]), .B(x[495]), .Z(n5661) );
  NAND U8225 ( .A(y[7717]), .B(x[492]), .Z(n5660) );
  XNOR U8226 ( .A(n5661), .B(n5660), .Z(n5709) );
  AND U8227 ( .A(x[494]), .B(y[7715]), .Z(n5708) );
  XOR U8228 ( .A(n5709), .B(n5708), .Z(n5732) );
  XOR U8229 ( .A(n5733), .B(n5732), .Z(n5734) );
  NANDN U8230 ( .A(n5663), .B(n5662), .Z(n5667) );
  NAND U8231 ( .A(n5665), .B(n5664), .Z(n5666) );
  AND U8232 ( .A(n5667), .B(n5666), .Z(n5745) );
  NAND U8233 ( .A(x[488]), .B(y[7727]), .Z(n6447) );
  AND U8234 ( .A(x[481]), .B(y[7720]), .Z(n5836) );
  NANDN U8235 ( .A(n6447), .B(n5836), .Z(n5671) );
  NAND U8236 ( .A(n5669), .B(n5668), .Z(n5670) );
  NAND U8237 ( .A(n5671), .B(n5670), .Z(n5744) );
  NANDN U8238 ( .A(n5673), .B(n5672), .Z(n5677) );
  NAND U8239 ( .A(n5675), .B(n5674), .Z(n5676) );
  AND U8240 ( .A(n5677), .B(n5676), .Z(n5741) );
  AND U8241 ( .A(x[480]), .B(y[7729]), .Z(n5723) );
  AND U8242 ( .A(x[497]), .B(y[7712]), .Z(n5722) );
  XOR U8243 ( .A(n5723), .B(n5722), .Z(n5725) );
  AND U8244 ( .A(x[496]), .B(y[7713]), .Z(n5719) );
  XOR U8245 ( .A(n5719), .B(o[49]), .Z(n5724) );
  XOR U8246 ( .A(n5725), .B(n5724), .Z(n5739) );
  AND U8247 ( .A(y[7727]), .B(x[482]), .Z(n5679) );
  NAND U8248 ( .A(y[7719]), .B(x[490]), .Z(n5678) );
  XNOR U8249 ( .A(n5679), .B(n5678), .Z(n5760) );
  NAND U8250 ( .A(x[483]), .B(y[7726]), .Z(n5761) );
  XOR U8251 ( .A(n5739), .B(n5738), .Z(n5740) );
  XOR U8252 ( .A(n5747), .B(n5746), .Z(n5784) );
  XOR U8253 ( .A(n5785), .B(n5784), .Z(n5786) );
  NAND U8254 ( .A(n5681), .B(n5680), .Z(n5685) );
  NANDN U8255 ( .A(n5683), .B(n5682), .Z(n5684) );
  AND U8256 ( .A(n5685), .B(n5684), .Z(n5703) );
  XOR U8257 ( .A(n5702), .B(n5703), .Z(n5704) );
  XOR U8258 ( .A(n5705), .B(n5704), .Z(n5793) );
  XOR U8259 ( .A(n5794), .B(n5793), .Z(n5795) );
  XOR U8260 ( .A(n5796), .B(n5795), .Z(n5792) );
  NANDN U8261 ( .A(n5687), .B(n5686), .Z(n5691) );
  NAND U8262 ( .A(n5689), .B(n5688), .Z(n5690) );
  NAND U8263 ( .A(n5691), .B(n5690), .Z(n5790) );
  XOR U8264 ( .A(n5790), .B(n5791), .Z(n5695) );
  XNOR U8265 ( .A(n5792), .B(n5695), .Z(N114) );
  NAND U8266 ( .A(n5697), .B(n5696), .Z(n5701) );
  NANDN U8267 ( .A(n5699), .B(n5698), .Z(n5700) );
  AND U8268 ( .A(n5701), .B(n5700), .Z(n5912) );
  NAND U8269 ( .A(n5703), .B(n5702), .Z(n5707) );
  NANDN U8270 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U8271 ( .A(n5707), .B(n5706), .Z(n5910) );
  AND U8272 ( .A(x[492]), .B(y[7714]), .Z(n6055) );
  AND U8273 ( .A(x[495]), .B(y[7717]), .Z(n5954) );
  NAND U8274 ( .A(n6055), .B(n5954), .Z(n5711) );
  NAND U8275 ( .A(n5709), .B(n5708), .Z(n5710) );
  NAND U8276 ( .A(n5711), .B(n5710), .Z(n5884) );
  NAND U8277 ( .A(n6976), .B(n5712), .Z(n5716) );
  NANDN U8278 ( .A(n5714), .B(n5713), .Z(n5715) );
  AND U8279 ( .A(n5716), .B(n5715), .Z(n5875) );
  AND U8280 ( .A(y[7729]), .B(x[481]), .Z(n5718) );
  NAND U8281 ( .A(y[7720]), .B(x[490]), .Z(n5717) );
  XNOR U8282 ( .A(n5718), .B(n5717), .Z(n5837) );
  NAND U8283 ( .A(n5719), .B(o[49]), .Z(n5838) );
  AND U8284 ( .A(y[7715]), .B(x[495]), .Z(n5721) );
  NAND U8285 ( .A(y[7721]), .B(x[489]), .Z(n5720) );
  XNOR U8286 ( .A(n5721), .B(n5720), .Z(n5828) );
  NAND U8287 ( .A(x[494]), .B(y[7716]), .Z(n5829) );
  XOR U8288 ( .A(n5873), .B(n5872), .Z(n5874) );
  XOR U8289 ( .A(n5884), .B(n5885), .Z(n5887) );
  NAND U8290 ( .A(n5723), .B(n5722), .Z(n5727) );
  NAND U8291 ( .A(n5725), .B(n5724), .Z(n5726) );
  NAND U8292 ( .A(n5727), .B(n5726), .Z(n5896) );
  AND U8293 ( .A(y[7714]), .B(x[496]), .Z(n5729) );
  NAND U8294 ( .A(y[7719]), .B(x[491]), .Z(n5728) );
  XNOR U8295 ( .A(n5729), .B(n5728), .Z(n5824) );
  NAND U8296 ( .A(x[482]), .B(y[7728]), .Z(n5825) );
  XOR U8297 ( .A(n5896), .B(n5897), .Z(n5899) );
  AND U8298 ( .A(x[485]), .B(y[7725]), .Z(n5962) );
  NAND U8299 ( .A(y[7724]), .B(x[486]), .Z(n5730) );
  XNOR U8300 ( .A(n5962), .B(n5730), .Z(n5821) );
  NAND U8301 ( .A(y[7726]), .B(x[484]), .Z(n5731) );
  XNOR U8302 ( .A(n6628), .B(n5731), .Z(n5859) );
  NAND U8303 ( .A(x[487]), .B(y[7723]), .Z(n5860) );
  XOR U8304 ( .A(n5821), .B(n5820), .Z(n5898) );
  XOR U8305 ( .A(n5899), .B(n5898), .Z(n5886) );
  XOR U8306 ( .A(n5887), .B(n5886), .Z(n5807) );
  NAND U8307 ( .A(n5733), .B(n5732), .Z(n5737) );
  NANDN U8308 ( .A(n5735), .B(n5734), .Z(n5736) );
  AND U8309 ( .A(n5737), .B(n5736), .Z(n5879) );
  NAND U8310 ( .A(n5739), .B(n5738), .Z(n5743) );
  NANDN U8311 ( .A(n5741), .B(n5740), .Z(n5742) );
  AND U8312 ( .A(n5743), .B(n5742), .Z(n5878) );
  XOR U8313 ( .A(n5879), .B(n5878), .Z(n5881) );
  NANDN U8314 ( .A(n5745), .B(n5744), .Z(n5749) );
  NAND U8315 ( .A(n5747), .B(n5746), .Z(n5748) );
  AND U8316 ( .A(n5749), .B(n5748), .Z(n5880) );
  XOR U8317 ( .A(n5881), .B(n5880), .Z(n5806) );
  AND U8318 ( .A(x[488]), .B(y[7724]), .Z(n6090) );
  NAND U8319 ( .A(n6090), .B(n5750), .Z(n5754) );
  NANDN U8320 ( .A(n5752), .B(n5751), .Z(n5753) );
  NAND U8321 ( .A(n5754), .B(n5753), .Z(n5891) );
  AND U8322 ( .A(x[489]), .B(y[7728]), .Z(n6734) );
  NAND U8323 ( .A(n6734), .B(n5836), .Z(n5758) );
  NAND U8324 ( .A(n5756), .B(n5755), .Z(n5757) );
  NAND U8325 ( .A(n5758), .B(n5757), .Z(n5890) );
  XOR U8326 ( .A(n5891), .B(n5890), .Z(n5893) );
  AND U8327 ( .A(x[490]), .B(y[7727]), .Z(n6651) );
  NANDN U8328 ( .A(n5759), .B(n6651), .Z(n5763) );
  NANDN U8329 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U8330 ( .A(n5763), .B(n5762), .Z(n5869) );
  AND U8331 ( .A(x[480]), .B(y[7730]), .Z(n5841) );
  NAND U8332 ( .A(x[498]), .B(y[7712]), .Z(n5842) );
  NAND U8333 ( .A(x[497]), .B(y[7713]), .Z(n5863) );
  XOR U8334 ( .A(n5844), .B(n5843), .Z(n5867) );
  AND U8335 ( .A(y[7717]), .B(x[493]), .Z(n5765) );
  NAND U8336 ( .A(y[7727]), .B(x[483]), .Z(n5764) );
  XNOR U8337 ( .A(n5765), .B(n5764), .Z(n5849) );
  NAND U8338 ( .A(x[492]), .B(y[7718]), .Z(n5850) );
  XOR U8339 ( .A(n5867), .B(n5866), .Z(n5868) );
  XOR U8340 ( .A(n5893), .B(n5892), .Z(n5813) );
  NANDN U8341 ( .A(n5767), .B(n5766), .Z(n5771) );
  NAND U8342 ( .A(n5769), .B(n5768), .Z(n5770) );
  AND U8343 ( .A(n5771), .B(n5770), .Z(n5812) );
  NANDN U8344 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U8345 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U8346 ( .A(n5777), .B(n5776), .Z(n5815) );
  XOR U8347 ( .A(n5809), .B(n5808), .Z(n5803) );
  NANDN U8348 ( .A(n5779), .B(n5778), .Z(n5783) );
  NANDN U8349 ( .A(n5781), .B(n5780), .Z(n5782) );
  AND U8350 ( .A(n5783), .B(n5782), .Z(n5801) );
  NAND U8351 ( .A(n5785), .B(n5784), .Z(n5789) );
  NANDN U8352 ( .A(n5787), .B(n5786), .Z(n5788) );
  NAND U8353 ( .A(n5789), .B(n5788), .Z(n5800) );
  XOR U8354 ( .A(n5910), .B(n5909), .Z(n5911) );
  XNOR U8355 ( .A(n5912), .B(n5911), .Z(n5905) );
  NAND U8356 ( .A(n5794), .B(n5793), .Z(n5798) );
  NANDN U8357 ( .A(n5796), .B(n5795), .Z(n5797) );
  NAND U8358 ( .A(n5798), .B(n5797), .Z(n5903) );
  IV U8359 ( .A(n5903), .Z(n5902) );
  XOR U8360 ( .A(n5904), .B(n5902), .Z(n5799) );
  XNOR U8361 ( .A(n5905), .B(n5799), .Z(N115) );
  NANDN U8362 ( .A(n5801), .B(n5800), .Z(n5805) );
  NANDN U8363 ( .A(n5803), .B(n5802), .Z(n5804) );
  AND U8364 ( .A(n5805), .B(n5804), .Z(n5919) );
  NANDN U8365 ( .A(n5807), .B(n5806), .Z(n5811) );
  NAND U8366 ( .A(n5809), .B(n5808), .Z(n5810) );
  AND U8367 ( .A(n5811), .B(n5810), .Z(n5917) );
  NANDN U8368 ( .A(n5813), .B(n5812), .Z(n5817) );
  NANDN U8369 ( .A(n5815), .B(n5814), .Z(n5816) );
  AND U8370 ( .A(n5817), .B(n5816), .Z(n6021) );
  AND U8371 ( .A(x[486]), .B(y[7725]), .Z(n5819) );
  NAND U8372 ( .A(n5819), .B(n5818), .Z(n5823) );
  NAND U8373 ( .A(n5821), .B(n5820), .Z(n5822) );
  AND U8374 ( .A(n5823), .B(n5822), .Z(n6015) );
  AND U8375 ( .A(x[496]), .B(y[7719]), .Z(n6382) );
  NAND U8376 ( .A(n6382), .B(n6206), .Z(n5827) );
  NANDN U8377 ( .A(n5825), .B(n5824), .Z(n5826) );
  AND U8378 ( .A(n5827), .B(n5826), .Z(n6013) );
  AND U8379 ( .A(x[495]), .B(y[7721]), .Z(n6654) );
  NAND U8380 ( .A(n6654), .B(n5941), .Z(n5831) );
  NANDN U8381 ( .A(n5829), .B(n5828), .Z(n5830) );
  AND U8382 ( .A(n5831), .B(n5830), .Z(n5932) );
  AND U8383 ( .A(y[7730]), .B(x[481]), .Z(n5833) );
  NAND U8384 ( .A(y[7723]), .B(x[488]), .Z(n5832) );
  XNOR U8385 ( .A(n5833), .B(n5832), .Z(n5979) );
  AND U8386 ( .A(y[7718]), .B(x[493]), .Z(n5835) );
  NAND U8387 ( .A(y[7729]), .B(x[482]), .Z(n5834) );
  XNOR U8388 ( .A(n5835), .B(n5834), .Z(n5947) );
  XOR U8389 ( .A(n5930), .B(n5929), .Z(n5931) );
  AND U8390 ( .A(x[490]), .B(y[7729]), .Z(n7058) );
  NAND U8391 ( .A(n7058), .B(n5836), .Z(n5840) );
  NANDN U8392 ( .A(n5838), .B(n5837), .Z(n5839) );
  AND U8393 ( .A(n5840), .B(n5839), .Z(n5991) );
  NANDN U8394 ( .A(n5842), .B(n5841), .Z(n5846) );
  NAND U8395 ( .A(n5844), .B(n5843), .Z(n5845) );
  AND U8396 ( .A(n5846), .B(n5845), .Z(n5989) );
  AND U8397 ( .A(y[7715]), .B(x[496]), .Z(n6592) );
  NAND U8398 ( .A(y[7722]), .B(x[489]), .Z(n5847) );
  XNOR U8399 ( .A(n6592), .B(n5847), .Z(n5942) );
  NAND U8400 ( .A(x[495]), .B(y[7716]), .Z(n5943) );
  AND U8401 ( .A(x[493]), .B(y[7727]), .Z(n7267) );
  NANDN U8402 ( .A(n5848), .B(n7267), .Z(n5852) );
  NANDN U8403 ( .A(n5850), .B(n5849), .Z(n5851) );
  AND U8404 ( .A(n5852), .B(n5851), .Z(n5997) );
  AND U8405 ( .A(y[7721]), .B(x[490]), .Z(n5854) );
  NAND U8406 ( .A(y[7714]), .B(x[497]), .Z(n5853) );
  XNOR U8407 ( .A(n5854), .B(n5853), .Z(n5985) );
  AND U8408 ( .A(x[498]), .B(y[7713]), .Z(n5961) );
  XOR U8409 ( .A(o[51]), .B(n5961), .Z(n5984) );
  XOR U8410 ( .A(n5985), .B(n5984), .Z(n5995) );
  NAND U8411 ( .A(y[7728]), .B(x[483]), .Z(n5855) );
  XNOR U8412 ( .A(n5856), .B(n5855), .Z(n5955) );
  XOR U8413 ( .A(n5995), .B(n5994), .Z(n5996) );
  NAND U8414 ( .A(n5858), .B(n5857), .Z(n5862) );
  NANDN U8415 ( .A(n5860), .B(n5859), .Z(n5861) );
  AND U8416 ( .A(n5862), .B(n5861), .Z(n5938) );
  AND U8417 ( .A(x[480]), .B(y[7731]), .Z(n5966) );
  NAND U8418 ( .A(x[499]), .B(y[7712]), .Z(n5967) );
  ANDN U8419 ( .B(o[50]), .A(n5863), .Z(n5968) );
  XOR U8420 ( .A(n5969), .B(n5968), .Z(n5936) );
  AND U8421 ( .A(x[484]), .B(y[7727]), .Z(n6103) );
  AND U8422 ( .A(y[7726]), .B(x[485]), .Z(n5865) );
  NAND U8423 ( .A(y[7725]), .B(x[486]), .Z(n5864) );
  XOR U8424 ( .A(n5865), .B(n5864), .Z(n5963) );
  XOR U8425 ( .A(n5936), .B(n5935), .Z(n5937) );
  XOR U8426 ( .A(n5938), .B(n5937), .Z(n6006) );
  XOR U8427 ( .A(n6007), .B(n6006), .Z(n6009) );
  XNOR U8428 ( .A(n6008), .B(n6009), .Z(n6002) );
  NAND U8429 ( .A(n5867), .B(n5866), .Z(n5871) );
  NANDN U8430 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U8431 ( .A(n5871), .B(n5870), .Z(n6001) );
  NAND U8432 ( .A(n5873), .B(n5872), .Z(n5877) );
  NANDN U8433 ( .A(n5875), .B(n5874), .Z(n5876) );
  NAND U8434 ( .A(n5877), .B(n5876), .Z(n6000) );
  XNOR U8435 ( .A(n6002), .B(n6003), .Z(n6018) );
  XOR U8436 ( .A(n6019), .B(n6018), .Z(n6020) );
  NAND U8437 ( .A(n5879), .B(n5878), .Z(n5883) );
  NAND U8438 ( .A(n5881), .B(n5880), .Z(n5882) );
  AND U8439 ( .A(n5883), .B(n5882), .Z(n6030) );
  NAND U8440 ( .A(n5885), .B(n5884), .Z(n5889) );
  NAND U8441 ( .A(n5887), .B(n5886), .Z(n5888) );
  NAND U8442 ( .A(n5889), .B(n5888), .Z(n6026) );
  NAND U8443 ( .A(n5891), .B(n5890), .Z(n5895) );
  NAND U8444 ( .A(n5893), .B(n5892), .Z(n5894) );
  NAND U8445 ( .A(n5895), .B(n5894), .Z(n6025) );
  NAND U8446 ( .A(n5897), .B(n5896), .Z(n5901) );
  NAND U8447 ( .A(n5899), .B(n5898), .Z(n5900) );
  NAND U8448 ( .A(n5901), .B(n5900), .Z(n6024) );
  XNOR U8449 ( .A(n6025), .B(n6024), .Z(n6027) );
  XNOR U8450 ( .A(n6030), .B(n6031), .Z(n6032) );
  XOR U8451 ( .A(n5917), .B(n5916), .Z(n5918) );
  XOR U8452 ( .A(n5919), .B(n5918), .Z(n5925) );
  OR U8453 ( .A(n5904), .B(n5902), .Z(n5908) );
  ANDN U8454 ( .B(n5904), .A(n5903), .Z(n5906) );
  OR U8455 ( .A(n5906), .B(n5905), .Z(n5907) );
  AND U8456 ( .A(n5908), .B(n5907), .Z(n5924) );
  NAND U8457 ( .A(n5910), .B(n5909), .Z(n5914) );
  NAND U8458 ( .A(n5912), .B(n5911), .Z(n5913) );
  NAND U8459 ( .A(n5914), .B(n5913), .Z(n5923) );
  IV U8460 ( .A(n5923), .Z(n5922) );
  XOR U8461 ( .A(n5924), .B(n5922), .Z(n5915) );
  XNOR U8462 ( .A(n5925), .B(n5915), .Z(N116) );
  NAND U8463 ( .A(n5917), .B(n5916), .Z(n5921) );
  NANDN U8464 ( .A(n5919), .B(n5918), .Z(n5920) );
  NAND U8465 ( .A(n5921), .B(n5920), .Z(n6151) );
  IV U8466 ( .A(n6151), .Z(n6150) );
  OR U8467 ( .A(n5924), .B(n5922), .Z(n5928) );
  ANDN U8468 ( .B(n5924), .A(n5923), .Z(n5926) );
  OR U8469 ( .A(n5926), .B(n5925), .Z(n5927) );
  AND U8470 ( .A(n5928), .B(n5927), .Z(n6152) );
  NAND U8471 ( .A(n5930), .B(n5929), .Z(n5934) );
  NANDN U8472 ( .A(n5932), .B(n5931), .Z(n5933) );
  AND U8473 ( .A(n5934), .B(n5933), .Z(n6038) );
  NAND U8474 ( .A(n5936), .B(n5935), .Z(n5940) );
  NANDN U8475 ( .A(n5938), .B(n5937), .Z(n5939) );
  NAND U8476 ( .A(n5940), .B(n5939), .Z(n6037) );
  AND U8477 ( .A(x[496]), .B(y[7722]), .Z(n6933) );
  NAND U8478 ( .A(n6933), .B(n5941), .Z(n5945) );
  NANDN U8479 ( .A(n5943), .B(n5942), .Z(n5944) );
  AND U8480 ( .A(n5945), .B(n5944), .Z(n6078) );
  AND U8481 ( .A(x[493]), .B(y[7729]), .Z(n7507) );
  NAND U8482 ( .A(n7507), .B(n5946), .Z(n5950) );
  NANDN U8483 ( .A(n5948), .B(n5947), .Z(n5949) );
  AND U8484 ( .A(n5950), .B(n5949), .Z(n6123) );
  AND U8485 ( .A(y[7716]), .B(x[496]), .Z(n5952) );
  NAND U8486 ( .A(y[7722]), .B(x[490]), .Z(n5951) );
  XNOR U8487 ( .A(n5952), .B(n5951), .Z(n6084) );
  AND U8488 ( .A(x[482]), .B(y[7730]), .Z(n6085) );
  XOR U8489 ( .A(n6084), .B(n6085), .Z(n6121) );
  NAND U8490 ( .A(y[7723]), .B(x[489]), .Z(n5953) );
  XNOR U8491 ( .A(n5954), .B(n5953), .Z(n6066) );
  AND U8492 ( .A(x[494]), .B(y[7718]), .Z(n6067) );
  XOR U8493 ( .A(n6066), .B(n6067), .Z(n6120) );
  XOR U8494 ( .A(n6121), .B(n6120), .Z(n6122) );
  AND U8495 ( .A(x[491]), .B(y[7728]), .Z(n7060) );
  IV U8496 ( .A(n7060), .Z(n6895) );
  NANDN U8497 ( .A(n6895), .B(n6233), .Z(n5958) );
  NANDN U8498 ( .A(n5956), .B(n5955), .Z(n5957) );
  AND U8499 ( .A(n5958), .B(n5957), .Z(n6129) );
  AND U8500 ( .A(y[7721]), .B(x[491]), .Z(n5960) );
  NAND U8501 ( .A(y[7731]), .B(x[481]), .Z(n5959) );
  XNOR U8502 ( .A(n5960), .B(n5959), .Z(n6062) );
  AND U8503 ( .A(x[499]), .B(y[7713]), .Z(n6070) );
  XOR U8504 ( .A(o[52]), .B(n6070), .Z(n6061) );
  XOR U8505 ( .A(n6062), .B(n6061), .Z(n6127) );
  AND U8506 ( .A(o[51]), .B(n5961), .Z(n6111) );
  AND U8507 ( .A(x[480]), .B(y[7732]), .Z(n6108) );
  AND U8508 ( .A(x[500]), .B(y[7712]), .Z(n6109) );
  XOR U8509 ( .A(n6108), .B(n6109), .Z(n6110) );
  XOR U8510 ( .A(n6111), .B(n6110), .Z(n6126) );
  XOR U8511 ( .A(n6127), .B(n6126), .Z(n6128) );
  XOR U8512 ( .A(n6080), .B(n6079), .Z(n6039) );
  XOR U8513 ( .A(n6040), .B(n6039), .Z(n6135) );
  NAND U8514 ( .A(x[486]), .B(y[7726]), .Z(n6071) );
  NANDN U8515 ( .A(n6071), .B(n5962), .Z(n5965) );
  NANDN U8516 ( .A(n5963), .B(n6103), .Z(n5964) );
  AND U8517 ( .A(n5965), .B(n5964), .Z(n6052) );
  NANDN U8518 ( .A(n5967), .B(n5966), .Z(n5971) );
  NAND U8519 ( .A(n5969), .B(n5968), .Z(n5970) );
  AND U8520 ( .A(n5971), .B(n5970), .Z(n6050) );
  AND U8521 ( .A(y[7714]), .B(x[498]), .Z(n5973) );
  NAND U8522 ( .A(y[7720]), .B(x[492]), .Z(n5972) );
  XNOR U8523 ( .A(n5973), .B(n5972), .Z(n6056) );
  AND U8524 ( .A(x[497]), .B(y[7715]), .Z(n6057) );
  XOR U8525 ( .A(n6056), .B(n6057), .Z(n6049) );
  AND U8526 ( .A(y[7719]), .B(x[493]), .Z(n5975) );
  NAND U8527 ( .A(y[7729]), .B(x[483]), .Z(n5974) );
  XNOR U8528 ( .A(n5975), .B(n5974), .Z(n6089) );
  XNOR U8529 ( .A(n6089), .B(n6090), .Z(n6073) );
  AND U8530 ( .A(y[7727]), .B(x[485]), .Z(n5977) );
  NAND U8531 ( .A(y[7728]), .B(x[484]), .Z(n5976) );
  XNOR U8532 ( .A(n5977), .B(n5976), .Z(n6104) );
  AND U8533 ( .A(x[487]), .B(y[7725]), .Z(n6105) );
  XOR U8534 ( .A(n6104), .B(n6105), .Z(n6072) );
  XOR U8535 ( .A(n6073), .B(n6074), .Z(n6116) );
  AND U8536 ( .A(x[488]), .B(y[7730]), .Z(n7220) );
  AND U8537 ( .A(x[481]), .B(y[7723]), .Z(n5978) );
  NAND U8538 ( .A(n7220), .B(n5978), .Z(n5982) );
  NANDN U8539 ( .A(n5980), .B(n5979), .Z(n5981) );
  AND U8540 ( .A(n5982), .B(n5981), .Z(n6115) );
  NAND U8541 ( .A(x[497]), .B(y[7721]), .Z(n6941) );
  NANDN U8542 ( .A(n6941), .B(n5983), .Z(n5987) );
  NAND U8543 ( .A(n5985), .B(n5984), .Z(n5986) );
  NAND U8544 ( .A(n5987), .B(n5986), .Z(n6114) );
  XNOR U8545 ( .A(n6116), .B(n6117), .Z(n6043) );
  XOR U8546 ( .A(n6044), .B(n6043), .Z(n6045) );
  NANDN U8547 ( .A(n5989), .B(n5988), .Z(n5993) );
  NANDN U8548 ( .A(n5991), .B(n5990), .Z(n5992) );
  NAND U8549 ( .A(n5993), .B(n5992), .Z(n6046) );
  NAND U8550 ( .A(n5995), .B(n5994), .Z(n5999) );
  NANDN U8551 ( .A(n5997), .B(n5996), .Z(n5998) );
  NAND U8552 ( .A(n5999), .B(n5998), .Z(n6133) );
  NANDN U8553 ( .A(n6001), .B(n6000), .Z(n6005) );
  NAND U8554 ( .A(n6003), .B(n6002), .Z(n6004) );
  AND U8555 ( .A(n6005), .B(n6004), .Z(n6147) );
  NAND U8556 ( .A(n6007), .B(n6006), .Z(n6011) );
  NAND U8557 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U8558 ( .A(n6011), .B(n6010), .Z(n6145) );
  NANDN U8559 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U8560 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U8561 ( .A(n6017), .B(n6016), .Z(n6144) );
  XNOR U8562 ( .A(n6147), .B(n6146), .Z(n6138) );
  XOR U8563 ( .A(n6139), .B(n6138), .Z(n6140) );
  NAND U8564 ( .A(n6019), .B(n6018), .Z(n6023) );
  NANDN U8565 ( .A(n6021), .B(n6020), .Z(n6022) );
  NAND U8566 ( .A(n6023), .B(n6022), .Z(n6141) );
  NAND U8567 ( .A(n6025), .B(n6024), .Z(n6029) );
  NANDN U8568 ( .A(n6027), .B(n6026), .Z(n6028) );
  AND U8569 ( .A(n6029), .B(n6028), .Z(n6158) );
  NANDN U8570 ( .A(n6031), .B(n6030), .Z(n6035) );
  NANDN U8571 ( .A(n6033), .B(n6032), .Z(n6034) );
  AND U8572 ( .A(n6035), .B(n6034), .Z(n6157) );
  XOR U8573 ( .A(n6158), .B(n6157), .Z(n6159) );
  XNOR U8574 ( .A(n6152), .B(n6153), .Z(n6036) );
  XOR U8575 ( .A(n6150), .B(n6036), .Z(N117) );
  NANDN U8576 ( .A(n6038), .B(n6037), .Z(n6042) );
  NAND U8577 ( .A(n6040), .B(n6039), .Z(n6041) );
  AND U8578 ( .A(n6042), .B(n6041), .Z(n6173) );
  NAND U8579 ( .A(n6044), .B(n6043), .Z(n6048) );
  NANDN U8580 ( .A(n6046), .B(n6045), .Z(n6047) );
  AND U8581 ( .A(n6048), .B(n6047), .Z(n6171) );
  NANDN U8582 ( .A(n6050), .B(n6049), .Z(n6054) );
  NANDN U8583 ( .A(n6052), .B(n6051), .Z(n6053) );
  AND U8584 ( .A(n6054), .B(n6053), .Z(n6258) );
  AND U8585 ( .A(x[498]), .B(y[7720]), .Z(n6940) );
  NAND U8586 ( .A(n6940), .B(n6055), .Z(n6059) );
  NAND U8587 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U8588 ( .A(n6059), .B(n6058), .Z(n6262) );
  AND U8589 ( .A(x[491]), .B(y[7731]), .Z(n7680) );
  AND U8590 ( .A(x[481]), .B(y[7721]), .Z(n6060) );
  NAND U8591 ( .A(n7680), .B(n6060), .Z(n6064) );
  NAND U8592 ( .A(n6062), .B(n6061), .Z(n6063) );
  NAND U8593 ( .A(n6064), .B(n6063), .Z(n6261) );
  XOR U8594 ( .A(n6262), .B(n6261), .Z(n6264) );
  AND U8595 ( .A(x[495]), .B(y[7723]), .Z(n6928) );
  NAND U8596 ( .A(n6928), .B(n6065), .Z(n6069) );
  NAND U8597 ( .A(n6067), .B(n6066), .Z(n6068) );
  NAND U8598 ( .A(n6069), .B(n6068), .Z(n6220) );
  AND U8599 ( .A(o[52]), .B(n6070), .Z(n6242) );
  AND U8600 ( .A(x[480]), .B(y[7733]), .Z(n6239) );
  AND U8601 ( .A(x[501]), .B(y[7712]), .Z(n6240) );
  XOR U8602 ( .A(n6239), .B(n6240), .Z(n6241) );
  XOR U8603 ( .A(n6242), .B(n6241), .Z(n6218) );
  AND U8604 ( .A(x[485]), .B(y[7728]), .Z(n6226) );
  AND U8605 ( .A(x[496]), .B(y[7717]), .Z(n6225) );
  XOR U8606 ( .A(n6226), .B(n6225), .Z(n6224) );
  AND U8607 ( .A(x[495]), .B(y[7718]), .Z(n6223) );
  XOR U8608 ( .A(n6224), .B(n6223), .Z(n6217) );
  XOR U8609 ( .A(n6218), .B(n6217), .Z(n6219) );
  XOR U8610 ( .A(n6220), .B(n6219), .Z(n6263) );
  XOR U8611 ( .A(n6264), .B(n6263), .Z(n6255) );
  NANDN U8612 ( .A(n6072), .B(n6071), .Z(n6076) );
  NANDN U8613 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U8614 ( .A(n6076), .B(n6075), .Z(n6256) );
  XOR U8615 ( .A(n6171), .B(n6170), .Z(n6172) );
  NANDN U8616 ( .A(n6078), .B(n6077), .Z(n6082) );
  NAND U8617 ( .A(n6080), .B(n6079), .Z(n6081) );
  AND U8618 ( .A(n6082), .B(n6081), .Z(n6179) );
  NAND U8619 ( .A(n6933), .B(n6083), .Z(n6087) );
  NAND U8620 ( .A(n6085), .B(n6084), .Z(n6086) );
  NAND U8621 ( .A(n6087), .B(n6086), .Z(n6189) );
  NAND U8622 ( .A(n7507), .B(n6088), .Z(n6092) );
  NAND U8623 ( .A(n6090), .B(n6089), .Z(n6091) );
  NAND U8624 ( .A(n6092), .B(n6091), .Z(n6276) );
  AND U8625 ( .A(y[7714]), .B(x[499]), .Z(n6094) );
  NAND U8626 ( .A(y[7722]), .B(x[491]), .Z(n6093) );
  XNOR U8627 ( .A(n6094), .B(n6093), .Z(n6207) );
  NAND U8628 ( .A(x[500]), .B(y[7713]), .Z(n6238) );
  XNOR U8629 ( .A(o[53]), .B(n6238), .Z(n6208) );
  XOR U8630 ( .A(n6207), .B(n6208), .Z(n6274) );
  AND U8631 ( .A(y[7715]), .B(x[498]), .Z(n6096) );
  NAND U8632 ( .A(y[7723]), .B(x[490]), .Z(n6095) );
  XNOR U8633 ( .A(n6096), .B(n6095), .Z(n6246) );
  AND U8634 ( .A(x[481]), .B(y[7732]), .Z(n6247) );
  XOR U8635 ( .A(n6246), .B(n6247), .Z(n6273) );
  XOR U8636 ( .A(n6274), .B(n6273), .Z(n6275) );
  XOR U8637 ( .A(n6276), .B(n6275), .Z(n6188) );
  XOR U8638 ( .A(n6189), .B(n6188), .Z(n6191) );
  AND U8639 ( .A(x[487]), .B(y[7726]), .Z(n6445) );
  AND U8640 ( .A(y[7727]), .B(x[486]), .Z(n6098) );
  NAND U8641 ( .A(y[7719]), .B(x[494]), .Z(n6097) );
  XNOR U8642 ( .A(n6098), .B(n6097), .Z(n6250) );
  XNOR U8643 ( .A(n6445), .B(n6250), .Z(n6197) );
  NAND U8644 ( .A(x[489]), .B(y[7724]), .Z(n6195) );
  NAND U8645 ( .A(x[488]), .B(y[7725]), .Z(n6194) );
  XOR U8646 ( .A(n6195), .B(n6194), .Z(n6196) );
  XNOR U8647 ( .A(n6197), .B(n6196), .Z(n6213) );
  AND U8648 ( .A(y[7721]), .B(x[492]), .Z(n6100) );
  NAND U8649 ( .A(y[7716]), .B(x[497]), .Z(n6099) );
  XNOR U8650 ( .A(n6100), .B(n6099), .Z(n6200) );
  AND U8651 ( .A(x[482]), .B(y[7731]), .Z(n6201) );
  XOR U8652 ( .A(n6200), .B(n6201), .Z(n6212) );
  AND U8653 ( .A(y[7720]), .B(x[493]), .Z(n6102) );
  NAND U8654 ( .A(y[7730]), .B(x[483]), .Z(n6101) );
  XNOR U8655 ( .A(n6102), .B(n6101), .Z(n6234) );
  AND U8656 ( .A(x[484]), .B(y[7729]), .Z(n6235) );
  XOR U8657 ( .A(n6234), .B(n6235), .Z(n6211) );
  XOR U8658 ( .A(n6212), .B(n6211), .Z(n6214) );
  XOR U8659 ( .A(n6213), .B(n6214), .Z(n6270) );
  NAND U8660 ( .A(n6226), .B(n6103), .Z(n6107) );
  NAND U8661 ( .A(n6105), .B(n6104), .Z(n6106) );
  NAND U8662 ( .A(n6107), .B(n6106), .Z(n6268) );
  NAND U8663 ( .A(n6109), .B(n6108), .Z(n6113) );
  NAND U8664 ( .A(n6111), .B(n6110), .Z(n6112) );
  NAND U8665 ( .A(n6113), .B(n6112), .Z(n6267) );
  XOR U8666 ( .A(n6268), .B(n6267), .Z(n6269) );
  XOR U8667 ( .A(n6270), .B(n6269), .Z(n6190) );
  XOR U8668 ( .A(n6191), .B(n6190), .Z(n6177) );
  NANDN U8669 ( .A(n6115), .B(n6114), .Z(n6119) );
  NAND U8670 ( .A(n6117), .B(n6116), .Z(n6118) );
  NAND U8671 ( .A(n6119), .B(n6118), .Z(n6184) );
  NAND U8672 ( .A(n6121), .B(n6120), .Z(n6125) );
  NANDN U8673 ( .A(n6123), .B(n6122), .Z(n6124) );
  NAND U8674 ( .A(n6125), .B(n6124), .Z(n6183) );
  NAND U8675 ( .A(n6127), .B(n6126), .Z(n6131) );
  NANDN U8676 ( .A(n6129), .B(n6128), .Z(n6130) );
  NAND U8677 ( .A(n6131), .B(n6130), .Z(n6182) );
  XOR U8678 ( .A(n6183), .B(n6182), .Z(n6185) );
  XOR U8679 ( .A(n6184), .B(n6185), .Z(n6176) );
  XOR U8680 ( .A(n6177), .B(n6176), .Z(n6178) );
  NANDN U8681 ( .A(n6133), .B(n6132), .Z(n6137) );
  NANDN U8682 ( .A(n6135), .B(n6134), .Z(n6136) );
  NAND U8683 ( .A(n6137), .B(n6136), .Z(n6164) );
  XOR U8684 ( .A(n6165), .B(n6164), .Z(n6167) );
  XNOR U8685 ( .A(n6166), .B(n6167), .Z(n6288) );
  NAND U8686 ( .A(n6139), .B(n6138), .Z(n6143) );
  NANDN U8687 ( .A(n6141), .B(n6140), .Z(n6142) );
  AND U8688 ( .A(n6143), .B(n6142), .Z(n6287) );
  NANDN U8689 ( .A(n6145), .B(n6144), .Z(n6149) );
  NAND U8690 ( .A(n6147), .B(n6146), .Z(n6148) );
  AND U8691 ( .A(n6149), .B(n6148), .Z(n6286) );
  XNOR U8692 ( .A(n6288), .B(n6289), .Z(n6282) );
  OR U8693 ( .A(n6152), .B(n6150), .Z(n6156) );
  ANDN U8694 ( .B(n6152), .A(n6151), .Z(n6154) );
  OR U8695 ( .A(n6154), .B(n6153), .Z(n6155) );
  AND U8696 ( .A(n6156), .B(n6155), .Z(n6281) );
  NAND U8697 ( .A(n6158), .B(n6157), .Z(n6162) );
  NANDN U8698 ( .A(n6160), .B(n6159), .Z(n6161) );
  AND U8699 ( .A(n6162), .B(n6161), .Z(n6280) );
  IV U8700 ( .A(n6280), .Z(n6279) );
  XOR U8701 ( .A(n6281), .B(n6279), .Z(n6163) );
  XNOR U8702 ( .A(n6282), .B(n6163), .Z(N118) );
  NAND U8703 ( .A(n6165), .B(n6164), .Z(n6169) );
  NAND U8704 ( .A(n6167), .B(n6166), .Z(n6168) );
  AND U8705 ( .A(n6169), .B(n6168), .Z(n6296) );
  NAND U8706 ( .A(n6171), .B(n6170), .Z(n6175) );
  NANDN U8707 ( .A(n6173), .B(n6172), .Z(n6174) );
  AND U8708 ( .A(n6175), .B(n6174), .Z(n6294) );
  NAND U8709 ( .A(n6177), .B(n6176), .Z(n6181) );
  NANDN U8710 ( .A(n6179), .B(n6178), .Z(n6180) );
  NAND U8711 ( .A(n6181), .B(n6180), .Z(n6307) );
  NAND U8712 ( .A(n6183), .B(n6182), .Z(n6187) );
  NAND U8713 ( .A(n6185), .B(n6184), .Z(n6186) );
  NAND U8714 ( .A(n6187), .B(n6186), .Z(n6306) );
  XOR U8715 ( .A(n6307), .B(n6306), .Z(n6309) );
  NAND U8716 ( .A(n6189), .B(n6188), .Z(n6193) );
  NAND U8717 ( .A(n6191), .B(n6190), .Z(n6192) );
  NAND U8718 ( .A(n6193), .B(n6192), .Z(n6421) );
  NAND U8719 ( .A(n6195), .B(n6194), .Z(n6199) );
  NAND U8720 ( .A(n6197), .B(n6196), .Z(n6198) );
  NAND U8721 ( .A(n6199), .B(n6198), .Z(n6415) );
  NANDN U8722 ( .A(n6941), .B(n6366), .Z(n6203) );
  NAND U8723 ( .A(n6201), .B(n6200), .Z(n6202) );
  NAND U8724 ( .A(n6203), .B(n6202), .Z(n6344) );
  AND U8725 ( .A(x[485]), .B(y[7729]), .Z(n6388) );
  AND U8726 ( .A(x[497]), .B(y[7717]), .Z(n6389) );
  XOR U8727 ( .A(n6388), .B(n6389), .Z(n6390) );
  AND U8728 ( .A(x[496]), .B(y[7718]), .Z(n6391) );
  XOR U8729 ( .A(n6390), .B(n6391), .Z(n6343) );
  AND U8730 ( .A(y[7716]), .B(x[498]), .Z(n6205) );
  NAND U8731 ( .A(y[7722]), .B(x[492]), .Z(n6204) );
  XNOR U8732 ( .A(n6205), .B(n6204), .Z(n6367) );
  AND U8733 ( .A(x[484]), .B(y[7730]), .Z(n6368) );
  XOR U8734 ( .A(n6367), .B(n6368), .Z(n6342) );
  XOR U8735 ( .A(n6343), .B(n6342), .Z(n6345) );
  XNOR U8736 ( .A(n6344), .B(n6345), .Z(n6412) );
  AND U8737 ( .A(x[499]), .B(y[7722]), .Z(n7398) );
  NAND U8738 ( .A(n7398), .B(n6206), .Z(n6210) );
  NAND U8739 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U8740 ( .A(n6210), .B(n6209), .Z(n6413) );
  XOR U8741 ( .A(n6412), .B(n6413), .Z(n6414) );
  XNOR U8742 ( .A(n6415), .B(n6414), .Z(n6418) );
  NAND U8743 ( .A(n6212), .B(n6211), .Z(n6216) );
  NAND U8744 ( .A(n6214), .B(n6213), .Z(n6215) );
  NAND U8745 ( .A(n6216), .B(n6215), .Z(n6401) );
  NAND U8746 ( .A(n6218), .B(n6217), .Z(n6222) );
  NAND U8747 ( .A(n6220), .B(n6219), .Z(n6221) );
  NAND U8748 ( .A(n6222), .B(n6221), .Z(n6400) );
  XOR U8749 ( .A(n6401), .B(n6400), .Z(n6403) );
  AND U8750 ( .A(n6224), .B(n6223), .Z(n6228) );
  NAND U8751 ( .A(n6226), .B(n6225), .Z(n6227) );
  NANDN U8752 ( .A(n6228), .B(n6227), .Z(n6363) );
  AND U8753 ( .A(y[7721]), .B(x[493]), .Z(n6230) );
  NAND U8754 ( .A(y[7714]), .B(x[500]), .Z(n6229) );
  XNOR U8755 ( .A(n6230), .B(n6229), .Z(n6384) );
  AND U8756 ( .A(x[482]), .B(y[7732]), .Z(n6385) );
  XOR U8757 ( .A(n6384), .B(n6385), .Z(n6361) );
  AND U8758 ( .A(y[7728]), .B(x[486]), .Z(n6232) );
  NAND U8759 ( .A(y[7719]), .B(x[495]), .Z(n6231) );
  XNOR U8760 ( .A(n6232), .B(n6231), .Z(n6396) );
  XOR U8761 ( .A(n6361), .B(n6360), .Z(n6362) );
  XOR U8762 ( .A(n6363), .B(n6362), .Z(n6407) );
  AND U8763 ( .A(x[493]), .B(y[7730]), .Z(n7682) );
  NAND U8764 ( .A(n6233), .B(n7682), .Z(n6237) );
  NAND U8765 ( .A(n6235), .B(n6234), .Z(n6236) );
  NAND U8766 ( .A(n6237), .B(n6236), .Z(n6333) );
  AND U8767 ( .A(x[481]), .B(y[7733]), .Z(n6356) );
  XOR U8768 ( .A(n6357), .B(n6356), .Z(n6355) );
  ANDN U8769 ( .B(o[53]), .A(n6238), .Z(n6354) );
  XOR U8770 ( .A(n6355), .B(n6354), .Z(n6330) );
  AND U8771 ( .A(x[494]), .B(y[7720]), .Z(n6348) );
  NAND U8772 ( .A(x[483]), .B(y[7731]), .Z(n6349) );
  XNOR U8773 ( .A(n6348), .B(n6349), .Z(n6350) );
  NAND U8774 ( .A(x[499]), .B(y[7715]), .Z(n6351) );
  XNOR U8775 ( .A(n6350), .B(n6351), .Z(n6331) );
  XOR U8776 ( .A(n6330), .B(n6331), .Z(n6332) );
  XOR U8777 ( .A(n6333), .B(n6332), .Z(n6406) );
  XOR U8778 ( .A(n6407), .B(n6406), .Z(n6409) );
  NAND U8779 ( .A(n6240), .B(n6239), .Z(n6244) );
  NAND U8780 ( .A(n6242), .B(n6241), .Z(n6243) );
  NAND U8781 ( .A(n6244), .B(n6243), .Z(n6325) );
  AND U8782 ( .A(x[498]), .B(y[7723]), .Z(n7401) );
  NAND U8783 ( .A(n7401), .B(n6245), .Z(n6249) );
  NAND U8784 ( .A(n6247), .B(n6246), .Z(n6248) );
  NAND U8785 ( .A(n6249), .B(n6248), .Z(n6324) );
  XOR U8786 ( .A(n6325), .B(n6324), .Z(n6327) );
  AND U8787 ( .A(x[494]), .B(y[7727]), .Z(n7441) );
  NAND U8788 ( .A(n7441), .B(n6395), .Z(n6252) );
  NAND U8789 ( .A(n6445), .B(n6250), .Z(n6251) );
  NAND U8790 ( .A(n6252), .B(n6251), .Z(n6339) );
  AND U8791 ( .A(x[480]), .B(y[7734]), .Z(n6371) );
  AND U8792 ( .A(x[502]), .B(y[7712]), .Z(n6372) );
  XOR U8793 ( .A(n6371), .B(n6372), .Z(n6373) );
  NAND U8794 ( .A(x[501]), .B(y[7713]), .Z(n6394) );
  XNOR U8795 ( .A(o[54]), .B(n6394), .Z(n6374) );
  XOR U8796 ( .A(n6373), .B(n6374), .Z(n6337) );
  AND U8797 ( .A(y[7727]), .B(x[487]), .Z(n6254) );
  NAND U8798 ( .A(y[7726]), .B(x[488]), .Z(n6253) );
  XNOR U8799 ( .A(n6254), .B(n6253), .Z(n6377) );
  XOR U8800 ( .A(n6337), .B(n6336), .Z(n6338) );
  XOR U8801 ( .A(n6339), .B(n6338), .Z(n6326) );
  XOR U8802 ( .A(n6327), .B(n6326), .Z(n6408) );
  XOR U8803 ( .A(n6409), .B(n6408), .Z(n6402) );
  XOR U8804 ( .A(n6403), .B(n6402), .Z(n6419) );
  XOR U8805 ( .A(n6418), .B(n6419), .Z(n6420) );
  XOR U8806 ( .A(n6421), .B(n6420), .Z(n6315) );
  NANDN U8807 ( .A(n6256), .B(n6255), .Z(n6260) );
  NANDN U8808 ( .A(n6258), .B(n6257), .Z(n6259) );
  NAND U8809 ( .A(n6260), .B(n6259), .Z(n6312) );
  NAND U8810 ( .A(n6262), .B(n6261), .Z(n6266) );
  NAND U8811 ( .A(n6264), .B(n6263), .Z(n6265) );
  NAND U8812 ( .A(n6266), .B(n6265), .Z(n6321) );
  NAND U8813 ( .A(n6268), .B(n6267), .Z(n6272) );
  NAND U8814 ( .A(n6270), .B(n6269), .Z(n6271) );
  NAND U8815 ( .A(n6272), .B(n6271), .Z(n6319) );
  NAND U8816 ( .A(n6274), .B(n6273), .Z(n6278) );
  NAND U8817 ( .A(n6276), .B(n6275), .Z(n6277) );
  NAND U8818 ( .A(n6278), .B(n6277), .Z(n6318) );
  XOR U8819 ( .A(n6319), .B(n6318), .Z(n6320) );
  XOR U8820 ( .A(n6321), .B(n6320), .Z(n6313) );
  XOR U8821 ( .A(n6312), .B(n6313), .Z(n6314) );
  XOR U8822 ( .A(n6315), .B(n6314), .Z(n6308) );
  XOR U8823 ( .A(n6309), .B(n6308), .Z(n6293) );
  XNOR U8824 ( .A(n6296), .B(n6295), .Z(n6302) );
  OR U8825 ( .A(n6281), .B(n6279), .Z(n6285) );
  ANDN U8826 ( .B(n6281), .A(n6280), .Z(n6283) );
  OR U8827 ( .A(n6283), .B(n6282), .Z(n6284) );
  AND U8828 ( .A(n6285), .B(n6284), .Z(n6301) );
  NANDN U8829 ( .A(n6287), .B(n6286), .Z(n6291) );
  NAND U8830 ( .A(n6289), .B(n6288), .Z(n6290) );
  NAND U8831 ( .A(n6291), .B(n6290), .Z(n6300) );
  IV U8832 ( .A(n6300), .Z(n6299) );
  XOR U8833 ( .A(n6301), .B(n6299), .Z(n6292) );
  XNOR U8834 ( .A(n6302), .B(n6292), .Z(N119) );
  NANDN U8835 ( .A(n6294), .B(n6293), .Z(n6298) );
  NAND U8836 ( .A(n6296), .B(n6295), .Z(n6297) );
  NAND U8837 ( .A(n6298), .B(n6297), .Z(n6555) );
  IV U8838 ( .A(n6555), .Z(n6554) );
  OR U8839 ( .A(n6301), .B(n6299), .Z(n6305) );
  ANDN U8840 ( .B(n6301), .A(n6300), .Z(n6303) );
  OR U8841 ( .A(n6303), .B(n6302), .Z(n6304) );
  AND U8842 ( .A(n6305), .B(n6304), .Z(n6556) );
  NAND U8843 ( .A(n6307), .B(n6306), .Z(n6311) );
  NAND U8844 ( .A(n6309), .B(n6308), .Z(n6310) );
  AND U8845 ( .A(n6311), .B(n6310), .Z(n6564) );
  NAND U8846 ( .A(n6313), .B(n6312), .Z(n6317) );
  NAND U8847 ( .A(n6315), .B(n6314), .Z(n6316) );
  AND U8848 ( .A(n6317), .B(n6316), .Z(n6562) );
  NAND U8849 ( .A(n6319), .B(n6318), .Z(n6323) );
  NAND U8850 ( .A(n6321), .B(n6320), .Z(n6322) );
  NAND U8851 ( .A(n6323), .B(n6322), .Z(n6539) );
  NAND U8852 ( .A(n6325), .B(n6324), .Z(n6329) );
  NAND U8853 ( .A(n6327), .B(n6326), .Z(n6328) );
  NAND U8854 ( .A(n6329), .B(n6328), .Z(n6533) );
  NAND U8855 ( .A(n6331), .B(n6330), .Z(n6335) );
  NAND U8856 ( .A(n6333), .B(n6332), .Z(n6334) );
  NAND U8857 ( .A(n6335), .B(n6334), .Z(n6531) );
  NAND U8858 ( .A(n6337), .B(n6336), .Z(n6341) );
  NAND U8859 ( .A(n6339), .B(n6338), .Z(n6340) );
  NAND U8860 ( .A(n6341), .B(n6340), .Z(n6530) );
  XOR U8861 ( .A(n6531), .B(n6530), .Z(n6532) );
  XOR U8862 ( .A(n6533), .B(n6532), .Z(n6551) );
  NAND U8863 ( .A(n6343), .B(n6342), .Z(n6347) );
  NAND U8864 ( .A(n6345), .B(n6344), .Z(n6346) );
  NAND U8865 ( .A(n6347), .B(n6346), .Z(n6549) );
  NANDN U8866 ( .A(n6349), .B(n6348), .Z(n6353) );
  NANDN U8867 ( .A(n6351), .B(n6350), .Z(n6352) );
  AND U8868 ( .A(n6353), .B(n6352), .Z(n6477) );
  XNOR U8869 ( .A(n6477), .B(n6476), .Z(n6478) );
  AND U8870 ( .A(y[7728]), .B(x[487]), .Z(n6359) );
  NAND U8871 ( .A(y[7726]), .B(x[489]), .Z(n6358) );
  XNOR U8872 ( .A(n6359), .B(n6358), .Z(n6446) );
  NAND U8873 ( .A(x[490]), .B(y[7725]), .Z(n6483) );
  XNOR U8874 ( .A(n6482), .B(n6483), .Z(n6484) );
  AND U8875 ( .A(x[486]), .B(y[7729]), .Z(n6437) );
  NAND U8876 ( .A(x[495]), .B(y[7720]), .Z(n6438) );
  XNOR U8877 ( .A(n6437), .B(n6438), .Z(n6439) );
  NAND U8878 ( .A(x[491]), .B(y[7724]), .Z(n6440) );
  XOR U8879 ( .A(n6439), .B(n6440), .Z(n6485) );
  XOR U8880 ( .A(n6484), .B(n6485), .Z(n6479) );
  XNOR U8881 ( .A(n6478), .B(n6479), .Z(n6548) );
  XOR U8882 ( .A(n6549), .B(n6548), .Z(n6550) );
  XOR U8883 ( .A(n6551), .B(n6550), .Z(n6537) );
  NAND U8884 ( .A(n6361), .B(n6360), .Z(n6365) );
  NAND U8885 ( .A(n6363), .B(n6362), .Z(n6364) );
  NAND U8886 ( .A(n6365), .B(n6364), .Z(n6471) );
  NAND U8887 ( .A(x[498]), .B(y[7722]), .Z(n7251) );
  NANDN U8888 ( .A(n7251), .B(n6366), .Z(n6370) );
  NAND U8889 ( .A(n6368), .B(n6367), .Z(n6369) );
  NAND U8890 ( .A(n6370), .B(n6369), .Z(n6507) );
  NAND U8891 ( .A(n6372), .B(n6371), .Z(n6376) );
  NAND U8892 ( .A(n6374), .B(n6373), .Z(n6375) );
  NAND U8893 ( .A(n6376), .B(n6375), .Z(n6506) );
  XOR U8894 ( .A(n6507), .B(n6506), .Z(n6509) );
  NANDN U8895 ( .A(n6447), .B(n6445), .Z(n6380) );
  NANDN U8896 ( .A(n6378), .B(n6377), .Z(n6379) );
  NAND U8897 ( .A(n6380), .B(n6379), .Z(n6520) );
  AND U8898 ( .A(x[480]), .B(y[7735]), .Z(n6454) );
  NAND U8899 ( .A(x[503]), .B(y[7712]), .Z(n6455) );
  XNOR U8900 ( .A(n6454), .B(n6455), .Z(n6456) );
  NAND U8901 ( .A(x[502]), .B(y[7713]), .Z(n6436) );
  XOR U8902 ( .A(o[55]), .B(n6436), .Z(n6457) );
  XNOR U8903 ( .A(n6456), .B(n6457), .Z(n6519) );
  NAND U8904 ( .A(y[7715]), .B(x[500]), .Z(n6381) );
  XNOR U8905 ( .A(n6382), .B(n6381), .Z(n6433) );
  AND U8906 ( .A(x[499]), .B(y[7716]), .Z(n6432) );
  XOR U8907 ( .A(n6433), .B(n6432), .Z(n6518) );
  XOR U8908 ( .A(n6519), .B(n6518), .Z(n6521) );
  XOR U8909 ( .A(n6520), .B(n6521), .Z(n6508) );
  XOR U8910 ( .A(n6509), .B(n6508), .Z(n6470) );
  XOR U8911 ( .A(n6471), .B(n6470), .Z(n6473) );
  NAND U8912 ( .A(x[500]), .B(y[7721]), .Z(n7453) );
  AND U8913 ( .A(x[493]), .B(y[7714]), .Z(n6383) );
  NANDN U8914 ( .A(n7453), .B(n6383), .Z(n6387) );
  NAND U8915 ( .A(n6385), .B(n6384), .Z(n6386) );
  NAND U8916 ( .A(n6387), .B(n6386), .Z(n6465) );
  NAND U8917 ( .A(n6389), .B(n6388), .Z(n6393) );
  NAND U8918 ( .A(n6391), .B(n6390), .Z(n6392) );
  NAND U8919 ( .A(n6393), .B(n6392), .Z(n6527) );
  AND U8920 ( .A(x[493]), .B(y[7722]), .Z(n6500) );
  NAND U8921 ( .A(x[482]), .B(y[7733]), .Z(n6501) );
  XNOR U8922 ( .A(n6500), .B(n6501), .Z(n6502) );
  NAND U8923 ( .A(x[501]), .B(y[7714]), .Z(n6503) );
  XNOR U8924 ( .A(n6502), .B(n6503), .Z(n6525) );
  AND U8925 ( .A(x[492]), .B(y[7723]), .Z(n6450) );
  NAND U8926 ( .A(x[481]), .B(y[7734]), .Z(n6451) );
  XNOR U8927 ( .A(n6450), .B(n6451), .Z(n6453) );
  ANDN U8928 ( .B(o[54]), .A(n6394), .Z(n6452) );
  XOR U8929 ( .A(n6453), .B(n6452), .Z(n6524) );
  XOR U8930 ( .A(n6525), .B(n6524), .Z(n6526) );
  XOR U8931 ( .A(n6527), .B(n6526), .Z(n6464) );
  XOR U8932 ( .A(n6465), .B(n6464), .Z(n6467) );
  AND U8933 ( .A(x[495]), .B(y[7728]), .Z(n7675) );
  NAND U8934 ( .A(n7675), .B(n6395), .Z(n6399) );
  NANDN U8935 ( .A(n6397), .B(n6396), .Z(n6398) );
  NAND U8936 ( .A(n6399), .B(n6398), .Z(n6515) );
  AND U8937 ( .A(x[494]), .B(y[7721]), .Z(n6494) );
  NAND U8938 ( .A(x[483]), .B(y[7732]), .Z(n6495) );
  XNOR U8939 ( .A(n6494), .B(n6495), .Z(n6496) );
  NAND U8940 ( .A(x[484]), .B(y[7731]), .Z(n6497) );
  XNOR U8941 ( .A(n6496), .B(n6497), .Z(n6512) );
  AND U8942 ( .A(x[485]), .B(y[7730]), .Z(n6488) );
  NAND U8943 ( .A(x[498]), .B(y[7717]), .Z(n6489) );
  XNOR U8944 ( .A(n6488), .B(n6489), .Z(n6490) );
  NAND U8945 ( .A(x[497]), .B(y[7718]), .Z(n6491) );
  XNOR U8946 ( .A(n6490), .B(n6491), .Z(n6513) );
  XOR U8947 ( .A(n6512), .B(n6513), .Z(n6514) );
  XOR U8948 ( .A(n6515), .B(n6514), .Z(n6466) );
  XOR U8949 ( .A(n6467), .B(n6466), .Z(n6472) );
  XOR U8950 ( .A(n6473), .B(n6472), .Z(n6536) );
  XOR U8951 ( .A(n6537), .B(n6536), .Z(n6538) );
  XNOR U8952 ( .A(n6539), .B(n6538), .Z(n6427) );
  NAND U8953 ( .A(n6401), .B(n6400), .Z(n6405) );
  NAND U8954 ( .A(n6403), .B(n6402), .Z(n6404) );
  NAND U8955 ( .A(n6405), .B(n6404), .Z(n6545) );
  NAND U8956 ( .A(n6407), .B(n6406), .Z(n6411) );
  NAND U8957 ( .A(n6409), .B(n6408), .Z(n6410) );
  NAND U8958 ( .A(n6411), .B(n6410), .Z(n6543) );
  NAND U8959 ( .A(n6413), .B(n6412), .Z(n6417) );
  NAND U8960 ( .A(n6415), .B(n6414), .Z(n6416) );
  AND U8961 ( .A(n6417), .B(n6416), .Z(n6542) );
  XOR U8962 ( .A(n6543), .B(n6542), .Z(n6544) );
  XNOR U8963 ( .A(n6545), .B(n6544), .Z(n6425) );
  NAND U8964 ( .A(n6419), .B(n6418), .Z(n6423) );
  NAND U8965 ( .A(n6421), .B(n6420), .Z(n6422) );
  AND U8966 ( .A(n6423), .B(n6422), .Z(n6426) );
  XOR U8967 ( .A(n6425), .B(n6426), .Z(n6428) );
  XOR U8968 ( .A(n6427), .B(n6428), .Z(n6561) );
  XOR U8969 ( .A(n6562), .B(n6561), .Z(n6563) );
  XOR U8970 ( .A(n6564), .B(n6563), .Z(n6557) );
  XNOR U8971 ( .A(n6556), .B(n6557), .Z(n6424) );
  XOR U8972 ( .A(n6554), .B(n6424), .Z(N120) );
  NAND U8973 ( .A(n6426), .B(n6425), .Z(n6430) );
  NAND U8974 ( .A(n6428), .B(n6427), .Z(n6429) );
  AND U8975 ( .A(n6430), .B(n6429), .Z(n6705) );
  AND U8976 ( .A(x[500]), .B(y[7719]), .Z(n6431) );
  NAND U8977 ( .A(n6431), .B(n6592), .Z(n6435) );
  NAND U8978 ( .A(n6433), .B(n6432), .Z(n6434) );
  AND U8979 ( .A(n6435), .B(n6434), .Z(n6616) );
  AND U8980 ( .A(x[502]), .B(y[7714]), .Z(n6633) );
  XOR U8981 ( .A(n6634), .B(n6633), .Z(n6636) );
  AND U8982 ( .A(x[482]), .B(y[7734]), .Z(n6635) );
  XOR U8983 ( .A(n6636), .B(n6635), .Z(n6614) );
  AND U8984 ( .A(x[481]), .B(y[7735]), .Z(n6641) );
  XOR U8985 ( .A(n6642), .B(n6641), .Z(n6640) );
  ANDN U8986 ( .B(o[55]), .A(n6436), .Z(n6639) );
  XOR U8987 ( .A(n6640), .B(n6639), .Z(n6613) );
  XOR U8988 ( .A(n6614), .B(n6613), .Z(n6615) );
  XNOR U8989 ( .A(n6616), .B(n6615), .Z(n6671) );
  NANDN U8990 ( .A(n6438), .B(n6437), .Z(n6442) );
  NANDN U8991 ( .A(n6440), .B(n6439), .Z(n6441) );
  AND U8992 ( .A(n6442), .B(n6441), .Z(n6610) );
  AND U8993 ( .A(y[7720]), .B(x[496]), .Z(n6444) );
  NAND U8994 ( .A(y[7715]), .B(x[501]), .Z(n6443) );
  XNOR U8995 ( .A(n6444), .B(n6443), .Z(n6593) );
  NAND U8996 ( .A(x[485]), .B(y[7731]), .Z(n6594) );
  XNOR U8997 ( .A(n6593), .B(n6594), .Z(n6607) );
  AND U8998 ( .A(x[486]), .B(y[7730]), .Z(n6987) );
  NAND U8999 ( .A(x[500]), .B(y[7716]), .Z(n6804) );
  NAND U9000 ( .A(x[499]), .B(y[7717]), .Z(n6600) );
  XOR U9001 ( .A(n6599), .B(n6600), .Z(n6608) );
  XNOR U9002 ( .A(n6607), .B(n6608), .Z(n6609) );
  XNOR U9003 ( .A(n6610), .B(n6609), .Z(n6588) );
  NAND U9004 ( .A(n6734), .B(n6445), .Z(n6449) );
  NANDN U9005 ( .A(n6447), .B(n6446), .Z(n6448) );
  AND U9006 ( .A(n6449), .B(n6448), .Z(n6587) );
  XOR U9007 ( .A(n6587), .B(n6586), .Z(n6589) );
  XOR U9008 ( .A(n6588), .B(n6589), .Z(n6672) );
  XNOR U9009 ( .A(n6671), .B(n6672), .Z(n6674) );
  NANDN U9010 ( .A(n6455), .B(n6454), .Z(n6459) );
  NANDN U9011 ( .A(n6457), .B(n6456), .Z(n6458) );
  AND U9012 ( .A(n6459), .B(n6458), .Z(n6666) );
  AND U9013 ( .A(x[483]), .B(y[7733]), .Z(n6653) );
  XOR U9014 ( .A(n6654), .B(n6653), .Z(n6656) );
  NAND U9015 ( .A(x[484]), .B(y[7732]), .Z(n6655) );
  XNOR U9016 ( .A(n6656), .B(n6655), .Z(n6665) );
  XNOR U9017 ( .A(n6666), .B(n6665), .Z(n6667) );
  AND U9018 ( .A(y[7727]), .B(x[489]), .Z(n6461) );
  NAND U9019 ( .A(y[7726]), .B(x[490]), .Z(n6460) );
  XNOR U9020 ( .A(n6461), .B(n6460), .Z(n6624) );
  AND U9021 ( .A(y[7722]), .B(x[494]), .Z(n6463) );
  NAND U9022 ( .A(y[7728]), .B(x[488]), .Z(n6462) );
  XNOR U9023 ( .A(n6463), .B(n6462), .Z(n6629) );
  NAND U9024 ( .A(x[491]), .B(y[7725]), .Z(n6630) );
  XOR U9025 ( .A(n6629), .B(n6630), .Z(n6625) );
  XOR U9026 ( .A(n6624), .B(n6625), .Z(n6668) );
  XNOR U9027 ( .A(n6667), .B(n6668), .Z(n6673) );
  XNOR U9028 ( .A(n6674), .B(n6673), .Z(n6684) );
  NAND U9029 ( .A(n6465), .B(n6464), .Z(n6469) );
  NAND U9030 ( .A(n6467), .B(n6466), .Z(n6468) );
  AND U9031 ( .A(n6469), .B(n6468), .Z(n6683) );
  XOR U9032 ( .A(n6684), .B(n6683), .Z(n6685) );
  NAND U9033 ( .A(n6471), .B(n6470), .Z(n6475) );
  NAND U9034 ( .A(n6473), .B(n6472), .Z(n6474) );
  AND U9035 ( .A(n6475), .B(n6474), .Z(n6686) );
  XOR U9036 ( .A(n6685), .B(n6686), .Z(n6692) );
  NANDN U9037 ( .A(n6477), .B(n6476), .Z(n6481) );
  NANDN U9038 ( .A(n6479), .B(n6478), .Z(n6480) );
  AND U9039 ( .A(n6481), .B(n6480), .Z(n6679) );
  NANDN U9040 ( .A(n6483), .B(n6482), .Z(n6487) );
  NANDN U9041 ( .A(n6485), .B(n6484), .Z(n6486) );
  AND U9042 ( .A(n6487), .B(n6486), .Z(n6678) );
  NANDN U9043 ( .A(n6489), .B(n6488), .Z(n6493) );
  NANDN U9044 ( .A(n6491), .B(n6490), .Z(n6492) );
  AND U9045 ( .A(n6493), .B(n6492), .Z(n6606) );
  AND U9046 ( .A(x[480]), .B(y[7736]), .Z(n6659) );
  NAND U9047 ( .A(x[504]), .B(y[7712]), .Z(n6660) );
  XNOR U9048 ( .A(n6659), .B(n6660), .Z(n6661) );
  NAND U9049 ( .A(x[503]), .B(y[7713]), .Z(n6652) );
  XOR U9050 ( .A(o[56]), .B(n6652), .Z(n6662) );
  XNOR U9051 ( .A(n6661), .B(n6662), .Z(n6604) );
  AND U9052 ( .A(x[487]), .B(y[7729]), .Z(n6646) );
  AND U9053 ( .A(x[498]), .B(y[7718]), .Z(n6645) );
  XOR U9054 ( .A(n6646), .B(n6645), .Z(n6648) );
  AND U9055 ( .A(x[497]), .B(y[7719]), .Z(n6647) );
  XOR U9056 ( .A(n6648), .B(n6647), .Z(n6603) );
  XOR U9057 ( .A(n6604), .B(n6603), .Z(n6605) );
  XNOR U9058 ( .A(n6606), .B(n6605), .Z(n6582) );
  NANDN U9059 ( .A(n6495), .B(n6494), .Z(n6499) );
  NANDN U9060 ( .A(n6497), .B(n6496), .Z(n6498) );
  AND U9061 ( .A(n6499), .B(n6498), .Z(n6581) );
  NANDN U9062 ( .A(n6501), .B(n6500), .Z(n6505) );
  NANDN U9063 ( .A(n6503), .B(n6502), .Z(n6504) );
  NAND U9064 ( .A(n6505), .B(n6504), .Z(n6580) );
  XOR U9065 ( .A(n6581), .B(n6580), .Z(n6583) );
  XNOR U9066 ( .A(n6582), .B(n6583), .Z(n6677) );
  XOR U9067 ( .A(n6678), .B(n6677), .Z(n6680) );
  XNOR U9068 ( .A(n6679), .B(n6680), .Z(n6577) );
  NAND U9069 ( .A(n6507), .B(n6506), .Z(n6511) );
  NAND U9070 ( .A(n6509), .B(n6508), .Z(n6510) );
  AND U9071 ( .A(n6511), .B(n6510), .Z(n6620) );
  NAND U9072 ( .A(n6513), .B(n6512), .Z(n6517) );
  NAND U9073 ( .A(n6515), .B(n6514), .Z(n6516) );
  AND U9074 ( .A(n6517), .B(n6516), .Z(n6618) );
  NAND U9075 ( .A(n6519), .B(n6518), .Z(n6523) );
  NAND U9076 ( .A(n6521), .B(n6520), .Z(n6522) );
  AND U9077 ( .A(n6523), .B(n6522), .Z(n6617) );
  XOR U9078 ( .A(n6618), .B(n6617), .Z(n6619) );
  XOR U9079 ( .A(n6620), .B(n6619), .Z(n6574) );
  NAND U9080 ( .A(n6525), .B(n6524), .Z(n6529) );
  NAND U9081 ( .A(n6527), .B(n6526), .Z(n6528) );
  AND U9082 ( .A(n6529), .B(n6528), .Z(n6575) );
  XOR U9083 ( .A(n6574), .B(n6575), .Z(n6576) );
  XOR U9084 ( .A(n6577), .B(n6576), .Z(n6689) );
  NAND U9085 ( .A(n6531), .B(n6530), .Z(n6535) );
  NAND U9086 ( .A(n6533), .B(n6532), .Z(n6534) );
  AND U9087 ( .A(n6535), .B(n6534), .Z(n6690) );
  XOR U9088 ( .A(n6689), .B(n6690), .Z(n6691) );
  XNOR U9089 ( .A(n6692), .B(n6691), .Z(n6703) );
  NAND U9090 ( .A(n6537), .B(n6536), .Z(n6541) );
  NAND U9091 ( .A(n6539), .B(n6538), .Z(n6540) );
  NAND U9092 ( .A(n6541), .B(n6540), .Z(n6571) );
  NAND U9093 ( .A(n6543), .B(n6542), .Z(n6547) );
  NAND U9094 ( .A(n6545), .B(n6544), .Z(n6546) );
  NAND U9095 ( .A(n6547), .B(n6546), .Z(n6569) );
  NAND U9096 ( .A(n6549), .B(n6548), .Z(n6553) );
  NAND U9097 ( .A(n6551), .B(n6550), .Z(n6552) );
  NAND U9098 ( .A(n6553), .B(n6552), .Z(n6568) );
  XOR U9099 ( .A(n6569), .B(n6568), .Z(n6570) );
  XOR U9100 ( .A(n6571), .B(n6570), .Z(n6702) );
  XOR U9101 ( .A(n6703), .B(n6702), .Z(n6704) );
  XNOR U9102 ( .A(n6705), .B(n6704), .Z(n6698) );
  OR U9103 ( .A(n6556), .B(n6554), .Z(n6560) );
  ANDN U9104 ( .B(n6556), .A(n6555), .Z(n6558) );
  OR U9105 ( .A(n6558), .B(n6557), .Z(n6559) );
  AND U9106 ( .A(n6560), .B(n6559), .Z(n6697) );
  NAND U9107 ( .A(n6562), .B(n6561), .Z(n6566) );
  NAND U9108 ( .A(n6564), .B(n6563), .Z(n6565) );
  AND U9109 ( .A(n6566), .B(n6565), .Z(n6696) );
  IV U9110 ( .A(n6696), .Z(n6695) );
  XOR U9111 ( .A(n6697), .B(n6695), .Z(n6567) );
  XNOR U9112 ( .A(n6698), .B(n6567), .Z(N121) );
  NAND U9113 ( .A(n6569), .B(n6568), .Z(n6573) );
  NAND U9114 ( .A(n6571), .B(n6570), .Z(n6572) );
  AND U9115 ( .A(n6573), .B(n6572), .Z(n6855) );
  NAND U9116 ( .A(n6575), .B(n6574), .Z(n6579) );
  NAND U9117 ( .A(n6577), .B(n6576), .Z(n6578) );
  NAND U9118 ( .A(n6579), .B(n6578), .Z(n6717) );
  NANDN U9119 ( .A(n6581), .B(n6580), .Z(n6585) );
  NANDN U9120 ( .A(n6583), .B(n6582), .Z(n6584) );
  AND U9121 ( .A(n6585), .B(n6584), .Z(n6722) );
  NANDN U9122 ( .A(n6587), .B(n6586), .Z(n6591) );
  NANDN U9123 ( .A(n6589), .B(n6588), .Z(n6590) );
  NAND U9124 ( .A(n6591), .B(n6590), .Z(n6721) );
  XNOR U9125 ( .A(n6722), .B(n6721), .Z(n6723) );
  NAND U9126 ( .A(x[501]), .B(y[7720]), .Z(n7689) );
  NANDN U9127 ( .A(n7689), .B(n6592), .Z(n6596) );
  NANDN U9128 ( .A(n6594), .B(n6593), .Z(n6595) );
  AND U9129 ( .A(n6596), .B(n6595), .Z(n6824) );
  AND U9130 ( .A(x[502]), .B(y[7715]), .Z(n6793) );
  AND U9131 ( .A(x[485]), .B(y[7732]), .Z(n6792) );
  NAND U9132 ( .A(x[497]), .B(y[7720]), .Z(n6791) );
  XOR U9133 ( .A(n6792), .B(n6791), .Z(n6794) );
  XOR U9134 ( .A(n6793), .B(n6794), .Z(n6822) );
  AND U9135 ( .A(y[7717]), .B(x[500]), .Z(n6598) );
  NAND U9136 ( .A(y[7716]), .B(x[501]), .Z(n6597) );
  XNOR U9137 ( .A(n6598), .B(n6597), .Z(n6805) );
  NAND U9138 ( .A(x[499]), .B(y[7718]), .Z(n6806) );
  XNOR U9139 ( .A(n6822), .B(n6821), .Z(n6823) );
  XOR U9140 ( .A(n6824), .B(n6823), .Z(n6748) );
  NANDN U9141 ( .A(n6804), .B(n6987), .Z(n6602) );
  NANDN U9142 ( .A(n6600), .B(n6599), .Z(n6601) );
  AND U9143 ( .A(n6602), .B(n6601), .Z(n6829) );
  AND U9144 ( .A(x[495]), .B(y[7722]), .Z(n6811) );
  AND U9145 ( .A(x[498]), .B(y[7719]), .Z(n6810) );
  NAND U9146 ( .A(x[486]), .B(y[7731]), .Z(n6809) );
  XOR U9147 ( .A(n6810), .B(n6809), .Z(n6812) );
  XOR U9148 ( .A(n6811), .B(n6812), .Z(n6828) );
  AND U9149 ( .A(x[503]), .B(y[7714]), .Z(n6787) );
  AND U9150 ( .A(x[484]), .B(y[7733]), .Z(n6786) );
  NAND U9151 ( .A(x[496]), .B(y[7721]), .Z(n6785) );
  XOR U9152 ( .A(n6786), .B(n6785), .Z(n6788) );
  XNOR U9153 ( .A(n6787), .B(n6788), .Z(n6827) );
  XOR U9154 ( .A(n6828), .B(n6827), .Z(n6830) );
  XNOR U9155 ( .A(n6829), .B(n6830), .Z(n6747) );
  XOR U9156 ( .A(n6748), .B(n6747), .Z(n6750) );
  XOR U9157 ( .A(n6750), .B(n6749), .Z(n6762) );
  NANDN U9158 ( .A(n6608), .B(n6607), .Z(n6612) );
  NANDN U9159 ( .A(n6610), .B(n6609), .Z(n6611) );
  AND U9160 ( .A(n6612), .B(n6611), .Z(n6760) );
  XNOR U9161 ( .A(n6760), .B(n6759), .Z(n6761) );
  XOR U9162 ( .A(n6762), .B(n6761), .Z(n6724) );
  XOR U9163 ( .A(n6723), .B(n6724), .Z(n6716) );
  NAND U9164 ( .A(n6618), .B(n6617), .Z(n6622) );
  NAND U9165 ( .A(n6620), .B(n6619), .Z(n6621) );
  NAND U9166 ( .A(n6622), .B(n6621), .Z(n6715) );
  XOR U9167 ( .A(n6716), .B(n6715), .Z(n6718) );
  XNOR U9168 ( .A(n6717), .B(n6718), .Z(n6711) );
  IV U9169 ( .A(n6651), .Z(n6733) );
  NANDN U9170 ( .A(n6733), .B(n6623), .Z(n6627) );
  NANDN U9171 ( .A(n6625), .B(n6624), .Z(n6626) );
  AND U9172 ( .A(n6627), .B(n6626), .Z(n6754) );
  AND U9173 ( .A(x[494]), .B(y[7728]), .Z(n7574) );
  NAND U9174 ( .A(n7574), .B(n6628), .Z(n6632) );
  NANDN U9175 ( .A(n6630), .B(n6629), .Z(n6631) );
  AND U9176 ( .A(n6632), .B(n6631), .Z(n6782) );
  AND U9177 ( .A(x[491]), .B(y[7726]), .Z(n6800) );
  AND U9178 ( .A(x[492]), .B(y[7725]), .Z(n6799) );
  NAND U9179 ( .A(x[487]), .B(y[7730]), .Z(n6798) );
  XOR U9180 ( .A(n6799), .B(n6798), .Z(n6801) );
  XOR U9181 ( .A(n6800), .B(n6801), .Z(n6780) );
  NAND U9182 ( .A(x[504]), .B(y[7713]), .Z(n6797) );
  XNOR U9183 ( .A(o[57]), .B(n6797), .Z(n6767) );
  NAND U9184 ( .A(x[481]), .B(y[7736]), .Z(n6768) );
  XNOR U9185 ( .A(n6767), .B(n6768), .Z(n6769) );
  NAND U9186 ( .A(x[493]), .B(y[7724]), .Z(n6770) );
  XNOR U9187 ( .A(n6769), .B(n6770), .Z(n6779) );
  XNOR U9188 ( .A(n6780), .B(n6779), .Z(n6781) );
  XNOR U9189 ( .A(n6782), .B(n6781), .Z(n6753) );
  XNOR U9190 ( .A(n6754), .B(n6753), .Z(n6755) );
  AND U9191 ( .A(n6634), .B(n6633), .Z(n6638) );
  NAND U9192 ( .A(n6636), .B(n6635), .Z(n6637) );
  NANDN U9193 ( .A(n6638), .B(n6637), .Z(n6743) );
  AND U9194 ( .A(n6640), .B(n6639), .Z(n6644) );
  NAND U9195 ( .A(n6642), .B(n6641), .Z(n6643) );
  NANDN U9196 ( .A(n6644), .B(n6643), .Z(n6744) );
  XOR U9197 ( .A(n6743), .B(n6744), .Z(n6745) );
  NAND U9198 ( .A(n6646), .B(n6645), .Z(n6650) );
  NAND U9199 ( .A(n6648), .B(n6647), .Z(n6649) );
  NAND U9200 ( .A(n6650), .B(n6649), .Z(n6741) );
  AND U9201 ( .A(x[488]), .B(y[7729]), .Z(n6736) );
  XOR U9202 ( .A(n6734), .B(n6651), .Z(n6735) );
  XOR U9203 ( .A(n6736), .B(n6735), .Z(n6739) );
  ANDN U9204 ( .B(o[56]), .A(n6652), .Z(n6730) );
  AND U9205 ( .A(x[505]), .B(y[7712]), .Z(n6728) );
  NAND U9206 ( .A(x[480]), .B(y[7737]), .Z(n6727) );
  XNOR U9207 ( .A(n6728), .B(n6727), .Z(n6729) );
  XOR U9208 ( .A(n6730), .B(n6729), .Z(n6740) );
  XNOR U9209 ( .A(n6739), .B(n6740), .Z(n6742) );
  XOR U9210 ( .A(n6741), .B(n6742), .Z(n6746) );
  XOR U9211 ( .A(n6745), .B(n6746), .Z(n6756) );
  XOR U9212 ( .A(n6755), .B(n6756), .Z(n6841) );
  NAND U9213 ( .A(n6654), .B(n6653), .Z(n6658) );
  ANDN U9214 ( .B(n6656), .A(n6655), .Z(n6657) );
  ANDN U9215 ( .B(n6658), .A(n6657), .Z(n6818) );
  NANDN U9216 ( .A(n6660), .B(n6659), .Z(n6664) );
  NANDN U9217 ( .A(n6662), .B(n6661), .Z(n6663) );
  AND U9218 ( .A(n6664), .B(n6663), .Z(n6816) );
  AND U9219 ( .A(x[494]), .B(y[7723]), .Z(n6773) );
  NAND U9220 ( .A(x[482]), .B(y[7735]), .Z(n6774) );
  NAND U9221 ( .A(x[483]), .B(y[7734]), .Z(n6776) );
  XNOR U9222 ( .A(n6816), .B(n6815), .Z(n6817) );
  XOR U9223 ( .A(n6818), .B(n6817), .Z(n6839) );
  NANDN U9224 ( .A(n6666), .B(n6665), .Z(n6670) );
  NANDN U9225 ( .A(n6668), .B(n6667), .Z(n6669) );
  AND U9226 ( .A(n6670), .B(n6669), .Z(n6840) );
  XOR U9227 ( .A(n6839), .B(n6840), .Z(n6842) );
  XOR U9228 ( .A(n6841), .B(n6842), .Z(n6833) );
  NANDN U9229 ( .A(n6672), .B(n6671), .Z(n6676) );
  NAND U9230 ( .A(n6674), .B(n6673), .Z(n6675) );
  NAND U9231 ( .A(n6676), .B(n6675), .Z(n6834) );
  XNOR U9232 ( .A(n6833), .B(n6834), .Z(n6835) );
  NANDN U9233 ( .A(n6678), .B(n6677), .Z(n6682) );
  OR U9234 ( .A(n6680), .B(n6679), .Z(n6681) );
  NAND U9235 ( .A(n6682), .B(n6681), .Z(n6836) );
  XOR U9236 ( .A(n6835), .B(n6836), .Z(n6709) );
  NAND U9237 ( .A(n6684), .B(n6683), .Z(n6688) );
  NAND U9238 ( .A(n6686), .B(n6685), .Z(n6687) );
  AND U9239 ( .A(n6688), .B(n6687), .Z(n6710) );
  XNOR U9240 ( .A(n6709), .B(n6710), .Z(n6712) );
  NAND U9241 ( .A(n6690), .B(n6689), .Z(n6694) );
  NAND U9242 ( .A(n6692), .B(n6691), .Z(n6693) );
  NAND U9243 ( .A(n6694), .B(n6693), .Z(n6852) );
  XOR U9244 ( .A(n6853), .B(n6852), .Z(n6854) );
  XNOR U9245 ( .A(n6855), .B(n6854), .Z(n6848) );
  OR U9246 ( .A(n6697), .B(n6695), .Z(n6701) );
  ANDN U9247 ( .B(n6697), .A(n6696), .Z(n6699) );
  OR U9248 ( .A(n6699), .B(n6698), .Z(n6700) );
  AND U9249 ( .A(n6701), .B(n6700), .Z(n6846) );
  NAND U9250 ( .A(n6703), .B(n6702), .Z(n6707) );
  NAND U9251 ( .A(n6705), .B(n6704), .Z(n6706) );
  AND U9252 ( .A(n6707), .B(n6706), .Z(n6847) );
  IV U9253 ( .A(n6847), .Z(n6845) );
  XOR U9254 ( .A(n6846), .B(n6845), .Z(n6708) );
  XNOR U9255 ( .A(n6848), .B(n6708), .Z(N122) );
  NAND U9256 ( .A(n6710), .B(n6709), .Z(n6714) );
  NANDN U9257 ( .A(n6712), .B(n6711), .Z(n6713) );
  NAND U9258 ( .A(n6714), .B(n6713), .Z(n7005) );
  NAND U9259 ( .A(n6716), .B(n6715), .Z(n6720) );
  NAND U9260 ( .A(n6718), .B(n6717), .Z(n6719) );
  AND U9261 ( .A(n6720), .B(n6719), .Z(n7006) );
  XOR U9262 ( .A(n7005), .B(n7006), .Z(n7008) );
  NANDN U9263 ( .A(n6722), .B(n6721), .Z(n6726) );
  NANDN U9264 ( .A(n6724), .B(n6723), .Z(n6725) );
  AND U9265 ( .A(n6726), .B(n6725), .Z(n6868) );
  AND U9266 ( .A(x[482]), .B(y[7736]), .Z(n6927) );
  XOR U9267 ( .A(n6928), .B(n6927), .Z(n6930) );
  NAND U9268 ( .A(x[504]), .B(y[7714]), .Z(n6929) );
  XNOR U9269 ( .A(n6930), .B(n6929), .Z(n6883) );
  NANDN U9270 ( .A(n6728), .B(n6727), .Z(n6732) );
  NANDN U9271 ( .A(n6730), .B(n6729), .Z(n6731) );
  NAND U9272 ( .A(n6732), .B(n6731), .Z(n6884) );
  XNOR U9273 ( .A(n6883), .B(n6884), .Z(n6885) );
  NANDN U9274 ( .A(n6734), .B(n6733), .Z(n6738) );
  NANDN U9275 ( .A(n6736), .B(n6735), .Z(n6737) );
  NAND U9276 ( .A(n6738), .B(n6737), .Z(n6886) );
  XOR U9277 ( .A(n6885), .B(n6886), .Z(n6957) );
  XOR U9278 ( .A(n6957), .B(n6958), .Z(n6960) );
  XOR U9279 ( .A(n6960), .B(n6959), .Z(n7002) );
  NAND U9280 ( .A(n6748), .B(n6747), .Z(n6752) );
  NAND U9281 ( .A(n6750), .B(n6749), .Z(n6751) );
  AND U9282 ( .A(n6752), .B(n6751), .Z(n7000) );
  NANDN U9283 ( .A(n6754), .B(n6753), .Z(n6758) );
  NANDN U9284 ( .A(n6756), .B(n6755), .Z(n6757) );
  AND U9285 ( .A(n6758), .B(n6757), .Z(n6999) );
  XNOR U9286 ( .A(n7000), .B(n6999), .Z(n7001) );
  XOR U9287 ( .A(n7002), .B(n7001), .Z(n6866) );
  NANDN U9288 ( .A(n6760), .B(n6759), .Z(n6764) );
  NANDN U9289 ( .A(n6762), .B(n6761), .Z(n6763) );
  AND U9290 ( .A(n6764), .B(n6763), .Z(n6874) );
  AND U9291 ( .A(y[7732]), .B(x[486]), .Z(n6766) );
  NAND U9292 ( .A(y[7730]), .B(x[488]), .Z(n6765) );
  XNOR U9293 ( .A(n6766), .B(n6765), .Z(n6988) );
  NAND U9294 ( .A(x[489]), .B(y[7729]), .Z(n6989) );
  XNOR U9295 ( .A(n6988), .B(n6989), .Z(n6962) );
  AND U9296 ( .A(x[487]), .B(y[7731]), .Z(n6961) );
  XOR U9297 ( .A(n6962), .B(n6961), .Z(n6964) );
  AND U9298 ( .A(x[492]), .B(y[7726]), .Z(n7069) );
  AND U9299 ( .A(x[485]), .B(y[7733]), .Z(n6898) );
  XOR U9300 ( .A(n7069), .B(n6898), .Z(n6900) );
  AND U9301 ( .A(x[490]), .B(y[7728]), .Z(n6899) );
  XOR U9302 ( .A(n6900), .B(n6899), .Z(n6963) );
  XOR U9303 ( .A(n6964), .B(n6963), .Z(n6954) );
  NANDN U9304 ( .A(n6768), .B(n6767), .Z(n6772) );
  NANDN U9305 ( .A(n6770), .B(n6769), .Z(n6771) );
  AND U9306 ( .A(n6772), .B(n6771), .Z(n6952) );
  NANDN U9307 ( .A(n6774), .B(n6773), .Z(n6778) );
  NANDN U9308 ( .A(n6776), .B(n6775), .Z(n6777) );
  NAND U9309 ( .A(n6778), .B(n6777), .Z(n6951) );
  XOR U9310 ( .A(n6954), .B(n6953), .Z(n6910) );
  NANDN U9311 ( .A(n6780), .B(n6779), .Z(n6784) );
  NANDN U9312 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U9313 ( .A(n6784), .B(n6783), .Z(n6909) );
  NANDN U9314 ( .A(n6786), .B(n6785), .Z(n6790) );
  OR U9315 ( .A(n6788), .B(n6787), .Z(n6789) );
  AND U9316 ( .A(n6790), .B(n6789), .Z(n6915) );
  NANDN U9317 ( .A(n6792), .B(n6791), .Z(n6796) );
  OR U9318 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U9319 ( .A(n6796), .B(n6795), .Z(n6916) );
  XNOR U9320 ( .A(n6915), .B(n6916), .Z(n6918) );
  ANDN U9321 ( .B(o[57]), .A(n6797), .Z(n6981) );
  NAND U9322 ( .A(x[494]), .B(y[7724]), .Z(n6982) );
  XNOR U9323 ( .A(n6981), .B(n6982), .Z(n6983) );
  NAND U9324 ( .A(x[481]), .B(y[7737]), .Z(n6984) );
  XNOR U9325 ( .A(n6983), .B(n6984), .Z(n6889) );
  NAND U9326 ( .A(x[505]), .B(y[7713]), .Z(n6992) );
  XNOR U9327 ( .A(o[58]), .B(n6992), .Z(n6903) );
  NAND U9328 ( .A(x[506]), .B(y[7712]), .Z(n6904) );
  XNOR U9329 ( .A(n6903), .B(n6904), .Z(n6905) );
  NAND U9330 ( .A(x[480]), .B(y[7738]), .Z(n6906) );
  XOR U9331 ( .A(n6905), .B(n6906), .Z(n6890) );
  XNOR U9332 ( .A(n6889), .B(n6890), .Z(n6891) );
  NANDN U9333 ( .A(n6799), .B(n6798), .Z(n6803) );
  OR U9334 ( .A(n6801), .B(n6800), .Z(n6802) );
  NAND U9335 ( .A(n6803), .B(n6802), .Z(n6892) );
  XNOR U9336 ( .A(n6891), .B(n6892), .Z(n6917) );
  XOR U9337 ( .A(n6918), .B(n6917), .Z(n6880) );
  AND U9338 ( .A(x[501]), .B(y[7717]), .Z(n6975) );
  NANDN U9339 ( .A(n6804), .B(n6975), .Z(n6808) );
  NANDN U9340 ( .A(n6806), .B(n6805), .Z(n6807) );
  AND U9341 ( .A(n6808), .B(n6807), .Z(n6948) );
  XOR U9342 ( .A(n6976), .B(n6975), .Z(n6978) );
  NAND U9343 ( .A(x[500]), .B(y[7718]), .Z(n6977) );
  XNOR U9344 ( .A(n6978), .B(n6977), .Z(n6945) );
  NAND U9345 ( .A(x[503]), .B(y[7715]), .Z(n6934) );
  XNOR U9346 ( .A(n6933), .B(n6934), .Z(n6935) );
  NAND U9347 ( .A(x[502]), .B(y[7716]), .Z(n6936) );
  XOR U9348 ( .A(n6935), .B(n6936), .Z(n6946) );
  AND U9349 ( .A(x[484]), .B(y[7734]), .Z(n6939) );
  XOR U9350 ( .A(n6940), .B(n6939), .Z(n6942) );
  AND U9351 ( .A(x[491]), .B(y[7727]), .Z(n6967) );
  NAND U9352 ( .A(x[483]), .B(y[7735]), .Z(n6968) );
  XNOR U9353 ( .A(n6967), .B(n6968), .Z(n6969) );
  NAND U9354 ( .A(x[499]), .B(y[7719]), .Z(n6970) );
  XOR U9355 ( .A(n6969), .B(n6970), .Z(n6922) );
  XNOR U9356 ( .A(n6921), .B(n6922), .Z(n6924) );
  NANDN U9357 ( .A(n6810), .B(n6809), .Z(n6814) );
  OR U9358 ( .A(n6812), .B(n6811), .Z(n6813) );
  AND U9359 ( .A(n6814), .B(n6813), .Z(n6923) );
  XNOR U9360 ( .A(n6924), .B(n6923), .Z(n6877) );
  XOR U9361 ( .A(n6878), .B(n6877), .Z(n6879) );
  XOR U9362 ( .A(n6912), .B(n6911), .Z(n6872) );
  NANDN U9363 ( .A(n6816), .B(n6815), .Z(n6820) );
  NANDN U9364 ( .A(n6818), .B(n6817), .Z(n6819) );
  NAND U9365 ( .A(n6820), .B(n6819), .Z(n6995) );
  NANDN U9366 ( .A(n6822), .B(n6821), .Z(n6826) );
  NANDN U9367 ( .A(n6824), .B(n6823), .Z(n6825) );
  NAND U9368 ( .A(n6826), .B(n6825), .Z(n6994) );
  NANDN U9369 ( .A(n6828), .B(n6827), .Z(n6832) );
  OR U9370 ( .A(n6830), .B(n6829), .Z(n6831) );
  NAND U9371 ( .A(n6832), .B(n6831), .Z(n6993) );
  XOR U9372 ( .A(n6994), .B(n6993), .Z(n6996) );
  XOR U9373 ( .A(n6995), .B(n6996), .Z(n6871) );
  XNOR U9374 ( .A(n6872), .B(n6871), .Z(n6873) );
  XNOR U9375 ( .A(n6874), .B(n6873), .Z(n6865) );
  XNOR U9376 ( .A(n6866), .B(n6865), .Z(n6867) );
  XNOR U9377 ( .A(n6868), .B(n6867), .Z(n6861) );
  NANDN U9378 ( .A(n6834), .B(n6833), .Z(n6838) );
  NANDN U9379 ( .A(n6836), .B(n6835), .Z(n6837) );
  AND U9380 ( .A(n6838), .B(n6837), .Z(n6859) );
  NAND U9381 ( .A(n6840), .B(n6839), .Z(n6844) );
  NAND U9382 ( .A(n6842), .B(n6841), .Z(n6843) );
  NAND U9383 ( .A(n6844), .B(n6843), .Z(n6860) );
  XOR U9384 ( .A(n6859), .B(n6860), .Z(n6862) );
  XNOR U9385 ( .A(n6861), .B(n6862), .Z(n7007) );
  XNOR U9386 ( .A(n7008), .B(n7007), .Z(n7013) );
  NANDN U9387 ( .A(n6845), .B(n6846), .Z(n6851) );
  NOR U9388 ( .A(n6847), .B(n6846), .Z(n6849) );
  OR U9389 ( .A(n6849), .B(n6848), .Z(n6850) );
  AND U9390 ( .A(n6851), .B(n6850), .Z(n7011) );
  NAND U9391 ( .A(n6853), .B(n6852), .Z(n6857) );
  NAND U9392 ( .A(n6855), .B(n6854), .Z(n6856) );
  AND U9393 ( .A(n6857), .B(n6856), .Z(n7012) );
  XOR U9394 ( .A(n7011), .B(n7012), .Z(n6858) );
  XNOR U9395 ( .A(n7013), .B(n6858), .Z(N123) );
  NANDN U9396 ( .A(n6860), .B(n6859), .Z(n6864) );
  NANDN U9397 ( .A(n6862), .B(n6861), .Z(n6863) );
  AND U9398 ( .A(n6864), .B(n6863), .Z(n7165) );
  NANDN U9399 ( .A(n6866), .B(n6865), .Z(n6870) );
  NANDN U9400 ( .A(n6868), .B(n6867), .Z(n6869) );
  AND U9401 ( .A(n6870), .B(n6869), .Z(n7163) );
  NANDN U9402 ( .A(n6872), .B(n6871), .Z(n6876) );
  NANDN U9403 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U9404 ( .A(n6876), .B(n6875), .Z(n7024) );
  NAND U9405 ( .A(n6878), .B(n6877), .Z(n6882) );
  NANDN U9406 ( .A(n6880), .B(n6879), .Z(n6881) );
  AND U9407 ( .A(n6882), .B(n6881), .Z(n7145) );
  NANDN U9408 ( .A(n6884), .B(n6883), .Z(n6888) );
  NANDN U9409 ( .A(n6886), .B(n6885), .Z(n6887) );
  AND U9410 ( .A(n6888), .B(n6887), .Z(n7134) );
  NANDN U9411 ( .A(n6890), .B(n6889), .Z(n6894) );
  NANDN U9412 ( .A(n6892), .B(n6891), .Z(n6893) );
  AND U9413 ( .A(n6894), .B(n6893), .Z(n7133) );
  AND U9414 ( .A(x[499]), .B(y[7720]), .Z(n7105) );
  NAND U9415 ( .A(x[505]), .B(y[7714]), .Z(n7106) );
  XNOR U9416 ( .A(n7105), .B(n7106), .Z(n7107) );
  NAND U9417 ( .A(x[486]), .B(y[7733]), .Z(n7108) );
  XNOR U9418 ( .A(n7107), .B(n7108), .Z(n7094) );
  AND U9419 ( .A(x[495]), .B(y[7724]), .Z(n7074) );
  NAND U9420 ( .A(x[482]), .B(y[7737]), .Z(n7075) );
  NAND U9421 ( .A(x[483]), .B(y[7736]), .Z(n7077) );
  XNOR U9422 ( .A(n7094), .B(n7095), .Z(n7096) );
  NAND U9423 ( .A(x[496]), .B(y[7723]), .Z(n7057) );
  XNOR U9424 ( .A(n7057), .B(n7058), .Z(n7059) );
  XNOR U9425 ( .A(n6895), .B(n7059), .Z(n7070) );
  AND U9426 ( .A(y[7726]), .B(x[493]), .Z(n6897) );
  NAND U9427 ( .A(y[7727]), .B(x[492]), .Z(n6896) );
  XNOR U9428 ( .A(n6897), .B(n6896), .Z(n7071) );
  XNOR U9429 ( .A(n7070), .B(n7071), .Z(n7097) );
  XNOR U9430 ( .A(n7096), .B(n7097), .Z(n7035) );
  NAND U9431 ( .A(n7069), .B(n6898), .Z(n6902) );
  AND U9432 ( .A(n6900), .B(n6899), .Z(n6901) );
  ANDN U9433 ( .B(n6902), .A(n6901), .Z(n7034) );
  NANDN U9434 ( .A(n6904), .B(n6903), .Z(n6908) );
  NANDN U9435 ( .A(n6906), .B(n6905), .Z(n6907) );
  NAND U9436 ( .A(n6908), .B(n6907), .Z(n7033) );
  XOR U9437 ( .A(n7034), .B(n7033), .Z(n7036) );
  XNOR U9438 ( .A(n7035), .B(n7036), .Z(n7132) );
  XOR U9439 ( .A(n7133), .B(n7132), .Z(n7135) );
  XOR U9440 ( .A(n7134), .B(n7135), .Z(n7144) );
  XOR U9441 ( .A(n7145), .B(n7144), .Z(n7147) );
  NANDN U9442 ( .A(n6910), .B(n6909), .Z(n6914) );
  NAND U9443 ( .A(n6912), .B(n6911), .Z(n6913) );
  AND U9444 ( .A(n6914), .B(n6913), .Z(n7146) );
  XOR U9445 ( .A(n7147), .B(n7146), .Z(n7022) );
  NANDN U9446 ( .A(n6916), .B(n6915), .Z(n6920) );
  NAND U9447 ( .A(n6918), .B(n6917), .Z(n6919) );
  AND U9448 ( .A(n6920), .B(n6919), .Z(n7141) );
  NANDN U9449 ( .A(n6922), .B(n6921), .Z(n6926) );
  NAND U9450 ( .A(n6924), .B(n6923), .Z(n6925) );
  AND U9451 ( .A(n6926), .B(n6925), .Z(n7139) );
  NAND U9452 ( .A(n6928), .B(n6927), .Z(n6932) );
  ANDN U9453 ( .B(n6930), .A(n6929), .Z(n6931) );
  ANDN U9454 ( .B(n6932), .A(n6931), .Z(n7040) );
  NANDN U9455 ( .A(n6934), .B(n6933), .Z(n6938) );
  NANDN U9456 ( .A(n6936), .B(n6935), .Z(n6937) );
  NAND U9457 ( .A(n6938), .B(n6937), .Z(n7039) );
  XNOR U9458 ( .A(n7040), .B(n7039), .Z(n7041) );
  NAND U9459 ( .A(n6940), .B(n6939), .Z(n6944) );
  ANDN U9460 ( .B(n6942), .A(n6941), .Z(n6943) );
  ANDN U9461 ( .B(n6944), .A(n6943), .Z(n7054) );
  AND U9462 ( .A(x[480]), .B(y[7739]), .Z(n7117) );
  NAND U9463 ( .A(x[507]), .B(y[7712]), .Z(n7118) );
  XNOR U9464 ( .A(n7117), .B(n7118), .Z(n7119) );
  AND U9465 ( .A(x[506]), .B(y[7713]), .Z(n7129) );
  XNOR U9466 ( .A(o[59]), .B(n7129), .Z(n7120) );
  XNOR U9467 ( .A(n7119), .B(n7120), .Z(n7051) );
  AND U9468 ( .A(x[489]), .B(y[7730]), .Z(n7123) );
  NAND U9469 ( .A(x[501]), .B(y[7718]), .Z(n7124) );
  XNOR U9470 ( .A(n7123), .B(n7124), .Z(n7125) );
  NAND U9471 ( .A(x[498]), .B(y[7721]), .Z(n7126) );
  XOR U9472 ( .A(n7125), .B(n7126), .Z(n7052) );
  XNOR U9473 ( .A(n7051), .B(n7052), .Z(n7053) );
  XOR U9474 ( .A(n7054), .B(n7053), .Z(n7042) );
  XNOR U9475 ( .A(n7041), .B(n7042), .Z(n7138) );
  XNOR U9476 ( .A(n7139), .B(n7138), .Z(n7140) );
  XOR U9477 ( .A(n7141), .B(n7140), .Z(n7152) );
  NANDN U9478 ( .A(n6946), .B(n6945), .Z(n6950) );
  NANDN U9479 ( .A(n6948), .B(n6947), .Z(n6949) );
  AND U9480 ( .A(n6950), .B(n6949), .Z(n7151) );
  NANDN U9481 ( .A(n6952), .B(n6951), .Z(n6956) );
  NAND U9482 ( .A(n6954), .B(n6953), .Z(n6955) );
  AND U9483 ( .A(n6956), .B(n6955), .Z(n7150) );
  XOR U9484 ( .A(n7151), .B(n7150), .Z(n7153) );
  XOR U9485 ( .A(n7152), .B(n7153), .Z(n7021) );
  XNOR U9486 ( .A(n7024), .B(n7023), .Z(n7018) );
  NAND U9487 ( .A(n6962), .B(n6961), .Z(n6966) );
  NAND U9488 ( .A(n6964), .B(n6963), .Z(n6965) );
  AND U9489 ( .A(n6966), .B(n6965), .Z(n7158) );
  NANDN U9490 ( .A(n6968), .B(n6967), .Z(n6972) );
  NANDN U9491 ( .A(n6970), .B(n6969), .Z(n6971) );
  AND U9492 ( .A(n6972), .B(n6971), .Z(n7093) );
  AND U9493 ( .A(y[7715]), .B(x[504]), .Z(n6974) );
  NAND U9494 ( .A(y[7719]), .B(x[500]), .Z(n6973) );
  XNOR U9495 ( .A(n6974), .B(n6973), .Z(n7101) );
  NAND U9496 ( .A(x[487]), .B(y[7732]), .Z(n7102) );
  XNOR U9497 ( .A(n7101), .B(n7102), .Z(n7091) );
  AND U9498 ( .A(x[488]), .B(y[7731]), .Z(n7063) );
  AND U9499 ( .A(x[503]), .B(y[7716]), .Z(n7064) );
  XOR U9500 ( .A(n7063), .B(n7064), .Z(n7065) );
  AND U9501 ( .A(x[502]), .B(y[7717]), .Z(n7066) );
  XOR U9502 ( .A(n7065), .B(n7066), .Z(n7090) );
  XOR U9503 ( .A(n7091), .B(n7090), .Z(n7092) );
  XOR U9504 ( .A(n7093), .B(n7092), .Z(n7156) );
  NAND U9505 ( .A(n6976), .B(n6975), .Z(n6980) );
  ANDN U9506 ( .B(n6978), .A(n6977), .Z(n6979) );
  ANDN U9507 ( .B(n6980), .A(n6979), .Z(n7087) );
  NANDN U9508 ( .A(n6982), .B(n6981), .Z(n6986) );
  NANDN U9509 ( .A(n6984), .B(n6983), .Z(n6985) );
  NAND U9510 ( .A(n6986), .B(n6985), .Z(n7086) );
  XNOR U9511 ( .A(n7087), .B(n7086), .Z(n7089) );
  AND U9512 ( .A(y[7732]), .B(x[488]), .Z(n7131) );
  NAND U9513 ( .A(n6987), .B(n7131), .Z(n6991) );
  NANDN U9514 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U9515 ( .A(n6991), .B(n6990), .Z(n7047) );
  AND U9516 ( .A(x[494]), .B(y[7725]), .Z(n7080) );
  NAND U9517 ( .A(x[481]), .B(y[7738]), .Z(n7081) );
  ANDN U9518 ( .B(o[58]), .A(n6992), .Z(n7082) );
  XOR U9519 ( .A(n7083), .B(n7082), .Z(n7046) );
  AND U9520 ( .A(x[497]), .B(y[7722]), .Z(n7111) );
  NAND U9521 ( .A(x[484]), .B(y[7735]), .Z(n7112) );
  XNOR U9522 ( .A(n7111), .B(n7112), .Z(n7114) );
  AND U9523 ( .A(x[485]), .B(y[7734]), .Z(n7113) );
  XOR U9524 ( .A(n7114), .B(n7113), .Z(n7045) );
  XOR U9525 ( .A(n7046), .B(n7045), .Z(n7048) );
  XOR U9526 ( .A(n7047), .B(n7048), .Z(n7088) );
  XOR U9527 ( .A(n7089), .B(n7088), .Z(n7157) );
  XNOR U9528 ( .A(n7158), .B(n7159), .Z(n7028) );
  XOR U9529 ( .A(n7027), .B(n7028), .Z(n7030) );
  NAND U9530 ( .A(n6994), .B(n6993), .Z(n6998) );
  NAND U9531 ( .A(n6996), .B(n6995), .Z(n6997) );
  AND U9532 ( .A(n6998), .B(n6997), .Z(n7029) );
  XNOR U9533 ( .A(n7030), .B(n7029), .Z(n7016) );
  NANDN U9534 ( .A(n7000), .B(n6999), .Z(n7004) );
  NAND U9535 ( .A(n7002), .B(n7001), .Z(n7003) );
  AND U9536 ( .A(n7004), .B(n7003), .Z(n7015) );
  XOR U9537 ( .A(n7016), .B(n7015), .Z(n7017) );
  XOR U9538 ( .A(n7018), .B(n7017), .Z(n7162) );
  XNOR U9539 ( .A(n7163), .B(n7162), .Z(n7164) );
  XNOR U9540 ( .A(n7165), .B(n7164), .Z(n7170) );
  NAND U9541 ( .A(n7006), .B(n7005), .Z(n7010) );
  NAND U9542 ( .A(n7008), .B(n7007), .Z(n7009) );
  AND U9543 ( .A(n7010), .B(n7009), .Z(n7169) );
  XNOR U9544 ( .A(n7169), .B(n7168), .Z(n7014) );
  XNOR U9545 ( .A(n7170), .B(n7014), .Z(N124) );
  NAND U9546 ( .A(n7016), .B(n7015), .Z(n7020) );
  NAND U9547 ( .A(n7018), .B(n7017), .Z(n7019) );
  NAND U9548 ( .A(n7020), .B(n7019), .Z(n7333) );
  NANDN U9549 ( .A(n7022), .B(n7021), .Z(n7026) );
  NAND U9550 ( .A(n7024), .B(n7023), .Z(n7025) );
  AND U9551 ( .A(n7026), .B(n7025), .Z(n7332) );
  XOR U9552 ( .A(n7333), .B(n7332), .Z(n7335) );
  NAND U9553 ( .A(n7028), .B(n7027), .Z(n7032) );
  NAND U9554 ( .A(n7030), .B(n7029), .Z(n7031) );
  AND U9555 ( .A(n7032), .B(n7031), .Z(n7173) );
  NANDN U9556 ( .A(n7034), .B(n7033), .Z(n7038) );
  NANDN U9557 ( .A(n7036), .B(n7035), .Z(n7037) );
  AND U9558 ( .A(n7038), .B(n7037), .Z(n7197) );
  NANDN U9559 ( .A(n7040), .B(n7039), .Z(n7044) );
  NANDN U9560 ( .A(n7042), .B(n7041), .Z(n7043) );
  AND U9561 ( .A(n7044), .B(n7043), .Z(n7302) );
  NAND U9562 ( .A(n7046), .B(n7045), .Z(n7050) );
  NAND U9563 ( .A(n7048), .B(n7047), .Z(n7049) );
  AND U9564 ( .A(n7050), .B(n7049), .Z(n7300) );
  NANDN U9565 ( .A(n7052), .B(n7051), .Z(n7056) );
  NANDN U9566 ( .A(n7054), .B(n7053), .Z(n7055) );
  NAND U9567 ( .A(n7056), .B(n7055), .Z(n7299) );
  XNOR U9568 ( .A(n7300), .B(n7299), .Z(n7301) );
  XNOR U9569 ( .A(n7302), .B(n7301), .Z(n7196) );
  XNOR U9570 ( .A(n7197), .B(n7196), .Z(n7199) );
  NANDN U9571 ( .A(n7058), .B(n7057), .Z(n7062) );
  NANDN U9572 ( .A(n7060), .B(n7059), .Z(n7061) );
  AND U9573 ( .A(n7062), .B(n7061), .Z(n7264) );
  AND U9574 ( .A(x[487]), .B(y[7733]), .Z(n7244) );
  AND U9575 ( .A(x[492]), .B(y[7728]), .Z(n7243) );
  XOR U9576 ( .A(n7244), .B(n7243), .Z(n7246) );
  AND U9577 ( .A(x[491]), .B(y[7729]), .Z(n7245) );
  XOR U9578 ( .A(n7246), .B(n7245), .Z(n7262) );
  AND U9579 ( .A(x[507]), .B(y[7713]), .Z(n7260) );
  XOR U9580 ( .A(o[60]), .B(n7260), .Z(n7274) );
  AND U9581 ( .A(x[506]), .B(y[7714]), .Z(n7273) );
  XOR U9582 ( .A(n7274), .B(n7273), .Z(n7276) );
  AND U9583 ( .A(x[495]), .B(y[7725]), .Z(n7275) );
  XNOR U9584 ( .A(n7276), .B(n7275), .Z(n7261) );
  NAND U9585 ( .A(n7064), .B(n7063), .Z(n7068) );
  NAND U9586 ( .A(n7066), .B(n7065), .Z(n7067) );
  AND U9587 ( .A(n7068), .B(n7067), .Z(n7284) );
  AND U9588 ( .A(x[497]), .B(y[7723]), .Z(n7209) );
  AND U9589 ( .A(x[502]), .B(y[7718]), .Z(n7208) );
  XOR U9590 ( .A(n7209), .B(n7208), .Z(n7211) );
  AND U9591 ( .A(x[484]), .B(y[7736]), .Z(n7210) );
  XOR U9592 ( .A(n7211), .B(n7210), .Z(n7282) );
  AND U9593 ( .A(x[486]), .B(y[7734]), .Z(n7427) );
  NAND U9594 ( .A(x[499]), .B(y[7721]), .Z(n7249) );
  XOR U9595 ( .A(n7282), .B(n7281), .Z(n7283) );
  XOR U9596 ( .A(n7306), .B(n7305), .Z(n7307) );
  NAND U9597 ( .A(n7267), .B(n7069), .Z(n7073) );
  NAND U9598 ( .A(n7071), .B(n7070), .Z(n7072) );
  AND U9599 ( .A(n7073), .B(n7072), .Z(n7205) );
  NANDN U9600 ( .A(n7075), .B(n7074), .Z(n7079) );
  NANDN U9601 ( .A(n7077), .B(n7076), .Z(n7078) );
  AND U9602 ( .A(n7079), .B(n7078), .Z(n7203) );
  NANDN U9603 ( .A(n7081), .B(n7080), .Z(n7085) );
  NAND U9604 ( .A(n7083), .B(n7082), .Z(n7084) );
  NAND U9605 ( .A(n7085), .B(n7084), .Z(n7202) );
  XNOR U9606 ( .A(n7307), .B(n7308), .Z(n7198) );
  XOR U9607 ( .A(n7199), .B(n7198), .Z(n7192) );
  NANDN U9608 ( .A(n7095), .B(n7094), .Z(n7099) );
  NANDN U9609 ( .A(n7097), .B(n7096), .Z(n7098) );
  NAND U9610 ( .A(n7099), .B(n7098), .Z(n7287) );
  XOR U9611 ( .A(n7288), .B(n7287), .Z(n7290) );
  XOR U9612 ( .A(n7289), .B(n7290), .Z(n7191) );
  AND U9613 ( .A(x[504]), .B(y[7719]), .Z(n7605) );
  AND U9614 ( .A(x[500]), .B(y[7715]), .Z(n7100) );
  NAND U9615 ( .A(n7605), .B(n7100), .Z(n7104) );
  NANDN U9616 ( .A(n7102), .B(n7101), .Z(n7103) );
  AND U9617 ( .A(n7104), .B(n7103), .Z(n7326) );
  AND U9618 ( .A(x[505]), .B(y[7715]), .Z(n7239) );
  XOR U9619 ( .A(n7240), .B(n7239), .Z(n7238) );
  NAND U9620 ( .A(x[481]), .B(y[7739]), .Z(n7237) );
  AND U9621 ( .A(x[496]), .B(y[7724]), .Z(n7231) );
  NAND U9622 ( .A(x[504]), .B(y[7716]), .Z(n7232) );
  NAND U9623 ( .A(x[482]), .B(y[7738]), .Z(n7234) );
  XOR U9624 ( .A(n7324), .B(n7323), .Z(n7325) );
  NANDN U9625 ( .A(n7106), .B(n7105), .Z(n7110) );
  NANDN U9626 ( .A(n7108), .B(n7107), .Z(n7109) );
  AND U9627 ( .A(n7110), .B(n7109), .Z(n7320) );
  NAND U9628 ( .A(x[483]), .B(y[7737]), .Z(n7268) );
  NAND U9629 ( .A(x[503]), .B(y[7717]), .Z(n7270) );
  AND U9630 ( .A(x[485]), .B(y[7735]), .Z(n7254) );
  NAND U9631 ( .A(x[501]), .B(y[7719]), .Z(n7255) );
  NAND U9632 ( .A(x[500]), .B(y[7720]), .Z(n7257) );
  XOR U9633 ( .A(n7318), .B(n7317), .Z(n7319) );
  NANDN U9634 ( .A(n7112), .B(n7111), .Z(n7116) );
  NAND U9635 ( .A(n7114), .B(n7113), .Z(n7115) );
  AND U9636 ( .A(n7116), .B(n7115), .Z(n7312) );
  NANDN U9637 ( .A(n7118), .B(n7117), .Z(n7122) );
  NANDN U9638 ( .A(n7120), .B(n7119), .Z(n7121) );
  NAND U9639 ( .A(n7122), .B(n7121), .Z(n7311) );
  NANDN U9640 ( .A(n7124), .B(n7123), .Z(n7128) );
  NANDN U9641 ( .A(n7126), .B(n7125), .Z(n7127) );
  NAND U9642 ( .A(n7128), .B(n7127), .Z(n7227) );
  AND U9643 ( .A(n7129), .B(o[59]), .Z(n7217) );
  AND U9644 ( .A(x[480]), .B(y[7740]), .Z(n7215) );
  AND U9645 ( .A(x[508]), .B(y[7712]), .Z(n7214) );
  XOR U9646 ( .A(n7215), .B(n7214), .Z(n7216) );
  XOR U9647 ( .A(n7217), .B(n7216), .Z(n7226) );
  NAND U9648 ( .A(y[7730]), .B(x[490]), .Z(n7130) );
  XNOR U9649 ( .A(n7131), .B(n7130), .Z(n7222) );
  AND U9650 ( .A(x[489]), .B(y[7731]), .Z(n7221) );
  XOR U9651 ( .A(n7222), .B(n7221), .Z(n7225) );
  XOR U9652 ( .A(n7226), .B(n7225), .Z(n7228) );
  XOR U9653 ( .A(n7227), .B(n7228), .Z(n7313) );
  XNOR U9654 ( .A(n7314), .B(n7313), .Z(n7293) );
  XOR U9655 ( .A(n7294), .B(n7293), .Z(n7295) );
  XOR U9656 ( .A(n7296), .B(n7295), .Z(n7190) );
  XOR U9657 ( .A(n7191), .B(n7190), .Z(n7193) );
  XOR U9658 ( .A(n7192), .B(n7193), .Z(n7186) );
  NANDN U9659 ( .A(n7133), .B(n7132), .Z(n7137) );
  OR U9660 ( .A(n7135), .B(n7134), .Z(n7136) );
  AND U9661 ( .A(n7137), .B(n7136), .Z(n7185) );
  NANDN U9662 ( .A(n7139), .B(n7138), .Z(n7143) );
  NANDN U9663 ( .A(n7141), .B(n7140), .Z(n7142) );
  NAND U9664 ( .A(n7143), .B(n7142), .Z(n7184) );
  XOR U9665 ( .A(n7185), .B(n7184), .Z(n7187) );
  XOR U9666 ( .A(n7186), .B(n7187), .Z(n7172) );
  XOR U9667 ( .A(n7173), .B(n7172), .Z(n7174) );
  NAND U9668 ( .A(n7145), .B(n7144), .Z(n7149) );
  NAND U9669 ( .A(n7147), .B(n7146), .Z(n7148) );
  NAND U9670 ( .A(n7149), .B(n7148), .Z(n7180) );
  NAND U9671 ( .A(n7151), .B(n7150), .Z(n7155) );
  NAND U9672 ( .A(n7153), .B(n7152), .Z(n7154) );
  AND U9673 ( .A(n7155), .B(n7154), .Z(n7179) );
  NANDN U9674 ( .A(n7157), .B(n7156), .Z(n7161) );
  NANDN U9675 ( .A(n7159), .B(n7158), .Z(n7160) );
  AND U9676 ( .A(n7161), .B(n7160), .Z(n7178) );
  XOR U9677 ( .A(n7179), .B(n7178), .Z(n7181) );
  XNOR U9678 ( .A(n7180), .B(n7181), .Z(n7175) );
  XNOR U9679 ( .A(n7335), .B(n7334), .Z(n7331) );
  NANDN U9680 ( .A(n7163), .B(n7162), .Z(n7167) );
  NANDN U9681 ( .A(n7165), .B(n7164), .Z(n7166) );
  NAND U9682 ( .A(n7167), .B(n7166), .Z(n7329) );
  XOR U9683 ( .A(n7329), .B(n7330), .Z(n7171) );
  XNOR U9684 ( .A(n7331), .B(n7171), .Z(N125) );
  NAND U9685 ( .A(n7173), .B(n7172), .Z(n7177) );
  NANDN U9686 ( .A(n7175), .B(n7174), .Z(n7176) );
  NAND U9687 ( .A(n7177), .B(n7176), .Z(n7348) );
  NAND U9688 ( .A(n7179), .B(n7178), .Z(n7183) );
  NAND U9689 ( .A(n7181), .B(n7180), .Z(n7182) );
  NAND U9690 ( .A(n7183), .B(n7182), .Z(n7346) );
  NANDN U9691 ( .A(n7185), .B(n7184), .Z(n7189) );
  OR U9692 ( .A(n7187), .B(n7186), .Z(n7188) );
  AND U9693 ( .A(n7189), .B(n7188), .Z(n7353) );
  NANDN U9694 ( .A(n7191), .B(n7190), .Z(n7195) );
  OR U9695 ( .A(n7193), .B(n7192), .Z(n7194) );
  AND U9696 ( .A(n7195), .B(n7194), .Z(n7352) );
  XNOR U9697 ( .A(n7353), .B(n7352), .Z(n7355) );
  NANDN U9698 ( .A(n7197), .B(n7196), .Z(n7201) );
  NAND U9699 ( .A(n7199), .B(n7198), .Z(n7200) );
  AND U9700 ( .A(n7201), .B(n7200), .Z(n7363) );
  NANDN U9701 ( .A(n7203), .B(n7202), .Z(n7207) );
  NANDN U9702 ( .A(n7205), .B(n7204), .Z(n7206) );
  AND U9703 ( .A(n7207), .B(n7206), .Z(n7474) );
  NAND U9704 ( .A(n7209), .B(n7208), .Z(n7213) );
  NAND U9705 ( .A(n7211), .B(n7210), .Z(n7212) );
  NAND U9706 ( .A(n7213), .B(n7212), .Z(n7511) );
  NAND U9707 ( .A(n7215), .B(n7214), .Z(n7219) );
  NAND U9708 ( .A(n7217), .B(n7216), .Z(n7218) );
  NAND U9709 ( .A(n7219), .B(n7218), .Z(n7510) );
  XOR U9710 ( .A(n7511), .B(n7510), .Z(n7512) );
  AND U9711 ( .A(y[7732]), .B(x[490]), .Z(n7508) );
  NAND U9712 ( .A(n7220), .B(n7508), .Z(n7224) );
  NAND U9713 ( .A(n7222), .B(n7221), .Z(n7223) );
  NAND U9714 ( .A(n7224), .B(n7223), .Z(n7479) );
  AND U9715 ( .A(x[502]), .B(y[7719]), .Z(n7448) );
  AND U9716 ( .A(x[492]), .B(y[7729]), .Z(n7683) );
  AND U9717 ( .A(x[481]), .B(y[7740]), .Z(n7446) );
  XOR U9718 ( .A(n7683), .B(n7446), .Z(n7447) );
  XOR U9719 ( .A(n7448), .B(n7447), .Z(n7478) );
  AND U9720 ( .A(x[495]), .B(y[7726]), .Z(n7451) );
  XOR U9721 ( .A(n7478), .B(n7477), .Z(n7480) );
  XNOR U9722 ( .A(n7479), .B(n7480), .Z(n7513) );
  NAND U9723 ( .A(n7226), .B(n7225), .Z(n7230) );
  NAND U9724 ( .A(n7228), .B(n7227), .Z(n7229) );
  AND U9725 ( .A(n7230), .B(n7229), .Z(n7471) );
  XOR U9726 ( .A(n7474), .B(n7473), .Z(n7468) );
  NANDN U9727 ( .A(n7232), .B(n7231), .Z(n7236) );
  NANDN U9728 ( .A(n7234), .B(n7233), .Z(n7235) );
  NAND U9729 ( .A(n7236), .B(n7235), .Z(n7484) );
  ANDN U9730 ( .B(n7238), .A(n7237), .Z(n7242) );
  NAND U9731 ( .A(n7240), .B(n7239), .Z(n7241) );
  NANDN U9732 ( .A(n7242), .B(n7241), .Z(n7483) );
  XOR U9733 ( .A(n7484), .B(n7483), .Z(n7485) );
  NAND U9734 ( .A(n7244), .B(n7243), .Z(n7248) );
  NAND U9735 ( .A(n7246), .B(n7245), .Z(n7247) );
  NAND U9736 ( .A(n7248), .B(n7247), .Z(n7388) );
  AND U9737 ( .A(x[491]), .B(y[7730]), .Z(n7424) );
  AND U9738 ( .A(x[483]), .B(y[7738]), .Z(n7422) );
  AND U9739 ( .A(x[497]), .B(y[7724]), .Z(n7421) );
  XOR U9740 ( .A(n7422), .B(n7421), .Z(n7423) );
  XOR U9741 ( .A(n7424), .B(n7423), .Z(n7387) );
  AND U9742 ( .A(x[503]), .B(y[7718]), .Z(n7418) );
  AND U9743 ( .A(x[493]), .B(y[7728]), .Z(n7416) );
  AND U9744 ( .A(x[504]), .B(y[7717]), .Z(n7653) );
  XOR U9745 ( .A(n7416), .B(n7653), .Z(n7417) );
  XOR U9746 ( .A(n7418), .B(n7417), .Z(n7386) );
  XOR U9747 ( .A(n7387), .B(n7386), .Z(n7389) );
  XNOR U9748 ( .A(n7388), .B(n7389), .Z(n7486) );
  NANDN U9749 ( .A(n7249), .B(n7427), .Z(n7253) );
  NANDN U9750 ( .A(n7251), .B(n7250), .Z(n7252) );
  AND U9751 ( .A(n7253), .B(n7252), .Z(n7491) );
  AND U9752 ( .A(x[505]), .B(y[7716]), .Z(n7443) );
  AND U9753 ( .A(x[506]), .B(y[7715]), .Z(n7440) );
  XOR U9754 ( .A(n7441), .B(n7440), .Z(n7442) );
  XOR U9755 ( .A(n7443), .B(n7442), .Z(n7490) );
  AND U9756 ( .A(x[508]), .B(y[7713]), .Z(n7458) );
  XOR U9757 ( .A(o[61]), .B(n7458), .Z(n7503) );
  AND U9758 ( .A(x[480]), .B(y[7741]), .Z(n7501) );
  AND U9759 ( .A(x[509]), .B(y[7712]), .Z(n7500) );
  XOR U9760 ( .A(n7501), .B(n7500), .Z(n7502) );
  XNOR U9761 ( .A(n7503), .B(n7502), .Z(n7489) );
  XNOR U9762 ( .A(n7491), .B(n7492), .Z(n7374) );
  NANDN U9763 ( .A(n7255), .B(n7254), .Z(n7259) );
  NANDN U9764 ( .A(n7257), .B(n7256), .Z(n7258) );
  NAND U9765 ( .A(n7259), .B(n7258), .Z(n7436) );
  AND U9766 ( .A(x[482]), .B(y[7739]), .Z(n7399) );
  XOR U9767 ( .A(n7399), .B(n7398), .Z(n7400) );
  XOR U9768 ( .A(n7401), .B(n7400), .Z(n7435) );
  AND U9769 ( .A(o[60]), .B(n7260), .Z(n7407) );
  AND U9770 ( .A(x[496]), .B(y[7725]), .Z(n7405) );
  AND U9771 ( .A(x[507]), .B(y[7714]), .Z(n7404) );
  XOR U9772 ( .A(n7405), .B(n7404), .Z(n7406) );
  XOR U9773 ( .A(n7407), .B(n7406), .Z(n7434) );
  XOR U9774 ( .A(n7435), .B(n7434), .Z(n7437) );
  XOR U9775 ( .A(n7436), .B(n7437), .Z(n7375) );
  NANDN U9776 ( .A(n7262), .B(n7261), .Z(n7266) );
  NANDN U9777 ( .A(n7264), .B(n7263), .Z(n7265) );
  AND U9778 ( .A(n7266), .B(n7265), .Z(n7381) );
  NANDN U9779 ( .A(n7268), .B(n7267), .Z(n7272) );
  NANDN U9780 ( .A(n7270), .B(n7269), .Z(n7271) );
  NAND U9781 ( .A(n7272), .B(n7271), .Z(n7411) );
  NAND U9782 ( .A(n7274), .B(n7273), .Z(n7278) );
  NAND U9783 ( .A(n7276), .B(n7275), .Z(n7277) );
  NAND U9784 ( .A(n7278), .B(n7277), .Z(n7410) );
  XOR U9785 ( .A(n7411), .B(n7410), .Z(n7413) );
  AND U9786 ( .A(x[485]), .B(y[7736]), .Z(n7395) );
  AND U9787 ( .A(x[484]), .B(y[7737]), .Z(n7393) );
  AND U9788 ( .A(x[490]), .B(y[7731]), .Z(n7392) );
  XOR U9789 ( .A(n7393), .B(n7392), .Z(n7394) );
  XOR U9790 ( .A(n7395), .B(n7394), .Z(n7497) );
  AND U9791 ( .A(x[489]), .B(y[7732]), .Z(n7621) );
  AND U9792 ( .A(x[488]), .B(y[7733]), .Z(n7429) );
  AND U9793 ( .A(x[486]), .B(y[7735]), .Z(n7280) );
  AND U9794 ( .A(y[7734]), .B(x[487]), .Z(n7279) );
  XOR U9795 ( .A(n7280), .B(n7279), .Z(n7428) );
  XOR U9796 ( .A(n7429), .B(n7428), .Z(n7495) );
  XOR U9797 ( .A(n7621), .B(n7495), .Z(n7496) );
  XOR U9798 ( .A(n7497), .B(n7496), .Z(n7412) );
  XNOR U9799 ( .A(n7413), .B(n7412), .Z(n7380) );
  XOR U9800 ( .A(n7383), .B(n7382), .Z(n7466) );
  NAND U9801 ( .A(n7282), .B(n7281), .Z(n7286) );
  NANDN U9802 ( .A(n7284), .B(n7283), .Z(n7285) );
  NAND U9803 ( .A(n7286), .B(n7285), .Z(n7465) );
  XNOR U9804 ( .A(n7363), .B(n7362), .Z(n7364) );
  NANDN U9805 ( .A(n7288), .B(n7287), .Z(n7292) );
  OR U9806 ( .A(n7290), .B(n7289), .Z(n7291) );
  AND U9807 ( .A(n7292), .B(n7291), .Z(n7357) );
  NAND U9808 ( .A(n7294), .B(n7293), .Z(n7298) );
  NAND U9809 ( .A(n7296), .B(n7295), .Z(n7297) );
  AND U9810 ( .A(n7298), .B(n7297), .Z(n7356) );
  XNOR U9811 ( .A(n7357), .B(n7356), .Z(n7358) );
  NANDN U9812 ( .A(n7300), .B(n7299), .Z(n7304) );
  NANDN U9813 ( .A(n7302), .B(n7301), .Z(n7303) );
  NAND U9814 ( .A(n7304), .B(n7303), .Z(n7370) );
  NAND U9815 ( .A(n7306), .B(n7305), .Z(n7310) );
  NANDN U9816 ( .A(n7308), .B(n7307), .Z(n7309) );
  NAND U9817 ( .A(n7310), .B(n7309), .Z(n7368) );
  NANDN U9818 ( .A(n7312), .B(n7311), .Z(n7316) );
  NAND U9819 ( .A(n7314), .B(n7313), .Z(n7315) );
  AND U9820 ( .A(n7316), .B(n7315), .Z(n7462) );
  NAND U9821 ( .A(n7318), .B(n7317), .Z(n7322) );
  NANDN U9822 ( .A(n7320), .B(n7319), .Z(n7321) );
  AND U9823 ( .A(n7322), .B(n7321), .Z(n7460) );
  NAND U9824 ( .A(n7324), .B(n7323), .Z(n7328) );
  NANDN U9825 ( .A(n7326), .B(n7325), .Z(n7327) );
  NAND U9826 ( .A(n7328), .B(n7327), .Z(n7459) );
  XOR U9827 ( .A(n7368), .B(n7369), .Z(n7371) );
  XNOR U9828 ( .A(n7370), .B(n7371), .Z(n7359) );
  XOR U9829 ( .A(n7358), .B(n7359), .Z(n7365) );
  XNOR U9830 ( .A(n7364), .B(n7365), .Z(n7354) );
  XOR U9831 ( .A(n7355), .B(n7354), .Z(n7347) );
  XOR U9832 ( .A(n7346), .B(n7347), .Z(n7349) );
  XOR U9833 ( .A(n7348), .B(n7349), .Z(n7342) );
  NAND U9834 ( .A(n7333), .B(n7332), .Z(n7337) );
  NAND U9835 ( .A(n7335), .B(n7334), .Z(n7336) );
  AND U9836 ( .A(n7337), .B(n7336), .Z(n7341) );
  IV U9837 ( .A(n7341), .Z(n7339) );
  XOR U9838 ( .A(n7340), .B(n7339), .Z(n7338) );
  XNOR U9839 ( .A(n7342), .B(n7338), .Z(N126) );
  NANDN U9840 ( .A(n7339), .B(n7340), .Z(n7345) );
  NOR U9841 ( .A(n7341), .B(n7340), .Z(n7343) );
  OR U9842 ( .A(n7343), .B(n7342), .Z(n7344) );
  AND U9843 ( .A(n7345), .B(n7344), .Z(n7804) );
  NAND U9844 ( .A(n7347), .B(n7346), .Z(n7351) );
  NAND U9845 ( .A(n7349), .B(n7348), .Z(n7350) );
  AND U9846 ( .A(n7351), .B(n7350), .Z(n7803) );
  XNOR U9847 ( .A(n7804), .B(n7803), .Z(n7802) );
  NANDN U9848 ( .A(n7357), .B(n7356), .Z(n7361) );
  NANDN U9849 ( .A(n7359), .B(n7358), .Z(n7360) );
  AND U9850 ( .A(n7361), .B(n7360), .Z(n7810) );
  NANDN U9851 ( .A(n7363), .B(n7362), .Z(n7367) );
  NANDN U9852 ( .A(n7365), .B(n7364), .Z(n7366) );
  AND U9853 ( .A(n7367), .B(n7366), .Z(n7809) );
  XOR U9854 ( .A(n7810), .B(n7809), .Z(n7808) );
  NAND U9855 ( .A(n7369), .B(n7368), .Z(n7373) );
  NAND U9856 ( .A(n7371), .B(n7370), .Z(n7372) );
  AND U9857 ( .A(n7373), .B(n7372), .Z(n7807) );
  XOR U9858 ( .A(n7808), .B(n7807), .Z(n7519) );
  NANDN U9859 ( .A(n7375), .B(n7374), .Z(n7379) );
  NANDN U9860 ( .A(n7377), .B(n7376), .Z(n7378) );
  AND U9861 ( .A(n7379), .B(n7378), .Z(n7793) );
  NANDN U9862 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U9863 ( .A(n7383), .B(n7382), .Z(n7384) );
  AND U9864 ( .A(n7385), .B(n7384), .Z(n7780) );
  NAND U9865 ( .A(n7387), .B(n7386), .Z(n7391) );
  NAND U9866 ( .A(n7389), .B(n7388), .Z(n7390) );
  AND U9867 ( .A(n7391), .B(n7390), .Z(n7525) );
  NAND U9868 ( .A(n7393), .B(n7392), .Z(n7397) );
  NAND U9869 ( .A(n7395), .B(n7394), .Z(n7396) );
  AND U9870 ( .A(n7397), .B(n7396), .Z(n7536) );
  AND U9871 ( .A(x[486]), .B(y[7736]), .Z(n7661) );
  AND U9872 ( .A(x[485]), .B(y[7737]), .Z(n7663) );
  AND U9873 ( .A(x[499]), .B(y[7723]), .Z(n7662) );
  XOR U9874 ( .A(n7663), .B(n7662), .Z(n7660) );
  XNOR U9875 ( .A(n7661), .B(n7660), .Z(n7540) );
  AND U9876 ( .A(x[484]), .B(y[7738]), .Z(n7701) );
  AND U9877 ( .A(x[483]), .B(y[7739]), .Z(n7703) );
  AND U9878 ( .A(x[498]), .B(y[7724]), .Z(n7702) );
  XOR U9879 ( .A(n7703), .B(n7702), .Z(n7700) );
  XOR U9880 ( .A(n7701), .B(n7700), .Z(n7543) );
  NAND U9881 ( .A(n7399), .B(n7398), .Z(n7403) );
  NAND U9882 ( .A(n7401), .B(n7400), .Z(n7402) );
  AND U9883 ( .A(n7403), .B(n7402), .Z(n7542) );
  XOR U9884 ( .A(n7540), .B(n7541), .Z(n7537) );
  XNOR U9885 ( .A(n7536), .B(n7537), .Z(n7535) );
  NAND U9886 ( .A(n7405), .B(n7404), .Z(n7409) );
  NAND U9887 ( .A(n7407), .B(n7406), .Z(n7408) );
  AND U9888 ( .A(n7409), .B(n7408), .Z(n7534) );
  XOR U9889 ( .A(n7535), .B(n7534), .Z(n7524) );
  XOR U9890 ( .A(n7525), .B(n7524), .Z(n7523) );
  NAND U9891 ( .A(n7411), .B(n7410), .Z(n7415) );
  NAND U9892 ( .A(n7413), .B(n7412), .Z(n7414) );
  AND U9893 ( .A(n7415), .B(n7414), .Z(n7522) );
  XOR U9894 ( .A(n7523), .B(n7522), .Z(n7783) );
  NAND U9895 ( .A(n7416), .B(n7653), .Z(n7420) );
  NAND U9896 ( .A(n7418), .B(n7417), .Z(n7419) );
  NAND U9897 ( .A(n7420), .B(n7419), .Z(n7531) );
  NAND U9898 ( .A(n7422), .B(n7421), .Z(n7426) );
  NAND U9899 ( .A(n7424), .B(n7423), .Z(n7425) );
  AND U9900 ( .A(n7426), .B(n7425), .Z(n7723) );
  AND U9901 ( .A(x[480]), .B(y[7742]), .Z(n7625) );
  AND U9902 ( .A(x[509]), .B(y[7713]), .Z(n7604) );
  XOR U9903 ( .A(o[62]), .B(n7604), .Z(n7627) );
  AND U9904 ( .A(x[510]), .B(y[7712]), .Z(n7626) );
  XOR U9905 ( .A(n7627), .B(n7626), .Z(n7624) );
  XOR U9906 ( .A(n7625), .B(n7624), .Z(n7725) );
  AND U9907 ( .A(x[500]), .B(y[7722]), .Z(n7575) );
  XOR U9908 ( .A(n7575), .B(n7574), .Z(n7573) );
  AND U9909 ( .A(x[488]), .B(y[7734]), .Z(n7572) );
  XNOR U9910 ( .A(n7573), .B(n7572), .Z(n7724) );
  XNOR U9911 ( .A(n7723), .B(n7722), .Z(n7530) );
  XOR U9912 ( .A(n7531), .B(n7530), .Z(n7528) );
  AND U9913 ( .A(x[487]), .B(y[7735]), .Z(n7687) );
  NAND U9914 ( .A(n7427), .B(n7687), .Z(n7431) );
  NAND U9915 ( .A(n7429), .B(n7428), .Z(n7430) );
  AND U9916 ( .A(n7431), .B(n7430), .Z(n7716) );
  AND U9917 ( .A(y[7721]), .B(x[501]), .Z(n7433) );
  AND U9918 ( .A(y[7720]), .B(x[502]), .Z(n7432) );
  XOR U9919 ( .A(n7433), .B(n7432), .Z(n7686) );
  XOR U9920 ( .A(n7687), .B(n7686), .Z(n7719) );
  AND U9921 ( .A(x[497]), .B(y[7725]), .Z(n7695) );
  AND U9922 ( .A(x[482]), .B(y[7740]), .Z(n7697) );
  AND U9923 ( .A(x[506]), .B(y[7716]), .Z(n7696) );
  XOR U9924 ( .A(n7697), .B(n7696), .Z(n7694) );
  XNOR U9925 ( .A(n7695), .B(n7694), .Z(n7718) );
  XNOR U9926 ( .A(n7716), .B(n7717), .Z(n7529) );
  NAND U9927 ( .A(n7435), .B(n7434), .Z(n7439) );
  NAND U9928 ( .A(n7437), .B(n7436), .Z(n7438) );
  NAND U9929 ( .A(n7439), .B(n7438), .Z(n7764) );
  XOR U9930 ( .A(n7765), .B(n7764), .Z(n7763) );
  AND U9931 ( .A(n7441), .B(n7440), .Z(n7445) );
  NAND U9932 ( .A(n7443), .B(n7442), .Z(n7444) );
  NANDN U9933 ( .A(n7445), .B(n7444), .Z(n7560) );
  AND U9934 ( .A(n7683), .B(n7446), .Z(n7450) );
  NAND U9935 ( .A(n7448), .B(n7447), .Z(n7449) );
  NANDN U9936 ( .A(n7450), .B(n7449), .Z(n7563) );
  NANDN U9937 ( .A(n7689), .B(n7451), .Z(n7455) );
  NANDN U9938 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U9939 ( .A(n7455), .B(n7454), .Z(n7553) );
  AND U9940 ( .A(x[503]), .B(y[7719]), .Z(n7651) );
  AND U9941 ( .A(y[7718]), .B(x[504]), .Z(n7457) );
  AND U9942 ( .A(y[7717]), .B(x[505]), .Z(n7456) );
  XOR U9943 ( .A(n7457), .B(n7456), .Z(n7650) );
  XOR U9944 ( .A(n7651), .B(n7650), .Z(n7555) );
  AND U9945 ( .A(n7458), .B(o[61]), .Z(n7645) );
  AND U9946 ( .A(x[508]), .B(y[7714]), .Z(n7647) );
  AND U9947 ( .A(x[496]), .B(y[7726]), .Z(n7646) );
  XOR U9948 ( .A(n7647), .B(n7646), .Z(n7644) );
  XNOR U9949 ( .A(n7645), .B(n7644), .Z(n7554) );
  XNOR U9950 ( .A(n7553), .B(n7552), .Z(n7562) );
  XOR U9951 ( .A(n7563), .B(n7562), .Z(n7561) );
  XOR U9952 ( .A(n7560), .B(n7561), .Z(n7762) );
  XOR U9953 ( .A(n7763), .B(n7762), .Z(n7782) );
  XNOR U9954 ( .A(n7780), .B(n7781), .Z(n7795) );
  NANDN U9955 ( .A(n7460), .B(n7459), .Z(n7464) );
  NANDN U9956 ( .A(n7462), .B(n7461), .Z(n7463) );
  AND U9957 ( .A(n7464), .B(n7463), .Z(n7794) );
  NANDN U9958 ( .A(n7466), .B(n7465), .Z(n7470) );
  NANDN U9959 ( .A(n7468), .B(n7467), .Z(n7469) );
  NAND U9960 ( .A(n7470), .B(n7469), .Z(n7776) );
  NANDN U9961 ( .A(n7472), .B(n7471), .Z(n7476) );
  NAND U9962 ( .A(n7474), .B(n7473), .Z(n7475) );
  AND U9963 ( .A(n7476), .B(n7475), .Z(n7757) );
  NAND U9964 ( .A(n7478), .B(n7477), .Z(n7482) );
  NAND U9965 ( .A(n7480), .B(n7479), .Z(n7481) );
  AND U9966 ( .A(n7482), .B(n7481), .Z(n7747) );
  NAND U9967 ( .A(n7484), .B(n7483), .Z(n7488) );
  NANDN U9968 ( .A(n7486), .B(n7485), .Z(n7487) );
  AND U9969 ( .A(n7488), .B(n7487), .Z(n7746) );
  XOR U9970 ( .A(n7747), .B(n7746), .Z(n7745) );
  NANDN U9971 ( .A(n7490), .B(n7489), .Z(n7494) );
  NANDN U9972 ( .A(n7492), .B(n7491), .Z(n7493) );
  NAND U9973 ( .A(n7494), .B(n7493), .Z(n7744) );
  XOR U9974 ( .A(n7745), .B(n7744), .Z(n7759) );
  NAND U9975 ( .A(n7621), .B(n7495), .Z(n7499) );
  NAND U9976 ( .A(n7497), .B(n7496), .Z(n7498) );
  AND U9977 ( .A(n7499), .B(n7498), .Z(n7740) );
  NAND U9978 ( .A(n7501), .B(n7500), .Z(n7505) );
  NAND U9979 ( .A(n7503), .B(n7502), .Z(n7504) );
  NAND U9980 ( .A(n7505), .B(n7504), .Z(n7546) );
  NAND U9981 ( .A(y[7730]), .B(x[492]), .Z(n7506) );
  XNOR U9982 ( .A(n7507), .B(n7506), .Z(n7681) );
  XOR U9983 ( .A(n7681), .B(n7680), .Z(n7619) );
  AND U9984 ( .A(y[7733]), .B(x[489]), .Z(n7509) );
  XOR U9985 ( .A(n7509), .B(n7508), .Z(n7618) );
  XOR U9986 ( .A(n7619), .B(n7618), .Z(n7549) );
  AND U9987 ( .A(x[507]), .B(y[7715]), .Z(n7569) );
  AND U9988 ( .A(x[481]), .B(y[7741]), .Z(n7568) );
  XOR U9989 ( .A(n7569), .B(n7568), .Z(n7567) );
  XOR U9990 ( .A(n7567), .B(n7566), .Z(n7548) );
  XOR U9991 ( .A(n7549), .B(n7548), .Z(n7547) );
  XOR U9992 ( .A(n7546), .B(n7547), .Z(n7741) );
  NAND U9993 ( .A(n7511), .B(n7510), .Z(n7515) );
  NANDN U9994 ( .A(n7513), .B(n7512), .Z(n7514) );
  AND U9995 ( .A(n7515), .B(n7514), .Z(n7738) );
  XNOR U9996 ( .A(n7739), .B(n7738), .Z(n7758) );
  XOR U9997 ( .A(n7757), .B(n7756), .Z(n7777) );
  XNOR U9998 ( .A(n7776), .B(n7777), .Z(n7775) );
  XOR U9999 ( .A(n7517), .B(n7516), .Z(n7801) );
  XNOR U10000 ( .A(n7802), .B(n7801), .Z(N127) );
  NANDN U10001 ( .A(n7517), .B(n7516), .Z(n7521) );
  NANDN U10002 ( .A(n7519), .B(n7518), .Z(n7520) );
  AND U10003 ( .A(n7521), .B(n7520), .Z(n7818) );
  NAND U10004 ( .A(n7523), .B(n7522), .Z(n7527) );
  NAND U10005 ( .A(n7525), .B(n7524), .Z(n7526) );
  AND U10006 ( .A(n7527), .B(n7526), .Z(n7791) );
  NANDN U10007 ( .A(n7529), .B(n7528), .Z(n7533) );
  NAND U10008 ( .A(n7531), .B(n7530), .Z(n7532) );
  AND U10009 ( .A(n7533), .B(n7532), .Z(n7773) );
  NAND U10010 ( .A(n7535), .B(n7534), .Z(n7539) );
  NANDN U10011 ( .A(n7537), .B(n7536), .Z(n7538) );
  AND U10012 ( .A(n7539), .B(n7538), .Z(n7755) );
  NANDN U10013 ( .A(n7541), .B(n7540), .Z(n7545) );
  NANDN U10014 ( .A(n7543), .B(n7542), .Z(n7544) );
  AND U10015 ( .A(n7545), .B(n7544), .Z(n7737) );
  NAND U10016 ( .A(n7547), .B(n7546), .Z(n7551) );
  NAND U10017 ( .A(n7549), .B(n7548), .Z(n7550) );
  AND U10018 ( .A(n7551), .B(n7550), .Z(n7559) );
  NAND U10019 ( .A(n7553), .B(n7552), .Z(n7557) );
  NANDN U10020 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U10021 ( .A(n7557), .B(n7556), .Z(n7558) );
  XNOR U10022 ( .A(n7559), .B(n7558), .Z(n7735) );
  NAND U10023 ( .A(n7561), .B(n7560), .Z(n7565) );
  NAND U10024 ( .A(n7563), .B(n7562), .Z(n7564) );
  AND U10025 ( .A(n7565), .B(n7564), .Z(n7733) );
  NAND U10026 ( .A(n7567), .B(n7566), .Z(n7571) );
  NAND U10027 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U10028 ( .A(n7571), .B(n7570), .Z(n7579) );
  NAND U10029 ( .A(n7573), .B(n7572), .Z(n7577) );
  NAND U10030 ( .A(n7575), .B(n7574), .Z(n7576) );
  NAND U10031 ( .A(n7577), .B(n7576), .Z(n7578) );
  XNOR U10032 ( .A(n7579), .B(n7578), .Z(n7643) );
  AND U10033 ( .A(y[7741]), .B(x[482]), .Z(n7581) );
  NAND U10034 ( .A(y[7726]), .B(x[497]), .Z(n7580) );
  XNOR U10035 ( .A(n7581), .B(n7580), .Z(n7585) );
  AND U10036 ( .A(y[7740]), .B(x[483]), .Z(n7583) );
  NAND U10037 ( .A(y[7725]), .B(x[498]), .Z(n7582) );
  XNOR U10038 ( .A(n7583), .B(n7582), .Z(n7584) );
  XOR U10039 ( .A(n7585), .B(n7584), .Z(n7587) );
  AND U10040 ( .A(x[490]), .B(y[7733]), .Z(n7620) );
  XNOR U10041 ( .A(n7682), .B(n7620), .Z(n7586) );
  XNOR U10042 ( .A(n7587), .B(n7586), .Z(n7603) );
  AND U10043 ( .A(y[7737]), .B(x[486]), .Z(n7589) );
  NAND U10044 ( .A(y[7720]), .B(x[503]), .Z(n7588) );
  XNOR U10045 ( .A(n7589), .B(n7588), .Z(n7593) );
  AND U10046 ( .A(y[7716]), .B(x[507]), .Z(n7591) );
  NAND U10047 ( .A(y[7724]), .B(x[499]), .Z(n7590) );
  XNOR U10048 ( .A(n7591), .B(n7590), .Z(n7592) );
  XOR U10049 ( .A(n7593), .B(n7592), .Z(n7601) );
  AND U10050 ( .A(y[7712]), .B(x[511]), .Z(n7595) );
  NAND U10051 ( .A(y[7739]), .B(x[484]), .Z(n7594) );
  XNOR U10052 ( .A(n7595), .B(n7594), .Z(n7599) );
  AND U10053 ( .A(y[7738]), .B(x[485]), .Z(n7597) );
  NAND U10054 ( .A(y[7736]), .B(x[487]), .Z(n7596) );
  XNOR U10055 ( .A(n7597), .B(n7596), .Z(n7598) );
  XNOR U10056 ( .A(n7599), .B(n7598), .Z(n7600) );
  XNOR U10057 ( .A(n7601), .B(n7600), .Z(n7602) );
  XOR U10058 ( .A(n7603), .B(n7602), .Z(n7617) );
  AND U10059 ( .A(y[7713]), .B(x[510]), .Z(n7611) );
  AND U10060 ( .A(n7604), .B(o[62]), .Z(n7609) );
  AND U10061 ( .A(x[505]), .B(y[7718]), .Z(n7652) );
  XOR U10062 ( .A(n7652), .B(o[63]), .Z(n7607) );
  AND U10063 ( .A(x[502]), .B(y[7721]), .Z(n7688) );
  XNOR U10064 ( .A(n7605), .B(n7688), .Z(n7606) );
  XNOR U10065 ( .A(n7607), .B(n7606), .Z(n7608) );
  XNOR U10066 ( .A(n7609), .B(n7608), .Z(n7610) );
  XNOR U10067 ( .A(n7611), .B(n7610), .Z(n7615) );
  AND U10068 ( .A(y[7722]), .B(x[501]), .Z(n7613) );
  NAND U10069 ( .A(y[7735]), .B(x[488]), .Z(n7612) );
  XNOR U10070 ( .A(n7613), .B(n7612), .Z(n7614) );
  XNOR U10071 ( .A(n7615), .B(n7614), .Z(n7616) );
  XNOR U10072 ( .A(n7617), .B(n7616), .Z(n7633) );
  NAND U10073 ( .A(n7619), .B(n7618), .Z(n7623) );
  NAND U10074 ( .A(n7621), .B(n7620), .Z(n7622) );
  AND U10075 ( .A(n7623), .B(n7622), .Z(n7631) );
  NAND U10076 ( .A(n7625), .B(n7624), .Z(n7629) );
  NAND U10077 ( .A(n7627), .B(n7626), .Z(n7628) );
  NAND U10078 ( .A(n7629), .B(n7628), .Z(n7630) );
  XNOR U10079 ( .A(n7631), .B(n7630), .Z(n7632) );
  XOR U10080 ( .A(n7633), .B(n7632), .Z(n7641) );
  AND U10081 ( .A(y[7714]), .B(x[509]), .Z(n7635) );
  NAND U10082 ( .A(y[7723]), .B(x[500]), .Z(n7634) );
  XNOR U10083 ( .A(n7635), .B(n7634), .Z(n7639) );
  AND U10084 ( .A(y[7727]), .B(x[496]), .Z(n7637) );
  NAND U10085 ( .A(y[7743]), .B(x[480]), .Z(n7636) );
  XNOR U10086 ( .A(n7637), .B(n7636), .Z(n7638) );
  XNOR U10087 ( .A(n7639), .B(n7638), .Z(n7640) );
  XNOR U10088 ( .A(n7641), .B(n7640), .Z(n7642) );
  XOR U10089 ( .A(n7643), .B(n7642), .Z(n7715) );
  NAND U10090 ( .A(n7645), .B(n7644), .Z(n7649) );
  NAND U10091 ( .A(n7647), .B(n7646), .Z(n7648) );
  AND U10092 ( .A(n7649), .B(n7648), .Z(n7657) );
  NAND U10093 ( .A(n7651), .B(n7650), .Z(n7655) );
  NAND U10094 ( .A(n7653), .B(n7652), .Z(n7654) );
  NAND U10095 ( .A(n7655), .B(n7654), .Z(n7656) );
  XNOR U10096 ( .A(n7657), .B(n7656), .Z(n7713) );
  AND U10097 ( .A(y[7742]), .B(x[481]), .Z(n7659) );
  NAND U10098 ( .A(y[7715]), .B(x[508]), .Z(n7658) );
  XNOR U10099 ( .A(n7659), .B(n7658), .Z(n7679) );
  AND U10100 ( .A(y[7734]), .B(x[489]), .Z(n7677) );
  NAND U10101 ( .A(n7661), .B(n7660), .Z(n7665) );
  NAND U10102 ( .A(n7663), .B(n7662), .Z(n7664) );
  AND U10103 ( .A(n7665), .B(n7664), .Z(n7673) );
  AND U10104 ( .A(y[7729]), .B(x[494]), .Z(n7667) );
  NAND U10105 ( .A(y[7717]), .B(x[506]), .Z(n7666) );
  XNOR U10106 ( .A(n7667), .B(n7666), .Z(n7671) );
  AND U10107 ( .A(y[7732]), .B(x[491]), .Z(n7669) );
  NAND U10108 ( .A(y[7731]), .B(x[492]), .Z(n7668) );
  XNOR U10109 ( .A(n7669), .B(n7668), .Z(n7670) );
  XNOR U10110 ( .A(n7671), .B(n7670), .Z(n7672) );
  XNOR U10111 ( .A(n7673), .B(n7672), .Z(n7674) );
  XNOR U10112 ( .A(n7675), .B(n7674), .Z(n7676) );
  XNOR U10113 ( .A(n7677), .B(n7676), .Z(n7678) );
  XOR U10114 ( .A(n7679), .B(n7678), .Z(n7711) );
  NAND U10115 ( .A(n7681), .B(n7680), .Z(n7685) );
  NAND U10116 ( .A(n7683), .B(n7682), .Z(n7684) );
  AND U10117 ( .A(n7685), .B(n7684), .Z(n7693) );
  NAND U10118 ( .A(n7687), .B(n7686), .Z(n7691) );
  NANDN U10119 ( .A(n7689), .B(n7688), .Z(n7690) );
  NAND U10120 ( .A(n7691), .B(n7690), .Z(n7692) );
  XNOR U10121 ( .A(n7693), .B(n7692), .Z(n7709) );
  NAND U10122 ( .A(n7695), .B(n7694), .Z(n7699) );
  NAND U10123 ( .A(n7697), .B(n7696), .Z(n7698) );
  AND U10124 ( .A(n7699), .B(n7698), .Z(n7707) );
  NAND U10125 ( .A(n7701), .B(n7700), .Z(n7705) );
  NAND U10126 ( .A(n7703), .B(n7702), .Z(n7704) );
  NAND U10127 ( .A(n7705), .B(n7704), .Z(n7706) );
  XNOR U10128 ( .A(n7707), .B(n7706), .Z(n7708) );
  XNOR U10129 ( .A(n7709), .B(n7708), .Z(n7710) );
  XNOR U10130 ( .A(n7711), .B(n7710), .Z(n7712) );
  XNOR U10131 ( .A(n7713), .B(n7712), .Z(n7714) );
  XNOR U10132 ( .A(n7715), .B(n7714), .Z(n7731) );
  NANDN U10133 ( .A(n7717), .B(n7716), .Z(n7721) );
  NANDN U10134 ( .A(n7719), .B(n7718), .Z(n7720) );
  AND U10135 ( .A(n7721), .B(n7720), .Z(n7729) );
  NAND U10136 ( .A(n7723), .B(n7722), .Z(n7727) );
  NANDN U10137 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U10138 ( .A(n7727), .B(n7726), .Z(n7728) );
  XNOR U10139 ( .A(n7729), .B(n7728), .Z(n7730) );
  XNOR U10140 ( .A(n7731), .B(n7730), .Z(n7732) );
  XNOR U10141 ( .A(n7733), .B(n7732), .Z(n7734) );
  XNOR U10142 ( .A(n7735), .B(n7734), .Z(n7736) );
  XNOR U10143 ( .A(n7737), .B(n7736), .Z(n7753) );
  NAND U10144 ( .A(n7739), .B(n7738), .Z(n7743) );
  NANDN U10145 ( .A(n7741), .B(n7740), .Z(n7742) );
  AND U10146 ( .A(n7743), .B(n7742), .Z(n7751) );
  NAND U10147 ( .A(n7745), .B(n7744), .Z(n7749) );
  NAND U10148 ( .A(n7747), .B(n7746), .Z(n7748) );
  NAND U10149 ( .A(n7749), .B(n7748), .Z(n7750) );
  XNOR U10150 ( .A(n7751), .B(n7750), .Z(n7752) );
  XNOR U10151 ( .A(n7753), .B(n7752), .Z(n7754) );
  XNOR U10152 ( .A(n7755), .B(n7754), .Z(n7771) );
  NAND U10153 ( .A(n7757), .B(n7756), .Z(n7761) );
  NANDN U10154 ( .A(n7759), .B(n7758), .Z(n7760) );
  AND U10155 ( .A(n7761), .B(n7760), .Z(n7769) );
  NAND U10156 ( .A(n7763), .B(n7762), .Z(n7767) );
  NAND U10157 ( .A(n7765), .B(n7764), .Z(n7766) );
  NAND U10158 ( .A(n7767), .B(n7766), .Z(n7768) );
  XNOR U10159 ( .A(n7769), .B(n7768), .Z(n7770) );
  XNOR U10160 ( .A(n7771), .B(n7770), .Z(n7772) );
  XNOR U10161 ( .A(n7773), .B(n7772), .Z(n7789) );
  NANDN U10162 ( .A(n7775), .B(n7774), .Z(n7779) );
  NAND U10163 ( .A(n7777), .B(n7776), .Z(n7778) );
  AND U10164 ( .A(n7779), .B(n7778), .Z(n7787) );
  NANDN U10165 ( .A(n7781), .B(n7780), .Z(n7785) );
  NANDN U10166 ( .A(n7783), .B(n7782), .Z(n7784) );
  NAND U10167 ( .A(n7785), .B(n7784), .Z(n7786) );
  XNOR U10168 ( .A(n7787), .B(n7786), .Z(n7788) );
  XNOR U10169 ( .A(n7789), .B(n7788), .Z(n7790) );
  XNOR U10170 ( .A(n7791), .B(n7790), .Z(n7800) );
  IV U10171 ( .A(n7793), .Z(n7792) );
  OR U10172 ( .A(n7794), .B(n7792), .Z(n7798) );
  ANDN U10173 ( .B(n7794), .A(n7793), .Z(n7796) );
  NANDN U10174 ( .A(n7796), .B(n7795), .Z(n7797) );
  NAND U10175 ( .A(n7798), .B(n7797), .Z(n7799) );
  XNOR U10176 ( .A(n7800), .B(n7799), .Z(n7816) );
  NAND U10177 ( .A(n7802), .B(n7801), .Z(n7806) );
  NANDN U10178 ( .A(n7804), .B(n7803), .Z(n7805) );
  AND U10179 ( .A(n7806), .B(n7805), .Z(n7814) );
  NAND U10180 ( .A(n7808), .B(n7807), .Z(n7812) );
  NAND U10181 ( .A(n7810), .B(n7809), .Z(n7811) );
  NAND U10182 ( .A(n7812), .B(n7811), .Z(n7813) );
  XNOR U10183 ( .A(n7814), .B(n7813), .Z(n7815) );
  XNOR U10184 ( .A(n7816), .B(n7815), .Z(n7817) );
  XNOR U10185 ( .A(n7818), .B(n7817), .Z(N128) );
  AND U10186 ( .A(x[480]), .B(y[7744]), .Z(n8465) );
  XOR U10187 ( .A(n8465), .B(o[64]), .Z(N161) );
  AND U10188 ( .A(x[481]), .B(y[7744]), .Z(n7827) );
  AND U10189 ( .A(x[480]), .B(y[7745]), .Z(n7826) );
  XNOR U10190 ( .A(n7826), .B(o[65]), .Z(n7819) );
  XNOR U10191 ( .A(n7827), .B(n7819), .Z(n7821) );
  NAND U10192 ( .A(n8465), .B(o[64]), .Z(n7820) );
  XNOR U10193 ( .A(n7821), .B(n7820), .Z(N162) );
  NANDN U10194 ( .A(n7827), .B(n7819), .Z(n7823) );
  NAND U10195 ( .A(n7821), .B(n7820), .Z(n7822) );
  AND U10196 ( .A(n7823), .B(n7822), .Z(n7833) );
  AND U10197 ( .A(x[480]), .B(y[7746]), .Z(n7840) );
  XNOR U10198 ( .A(n7840), .B(o[66]), .Z(n7832) );
  XNOR U10199 ( .A(n7833), .B(n7832), .Z(n7835) );
  AND U10200 ( .A(y[7744]), .B(x[482]), .Z(n7825) );
  NAND U10201 ( .A(y[7745]), .B(x[481]), .Z(n7824) );
  XNOR U10202 ( .A(n7825), .B(n7824), .Z(n7829) );
  AND U10203 ( .A(n7826), .B(o[65]), .Z(n7828) );
  XNOR U10204 ( .A(n7829), .B(n7828), .Z(n7834) );
  XNOR U10205 ( .A(n7835), .B(n7834), .Z(N163) );
  AND U10206 ( .A(x[482]), .B(y[7745]), .Z(n7847) );
  NAND U10207 ( .A(n7847), .B(n7827), .Z(n7831) );
  NAND U10208 ( .A(n7829), .B(n7828), .Z(n7830) );
  AND U10209 ( .A(n7831), .B(n7830), .Z(n7850) );
  NANDN U10210 ( .A(n7833), .B(n7832), .Z(n7837) );
  NAND U10211 ( .A(n7835), .B(n7834), .Z(n7836) );
  AND U10212 ( .A(n7837), .B(n7836), .Z(n7849) );
  XNOR U10213 ( .A(n7850), .B(n7849), .Z(n7852) );
  AND U10214 ( .A(x[481]), .B(y[7746]), .Z(n7956) );
  XOR U10215 ( .A(n7847), .B(o[67]), .Z(n7855) );
  XOR U10216 ( .A(n7956), .B(n7855), .Z(n7857) );
  AND U10217 ( .A(y[7744]), .B(x[483]), .Z(n7839) );
  NAND U10218 ( .A(y[7747]), .B(x[480]), .Z(n7838) );
  XNOR U10219 ( .A(n7839), .B(n7838), .Z(n7842) );
  AND U10220 ( .A(n7840), .B(o[66]), .Z(n7841) );
  XOR U10221 ( .A(n7842), .B(n7841), .Z(n7856) );
  XOR U10222 ( .A(n7857), .B(n7856), .Z(n7851) );
  XOR U10223 ( .A(n7852), .B(n7851), .Z(N164) );
  AND U10224 ( .A(x[483]), .B(y[7747]), .Z(n7900) );
  NAND U10225 ( .A(n8465), .B(n7900), .Z(n7844) );
  NAND U10226 ( .A(n7842), .B(n7841), .Z(n7843) );
  NAND U10227 ( .A(n7844), .B(n7843), .Z(n7878) );
  AND U10228 ( .A(y[7748]), .B(x[480]), .Z(n7846) );
  NAND U10229 ( .A(y[7744]), .B(x[484]), .Z(n7845) );
  XNOR U10230 ( .A(n7846), .B(n7845), .Z(n7871) );
  NAND U10231 ( .A(n7847), .B(o[67]), .Z(n7872) );
  AND U10232 ( .A(x[482]), .B(y[7746]), .Z(n8015) );
  NAND U10233 ( .A(y[7747]), .B(x[481]), .Z(n7848) );
  XNOR U10234 ( .A(n8015), .B(n7848), .Z(n7868) );
  AND U10235 ( .A(x[483]), .B(y[7745]), .Z(n7865) );
  XOR U10236 ( .A(o[68]), .B(n7865), .Z(n7867) );
  XOR U10237 ( .A(n7868), .B(n7867), .Z(n7875) );
  XOR U10238 ( .A(n7876), .B(n7875), .Z(n7877) );
  XOR U10239 ( .A(n7878), .B(n7877), .Z(n7882) );
  NANDN U10240 ( .A(n7850), .B(n7849), .Z(n7854) );
  NAND U10241 ( .A(n7852), .B(n7851), .Z(n7853) );
  NAND U10242 ( .A(n7854), .B(n7853), .Z(n7883) );
  NAND U10243 ( .A(n7956), .B(n7855), .Z(n7859) );
  NAND U10244 ( .A(n7857), .B(n7856), .Z(n7858) );
  NAND U10245 ( .A(n7859), .B(n7858), .Z(n7884) );
  IV U10246 ( .A(n7884), .Z(n7881) );
  XOR U10247 ( .A(n7883), .B(n7881), .Z(n7860) );
  XNOR U10248 ( .A(n7882), .B(n7860), .Z(N165) );
  AND U10249 ( .A(y[7746]), .B(x[483]), .Z(n7862) );
  NAND U10250 ( .A(y[7748]), .B(x[481]), .Z(n7861) );
  XNOR U10251 ( .A(n7862), .B(n7861), .Z(n7887) );
  AND U10252 ( .A(x[484]), .B(y[7745]), .Z(n7898) );
  XOR U10253 ( .A(n7898), .B(o[69]), .Z(n7886) );
  XNOR U10254 ( .A(n7887), .B(n7886), .Z(n7890) );
  NAND U10255 ( .A(x[482]), .B(y[7747]), .Z(n7964) );
  AND U10256 ( .A(y[7744]), .B(x[485]), .Z(n7864) );
  NAND U10257 ( .A(y[7749]), .B(x[480]), .Z(n7863) );
  XNOR U10258 ( .A(n7864), .B(n7863), .Z(n7893) );
  AND U10259 ( .A(o[68]), .B(n7865), .Z(n7892) );
  XOR U10260 ( .A(n7893), .B(n7892), .Z(n7891) );
  XOR U10261 ( .A(n7964), .B(n7891), .Z(n7866) );
  XOR U10262 ( .A(n7890), .B(n7866), .Z(n7908) );
  NANDN U10263 ( .A(n7964), .B(n7956), .Z(n7870) );
  NAND U10264 ( .A(n7868), .B(n7867), .Z(n7869) );
  AND U10265 ( .A(n7870), .B(n7869), .Z(n7906) );
  AND U10266 ( .A(x[484]), .B(y[7748]), .Z(n8671) );
  NAND U10267 ( .A(n8671), .B(n8465), .Z(n7874) );
  NANDN U10268 ( .A(n7872), .B(n7871), .Z(n7873) );
  NAND U10269 ( .A(n7874), .B(n7873), .Z(n7905) );
  XNOR U10270 ( .A(n7908), .B(n7907), .Z(n7904) );
  NAND U10271 ( .A(n7876), .B(n7875), .Z(n7880) );
  NAND U10272 ( .A(n7878), .B(n7877), .Z(n7879) );
  NAND U10273 ( .A(n7880), .B(n7879), .Z(n7903) );
  XOR U10274 ( .A(n7903), .B(n7902), .Z(n7885) );
  XNOR U10275 ( .A(n7904), .B(n7885), .Z(N166) );
  AND U10276 ( .A(x[483]), .B(y[7748]), .Z(n7965) );
  NAND U10277 ( .A(n7965), .B(n7956), .Z(n7889) );
  NAND U10278 ( .A(n7887), .B(n7886), .Z(n7888) );
  NAND U10279 ( .A(n7889), .B(n7888), .Z(n7944) );
  XOR U10280 ( .A(n7944), .B(n7943), .Z(n7946) );
  AND U10281 ( .A(x[485]), .B(y[7749]), .Z(n8142) );
  NAND U10282 ( .A(n8465), .B(n8142), .Z(n7895) );
  NAND U10283 ( .A(n7893), .B(n7892), .Z(n7894) );
  AND U10284 ( .A(n7895), .B(n7894), .Z(n7913) );
  AND U10285 ( .A(y[7744]), .B(x[486]), .Z(n7897) );
  NAND U10286 ( .A(y[7750]), .B(x[480]), .Z(n7896) );
  XNOR U10287 ( .A(n7897), .B(n7896), .Z(n7919) );
  NAND U10288 ( .A(n7898), .B(o[69]), .Z(n7920) );
  NAND U10289 ( .A(y[7748]), .B(x[482]), .Z(n7899) );
  XNOR U10290 ( .A(n7900), .B(n7899), .Z(n7924) );
  AND U10291 ( .A(x[481]), .B(y[7749]), .Z(n8172) );
  NAND U10292 ( .A(y[7746]), .B(x[484]), .Z(n7901) );
  XNOR U10293 ( .A(n8172), .B(n7901), .Z(n7928) );
  NAND U10294 ( .A(x[485]), .B(y[7745]), .Z(n7935) );
  XOR U10295 ( .A(n7928), .B(n7927), .Z(n7923) );
  XOR U10296 ( .A(n7924), .B(n7923), .Z(n7914) );
  XOR U10297 ( .A(n7915), .B(n7914), .Z(n7945) );
  XNOR U10298 ( .A(n7946), .B(n7945), .Z(n7939) );
  NANDN U10299 ( .A(n7906), .B(n7905), .Z(n7910) );
  NAND U10300 ( .A(n7908), .B(n7907), .Z(n7909) );
  NAND U10301 ( .A(n7910), .B(n7909), .Z(n7937) );
  IV U10302 ( .A(n7937), .Z(n7936) );
  XOR U10303 ( .A(n7938), .B(n7936), .Z(n7911) );
  XNOR U10304 ( .A(n7939), .B(n7911), .Z(N167) );
  NANDN U10305 ( .A(n7913), .B(n7912), .Z(n7917) );
  NAND U10306 ( .A(n7915), .B(n7914), .Z(n7916) );
  AND U10307 ( .A(n7917), .B(n7916), .Z(n7984) );
  AND U10308 ( .A(y[7746]), .B(x[485]), .Z(n8047) );
  NAND U10309 ( .A(y[7750]), .B(x[481]), .Z(n7918) );
  XNOR U10310 ( .A(n8047), .B(n7918), .Z(n7957) );
  NAND U10311 ( .A(x[486]), .B(y[7745]), .Z(n7962) );
  XOR U10312 ( .A(o[71]), .B(n7962), .Z(n7958) );
  AND U10313 ( .A(y[7750]), .B(x[486]), .Z(n8192) );
  NAND U10314 ( .A(n8465), .B(n8192), .Z(n7922) );
  NANDN U10315 ( .A(n7920), .B(n7919), .Z(n7921) );
  AND U10316 ( .A(n7922), .B(n7921), .Z(n7975) );
  NANDN U10317 ( .A(n7964), .B(n7965), .Z(n7926) );
  NAND U10318 ( .A(n7924), .B(n7923), .Z(n7925) );
  AND U10319 ( .A(n7926), .B(n7925), .Z(n7977) );
  XOR U10320 ( .A(n7978), .B(n7977), .Z(n7982) );
  AND U10321 ( .A(x[484]), .B(y[7749]), .Z(n8470) );
  NAND U10322 ( .A(n8470), .B(n7956), .Z(n7930) );
  NAND U10323 ( .A(n7928), .B(n7927), .Z(n7929) );
  AND U10324 ( .A(n7930), .B(n7929), .Z(n7953) );
  AND U10325 ( .A(y[7749]), .B(x[482]), .Z(n7932) );
  NAND U10326 ( .A(y[7747]), .B(x[484]), .Z(n7931) );
  XNOR U10327 ( .A(n7932), .B(n7931), .Z(n7966) );
  XOR U10328 ( .A(n7966), .B(n7965), .Z(n7951) );
  AND U10329 ( .A(y[7744]), .B(x[487]), .Z(n7934) );
  NAND U10330 ( .A(y[7751]), .B(x[480]), .Z(n7933) );
  XNOR U10331 ( .A(n7934), .B(n7933), .Z(n7970) );
  ANDN U10332 ( .B(o[70]), .A(n7935), .Z(n7969) );
  XNOR U10333 ( .A(n7970), .B(n7969), .Z(n7950) );
  XOR U10334 ( .A(n7953), .B(n7952), .Z(n7981) );
  XOR U10335 ( .A(n7982), .B(n7981), .Z(n7983) );
  XNOR U10336 ( .A(n7984), .B(n7983), .Z(n7990) );
  OR U10337 ( .A(n7938), .B(n7936), .Z(n7942) );
  ANDN U10338 ( .B(n7938), .A(n7937), .Z(n7940) );
  OR U10339 ( .A(n7940), .B(n7939), .Z(n7941) );
  AND U10340 ( .A(n7942), .B(n7941), .Z(n7988) );
  NAND U10341 ( .A(n7944), .B(n7943), .Z(n7948) );
  NAND U10342 ( .A(n7946), .B(n7945), .Z(n7947) );
  AND U10343 ( .A(n7948), .B(n7947), .Z(n7989) );
  IV U10344 ( .A(n7989), .Z(n7987) );
  XOR U10345 ( .A(n7988), .B(n7987), .Z(n7949) );
  XNOR U10346 ( .A(n7990), .B(n7949), .Z(N168) );
  NANDN U10347 ( .A(n7951), .B(n7950), .Z(n7955) );
  NAND U10348 ( .A(n7953), .B(n7952), .Z(n7954) );
  AND U10349 ( .A(n7955), .B(n7954), .Z(n8028) );
  AND U10350 ( .A(x[485]), .B(y[7750]), .Z(n8134) );
  NAND U10351 ( .A(n8134), .B(n7956), .Z(n7960) );
  NANDN U10352 ( .A(n7958), .B(n7957), .Z(n7959) );
  AND U10353 ( .A(n7960), .B(n7959), .Z(n8026) );
  AND U10354 ( .A(y[7747]), .B(x[485]), .Z(n8574) );
  NAND U10355 ( .A(y[7751]), .B(x[481]), .Z(n7961) );
  XNOR U10356 ( .A(n8574), .B(n7961), .Z(n8006) );
  ANDN U10357 ( .B(o[71]), .A(n7962), .Z(n8007) );
  XNOR U10358 ( .A(n8006), .B(n8007), .Z(n8011) );
  AND U10359 ( .A(x[483]), .B(y[7749]), .Z(n8811) );
  AND U10360 ( .A(x[486]), .B(y[7746]), .Z(n7963) );
  AND U10361 ( .A(y[7750]), .B(x[482]), .Z(n8905) );
  XOR U10362 ( .A(n7963), .B(n8905), .Z(n8016) );
  XNOR U10363 ( .A(n8671), .B(n8016), .Z(n8010) );
  XOR U10364 ( .A(n8811), .B(n8010), .Z(n8012) );
  XOR U10365 ( .A(n8011), .B(n8012), .Z(n8025) );
  XNOR U10366 ( .A(n8028), .B(n8027), .Z(n8036) );
  NANDN U10367 ( .A(n7964), .B(n8470), .Z(n7968) );
  NAND U10368 ( .A(n7966), .B(n7965), .Z(n7967) );
  AND U10369 ( .A(n7968), .B(n7967), .Z(n8022) );
  AND U10370 ( .A(x[487]), .B(y[7751]), .Z(n8340) );
  NAND U10371 ( .A(n8465), .B(n8340), .Z(n7972) );
  NAND U10372 ( .A(n7970), .B(n7969), .Z(n7971) );
  AND U10373 ( .A(n7972), .B(n7971), .Z(n8020) );
  AND U10374 ( .A(y[7744]), .B(x[488]), .Z(n7974) );
  NAND U10375 ( .A(y[7752]), .B(x[480]), .Z(n7973) );
  XNOR U10376 ( .A(n7974), .B(n7973), .Z(n7996) );
  NAND U10377 ( .A(x[487]), .B(y[7745]), .Z(n8002) );
  XOR U10378 ( .A(o[72]), .B(n8002), .Z(n7997) );
  XNOR U10379 ( .A(n7996), .B(n7997), .Z(n8019) );
  NANDN U10380 ( .A(n7976), .B(n7975), .Z(n7980) );
  NAND U10381 ( .A(n7978), .B(n7977), .Z(n7979) );
  NAND U10382 ( .A(n7980), .B(n7979), .Z(n8034) );
  XOR U10383 ( .A(n8036), .B(n8037), .Z(n8033) );
  NAND U10384 ( .A(n7982), .B(n7981), .Z(n7986) );
  NAND U10385 ( .A(n7984), .B(n7983), .Z(n7985) );
  NAND U10386 ( .A(n7986), .B(n7985), .Z(n8031) );
  NANDN U10387 ( .A(n7987), .B(n7988), .Z(n7993) );
  NOR U10388 ( .A(n7989), .B(n7988), .Z(n7991) );
  OR U10389 ( .A(n7991), .B(n7990), .Z(n7992) );
  AND U10390 ( .A(n7993), .B(n7992), .Z(n8032) );
  XOR U10391 ( .A(n8031), .B(n8032), .Z(n7994) );
  XNOR U10392 ( .A(n8033), .B(n7994), .Z(N169) );
  AND U10393 ( .A(x[488]), .B(y[7752]), .Z(n7995) );
  NAND U10394 ( .A(n7995), .B(n8465), .Z(n7999) );
  NANDN U10395 ( .A(n7997), .B(n7996), .Z(n7998) );
  AND U10396 ( .A(n7999), .B(n7998), .Z(n8074) );
  AND U10397 ( .A(y[7748]), .B(x[485]), .Z(n8001) );
  NAND U10398 ( .A(y[7746]), .B(x[487]), .Z(n8000) );
  XNOR U10399 ( .A(n8001), .B(n8000), .Z(n8049) );
  ANDN U10400 ( .B(o[72]), .A(n8002), .Z(n8048) );
  XOR U10401 ( .A(n8049), .B(n8048), .Z(n8072) );
  AND U10402 ( .A(y[7744]), .B(x[489]), .Z(n8004) );
  NAND U10403 ( .A(y[7753]), .B(x[480]), .Z(n8003) );
  XNOR U10404 ( .A(n8004), .B(n8003), .Z(n8056) );
  NAND U10405 ( .A(x[488]), .B(y[7745]), .Z(n8063) );
  XNOR U10406 ( .A(o[73]), .B(n8063), .Z(n8055) );
  XNOR U10407 ( .A(n8056), .B(n8055), .Z(n8071) );
  XNOR U10408 ( .A(n8072), .B(n8071), .Z(n8073) );
  XOR U10409 ( .A(n8074), .B(n8073), .Z(n8070) );
  AND U10410 ( .A(y[7747]), .B(x[486]), .Z(n8409) );
  NAND U10411 ( .A(y[7752]), .B(x[481]), .Z(n8005) );
  XNOR U10412 ( .A(n8409), .B(n8005), .Z(n8060) );
  XOR U10413 ( .A(n8470), .B(n8060), .Z(n8078) );
  NAND U10414 ( .A(x[482]), .B(y[7751]), .Z(n8718) );
  AND U10415 ( .A(x[483]), .B(y[7750]), .Z(n8419) );
  XNOR U10416 ( .A(n8718), .B(n8419), .Z(n8077) );
  XOR U10417 ( .A(n8078), .B(n8077), .Z(n8067) );
  NAND U10418 ( .A(x[485]), .B(y[7751]), .Z(n8246) );
  AND U10419 ( .A(x[481]), .B(y[7747]), .Z(n8059) );
  NANDN U10420 ( .A(n8246), .B(n8059), .Z(n8009) );
  NAND U10421 ( .A(n8007), .B(n8006), .Z(n8008) );
  NAND U10422 ( .A(n8009), .B(n8008), .Z(n8068) );
  XOR U10423 ( .A(n8067), .B(n8068), .Z(n8069) );
  XOR U10424 ( .A(n8070), .B(n8069), .Z(n8043) );
  NANDN U10425 ( .A(n8811), .B(n8010), .Z(n8014) );
  NANDN U10426 ( .A(n8012), .B(n8011), .Z(n8013) );
  NAND U10427 ( .A(n8014), .B(n8013), .Z(n8041) );
  NAND U10428 ( .A(n8192), .B(n8015), .Z(n8018) );
  NAND U10429 ( .A(n8671), .B(n8016), .Z(n8017) );
  AND U10430 ( .A(n8018), .B(n8017), .Z(n8042) );
  XNOR U10431 ( .A(n8041), .B(n8042), .Z(n8044) );
  NANDN U10432 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U10433 ( .A(n8022), .B(n8021), .Z(n8023) );
  AND U10434 ( .A(n8024), .B(n8023), .Z(n8082) );
  NANDN U10435 ( .A(n8026), .B(n8025), .Z(n8030) );
  NAND U10436 ( .A(n8028), .B(n8027), .Z(n8029) );
  NAND U10437 ( .A(n8030), .B(n8029), .Z(n8081) );
  XNOR U10438 ( .A(n8083), .B(n8084), .Z(n8089) );
  NANDN U10439 ( .A(n8035), .B(n8034), .Z(n8039) );
  NANDN U10440 ( .A(n8037), .B(n8036), .Z(n8038) );
  AND U10441 ( .A(n8039), .B(n8038), .Z(n8087) );
  XOR U10442 ( .A(n8088), .B(n8087), .Z(n8040) );
  XNOR U10443 ( .A(n8089), .B(n8040), .Z(N170) );
  NAND U10444 ( .A(n8042), .B(n8041), .Z(n8046) );
  NANDN U10445 ( .A(n8044), .B(n8043), .Z(n8045) );
  NAND U10446 ( .A(n8046), .B(n8045), .Z(n8093) );
  AND U10447 ( .A(y[7748]), .B(x[487]), .Z(n8136) );
  NAND U10448 ( .A(n8136), .B(n8047), .Z(n8051) );
  NAND U10449 ( .A(n8049), .B(n8048), .Z(n8050) );
  AND U10450 ( .A(n8051), .B(n8050), .Z(n8149) );
  AND U10451 ( .A(y[7747]), .B(x[487]), .Z(n8053) );
  NAND U10452 ( .A(y[7750]), .B(x[484]), .Z(n8052) );
  XNOR U10453 ( .A(n8053), .B(n8052), .Z(n8120) );
  AND U10454 ( .A(x[486]), .B(y[7748]), .Z(n8119) );
  XOR U10455 ( .A(n8120), .B(n8119), .Z(n8147) );
  AND U10456 ( .A(x[488]), .B(y[7746]), .Z(n8314) );
  AND U10457 ( .A(x[489]), .B(y[7745]), .Z(n8130) );
  XOR U10458 ( .A(n8130), .B(o[74]), .Z(n8141) );
  XOR U10459 ( .A(n8314), .B(n8141), .Z(n8143) );
  XNOR U10460 ( .A(n8143), .B(n8142), .Z(n8146) );
  XOR U10461 ( .A(n8149), .B(n8148), .Z(n8109) );
  AND U10462 ( .A(x[489]), .B(y[7753]), .Z(n8054) );
  NAND U10463 ( .A(n8054), .B(n8465), .Z(n8058) );
  NAND U10464 ( .A(n8056), .B(n8055), .Z(n8057) );
  AND U10465 ( .A(n8058), .B(n8057), .Z(n8107) );
  AND U10466 ( .A(x[486]), .B(y[7752]), .Z(n8350) );
  NAND U10467 ( .A(n8350), .B(n8059), .Z(n8062) );
  NAND U10468 ( .A(n8470), .B(n8060), .Z(n8061) );
  NAND U10469 ( .A(n8062), .B(n8061), .Z(n8114) );
  ANDN U10470 ( .B(o[73]), .A(n8063), .Z(n8125) );
  AND U10471 ( .A(y[7744]), .B(x[490]), .Z(n8065) );
  AND U10472 ( .A(y[7754]), .B(x[480]), .Z(n8064) );
  XOR U10473 ( .A(n8065), .B(n8064), .Z(n8124) );
  XOR U10474 ( .A(n8125), .B(n8124), .Z(n8113) );
  AND U10475 ( .A(y[7751]), .B(x[483]), .Z(n9061) );
  NAND U10476 ( .A(y[7753]), .B(x[481]), .Z(n8066) );
  XNOR U10477 ( .A(n9061), .B(n8066), .Z(n8138) );
  AND U10478 ( .A(x[482]), .B(y[7752]), .Z(n8137) );
  XOR U10479 ( .A(n8138), .B(n8137), .Z(n8112) );
  XOR U10480 ( .A(n8113), .B(n8112), .Z(n8115) );
  XOR U10481 ( .A(n8114), .B(n8115), .Z(n8106) );
  XNOR U10482 ( .A(n8107), .B(n8106), .Z(n8108) );
  XOR U10483 ( .A(n8109), .B(n8108), .Z(n8092) );
  NANDN U10484 ( .A(n8072), .B(n8071), .Z(n8076) );
  NAND U10485 ( .A(n8074), .B(n8073), .Z(n8075) );
  AND U10486 ( .A(n8076), .B(n8075), .Z(n8100) );
  ANDN U10487 ( .B(n8718), .A(n8419), .Z(n8080) );
  NANDN U10488 ( .A(n8078), .B(n8077), .Z(n8079) );
  NANDN U10489 ( .A(n8080), .B(n8079), .Z(n8101) );
  XOR U10490 ( .A(n8100), .B(n8101), .Z(n8103) );
  XNOR U10491 ( .A(n8102), .B(n8103), .Z(n8091) );
  XOR U10492 ( .A(n8092), .B(n8091), .Z(n8094) );
  XOR U10493 ( .A(n8093), .B(n8094), .Z(n8099) );
  NANDN U10494 ( .A(n8082), .B(n8081), .Z(n8086) );
  NAND U10495 ( .A(n8084), .B(n8083), .Z(n8085) );
  NAND U10496 ( .A(n8086), .B(n8085), .Z(n8097) );
  XOR U10497 ( .A(n8097), .B(n8098), .Z(n8090) );
  XNOR U10498 ( .A(n8099), .B(n8090), .Z(N171) );
  NAND U10499 ( .A(n8092), .B(n8091), .Z(n8096) );
  NAND U10500 ( .A(n8094), .B(n8093), .Z(n8095) );
  NAND U10501 ( .A(n8096), .B(n8095), .Z(n8153) );
  NANDN U10502 ( .A(n8101), .B(n8100), .Z(n8105) );
  OR U10503 ( .A(n8103), .B(n8102), .Z(n8104) );
  AND U10504 ( .A(n8105), .B(n8104), .Z(n8159) );
  NANDN U10505 ( .A(n8107), .B(n8106), .Z(n8111) );
  NANDN U10506 ( .A(n8109), .B(n8108), .Z(n8110) );
  AND U10507 ( .A(n8111), .B(n8110), .Z(n8157) );
  NAND U10508 ( .A(n8113), .B(n8112), .Z(n8117) );
  NAND U10509 ( .A(n8115), .B(n8114), .Z(n8116) );
  NAND U10510 ( .A(n8117), .B(n8116), .Z(n8213) );
  AND U10511 ( .A(x[487]), .B(y[7750]), .Z(n8241) );
  AND U10512 ( .A(x[484]), .B(y[7747]), .Z(n8118) );
  NAND U10513 ( .A(n8241), .B(n8118), .Z(n8122) );
  NAND U10514 ( .A(n8120), .B(n8119), .Z(n8121) );
  NAND U10515 ( .A(n8122), .B(n8121), .Z(n8211) );
  AND U10516 ( .A(x[490]), .B(y[7754]), .Z(n8123) );
  NAND U10517 ( .A(n8123), .B(n8465), .Z(n8127) );
  NAND U10518 ( .A(n8125), .B(n8124), .Z(n8126) );
  NAND U10519 ( .A(n8127), .B(n8126), .Z(n8207) );
  AND U10520 ( .A(y[7744]), .B(x[491]), .Z(n8129) );
  NAND U10521 ( .A(y[7755]), .B(x[480]), .Z(n8128) );
  XNOR U10522 ( .A(n8129), .B(n8128), .Z(n8182) );
  NAND U10523 ( .A(n8130), .B(o[74]), .Z(n8183) );
  AND U10524 ( .A(y[7749]), .B(x[486]), .Z(n8132) );
  NAND U10525 ( .A(y[7754]), .B(x[481]), .Z(n8131) );
  XNOR U10526 ( .A(n8132), .B(n8131), .Z(n8174) );
  NAND U10527 ( .A(x[490]), .B(y[7745]), .Z(n8193) );
  XOR U10528 ( .A(n8174), .B(n8173), .Z(n8205) );
  XOR U10529 ( .A(n8206), .B(n8205), .Z(n8208) );
  XOR U10530 ( .A(n8207), .B(n8208), .Z(n8212) );
  XOR U10531 ( .A(n8211), .B(n8212), .Z(n8214) );
  XNOR U10532 ( .A(n8213), .B(n8214), .Z(n8196) );
  AND U10533 ( .A(x[483]), .B(y[7752]), .Z(n9194) );
  NAND U10534 ( .A(y[7753]), .B(x[482]), .Z(n8133) );
  XNOR U10535 ( .A(n8134), .B(n8133), .Z(n8169) );
  AND U10536 ( .A(x[484]), .B(y[7751]), .Z(n8168) );
  XNOR U10537 ( .A(n8169), .B(n8168), .Z(n8200) );
  XNOR U10538 ( .A(n9194), .B(n8200), .Z(n8201) );
  NAND U10539 ( .A(y[7746]), .B(x[489]), .Z(n8135) );
  XNOR U10540 ( .A(n8136), .B(n8135), .Z(n8187) );
  NAND U10541 ( .A(x[488]), .B(y[7747]), .Z(n8188) );
  NAND U10542 ( .A(x[483]), .B(y[7753]), .Z(n8237) );
  AND U10543 ( .A(x[481]), .B(y[7751]), .Z(n8460) );
  NANDN U10544 ( .A(n8237), .B(n8460), .Z(n8140) );
  NAND U10545 ( .A(n8138), .B(n8137), .Z(n8139) );
  NAND U10546 ( .A(n8140), .B(n8139), .Z(n8163) );
  NAND U10547 ( .A(n8314), .B(n8141), .Z(n8145) );
  NAND U10548 ( .A(n8143), .B(n8142), .Z(n8144) );
  NAND U10549 ( .A(n8145), .B(n8144), .Z(n8162) );
  XOR U10550 ( .A(n8163), .B(n8162), .Z(n8164) );
  NANDN U10551 ( .A(n8147), .B(n8146), .Z(n8151) );
  NAND U10552 ( .A(n8149), .B(n8148), .Z(n8150) );
  NAND U10553 ( .A(n8151), .B(n8150), .Z(n8194) );
  XOR U10554 ( .A(n8196), .B(n8197), .Z(n8156) );
  XNOR U10555 ( .A(n8157), .B(n8156), .Z(n8158) );
  XNOR U10556 ( .A(n8159), .B(n8158), .Z(n8155) );
  XNOR U10557 ( .A(n8154), .B(n8155), .Z(n8152) );
  XNOR U10558 ( .A(n8153), .B(n8152), .Z(N172) );
  NANDN U10559 ( .A(n8157), .B(n8156), .Z(n8161) );
  NANDN U10560 ( .A(n8159), .B(n8158), .Z(n8160) );
  NAND U10561 ( .A(n8161), .B(n8160), .Z(n8280) );
  NAND U10562 ( .A(n8163), .B(n8162), .Z(n8167) );
  NANDN U10563 ( .A(n8165), .B(n8164), .Z(n8166) );
  NAND U10564 ( .A(n8167), .B(n8166), .Z(n8276) );
  AND U10565 ( .A(x[485]), .B(y[7753]), .Z(n8709) );
  NAND U10566 ( .A(n8905), .B(n8709), .Z(n8171) );
  NAND U10567 ( .A(n8169), .B(n8168), .Z(n8170) );
  AND U10568 ( .A(n8171), .B(n8170), .Z(n8225) );
  AND U10569 ( .A(x[486]), .B(y[7754]), .Z(n8477) );
  NAND U10570 ( .A(n8477), .B(n8172), .Z(n8176) );
  NAND U10571 ( .A(n8174), .B(n8173), .Z(n8175) );
  NAND U10572 ( .A(n8176), .B(n8175), .Z(n8224) );
  AND U10573 ( .A(x[489]), .B(y[7747]), .Z(n8900) );
  AND U10574 ( .A(y[7746]), .B(x[490]), .Z(n8943) );
  NAND U10575 ( .A(y[7752]), .B(x[484]), .Z(n8177) );
  XOR U10576 ( .A(n8943), .B(n8177), .Z(n8267) );
  NAND U10577 ( .A(x[487]), .B(y[7749]), .Z(n8245) );
  XOR U10578 ( .A(n8246), .B(n8245), .Z(n8248) );
  AND U10579 ( .A(y[7744]), .B(x[492]), .Z(n8179) );
  NAND U10580 ( .A(y[7756]), .B(x[480]), .Z(n8178) );
  XNOR U10581 ( .A(n8179), .B(n8178), .Z(n8262) );
  AND U10582 ( .A(x[491]), .B(y[7745]), .Z(n8242) );
  XOR U10583 ( .A(o[76]), .B(n8242), .Z(n8261) );
  XOR U10584 ( .A(n8262), .B(n8261), .Z(n8231) );
  AND U10585 ( .A(y[7754]), .B(x[482]), .Z(n8181) );
  NAND U10586 ( .A(y[7748]), .B(x[488]), .Z(n8180) );
  XNOR U10587 ( .A(n8181), .B(n8180), .Z(n8236) );
  XOR U10588 ( .A(n8231), .B(n8230), .Z(n8233) );
  XOR U10589 ( .A(n8232), .B(n8233), .Z(n8226) );
  XOR U10590 ( .A(n8227), .B(n8226), .Z(n8274) );
  AND U10591 ( .A(x[491]), .B(y[7755]), .Z(n9304) );
  NAND U10592 ( .A(n9304), .B(n8465), .Z(n8185) );
  NANDN U10593 ( .A(n8183), .B(n8182), .Z(n8184) );
  AND U10594 ( .A(n8185), .B(n8184), .Z(n8254) );
  AND U10595 ( .A(x[487]), .B(y[7746]), .Z(n8395) );
  AND U10596 ( .A(x[489]), .B(y[7748]), .Z(n8186) );
  NAND U10597 ( .A(n8395), .B(n8186), .Z(n8190) );
  NANDN U10598 ( .A(n8188), .B(n8187), .Z(n8189) );
  AND U10599 ( .A(n8190), .B(n8189), .Z(n8252) );
  NAND U10600 ( .A(y[7755]), .B(x[481]), .Z(n8191) );
  XNOR U10601 ( .A(n8192), .B(n8191), .Z(n8258) );
  ANDN U10602 ( .B(o[75]), .A(n8193), .Z(n8257) );
  XOR U10603 ( .A(n8258), .B(n8257), .Z(n8251) );
  XNOR U10604 ( .A(n8274), .B(n8275), .Z(n8277) );
  XOR U10605 ( .A(n8276), .B(n8277), .Z(n8284) );
  NANDN U10606 ( .A(n8195), .B(n8194), .Z(n8199) );
  NANDN U10607 ( .A(n8197), .B(n8196), .Z(n8198) );
  NAND U10608 ( .A(n8199), .B(n8198), .Z(n8283) );
  NANDN U10609 ( .A(n9194), .B(n8200), .Z(n8204) );
  NANDN U10610 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U10611 ( .A(n8204), .B(n8203), .Z(n8218) );
  NAND U10612 ( .A(n8206), .B(n8205), .Z(n8210) );
  NAND U10613 ( .A(n8208), .B(n8207), .Z(n8209) );
  AND U10614 ( .A(n8210), .B(n8209), .Z(n8219) );
  XOR U10615 ( .A(n8218), .B(n8219), .Z(n8221) );
  NAND U10616 ( .A(n8212), .B(n8211), .Z(n8216) );
  NAND U10617 ( .A(n8214), .B(n8213), .Z(n8215) );
  AND U10618 ( .A(n8216), .B(n8215), .Z(n8220) );
  XOR U10619 ( .A(n8221), .B(n8220), .Z(n8285) );
  XOR U10620 ( .A(n8286), .B(n8285), .Z(n8282) );
  XOR U10621 ( .A(n8280), .B(n8282), .Z(n8217) );
  XNOR U10622 ( .A(n8281), .B(n8217), .Z(N173) );
  NAND U10623 ( .A(n8219), .B(n8218), .Z(n8223) );
  NAND U10624 ( .A(n8221), .B(n8220), .Z(n8222) );
  NAND U10625 ( .A(n8223), .B(n8222), .Z(n8366) );
  NANDN U10626 ( .A(n8225), .B(n8224), .Z(n8229) );
  NAND U10627 ( .A(n8227), .B(n8226), .Z(n8228) );
  AND U10628 ( .A(n8229), .B(n8228), .Z(n8291) );
  NAND U10629 ( .A(n8231), .B(n8230), .Z(n8235) );
  NAND U10630 ( .A(n8233), .B(n8232), .Z(n8234) );
  NAND U10631 ( .A(n8235), .B(n8234), .Z(n8298) );
  AND U10632 ( .A(y[7754]), .B(x[488]), .Z(n9548) );
  AND U10633 ( .A(x[482]), .B(y[7748]), .Z(n8405) );
  NAND U10634 ( .A(n9548), .B(n8405), .Z(n8239) );
  NANDN U10635 ( .A(n8237), .B(n8236), .Z(n8238) );
  AND U10636 ( .A(n8239), .B(n8238), .Z(n8329) );
  NAND U10637 ( .A(y[7756]), .B(x[481]), .Z(n8240) );
  XNOR U10638 ( .A(n8241), .B(n8240), .Z(n8320) );
  AND U10639 ( .A(o[76]), .B(n8242), .Z(n8319) );
  XOR U10640 ( .A(n8320), .B(n8319), .Z(n8327) );
  AND U10641 ( .A(x[486]), .B(y[7751]), .Z(n9344) );
  AND U10642 ( .A(y[7755]), .B(x[482]), .Z(n8244) );
  NAND U10643 ( .A(y[7748]), .B(x[489]), .Z(n8243) );
  XNOR U10644 ( .A(n8244), .B(n8243), .Z(n8333) );
  XOR U10645 ( .A(n9344), .B(n8333), .Z(n8326) );
  XOR U10646 ( .A(n8327), .B(n8326), .Z(n8328) );
  NAND U10647 ( .A(n8246), .B(n8245), .Z(n8250) );
  ANDN U10648 ( .B(n8248), .A(n8247), .Z(n8249) );
  ANDN U10649 ( .B(n8250), .A(n8249), .Z(n8296) );
  XOR U10650 ( .A(n8297), .B(n8296), .Z(n8299) );
  XOR U10651 ( .A(n8298), .B(n8299), .Z(n8290) );
  NANDN U10652 ( .A(n8252), .B(n8251), .Z(n8256) );
  NANDN U10653 ( .A(n8254), .B(n8253), .Z(n8255) );
  AND U10654 ( .A(n8256), .B(n8255), .Z(n8305) );
  NAND U10655 ( .A(x[486]), .B(y[7755]), .Z(n8711) );
  AND U10656 ( .A(x[481]), .B(y[7750]), .Z(n8318) );
  NANDN U10657 ( .A(n8711), .B(n8318), .Z(n8260) );
  NAND U10658 ( .A(n8258), .B(n8257), .Z(n8259) );
  AND U10659 ( .A(n8260), .B(n8259), .Z(n8311) );
  AND U10660 ( .A(x[492]), .B(y[7756]), .Z(n9556) );
  NAND U10661 ( .A(n9556), .B(n8465), .Z(n8264) );
  NAND U10662 ( .A(n8262), .B(n8261), .Z(n8263) );
  AND U10663 ( .A(n8264), .B(n8263), .Z(n8309) );
  AND U10664 ( .A(x[490]), .B(y[7747]), .Z(n9206) );
  AND U10665 ( .A(y[7746]), .B(x[491]), .Z(n9167) );
  NAND U10666 ( .A(y[7749]), .B(x[488]), .Z(n8265) );
  XNOR U10667 ( .A(n9167), .B(n8265), .Z(n8315) );
  XOR U10668 ( .A(n9206), .B(n8315), .Z(n8308) );
  AND U10669 ( .A(x[490]), .B(y[7752]), .Z(n8677) );
  AND U10670 ( .A(x[484]), .B(y[7746]), .Z(n8266) );
  NAND U10671 ( .A(n8677), .B(n8266), .Z(n8269) );
  NANDN U10672 ( .A(n8267), .B(n8900), .Z(n8268) );
  AND U10673 ( .A(n8269), .B(n8268), .Z(n8354) );
  AND U10674 ( .A(y[7744]), .B(x[493]), .Z(n8271) );
  NAND U10675 ( .A(y[7757]), .B(x[480]), .Z(n8270) );
  XNOR U10676 ( .A(n8271), .B(n8270), .Z(n8346) );
  AND U10677 ( .A(x[492]), .B(y[7745]), .Z(n8338) );
  XOR U10678 ( .A(o[77]), .B(n8338), .Z(n8345) );
  XOR U10679 ( .A(n8346), .B(n8345), .Z(n8352) );
  AND U10680 ( .A(y[7752]), .B(x[485]), .Z(n8273) );
  NAND U10681 ( .A(y[7754]), .B(x[483]), .Z(n8272) );
  XNOR U10682 ( .A(n8273), .B(n8272), .Z(n8341) );
  AND U10683 ( .A(x[484]), .B(y[7753]), .Z(n8342) );
  XOR U10684 ( .A(n8341), .B(n8342), .Z(n8351) );
  XOR U10685 ( .A(n8352), .B(n8351), .Z(n8353) );
  XOR U10686 ( .A(n8303), .B(n8302), .Z(n8304) );
  XOR U10687 ( .A(n8293), .B(n8292), .Z(n8365) );
  NANDN U10688 ( .A(n8275), .B(n8274), .Z(n8279) );
  NAND U10689 ( .A(n8277), .B(n8276), .Z(n8278) );
  AND U10690 ( .A(n8279), .B(n8278), .Z(n8364) );
  XOR U10691 ( .A(n8366), .B(n8367), .Z(n8360) );
  NANDN U10692 ( .A(n8284), .B(n8283), .Z(n8288) );
  NAND U10693 ( .A(n8286), .B(n8285), .Z(n8287) );
  AND U10694 ( .A(n8288), .B(n8287), .Z(n8358) );
  IV U10695 ( .A(n8358), .Z(n8357) );
  XOR U10696 ( .A(n8359), .B(n8357), .Z(n8289) );
  XNOR U10697 ( .A(n8360), .B(n8289), .Z(N174) );
  NANDN U10698 ( .A(n8291), .B(n8290), .Z(n8295) );
  NAND U10699 ( .A(n8293), .B(n8292), .Z(n8294) );
  AND U10700 ( .A(n8295), .B(n8294), .Z(n8454) );
  NAND U10701 ( .A(n8297), .B(n8296), .Z(n8301) );
  NAND U10702 ( .A(n8299), .B(n8298), .Z(n8300) );
  NAND U10703 ( .A(n8301), .B(n8300), .Z(n8453) );
  NAND U10704 ( .A(n8303), .B(n8302), .Z(n8307) );
  NANDN U10705 ( .A(n8305), .B(n8304), .Z(n8306) );
  AND U10706 ( .A(n8307), .B(n8306), .Z(n8374) );
  NANDN U10707 ( .A(n8309), .B(n8308), .Z(n8313) );
  NANDN U10708 ( .A(n8311), .B(n8310), .Z(n8312) );
  AND U10709 ( .A(n8313), .B(n8312), .Z(n8380) );
  AND U10710 ( .A(x[491]), .B(y[7749]), .Z(n8491) );
  NAND U10711 ( .A(n8491), .B(n8314), .Z(n8317) );
  NAND U10712 ( .A(n8315), .B(n9206), .Z(n8316) );
  NAND U10713 ( .A(n8317), .B(n8316), .Z(n8435) );
  AND U10714 ( .A(x[487]), .B(y[7756]), .Z(n8914) );
  NAND U10715 ( .A(n8914), .B(n8318), .Z(n8322) );
  NAND U10716 ( .A(n8320), .B(n8319), .Z(n8321) );
  NAND U10717 ( .A(n8322), .B(n8321), .Z(n8434) );
  XOR U10718 ( .A(n8435), .B(n8434), .Z(n8437) );
  AND U10719 ( .A(x[484]), .B(y[7754]), .Z(n8820) );
  AND U10720 ( .A(y[7755]), .B(x[483]), .Z(n8324) );
  NAND U10721 ( .A(y[7750]), .B(x[488]), .Z(n8323) );
  XNOR U10722 ( .A(n8324), .B(n8323), .Z(n8420) );
  XOR U10723 ( .A(n8709), .B(n8420), .Z(n8429) );
  XOR U10724 ( .A(n8820), .B(n8429), .Z(n8431) );
  AND U10725 ( .A(x[489]), .B(y[7749]), .Z(n9032) );
  AND U10726 ( .A(y[7756]), .B(x[482]), .Z(n8325) );
  AND U10727 ( .A(x[490]), .B(y[7748]), .Z(n9056) );
  XOR U10728 ( .A(n8325), .B(n9056), .Z(n8406) );
  XOR U10729 ( .A(n9032), .B(n8406), .Z(n8430) );
  XOR U10730 ( .A(n8431), .B(n8430), .Z(n8436) );
  XOR U10731 ( .A(n8437), .B(n8436), .Z(n8378) );
  NAND U10732 ( .A(n8327), .B(n8326), .Z(n8331) );
  NANDN U10733 ( .A(n8329), .B(n8328), .Z(n8330) );
  AND U10734 ( .A(n8331), .B(n8330), .Z(n8377) );
  XOR U10735 ( .A(n8380), .B(n8379), .Z(n8372) );
  AND U10736 ( .A(x[489]), .B(y[7755]), .Z(n8332) );
  NAND U10737 ( .A(n8332), .B(n8405), .Z(n8335) );
  NAND U10738 ( .A(n8333), .B(n9344), .Z(n8334) );
  NAND U10739 ( .A(n8335), .B(n8334), .Z(n8392) );
  AND U10740 ( .A(y[7744]), .B(x[494]), .Z(n8337) );
  NAND U10741 ( .A(y[7758]), .B(x[480]), .Z(n8336) );
  XNOR U10742 ( .A(n8337), .B(n8336), .Z(n8415) );
  AND U10743 ( .A(o[77]), .B(n8338), .Z(n8414) );
  XOR U10744 ( .A(n8415), .B(n8414), .Z(n8390) );
  NAND U10745 ( .A(y[7746]), .B(x[492]), .Z(n8339) );
  XNOR U10746 ( .A(n8340), .B(n8339), .Z(n8397) );
  AND U10747 ( .A(x[493]), .B(y[7745]), .Z(n8404) );
  XOR U10748 ( .A(o[78]), .B(n8404), .Z(n8396) );
  XOR U10749 ( .A(n8397), .B(n8396), .Z(n8389) );
  XOR U10750 ( .A(n8390), .B(n8389), .Z(n8391) );
  XNOR U10751 ( .A(n8392), .B(n8391), .Z(n8441) );
  AND U10752 ( .A(x[485]), .B(y[7754]), .Z(n8478) );
  NAND U10753 ( .A(n9194), .B(n8478), .Z(n8344) );
  NAND U10754 ( .A(n8342), .B(n8341), .Z(n8343) );
  AND U10755 ( .A(n8344), .B(n8343), .Z(n8386) );
  AND U10756 ( .A(x[493]), .B(y[7757]), .Z(n9945) );
  NAND U10757 ( .A(n9945), .B(n8465), .Z(n8348) );
  NAND U10758 ( .A(n8346), .B(n8345), .Z(n8347) );
  NAND U10759 ( .A(n8348), .B(n8347), .Z(n8384) );
  NAND U10760 ( .A(y[7747]), .B(x[491]), .Z(n8349) );
  XNOR U10761 ( .A(n8350), .B(n8349), .Z(n8410) );
  AND U10762 ( .A(x[481]), .B(y[7757]), .Z(n8411) );
  XOR U10763 ( .A(n8410), .B(n8411), .Z(n8383) );
  XOR U10764 ( .A(n8384), .B(n8383), .Z(n8385) );
  XOR U10765 ( .A(n8386), .B(n8385), .Z(n8440) );
  XOR U10766 ( .A(n8441), .B(n8440), .Z(n8443) );
  NAND U10767 ( .A(n8352), .B(n8351), .Z(n8356) );
  NANDN U10768 ( .A(n8354), .B(n8353), .Z(n8355) );
  AND U10769 ( .A(n8356), .B(n8355), .Z(n8442) );
  XNOR U10770 ( .A(n8443), .B(n8442), .Z(n8371) );
  XNOR U10771 ( .A(n8456), .B(n8455), .Z(n8449) );
  OR U10772 ( .A(n8359), .B(n8357), .Z(n8363) );
  ANDN U10773 ( .B(n8359), .A(n8358), .Z(n8361) );
  OR U10774 ( .A(n8361), .B(n8360), .Z(n8362) );
  AND U10775 ( .A(n8363), .B(n8362), .Z(n8448) );
  NANDN U10776 ( .A(n8365), .B(n8364), .Z(n8369) );
  NAND U10777 ( .A(n8367), .B(n8366), .Z(n8368) );
  AND U10778 ( .A(n8369), .B(n8368), .Z(n8447) );
  IV U10779 ( .A(n8447), .Z(n8446) );
  XOR U10780 ( .A(n8448), .B(n8446), .Z(n8370) );
  XNOR U10781 ( .A(n8449), .B(n8370), .Z(N175) );
  NANDN U10782 ( .A(n8372), .B(n8371), .Z(n8376) );
  NANDN U10783 ( .A(n8374), .B(n8373), .Z(n8375) );
  AND U10784 ( .A(n8376), .B(n8375), .Z(n8552) );
  NANDN U10785 ( .A(n8378), .B(n8377), .Z(n8382) );
  NAND U10786 ( .A(n8380), .B(n8379), .Z(n8381) );
  AND U10787 ( .A(n8382), .B(n8381), .Z(n8521) );
  NAND U10788 ( .A(n8384), .B(n8383), .Z(n8388) );
  NANDN U10789 ( .A(n8386), .B(n8385), .Z(n8387) );
  NAND U10790 ( .A(n8388), .B(n8387), .Z(n8527) );
  NAND U10791 ( .A(n8390), .B(n8389), .Z(n8394) );
  NAND U10792 ( .A(n8392), .B(n8391), .Z(n8393) );
  NAND U10793 ( .A(n8394), .B(n8393), .Z(n8525) );
  AND U10794 ( .A(x[492]), .B(y[7751]), .Z(n8906) );
  NAND U10795 ( .A(n8906), .B(n8395), .Z(n8399) );
  NAND U10796 ( .A(n8397), .B(n8396), .Z(n8398) );
  AND U10797 ( .A(n8399), .B(n8398), .Z(n8501) );
  AND U10798 ( .A(y[7748]), .B(x[491]), .Z(n8401) );
  NAND U10799 ( .A(y[7746]), .B(x[493]), .Z(n8400) );
  XNOR U10800 ( .A(n8401), .B(n8400), .Z(n8505) );
  AND U10801 ( .A(x[492]), .B(y[7747]), .Z(n8504) );
  XNOR U10802 ( .A(n8505), .B(n8504), .Z(n8499) );
  AND U10803 ( .A(y[7744]), .B(x[495]), .Z(n8403) );
  NAND U10804 ( .A(y[7759]), .B(x[480]), .Z(n8402) );
  XNOR U10805 ( .A(n8403), .B(n8402), .Z(n8467) );
  AND U10806 ( .A(o[78]), .B(n8404), .Z(n8466) );
  XNOR U10807 ( .A(n8467), .B(n8466), .Z(n8498) );
  XOR U10808 ( .A(n8499), .B(n8498), .Z(n8500) );
  XNOR U10809 ( .A(n8501), .B(n8500), .Z(n8533) );
  NAND U10810 ( .A(x[490]), .B(y[7756]), .Z(n9346) );
  NANDN U10811 ( .A(n9346), .B(n8405), .Z(n8408) );
  NAND U10812 ( .A(n9032), .B(n8406), .Z(n8407) );
  NAND U10813 ( .A(n8408), .B(n8407), .Z(n8531) );
  AND U10814 ( .A(x[491]), .B(y[7752]), .Z(n8819) );
  NAND U10815 ( .A(n8819), .B(n8409), .Z(n8413) );
  NAND U10816 ( .A(n8411), .B(n8410), .Z(n8412) );
  NAND U10817 ( .A(n8413), .B(n8412), .Z(n8530) );
  XOR U10818 ( .A(n8531), .B(n8530), .Z(n8532) );
  XOR U10819 ( .A(n8533), .B(n8532), .Z(n8524) );
  XOR U10820 ( .A(n8525), .B(n8524), .Z(n8526) );
  XNOR U10821 ( .A(n8527), .B(n8526), .Z(n8518) );
  AND U10822 ( .A(x[494]), .B(y[7758]), .Z(n10203) );
  NAND U10823 ( .A(n10203), .B(n8465), .Z(n8417) );
  NAND U10824 ( .A(n8415), .B(n8414), .Z(n8416) );
  NAND U10825 ( .A(n8417), .B(n8416), .Z(n8493) );
  AND U10826 ( .A(x[488]), .B(y[7755]), .Z(n8418) );
  NAND U10827 ( .A(n8419), .B(n8418), .Z(n8422) );
  NAND U10828 ( .A(n8420), .B(n8709), .Z(n8421) );
  NAND U10829 ( .A(n8422), .B(n8421), .Z(n8492) );
  XOR U10830 ( .A(n8493), .B(n8492), .Z(n8495) );
  AND U10831 ( .A(y[7749]), .B(x[490]), .Z(n8424) );
  NAND U10832 ( .A(y[7755]), .B(x[484]), .Z(n8423) );
  XNOR U10833 ( .A(n8424), .B(n8423), .Z(n8473) );
  AND U10834 ( .A(x[487]), .B(y[7752]), .Z(n8472) );
  XNOR U10835 ( .A(n8473), .B(n8472), .Z(n8480) );
  NAND U10836 ( .A(x[486]), .B(y[7753]), .Z(n8583) );
  XNOR U10837 ( .A(n8583), .B(n8478), .Z(n8479) );
  XNOR U10838 ( .A(n8480), .B(n8479), .Z(n8514) );
  AND U10839 ( .A(y[7757]), .B(x[482]), .Z(n8426) );
  NAND U10840 ( .A(y[7750]), .B(x[489]), .Z(n8425) );
  XNOR U10841 ( .A(n8426), .B(n8425), .Z(n8483) );
  AND U10842 ( .A(x[483]), .B(y[7756]), .Z(n8484) );
  XOR U10843 ( .A(n8483), .B(n8484), .Z(n8513) );
  AND U10844 ( .A(y[7758]), .B(x[481]), .Z(n8428) );
  NAND U10845 ( .A(y[7751]), .B(x[488]), .Z(n8427) );
  XNOR U10846 ( .A(n8428), .B(n8427), .Z(n8462) );
  AND U10847 ( .A(x[494]), .B(y[7745]), .Z(n8489) );
  XOR U10848 ( .A(o[79]), .B(n8489), .Z(n8461) );
  XOR U10849 ( .A(n8462), .B(n8461), .Z(n8512) );
  XOR U10850 ( .A(n8513), .B(n8512), .Z(n8515) );
  XOR U10851 ( .A(n8514), .B(n8515), .Z(n8494) );
  XNOR U10852 ( .A(n8495), .B(n8494), .Z(n8537) );
  NAND U10853 ( .A(n8820), .B(n8429), .Z(n8433) );
  NAND U10854 ( .A(n8431), .B(n8430), .Z(n8432) );
  AND U10855 ( .A(n8433), .B(n8432), .Z(n8536) );
  XOR U10856 ( .A(n8537), .B(n8536), .Z(n8538) );
  NAND U10857 ( .A(n8435), .B(n8434), .Z(n8439) );
  NAND U10858 ( .A(n8437), .B(n8436), .Z(n8438) );
  AND U10859 ( .A(n8439), .B(n8438), .Z(n8539) );
  XOR U10860 ( .A(n8538), .B(n8539), .Z(n8519) );
  XOR U10861 ( .A(n8518), .B(n8519), .Z(n8520) );
  NAND U10862 ( .A(n8441), .B(n8440), .Z(n8445) );
  NAND U10863 ( .A(n8443), .B(n8442), .Z(n8444) );
  AND U10864 ( .A(n8445), .B(n8444), .Z(n8550) );
  XOR U10865 ( .A(n8549), .B(n8550), .Z(n8551) );
  XOR U10866 ( .A(n8552), .B(n8551), .Z(n8545) );
  OR U10867 ( .A(n8448), .B(n8446), .Z(n8452) );
  ANDN U10868 ( .B(n8448), .A(n8447), .Z(n8450) );
  OR U10869 ( .A(n8450), .B(n8449), .Z(n8451) );
  AND U10870 ( .A(n8452), .B(n8451), .Z(n8544) );
  NANDN U10871 ( .A(n8454), .B(n8453), .Z(n8458) );
  NAND U10872 ( .A(n8456), .B(n8455), .Z(n8457) );
  NAND U10873 ( .A(n8458), .B(n8457), .Z(n8543) );
  IV U10874 ( .A(n8543), .Z(n8542) );
  XOR U10875 ( .A(n8544), .B(n8542), .Z(n8459) );
  XNOR U10876 ( .A(n8545), .B(n8459), .Z(N176) );
  AND U10877 ( .A(x[488]), .B(y[7758]), .Z(n8821) );
  NAND U10878 ( .A(n8821), .B(n8460), .Z(n8464) );
  NAND U10879 ( .A(n8462), .B(n8461), .Z(n8463) );
  AND U10880 ( .A(n8464), .B(n8463), .Z(n8613) );
  AND U10881 ( .A(x[495]), .B(y[7759]), .Z(n10643) );
  NAND U10882 ( .A(n10643), .B(n8465), .Z(n8469) );
  NAND U10883 ( .A(n8467), .B(n8466), .Z(n8468) );
  NAND U10884 ( .A(n8469), .B(n8468), .Z(n8612) );
  AND U10885 ( .A(x[490]), .B(y[7755]), .Z(n8471) );
  NAND U10886 ( .A(n8471), .B(n8470), .Z(n8475) );
  NAND U10887 ( .A(n8473), .B(n8472), .Z(n8474) );
  NAND U10888 ( .A(n8475), .B(n8474), .Z(n8570) );
  AND U10889 ( .A(x[480]), .B(y[7760]), .Z(n8592) );
  AND U10890 ( .A(x[496]), .B(y[7744]), .Z(n8593) );
  XOR U10891 ( .A(n8592), .B(n8593), .Z(n8595) );
  NAND U10892 ( .A(x[495]), .B(y[7745]), .Z(n8580) );
  XOR U10893 ( .A(n8595), .B(n8594), .Z(n8569) );
  NAND U10894 ( .A(y[7753]), .B(x[487]), .Z(n8476) );
  XNOR U10895 ( .A(n8477), .B(n8476), .Z(n8585) );
  AND U10896 ( .A(x[490]), .B(y[7750]), .Z(n8584) );
  XOR U10897 ( .A(n8585), .B(n8584), .Z(n8568) );
  XOR U10898 ( .A(n8569), .B(n8568), .Z(n8571) );
  XOR U10899 ( .A(n8570), .B(n8571), .Z(n8614) );
  XNOR U10900 ( .A(n8615), .B(n8614), .Z(n8565) );
  NANDN U10901 ( .A(n8478), .B(n8583), .Z(n8482) );
  NAND U10902 ( .A(n8480), .B(n8479), .Z(n8481) );
  NAND U10903 ( .A(n8482), .B(n8481), .Z(n8563) );
  NAND U10904 ( .A(x[489]), .B(y[7757]), .Z(n9327) );
  NANDN U10905 ( .A(n9327), .B(n8905), .Z(n8486) );
  NAND U10906 ( .A(n8484), .B(n8483), .Z(n8485) );
  AND U10907 ( .A(n8486), .B(n8485), .Z(n8603) );
  AND U10908 ( .A(y[7759]), .B(x[481]), .Z(n8488) );
  NAND U10909 ( .A(y[7752]), .B(x[488]), .Z(n8487) );
  XNOR U10910 ( .A(n8488), .B(n8487), .Z(n8589) );
  AND U10911 ( .A(o[79]), .B(n8489), .Z(n8588) );
  XOR U10912 ( .A(n8589), .B(n8588), .Z(n8601) );
  NAND U10913 ( .A(y[7746]), .B(x[494]), .Z(n8490) );
  XNOR U10914 ( .A(n8491), .B(n8490), .Z(n8624) );
  AND U10915 ( .A(x[484]), .B(y[7756]), .Z(n8625) );
  XOR U10916 ( .A(n8624), .B(n8625), .Z(n8600) );
  XOR U10917 ( .A(n8601), .B(n8600), .Z(n8602) );
  XOR U10918 ( .A(n8603), .B(n8602), .Z(n8562) );
  XOR U10919 ( .A(n8563), .B(n8562), .Z(n8564) );
  XOR U10920 ( .A(n8565), .B(n8564), .Z(n8606) );
  NAND U10921 ( .A(n8493), .B(n8492), .Z(n8497) );
  NAND U10922 ( .A(n8495), .B(n8494), .Z(n8496) );
  AND U10923 ( .A(n8497), .B(n8496), .Z(n8607) );
  XOR U10924 ( .A(n8606), .B(n8607), .Z(n8609) );
  NAND U10925 ( .A(n8499), .B(n8498), .Z(n8503) );
  NAND U10926 ( .A(n8501), .B(n8500), .Z(n8502) );
  NAND U10927 ( .A(n8503), .B(n8502), .Z(n8638) );
  AND U10928 ( .A(x[493]), .B(y[7748]), .Z(n8634) );
  NAND U10929 ( .A(n9167), .B(n8634), .Z(n8507) );
  NAND U10930 ( .A(n8505), .B(n8504), .Z(n8506) );
  NAND U10931 ( .A(n8507), .B(n8506), .Z(n8621) );
  AND U10932 ( .A(y[7758]), .B(x[482]), .Z(n8509) );
  NAND U10933 ( .A(y[7751]), .B(x[489]), .Z(n8508) );
  XNOR U10934 ( .A(n8509), .B(n8508), .Z(n8628) );
  AND U10935 ( .A(x[483]), .B(y[7757]), .Z(n8629) );
  XOR U10936 ( .A(n8628), .B(n8629), .Z(n8619) );
  AND U10937 ( .A(x[492]), .B(y[7748]), .Z(n9315) );
  AND U10938 ( .A(y[7755]), .B(x[485]), .Z(n8511) );
  NAND U10939 ( .A(y[7747]), .B(x[493]), .Z(n8510) );
  XNOR U10940 ( .A(n8511), .B(n8510), .Z(n8575) );
  XOR U10941 ( .A(n9315), .B(n8575), .Z(n8618) );
  XOR U10942 ( .A(n8619), .B(n8618), .Z(n8620) );
  XNOR U10943 ( .A(n8621), .B(n8620), .Z(n8635) );
  NAND U10944 ( .A(n8513), .B(n8512), .Z(n8517) );
  NAND U10945 ( .A(n8515), .B(n8514), .Z(n8516) );
  AND U10946 ( .A(n8517), .B(n8516), .Z(n8636) );
  XOR U10947 ( .A(n8635), .B(n8636), .Z(n8637) );
  XOR U10948 ( .A(n8638), .B(n8637), .Z(n8608) );
  XOR U10949 ( .A(n8609), .B(n8608), .Z(n8649) );
  NAND U10950 ( .A(n8519), .B(n8518), .Z(n8523) );
  NANDN U10951 ( .A(n8521), .B(n8520), .Z(n8522) );
  AND U10952 ( .A(n8523), .B(n8522), .Z(n8648) );
  NAND U10953 ( .A(n8525), .B(n8524), .Z(n8529) );
  NAND U10954 ( .A(n8527), .B(n8526), .Z(n8528) );
  NAND U10955 ( .A(n8529), .B(n8528), .Z(n8559) );
  NAND U10956 ( .A(n8531), .B(n8530), .Z(n8535) );
  NAND U10957 ( .A(n8533), .B(n8532), .Z(n8534) );
  NAND U10958 ( .A(n8535), .B(n8534), .Z(n8557) );
  NAND U10959 ( .A(n8537), .B(n8536), .Z(n8541) );
  NAND U10960 ( .A(n8539), .B(n8538), .Z(n8540) );
  AND U10961 ( .A(n8541), .B(n8540), .Z(n8556) );
  XOR U10962 ( .A(n8557), .B(n8556), .Z(n8558) );
  XOR U10963 ( .A(n8559), .B(n8558), .Z(n8650) );
  XNOR U10964 ( .A(n8651), .B(n8650), .Z(n8644) );
  OR U10965 ( .A(n8544), .B(n8542), .Z(n8548) );
  ANDN U10966 ( .B(n8544), .A(n8543), .Z(n8546) );
  OR U10967 ( .A(n8546), .B(n8545), .Z(n8547) );
  AND U10968 ( .A(n8548), .B(n8547), .Z(n8643) );
  NAND U10969 ( .A(n8550), .B(n8549), .Z(n8554) );
  NANDN U10970 ( .A(n8552), .B(n8551), .Z(n8553) );
  NAND U10971 ( .A(n8554), .B(n8553), .Z(n8642) );
  IV U10972 ( .A(n8642), .Z(n8641) );
  XOR U10973 ( .A(n8643), .B(n8641), .Z(n8555) );
  XNOR U10974 ( .A(n8644), .B(n8555), .Z(N177) );
  NAND U10975 ( .A(n8557), .B(n8556), .Z(n8561) );
  NAND U10976 ( .A(n8559), .B(n8558), .Z(n8560) );
  AND U10977 ( .A(n8561), .B(n8560), .Z(n8759) );
  NAND U10978 ( .A(n8563), .B(n8562), .Z(n8567) );
  NAND U10979 ( .A(n8565), .B(n8564), .Z(n8566) );
  NAND U10980 ( .A(n8567), .B(n8566), .Z(n8664) );
  NAND U10981 ( .A(n8569), .B(n8568), .Z(n8573) );
  NAND U10982 ( .A(n8571), .B(n8570), .Z(n8572) );
  AND U10983 ( .A(n8573), .B(n8572), .Z(n8746) );
  AND U10984 ( .A(x[493]), .B(y[7755]), .Z(n9562) );
  NAND U10985 ( .A(n9562), .B(n8574), .Z(n8577) );
  NAND U10986 ( .A(n8575), .B(n9315), .Z(n8576) );
  NAND U10987 ( .A(n8577), .B(n8576), .Z(n8694) );
  AND U10988 ( .A(y[7760]), .B(x[481]), .Z(n8579) );
  NAND U10989 ( .A(y[7752]), .B(x[489]), .Z(n8578) );
  XNOR U10990 ( .A(n8579), .B(n8578), .Z(n8715) );
  ANDN U10991 ( .B(o[80]), .A(n8580), .Z(n8714) );
  XOR U10992 ( .A(n8715), .B(n8714), .Z(n8692) );
  AND U10993 ( .A(y[7746]), .B(x[495]), .Z(n8582) );
  NAND U10994 ( .A(y[7749]), .B(x[492]), .Z(n8581) );
  XNOR U10995 ( .A(n8582), .B(n8581), .Z(n8667) );
  NAND U10996 ( .A(x[494]), .B(y[7747]), .Z(n8668) );
  XOR U10997 ( .A(n8692), .B(n8691), .Z(n8693) );
  XOR U10998 ( .A(n8694), .B(n8693), .Z(n8744) );
  AND U10999 ( .A(x[487]), .B(y[7754]), .Z(n8726) );
  NANDN U11000 ( .A(n8583), .B(n8726), .Z(n8587) );
  NAND U11001 ( .A(n8585), .B(n8584), .Z(n8586) );
  NAND U11002 ( .A(n8587), .B(n8586), .Z(n8704) );
  NAND U11003 ( .A(x[488]), .B(y[7759]), .Z(n9465) );
  AND U11004 ( .A(x[481]), .B(y[7752]), .Z(n8799) );
  NANDN U11005 ( .A(n9465), .B(n8799), .Z(n8591) );
  NAND U11006 ( .A(n8589), .B(n8588), .Z(n8590) );
  NAND U11007 ( .A(n8591), .B(n8590), .Z(n8703) );
  XOR U11008 ( .A(n8704), .B(n8703), .Z(n8706) );
  NAND U11009 ( .A(n8593), .B(n8592), .Z(n8597) );
  NAND U11010 ( .A(n8595), .B(n8594), .Z(n8596) );
  NAND U11011 ( .A(n8597), .B(n8596), .Z(n8700) );
  AND U11012 ( .A(x[480]), .B(y[7761]), .Z(n8681) );
  NAND U11013 ( .A(x[497]), .B(y[7744]), .Z(n8682) );
  AND U11014 ( .A(x[496]), .B(y[7745]), .Z(n8676) );
  XOR U11015 ( .A(o[81]), .B(n8676), .Z(n8683) );
  XOR U11016 ( .A(n8684), .B(n8683), .Z(n8698) );
  AND U11017 ( .A(y[7759]), .B(x[482]), .Z(n8599) );
  NAND U11018 ( .A(y[7751]), .B(x[490]), .Z(n8598) );
  XNOR U11019 ( .A(n8599), .B(n8598), .Z(n8719) );
  NAND U11020 ( .A(x[483]), .B(y[7758]), .Z(n8720) );
  XOR U11021 ( .A(n8698), .B(n8697), .Z(n8699) );
  XOR U11022 ( .A(n8700), .B(n8699), .Z(n8705) );
  XOR U11023 ( .A(n8706), .B(n8705), .Z(n8743) );
  XOR U11024 ( .A(n8744), .B(n8743), .Z(n8745) );
  NAND U11025 ( .A(n8601), .B(n8600), .Z(n8605) );
  NANDN U11026 ( .A(n8603), .B(n8602), .Z(n8604) );
  AND U11027 ( .A(n8605), .B(n8604), .Z(n8662) );
  XOR U11028 ( .A(n8661), .B(n8662), .Z(n8663) );
  XNOR U11029 ( .A(n8664), .B(n8663), .Z(n8757) );
  NAND U11030 ( .A(n8607), .B(n8606), .Z(n8611) );
  NAND U11031 ( .A(n8609), .B(n8608), .Z(n8610) );
  AND U11032 ( .A(n8611), .B(n8610), .Z(n8658) );
  NANDN U11033 ( .A(n8613), .B(n8612), .Z(n8617) );
  NAND U11034 ( .A(n8615), .B(n8614), .Z(n8616) );
  NAND U11035 ( .A(n8617), .B(n8616), .Z(n8740) );
  NAND U11036 ( .A(n8619), .B(n8618), .Z(n8623) );
  NAND U11037 ( .A(n8621), .B(n8620), .Z(n8622) );
  NAND U11038 ( .A(n8623), .B(n8622), .Z(n8738) );
  NAND U11039 ( .A(x[494]), .B(y[7749]), .Z(n8940) );
  NANDN U11040 ( .A(n8940), .B(n9167), .Z(n8627) );
  NAND U11041 ( .A(n8625), .B(n8624), .Z(n8626) );
  NAND U11042 ( .A(n8627), .B(n8626), .Z(n8732) );
  AND U11043 ( .A(x[489]), .B(y[7758]), .Z(n9545) );
  NANDN U11044 ( .A(n8718), .B(n9545), .Z(n8631) );
  NAND U11045 ( .A(n8629), .B(n8628), .Z(n8630) );
  NAND U11046 ( .A(n8631), .B(n8630), .Z(n8731) );
  XOR U11047 ( .A(n8732), .B(n8731), .Z(n8734) );
  AND U11048 ( .A(x[485]), .B(y[7756]), .Z(n8781) );
  NAND U11049 ( .A(y[7753]), .B(x[488]), .Z(n8632) );
  XNOR U11050 ( .A(n8781), .B(n8632), .Z(n8710) );
  XOR U11051 ( .A(n8726), .B(n8725), .Z(n8728) );
  NAND U11052 ( .A(y[7757]), .B(x[484]), .Z(n8633) );
  XNOR U11053 ( .A(n8634), .B(n8633), .Z(n8672) );
  AND U11054 ( .A(x[491]), .B(y[7750]), .Z(n8673) );
  XOR U11055 ( .A(n8672), .B(n8673), .Z(n8727) );
  XOR U11056 ( .A(n8728), .B(n8727), .Z(n8733) );
  XOR U11057 ( .A(n8734), .B(n8733), .Z(n8737) );
  XOR U11058 ( .A(n8738), .B(n8737), .Z(n8739) );
  XNOR U11059 ( .A(n8740), .B(n8739), .Z(n8656) );
  NAND U11060 ( .A(n8636), .B(n8635), .Z(n8640) );
  NAND U11061 ( .A(n8638), .B(n8637), .Z(n8639) );
  NAND U11062 ( .A(n8640), .B(n8639), .Z(n8655) );
  XOR U11063 ( .A(n8656), .B(n8655), .Z(n8657) );
  XOR U11064 ( .A(n8658), .B(n8657), .Z(n8756) );
  XOR U11065 ( .A(n8757), .B(n8756), .Z(n8758) );
  XOR U11066 ( .A(n8759), .B(n8758), .Z(n8752) );
  OR U11067 ( .A(n8643), .B(n8641), .Z(n8647) );
  ANDN U11068 ( .B(n8643), .A(n8642), .Z(n8645) );
  OR U11069 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U11070 ( .A(n8647), .B(n8646), .Z(n8751) );
  NANDN U11071 ( .A(n8649), .B(n8648), .Z(n8653) );
  NAND U11072 ( .A(n8651), .B(n8650), .Z(n8652) );
  NAND U11073 ( .A(n8653), .B(n8652), .Z(n8750) );
  IV U11074 ( .A(n8750), .Z(n8749) );
  XOR U11075 ( .A(n8751), .B(n8749), .Z(n8654) );
  XNOR U11076 ( .A(n8752), .B(n8654), .Z(N178) );
  NAND U11077 ( .A(n8656), .B(n8655), .Z(n8660) );
  NANDN U11078 ( .A(n8658), .B(n8657), .Z(n8659) );
  AND U11079 ( .A(n8660), .B(n8659), .Z(n8868) );
  NAND U11080 ( .A(n8662), .B(n8661), .Z(n8666) );
  NAND U11081 ( .A(n8664), .B(n8663), .Z(n8665) );
  AND U11082 ( .A(n8666), .B(n8665), .Z(n8866) );
  AND U11083 ( .A(x[495]), .B(y[7749]), .Z(n8913) );
  AND U11084 ( .A(x[492]), .B(y[7746]), .Z(n9022) );
  NAND U11085 ( .A(n8913), .B(n9022), .Z(n8670) );
  NANDN U11086 ( .A(n8668), .B(n8667), .Z(n8669) );
  NAND U11087 ( .A(n8670), .B(n8669), .Z(n8848) );
  NAND U11088 ( .A(n9945), .B(n8671), .Z(n8675) );
  NAND U11089 ( .A(n8673), .B(n8672), .Z(n8674) );
  NAND U11090 ( .A(n8675), .B(n8674), .Z(n8837) );
  AND U11091 ( .A(n8676), .B(o[81]), .Z(n8801) );
  AND U11092 ( .A(y[7761]), .B(x[481]), .Z(n8678) );
  XOR U11093 ( .A(n8678), .B(n8677), .Z(n8800) );
  XOR U11094 ( .A(n8801), .B(n8800), .Z(n8836) );
  AND U11095 ( .A(y[7747]), .B(x[495]), .Z(n8680) );
  NAND U11096 ( .A(y[7753]), .B(x[489]), .Z(n8679) );
  XNOR U11097 ( .A(n8680), .B(n8679), .Z(n8792) );
  AND U11098 ( .A(x[494]), .B(y[7748]), .Z(n8791) );
  XOR U11099 ( .A(n8792), .B(n8791), .Z(n8835) );
  XOR U11100 ( .A(n8836), .B(n8835), .Z(n8838) );
  XOR U11101 ( .A(n8837), .B(n8838), .Z(n8847) );
  XOR U11102 ( .A(n8848), .B(n8847), .Z(n8850) );
  NANDN U11103 ( .A(n8682), .B(n8681), .Z(n8686) );
  NAND U11104 ( .A(n8684), .B(n8683), .Z(n8685) );
  AND U11105 ( .A(n8686), .B(n8685), .Z(n8860) );
  AND U11106 ( .A(y[7746]), .B(x[496]), .Z(n8688) );
  NAND U11107 ( .A(y[7751]), .B(x[491]), .Z(n8687) );
  XNOR U11108 ( .A(n8688), .B(n8687), .Z(n8788) );
  AND U11109 ( .A(x[482]), .B(y[7760]), .Z(n8787) );
  XOR U11110 ( .A(n8788), .B(n8787), .Z(n8859) );
  AND U11111 ( .A(x[485]), .B(y[7757]), .Z(n8921) );
  NAND U11112 ( .A(y[7756]), .B(x[486]), .Z(n8689) );
  XNOR U11113 ( .A(n8921), .B(n8689), .Z(n8784) );
  NAND U11114 ( .A(y[7758]), .B(x[484]), .Z(n8690) );
  XNOR U11115 ( .A(n9548), .B(n8690), .Z(n8823) );
  AND U11116 ( .A(x[487]), .B(y[7755]), .Z(n8822) );
  XOR U11117 ( .A(n8823), .B(n8822), .Z(n8783) );
  XOR U11118 ( .A(n8784), .B(n8783), .Z(n8861) );
  XOR U11119 ( .A(n8862), .B(n8861), .Z(n8849) );
  XOR U11120 ( .A(n8850), .B(n8849), .Z(n8770) );
  NAND U11121 ( .A(n8692), .B(n8691), .Z(n8696) );
  NAND U11122 ( .A(n8694), .B(n8693), .Z(n8695) );
  AND U11123 ( .A(n8696), .B(n8695), .Z(n8841) );
  NAND U11124 ( .A(n8698), .B(n8697), .Z(n8702) );
  NAND U11125 ( .A(n8700), .B(n8699), .Z(n8701) );
  AND U11126 ( .A(n8702), .B(n8701), .Z(n8842) );
  XOR U11127 ( .A(n8841), .B(n8842), .Z(n8843) );
  NAND U11128 ( .A(n8704), .B(n8703), .Z(n8708) );
  NAND U11129 ( .A(n8706), .B(n8705), .Z(n8707) );
  AND U11130 ( .A(n8708), .B(n8707), .Z(n8844) );
  XOR U11131 ( .A(n8843), .B(n8844), .Z(n8769) );
  AND U11132 ( .A(x[488]), .B(y[7756]), .Z(n9062) );
  NAND U11133 ( .A(n9062), .B(n8709), .Z(n8713) );
  NANDN U11134 ( .A(n8711), .B(n8710), .Z(n8712) );
  NAND U11135 ( .A(n8713), .B(n8712), .Z(n8854) );
  NAND U11136 ( .A(x[489]), .B(y[7760]), .Z(n9686) );
  NANDN U11137 ( .A(n9686), .B(n8799), .Z(n8717) );
  NAND U11138 ( .A(n8715), .B(n8714), .Z(n8716) );
  NAND U11139 ( .A(n8717), .B(n8716), .Z(n8853) );
  XOR U11140 ( .A(n8854), .B(n8853), .Z(n8856) );
  AND U11141 ( .A(x[490]), .B(y[7759]), .Z(n9687) );
  NANDN U11142 ( .A(n8718), .B(n9687), .Z(n8722) );
  NANDN U11143 ( .A(n8720), .B(n8719), .Z(n8721) );
  NAND U11144 ( .A(n8722), .B(n8721), .Z(n8831) );
  AND U11145 ( .A(x[480]), .B(y[7762]), .Z(n8805) );
  AND U11146 ( .A(x[498]), .B(y[7744]), .Z(n8804) );
  XOR U11147 ( .A(n8805), .B(n8804), .Z(n8807) );
  AND U11148 ( .A(x[497]), .B(y[7745]), .Z(n8826) );
  XOR U11149 ( .A(n8826), .B(o[82]), .Z(n8806) );
  XOR U11150 ( .A(n8807), .B(n8806), .Z(n8830) );
  AND U11151 ( .A(y[7749]), .B(x[493]), .Z(n8724) );
  NAND U11152 ( .A(y[7759]), .B(x[483]), .Z(n8723) );
  XNOR U11153 ( .A(n8724), .B(n8723), .Z(n8813) );
  AND U11154 ( .A(x[492]), .B(y[7750]), .Z(n8812) );
  XOR U11155 ( .A(n8813), .B(n8812), .Z(n8829) );
  XOR U11156 ( .A(n8830), .B(n8829), .Z(n8832) );
  XOR U11157 ( .A(n8831), .B(n8832), .Z(n8855) );
  XNOR U11158 ( .A(n8856), .B(n8855), .Z(n8776) );
  NAND U11159 ( .A(n8726), .B(n8725), .Z(n8730) );
  NAND U11160 ( .A(n8728), .B(n8727), .Z(n8729) );
  AND U11161 ( .A(n8730), .B(n8729), .Z(n8775) );
  XOR U11162 ( .A(n8776), .B(n8775), .Z(n8777) );
  NAND U11163 ( .A(n8732), .B(n8731), .Z(n8736) );
  NAND U11164 ( .A(n8734), .B(n8733), .Z(n8735) );
  AND U11165 ( .A(n8736), .B(n8735), .Z(n8778) );
  XOR U11166 ( .A(n8777), .B(n8778), .Z(n8771) );
  XOR U11167 ( .A(n8772), .B(n8771), .Z(n8766) );
  NAND U11168 ( .A(n8738), .B(n8737), .Z(n8742) );
  NAND U11169 ( .A(n8740), .B(n8739), .Z(n8741) );
  AND U11170 ( .A(n8742), .B(n8741), .Z(n8764) );
  NAND U11171 ( .A(n8744), .B(n8743), .Z(n8748) );
  NANDN U11172 ( .A(n8746), .B(n8745), .Z(n8747) );
  NAND U11173 ( .A(n8748), .B(n8747), .Z(n8763) );
  XOR U11174 ( .A(n8866), .B(n8865), .Z(n8867) );
  XOR U11175 ( .A(n8868), .B(n8867), .Z(n8874) );
  OR U11176 ( .A(n8751), .B(n8749), .Z(n8755) );
  ANDN U11177 ( .B(n8751), .A(n8750), .Z(n8753) );
  OR U11178 ( .A(n8753), .B(n8752), .Z(n8754) );
  AND U11179 ( .A(n8755), .B(n8754), .Z(n8872) );
  NAND U11180 ( .A(n8757), .B(n8756), .Z(n8761) );
  NANDN U11181 ( .A(n8759), .B(n8758), .Z(n8760) );
  AND U11182 ( .A(n8761), .B(n8760), .Z(n8873) );
  IV U11183 ( .A(n8873), .Z(n8871) );
  XOR U11184 ( .A(n8872), .B(n8871), .Z(n8762) );
  XNOR U11185 ( .A(n8874), .B(n8762), .Z(N179) );
  NANDN U11186 ( .A(n8764), .B(n8763), .Z(n8768) );
  NANDN U11187 ( .A(n8766), .B(n8765), .Z(n8767) );
  AND U11188 ( .A(n8768), .B(n8767), .Z(n8882) );
  NANDN U11189 ( .A(n8770), .B(n8769), .Z(n8774) );
  NAND U11190 ( .A(n8772), .B(n8771), .Z(n8773) );
  AND U11191 ( .A(n8774), .B(n8773), .Z(n8880) );
  NAND U11192 ( .A(n8776), .B(n8775), .Z(n8780) );
  NAND U11193 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U11194 ( .A(n8780), .B(n8779), .Z(n8980) );
  AND U11195 ( .A(x[486]), .B(y[7757]), .Z(n8782) );
  NAND U11196 ( .A(n8782), .B(n8781), .Z(n8786) );
  NAND U11197 ( .A(n8784), .B(n8783), .Z(n8785) );
  NAND U11198 ( .A(n8786), .B(n8785), .Z(n8974) );
  AND U11199 ( .A(x[496]), .B(y[7751]), .Z(n9331) );
  NAND U11200 ( .A(n9331), .B(n9167), .Z(n8790) );
  NAND U11201 ( .A(n8788), .B(n8787), .Z(n8789) );
  NAND U11202 ( .A(n8790), .B(n8789), .Z(n8972) );
  AND U11203 ( .A(x[495]), .B(y[7753]), .Z(n9575) );
  NAND U11204 ( .A(n9575), .B(n8900), .Z(n8794) );
  NAND U11205 ( .A(n8792), .B(n8791), .Z(n8793) );
  NAND U11206 ( .A(n8794), .B(n8793), .Z(n8890) );
  AND U11207 ( .A(y[7762]), .B(x[481]), .Z(n8796) );
  NAND U11208 ( .A(y[7755]), .B(x[488]), .Z(n8795) );
  XNOR U11209 ( .A(n8796), .B(n8795), .Z(n8939) );
  AND U11210 ( .A(y[7750]), .B(x[493]), .Z(n8798) );
  NAND U11211 ( .A(y[7761]), .B(x[482]), .Z(n8797) );
  XNOR U11212 ( .A(n8798), .B(n8797), .Z(n8907) );
  XOR U11213 ( .A(n8907), .B(n8906), .Z(n8888) );
  XOR U11214 ( .A(n8889), .B(n8888), .Z(n8891) );
  XOR U11215 ( .A(n8890), .B(n8891), .Z(n8973) );
  XOR U11216 ( .A(n8972), .B(n8973), .Z(n8975) );
  XOR U11217 ( .A(n8974), .B(n8975), .Z(n8979) );
  NAND U11218 ( .A(x[490]), .B(y[7761]), .Z(n10025) );
  NANDN U11219 ( .A(n10025), .B(n8799), .Z(n8803) );
  NAND U11220 ( .A(n8801), .B(n8800), .Z(n8802) );
  NAND U11221 ( .A(n8803), .B(n8802), .Z(n8950) );
  NAND U11222 ( .A(n8805), .B(n8804), .Z(n8809) );
  NAND U11223 ( .A(n8807), .B(n8806), .Z(n8808) );
  NAND U11224 ( .A(n8809), .B(n8808), .Z(n8948) );
  AND U11225 ( .A(y[7747]), .B(x[496]), .Z(n9620) );
  NAND U11226 ( .A(y[7754]), .B(x[489]), .Z(n8810) );
  XNOR U11227 ( .A(n9620), .B(n8810), .Z(n8901) );
  NAND U11228 ( .A(x[495]), .B(y[7748]), .Z(n8902) );
  XOR U11229 ( .A(n8948), .B(n8949), .Z(n8951) );
  XOR U11230 ( .A(n8950), .B(n8951), .Z(n8969) );
  AND U11231 ( .A(x[493]), .B(y[7759]), .Z(n10231) );
  NAND U11232 ( .A(n8811), .B(n10231), .Z(n8815) );
  NAND U11233 ( .A(n8813), .B(n8812), .Z(n8814) );
  NAND U11234 ( .A(n8815), .B(n8814), .Z(n8956) );
  AND U11235 ( .A(y[7753]), .B(x[490]), .Z(n8817) );
  NAND U11236 ( .A(y[7746]), .B(x[497]), .Z(n8816) );
  XNOR U11237 ( .A(n8817), .B(n8816), .Z(n8945) );
  AND U11238 ( .A(x[498]), .B(y[7745]), .Z(n8920) );
  XOR U11239 ( .A(o[83]), .B(n8920), .Z(n8944) );
  XOR U11240 ( .A(n8945), .B(n8944), .Z(n8955) );
  NAND U11241 ( .A(y[7760]), .B(x[483]), .Z(n8818) );
  XNOR U11242 ( .A(n8819), .B(n8818), .Z(n8915) );
  XOR U11243 ( .A(n8915), .B(n8914), .Z(n8954) );
  XOR U11244 ( .A(n8955), .B(n8954), .Z(n8957) );
  XOR U11245 ( .A(n8956), .B(n8957), .Z(n8967) );
  NAND U11246 ( .A(n8821), .B(n8820), .Z(n8825) );
  NAND U11247 ( .A(n8823), .B(n8822), .Z(n8824) );
  NAND U11248 ( .A(n8825), .B(n8824), .Z(n8896) );
  AND U11249 ( .A(x[480]), .B(y[7763]), .Z(n8925) );
  NAND U11250 ( .A(x[499]), .B(y[7744]), .Z(n8926) );
  NAND U11251 ( .A(n8826), .B(o[82]), .Z(n8928) );
  AND U11252 ( .A(x[484]), .B(y[7759]), .Z(n9076) );
  AND U11253 ( .A(y[7758]), .B(x[485]), .Z(n8828) );
  NAND U11254 ( .A(y[7757]), .B(x[486]), .Z(n8827) );
  XOR U11255 ( .A(n8828), .B(n8827), .Z(n8922) );
  XOR U11256 ( .A(n8895), .B(n8894), .Z(n8897) );
  XNOR U11257 ( .A(n8896), .B(n8897), .Z(n8966) );
  NAND U11258 ( .A(n8830), .B(n8829), .Z(n8834) );
  NAND U11259 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U11260 ( .A(n8834), .B(n8833), .Z(n8961) );
  NAND U11261 ( .A(n8836), .B(n8835), .Z(n8840) );
  NAND U11262 ( .A(n8838), .B(n8837), .Z(n8839) );
  NAND U11263 ( .A(n8840), .B(n8839), .Z(n8960) );
  XOR U11264 ( .A(n8961), .B(n8960), .Z(n8962) );
  XNOR U11265 ( .A(n8963), .B(n8962), .Z(n8978) );
  XOR U11266 ( .A(n8980), .B(n8981), .Z(n8992) );
  NAND U11267 ( .A(n8842), .B(n8841), .Z(n8846) );
  NAND U11268 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U11269 ( .A(n8846), .B(n8845), .Z(n8991) );
  NAND U11270 ( .A(n8848), .B(n8847), .Z(n8852) );
  NAND U11271 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U11272 ( .A(n8852), .B(n8851), .Z(n8987) );
  NAND U11273 ( .A(n8854), .B(n8853), .Z(n8858) );
  NAND U11274 ( .A(n8856), .B(n8855), .Z(n8857) );
  AND U11275 ( .A(n8858), .B(n8857), .Z(n8985) );
  NANDN U11276 ( .A(n8860), .B(n8859), .Z(n8864) );
  NAND U11277 ( .A(n8862), .B(n8861), .Z(n8863) );
  NAND U11278 ( .A(n8864), .B(n8863), .Z(n8984) );
  XOR U11279 ( .A(n8991), .B(n8990), .Z(n8993) );
  XOR U11280 ( .A(n8992), .B(n8993), .Z(n8879) );
  XOR U11281 ( .A(n8880), .B(n8879), .Z(n8881) );
  XOR U11282 ( .A(n8882), .B(n8881), .Z(n8887) );
  NAND U11283 ( .A(n8866), .B(n8865), .Z(n8870) );
  NAND U11284 ( .A(n8868), .B(n8867), .Z(n8869) );
  NAND U11285 ( .A(n8870), .B(n8869), .Z(n8886) );
  NANDN U11286 ( .A(n8871), .B(n8872), .Z(n8877) );
  NOR U11287 ( .A(n8873), .B(n8872), .Z(n8875) );
  OR U11288 ( .A(n8875), .B(n8874), .Z(n8876) );
  AND U11289 ( .A(n8877), .B(n8876), .Z(n8885) );
  XOR U11290 ( .A(n8886), .B(n8885), .Z(n8878) );
  XNOR U11291 ( .A(n8887), .B(n8878), .Z(N180) );
  NAND U11292 ( .A(n8880), .B(n8879), .Z(n8884) );
  NANDN U11293 ( .A(n8882), .B(n8881), .Z(n8883) );
  NAND U11294 ( .A(n8884), .B(n8883), .Z(n9004) );
  IV U11295 ( .A(n9004), .Z(n9003) );
  NAND U11296 ( .A(n8889), .B(n8888), .Z(n8893) );
  NAND U11297 ( .A(n8891), .B(n8890), .Z(n8892) );
  NAND U11298 ( .A(n8893), .B(n8892), .Z(n9011) );
  NAND U11299 ( .A(n8895), .B(n8894), .Z(n8899) );
  NAND U11300 ( .A(n8897), .B(n8896), .Z(n8898) );
  NAND U11301 ( .A(n8899), .B(n8898), .Z(n9010) );
  XOR U11302 ( .A(n9011), .B(n9010), .Z(n9013) );
  AND U11303 ( .A(x[496]), .B(y[7754]), .Z(n9857) );
  NAND U11304 ( .A(n9857), .B(n8900), .Z(n8904) );
  NANDN U11305 ( .A(n8902), .B(n8901), .Z(n8903) );
  AND U11306 ( .A(n8904), .B(n8903), .Z(n9051) );
  AND U11307 ( .A(x[493]), .B(y[7761]), .Z(n10459) );
  NAND U11308 ( .A(n10459), .B(n8905), .Z(n8909) );
  NAND U11309 ( .A(n8907), .B(n8906), .Z(n8908) );
  AND U11310 ( .A(n8909), .B(n8908), .Z(n9096) );
  AND U11311 ( .A(y[7748]), .B(x[496]), .Z(n8911) );
  NAND U11312 ( .A(y[7754]), .B(x[490]), .Z(n8910) );
  XNOR U11313 ( .A(n8911), .B(n8910), .Z(n9057) );
  NAND U11314 ( .A(x[482]), .B(y[7762]), .Z(n9058) );
  NAND U11315 ( .A(y[7755]), .B(x[489]), .Z(n8912) );
  XNOR U11316 ( .A(n8913), .B(n8912), .Z(n9033) );
  AND U11317 ( .A(x[494]), .B(y[7750]), .Z(n9034) );
  XOR U11318 ( .A(n9033), .B(n9034), .Z(n9093) );
  XOR U11319 ( .A(n9094), .B(n9093), .Z(n9095) );
  NAND U11320 ( .A(x[491]), .B(y[7760]), .Z(n10026) );
  NANDN U11321 ( .A(n10026), .B(n9194), .Z(n8917) );
  NAND U11322 ( .A(n8915), .B(n8914), .Z(n8916) );
  AND U11323 ( .A(n8917), .B(n8916), .Z(n9102) );
  AND U11324 ( .A(y[7753]), .B(x[491]), .Z(n8919) );
  NAND U11325 ( .A(y[7763]), .B(x[481]), .Z(n8918) );
  XNOR U11326 ( .A(n8919), .B(n8918), .Z(n9029) );
  AND U11327 ( .A(x[499]), .B(y[7745]), .Z(n9037) );
  XOR U11328 ( .A(o[84]), .B(n9037), .Z(n9028) );
  XOR U11329 ( .A(n9029), .B(n9028), .Z(n9100) );
  AND U11330 ( .A(x[480]), .B(y[7764]), .Z(n9081) );
  AND U11331 ( .A(x[500]), .B(y[7744]), .Z(n9082) );
  XOR U11332 ( .A(n9081), .B(n9082), .Z(n9084) );
  AND U11333 ( .A(o[83]), .B(n8920), .Z(n9083) );
  XOR U11334 ( .A(n9084), .B(n9083), .Z(n9099) );
  XOR U11335 ( .A(n9100), .B(n9099), .Z(n9101) );
  XOR U11336 ( .A(n9053), .B(n9052), .Z(n9012) );
  XOR U11337 ( .A(n9013), .B(n9012), .Z(n9108) );
  AND U11338 ( .A(x[486]), .B(y[7758]), .Z(n9017) );
  IV U11339 ( .A(n9017), .Z(n8937) );
  NANDN U11340 ( .A(n8937), .B(n8921), .Z(n8924) );
  NANDN U11341 ( .A(n8922), .B(n9076), .Z(n8923) );
  AND U11342 ( .A(n8924), .B(n8923), .Z(n9041) );
  NANDN U11343 ( .A(n8926), .B(n8925), .Z(n8930) );
  NANDN U11344 ( .A(n8928), .B(n8927), .Z(n8929) );
  AND U11345 ( .A(n8930), .B(n8929), .Z(n9039) );
  AND U11346 ( .A(y[7746]), .B(x[498]), .Z(n8932) );
  NAND U11347 ( .A(y[7752]), .B(x[492]), .Z(n8931) );
  XNOR U11348 ( .A(n8932), .B(n8931), .Z(n9023) );
  AND U11349 ( .A(x[497]), .B(y[7747]), .Z(n9024) );
  XOR U11350 ( .A(n9023), .B(n9024), .Z(n9038) );
  AND U11351 ( .A(y[7751]), .B(x[493]), .Z(n8934) );
  NAND U11352 ( .A(y[7761]), .B(x[483]), .Z(n8933) );
  XNOR U11353 ( .A(n8934), .B(n8933), .Z(n9063) );
  XOR U11354 ( .A(n9063), .B(n9062), .Z(n9019) );
  AND U11355 ( .A(y[7759]), .B(x[485]), .Z(n8936) );
  NAND U11356 ( .A(y[7760]), .B(x[484]), .Z(n8935) );
  XNOR U11357 ( .A(n8936), .B(n8935), .Z(n9078) );
  AND U11358 ( .A(x[487]), .B(y[7757]), .Z(n9077) );
  XNOR U11359 ( .A(n9078), .B(n9077), .Z(n9016) );
  XOR U11360 ( .A(n8937), .B(n9016), .Z(n9018) );
  AND U11361 ( .A(x[488]), .B(y[7762]), .Z(n10183) );
  AND U11362 ( .A(x[481]), .B(y[7755]), .Z(n8938) );
  NAND U11363 ( .A(n10183), .B(n8938), .Z(n8942) );
  NANDN U11364 ( .A(n8940), .B(n8939), .Z(n8941) );
  AND U11365 ( .A(n8942), .B(n8941), .Z(n9088) );
  AND U11366 ( .A(x[497]), .B(y[7753]), .Z(n9865) );
  NAND U11367 ( .A(n9865), .B(n8943), .Z(n8947) );
  NAND U11368 ( .A(n8945), .B(n8944), .Z(n8946) );
  NAND U11369 ( .A(n8947), .B(n8946), .Z(n9087) );
  XNOR U11370 ( .A(n9089), .B(n9090), .Z(n9044) );
  NAND U11371 ( .A(n8949), .B(n8948), .Z(n8953) );
  NAND U11372 ( .A(n8951), .B(n8950), .Z(n8952) );
  AND U11373 ( .A(n8953), .B(n8952), .Z(n9046) );
  XOR U11374 ( .A(n9047), .B(n9046), .Z(n9106) );
  NAND U11375 ( .A(n8955), .B(n8954), .Z(n8959) );
  NAND U11376 ( .A(n8957), .B(n8956), .Z(n8958) );
  AND U11377 ( .A(n8959), .B(n8958), .Z(n9105) );
  XOR U11378 ( .A(n9106), .B(n9105), .Z(n9107) );
  NAND U11379 ( .A(n8961), .B(n8960), .Z(n8965) );
  NAND U11380 ( .A(n8963), .B(n8962), .Z(n8964) );
  AND U11381 ( .A(n8965), .B(n8964), .Z(n9120) );
  NANDN U11382 ( .A(n8967), .B(n8966), .Z(n8971) );
  NANDN U11383 ( .A(n8969), .B(n8968), .Z(n8970) );
  NAND U11384 ( .A(n8971), .B(n8970), .Z(n9117) );
  NAND U11385 ( .A(n8973), .B(n8972), .Z(n8977) );
  NAND U11386 ( .A(n8975), .B(n8974), .Z(n8976) );
  AND U11387 ( .A(n8977), .B(n8976), .Z(n9118) );
  XOR U11388 ( .A(n9117), .B(n9118), .Z(n9119) );
  XNOR U11389 ( .A(n9120), .B(n9119), .Z(n9111) );
  NANDN U11390 ( .A(n8979), .B(n8978), .Z(n8983) );
  NANDN U11391 ( .A(n8981), .B(n8980), .Z(n8982) );
  AND U11392 ( .A(n8983), .B(n8982), .Z(n9113) );
  XNOR U11393 ( .A(n9114), .B(n9113), .Z(n9000) );
  NANDN U11394 ( .A(n8985), .B(n8984), .Z(n8989) );
  NANDN U11395 ( .A(n8987), .B(n8986), .Z(n8988) );
  AND U11396 ( .A(n8989), .B(n8988), .Z(n8997) );
  NAND U11397 ( .A(n8991), .B(n8990), .Z(n8995) );
  NAND U11398 ( .A(n8993), .B(n8992), .Z(n8994) );
  AND U11399 ( .A(n8995), .B(n8994), .Z(n8998) );
  XOR U11400 ( .A(n8997), .B(n8998), .Z(n8999) );
  XOR U11401 ( .A(n9000), .B(n8999), .Z(n9006) );
  XNOR U11402 ( .A(n9005), .B(n9006), .Z(n8996) );
  XOR U11403 ( .A(n9003), .B(n8996), .Z(N181) );
  NAND U11404 ( .A(n8998), .B(n8997), .Z(n9002) );
  NAND U11405 ( .A(n9000), .B(n8999), .Z(n9001) );
  NAND U11406 ( .A(n9002), .B(n9001), .Z(n9132) );
  IV U11407 ( .A(n9132), .Z(n9130) );
  OR U11408 ( .A(n9005), .B(n9003), .Z(n9009) );
  ANDN U11409 ( .B(n9005), .A(n9004), .Z(n9007) );
  OR U11410 ( .A(n9007), .B(n9006), .Z(n9008) );
  AND U11411 ( .A(n9009), .B(n9008), .Z(n9131) );
  NAND U11412 ( .A(n9011), .B(n9010), .Z(n9015) );
  NAND U11413 ( .A(n9013), .B(n9012), .Z(n9014) );
  NAND U11414 ( .A(n9015), .B(n9014), .Z(n9145) );
  NANDN U11415 ( .A(n9017), .B(n9016), .Z(n9021) );
  NANDN U11416 ( .A(n9019), .B(n9018), .Z(n9020) );
  AND U11417 ( .A(n9021), .B(n9020), .Z(n9235) );
  AND U11418 ( .A(x[498]), .B(y[7752]), .Z(n9864) );
  NAND U11419 ( .A(n9864), .B(n9022), .Z(n9026) );
  NAND U11420 ( .A(n9024), .B(n9023), .Z(n9025) );
  NAND U11421 ( .A(n9026), .B(n9025), .Z(n9217) );
  AND U11422 ( .A(x[491]), .B(y[7763]), .Z(n10524) );
  AND U11423 ( .A(x[481]), .B(y[7753]), .Z(n9027) );
  NAND U11424 ( .A(n10524), .B(n9027), .Z(n9031) );
  NAND U11425 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U11426 ( .A(n9031), .B(n9030), .Z(n9216) );
  XOR U11427 ( .A(n9217), .B(n9216), .Z(n9219) );
  AND U11428 ( .A(x[495]), .B(y[7755]), .Z(n9852) );
  NAND U11429 ( .A(n9852), .B(n9032), .Z(n9036) );
  NAND U11430 ( .A(n9034), .B(n9033), .Z(n9035) );
  NAND U11431 ( .A(n9036), .B(n9035), .Z(n9181) );
  AND U11432 ( .A(x[480]), .B(y[7765]), .Z(n9200) );
  AND U11433 ( .A(x[501]), .B(y[7744]), .Z(n9201) );
  XOR U11434 ( .A(n9200), .B(n9201), .Z(n9203) );
  AND U11435 ( .A(o[84]), .B(n9037), .Z(n9202) );
  XOR U11436 ( .A(n9203), .B(n9202), .Z(n9179) );
  AND U11437 ( .A(x[485]), .B(y[7760]), .Z(n9187) );
  AND U11438 ( .A(x[496]), .B(y[7749]), .Z(n9186) );
  XOR U11439 ( .A(n9187), .B(n9186), .Z(n9185) );
  AND U11440 ( .A(x[495]), .B(y[7750]), .Z(n9184) );
  XOR U11441 ( .A(n9185), .B(n9184), .Z(n9178) );
  XOR U11442 ( .A(n9179), .B(n9178), .Z(n9180) );
  XOR U11443 ( .A(n9181), .B(n9180), .Z(n9218) );
  XNOR U11444 ( .A(n9219), .B(n9218), .Z(n9234) );
  NANDN U11445 ( .A(n9039), .B(n9038), .Z(n9043) );
  NANDN U11446 ( .A(n9041), .B(n9040), .Z(n9042) );
  NAND U11447 ( .A(n9043), .B(n9042), .Z(n9237) );
  NANDN U11448 ( .A(n9045), .B(n9044), .Z(n9049) );
  NAND U11449 ( .A(n9047), .B(n9046), .Z(n9048) );
  AND U11450 ( .A(n9049), .B(n9048), .Z(n9143) );
  XOR U11451 ( .A(n9145), .B(n9146), .Z(n9140) );
  NANDN U11452 ( .A(n9051), .B(n9050), .Z(n9055) );
  NAND U11453 ( .A(n9053), .B(n9052), .Z(n9054) );
  AND U11454 ( .A(n9055), .B(n9054), .Z(n9243) );
  NAND U11455 ( .A(n9857), .B(n9056), .Z(n9060) );
  NANDN U11456 ( .A(n9058), .B(n9057), .Z(n9059) );
  AND U11457 ( .A(n9060), .B(n9059), .Z(n9150) );
  NAND U11458 ( .A(n10459), .B(n9061), .Z(n9065) );
  NAND U11459 ( .A(n9063), .B(n9062), .Z(n9064) );
  NAND U11460 ( .A(n9065), .B(n9064), .Z(n9231) );
  AND U11461 ( .A(y[7746]), .B(x[499]), .Z(n9067) );
  NAND U11462 ( .A(y[7754]), .B(x[491]), .Z(n9066) );
  XNOR U11463 ( .A(n9067), .B(n9066), .Z(n9169) );
  AND U11464 ( .A(x[500]), .B(y[7745]), .Z(n9199) );
  XOR U11465 ( .A(o[85]), .B(n9199), .Z(n9168) );
  XOR U11466 ( .A(n9169), .B(n9168), .Z(n9229) );
  AND U11467 ( .A(y[7747]), .B(x[498]), .Z(n9069) );
  NAND U11468 ( .A(y[7755]), .B(x[490]), .Z(n9068) );
  XNOR U11469 ( .A(n9069), .B(n9068), .Z(n9207) );
  AND U11470 ( .A(x[481]), .B(y[7764]), .Z(n9208) );
  XOR U11471 ( .A(n9207), .B(n9208), .Z(n9228) );
  XOR U11472 ( .A(n9229), .B(n9228), .Z(n9230) );
  XOR U11473 ( .A(n9231), .B(n9230), .Z(n9149) );
  AND U11474 ( .A(x[487]), .B(y[7758]), .Z(n9463) );
  AND U11475 ( .A(y[7759]), .B(x[486]), .Z(n9071) );
  NAND U11476 ( .A(y[7751]), .B(x[494]), .Z(n9070) );
  XNOR U11477 ( .A(n9071), .B(n9070), .Z(n9211) );
  XNOR U11478 ( .A(n9463), .B(n9211), .Z(n9158) );
  NAND U11479 ( .A(x[489]), .B(y[7756]), .Z(n9156) );
  NAND U11480 ( .A(x[488]), .B(y[7757]), .Z(n9155) );
  XOR U11481 ( .A(n9156), .B(n9155), .Z(n9157) );
  XNOR U11482 ( .A(n9158), .B(n9157), .Z(n9174) );
  AND U11483 ( .A(y[7753]), .B(x[492]), .Z(n9073) );
  NAND U11484 ( .A(y[7748]), .B(x[497]), .Z(n9072) );
  XNOR U11485 ( .A(n9073), .B(n9072), .Z(n9161) );
  AND U11486 ( .A(x[482]), .B(y[7763]), .Z(n9162) );
  XOR U11487 ( .A(n9161), .B(n9162), .Z(n9173) );
  AND U11488 ( .A(y[7752]), .B(x[493]), .Z(n9075) );
  NAND U11489 ( .A(y[7762]), .B(x[483]), .Z(n9074) );
  XNOR U11490 ( .A(n9075), .B(n9074), .Z(n9195) );
  AND U11491 ( .A(x[484]), .B(y[7761]), .Z(n9196) );
  XOR U11492 ( .A(n9195), .B(n9196), .Z(n9172) );
  XOR U11493 ( .A(n9173), .B(n9172), .Z(n9175) );
  XOR U11494 ( .A(n9174), .B(n9175), .Z(n9225) );
  NAND U11495 ( .A(n9187), .B(n9076), .Z(n9080) );
  NAND U11496 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U11497 ( .A(n9080), .B(n9079), .Z(n9223) );
  NAND U11498 ( .A(n9082), .B(n9081), .Z(n9086) );
  NAND U11499 ( .A(n9084), .B(n9083), .Z(n9085) );
  NAND U11500 ( .A(n9086), .B(n9085), .Z(n9222) );
  XOR U11501 ( .A(n9223), .B(n9222), .Z(n9224) );
  XOR U11502 ( .A(n9225), .B(n9224), .Z(n9151) );
  XOR U11503 ( .A(n9152), .B(n9151), .Z(n9241) );
  NANDN U11504 ( .A(n9088), .B(n9087), .Z(n9092) );
  NAND U11505 ( .A(n9090), .B(n9089), .Z(n9091) );
  NAND U11506 ( .A(n9092), .B(n9091), .Z(n9248) );
  NAND U11507 ( .A(n9094), .B(n9093), .Z(n9098) );
  NANDN U11508 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U11509 ( .A(n9098), .B(n9097), .Z(n9247) );
  NAND U11510 ( .A(n9100), .B(n9099), .Z(n9104) );
  NANDN U11511 ( .A(n9102), .B(n9101), .Z(n9103) );
  NAND U11512 ( .A(n9104), .B(n9103), .Z(n9246) );
  XOR U11513 ( .A(n9247), .B(n9246), .Z(n9249) );
  XOR U11514 ( .A(n9248), .B(n9249), .Z(n9240) );
  XOR U11515 ( .A(n9241), .B(n9240), .Z(n9242) );
  NAND U11516 ( .A(n9106), .B(n9105), .Z(n9110) );
  NANDN U11517 ( .A(n9108), .B(n9107), .Z(n9109) );
  NAND U11518 ( .A(n9110), .B(n9109), .Z(n9137) );
  NANDN U11519 ( .A(n9112), .B(n9111), .Z(n9116) );
  NAND U11520 ( .A(n9114), .B(n9113), .Z(n9115) );
  NAND U11521 ( .A(n9116), .B(n9115), .Z(n9124) );
  NAND U11522 ( .A(n9118), .B(n9117), .Z(n9122) );
  NAND U11523 ( .A(n9120), .B(n9119), .Z(n9121) );
  AND U11524 ( .A(n9122), .B(n9121), .Z(n9125) );
  XOR U11525 ( .A(n9124), .B(n9125), .Z(n9126) );
  XNOR U11526 ( .A(n9131), .B(n9133), .Z(n9123) );
  XOR U11527 ( .A(n9130), .B(n9123), .Z(N182) );
  NAND U11528 ( .A(n9125), .B(n9124), .Z(n9129) );
  NANDN U11529 ( .A(n9127), .B(n9126), .Z(n9128) );
  AND U11530 ( .A(n9129), .B(n9128), .Z(n9373) );
  NANDN U11531 ( .A(n9130), .B(n9131), .Z(n9136) );
  NOR U11532 ( .A(n9132), .B(n9131), .Z(n9134) );
  OR U11533 ( .A(n9134), .B(n9133), .Z(n9135) );
  AND U11534 ( .A(n9136), .B(n9135), .Z(n9374) );
  NANDN U11535 ( .A(n9138), .B(n9137), .Z(n9142) );
  NANDN U11536 ( .A(n9140), .B(n9139), .Z(n9141) );
  AND U11537 ( .A(n9142), .B(n9141), .Z(n9378) );
  NANDN U11538 ( .A(n9144), .B(n9143), .Z(n9148) );
  NAND U11539 ( .A(n9146), .B(n9145), .Z(n9147) );
  NAND U11540 ( .A(n9148), .B(n9147), .Z(n9376) );
  NANDN U11541 ( .A(n9150), .B(n9149), .Z(n9154) );
  NAND U11542 ( .A(n9152), .B(n9151), .Z(n9153) );
  AND U11543 ( .A(n9154), .B(n9153), .Z(n9370) );
  NAND U11544 ( .A(n9156), .B(n9155), .Z(n9160) );
  NAND U11545 ( .A(n9158), .B(n9157), .Z(n9159) );
  NAND U11546 ( .A(n9160), .B(n9159), .Z(n9364) );
  NAND U11547 ( .A(n9865), .B(n9315), .Z(n9164) );
  NAND U11548 ( .A(n9162), .B(n9161), .Z(n9163) );
  NAND U11549 ( .A(n9164), .B(n9163), .Z(n9291) );
  AND U11550 ( .A(x[485]), .B(y[7761]), .Z(n9337) );
  AND U11551 ( .A(x[497]), .B(y[7749]), .Z(n9338) );
  XOR U11552 ( .A(n9337), .B(n9338), .Z(n9339) );
  AND U11553 ( .A(x[496]), .B(y[7750]), .Z(n9340) );
  XOR U11554 ( .A(n9339), .B(n9340), .Z(n9290) );
  AND U11555 ( .A(y[7748]), .B(x[498]), .Z(n9166) );
  NAND U11556 ( .A(y[7754]), .B(x[492]), .Z(n9165) );
  XNOR U11557 ( .A(n9166), .B(n9165), .Z(n9316) );
  AND U11558 ( .A(x[484]), .B(y[7762]), .Z(n9317) );
  XOR U11559 ( .A(n9316), .B(n9317), .Z(n9289) );
  XOR U11560 ( .A(n9290), .B(n9289), .Z(n9292) );
  XNOR U11561 ( .A(n9291), .B(n9292), .Z(n9361) );
  AND U11562 ( .A(x[499]), .B(y[7754]), .Z(n10344) );
  NAND U11563 ( .A(n10344), .B(n9167), .Z(n9171) );
  NAND U11564 ( .A(n9169), .B(n9168), .Z(n9170) );
  AND U11565 ( .A(n9171), .B(n9170), .Z(n9362) );
  XOR U11566 ( .A(n9361), .B(n9362), .Z(n9363) );
  XNOR U11567 ( .A(n9364), .B(n9363), .Z(n9367) );
  NAND U11568 ( .A(n9173), .B(n9172), .Z(n9177) );
  NAND U11569 ( .A(n9175), .B(n9174), .Z(n9176) );
  NAND U11570 ( .A(n9177), .B(n9176), .Z(n9350) );
  NAND U11571 ( .A(n9179), .B(n9178), .Z(n9183) );
  NAND U11572 ( .A(n9181), .B(n9180), .Z(n9182) );
  NAND U11573 ( .A(n9183), .B(n9182), .Z(n9349) );
  XOR U11574 ( .A(n9350), .B(n9349), .Z(n9352) );
  AND U11575 ( .A(n9185), .B(n9184), .Z(n9189) );
  NAND U11576 ( .A(n9187), .B(n9186), .Z(n9188) );
  NANDN U11577 ( .A(n9189), .B(n9188), .Z(n9312) );
  AND U11578 ( .A(y[7753]), .B(x[493]), .Z(n9191) );
  NAND U11579 ( .A(y[7746]), .B(x[500]), .Z(n9190) );
  XNOR U11580 ( .A(n9191), .B(n9190), .Z(n9333) );
  AND U11581 ( .A(x[482]), .B(y[7764]), .Z(n9334) );
  XOR U11582 ( .A(n9333), .B(n9334), .Z(n9310) );
  AND U11583 ( .A(y[7760]), .B(x[486]), .Z(n9193) );
  NAND U11584 ( .A(y[7751]), .B(x[495]), .Z(n9192) );
  XNOR U11585 ( .A(n9193), .B(n9192), .Z(n9345) );
  XOR U11586 ( .A(n9310), .B(n9309), .Z(n9311) );
  XOR U11587 ( .A(n9312), .B(n9311), .Z(n9356) );
  AND U11588 ( .A(x[493]), .B(y[7762]), .Z(n10591) );
  NAND U11589 ( .A(n9194), .B(n10591), .Z(n9198) );
  NAND U11590 ( .A(n9196), .B(n9195), .Z(n9197) );
  NAND U11591 ( .A(n9198), .B(n9197), .Z(n9280) );
  AND U11592 ( .A(x[481]), .B(y[7765]), .Z(n9303) );
  XOR U11593 ( .A(n9304), .B(n9303), .Z(n9302) );
  AND U11594 ( .A(o[85]), .B(n9199), .Z(n9301) );
  XOR U11595 ( .A(n9302), .B(n9301), .Z(n9278) );
  AND U11596 ( .A(x[494]), .B(y[7752]), .Z(n9295) );
  AND U11597 ( .A(x[483]), .B(y[7763]), .Z(n9296) );
  XOR U11598 ( .A(n9295), .B(n9296), .Z(n9297) );
  AND U11599 ( .A(x[499]), .B(y[7747]), .Z(n9298) );
  XOR U11600 ( .A(n9297), .B(n9298), .Z(n9277) );
  XOR U11601 ( .A(n9278), .B(n9277), .Z(n9279) );
  XOR U11602 ( .A(n9280), .B(n9279), .Z(n9355) );
  XOR U11603 ( .A(n9356), .B(n9355), .Z(n9358) );
  NAND U11604 ( .A(n9201), .B(n9200), .Z(n9205) );
  NAND U11605 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U11606 ( .A(n9205), .B(n9204), .Z(n9272) );
  AND U11607 ( .A(x[498]), .B(y[7755]), .Z(n10347) );
  NAND U11608 ( .A(n10347), .B(n9206), .Z(n9210) );
  NAND U11609 ( .A(n9208), .B(n9207), .Z(n9209) );
  NAND U11610 ( .A(n9210), .B(n9209), .Z(n9271) );
  XOR U11611 ( .A(n9272), .B(n9271), .Z(n9274) );
  AND U11612 ( .A(x[494]), .B(y[7759]), .Z(n10357) );
  NAND U11613 ( .A(n10357), .B(n9344), .Z(n9213) );
  NAND U11614 ( .A(n9463), .B(n9211), .Z(n9212) );
  NAND U11615 ( .A(n9213), .B(n9212), .Z(n9286) );
  AND U11616 ( .A(x[480]), .B(y[7766]), .Z(n9320) );
  AND U11617 ( .A(x[502]), .B(y[7744]), .Z(n9321) );
  XOR U11618 ( .A(n9320), .B(n9321), .Z(n9323) );
  AND U11619 ( .A(x[501]), .B(y[7745]), .Z(n9343) );
  XOR U11620 ( .A(o[86]), .B(n9343), .Z(n9322) );
  XOR U11621 ( .A(n9323), .B(n9322), .Z(n9284) );
  AND U11622 ( .A(y[7759]), .B(x[487]), .Z(n9215) );
  NAND U11623 ( .A(y[7758]), .B(x[488]), .Z(n9214) );
  XNOR U11624 ( .A(n9215), .B(n9214), .Z(n9326) );
  XOR U11625 ( .A(n9284), .B(n9283), .Z(n9285) );
  XOR U11626 ( .A(n9286), .B(n9285), .Z(n9273) );
  XOR U11627 ( .A(n9274), .B(n9273), .Z(n9357) );
  XOR U11628 ( .A(n9358), .B(n9357), .Z(n9351) );
  XOR U11629 ( .A(n9352), .B(n9351), .Z(n9368) );
  XOR U11630 ( .A(n9367), .B(n9368), .Z(n9369) );
  NAND U11631 ( .A(n9217), .B(n9216), .Z(n9221) );
  NAND U11632 ( .A(n9219), .B(n9218), .Z(n9220) );
  NAND U11633 ( .A(n9221), .B(n9220), .Z(n9268) );
  NAND U11634 ( .A(n9223), .B(n9222), .Z(n9227) );
  NAND U11635 ( .A(n9225), .B(n9224), .Z(n9226) );
  NAND U11636 ( .A(n9227), .B(n9226), .Z(n9266) );
  NAND U11637 ( .A(n9229), .B(n9228), .Z(n9233) );
  NAND U11638 ( .A(n9231), .B(n9230), .Z(n9232) );
  NAND U11639 ( .A(n9233), .B(n9232), .Z(n9265) );
  XOR U11640 ( .A(n9266), .B(n9265), .Z(n9267) );
  XNOR U11641 ( .A(n9268), .B(n9267), .Z(n9260) );
  NANDN U11642 ( .A(n9235), .B(n9234), .Z(n9239) );
  NANDN U11643 ( .A(n9237), .B(n9236), .Z(n9238) );
  NAND U11644 ( .A(n9239), .B(n9238), .Z(n9259) );
  XOR U11645 ( .A(n9260), .B(n9259), .Z(n9262) );
  XNOR U11646 ( .A(n9261), .B(n9262), .Z(n9255) );
  NAND U11647 ( .A(n9241), .B(n9240), .Z(n9245) );
  NANDN U11648 ( .A(n9243), .B(n9242), .Z(n9244) );
  AND U11649 ( .A(n9245), .B(n9244), .Z(n9254) );
  NAND U11650 ( .A(n9247), .B(n9246), .Z(n9251) );
  NAND U11651 ( .A(n9249), .B(n9248), .Z(n9250) );
  NAND U11652 ( .A(n9251), .B(n9250), .Z(n9253) );
  XNOR U11653 ( .A(n9255), .B(n9256), .Z(n9377) );
  XNOR U11654 ( .A(n9378), .B(n9379), .Z(n9375) );
  XNOR U11655 ( .A(n9374), .B(n9375), .Z(n9252) );
  XOR U11656 ( .A(n9373), .B(n9252), .Z(N183) );
  NANDN U11657 ( .A(n9254), .B(n9253), .Z(n9258) );
  NAND U11658 ( .A(n9256), .B(n9255), .Z(n9257) );
  AND U11659 ( .A(n9258), .B(n9257), .Z(n9517) );
  NAND U11660 ( .A(n9260), .B(n9259), .Z(n9264) );
  NAND U11661 ( .A(n9262), .B(n9261), .Z(n9263) );
  AND U11662 ( .A(n9264), .B(n9263), .Z(n9515) );
  NAND U11663 ( .A(n9266), .B(n9265), .Z(n9270) );
  NAND U11664 ( .A(n9268), .B(n9267), .Z(n9269) );
  NAND U11665 ( .A(n9270), .B(n9269), .Z(n9499) );
  NAND U11666 ( .A(n9272), .B(n9271), .Z(n9276) );
  NAND U11667 ( .A(n9274), .B(n9273), .Z(n9275) );
  NAND U11668 ( .A(n9276), .B(n9275), .Z(n9446) );
  NAND U11669 ( .A(n9278), .B(n9277), .Z(n9282) );
  NAND U11670 ( .A(n9280), .B(n9279), .Z(n9281) );
  NAND U11671 ( .A(n9282), .B(n9281), .Z(n9444) );
  NAND U11672 ( .A(n9284), .B(n9283), .Z(n9288) );
  NAND U11673 ( .A(n9286), .B(n9285), .Z(n9287) );
  NAND U11674 ( .A(n9288), .B(n9287), .Z(n9443) );
  XOR U11675 ( .A(n9444), .B(n9443), .Z(n9445) );
  XOR U11676 ( .A(n9446), .B(n9445), .Z(n9511) );
  NAND U11677 ( .A(n9290), .B(n9289), .Z(n9294) );
  NAND U11678 ( .A(n9292), .B(n9291), .Z(n9293) );
  NAND U11679 ( .A(n9294), .B(n9293), .Z(n9509) );
  NAND U11680 ( .A(n9296), .B(n9295), .Z(n9300) );
  NAND U11681 ( .A(n9298), .B(n9297), .Z(n9299) );
  NAND U11682 ( .A(n9300), .B(n9299), .Z(n9390) );
  AND U11683 ( .A(n9302), .B(n9301), .Z(n9306) );
  NAND U11684 ( .A(n9304), .B(n9303), .Z(n9305) );
  NANDN U11685 ( .A(n9306), .B(n9305), .Z(n9389) );
  XOR U11686 ( .A(n9390), .B(n9389), .Z(n9392) );
  AND U11687 ( .A(y[7760]), .B(x[487]), .Z(n9308) );
  NAND U11688 ( .A(y[7758]), .B(x[489]), .Z(n9307) );
  XNOR U11689 ( .A(n9308), .B(n9307), .Z(n9464) );
  AND U11690 ( .A(x[490]), .B(y[7757]), .Z(n9396) );
  XOR U11691 ( .A(n9395), .B(n9396), .Z(n9398) );
  AND U11692 ( .A(x[486]), .B(y[7761]), .Z(n9455) );
  AND U11693 ( .A(x[495]), .B(y[7752]), .Z(n9456) );
  XOR U11694 ( .A(n9455), .B(n9456), .Z(n9457) );
  AND U11695 ( .A(x[491]), .B(y[7756]), .Z(n9458) );
  XOR U11696 ( .A(n9457), .B(n9458), .Z(n9397) );
  XOR U11697 ( .A(n9398), .B(n9397), .Z(n9391) );
  XOR U11698 ( .A(n9392), .B(n9391), .Z(n9508) );
  XOR U11699 ( .A(n9509), .B(n9508), .Z(n9510) );
  XOR U11700 ( .A(n9511), .B(n9510), .Z(n9497) );
  NAND U11701 ( .A(n9310), .B(n9309), .Z(n9314) );
  NAND U11702 ( .A(n9312), .B(n9311), .Z(n9313) );
  NAND U11703 ( .A(n9314), .B(n9313), .Z(n9491) );
  AND U11704 ( .A(x[498]), .B(y[7754]), .Z(n10213) );
  NAND U11705 ( .A(n10213), .B(n9315), .Z(n9319) );
  NAND U11706 ( .A(n9317), .B(n9316), .Z(n9318) );
  NAND U11707 ( .A(n9319), .B(n9318), .Z(n9432) );
  NAND U11708 ( .A(n9321), .B(n9320), .Z(n9325) );
  NAND U11709 ( .A(n9323), .B(n9322), .Z(n9324) );
  NAND U11710 ( .A(n9325), .B(n9324), .Z(n9431) );
  XOR U11711 ( .A(n9432), .B(n9431), .Z(n9433) );
  NANDN U11712 ( .A(n9465), .B(n9463), .Z(n9329) );
  NANDN U11713 ( .A(n9327), .B(n9326), .Z(n9328) );
  NAND U11714 ( .A(n9329), .B(n9328), .Z(n9427) );
  AND U11715 ( .A(x[480]), .B(y[7767]), .Z(n9474) );
  AND U11716 ( .A(x[503]), .B(y[7744]), .Z(n9475) );
  XOR U11717 ( .A(n9474), .B(n9475), .Z(n9477) );
  AND U11718 ( .A(x[502]), .B(y[7745]), .Z(n9454) );
  XOR U11719 ( .A(o[87]), .B(n9454), .Z(n9476) );
  XOR U11720 ( .A(n9477), .B(n9476), .Z(n9426) );
  NAND U11721 ( .A(y[7747]), .B(x[500]), .Z(n9330) );
  XNOR U11722 ( .A(n9331), .B(n9330), .Z(n9450) );
  AND U11723 ( .A(x[499]), .B(y[7748]), .Z(n9451) );
  XOR U11724 ( .A(n9450), .B(n9451), .Z(n9425) );
  XOR U11725 ( .A(n9426), .B(n9425), .Z(n9428) );
  XNOR U11726 ( .A(n9427), .B(n9428), .Z(n9434) );
  XOR U11727 ( .A(n9491), .B(n9490), .Z(n9493) );
  AND U11728 ( .A(x[500]), .B(y[7753]), .Z(n10368) );
  AND U11729 ( .A(x[493]), .B(y[7746]), .Z(n9332) );
  NAND U11730 ( .A(n10368), .B(n9332), .Z(n9336) );
  NAND U11731 ( .A(n9334), .B(n9333), .Z(n9335) );
  NAND U11732 ( .A(n9336), .B(n9335), .Z(n9485) );
  NAND U11733 ( .A(n9338), .B(n9337), .Z(n9342) );
  NAND U11734 ( .A(n9340), .B(n9339), .Z(n9341) );
  NAND U11735 ( .A(n9342), .B(n9341), .Z(n9439) );
  AND U11736 ( .A(x[493]), .B(y[7754]), .Z(n9413) );
  AND U11737 ( .A(x[482]), .B(y[7765]), .Z(n9414) );
  XOR U11738 ( .A(n9413), .B(n9414), .Z(n9415) );
  AND U11739 ( .A(x[501]), .B(y[7746]), .Z(n9416) );
  XOR U11740 ( .A(n9415), .B(n9416), .Z(n9438) );
  AND U11741 ( .A(x[492]), .B(y[7755]), .Z(n9468) );
  AND U11742 ( .A(x[481]), .B(y[7766]), .Z(n9469) );
  XOR U11743 ( .A(n9468), .B(n9469), .Z(n9471) );
  AND U11744 ( .A(o[86]), .B(n9343), .Z(n9470) );
  XOR U11745 ( .A(n9471), .B(n9470), .Z(n9437) );
  XOR U11746 ( .A(n9438), .B(n9437), .Z(n9440) );
  XOR U11747 ( .A(n9439), .B(n9440), .Z(n9484) );
  XOR U11748 ( .A(n9485), .B(n9484), .Z(n9487) );
  AND U11749 ( .A(x[495]), .B(y[7760]), .Z(n10585) );
  NAND U11750 ( .A(n10585), .B(n9344), .Z(n9348) );
  NANDN U11751 ( .A(n9346), .B(n9345), .Z(n9347) );
  NAND U11752 ( .A(n9348), .B(n9347), .Z(n9421) );
  AND U11753 ( .A(x[494]), .B(y[7753]), .Z(n9407) );
  AND U11754 ( .A(x[483]), .B(y[7764]), .Z(n9408) );
  XOR U11755 ( .A(n9407), .B(n9408), .Z(n9409) );
  AND U11756 ( .A(x[484]), .B(y[7763]), .Z(n9410) );
  XOR U11757 ( .A(n9409), .B(n9410), .Z(n9420) );
  AND U11758 ( .A(x[485]), .B(y[7762]), .Z(n9401) );
  AND U11759 ( .A(x[498]), .B(y[7749]), .Z(n9402) );
  XOR U11760 ( .A(n9401), .B(n9402), .Z(n9404) );
  AND U11761 ( .A(x[497]), .B(y[7750]), .Z(n9403) );
  XOR U11762 ( .A(n9404), .B(n9403), .Z(n9419) );
  XOR U11763 ( .A(n9420), .B(n9419), .Z(n9422) );
  XOR U11764 ( .A(n9421), .B(n9422), .Z(n9486) );
  XOR U11765 ( .A(n9487), .B(n9486), .Z(n9492) );
  XOR U11766 ( .A(n9493), .B(n9492), .Z(n9496) );
  XOR U11767 ( .A(n9497), .B(n9496), .Z(n9498) );
  XOR U11768 ( .A(n9499), .B(n9498), .Z(n9386) );
  NAND U11769 ( .A(n9350), .B(n9349), .Z(n9354) );
  NAND U11770 ( .A(n9352), .B(n9351), .Z(n9353) );
  NAND U11771 ( .A(n9354), .B(n9353), .Z(n9505) );
  NAND U11772 ( .A(n9356), .B(n9355), .Z(n9360) );
  NAND U11773 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U11774 ( .A(n9360), .B(n9359), .Z(n9503) );
  NAND U11775 ( .A(n9362), .B(n9361), .Z(n9366) );
  NAND U11776 ( .A(n9364), .B(n9363), .Z(n9365) );
  AND U11777 ( .A(n9366), .B(n9365), .Z(n9502) );
  XOR U11778 ( .A(n9503), .B(n9502), .Z(n9504) );
  XOR U11779 ( .A(n9505), .B(n9504), .Z(n9384) );
  NAND U11780 ( .A(n9368), .B(n9367), .Z(n9372) );
  NANDN U11781 ( .A(n9370), .B(n9369), .Z(n9371) );
  AND U11782 ( .A(n9372), .B(n9371), .Z(n9383) );
  XNOR U11783 ( .A(n9517), .B(n9516), .Z(n9522) );
  NANDN U11784 ( .A(n9377), .B(n9376), .Z(n9381) );
  NANDN U11785 ( .A(n9379), .B(n9378), .Z(n9380) );
  AND U11786 ( .A(n9381), .B(n9380), .Z(n9520) );
  XOR U11787 ( .A(n9521), .B(n9520), .Z(n9382) );
  XNOR U11788 ( .A(n9522), .B(n9382), .Z(N184) );
  NANDN U11789 ( .A(n9384), .B(n9383), .Z(n9388) );
  NANDN U11790 ( .A(n9386), .B(n9385), .Z(n9387) );
  AND U11791 ( .A(n9388), .B(n9387), .Z(n9526) );
  NAND U11792 ( .A(n9390), .B(n9389), .Z(n9394) );
  NAND U11793 ( .A(n9392), .B(n9391), .Z(n9393) );
  NAND U11794 ( .A(n9394), .B(n9393), .Z(n9599) );
  NAND U11795 ( .A(n9396), .B(n9395), .Z(n9400) );
  NAND U11796 ( .A(n9398), .B(n9397), .Z(n9399) );
  NAND U11797 ( .A(n9400), .B(n9399), .Z(n9597) );
  NAND U11798 ( .A(n9402), .B(n9401), .Z(n9406) );
  NAND U11799 ( .A(n9404), .B(n9403), .Z(n9405) );
  NAND U11800 ( .A(n9406), .B(n9405), .Z(n9634) );
  AND U11801 ( .A(x[480]), .B(y[7768]), .Z(n9579) );
  AND U11802 ( .A(x[504]), .B(y[7744]), .Z(n9578) );
  XOR U11803 ( .A(n9579), .B(n9578), .Z(n9581) );
  AND U11804 ( .A(x[503]), .B(y[7745]), .Z(n9571) );
  XOR U11805 ( .A(n9571), .B(o[88]), .Z(n9580) );
  XOR U11806 ( .A(n9581), .B(n9580), .Z(n9632) );
  AND U11807 ( .A(x[487]), .B(y[7761]), .Z(n9566) );
  AND U11808 ( .A(x[498]), .B(y[7750]), .Z(n9565) );
  XOR U11809 ( .A(n9566), .B(n9565), .Z(n9568) );
  AND U11810 ( .A(x[497]), .B(y[7751]), .Z(n9567) );
  XOR U11811 ( .A(n9568), .B(n9567), .Z(n9631) );
  XOR U11812 ( .A(n9632), .B(n9631), .Z(n9633) );
  XOR U11813 ( .A(n9634), .B(n9633), .Z(n9611) );
  NAND U11814 ( .A(n9408), .B(n9407), .Z(n9412) );
  NAND U11815 ( .A(n9410), .B(n9409), .Z(n9411) );
  NAND U11816 ( .A(n9412), .B(n9411), .Z(n9609) );
  NAND U11817 ( .A(n9414), .B(n9413), .Z(n9418) );
  NAND U11818 ( .A(n9416), .B(n9415), .Z(n9417) );
  NAND U11819 ( .A(n9418), .B(n9417), .Z(n9608) );
  XOR U11820 ( .A(n9609), .B(n9608), .Z(n9610) );
  XOR U11821 ( .A(n9611), .B(n9610), .Z(n9596) );
  XOR U11822 ( .A(n9597), .B(n9596), .Z(n9598) );
  XNOR U11823 ( .A(n9599), .B(n9598), .Z(n9604) );
  NAND U11824 ( .A(n9420), .B(n9419), .Z(n9424) );
  NAND U11825 ( .A(n9422), .B(n9421), .Z(n9423) );
  AND U11826 ( .A(n9424), .B(n9423), .Z(n9650) );
  NAND U11827 ( .A(n9426), .B(n9425), .Z(n9430) );
  NAND U11828 ( .A(n9428), .B(n9427), .Z(n9429) );
  AND U11829 ( .A(n9430), .B(n9429), .Z(n9649) );
  XOR U11830 ( .A(n9650), .B(n9649), .Z(n9652) );
  NAND U11831 ( .A(n9432), .B(n9431), .Z(n9436) );
  NANDN U11832 ( .A(n9434), .B(n9433), .Z(n9435) );
  AND U11833 ( .A(n9436), .B(n9435), .Z(n9651) );
  XOR U11834 ( .A(n9652), .B(n9651), .Z(n9602) );
  NAND U11835 ( .A(n9438), .B(n9437), .Z(n9442) );
  NAND U11836 ( .A(n9440), .B(n9439), .Z(n9441) );
  AND U11837 ( .A(n9442), .B(n9441), .Z(n9603) );
  XOR U11838 ( .A(n9602), .B(n9603), .Z(n9605) );
  XOR U11839 ( .A(n9604), .B(n9605), .Z(n9655) );
  NAND U11840 ( .A(n9444), .B(n9443), .Z(n9448) );
  NAND U11841 ( .A(n9446), .B(n9445), .Z(n9447) );
  AND U11842 ( .A(n9448), .B(n9447), .Z(n9656) );
  XOR U11843 ( .A(n9655), .B(n9656), .Z(n9658) );
  AND U11844 ( .A(x[500]), .B(y[7751]), .Z(n9449) );
  NAND U11845 ( .A(n9449), .B(n9620), .Z(n9453) );
  NAND U11846 ( .A(n9451), .B(n9450), .Z(n9452) );
  NAND U11847 ( .A(n9453), .B(n9452), .Z(n9646) );
  AND U11848 ( .A(x[502]), .B(y[7746]), .Z(n9555) );
  XOR U11849 ( .A(n9556), .B(n9555), .Z(n9554) );
  AND U11850 ( .A(x[482]), .B(y[7766]), .Z(n9553) );
  XOR U11851 ( .A(n9554), .B(n9553), .Z(n9644) );
  AND U11852 ( .A(x[481]), .B(y[7767]), .Z(n9561) );
  XOR U11853 ( .A(n9562), .B(n9561), .Z(n9560) );
  AND U11854 ( .A(o[87]), .B(n9454), .Z(n9559) );
  XOR U11855 ( .A(n9560), .B(n9559), .Z(n9643) );
  XOR U11856 ( .A(n9644), .B(n9643), .Z(n9645) );
  XOR U11857 ( .A(n9646), .B(n9645), .Z(n9591) );
  NAND U11858 ( .A(n9456), .B(n9455), .Z(n9460) );
  NAND U11859 ( .A(n9458), .B(n9457), .Z(n9459) );
  NAND U11860 ( .A(n9460), .B(n9459), .Z(n9640) );
  AND U11861 ( .A(y[7752]), .B(x[496]), .Z(n9462) );
  NAND U11862 ( .A(y[7747]), .B(x[501]), .Z(n9461) );
  XNOR U11863 ( .A(n9462), .B(n9461), .Z(n9622) );
  AND U11864 ( .A(x[485]), .B(y[7763]), .Z(n9621) );
  XOR U11865 ( .A(n9622), .B(n9621), .Z(n9638) );
  AND U11866 ( .A(x[486]), .B(y[7762]), .Z(n9956) );
  AND U11867 ( .A(x[500]), .B(y[7748]), .Z(n9761) );
  XOR U11868 ( .A(n9956), .B(n9761), .Z(n9628) );
  AND U11869 ( .A(x[499]), .B(y[7749]), .Z(n9627) );
  XOR U11870 ( .A(n9628), .B(n9627), .Z(n9637) );
  XOR U11871 ( .A(n9638), .B(n9637), .Z(n9639) );
  XOR U11872 ( .A(n9640), .B(n9639), .Z(n9617) );
  NANDN U11873 ( .A(n9686), .B(n9463), .Z(n9467) );
  NANDN U11874 ( .A(n9465), .B(n9464), .Z(n9466) );
  NAND U11875 ( .A(n9467), .B(n9466), .Z(n9615) );
  NAND U11876 ( .A(n9469), .B(n9468), .Z(n9473) );
  NAND U11877 ( .A(n9471), .B(n9470), .Z(n9472) );
  NAND U11878 ( .A(n9473), .B(n9472), .Z(n9614) );
  XOR U11879 ( .A(n9615), .B(n9614), .Z(n9616) );
  XOR U11880 ( .A(n9617), .B(n9616), .Z(n9590) );
  XOR U11881 ( .A(n9591), .B(n9590), .Z(n9593) );
  NAND U11882 ( .A(n9475), .B(n9474), .Z(n9479) );
  NAND U11883 ( .A(n9477), .B(n9476), .Z(n9478) );
  NAND U11884 ( .A(n9479), .B(n9478), .Z(n9585) );
  AND U11885 ( .A(x[483]), .B(y[7765]), .Z(n9574) );
  XOR U11886 ( .A(n9575), .B(n9574), .Z(n9573) );
  AND U11887 ( .A(x[484]), .B(y[7764]), .Z(n9572) );
  XOR U11888 ( .A(n9573), .B(n9572), .Z(n9584) );
  XOR U11889 ( .A(n9585), .B(n9584), .Z(n9587) );
  AND U11890 ( .A(y[7759]), .B(x[489]), .Z(n9481) );
  NAND U11891 ( .A(y[7758]), .B(x[490]), .Z(n9480) );
  XNOR U11892 ( .A(n9481), .B(n9480), .Z(n9547) );
  AND U11893 ( .A(y[7754]), .B(x[494]), .Z(n9483) );
  NAND U11894 ( .A(y[7760]), .B(x[488]), .Z(n9482) );
  XNOR U11895 ( .A(n9483), .B(n9482), .Z(n9549) );
  NAND U11896 ( .A(x[491]), .B(y[7757]), .Z(n9550) );
  XOR U11897 ( .A(n9547), .B(n9546), .Z(n9586) );
  XOR U11898 ( .A(n9587), .B(n9586), .Z(n9592) );
  XNOR U11899 ( .A(n9593), .B(n9592), .Z(n9540) );
  NAND U11900 ( .A(n9485), .B(n9484), .Z(n9489) );
  NAND U11901 ( .A(n9487), .B(n9486), .Z(n9488) );
  AND U11902 ( .A(n9489), .B(n9488), .Z(n9539) );
  XOR U11903 ( .A(n9540), .B(n9539), .Z(n9541) );
  NAND U11904 ( .A(n9491), .B(n9490), .Z(n9495) );
  NAND U11905 ( .A(n9493), .B(n9492), .Z(n9494) );
  AND U11906 ( .A(n9495), .B(n9494), .Z(n9542) );
  XOR U11907 ( .A(n9541), .B(n9542), .Z(n9657) );
  XNOR U11908 ( .A(n9658), .B(n9657), .Z(n9524) );
  NAND U11909 ( .A(n9497), .B(n9496), .Z(n9501) );
  NAND U11910 ( .A(n9499), .B(n9498), .Z(n9500) );
  NAND U11911 ( .A(n9501), .B(n9500), .Z(n9536) );
  NAND U11912 ( .A(n9503), .B(n9502), .Z(n9507) );
  NAND U11913 ( .A(n9505), .B(n9504), .Z(n9506) );
  NAND U11914 ( .A(n9507), .B(n9506), .Z(n9534) );
  NAND U11915 ( .A(n9509), .B(n9508), .Z(n9513) );
  NAND U11916 ( .A(n9511), .B(n9510), .Z(n9512) );
  NAND U11917 ( .A(n9513), .B(n9512), .Z(n9533) );
  XOR U11918 ( .A(n9534), .B(n9533), .Z(n9535) );
  XNOR U11919 ( .A(n9536), .B(n9535), .Z(n9525) );
  XOR U11920 ( .A(n9524), .B(n9525), .Z(n9527) );
  XNOR U11921 ( .A(n9526), .B(n9527), .Z(n9532) );
  NANDN U11922 ( .A(n9515), .B(n9514), .Z(n9519) );
  NAND U11923 ( .A(n9517), .B(n9516), .Z(n9518) );
  NAND U11924 ( .A(n9519), .B(n9518), .Z(n9530) );
  XOR U11925 ( .A(n9530), .B(n9531), .Z(n9523) );
  XNOR U11926 ( .A(n9532), .B(n9523), .Z(N185) );
  NANDN U11927 ( .A(n9525), .B(n9524), .Z(n9529) );
  NANDN U11928 ( .A(n9527), .B(n9526), .Z(n9528) );
  AND U11929 ( .A(n9529), .B(n9528), .Z(n9808) );
  NAND U11930 ( .A(n9534), .B(n9533), .Z(n9538) );
  NAND U11931 ( .A(n9536), .B(n9535), .Z(n9537) );
  NAND U11932 ( .A(n9538), .B(n9537), .Z(n9805) );
  NAND U11933 ( .A(n9540), .B(n9539), .Z(n9544) );
  NAND U11934 ( .A(n9542), .B(n9541), .Z(n9543) );
  AND U11935 ( .A(n9544), .B(n9543), .Z(n9663) );
  AND U11936 ( .A(x[494]), .B(y[7760]), .Z(n10637) );
  NAND U11937 ( .A(n10637), .B(n9548), .Z(n9552) );
  NANDN U11938 ( .A(n9550), .B(n9549), .Z(n9551) );
  AND U11939 ( .A(n9552), .B(n9551), .Z(n9739) );
  NAND U11940 ( .A(x[491]), .B(y[7758]), .Z(n9757) );
  NAND U11941 ( .A(x[492]), .B(y[7757]), .Z(n9756) );
  NAND U11942 ( .A(x[487]), .B(y[7762]), .Z(n9755) );
  XNOR U11943 ( .A(n9756), .B(n9755), .Z(n9758) );
  NAND U11944 ( .A(x[504]), .B(y[7745]), .Z(n9754) );
  XNOR U11945 ( .A(o[89]), .B(n9754), .Z(n9724) );
  NAND U11946 ( .A(x[481]), .B(y[7768]), .Z(n9725) );
  NAND U11947 ( .A(x[493]), .B(y[7756]), .Z(n9727) );
  XOR U11948 ( .A(n9736), .B(n9737), .Z(n9738) );
  XOR U11949 ( .A(n9711), .B(n9710), .Z(n9713) );
  AND U11950 ( .A(n9554), .B(n9553), .Z(n9558) );
  NAND U11951 ( .A(n9556), .B(n9555), .Z(n9557) );
  NANDN U11952 ( .A(n9558), .B(n9557), .Z(n9699) );
  AND U11953 ( .A(n9560), .B(n9559), .Z(n9564) );
  NAND U11954 ( .A(n9562), .B(n9561), .Z(n9563) );
  NANDN U11955 ( .A(n9564), .B(n9563), .Z(n9698) );
  XOR U11956 ( .A(n9699), .B(n9698), .Z(n9701) );
  NAND U11957 ( .A(n9566), .B(n9565), .Z(n9570) );
  NAND U11958 ( .A(n9568), .B(n9567), .Z(n9569) );
  NAND U11959 ( .A(n9570), .B(n9569), .Z(n9695) );
  NAND U11960 ( .A(x[488]), .B(y[7761]), .Z(n9689) );
  XNOR U11961 ( .A(n9686), .B(n9687), .Z(n9688) );
  XNOR U11962 ( .A(n9689), .B(n9688), .Z(n9693) );
  AND U11963 ( .A(n9571), .B(o[88]), .Z(n9683) );
  NAND U11964 ( .A(x[505]), .B(y[7744]), .Z(n9681) );
  NAND U11965 ( .A(x[480]), .B(y[7769]), .Z(n9680) );
  XOR U11966 ( .A(n9681), .B(n9680), .Z(n9682) );
  XOR U11967 ( .A(n9683), .B(n9682), .Z(n9692) );
  XOR U11968 ( .A(n9693), .B(n9692), .Z(n9694) );
  XOR U11969 ( .A(n9695), .B(n9694), .Z(n9700) );
  XOR U11970 ( .A(n9701), .B(n9700), .Z(n9712) );
  XNOR U11971 ( .A(n9713), .B(n9712), .Z(n9799) );
  AND U11972 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U11973 ( .A(n9575), .B(n9574), .Z(n9576) );
  NANDN U11974 ( .A(n9577), .B(n9576), .Z(n9775) );
  NAND U11975 ( .A(n9579), .B(n9578), .Z(n9583) );
  NAND U11976 ( .A(n9581), .B(n9580), .Z(n9582) );
  NAND U11977 ( .A(n9583), .B(n9582), .Z(n9773) );
  AND U11978 ( .A(x[494]), .B(y[7755]), .Z(n9730) );
  AND U11979 ( .A(x[482]), .B(y[7767]), .Z(n9731) );
  XOR U11980 ( .A(n9730), .B(n9731), .Z(n9732) );
  AND U11981 ( .A(x[483]), .B(y[7766]), .Z(n9733) );
  XOR U11982 ( .A(n9732), .B(n9733), .Z(n9772) );
  XOR U11983 ( .A(n9773), .B(n9772), .Z(n9774) );
  XNOR U11984 ( .A(n9775), .B(n9774), .Z(n9797) );
  NAND U11985 ( .A(n9585), .B(n9584), .Z(n9589) );
  NAND U11986 ( .A(n9587), .B(n9586), .Z(n9588) );
  AND U11987 ( .A(n9589), .B(n9588), .Z(n9796) );
  XOR U11988 ( .A(n9797), .B(n9796), .Z(n9798) );
  XOR U11989 ( .A(n9799), .B(n9798), .Z(n9790) );
  NAND U11990 ( .A(n9591), .B(n9590), .Z(n9595) );
  NAND U11991 ( .A(n9593), .B(n9592), .Z(n9594) );
  AND U11992 ( .A(n9595), .B(n9594), .Z(n9791) );
  XOR U11993 ( .A(n9790), .B(n9791), .Z(n9792) );
  NAND U11994 ( .A(n9597), .B(n9596), .Z(n9601) );
  NAND U11995 ( .A(n9599), .B(n9598), .Z(n9600) );
  AND U11996 ( .A(n9601), .B(n9600), .Z(n9793) );
  XOR U11997 ( .A(n9792), .B(n9793), .Z(n9662) );
  NAND U11998 ( .A(n9603), .B(n9602), .Z(n9607) );
  NAND U11999 ( .A(n9605), .B(n9604), .Z(n9606) );
  NAND U12000 ( .A(n9607), .B(n9606), .Z(n9670) );
  NAND U12001 ( .A(n9609), .B(n9608), .Z(n9613) );
  NAND U12002 ( .A(n9611), .B(n9610), .Z(n9612) );
  NAND U12003 ( .A(n9613), .B(n9612), .Z(n9675) );
  NAND U12004 ( .A(n9615), .B(n9614), .Z(n9619) );
  NAND U12005 ( .A(n9617), .B(n9616), .Z(n9618) );
  NAND U12006 ( .A(n9619), .B(n9618), .Z(n9674) );
  XOR U12007 ( .A(n9675), .B(n9674), .Z(n9677) );
  AND U12008 ( .A(x[501]), .B(y[7752]), .Z(n10651) );
  NAND U12009 ( .A(n10651), .B(n9620), .Z(n9624) );
  NAND U12010 ( .A(n9622), .B(n9621), .Z(n9623) );
  NAND U12011 ( .A(n9624), .B(n9623), .Z(n9780) );
  NAND U12012 ( .A(x[502]), .B(y[7747]), .Z(n9750) );
  NAND U12013 ( .A(x[485]), .B(y[7764]), .Z(n9749) );
  NAND U12014 ( .A(x[497]), .B(y[7752]), .Z(n9748) );
  XOR U12015 ( .A(n9749), .B(n9748), .Z(n9751) );
  XOR U12016 ( .A(n9750), .B(n9751), .Z(n9779) );
  AND U12017 ( .A(y[7749]), .B(x[500]), .Z(n9626) );
  NAND U12018 ( .A(y[7748]), .B(x[501]), .Z(n9625) );
  XNOR U12019 ( .A(n9626), .B(n9625), .Z(n9763) );
  AND U12020 ( .A(x[499]), .B(y[7750]), .Z(n9762) );
  XOR U12021 ( .A(n9763), .B(n9762), .Z(n9778) );
  XNOR U12022 ( .A(n9780), .B(n9781), .Z(n9705) );
  NAND U12023 ( .A(n9956), .B(n9761), .Z(n9630) );
  NAND U12024 ( .A(n9628), .B(n9627), .Z(n9629) );
  NAND U12025 ( .A(n9630), .B(n9629), .Z(n9786) );
  NAND U12026 ( .A(x[495]), .B(y[7754]), .Z(n9768) );
  NAND U12027 ( .A(x[498]), .B(y[7751]), .Z(n9767) );
  NAND U12028 ( .A(x[486]), .B(y[7763]), .Z(n9766) );
  XOR U12029 ( .A(n9767), .B(n9766), .Z(n9769) );
  XOR U12030 ( .A(n9768), .B(n9769), .Z(n9785) );
  NAND U12031 ( .A(x[503]), .B(y[7746]), .Z(n9744) );
  NAND U12032 ( .A(x[484]), .B(y[7765]), .Z(n9743) );
  NAND U12033 ( .A(x[496]), .B(y[7753]), .Z(n9742) );
  XOR U12034 ( .A(n9743), .B(n9742), .Z(n9745) );
  XNOR U12035 ( .A(n9744), .B(n9745), .Z(n9784) );
  XOR U12036 ( .A(n9786), .B(n9787), .Z(n9704) );
  XOR U12037 ( .A(n9705), .B(n9704), .Z(n9707) );
  NAND U12038 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U12039 ( .A(n9634), .B(n9633), .Z(n9635) );
  AND U12040 ( .A(n9636), .B(n9635), .Z(n9706) );
  XNOR U12041 ( .A(n9707), .B(n9706), .Z(n9719) );
  NAND U12042 ( .A(n9638), .B(n9637), .Z(n9642) );
  NAND U12043 ( .A(n9640), .B(n9639), .Z(n9641) );
  NAND U12044 ( .A(n9642), .B(n9641), .Z(n9717) );
  NAND U12045 ( .A(n9644), .B(n9643), .Z(n9648) );
  NAND U12046 ( .A(n9646), .B(n9645), .Z(n9647) );
  NAND U12047 ( .A(n9648), .B(n9647), .Z(n9716) );
  XOR U12048 ( .A(n9717), .B(n9716), .Z(n9718) );
  XOR U12049 ( .A(n9719), .B(n9718), .Z(n9676) );
  XOR U12050 ( .A(n9677), .B(n9676), .Z(n9669) );
  NAND U12051 ( .A(n9650), .B(n9649), .Z(n9654) );
  NAND U12052 ( .A(n9652), .B(n9651), .Z(n9653) );
  NAND U12053 ( .A(n9654), .B(n9653), .Z(n9668) );
  XOR U12054 ( .A(n9670), .B(n9671), .Z(n9664) );
  XNOR U12055 ( .A(n9665), .B(n9664), .Z(n9803) );
  NAND U12056 ( .A(n9656), .B(n9655), .Z(n9660) );
  NAND U12057 ( .A(n9658), .B(n9657), .Z(n9659) );
  AND U12058 ( .A(n9660), .B(n9659), .Z(n9802) );
  XOR U12059 ( .A(n9803), .B(n9802), .Z(n9804) );
  XOR U12060 ( .A(n9805), .B(n9804), .Z(n9810) );
  XNOR U12061 ( .A(n9809), .B(n9810), .Z(n9661) );
  XOR U12062 ( .A(n9808), .B(n9661), .Z(N186) );
  NANDN U12063 ( .A(n9663), .B(n9662), .Z(n9667) );
  NAND U12064 ( .A(n9665), .B(n9664), .Z(n9666) );
  AND U12065 ( .A(n9667), .B(n9666), .Z(n9812) );
  NANDN U12066 ( .A(n9669), .B(n9668), .Z(n9673) );
  NAND U12067 ( .A(n9671), .B(n9670), .Z(n9672) );
  NAND U12068 ( .A(n9673), .B(n9672), .Z(n9813) );
  NAND U12069 ( .A(n9675), .B(n9674), .Z(n9679) );
  NAND U12070 ( .A(n9677), .B(n9676), .Z(n9678) );
  NAND U12071 ( .A(n9679), .B(n9678), .Z(n9830) );
  AND U12072 ( .A(x[482]), .B(y[7768]), .Z(n9851) );
  XOR U12073 ( .A(n9852), .B(n9851), .Z(n9854) );
  NAND U12074 ( .A(x[504]), .B(y[7746]), .Z(n9853) );
  XNOR U12075 ( .A(n9854), .B(n9853), .Z(n9888) );
  NAND U12076 ( .A(n9681), .B(n9680), .Z(n9685) );
  NANDN U12077 ( .A(n9683), .B(n9682), .Z(n9684) );
  AND U12078 ( .A(n9685), .B(n9684), .Z(n9887) );
  XOR U12079 ( .A(n9888), .B(n9887), .Z(n9890) );
  NANDN U12080 ( .A(n9687), .B(n9686), .Z(n9691) );
  NAND U12081 ( .A(n9689), .B(n9688), .Z(n9690) );
  AND U12082 ( .A(n9691), .B(n9690), .Z(n9889) );
  XOR U12083 ( .A(n9890), .B(n9889), .Z(n9925) );
  NAND U12084 ( .A(n9693), .B(n9692), .Z(n9697) );
  NAND U12085 ( .A(n9695), .B(n9694), .Z(n9696) );
  AND U12086 ( .A(n9697), .B(n9696), .Z(n9924) );
  NAND U12087 ( .A(n9699), .B(n9698), .Z(n9703) );
  NAND U12088 ( .A(n9701), .B(n9700), .Z(n9702) );
  AND U12089 ( .A(n9703), .B(n9702), .Z(n9926) );
  XOR U12090 ( .A(n9927), .B(n9926), .Z(n9921) );
  NAND U12091 ( .A(n9705), .B(n9704), .Z(n9709) );
  NAND U12092 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U12093 ( .A(n9709), .B(n9708), .Z(n9918) );
  NAND U12094 ( .A(n9711), .B(n9710), .Z(n9715) );
  NAND U12095 ( .A(n9713), .B(n9712), .Z(n9714) );
  AND U12096 ( .A(n9715), .B(n9714), .Z(n9919) );
  XOR U12097 ( .A(n9918), .B(n9919), .Z(n9920) );
  XNOR U12098 ( .A(n9921), .B(n9920), .Z(n9828) );
  NAND U12099 ( .A(n9717), .B(n9716), .Z(n9721) );
  NAND U12100 ( .A(n9719), .B(n9718), .Z(n9720) );
  NAND U12101 ( .A(n9721), .B(n9720), .Z(n9835) );
  AND U12102 ( .A(x[492]), .B(y[7758]), .Z(n10034) );
  AND U12103 ( .A(x[485]), .B(y[7765]), .Z(n9901) );
  XOR U12104 ( .A(n10034), .B(n9901), .Z(n9903) );
  NAND U12105 ( .A(x[490]), .B(y[7760]), .Z(n9902) );
  XNOR U12106 ( .A(n9903), .B(n9902), .Z(n9933) );
  AND U12107 ( .A(x[487]), .B(y[7763]), .Z(n9931) );
  AND U12108 ( .A(y[7764]), .B(x[486]), .Z(n9723) );
  NAND U12109 ( .A(y[7762]), .B(x[488]), .Z(n9722) );
  XNOR U12110 ( .A(n9723), .B(n9722), .Z(n9957) );
  NAND U12111 ( .A(x[489]), .B(y[7761]), .Z(n9958) );
  XNOR U12112 ( .A(n9957), .B(n9958), .Z(n9930) );
  XOR U12113 ( .A(n9931), .B(n9930), .Z(n9932) );
  XOR U12114 ( .A(n9933), .B(n9932), .Z(n9877) );
  NANDN U12115 ( .A(n9725), .B(n9724), .Z(n9729) );
  NANDN U12116 ( .A(n9727), .B(n9726), .Z(n9728) );
  NAND U12117 ( .A(n9729), .B(n9728), .Z(n9876) );
  NAND U12118 ( .A(n9731), .B(n9730), .Z(n9735) );
  NAND U12119 ( .A(n9733), .B(n9732), .Z(n9734) );
  NAND U12120 ( .A(n9735), .B(n9734), .Z(n9875) );
  XNOR U12121 ( .A(n9876), .B(n9875), .Z(n9878) );
  NAND U12122 ( .A(n9737), .B(n9736), .Z(n9741) );
  NANDN U12123 ( .A(n9739), .B(n9738), .Z(n9740) );
  AND U12124 ( .A(n9741), .B(n9740), .Z(n9912) );
  NAND U12125 ( .A(n9743), .B(n9742), .Z(n9747) );
  NAND U12126 ( .A(n9745), .B(n9744), .Z(n9746) );
  AND U12127 ( .A(n9747), .B(n9746), .Z(n9840) );
  NAND U12128 ( .A(n9749), .B(n9748), .Z(n9753) );
  NAND U12129 ( .A(n9751), .B(n9750), .Z(n9752) );
  AND U12130 ( .A(n9753), .B(n9752), .Z(n9839) );
  XOR U12131 ( .A(n9840), .B(n9839), .Z(n9842) );
  ANDN U12132 ( .B(o[89]), .A(n9754), .Z(n9950) );
  NAND U12133 ( .A(x[494]), .B(y[7756]), .Z(n9951) );
  XNOR U12134 ( .A(n9950), .B(n9951), .Z(n9952) );
  NAND U12135 ( .A(x[481]), .B(y[7769]), .Z(n9953) );
  XNOR U12136 ( .A(n9952), .B(n9953), .Z(n9894) );
  NAND U12137 ( .A(x[505]), .B(y[7745]), .Z(n9961) );
  XNOR U12138 ( .A(o[90]), .B(n9961), .Z(n9906) );
  NAND U12139 ( .A(x[506]), .B(y[7744]), .Z(n9907) );
  XNOR U12140 ( .A(n9906), .B(n9907), .Z(n9909) );
  AND U12141 ( .A(x[480]), .B(y[7770]), .Z(n9908) );
  XOR U12142 ( .A(n9909), .B(n9908), .Z(n9893) );
  XOR U12143 ( .A(n9894), .B(n9893), .Z(n9896) );
  NAND U12144 ( .A(n9756), .B(n9755), .Z(n9760) );
  NANDN U12145 ( .A(n9758), .B(n9757), .Z(n9759) );
  AND U12146 ( .A(n9760), .B(n9759), .Z(n9895) );
  XOR U12147 ( .A(n9896), .B(n9895), .Z(n9841) );
  XNOR U12148 ( .A(n9842), .B(n9841), .Z(n9883) );
  AND U12149 ( .A(x[501]), .B(y[7749]), .Z(n9944) );
  NAND U12150 ( .A(n9944), .B(n9761), .Z(n9765) );
  NAND U12151 ( .A(n9763), .B(n9762), .Z(n9764) );
  NAND U12152 ( .A(n9765), .B(n9764), .Z(n9871) );
  XOR U12153 ( .A(n9945), .B(n9944), .Z(n9947) );
  NAND U12154 ( .A(x[500]), .B(y[7750]), .Z(n9946) );
  XNOR U12155 ( .A(n9947), .B(n9946), .Z(n9870) );
  NAND U12156 ( .A(x[503]), .B(y[7747]), .Z(n9858) );
  XNOR U12157 ( .A(n9857), .B(n9858), .Z(n9860) );
  AND U12158 ( .A(x[502]), .B(y[7748]), .Z(n9859) );
  XOR U12159 ( .A(n9860), .B(n9859), .Z(n9869) );
  XOR U12160 ( .A(n9870), .B(n9869), .Z(n9872) );
  XOR U12161 ( .A(n9871), .B(n9872), .Z(n9882) );
  AND U12162 ( .A(x[483]), .B(y[7767]), .Z(n9936) );
  NAND U12163 ( .A(x[499]), .B(y[7751]), .Z(n9937) );
  XNOR U12164 ( .A(n9936), .B(n9937), .Z(n9938) );
  NAND U12165 ( .A(x[491]), .B(y[7759]), .Z(n9939) );
  XNOR U12166 ( .A(n9938), .B(n9939), .Z(n9846) );
  AND U12167 ( .A(x[484]), .B(y[7766]), .Z(n9863) );
  XOR U12168 ( .A(n9864), .B(n9863), .Z(n9866) );
  XOR U12169 ( .A(n9866), .B(n9865), .Z(n9845) );
  XOR U12170 ( .A(n9846), .B(n9845), .Z(n9848) );
  NAND U12171 ( .A(n9767), .B(n9766), .Z(n9771) );
  NAND U12172 ( .A(n9769), .B(n9768), .Z(n9770) );
  AND U12173 ( .A(n9771), .B(n9770), .Z(n9847) );
  XNOR U12174 ( .A(n9848), .B(n9847), .Z(n9881) );
  XOR U12175 ( .A(n9883), .B(n9884), .Z(n9915) );
  XNOR U12176 ( .A(n9914), .B(n9915), .Z(n9834) );
  NAND U12177 ( .A(n9773), .B(n9772), .Z(n9777) );
  NAND U12178 ( .A(n9775), .B(n9774), .Z(n9776) );
  NAND U12179 ( .A(n9777), .B(n9776), .Z(n9964) );
  NANDN U12180 ( .A(n9779), .B(n9778), .Z(n9783) );
  NAND U12181 ( .A(n9781), .B(n9780), .Z(n9782) );
  NAND U12182 ( .A(n9783), .B(n9782), .Z(n9963) );
  NANDN U12183 ( .A(n9785), .B(n9784), .Z(n9789) );
  NANDN U12184 ( .A(n9787), .B(n9786), .Z(n9788) );
  NAND U12185 ( .A(n9789), .B(n9788), .Z(n9962) );
  XOR U12186 ( .A(n9963), .B(n9962), .Z(n9965) );
  XOR U12187 ( .A(n9964), .B(n9965), .Z(n9833) );
  XOR U12188 ( .A(n9835), .B(n9836), .Z(n9827) );
  XOR U12189 ( .A(n9828), .B(n9827), .Z(n9829) );
  XOR U12190 ( .A(n9830), .B(n9829), .Z(n9824) );
  NAND U12191 ( .A(n9791), .B(n9790), .Z(n9795) );
  NAND U12192 ( .A(n9793), .B(n9792), .Z(n9794) );
  AND U12193 ( .A(n9795), .B(n9794), .Z(n9821) );
  NAND U12194 ( .A(n9797), .B(n9796), .Z(n9801) );
  NAND U12195 ( .A(n9799), .B(n9798), .Z(n9800) );
  AND U12196 ( .A(n9801), .B(n9800), .Z(n9822) );
  XOR U12197 ( .A(n9821), .B(n9822), .Z(n9823) );
  XOR U12198 ( .A(n9824), .B(n9823), .Z(n9814) );
  XNOR U12199 ( .A(n9815), .B(n9814), .Z(n9820) );
  NAND U12200 ( .A(n9803), .B(n9802), .Z(n9807) );
  NAND U12201 ( .A(n9805), .B(n9804), .Z(n9806) );
  NAND U12202 ( .A(n9807), .B(n9806), .Z(n9819) );
  XOR U12203 ( .A(n9819), .B(n9818), .Z(n9811) );
  XNOR U12204 ( .A(n9820), .B(n9811), .Z(N187) );
  NANDN U12205 ( .A(n9813), .B(n9812), .Z(n9817) );
  NAND U12206 ( .A(n9815), .B(n9814), .Z(n9816) );
  NAND U12207 ( .A(n9817), .B(n9816), .Z(n9976) );
  IV U12208 ( .A(n9976), .Z(n9975) );
  NAND U12209 ( .A(n9822), .B(n9821), .Z(n9826) );
  NAND U12210 ( .A(n9824), .B(n9823), .Z(n9825) );
  AND U12211 ( .A(n9826), .B(n9825), .Z(n9972) );
  NAND U12212 ( .A(n9828), .B(n9827), .Z(n9832) );
  NAND U12213 ( .A(n9830), .B(n9829), .Z(n9831) );
  AND U12214 ( .A(n9832), .B(n9831), .Z(n9970) );
  NANDN U12215 ( .A(n9834), .B(n9833), .Z(n9838) );
  NAND U12216 ( .A(n9836), .B(n9835), .Z(n9837) );
  NAND U12217 ( .A(n9838), .B(n9837), .Z(n9984) );
  NAND U12218 ( .A(n9840), .B(n9839), .Z(n9844) );
  NAND U12219 ( .A(n9842), .B(n9841), .Z(n9843) );
  NAND U12220 ( .A(n9844), .B(n9843), .Z(n10101) );
  NAND U12221 ( .A(n9846), .B(n9845), .Z(n9850) );
  NAND U12222 ( .A(n9848), .B(n9847), .Z(n9849) );
  NAND U12223 ( .A(n9850), .B(n9849), .Z(n10099) );
  NAND U12224 ( .A(n9852), .B(n9851), .Z(n9856) );
  ANDN U12225 ( .B(n9854), .A(n9853), .Z(n9855) );
  ANDN U12226 ( .B(n9856), .A(n9855), .Z(n10007) );
  NANDN U12227 ( .A(n9858), .B(n9857), .Z(n9862) );
  NAND U12228 ( .A(n9860), .B(n9859), .Z(n9861) );
  NAND U12229 ( .A(n9862), .B(n9861), .Z(n10006) );
  XNOR U12230 ( .A(n10007), .B(n10006), .Z(n10008) );
  NAND U12231 ( .A(n9864), .B(n9863), .Z(n9868) );
  AND U12232 ( .A(n9866), .B(n9865), .Z(n9867) );
  ANDN U12233 ( .B(n9868), .A(n9867), .Z(n10021) );
  AND U12234 ( .A(x[480]), .B(y[7771]), .Z(n10080) );
  NAND U12235 ( .A(x[507]), .B(y[7744]), .Z(n10081) );
  XNOR U12236 ( .A(n10080), .B(n10081), .Z(n10083) );
  AND U12237 ( .A(x[506]), .B(y[7745]), .Z(n10084) );
  XOR U12238 ( .A(o[91]), .B(n10084), .Z(n10082) );
  XOR U12239 ( .A(n10083), .B(n10082), .Z(n10018) );
  AND U12240 ( .A(x[489]), .B(y[7762]), .Z(n10087) );
  NAND U12241 ( .A(x[501]), .B(y[7750]), .Z(n10088) );
  XNOR U12242 ( .A(n10087), .B(n10088), .Z(n10089) );
  NAND U12243 ( .A(x[498]), .B(y[7753]), .Z(n10090) );
  XOR U12244 ( .A(n10089), .B(n10090), .Z(n10019) );
  XNOR U12245 ( .A(n10018), .B(n10019), .Z(n10020) );
  XOR U12246 ( .A(n10021), .B(n10020), .Z(n10009) );
  XNOR U12247 ( .A(n10008), .B(n10009), .Z(n10100) );
  XOR U12248 ( .A(n10099), .B(n10100), .Z(n10102) );
  XOR U12249 ( .A(n10101), .B(n10102), .Z(n10120) );
  NAND U12250 ( .A(n9870), .B(n9869), .Z(n9874) );
  NAND U12251 ( .A(n9872), .B(n9871), .Z(n9873) );
  AND U12252 ( .A(n9874), .B(n9873), .Z(n10118) );
  NAND U12253 ( .A(n9876), .B(n9875), .Z(n9880) );
  NANDN U12254 ( .A(n9878), .B(n9877), .Z(n9879) );
  AND U12255 ( .A(n9880), .B(n9879), .Z(n10117) );
  XOR U12256 ( .A(n10118), .B(n10117), .Z(n10119) );
  NANDN U12257 ( .A(n9882), .B(n9881), .Z(n9886) );
  NANDN U12258 ( .A(n9884), .B(n9883), .Z(n9885) );
  AND U12259 ( .A(n9886), .B(n9885), .Z(n10105) );
  NAND U12260 ( .A(n9888), .B(n9887), .Z(n9892) );
  NAND U12261 ( .A(n9890), .B(n9889), .Z(n9891) );
  NAND U12262 ( .A(n9892), .B(n9891), .Z(n10095) );
  NAND U12263 ( .A(n9894), .B(n9893), .Z(n9898) );
  NAND U12264 ( .A(n9896), .B(n9895), .Z(n9897) );
  NAND U12265 ( .A(n9898), .B(n9897), .Z(n10093) );
  AND U12266 ( .A(x[499]), .B(y[7752]), .Z(n10068) );
  NAND U12267 ( .A(x[505]), .B(y[7746]), .Z(n10069) );
  XNOR U12268 ( .A(n10068), .B(n10069), .Z(n10070) );
  NAND U12269 ( .A(x[486]), .B(y[7765]), .Z(n10071) );
  XNOR U12270 ( .A(n10070), .B(n10071), .Z(n10060) );
  AND U12271 ( .A(x[495]), .B(y[7756]), .Z(n10040) );
  AND U12272 ( .A(x[482]), .B(y[7769]), .Z(n10039) );
  XOR U12273 ( .A(n10040), .B(n10039), .Z(n10042) );
  AND U12274 ( .A(x[483]), .B(y[7768]), .Z(n10041) );
  XOR U12275 ( .A(n10042), .B(n10041), .Z(n10059) );
  XOR U12276 ( .A(n10060), .B(n10059), .Z(n10062) );
  NAND U12277 ( .A(x[496]), .B(y[7755]), .Z(n10024) );
  XOR U12278 ( .A(n10024), .B(n10025), .Z(n10027) );
  XNOR U12279 ( .A(n10026), .B(n10027), .Z(n10036) );
  AND U12280 ( .A(y[7758]), .B(x[493]), .Z(n9900) );
  NAND U12281 ( .A(y[7759]), .B(x[492]), .Z(n9899) );
  XNOR U12282 ( .A(n9900), .B(n9899), .Z(n10035) );
  XOR U12283 ( .A(n10036), .B(n10035), .Z(n10061) );
  XOR U12284 ( .A(n10062), .B(n10061), .Z(n10003) );
  NAND U12285 ( .A(n10034), .B(n9901), .Z(n9905) );
  ANDN U12286 ( .B(n9903), .A(n9902), .Z(n9904) );
  ANDN U12287 ( .B(n9905), .A(n9904), .Z(n10001) );
  NANDN U12288 ( .A(n9907), .B(n9906), .Z(n9911) );
  NAND U12289 ( .A(n9909), .B(n9908), .Z(n9910) );
  NAND U12290 ( .A(n9911), .B(n9910), .Z(n10000) );
  XNOR U12291 ( .A(n10001), .B(n10000), .Z(n10002) );
  XOR U12292 ( .A(n10003), .B(n10002), .Z(n10094) );
  XNOR U12293 ( .A(n10093), .B(n10094), .Z(n10096) );
  XNOR U12294 ( .A(n10105), .B(n10106), .Z(n10108) );
  NANDN U12295 ( .A(n9913), .B(n9912), .Z(n9917) );
  NANDN U12296 ( .A(n9915), .B(n9914), .Z(n9916) );
  AND U12297 ( .A(n9917), .B(n9916), .Z(n10107) );
  XOR U12298 ( .A(n10108), .B(n10107), .Z(n9982) );
  XOR U12299 ( .A(n9984), .B(n9985), .Z(n9991) );
  NAND U12300 ( .A(n9919), .B(n9918), .Z(n9923) );
  NAND U12301 ( .A(n9921), .B(n9920), .Z(n9922) );
  NAND U12302 ( .A(n9923), .B(n9922), .Z(n9988) );
  NANDN U12303 ( .A(n9925), .B(n9924), .Z(n9929) );
  NAND U12304 ( .A(n9927), .B(n9926), .Z(n9928) );
  NAND U12305 ( .A(n9929), .B(n9928), .Z(n9994) );
  NAND U12306 ( .A(n9931), .B(n9930), .Z(n9935) );
  NAND U12307 ( .A(n9933), .B(n9932), .Z(n9934) );
  AND U12308 ( .A(n9935), .B(n9934), .Z(n10113) );
  NANDN U12309 ( .A(n9937), .B(n9936), .Z(n9941) );
  NANDN U12310 ( .A(n9939), .B(n9938), .Z(n9940) );
  AND U12311 ( .A(n9941), .B(n9940), .Z(n10058) );
  AND U12312 ( .A(y[7747]), .B(x[504]), .Z(n9943) );
  NAND U12313 ( .A(y[7751]), .B(x[500]), .Z(n9942) );
  XNOR U12314 ( .A(n9943), .B(n9942), .Z(n10064) );
  NAND U12315 ( .A(x[487]), .B(y[7764]), .Z(n10065) );
  XNOR U12316 ( .A(n10064), .B(n10065), .Z(n10056) );
  AND U12317 ( .A(x[488]), .B(y[7763]), .Z(n10029) );
  AND U12318 ( .A(x[503]), .B(y[7748]), .Z(n10028) );
  XOR U12319 ( .A(n10029), .B(n10028), .Z(n10031) );
  AND U12320 ( .A(x[502]), .B(y[7749]), .Z(n10030) );
  XOR U12321 ( .A(n10031), .B(n10030), .Z(n10055) );
  XOR U12322 ( .A(n10056), .B(n10055), .Z(n10057) );
  XOR U12323 ( .A(n10058), .B(n10057), .Z(n10111) );
  NAND U12324 ( .A(n9945), .B(n9944), .Z(n9949) );
  ANDN U12325 ( .B(n9947), .A(n9946), .Z(n9948) );
  ANDN U12326 ( .B(n9949), .A(n9948), .Z(n10052) );
  NANDN U12327 ( .A(n9951), .B(n9950), .Z(n9955) );
  NANDN U12328 ( .A(n9953), .B(n9952), .Z(n9954) );
  NAND U12329 ( .A(n9955), .B(n9954), .Z(n10051) );
  XNOR U12330 ( .A(n10052), .B(n10051), .Z(n10054) );
  AND U12331 ( .A(x[488]), .B(y[7764]), .Z(n10086) );
  NAND U12332 ( .A(n9956), .B(n10086), .Z(n9960) );
  NANDN U12333 ( .A(n9958), .B(n9957), .Z(n9959) );
  NAND U12334 ( .A(n9960), .B(n9959), .Z(n10014) );
  AND U12335 ( .A(x[494]), .B(y[7757]), .Z(n10046) );
  AND U12336 ( .A(x[481]), .B(y[7770]), .Z(n10045) );
  XOR U12337 ( .A(n10046), .B(n10045), .Z(n10048) );
  ANDN U12338 ( .B(o[90]), .A(n9961), .Z(n10047) );
  XOR U12339 ( .A(n10048), .B(n10047), .Z(n10013) );
  AND U12340 ( .A(x[497]), .B(y[7754]), .Z(n10074) );
  NAND U12341 ( .A(x[484]), .B(y[7767]), .Z(n10075) );
  XNOR U12342 ( .A(n10074), .B(n10075), .Z(n10077) );
  AND U12343 ( .A(x[485]), .B(y[7766]), .Z(n10076) );
  XOR U12344 ( .A(n10077), .B(n10076), .Z(n10012) );
  XOR U12345 ( .A(n10013), .B(n10012), .Z(n10015) );
  XOR U12346 ( .A(n10014), .B(n10015), .Z(n10053) );
  XOR U12347 ( .A(n10054), .B(n10053), .Z(n10112) );
  XNOR U12348 ( .A(n10113), .B(n10114), .Z(n9995) );
  XOR U12349 ( .A(n9994), .B(n9995), .Z(n9997) );
  NAND U12350 ( .A(n9963), .B(n9962), .Z(n9967) );
  NAND U12351 ( .A(n9965), .B(n9964), .Z(n9966) );
  AND U12352 ( .A(n9967), .B(n9966), .Z(n9996) );
  XOR U12353 ( .A(n9997), .B(n9996), .Z(n9989) );
  XOR U12354 ( .A(n9988), .B(n9989), .Z(n9990) );
  XOR U12355 ( .A(n9970), .B(n9969), .Z(n9971) );
  XOR U12356 ( .A(n9972), .B(n9971), .Z(n9978) );
  XNOR U12357 ( .A(n9977), .B(n9978), .Z(n9968) );
  XOR U12358 ( .A(n9975), .B(n9968), .Z(N188) );
  NAND U12359 ( .A(n9970), .B(n9969), .Z(n9974) );
  NAND U12360 ( .A(n9972), .B(n9971), .Z(n9973) );
  NAND U12361 ( .A(n9974), .B(n9973), .Z(n10132) );
  IV U12362 ( .A(n10132), .Z(n10130) );
  OR U12363 ( .A(n9977), .B(n9975), .Z(n9981) );
  ANDN U12364 ( .B(n9977), .A(n9976), .Z(n9979) );
  OR U12365 ( .A(n9979), .B(n9978), .Z(n9980) );
  AND U12366 ( .A(n9981), .B(n9980), .Z(n10131) );
  NANDN U12367 ( .A(n9983), .B(n9982), .Z(n9987) );
  NAND U12368 ( .A(n9985), .B(n9984), .Z(n9986) );
  NAND U12369 ( .A(n9987), .B(n9986), .Z(n10124) );
  NAND U12370 ( .A(n9989), .B(n9988), .Z(n9993) );
  NANDN U12371 ( .A(n9991), .B(n9990), .Z(n9992) );
  AND U12372 ( .A(n9993), .B(n9992), .Z(n10125) );
  XOR U12373 ( .A(n10124), .B(n10125), .Z(n10127) );
  NAND U12374 ( .A(n9995), .B(n9994), .Z(n9999) );
  NAND U12375 ( .A(n9997), .B(n9996), .Z(n9998) );
  AND U12376 ( .A(n9999), .B(n9998), .Z(n10137) );
  NANDN U12377 ( .A(n10001), .B(n10000), .Z(n10005) );
  NAND U12378 ( .A(n10003), .B(n10002), .Z(n10004) );
  AND U12379 ( .A(n10005), .B(n10004), .Z(n10162) );
  NANDN U12380 ( .A(n10007), .B(n10006), .Z(n10011) );
  NANDN U12381 ( .A(n10009), .B(n10008), .Z(n10010) );
  AND U12382 ( .A(n10011), .B(n10010), .Z(n10263) );
  NAND U12383 ( .A(n10013), .B(n10012), .Z(n10017) );
  NAND U12384 ( .A(n10015), .B(n10014), .Z(n10016) );
  AND U12385 ( .A(n10017), .B(n10016), .Z(n10261) );
  NANDN U12386 ( .A(n10019), .B(n10018), .Z(n10023) );
  NANDN U12387 ( .A(n10021), .B(n10020), .Z(n10022) );
  NAND U12388 ( .A(n10023), .B(n10022), .Z(n10260) );
  XNOR U12389 ( .A(n10261), .B(n10260), .Z(n10262) );
  XNOR U12390 ( .A(n10263), .B(n10262), .Z(n10161) );
  XNOR U12391 ( .A(n10162), .B(n10161), .Z(n10164) );
  AND U12392 ( .A(x[495]), .B(y[7757]), .Z(n10239) );
  AND U12393 ( .A(x[507]), .B(y[7745]), .Z(n10223) );
  XOR U12394 ( .A(o[92]), .B(n10223), .Z(n10237) );
  AND U12395 ( .A(x[506]), .B(y[7746]), .Z(n10236) );
  XOR U12396 ( .A(n10237), .B(n10236), .Z(n10238) );
  XOR U12397 ( .A(n10239), .B(n10238), .Z(n10225) );
  AND U12398 ( .A(x[487]), .B(y[7765]), .Z(n10207) );
  AND U12399 ( .A(x[492]), .B(y[7760]), .Z(n10206) );
  XOR U12400 ( .A(n10207), .B(n10206), .Z(n10209) );
  AND U12401 ( .A(x[491]), .B(y[7761]), .Z(n10208) );
  XNOR U12402 ( .A(n10209), .B(n10208), .Z(n10224) );
  XOR U12403 ( .A(n10226), .B(n10227), .Z(n10267) );
  AND U12404 ( .A(x[497]), .B(y[7755]), .Z(n10172) );
  AND U12405 ( .A(x[502]), .B(y[7750]), .Z(n10171) );
  XOR U12406 ( .A(n10172), .B(n10171), .Z(n10174) );
  AND U12407 ( .A(x[484]), .B(y[7768]), .Z(n10173) );
  XOR U12408 ( .A(n10174), .B(n10173), .Z(n10245) );
  AND U12409 ( .A(x[486]), .B(y[7766]), .Z(n10386) );
  AND U12410 ( .A(x[499]), .B(y[7753]), .Z(n10212) );
  XOR U12411 ( .A(n10386), .B(n10212), .Z(n10214) );
  XOR U12412 ( .A(n10214), .B(n10213), .Z(n10244) );
  XOR U12413 ( .A(n10245), .B(n10244), .Z(n10247) );
  NAND U12414 ( .A(n10029), .B(n10028), .Z(n10033) );
  NAND U12415 ( .A(n10031), .B(n10030), .Z(n10032) );
  NAND U12416 ( .A(n10033), .B(n10032), .Z(n10246) );
  XOR U12417 ( .A(n10247), .B(n10246), .Z(n10266) );
  XOR U12418 ( .A(n10267), .B(n10266), .Z(n10269) );
  NAND U12419 ( .A(n10231), .B(n10034), .Z(n10038) );
  NAND U12420 ( .A(n10036), .B(n10035), .Z(n10037) );
  NAND U12421 ( .A(n10038), .B(n10037), .Z(n10190) );
  NAND U12422 ( .A(n10040), .B(n10039), .Z(n10044) );
  NAND U12423 ( .A(n10042), .B(n10041), .Z(n10043) );
  NAND U12424 ( .A(n10044), .B(n10043), .Z(n10189) );
  NAND U12425 ( .A(n10046), .B(n10045), .Z(n10050) );
  NAND U12426 ( .A(n10048), .B(n10047), .Z(n10049) );
  NAND U12427 ( .A(n10050), .B(n10049), .Z(n10188) );
  XOR U12428 ( .A(n10189), .B(n10188), .Z(n10191) );
  XOR U12429 ( .A(n10190), .B(n10191), .Z(n10268) );
  XOR U12430 ( .A(n10269), .B(n10268), .Z(n10163) );
  XNOR U12431 ( .A(n10164), .B(n10163), .Z(n10158) );
  XNOR U12432 ( .A(n10251), .B(n10250), .Z(n10252) );
  XOR U12433 ( .A(n10253), .B(n10252), .Z(n10155) );
  AND U12434 ( .A(x[504]), .B(y[7751]), .Z(n10573) );
  AND U12435 ( .A(x[500]), .B(y[7747]), .Z(n10063) );
  NAND U12436 ( .A(n10573), .B(n10063), .Z(n10067) );
  NANDN U12437 ( .A(n10065), .B(n10064), .Z(n10066) );
  NAND U12438 ( .A(n10067), .B(n10066), .Z(n10284) );
  AND U12439 ( .A(x[505]), .B(y[7747]), .Z(n10202) );
  XOR U12440 ( .A(n10203), .B(n10202), .Z(n10201) );
  AND U12441 ( .A(x[481]), .B(y[7771]), .Z(n10200) );
  XOR U12442 ( .A(n10201), .B(n10200), .Z(n10283) );
  AND U12443 ( .A(x[496]), .B(y[7756]), .Z(n10195) );
  AND U12444 ( .A(x[504]), .B(y[7748]), .Z(n10194) );
  XOR U12445 ( .A(n10195), .B(n10194), .Z(n10197) );
  AND U12446 ( .A(x[482]), .B(y[7770]), .Z(n10196) );
  XOR U12447 ( .A(n10197), .B(n10196), .Z(n10282) );
  XOR U12448 ( .A(n10283), .B(n10282), .Z(n10285) );
  XNOR U12449 ( .A(n10284), .B(n10285), .Z(n10258) );
  NANDN U12450 ( .A(n10069), .B(n10068), .Z(n10073) );
  NANDN U12451 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U12452 ( .A(n10073), .B(n10072), .Z(n10278) );
  AND U12453 ( .A(x[483]), .B(y[7769]), .Z(n10230) );
  XOR U12454 ( .A(n10231), .B(n10230), .Z(n10233) );
  AND U12455 ( .A(x[503]), .B(y[7749]), .Z(n10232) );
  XOR U12456 ( .A(n10233), .B(n10232), .Z(n10277) );
  AND U12457 ( .A(x[485]), .B(y[7767]), .Z(n10218) );
  AND U12458 ( .A(x[501]), .B(y[7751]), .Z(n10217) );
  XOR U12459 ( .A(n10218), .B(n10217), .Z(n10220) );
  AND U12460 ( .A(x[500]), .B(y[7752]), .Z(n10219) );
  XOR U12461 ( .A(n10220), .B(n10219), .Z(n10276) );
  XOR U12462 ( .A(n10277), .B(n10276), .Z(n10279) );
  XNOR U12463 ( .A(n10278), .B(n10279), .Z(n10256) );
  NANDN U12464 ( .A(n10075), .B(n10074), .Z(n10079) );
  NAND U12465 ( .A(n10077), .B(n10076), .Z(n10078) );
  NAND U12466 ( .A(n10079), .B(n10078), .Z(n10271) );
  XOR U12467 ( .A(n10271), .B(n10270), .Z(n10273) );
  AND U12468 ( .A(n10084), .B(o[91]), .Z(n10180) );
  AND U12469 ( .A(x[480]), .B(y[7772]), .Z(n10178) );
  AND U12470 ( .A(x[508]), .B(y[7744]), .Z(n10177) );
  XOR U12471 ( .A(n10178), .B(n10177), .Z(n10179) );
  XOR U12472 ( .A(n10180), .B(n10179), .Z(n10166) );
  NAND U12473 ( .A(y[7762]), .B(x[490]), .Z(n10085) );
  XNOR U12474 ( .A(n10086), .B(n10085), .Z(n10185) );
  AND U12475 ( .A(x[489]), .B(y[7763]), .Z(n10184) );
  XOR U12476 ( .A(n10185), .B(n10184), .Z(n10165) );
  XOR U12477 ( .A(n10166), .B(n10165), .Z(n10168) );
  NANDN U12478 ( .A(n10088), .B(n10087), .Z(n10092) );
  NANDN U12479 ( .A(n10090), .B(n10089), .Z(n10091) );
  NAND U12480 ( .A(n10092), .B(n10091), .Z(n10167) );
  XOR U12481 ( .A(n10168), .B(n10167), .Z(n10272) );
  XNOR U12482 ( .A(n10273), .B(n10272), .Z(n10257) );
  XOR U12483 ( .A(n10256), .B(n10257), .Z(n10259) );
  XOR U12484 ( .A(n10258), .B(n10259), .Z(n10156) );
  XOR U12485 ( .A(n10155), .B(n10156), .Z(n10157) );
  XNOR U12486 ( .A(n10158), .B(n10157), .Z(n10151) );
  NAND U12487 ( .A(n10094), .B(n10093), .Z(n10098) );
  NANDN U12488 ( .A(n10096), .B(n10095), .Z(n10097) );
  NAND U12489 ( .A(n10098), .B(n10097), .Z(n10150) );
  NAND U12490 ( .A(n10100), .B(n10099), .Z(n10104) );
  NAND U12491 ( .A(n10102), .B(n10101), .Z(n10103) );
  NAND U12492 ( .A(n10104), .B(n10103), .Z(n10149) );
  XNOR U12493 ( .A(n10150), .B(n10149), .Z(n10152) );
  XNOR U12494 ( .A(n10137), .B(n10138), .Z(n10140) );
  NANDN U12495 ( .A(n10106), .B(n10105), .Z(n10110) );
  NAND U12496 ( .A(n10108), .B(n10107), .Z(n10109) );
  NAND U12497 ( .A(n10110), .B(n10109), .Z(n10145) );
  NANDN U12498 ( .A(n10112), .B(n10111), .Z(n10116) );
  NANDN U12499 ( .A(n10114), .B(n10113), .Z(n10115) );
  AND U12500 ( .A(n10116), .B(n10115), .Z(n10144) );
  NAND U12501 ( .A(n10118), .B(n10117), .Z(n10122) );
  NANDN U12502 ( .A(n10120), .B(n10119), .Z(n10121) );
  AND U12503 ( .A(n10122), .B(n10121), .Z(n10143) );
  XOR U12504 ( .A(n10144), .B(n10143), .Z(n10146) );
  XOR U12505 ( .A(n10145), .B(n10146), .Z(n10139) );
  XOR U12506 ( .A(n10140), .B(n10139), .Z(n10126) );
  XOR U12507 ( .A(n10127), .B(n10126), .Z(n10133) );
  XNOR U12508 ( .A(n10131), .B(n10133), .Z(n10123) );
  XOR U12509 ( .A(n10130), .B(n10123), .Z(N189) );
  NAND U12510 ( .A(n10125), .B(n10124), .Z(n10129) );
  NAND U12511 ( .A(n10127), .B(n10126), .Z(n10128) );
  AND U12512 ( .A(n10129), .B(n10128), .Z(n10289) );
  NANDN U12513 ( .A(n10130), .B(n10131), .Z(n10136) );
  NOR U12514 ( .A(n10132), .B(n10131), .Z(n10134) );
  OR U12515 ( .A(n10134), .B(n10133), .Z(n10135) );
  AND U12516 ( .A(n10136), .B(n10135), .Z(n10290) );
  NANDN U12517 ( .A(n10138), .B(n10137), .Z(n10142) );
  NAND U12518 ( .A(n10140), .B(n10139), .Z(n10141) );
  NAND U12519 ( .A(n10142), .B(n10141), .Z(n10294) );
  NAND U12520 ( .A(n10144), .B(n10143), .Z(n10148) );
  NAND U12521 ( .A(n10146), .B(n10145), .Z(n10147) );
  NAND U12522 ( .A(n10148), .B(n10147), .Z(n10292) );
  NAND U12523 ( .A(n10150), .B(n10149), .Z(n10154) );
  NANDN U12524 ( .A(n10152), .B(n10151), .Z(n10153) );
  NAND U12525 ( .A(n10154), .B(n10153), .Z(n10298) );
  NAND U12526 ( .A(n10156), .B(n10155), .Z(n10160) );
  NAND U12527 ( .A(n10158), .B(n10157), .Z(n10159) );
  AND U12528 ( .A(n10160), .B(n10159), .Z(n10299) );
  XOR U12529 ( .A(n10298), .B(n10299), .Z(n10301) );
  NAND U12530 ( .A(n10166), .B(n10165), .Z(n10170) );
  NAND U12531 ( .A(n10168), .B(n10167), .Z(n10169) );
  AND U12532 ( .A(n10170), .B(n10169), .Z(n10417) );
  NAND U12533 ( .A(n10172), .B(n10171), .Z(n10176) );
  NAND U12534 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U12535 ( .A(n10176), .B(n10175), .Z(n10442) );
  NAND U12536 ( .A(n10178), .B(n10177), .Z(n10182) );
  NAND U12537 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U12538 ( .A(n10182), .B(n10181), .Z(n10441) );
  XOR U12539 ( .A(n10442), .B(n10441), .Z(n10443) );
  AND U12540 ( .A(y[7764]), .B(x[490]), .Z(n10460) );
  NAND U12541 ( .A(n10183), .B(n10460), .Z(n10187) );
  NAND U12542 ( .A(n10185), .B(n10184), .Z(n10186) );
  NAND U12543 ( .A(n10187), .B(n10186), .Z(n10425) );
  AND U12544 ( .A(x[502]), .B(y[7751]), .Z(n10364) );
  AND U12545 ( .A(x[492]), .B(y[7761]), .Z(n10522) );
  AND U12546 ( .A(x[481]), .B(y[7772]), .Z(n10362) );
  XOR U12547 ( .A(n10522), .B(n10362), .Z(n10363) );
  XOR U12548 ( .A(n10364), .B(n10363), .Z(n10424) );
  AND U12549 ( .A(x[495]), .B(y[7758]), .Z(n10367) );
  XOR U12550 ( .A(n10367), .B(n10651), .Z(n10369) );
  XOR U12551 ( .A(n10369), .B(n10368), .Z(n10423) );
  XOR U12552 ( .A(n10424), .B(n10423), .Z(n10426) );
  XNOR U12553 ( .A(n10425), .B(n10426), .Z(n10444) );
  NAND U12554 ( .A(n10189), .B(n10188), .Z(n10193) );
  NAND U12555 ( .A(n10191), .B(n10190), .Z(n10192) );
  AND U12556 ( .A(n10193), .B(n10192), .Z(n10419) );
  XOR U12557 ( .A(n10420), .B(n10419), .Z(n10414) );
  NAND U12558 ( .A(n10195), .B(n10194), .Z(n10199) );
  NAND U12559 ( .A(n10197), .B(n10196), .Z(n10198) );
  NAND U12560 ( .A(n10199), .B(n10198), .Z(n10430) );
  AND U12561 ( .A(n10201), .B(n10200), .Z(n10205) );
  NAND U12562 ( .A(n10203), .B(n10202), .Z(n10204) );
  NANDN U12563 ( .A(n10205), .B(n10204), .Z(n10429) );
  XOR U12564 ( .A(n10430), .B(n10429), .Z(n10431) );
  NAND U12565 ( .A(n10207), .B(n10206), .Z(n10211) );
  NAND U12566 ( .A(n10209), .B(n10208), .Z(n10210) );
  NAND U12567 ( .A(n10211), .B(n10210), .Z(n10328) );
  AND U12568 ( .A(x[491]), .B(y[7762]), .Z(n10383) );
  AND U12569 ( .A(x[483]), .B(y[7770]), .Z(n10381) );
  AND U12570 ( .A(x[497]), .B(y[7756]), .Z(n10380) );
  XOR U12571 ( .A(n10381), .B(n10380), .Z(n10382) );
  XOR U12572 ( .A(n10383), .B(n10382), .Z(n10327) );
  AND U12573 ( .A(x[503]), .B(y[7750]), .Z(n10377) );
  AND U12574 ( .A(x[493]), .B(y[7760]), .Z(n10375) );
  AND U12575 ( .A(x[504]), .B(y[7749]), .Z(n10555) );
  XOR U12576 ( .A(n10375), .B(n10555), .Z(n10376) );
  XOR U12577 ( .A(n10377), .B(n10376), .Z(n10326) );
  XOR U12578 ( .A(n10327), .B(n10326), .Z(n10329) );
  XNOR U12579 ( .A(n10328), .B(n10329), .Z(n10432) );
  NAND U12580 ( .A(n10386), .B(n10212), .Z(n10216) );
  NAND U12581 ( .A(n10214), .B(n10213), .Z(n10215) );
  NAND U12582 ( .A(n10216), .B(n10215), .Z(n10438) );
  AND U12583 ( .A(x[505]), .B(y[7748]), .Z(n10359) );
  AND U12584 ( .A(x[506]), .B(y[7747]), .Z(n10356) );
  XOR U12585 ( .A(n10357), .B(n10356), .Z(n10358) );
  XOR U12586 ( .A(n10359), .B(n10358), .Z(n10436) );
  AND U12587 ( .A(x[508]), .B(y[7745]), .Z(n10374) );
  XOR U12588 ( .A(o[93]), .B(n10374), .Z(n10455) );
  AND U12589 ( .A(x[480]), .B(y[7773]), .Z(n10453) );
  AND U12590 ( .A(x[509]), .B(y[7744]), .Z(n10452) );
  XOR U12591 ( .A(n10453), .B(n10452), .Z(n10454) );
  XNOR U12592 ( .A(n10455), .B(n10454), .Z(n10435) );
  XOR U12593 ( .A(n10438), .B(n10437), .Z(n10405) );
  NAND U12594 ( .A(n10218), .B(n10217), .Z(n10222) );
  NAND U12595 ( .A(n10220), .B(n10219), .Z(n10221) );
  NAND U12596 ( .A(n10222), .B(n10221), .Z(n10395) );
  AND U12597 ( .A(o[92]), .B(n10223), .Z(n10335) );
  AND U12598 ( .A(x[496]), .B(y[7757]), .Z(n10333) );
  AND U12599 ( .A(x[507]), .B(y[7746]), .Z(n10332) );
  XOR U12600 ( .A(n10333), .B(n10332), .Z(n10334) );
  XOR U12601 ( .A(n10335), .B(n10334), .Z(n10394) );
  AND U12602 ( .A(x[482]), .B(y[7771]), .Z(n10345) );
  XOR U12603 ( .A(n10345), .B(n10344), .Z(n10346) );
  XOR U12604 ( .A(n10347), .B(n10346), .Z(n10393) );
  XOR U12605 ( .A(n10394), .B(n10393), .Z(n10396) );
  XOR U12606 ( .A(n10395), .B(n10396), .Z(n10406) );
  NANDN U12607 ( .A(n10225), .B(n10224), .Z(n10229) );
  NANDN U12608 ( .A(n10227), .B(n10226), .Z(n10228) );
  NAND U12609 ( .A(n10229), .B(n10228), .Z(n10320) );
  NAND U12610 ( .A(n10231), .B(n10230), .Z(n10235) );
  NAND U12611 ( .A(n10233), .B(n10232), .Z(n10234) );
  NAND U12612 ( .A(n10235), .B(n10234), .Z(n10351) );
  NAND U12613 ( .A(n10237), .B(n10236), .Z(n10241) );
  NAND U12614 ( .A(n10239), .B(n10238), .Z(n10240) );
  NAND U12615 ( .A(n10241), .B(n10240), .Z(n10350) );
  XOR U12616 ( .A(n10351), .B(n10350), .Z(n10353) );
  AND U12617 ( .A(x[488]), .B(y[7765]), .Z(n10388) );
  AND U12618 ( .A(x[486]), .B(y[7767]), .Z(n10243) );
  AND U12619 ( .A(y[7766]), .B(x[487]), .Z(n10242) );
  XOR U12620 ( .A(n10243), .B(n10242), .Z(n10387) );
  XOR U12621 ( .A(n10388), .B(n10387), .Z(n10447) );
  AND U12622 ( .A(x[489]), .B(y[7764]), .Z(n10568) );
  XOR U12623 ( .A(n10447), .B(n10568), .Z(n10449) );
  AND U12624 ( .A(x[485]), .B(y[7768]), .Z(n10341) );
  AND U12625 ( .A(x[484]), .B(y[7769]), .Z(n10339) );
  AND U12626 ( .A(x[490]), .B(y[7763]), .Z(n10338) );
  XOR U12627 ( .A(n10339), .B(n10338), .Z(n10340) );
  XOR U12628 ( .A(n10341), .B(n10340), .Z(n10448) );
  XOR U12629 ( .A(n10449), .B(n10448), .Z(n10352) );
  XOR U12630 ( .A(n10353), .B(n10352), .Z(n10321) );
  XNOR U12631 ( .A(n10322), .B(n10323), .Z(n10412) );
  NAND U12632 ( .A(n10245), .B(n10244), .Z(n10249) );
  NAND U12633 ( .A(n10247), .B(n10246), .Z(n10248) );
  NAND U12634 ( .A(n10249), .B(n10248), .Z(n10411) );
  XNOR U12635 ( .A(n10309), .B(n10308), .Z(n10311) );
  NANDN U12636 ( .A(n10251), .B(n10250), .Z(n10255) );
  NANDN U12637 ( .A(n10253), .B(n10252), .Z(n10254) );
  AND U12638 ( .A(n10255), .B(n10254), .Z(n10305) );
  XNOR U12639 ( .A(n10305), .B(n10304), .Z(n10307) );
  NANDN U12640 ( .A(n10261), .B(n10260), .Z(n10265) );
  NANDN U12641 ( .A(n10263), .B(n10262), .Z(n10264) );
  NAND U12642 ( .A(n10265), .B(n10264), .Z(n10316) );
  NAND U12643 ( .A(n10271), .B(n10270), .Z(n10275) );
  NAND U12644 ( .A(n10273), .B(n10272), .Z(n10274) );
  NAND U12645 ( .A(n10275), .B(n10274), .Z(n10401) );
  NAND U12646 ( .A(n10277), .B(n10276), .Z(n10281) );
  NAND U12647 ( .A(n10279), .B(n10278), .Z(n10280) );
  NAND U12648 ( .A(n10281), .B(n10280), .Z(n10400) );
  NAND U12649 ( .A(n10283), .B(n10282), .Z(n10287) );
  NAND U12650 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U12651 ( .A(n10287), .B(n10286), .Z(n10399) );
  XOR U12652 ( .A(n10400), .B(n10399), .Z(n10402) );
  XOR U12653 ( .A(n10401), .B(n10402), .Z(n10315) );
  XOR U12654 ( .A(n10314), .B(n10315), .Z(n10317) );
  XOR U12655 ( .A(n10316), .B(n10317), .Z(n10306) );
  XOR U12656 ( .A(n10307), .B(n10306), .Z(n10310) );
  XOR U12657 ( .A(n10311), .B(n10310), .Z(n10300) );
  XOR U12658 ( .A(n10301), .B(n10300), .Z(n10293) );
  XOR U12659 ( .A(n10292), .B(n10293), .Z(n10295) );
  XOR U12660 ( .A(n10294), .B(n10295), .Z(n10291) );
  XNOR U12661 ( .A(n10290), .B(n10291), .Z(n10288) );
  XOR U12662 ( .A(n10289), .B(n10288), .Z(N190) );
  NAND U12663 ( .A(n10293), .B(n10292), .Z(n10297) );
  NAND U12664 ( .A(n10295), .B(n10294), .Z(n10296) );
  AND U12665 ( .A(n10297), .B(n10296), .Z(n10723) );
  XNOR U12666 ( .A(n10724), .B(n10723), .Z(n10722) );
  NAND U12667 ( .A(n10299), .B(n10298), .Z(n10303) );
  NAND U12668 ( .A(n10301), .B(n10300), .Z(n10302) );
  NAND U12669 ( .A(n10303), .B(n10302), .Z(n10742) );
  NANDN U12670 ( .A(n10309), .B(n10308), .Z(n10313) );
  NAND U12671 ( .A(n10311), .B(n10310), .Z(n10312) );
  NAND U12672 ( .A(n10313), .B(n10312), .Z(n10465) );
  NAND U12673 ( .A(n10315), .B(n10314), .Z(n10319) );
  NAND U12674 ( .A(n10317), .B(n10316), .Z(n10318) );
  NAND U12675 ( .A(n10319), .B(n10318), .Z(n10463) );
  XOR U12676 ( .A(n10462), .B(n10463), .Z(n10740) );
  NANDN U12677 ( .A(n10321), .B(n10320), .Z(n10325) );
  NANDN U12678 ( .A(n10323), .B(n10322), .Z(n10324) );
  AND U12679 ( .A(n10325), .B(n10324), .Z(n10710) );
  NAND U12680 ( .A(n10327), .B(n10326), .Z(n10331) );
  NAND U12681 ( .A(n10329), .B(n10328), .Z(n10330) );
  AND U12682 ( .A(n10331), .B(n10330), .Z(n10471) );
  NAND U12683 ( .A(n10333), .B(n10332), .Z(n10337) );
  NAND U12684 ( .A(n10335), .B(n10334), .Z(n10336) );
  NAND U12685 ( .A(n10337), .B(n10336), .Z(n10480) );
  NAND U12686 ( .A(n10339), .B(n10338), .Z(n10343) );
  NAND U12687 ( .A(n10341), .B(n10340), .Z(n10342) );
  NAND U12688 ( .A(n10343), .B(n10342), .Z(n10483) );
  AND U12689 ( .A(x[486]), .B(y[7768]), .Z(n10559) );
  AND U12690 ( .A(x[485]), .B(y[7769]), .Z(n10561) );
  AND U12691 ( .A(x[499]), .B(y[7755]), .Z(n10560) );
  XOR U12692 ( .A(n10561), .B(n10560), .Z(n10558) );
  XNOR U12693 ( .A(n10559), .B(n10558), .Z(n10484) );
  AND U12694 ( .A(x[484]), .B(y[7770]), .Z(n10517) );
  AND U12695 ( .A(x[483]), .B(y[7771]), .Z(n10519) );
  AND U12696 ( .A(x[498]), .B(y[7756]), .Z(n10518) );
  XOR U12697 ( .A(n10519), .B(n10518), .Z(n10516) );
  XOR U12698 ( .A(n10517), .B(n10516), .Z(n10487) );
  NAND U12699 ( .A(n10345), .B(n10344), .Z(n10349) );
  NAND U12700 ( .A(n10347), .B(n10346), .Z(n10348) );
  AND U12701 ( .A(n10349), .B(n10348), .Z(n10486) );
  XOR U12702 ( .A(n10484), .B(n10485), .Z(n10482) );
  XOR U12703 ( .A(n10483), .B(n10482), .Z(n10481) );
  XOR U12704 ( .A(n10480), .B(n10481), .Z(n10470) );
  NAND U12705 ( .A(n10351), .B(n10350), .Z(n10355) );
  NAND U12706 ( .A(n10353), .B(n10352), .Z(n10354) );
  AND U12707 ( .A(n10355), .B(n10354), .Z(n10469) );
  XNOR U12708 ( .A(n10468), .B(n10469), .Z(n10712) );
  NAND U12709 ( .A(n10357), .B(n10356), .Z(n10361) );
  AND U12710 ( .A(n10359), .B(n10358), .Z(n10360) );
  ANDN U12711 ( .B(n10361), .A(n10360), .Z(n10505) );
  NAND U12712 ( .A(n10522), .B(n10362), .Z(n10366) );
  AND U12713 ( .A(n10364), .B(n10363), .Z(n10365) );
  ANDN U12714 ( .B(n10366), .A(n10365), .Z(n10507) );
  NAND U12715 ( .A(n10367), .B(n10651), .Z(n10371) );
  NAND U12716 ( .A(n10369), .B(n10368), .Z(n10370) );
  AND U12717 ( .A(n10371), .B(n10370), .Z(n10667) );
  AND U12718 ( .A(x[503]), .B(y[7751]), .Z(n10554) );
  AND U12719 ( .A(y[7750]), .B(x[504]), .Z(n10373) );
  AND U12720 ( .A(y[7749]), .B(x[505]), .Z(n10372) );
  XOR U12721 ( .A(n10373), .B(n10372), .Z(n10553) );
  XOR U12722 ( .A(n10554), .B(n10553), .Z(n10669) );
  AND U12723 ( .A(n10374), .B(o[93]), .Z(n10513) );
  AND U12724 ( .A(x[508]), .B(y[7746]), .Z(n10511) );
  AND U12725 ( .A(x[496]), .B(y[7758]), .Z(n10510) );
  XOR U12726 ( .A(n10511), .B(n10510), .Z(n10512) );
  XNOR U12727 ( .A(n10513), .B(n10512), .Z(n10668) );
  XNOR U12728 ( .A(n10667), .B(n10666), .Z(n10506) );
  XNOR U12729 ( .A(n10505), .B(n10504), .Z(n10697) );
  NAND U12730 ( .A(n10375), .B(n10555), .Z(n10379) );
  NAND U12731 ( .A(n10377), .B(n10376), .Z(n10378) );
  AND U12732 ( .A(n10379), .B(n10378), .Z(n10477) );
  NAND U12733 ( .A(n10381), .B(n10380), .Z(n10385) );
  NAND U12734 ( .A(n10383), .B(n10382), .Z(n10384) );
  AND U12735 ( .A(n10385), .B(n10384), .Z(n10661) );
  AND U12736 ( .A(x[480]), .B(y[7774]), .Z(n10548) );
  AND U12737 ( .A(x[509]), .B(y[7745]), .Z(n10571) );
  XOR U12738 ( .A(o[94]), .B(n10571), .Z(n10550) );
  AND U12739 ( .A(x[510]), .B(y[7744]), .Z(n10549) );
  XOR U12740 ( .A(n10550), .B(n10549), .Z(n10547) );
  XOR U12741 ( .A(n10548), .B(n10547), .Z(n10663) );
  AND U12742 ( .A(x[500]), .B(y[7754]), .Z(n10636) );
  XOR U12743 ( .A(n10637), .B(n10636), .Z(n10635) );
  AND U12744 ( .A(x[488]), .B(y[7766]), .Z(n10634) );
  XNOR U12745 ( .A(n10635), .B(n10634), .Z(n10662) );
  XNOR U12746 ( .A(n10661), .B(n10660), .Z(n10476) );
  AND U12747 ( .A(x[487]), .B(y[7767]), .Z(n10649) );
  NAND U12748 ( .A(n10386), .B(n10649), .Z(n10390) );
  NAND U12749 ( .A(n10388), .B(n10387), .Z(n10389) );
  AND U12750 ( .A(n10390), .B(n10389), .Z(n10497) );
  AND U12751 ( .A(y[7753]), .B(x[501]), .Z(n10392) );
  AND U12752 ( .A(y[7752]), .B(x[502]), .Z(n10391) );
  XOR U12753 ( .A(n10392), .B(n10391), .Z(n10648) );
  XOR U12754 ( .A(n10649), .B(n10648), .Z(n10499) );
  AND U12755 ( .A(x[497]), .B(y[7757]), .Z(n10629) );
  AND U12756 ( .A(x[482]), .B(y[7772]), .Z(n10631) );
  AND U12757 ( .A(x[506]), .B(y[7748]), .Z(n10630) );
  XOR U12758 ( .A(n10631), .B(n10630), .Z(n10628) );
  XNOR U12759 ( .A(n10629), .B(n10628), .Z(n10498) );
  XOR U12760 ( .A(n10497), .B(n10496), .Z(n10475) );
  XNOR U12761 ( .A(n10474), .B(n10475), .Z(n10699) );
  NAND U12762 ( .A(n10394), .B(n10393), .Z(n10398) );
  NAND U12763 ( .A(n10396), .B(n10395), .Z(n10397) );
  AND U12764 ( .A(n10398), .B(n10397), .Z(n10700) );
  XOR U12765 ( .A(n10697), .B(n10696), .Z(n10711) );
  XOR U12766 ( .A(n10712), .B(n10711), .Z(n10709) );
  XOR U12767 ( .A(n10710), .B(n10709), .Z(n10704) );
  NAND U12768 ( .A(n10400), .B(n10399), .Z(n10404) );
  NAND U12769 ( .A(n10402), .B(n10401), .Z(n10403) );
  AND U12770 ( .A(n10404), .B(n10403), .Z(n10705) );
  NANDN U12771 ( .A(n10406), .B(n10405), .Z(n10410) );
  NANDN U12772 ( .A(n10408), .B(n10407), .Z(n10409) );
  AND U12773 ( .A(n10410), .B(n10409), .Z(n10706) );
  XOR U12774 ( .A(n10704), .B(n10703), .Z(n10727) );
  NANDN U12775 ( .A(n10412), .B(n10411), .Z(n10416) );
  NANDN U12776 ( .A(n10414), .B(n10413), .Z(n10415) );
  AND U12777 ( .A(n10416), .B(n10415), .Z(n10730) );
  NANDN U12778 ( .A(n10418), .B(n10417), .Z(n10422) );
  NAND U12779 ( .A(n10420), .B(n10419), .Z(n10421) );
  AND U12780 ( .A(n10422), .B(n10421), .Z(n10693) );
  NAND U12781 ( .A(n10424), .B(n10423), .Z(n10428) );
  NAND U12782 ( .A(n10426), .B(n10425), .Z(n10427) );
  AND U12783 ( .A(n10428), .B(n10427), .Z(n10688) );
  NAND U12784 ( .A(n10430), .B(n10429), .Z(n10434) );
  NANDN U12785 ( .A(n10432), .B(n10431), .Z(n10433) );
  NAND U12786 ( .A(n10434), .B(n10433), .Z(n10689) );
  NANDN U12787 ( .A(n10436), .B(n10435), .Z(n10440) );
  OR U12788 ( .A(n10438), .B(n10437), .Z(n10439) );
  NAND U12789 ( .A(n10440), .B(n10439), .Z(n10686) );
  XOR U12790 ( .A(n10687), .B(n10686), .Z(n10695) );
  NAND U12791 ( .A(n10442), .B(n10441), .Z(n10446) );
  NANDN U12792 ( .A(n10444), .B(n10443), .Z(n10445) );
  AND U12793 ( .A(n10446), .B(n10445), .Z(n10681) );
  NAND U12794 ( .A(n10447), .B(n10568), .Z(n10451) );
  NAND U12795 ( .A(n10449), .B(n10448), .Z(n10450) );
  AND U12796 ( .A(n10451), .B(n10450), .Z(n10683) );
  NAND U12797 ( .A(n10453), .B(n10452), .Z(n10457) );
  NAND U12798 ( .A(n10455), .B(n10454), .Z(n10456) );
  AND U12799 ( .A(n10457), .B(n10456), .Z(n10491) );
  AND U12800 ( .A(y[7762]), .B(x[492]), .Z(n10458) );
  XOR U12801 ( .A(n10459), .B(n10458), .Z(n10523) );
  XOR U12802 ( .A(n10524), .B(n10523), .Z(n10567) );
  AND U12803 ( .A(y[7765]), .B(x[489]), .Z(n10461) );
  XOR U12804 ( .A(n10461), .B(n10460), .Z(n10566) );
  XOR U12805 ( .A(n10567), .B(n10566), .Z(n10493) );
  AND U12806 ( .A(x[507]), .B(y[7747]), .Z(n10645) );
  AND U12807 ( .A(x[481]), .B(y[7773]), .Z(n10644) );
  XOR U12808 ( .A(n10645), .B(n10644), .Z(n10642) );
  XOR U12809 ( .A(n10643), .B(n10642), .Z(n10492) );
  XOR U12810 ( .A(n10493), .B(n10492), .Z(n10490) );
  XOR U12811 ( .A(n10491), .B(n10490), .Z(n10682) );
  XOR U12812 ( .A(n10683), .B(n10682), .Z(n10680) );
  XNOR U12813 ( .A(n10681), .B(n10680), .Z(n10694) );
  XOR U12814 ( .A(n10693), .B(n10692), .Z(n10729) );
  XOR U12815 ( .A(n10727), .B(n10728), .Z(n10739) );
  XOR U12816 ( .A(n10740), .B(n10739), .Z(n10741) );
  XOR U12817 ( .A(n10742), .B(n10741), .Z(n10721) );
  XNOR U12818 ( .A(n10722), .B(n10721), .Z(N191) );
  NANDN U12819 ( .A(n10463), .B(n10462), .Z(n10467) );
  NANDN U12820 ( .A(n10465), .B(n10464), .Z(n10466) );
  AND U12821 ( .A(n10467), .B(n10466), .Z(n10738) );
  NANDN U12822 ( .A(n10469), .B(n10468), .Z(n10473) );
  NANDN U12823 ( .A(n10471), .B(n10470), .Z(n10472) );
  AND U12824 ( .A(n10473), .B(n10472), .Z(n10720) );
  NANDN U12825 ( .A(n10475), .B(n10474), .Z(n10479) );
  NANDN U12826 ( .A(n10477), .B(n10476), .Z(n10478) );
  AND U12827 ( .A(n10479), .B(n10478), .Z(n10702) );
  NANDN U12828 ( .A(n10485), .B(n10484), .Z(n10489) );
  NANDN U12829 ( .A(n10487), .B(n10486), .Z(n10488) );
  NANDN U12830 ( .A(n10491), .B(n10490), .Z(n10495) );
  NAND U12831 ( .A(n10493), .B(n10492), .Z(n10494) );
  AND U12832 ( .A(n10495), .B(n10494), .Z(n10503) );
  NAND U12833 ( .A(n10497), .B(n10496), .Z(n10501) );
  NANDN U12834 ( .A(n10499), .B(n10498), .Z(n10500) );
  NAND U12835 ( .A(n10501), .B(n10500), .Z(n10502) );
  XNOR U12836 ( .A(n10503), .B(n10502), .Z(n10679) );
  NANDN U12837 ( .A(n10505), .B(n10504), .Z(n10509) );
  NANDN U12838 ( .A(n10507), .B(n10506), .Z(n10508) );
  AND U12839 ( .A(n10509), .B(n10508), .Z(n10677) );
  AND U12840 ( .A(n10511), .B(n10510), .Z(n10515) );
  AND U12841 ( .A(n10513), .B(n10512), .Z(n10514) );
  NOR U12842 ( .A(n10515), .B(n10514), .Z(n10546) );
  NAND U12843 ( .A(n10517), .B(n10516), .Z(n10521) );
  NAND U12844 ( .A(n10519), .B(n10518), .Z(n10520) );
  AND U12845 ( .A(n10521), .B(n10520), .Z(n10528) );
  NAND U12846 ( .A(n10522), .B(n10591), .Z(n10526) );
  NAND U12847 ( .A(n10524), .B(n10523), .Z(n10525) );
  AND U12848 ( .A(n10526), .B(n10525), .Z(n10527) );
  XNOR U12849 ( .A(n10528), .B(n10527), .Z(n10544) );
  AND U12850 ( .A(y[7744]), .B(x[511]), .Z(n10530) );
  NAND U12851 ( .A(y[7768]), .B(x[487]), .Z(n10529) );
  XNOR U12852 ( .A(n10530), .B(n10529), .Z(n10534) );
  AND U12853 ( .A(y[7748]), .B(x[507]), .Z(n10532) );
  NAND U12854 ( .A(y[7758]), .B(x[497]), .Z(n10531) );
  XNOR U12855 ( .A(n10532), .B(n10531), .Z(n10533) );
  XOR U12856 ( .A(n10534), .B(n10533), .Z(n10542) );
  AND U12857 ( .A(y[7769]), .B(x[486]), .Z(n10536) );
  NAND U12858 ( .A(y[7772]), .B(x[483]), .Z(n10535) );
  XNOR U12859 ( .A(n10536), .B(n10535), .Z(n10540) );
  AND U12860 ( .A(y[7770]), .B(x[485]), .Z(n10538) );
  NAND U12861 ( .A(y[7773]), .B(x[482]), .Z(n10537) );
  XNOR U12862 ( .A(n10538), .B(n10537), .Z(n10539) );
  XNOR U12863 ( .A(n10540), .B(n10539), .Z(n10541) );
  XNOR U12864 ( .A(n10542), .B(n10541), .Z(n10543) );
  XOR U12865 ( .A(n10544), .B(n10543), .Z(n10545) );
  XNOR U12866 ( .A(n10546), .B(n10545), .Z(n10627) );
  NAND U12867 ( .A(n10548), .B(n10547), .Z(n10552) );
  NAND U12868 ( .A(n10550), .B(n10549), .Z(n10551) );
  AND U12869 ( .A(n10552), .B(n10551), .Z(n10625) );
  NAND U12870 ( .A(n10554), .B(n10553), .Z(n10557) );
  AND U12871 ( .A(x[505]), .B(y[7750]), .Z(n10572) );
  NAND U12872 ( .A(n10555), .B(n10572), .Z(n10556) );
  AND U12873 ( .A(n10557), .B(n10556), .Z(n10565) );
  NAND U12874 ( .A(n10559), .B(n10558), .Z(n10563) );
  NAND U12875 ( .A(n10561), .B(n10560), .Z(n10562) );
  NAND U12876 ( .A(n10563), .B(n10562), .Z(n10564) );
  XNOR U12877 ( .A(n10565), .B(n10564), .Z(n10623) );
  NAND U12878 ( .A(n10567), .B(n10566), .Z(n10570) );
  AND U12879 ( .A(x[490]), .B(y[7765]), .Z(n10590) );
  NAND U12880 ( .A(n10568), .B(n10590), .Z(n10569) );
  AND U12881 ( .A(n10570), .B(n10569), .Z(n10621) );
  AND U12882 ( .A(y[7757]), .B(x[498]), .Z(n10579) );
  AND U12883 ( .A(n10571), .B(o[94]), .Z(n10577) );
  AND U12884 ( .A(x[502]), .B(y[7753]), .Z(n10650) );
  XOR U12885 ( .A(n10650), .B(o[95]), .Z(n10575) );
  XNOR U12886 ( .A(n10573), .B(n10572), .Z(n10574) );
  XNOR U12887 ( .A(n10575), .B(n10574), .Z(n10576) );
  XNOR U12888 ( .A(n10577), .B(n10576), .Z(n10578) );
  XNOR U12889 ( .A(n10579), .B(n10578), .Z(n10619) );
  AND U12890 ( .A(y[7774]), .B(x[481]), .Z(n10581) );
  NAND U12891 ( .A(y[7747]), .B(x[508]), .Z(n10580) );
  XNOR U12892 ( .A(n10581), .B(n10580), .Z(n10589) );
  AND U12893 ( .A(y[7775]), .B(x[480]), .Z(n10587) );
  AND U12894 ( .A(y[7764]), .B(x[491]), .Z(n10583) );
  NAND U12895 ( .A(y[7763]), .B(x[492]), .Z(n10582) );
  XNOR U12896 ( .A(n10583), .B(n10582), .Z(n10584) );
  XNOR U12897 ( .A(n10585), .B(n10584), .Z(n10586) );
  XNOR U12898 ( .A(n10587), .B(n10586), .Z(n10588) );
  XOR U12899 ( .A(n10589), .B(n10588), .Z(n10593) );
  XNOR U12900 ( .A(n10591), .B(n10590), .Z(n10592) );
  XNOR U12901 ( .A(n10593), .B(n10592), .Z(n10609) );
  AND U12902 ( .A(y[7745]), .B(x[510]), .Z(n10595) );
  NAND U12903 ( .A(y[7759]), .B(x[496]), .Z(n10594) );
  XNOR U12904 ( .A(n10595), .B(n10594), .Z(n10599) );
  AND U12905 ( .A(y[7752]), .B(x[503]), .Z(n10597) );
  NAND U12906 ( .A(y[7755]), .B(x[500]), .Z(n10596) );
  XNOR U12907 ( .A(n10597), .B(n10596), .Z(n10598) );
  XOR U12908 ( .A(n10599), .B(n10598), .Z(n10607) );
  AND U12909 ( .A(y[7761]), .B(x[494]), .Z(n10601) );
  NAND U12910 ( .A(y[7749]), .B(x[506]), .Z(n10600) );
  XNOR U12911 ( .A(n10601), .B(n10600), .Z(n10605) );
  AND U12912 ( .A(y[7746]), .B(x[509]), .Z(n10603) );
  NAND U12913 ( .A(y[7766]), .B(x[489]), .Z(n10602) );
  XNOR U12914 ( .A(n10603), .B(n10602), .Z(n10604) );
  XNOR U12915 ( .A(n10605), .B(n10604), .Z(n10606) );
  XNOR U12916 ( .A(n10607), .B(n10606), .Z(n10608) );
  XOR U12917 ( .A(n10609), .B(n10608), .Z(n10617) );
  AND U12918 ( .A(y[7756]), .B(x[499]), .Z(n10611) );
  NAND U12919 ( .A(y[7771]), .B(x[484]), .Z(n10610) );
  XNOR U12920 ( .A(n10611), .B(n10610), .Z(n10615) );
  AND U12921 ( .A(y[7754]), .B(x[501]), .Z(n10613) );
  NAND U12922 ( .A(y[7767]), .B(x[488]), .Z(n10612) );
  XNOR U12923 ( .A(n10613), .B(n10612), .Z(n10614) );
  XNOR U12924 ( .A(n10615), .B(n10614), .Z(n10616) );
  XNOR U12925 ( .A(n10617), .B(n10616), .Z(n10618) );
  XNOR U12926 ( .A(n10619), .B(n10618), .Z(n10620) );
  XNOR U12927 ( .A(n10621), .B(n10620), .Z(n10622) );
  XNOR U12928 ( .A(n10623), .B(n10622), .Z(n10624) );
  XNOR U12929 ( .A(n10625), .B(n10624), .Z(n10626) );
  XOR U12930 ( .A(n10627), .B(n10626), .Z(n10659) );
  NAND U12931 ( .A(n10629), .B(n10628), .Z(n10633) );
  NAND U12932 ( .A(n10631), .B(n10630), .Z(n10632) );
  AND U12933 ( .A(n10633), .B(n10632), .Z(n10641) );
  NAND U12934 ( .A(n10635), .B(n10634), .Z(n10639) );
  NAND U12935 ( .A(n10637), .B(n10636), .Z(n10638) );
  NAND U12936 ( .A(n10639), .B(n10638), .Z(n10640) );
  XNOR U12937 ( .A(n10641), .B(n10640), .Z(n10657) );
  NAND U12938 ( .A(n10643), .B(n10642), .Z(n10647) );
  NAND U12939 ( .A(n10645), .B(n10644), .Z(n10646) );
  AND U12940 ( .A(n10647), .B(n10646), .Z(n10655) );
  NAND U12941 ( .A(n10649), .B(n10648), .Z(n10653) );
  NAND U12942 ( .A(n10651), .B(n10650), .Z(n10652) );
  NAND U12943 ( .A(n10653), .B(n10652), .Z(n10654) );
  XNOR U12944 ( .A(n10655), .B(n10654), .Z(n10656) );
  XNOR U12945 ( .A(n10657), .B(n10656), .Z(n10658) );
  XNOR U12946 ( .A(n10659), .B(n10658), .Z(n10675) );
  NAND U12947 ( .A(n10661), .B(n10660), .Z(n10665) );
  NANDN U12948 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U12949 ( .A(n10665), .B(n10664), .Z(n10673) );
  NAND U12950 ( .A(n10667), .B(n10666), .Z(n10671) );
  NANDN U12951 ( .A(n10669), .B(n10668), .Z(n10670) );
  NAND U12952 ( .A(n10671), .B(n10670), .Z(n10672) );
  XNOR U12953 ( .A(n10673), .B(n10672), .Z(n10674) );
  XNOR U12954 ( .A(n10675), .B(n10674), .Z(n10676) );
  XNOR U12955 ( .A(n10677), .B(n10676), .Z(n10678) );
  NAND U12956 ( .A(n10681), .B(n10680), .Z(n10685) );
  NAND U12957 ( .A(n10683), .B(n10682), .Z(n10684) );
  NAND U12958 ( .A(n10687), .B(n10686), .Z(n10691) );
  NANDN U12959 ( .A(n10689), .B(n10688), .Z(n10690) );
  IV U12960 ( .A(n10696), .Z(n10698) );
  XNOR U12961 ( .A(n10702), .B(n10701), .Z(n10718) );
  NANDN U12962 ( .A(n10704), .B(n10703), .Z(n10708) );
  NANDN U12963 ( .A(n10706), .B(n10705), .Z(n10707) );
  AND U12964 ( .A(n10708), .B(n10707), .Z(n10716) );
  NAND U12965 ( .A(n10710), .B(n10709), .Z(n10714) );
  NAND U12966 ( .A(n10712), .B(n10711), .Z(n10713) );
  NAND U12967 ( .A(n10714), .B(n10713), .Z(n10715) );
  XNOR U12968 ( .A(n10716), .B(n10715), .Z(n10717) );
  XNOR U12969 ( .A(n10718), .B(n10717), .Z(n10719) );
  XNOR U12970 ( .A(n10720), .B(n10719), .Z(n10736) );
  NAND U12971 ( .A(n10722), .B(n10721), .Z(n10726) );
  NANDN U12972 ( .A(n10724), .B(n10723), .Z(n10725) );
  AND U12973 ( .A(n10726), .B(n10725), .Z(n10734) );
  NANDN U12974 ( .A(n10728), .B(n10727), .Z(n10732) );
  NANDN U12975 ( .A(n10730), .B(n10729), .Z(n10731) );
  NAND U12976 ( .A(n10732), .B(n10731), .Z(n10733) );
  XNOR U12977 ( .A(n10734), .B(n10733), .Z(n10735) );
  XNOR U12978 ( .A(n10736), .B(n10735), .Z(n10737) );
  XNOR U12979 ( .A(n10738), .B(n10737), .Z(n10746) );
  ANDN U12980 ( .B(n10740), .A(n10739), .Z(n10744) );
  ANDN U12981 ( .B(n10742), .A(n10741), .Z(n10743) );
  NOR U12982 ( .A(n10744), .B(n10743), .Z(n10745) );
  XNOR U12983 ( .A(n10746), .B(n10745), .Z(N192) );
  AND U12984 ( .A(x[480]), .B(y[7776]), .Z(n11395) );
  XOR U12985 ( .A(n11395), .B(o[96]), .Z(N225) );
  AND U12986 ( .A(x[481]), .B(y[7776]), .Z(n10755) );
  AND U12987 ( .A(x[480]), .B(y[7777]), .Z(n10754) );
  XNOR U12988 ( .A(n10754), .B(o[97]), .Z(n10747) );
  XNOR U12989 ( .A(n10755), .B(n10747), .Z(n10749) );
  NAND U12990 ( .A(n11395), .B(o[96]), .Z(n10748) );
  XNOR U12991 ( .A(n10749), .B(n10748), .Z(N226) );
  NANDN U12992 ( .A(n10755), .B(n10747), .Z(n10751) );
  NAND U12993 ( .A(n10749), .B(n10748), .Z(n10750) );
  AND U12994 ( .A(n10751), .B(n10750), .Z(n10761) );
  AND U12995 ( .A(x[480]), .B(y[7778]), .Z(n10768) );
  XNOR U12996 ( .A(n10768), .B(o[98]), .Z(n10760) );
  XNOR U12997 ( .A(n10761), .B(n10760), .Z(n10763) );
  AND U12998 ( .A(y[7776]), .B(x[482]), .Z(n10753) );
  NAND U12999 ( .A(y[7777]), .B(x[481]), .Z(n10752) );
  XNOR U13000 ( .A(n10753), .B(n10752), .Z(n10757) );
  AND U13001 ( .A(n10754), .B(o[97]), .Z(n10756) );
  XNOR U13002 ( .A(n10757), .B(n10756), .Z(n10762) );
  XNOR U13003 ( .A(n10763), .B(n10762), .Z(N227) );
  AND U13004 ( .A(x[482]), .B(y[7777]), .Z(n10775) );
  NAND U13005 ( .A(n10775), .B(n10755), .Z(n10759) );
  NAND U13006 ( .A(n10757), .B(n10756), .Z(n10758) );
  AND U13007 ( .A(n10759), .B(n10758), .Z(n10778) );
  NANDN U13008 ( .A(n10761), .B(n10760), .Z(n10765) );
  NAND U13009 ( .A(n10763), .B(n10762), .Z(n10764) );
  AND U13010 ( .A(n10765), .B(n10764), .Z(n10777) );
  XNOR U13011 ( .A(n10778), .B(n10777), .Z(n10780) );
  AND U13012 ( .A(x[481]), .B(y[7778]), .Z(n10893) );
  XOR U13013 ( .A(n10775), .B(o[99]), .Z(n10783) );
  XOR U13014 ( .A(n10893), .B(n10783), .Z(n10785) );
  AND U13015 ( .A(y[7776]), .B(x[483]), .Z(n10767) );
  NAND U13016 ( .A(y[7779]), .B(x[480]), .Z(n10766) );
  XNOR U13017 ( .A(n10767), .B(n10766), .Z(n10770) );
  AND U13018 ( .A(n10768), .B(o[98]), .Z(n10769) );
  XOR U13019 ( .A(n10770), .B(n10769), .Z(n10784) );
  XOR U13020 ( .A(n10785), .B(n10784), .Z(n10779) );
  XOR U13021 ( .A(n10780), .B(n10779), .Z(N228) );
  AND U13022 ( .A(x[483]), .B(y[7779]), .Z(n10828) );
  NAND U13023 ( .A(n11395), .B(n10828), .Z(n10772) );
  NAND U13024 ( .A(n10770), .B(n10769), .Z(n10771) );
  NAND U13025 ( .A(n10772), .B(n10771), .Z(n10806) );
  AND U13026 ( .A(y[7780]), .B(x[480]), .Z(n10774) );
  NAND U13027 ( .A(y[7776]), .B(x[484]), .Z(n10773) );
  XNOR U13028 ( .A(n10774), .B(n10773), .Z(n10799) );
  AND U13029 ( .A(n10775), .B(o[99]), .Z(n10800) );
  XOR U13030 ( .A(n10799), .B(n10800), .Z(n10804) );
  AND U13031 ( .A(x[482]), .B(y[7778]), .Z(n10937) );
  NAND U13032 ( .A(y[7779]), .B(x[481]), .Z(n10776) );
  XNOR U13033 ( .A(n10937), .B(n10776), .Z(n10796) );
  AND U13034 ( .A(x[483]), .B(y[7777]), .Z(n10791) );
  XOR U13035 ( .A(o[100]), .B(n10791), .Z(n10795) );
  XOR U13036 ( .A(n10796), .B(n10795), .Z(n10803) );
  XOR U13037 ( .A(n10804), .B(n10803), .Z(n10805) );
  XOR U13038 ( .A(n10806), .B(n10805), .Z(n10810) );
  NANDN U13039 ( .A(n10778), .B(n10777), .Z(n10782) );
  NAND U13040 ( .A(n10780), .B(n10779), .Z(n10781) );
  NAND U13041 ( .A(n10782), .B(n10781), .Z(n10811) );
  NAND U13042 ( .A(n10893), .B(n10783), .Z(n10787) );
  NAND U13043 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U13044 ( .A(n10787), .B(n10786), .Z(n10812) );
  IV U13045 ( .A(n10812), .Z(n10809) );
  XOR U13046 ( .A(n10811), .B(n10809), .Z(n10788) );
  XNOR U13047 ( .A(n10810), .B(n10788), .Z(N229) );
  AND U13048 ( .A(y[7778]), .B(x[483]), .Z(n10790) );
  NAND U13049 ( .A(y[7780]), .B(x[481]), .Z(n10789) );
  XNOR U13050 ( .A(n10790), .B(n10789), .Z(n10815) );
  AND U13051 ( .A(x[484]), .B(y[7777]), .Z(n10824) );
  XOR U13052 ( .A(n10824), .B(o[101]), .Z(n10814) );
  XNOR U13053 ( .A(n10815), .B(n10814), .Z(n10818) );
  NAND U13054 ( .A(x[482]), .B(y[7779]), .Z(n10901) );
  AND U13055 ( .A(o[100]), .B(n10791), .Z(n10820) );
  AND U13056 ( .A(y[7776]), .B(x[485]), .Z(n10793) );
  NAND U13057 ( .A(y[7781]), .B(x[480]), .Z(n10792) );
  XNOR U13058 ( .A(n10793), .B(n10792), .Z(n10821) );
  XOR U13059 ( .A(n10820), .B(n10821), .Z(n10819) );
  XOR U13060 ( .A(n10901), .B(n10819), .Z(n10794) );
  XOR U13061 ( .A(n10818), .B(n10794), .Z(n10836) );
  NANDN U13062 ( .A(n10901), .B(n10893), .Z(n10798) );
  NAND U13063 ( .A(n10796), .B(n10795), .Z(n10797) );
  NAND U13064 ( .A(n10798), .B(n10797), .Z(n10834) );
  AND U13065 ( .A(x[484]), .B(y[7780]), .Z(n11590) );
  NAND U13066 ( .A(n11590), .B(n11395), .Z(n10802) );
  NAND U13067 ( .A(n10800), .B(n10799), .Z(n10801) );
  NAND U13068 ( .A(n10802), .B(n10801), .Z(n10833) );
  XOR U13069 ( .A(n10834), .B(n10833), .Z(n10835) );
  XNOR U13070 ( .A(n10836), .B(n10835), .Z(n10832) );
  NAND U13071 ( .A(n10804), .B(n10803), .Z(n10808) );
  NAND U13072 ( .A(n10806), .B(n10805), .Z(n10807) );
  NAND U13073 ( .A(n10808), .B(n10807), .Z(n10831) );
  XOR U13074 ( .A(n10831), .B(n10830), .Z(n10813) );
  XNOR U13075 ( .A(n10832), .B(n10813), .Z(N230) );
  AND U13076 ( .A(x[483]), .B(y[7780]), .Z(n10902) );
  NAND U13077 ( .A(n10902), .B(n10893), .Z(n10817) );
  NAND U13078 ( .A(n10815), .B(n10814), .Z(n10816) );
  NAND U13079 ( .A(n10817), .B(n10816), .Z(n10871) );
  XOR U13080 ( .A(n10871), .B(n10872), .Z(n10874) );
  AND U13081 ( .A(x[485]), .B(y[7781]), .Z(n11061) );
  NAND U13082 ( .A(n11395), .B(n11061), .Z(n10823) );
  NAND U13083 ( .A(n10821), .B(n10820), .Z(n10822) );
  NAND U13084 ( .A(n10823), .B(n10822), .Z(n10841) );
  AND U13085 ( .A(n10824), .B(o[101]), .Z(n10847) );
  AND U13086 ( .A(y[7776]), .B(x[486]), .Z(n10826) );
  NAND U13087 ( .A(y[7782]), .B(x[480]), .Z(n10825) );
  XNOR U13088 ( .A(n10826), .B(n10825), .Z(n10848) );
  XOR U13089 ( .A(n10847), .B(n10848), .Z(n10840) );
  XOR U13090 ( .A(n10841), .B(n10840), .Z(n10843) );
  NAND U13091 ( .A(y[7780]), .B(x[482]), .Z(n10827) );
  XNOR U13092 ( .A(n10828), .B(n10827), .Z(n10852) );
  AND U13093 ( .A(y[7781]), .B(x[481]), .Z(n11095) );
  NAND U13094 ( .A(y[7778]), .B(x[484]), .Z(n10829) );
  XNOR U13095 ( .A(n11095), .B(n10829), .Z(n10856) );
  NAND U13096 ( .A(x[485]), .B(y[7777]), .Z(n10863) );
  XOR U13097 ( .A(n10856), .B(n10855), .Z(n10851) );
  XOR U13098 ( .A(n10852), .B(n10851), .Z(n10842) );
  XOR U13099 ( .A(n10843), .B(n10842), .Z(n10873) );
  XOR U13100 ( .A(n10874), .B(n10873), .Z(n10867) );
  NAND U13101 ( .A(n10834), .B(n10833), .Z(n10838) );
  NAND U13102 ( .A(n10836), .B(n10835), .Z(n10837) );
  AND U13103 ( .A(n10838), .B(n10837), .Z(n10866) );
  IV U13104 ( .A(n10866), .Z(n10864) );
  XOR U13105 ( .A(n10865), .B(n10864), .Z(n10839) );
  XNOR U13106 ( .A(n10867), .B(n10839), .Z(N231) );
  NAND U13107 ( .A(n10841), .B(n10840), .Z(n10845) );
  NAND U13108 ( .A(n10843), .B(n10842), .Z(n10844) );
  AND U13109 ( .A(n10845), .B(n10844), .Z(n10881) );
  AND U13110 ( .A(y[7778]), .B(x[485]), .Z(n10982) );
  NAND U13111 ( .A(y[7782]), .B(x[481]), .Z(n10846) );
  XNOR U13112 ( .A(n10982), .B(n10846), .Z(n10895) );
  AND U13113 ( .A(x[486]), .B(y[7777]), .Z(n10898) );
  XOR U13114 ( .A(o[103]), .B(n10898), .Z(n10894) );
  XOR U13115 ( .A(n10895), .B(n10894), .Z(n10913) );
  AND U13116 ( .A(x[486]), .B(y[7782]), .Z(n11116) );
  NAND U13117 ( .A(n11395), .B(n11116), .Z(n10850) );
  NAND U13118 ( .A(n10848), .B(n10847), .Z(n10849) );
  AND U13119 ( .A(n10850), .B(n10849), .Z(n10912) );
  NANDN U13120 ( .A(n10901), .B(n10902), .Z(n10854) );
  NAND U13121 ( .A(n10852), .B(n10851), .Z(n10853) );
  AND U13122 ( .A(n10854), .B(n10853), .Z(n10914) );
  XOR U13123 ( .A(n10915), .B(n10914), .Z(n10879) );
  AND U13124 ( .A(x[484]), .B(y[7781]), .Z(n11400) );
  NAND U13125 ( .A(n11400), .B(n10893), .Z(n10858) );
  NAND U13126 ( .A(n10856), .B(n10855), .Z(n10857) );
  AND U13127 ( .A(n10858), .B(n10857), .Z(n10890) );
  AND U13128 ( .A(y[7781]), .B(x[482]), .Z(n10860) );
  NAND U13129 ( .A(y[7779]), .B(x[484]), .Z(n10859) );
  XNOR U13130 ( .A(n10860), .B(n10859), .Z(n10903) );
  XOR U13131 ( .A(n10903), .B(n10902), .Z(n10888) );
  AND U13132 ( .A(y[7776]), .B(x[487]), .Z(n10862) );
  NAND U13133 ( .A(y[7783]), .B(x[480]), .Z(n10861) );
  XNOR U13134 ( .A(n10862), .B(n10861), .Z(n10907) );
  ANDN U13135 ( .B(o[102]), .A(n10863), .Z(n10906) );
  XNOR U13136 ( .A(n10907), .B(n10906), .Z(n10887) );
  XOR U13137 ( .A(n10890), .B(n10889), .Z(n10878) );
  XOR U13138 ( .A(n10879), .B(n10878), .Z(n10880) );
  XNOR U13139 ( .A(n10881), .B(n10880), .Z(n10886) );
  NANDN U13140 ( .A(n10864), .B(n10865), .Z(n10870) );
  NOR U13141 ( .A(n10866), .B(n10865), .Z(n10868) );
  OR U13142 ( .A(n10868), .B(n10867), .Z(n10869) );
  AND U13143 ( .A(n10870), .B(n10869), .Z(n10885) );
  NAND U13144 ( .A(n10872), .B(n10871), .Z(n10876) );
  NAND U13145 ( .A(n10874), .B(n10873), .Z(n10875) );
  AND U13146 ( .A(n10876), .B(n10875), .Z(n10884) );
  XOR U13147 ( .A(n10885), .B(n10884), .Z(n10877) );
  XNOR U13148 ( .A(n10886), .B(n10877), .Z(N232) );
  NAND U13149 ( .A(n10879), .B(n10878), .Z(n10883) );
  NAND U13150 ( .A(n10881), .B(n10880), .Z(n10882) );
  AND U13151 ( .A(n10883), .B(n10882), .Z(n10954) );
  NANDN U13152 ( .A(n10888), .B(n10887), .Z(n10892) );
  NAND U13153 ( .A(n10890), .B(n10889), .Z(n10891) );
  AND U13154 ( .A(n10892), .B(n10891), .Z(n10950) );
  AND U13155 ( .A(x[485]), .B(y[7782]), .Z(n11053) );
  NAND U13156 ( .A(n11053), .B(n10893), .Z(n10897) );
  NAND U13157 ( .A(n10895), .B(n10894), .Z(n10896) );
  AND U13158 ( .A(n10897), .B(n10896), .Z(n10948) );
  AND U13159 ( .A(o[103]), .B(n10898), .Z(n10930) );
  AND U13160 ( .A(x[485]), .B(y[7779]), .Z(n11531) );
  NAND U13161 ( .A(y[7783]), .B(x[481]), .Z(n10899) );
  XNOR U13162 ( .A(n11531), .B(n10899), .Z(n10931) );
  XNOR U13163 ( .A(n10930), .B(n10931), .Z(n10935) );
  NAND U13164 ( .A(x[483]), .B(y[7781]), .Z(n11726) );
  AND U13165 ( .A(x[486]), .B(y[7778]), .Z(n10900) );
  AND U13166 ( .A(y[7782]), .B(x[482]), .Z(n11824) );
  XOR U13167 ( .A(n10900), .B(n11824), .Z(n10938) );
  XNOR U13168 ( .A(n11590), .B(n10938), .Z(n10934) );
  XNOR U13169 ( .A(n11726), .B(n10934), .Z(n10936) );
  XOR U13170 ( .A(n10935), .B(n10936), .Z(n10947) );
  XOR U13171 ( .A(n10950), .B(n10949), .Z(n10959) );
  NANDN U13172 ( .A(n10901), .B(n11400), .Z(n10905) );
  NAND U13173 ( .A(n10903), .B(n10902), .Z(n10904) );
  AND U13174 ( .A(n10905), .B(n10904), .Z(n10944) );
  AND U13175 ( .A(x[487]), .B(y[7783]), .Z(n11293) );
  NAND U13176 ( .A(n11395), .B(n11293), .Z(n10909) );
  NAND U13177 ( .A(n10907), .B(n10906), .Z(n10908) );
  AND U13178 ( .A(n10909), .B(n10908), .Z(n10942) );
  AND U13179 ( .A(y[7776]), .B(x[488]), .Z(n10911) );
  NAND U13180 ( .A(y[7784]), .B(x[480]), .Z(n10910) );
  XNOR U13181 ( .A(n10911), .B(n10910), .Z(n10921) );
  AND U13182 ( .A(x[487]), .B(y[7777]), .Z(n10924) );
  XOR U13183 ( .A(o[104]), .B(n10924), .Z(n10920) );
  XOR U13184 ( .A(n10921), .B(n10920), .Z(n10941) );
  NANDN U13185 ( .A(n10913), .B(n10912), .Z(n10917) );
  NAND U13186 ( .A(n10915), .B(n10914), .Z(n10916) );
  NAND U13187 ( .A(n10917), .B(n10916), .Z(n10956) );
  XNOR U13188 ( .A(n10953), .B(n10955), .Z(n10918) );
  XOR U13189 ( .A(n10954), .B(n10918), .Z(N233) );
  AND U13190 ( .A(x[488]), .B(y[7784]), .Z(n10919) );
  NAND U13191 ( .A(n10919), .B(n11395), .Z(n10923) );
  NAND U13192 ( .A(n10921), .B(n10920), .Z(n10922) );
  AND U13193 ( .A(n10923), .B(n10922), .Z(n11011) );
  AND U13194 ( .A(o[104]), .B(n10924), .Z(n10984) );
  AND U13195 ( .A(y[7780]), .B(x[485]), .Z(n10926) );
  NAND U13196 ( .A(y[7778]), .B(x[487]), .Z(n10925) );
  XNOR U13197 ( .A(n10926), .B(n10925), .Z(n10983) );
  XNOR U13198 ( .A(n10984), .B(n10983), .Z(n11009) );
  AND U13199 ( .A(y[7776]), .B(x[489]), .Z(n10928) );
  NAND U13200 ( .A(y[7785]), .B(x[480]), .Z(n10927) );
  XNOR U13201 ( .A(n10928), .B(n10927), .Z(n10991) );
  AND U13202 ( .A(x[488]), .B(y[7777]), .Z(n11000) );
  XOR U13203 ( .A(o[105]), .B(n11000), .Z(n10990) );
  XNOR U13204 ( .A(n10991), .B(n10990), .Z(n11008) );
  XOR U13205 ( .A(n11009), .B(n11008), .Z(n11010) );
  XNOR U13206 ( .A(n11011), .B(n11010), .Z(n11005) );
  AND U13207 ( .A(y[7779]), .B(x[486]), .Z(n11365) );
  NAND U13208 ( .A(y[7784]), .B(x[481]), .Z(n10929) );
  XNOR U13209 ( .A(n11365), .B(n10929), .Z(n10995) );
  XNOR U13210 ( .A(n11400), .B(n10995), .Z(n11015) );
  NAND U13211 ( .A(x[482]), .B(y[7783]), .Z(n11504) );
  NAND U13212 ( .A(x[483]), .B(y[7782]), .Z(n11318) );
  XOR U13213 ( .A(n11504), .B(n11318), .Z(n11014) );
  XNOR U13214 ( .A(n11015), .B(n11014), .Z(n11003) );
  NAND U13215 ( .A(x[485]), .B(y[7783]), .Z(n11183) );
  AND U13216 ( .A(x[481]), .B(y[7779]), .Z(n10994) );
  NANDN U13217 ( .A(n11183), .B(n10994), .Z(n10933) );
  NAND U13218 ( .A(n10931), .B(n10930), .Z(n10932) );
  NAND U13219 ( .A(n10933), .B(n10932), .Z(n11002) );
  XOR U13220 ( .A(n11003), .B(n11002), .Z(n11004) );
  XNOR U13221 ( .A(n11005), .B(n11004), .Z(n10978) );
  NAND U13222 ( .A(n11116), .B(n10937), .Z(n10940) );
  NAND U13223 ( .A(n11590), .B(n10938), .Z(n10939) );
  AND U13224 ( .A(n10940), .B(n10939), .Z(n10977) );
  XNOR U13225 ( .A(n10976), .B(n10977), .Z(n10979) );
  NANDN U13226 ( .A(n10942), .B(n10941), .Z(n10946) );
  NANDN U13227 ( .A(n10944), .B(n10943), .Z(n10945) );
  AND U13228 ( .A(n10946), .B(n10945), .Z(n10964) );
  NANDN U13229 ( .A(n10948), .B(n10947), .Z(n10952) );
  NAND U13230 ( .A(n10950), .B(n10949), .Z(n10951) );
  NAND U13231 ( .A(n10952), .B(n10951), .Z(n10963) );
  XNOR U13232 ( .A(n10965), .B(n10966), .Z(n10972) );
  NANDN U13233 ( .A(n10957), .B(n10956), .Z(n10961) );
  NANDN U13234 ( .A(n10959), .B(n10958), .Z(n10960) );
  AND U13235 ( .A(n10961), .B(n10960), .Z(n10970) );
  IV U13236 ( .A(n10970), .Z(n10969) );
  XOR U13237 ( .A(n10971), .B(n10969), .Z(n10962) );
  XNOR U13238 ( .A(n10972), .B(n10962), .Z(N234) );
  NANDN U13239 ( .A(n10964), .B(n10963), .Z(n10968) );
  NAND U13240 ( .A(n10966), .B(n10965), .Z(n10967) );
  NAND U13241 ( .A(n10968), .B(n10967), .Z(n11072) );
  IV U13242 ( .A(n11072), .Z(n11071) );
  OR U13243 ( .A(n10971), .B(n10969), .Z(n10975) );
  ANDN U13244 ( .B(n10971), .A(n10970), .Z(n10973) );
  OR U13245 ( .A(n10973), .B(n10972), .Z(n10974) );
  AND U13246 ( .A(n10975), .B(n10974), .Z(n11073) );
  NAND U13247 ( .A(n10977), .B(n10976), .Z(n10981) );
  NANDN U13248 ( .A(n10979), .B(n10978), .Z(n10980) );
  NAND U13249 ( .A(n10981), .B(n10980), .Z(n11080) );
  AND U13250 ( .A(x[487]), .B(y[7780]), .Z(n11055) );
  NAND U13251 ( .A(n11055), .B(n10982), .Z(n10986) );
  NAND U13252 ( .A(n10984), .B(n10983), .Z(n10985) );
  AND U13253 ( .A(n10986), .B(n10985), .Z(n11068) );
  AND U13254 ( .A(y[7779]), .B(x[487]), .Z(n10988) );
  NAND U13255 ( .A(y[7782]), .B(x[484]), .Z(n10987) );
  XNOR U13256 ( .A(n10988), .B(n10987), .Z(n11038) );
  NAND U13257 ( .A(x[486]), .B(y[7780]), .Z(n11039) );
  AND U13258 ( .A(x[488]), .B(y[7778]), .Z(n11261) );
  AND U13259 ( .A(x[489]), .B(y[7777]), .Z(n11049) );
  XOR U13260 ( .A(o[106]), .B(n11049), .Z(n11060) );
  XOR U13261 ( .A(n11261), .B(n11060), .Z(n11062) );
  XNOR U13262 ( .A(n11062), .B(n11061), .Z(n11065) );
  XOR U13263 ( .A(n11066), .B(n11065), .Z(n11067) );
  XNOR U13264 ( .A(n11068), .B(n11067), .Z(n11028) );
  AND U13265 ( .A(x[489]), .B(y[7785]), .Z(n10989) );
  NAND U13266 ( .A(n10989), .B(n11395), .Z(n10993) );
  NAND U13267 ( .A(n10991), .B(n10990), .Z(n10992) );
  NAND U13268 ( .A(n10993), .B(n10992), .Z(n11026) );
  AND U13269 ( .A(x[486]), .B(y[7784]), .Z(n11284) );
  NAND U13270 ( .A(n11284), .B(n10994), .Z(n10997) );
  NAND U13271 ( .A(n11400), .B(n10995), .Z(n10996) );
  NAND U13272 ( .A(n10997), .B(n10996), .Z(n11034) );
  AND U13273 ( .A(y[7776]), .B(x[490]), .Z(n10999) );
  NAND U13274 ( .A(y[7786]), .B(x[480]), .Z(n10998) );
  XNOR U13275 ( .A(n10999), .B(n10998), .Z(n11044) );
  AND U13276 ( .A(o[105]), .B(n11000), .Z(n11043) );
  XOR U13277 ( .A(n11044), .B(n11043), .Z(n11032) );
  AND U13278 ( .A(y[7783]), .B(x[483]), .Z(n11966) );
  NAND U13279 ( .A(y[7785]), .B(x[481]), .Z(n11001) );
  XNOR U13280 ( .A(n11966), .B(n11001), .Z(n11056) );
  AND U13281 ( .A(x[482]), .B(y[7784]), .Z(n11057) );
  XOR U13282 ( .A(n11056), .B(n11057), .Z(n11031) );
  XOR U13283 ( .A(n11032), .B(n11031), .Z(n11033) );
  XOR U13284 ( .A(n11034), .B(n11033), .Z(n11025) );
  XOR U13285 ( .A(n11026), .B(n11025), .Z(n11027) );
  XOR U13286 ( .A(n11028), .B(n11027), .Z(n11079) );
  NAND U13287 ( .A(n11003), .B(n11002), .Z(n11007) );
  NAND U13288 ( .A(n11005), .B(n11004), .Z(n11006) );
  AND U13289 ( .A(n11007), .B(n11006), .Z(n11022) );
  NAND U13290 ( .A(n11009), .B(n11008), .Z(n11013) );
  NAND U13291 ( .A(n11011), .B(n11010), .Z(n11012) );
  AND U13292 ( .A(n11013), .B(n11012), .Z(n11019) );
  NAND U13293 ( .A(n11015), .B(n11014), .Z(n11017) );
  IV U13294 ( .A(n11504), .Z(n11637) );
  ANDN U13295 ( .B(n11318), .A(n11637), .Z(n11016) );
  ANDN U13296 ( .B(n11017), .A(n11016), .Z(n11020) );
  XOR U13297 ( .A(n11019), .B(n11020), .Z(n11021) );
  XOR U13298 ( .A(n11022), .B(n11021), .Z(n11078) );
  XOR U13299 ( .A(n11080), .B(n11081), .Z(n11074) );
  XNOR U13300 ( .A(n11073), .B(n11074), .Z(n11018) );
  XOR U13301 ( .A(n11071), .B(n11018), .Z(N235) );
  NAND U13302 ( .A(n11020), .B(n11019), .Z(n11024) );
  NANDN U13303 ( .A(n11022), .B(n11021), .Z(n11023) );
  AND U13304 ( .A(n11024), .B(n11023), .Z(n11151) );
  NAND U13305 ( .A(n11026), .B(n11025), .Z(n11030) );
  NAND U13306 ( .A(n11028), .B(n11027), .Z(n11029) );
  NAND U13307 ( .A(n11030), .B(n11029), .Z(n11149) );
  NAND U13308 ( .A(n11032), .B(n11031), .Z(n11036) );
  NAND U13309 ( .A(n11034), .B(n11033), .Z(n11035) );
  NAND U13310 ( .A(n11036), .B(n11035), .Z(n11138) );
  AND U13311 ( .A(x[487]), .B(y[7782]), .Z(n11178) );
  AND U13312 ( .A(x[484]), .B(y[7779]), .Z(n11037) );
  NAND U13313 ( .A(n11178), .B(n11037), .Z(n11041) );
  NANDN U13314 ( .A(n11039), .B(n11038), .Z(n11040) );
  AND U13315 ( .A(n11041), .B(n11040), .Z(n11136) );
  AND U13316 ( .A(x[490]), .B(y[7786]), .Z(n11042) );
  NAND U13317 ( .A(n11042), .B(n11395), .Z(n11046) );
  NAND U13318 ( .A(n11044), .B(n11043), .Z(n11045) );
  AND U13319 ( .A(n11046), .B(n11045), .Z(n11132) );
  AND U13320 ( .A(y[7776]), .B(x[491]), .Z(n11048) );
  NAND U13321 ( .A(y[7787]), .B(x[480]), .Z(n11047) );
  XNOR U13322 ( .A(n11048), .B(n11047), .Z(n11107) );
  AND U13323 ( .A(o[106]), .B(n11049), .Z(n11106) );
  XOR U13324 ( .A(n11107), .B(n11106), .Z(n11130) );
  AND U13325 ( .A(y[7781]), .B(x[486]), .Z(n11051) );
  NAND U13326 ( .A(y[7786]), .B(x[481]), .Z(n11050) );
  XNOR U13327 ( .A(n11051), .B(n11050), .Z(n11097) );
  AND U13328 ( .A(x[490]), .B(y[7777]), .Z(n11117) );
  XOR U13329 ( .A(o[107]), .B(n11117), .Z(n11096) );
  XOR U13330 ( .A(n11097), .B(n11096), .Z(n11129) );
  XOR U13331 ( .A(n11130), .B(n11129), .Z(n11131) );
  XNOR U13332 ( .A(n11138), .B(n11137), .Z(n11120) );
  AND U13333 ( .A(x[483]), .B(y[7784]), .Z(n12099) );
  NAND U13334 ( .A(y[7785]), .B(x[482]), .Z(n11052) );
  XNOR U13335 ( .A(n11053), .B(n11052), .Z(n11092) );
  AND U13336 ( .A(x[484]), .B(y[7783]), .Z(n11091) );
  XNOR U13337 ( .A(n11092), .B(n11091), .Z(n11124) );
  XNOR U13338 ( .A(n12099), .B(n11124), .Z(n11126) );
  NAND U13339 ( .A(y[7778]), .B(x[489]), .Z(n11054) );
  XNOR U13340 ( .A(n11055), .B(n11054), .Z(n11112) );
  AND U13341 ( .A(x[488]), .B(y[7779]), .Z(n11111) );
  XNOR U13342 ( .A(n11112), .B(n11111), .Z(n11125) );
  XNOR U13343 ( .A(n11126), .B(n11125), .Z(n11088) );
  AND U13344 ( .A(x[483]), .B(y[7785]), .Z(n11105) );
  IV U13345 ( .A(n11105), .Z(n11174) );
  AND U13346 ( .A(x[481]), .B(y[7783]), .Z(n11390) );
  NANDN U13347 ( .A(n11174), .B(n11390), .Z(n11059) );
  NAND U13348 ( .A(n11057), .B(n11056), .Z(n11058) );
  NAND U13349 ( .A(n11059), .B(n11058), .Z(n11086) );
  NAND U13350 ( .A(n11261), .B(n11060), .Z(n11064) );
  NAND U13351 ( .A(n11062), .B(n11061), .Z(n11063) );
  NAND U13352 ( .A(n11064), .B(n11063), .Z(n11085) );
  XOR U13353 ( .A(n11086), .B(n11085), .Z(n11087) );
  XNOR U13354 ( .A(n11088), .B(n11087), .Z(n11119) );
  NAND U13355 ( .A(n11066), .B(n11065), .Z(n11070) );
  NAND U13356 ( .A(n11068), .B(n11067), .Z(n11069) );
  NAND U13357 ( .A(n11070), .B(n11069), .Z(n11118) );
  XNOR U13358 ( .A(n11119), .B(n11118), .Z(n11121) );
  XOR U13359 ( .A(n11120), .B(n11121), .Z(n11148) );
  XOR U13360 ( .A(n11149), .B(n11148), .Z(n11150) );
  XOR U13361 ( .A(n11151), .B(n11150), .Z(n11144) );
  OR U13362 ( .A(n11073), .B(n11071), .Z(n11077) );
  ANDN U13363 ( .B(n11073), .A(n11072), .Z(n11075) );
  OR U13364 ( .A(n11075), .B(n11074), .Z(n11076) );
  AND U13365 ( .A(n11077), .B(n11076), .Z(n11143) );
  NANDN U13366 ( .A(n11079), .B(n11078), .Z(n11083) );
  NAND U13367 ( .A(n11081), .B(n11080), .Z(n11082) );
  AND U13368 ( .A(n11083), .B(n11082), .Z(n11142) );
  IV U13369 ( .A(n11142), .Z(n11141) );
  XOR U13370 ( .A(n11143), .B(n11141), .Z(n11084) );
  XNOR U13371 ( .A(n11144), .B(n11084), .Z(N236) );
  NAND U13372 ( .A(n11086), .B(n11085), .Z(n11090) );
  NAND U13373 ( .A(n11088), .B(n11087), .Z(n11089) );
  AND U13374 ( .A(n11090), .B(n11089), .Z(n11213) );
  AND U13375 ( .A(x[485]), .B(y[7785]), .Z(n11628) );
  NAND U13376 ( .A(n11824), .B(n11628), .Z(n11094) );
  NAND U13377 ( .A(n11092), .B(n11091), .Z(n11093) );
  NAND U13378 ( .A(n11094), .B(n11093), .Z(n11162) );
  AND U13379 ( .A(x[486]), .B(y[7786]), .Z(n11407) );
  NAND U13380 ( .A(n11407), .B(n11095), .Z(n11099) );
  NAND U13381 ( .A(n11097), .B(n11096), .Z(n11098) );
  NAND U13382 ( .A(n11099), .B(n11098), .Z(n11161) );
  XOR U13383 ( .A(n11162), .B(n11161), .Z(n11164) );
  AND U13384 ( .A(x[489]), .B(y[7779]), .Z(n11819) );
  AND U13385 ( .A(x[490]), .B(y[7778]), .Z(n11873) );
  AND U13386 ( .A(y[7784]), .B(x[484]), .Z(n11100) );
  XOR U13387 ( .A(n11873), .B(n11100), .Z(n11203) );
  XOR U13388 ( .A(n11819), .B(n11203), .Z(n11184) );
  NAND U13389 ( .A(x[487]), .B(y[7781]), .Z(n11182) );
  XOR U13390 ( .A(n11183), .B(n11182), .Z(n11185) );
  AND U13391 ( .A(y[7776]), .B(x[492]), .Z(n11102) );
  NAND U13392 ( .A(y[7788]), .B(x[480]), .Z(n11101) );
  XNOR U13393 ( .A(n11102), .B(n11101), .Z(n11199) );
  AND U13394 ( .A(x[491]), .B(y[7777]), .Z(n11179) );
  XOR U13395 ( .A(n11179), .B(o[108]), .Z(n11198) );
  XOR U13396 ( .A(n11199), .B(n11198), .Z(n11168) );
  AND U13397 ( .A(y[7786]), .B(x[482]), .Z(n11104) );
  NAND U13398 ( .A(y[7780]), .B(x[488]), .Z(n11103) );
  XNOR U13399 ( .A(n11104), .B(n11103), .Z(n11173) );
  XOR U13400 ( .A(n11173), .B(n11105), .Z(n11167) );
  XOR U13401 ( .A(n11168), .B(n11167), .Z(n11170) );
  XOR U13402 ( .A(n11169), .B(n11170), .Z(n11163) );
  XOR U13403 ( .A(n11164), .B(n11163), .Z(n11211) );
  AND U13404 ( .A(x[491]), .B(y[7787]), .Z(n12235) );
  NAND U13405 ( .A(n12235), .B(n11395), .Z(n11109) );
  NAND U13406 ( .A(n11107), .B(n11106), .Z(n11108) );
  NAND U13407 ( .A(n11109), .B(n11108), .Z(n11191) );
  AND U13408 ( .A(x[487]), .B(y[7778]), .Z(n11351) );
  AND U13409 ( .A(x[489]), .B(y[7780]), .Z(n11110) );
  NAND U13410 ( .A(n11351), .B(n11110), .Z(n11114) );
  NAND U13411 ( .A(n11112), .B(n11111), .Z(n11113) );
  NAND U13412 ( .A(n11114), .B(n11113), .Z(n11189) );
  NAND U13413 ( .A(y[7787]), .B(x[481]), .Z(n11115) );
  XNOR U13414 ( .A(n11116), .B(n11115), .Z(n11194) );
  XOR U13415 ( .A(n11194), .B(n11195), .Z(n11188) );
  XOR U13416 ( .A(n11189), .B(n11188), .Z(n11190) );
  XOR U13417 ( .A(n11191), .B(n11190), .Z(n11210) );
  XOR U13418 ( .A(n11211), .B(n11210), .Z(n11212) );
  NAND U13419 ( .A(n11119), .B(n11118), .Z(n11123) );
  NANDN U13420 ( .A(n11121), .B(n11120), .Z(n11122) );
  NAND U13421 ( .A(n11123), .B(n11122), .Z(n11223) );
  XOR U13422 ( .A(n11224), .B(n11223), .Z(n11226) );
  NANDN U13423 ( .A(n12099), .B(n11124), .Z(n11128) );
  NAND U13424 ( .A(n11126), .B(n11125), .Z(n11127) );
  AND U13425 ( .A(n11128), .B(n11127), .Z(n11156) );
  NAND U13426 ( .A(n11130), .B(n11129), .Z(n11134) );
  NANDN U13427 ( .A(n11132), .B(n11131), .Z(n11133) );
  AND U13428 ( .A(n11134), .B(n11133), .Z(n11155) );
  NANDN U13429 ( .A(n11136), .B(n11135), .Z(n11140) );
  NAND U13430 ( .A(n11138), .B(n11137), .Z(n11139) );
  NAND U13431 ( .A(n11140), .B(n11139), .Z(n11158) );
  XNOR U13432 ( .A(n11226), .B(n11225), .Z(n11219) );
  OR U13433 ( .A(n11143), .B(n11141), .Z(n11147) );
  ANDN U13434 ( .B(n11143), .A(n11142), .Z(n11145) );
  OR U13435 ( .A(n11145), .B(n11144), .Z(n11146) );
  AND U13436 ( .A(n11147), .B(n11146), .Z(n11217) );
  NAND U13437 ( .A(n11149), .B(n11148), .Z(n11153) );
  NANDN U13438 ( .A(n11151), .B(n11150), .Z(n11152) );
  AND U13439 ( .A(n11153), .B(n11152), .Z(n11218) );
  IV U13440 ( .A(n11218), .Z(n11216) );
  XOR U13441 ( .A(n11217), .B(n11216), .Z(n11154) );
  XNOR U13442 ( .A(n11219), .B(n11154), .Z(N237) );
  NANDN U13443 ( .A(n11156), .B(n11155), .Z(n11160) );
  NANDN U13444 ( .A(n11158), .B(n11157), .Z(n11159) );
  AND U13445 ( .A(n11160), .B(n11159), .Z(n11236) );
  NAND U13446 ( .A(n11162), .B(n11161), .Z(n11166) );
  NAND U13447 ( .A(n11164), .B(n11163), .Z(n11165) );
  NAND U13448 ( .A(n11166), .B(n11165), .Z(n11240) );
  NAND U13449 ( .A(n11168), .B(n11167), .Z(n11172) );
  NAND U13450 ( .A(n11170), .B(n11169), .Z(n11171) );
  NAND U13451 ( .A(n11172), .B(n11171), .Z(n11247) );
  AND U13452 ( .A(y[7786]), .B(x[488]), .Z(n12501) );
  AND U13453 ( .A(x[482]), .B(y[7780]), .Z(n11361) );
  NAND U13454 ( .A(n12501), .B(n11361), .Z(n11176) );
  NANDN U13455 ( .A(n11174), .B(n11173), .Z(n11175) );
  NAND U13456 ( .A(n11176), .B(n11175), .Z(n11275) );
  NAND U13457 ( .A(y[7788]), .B(x[481]), .Z(n11177) );
  XNOR U13458 ( .A(n11178), .B(n11177), .Z(n11266) );
  NAND U13459 ( .A(n11179), .B(o[108]), .Z(n11267) );
  XNOR U13460 ( .A(n11266), .B(n11267), .Z(n11274) );
  AND U13461 ( .A(x[486]), .B(y[7783]), .Z(n12275) );
  AND U13462 ( .A(y[7787]), .B(x[482]), .Z(n11181) );
  NAND U13463 ( .A(y[7780]), .B(x[489]), .Z(n11180) );
  XNOR U13464 ( .A(n11181), .B(n11180), .Z(n11286) );
  XOR U13465 ( .A(n12275), .B(n11286), .Z(n11273) );
  XOR U13466 ( .A(n11274), .B(n11273), .Z(n11276) );
  XOR U13467 ( .A(n11275), .B(n11276), .Z(n11246) );
  NAND U13468 ( .A(n11183), .B(n11182), .Z(n11187) );
  ANDN U13469 ( .B(n11185), .A(n11184), .Z(n11186) );
  ANDN U13470 ( .B(n11187), .A(n11186), .Z(n11245) );
  XOR U13471 ( .A(n11246), .B(n11245), .Z(n11248) );
  XOR U13472 ( .A(n11247), .B(n11248), .Z(n11239) );
  XOR U13473 ( .A(n11240), .B(n11239), .Z(n11242) );
  NAND U13474 ( .A(n11189), .B(n11188), .Z(n11193) );
  NAND U13475 ( .A(n11191), .B(n11190), .Z(n11192) );
  NAND U13476 ( .A(n11193), .B(n11192), .Z(n11253) );
  AND U13477 ( .A(x[486]), .B(y[7787]), .Z(n11510) );
  IV U13478 ( .A(n11510), .Z(n11630) );
  AND U13479 ( .A(x[481]), .B(y[7782]), .Z(n11265) );
  NANDN U13480 ( .A(n11630), .B(n11265), .Z(n11197) );
  NAND U13481 ( .A(n11195), .B(n11194), .Z(n11196) );
  NAND U13482 ( .A(n11197), .B(n11196), .Z(n11259) );
  AND U13483 ( .A(x[492]), .B(y[7788]), .Z(n12507) );
  AND U13484 ( .A(x[490]), .B(y[7779]), .Z(n12111) );
  AND U13485 ( .A(y[7778]), .B(x[491]), .Z(n12072) );
  NAND U13486 ( .A(y[7781]), .B(x[488]), .Z(n11200) );
  XOR U13487 ( .A(n12072), .B(n11200), .Z(n11262) );
  XNOR U13488 ( .A(n12111), .B(n11262), .Z(n11258) );
  XOR U13489 ( .A(n11257), .B(n11258), .Z(n11260) );
  XOR U13490 ( .A(n11259), .B(n11260), .Z(n11251) );
  AND U13491 ( .A(x[490]), .B(y[7784]), .Z(n11202) );
  AND U13492 ( .A(x[484]), .B(y[7778]), .Z(n11201) );
  NAND U13493 ( .A(n11202), .B(n11201), .Z(n11205) );
  NAND U13494 ( .A(n11819), .B(n11203), .Z(n11204) );
  NAND U13495 ( .A(n11205), .B(n11204), .Z(n11296) );
  AND U13496 ( .A(y[7776]), .B(x[493]), .Z(n11207) );
  NAND U13497 ( .A(y[7789]), .B(x[480]), .Z(n11206) );
  XNOR U13498 ( .A(n11207), .B(n11206), .Z(n11282) );
  AND U13499 ( .A(x[492]), .B(y[7777]), .Z(n11291) );
  XOR U13500 ( .A(o[109]), .B(n11291), .Z(n11281) );
  XOR U13501 ( .A(n11282), .B(n11281), .Z(n11295) );
  AND U13502 ( .A(y[7784]), .B(x[485]), .Z(n11209) );
  NAND U13503 ( .A(y[7786]), .B(x[483]), .Z(n11208) );
  XNOR U13504 ( .A(n11209), .B(n11208), .Z(n11277) );
  NAND U13505 ( .A(x[484]), .B(y[7785]), .Z(n11278) );
  XNOR U13506 ( .A(n11277), .B(n11278), .Z(n11294) );
  XOR U13507 ( .A(n11295), .B(n11294), .Z(n11297) );
  XOR U13508 ( .A(n11296), .B(n11297), .Z(n11252) );
  XOR U13509 ( .A(n11251), .B(n11252), .Z(n11254) );
  XOR U13510 ( .A(n11253), .B(n11254), .Z(n11241) );
  XOR U13511 ( .A(n11242), .B(n11241), .Z(n11234) );
  NAND U13512 ( .A(n11211), .B(n11210), .Z(n11215) );
  NANDN U13513 ( .A(n11213), .B(n11212), .Z(n11214) );
  AND U13514 ( .A(n11215), .B(n11214), .Z(n11233) );
  XOR U13515 ( .A(n11236), .B(n11235), .Z(n11232) );
  NANDN U13516 ( .A(n11216), .B(n11217), .Z(n11222) );
  NOR U13517 ( .A(n11218), .B(n11217), .Z(n11220) );
  OR U13518 ( .A(n11220), .B(n11219), .Z(n11221) );
  AND U13519 ( .A(n11222), .B(n11221), .Z(n11231) );
  NAND U13520 ( .A(n11224), .B(n11223), .Z(n11228) );
  NAND U13521 ( .A(n11226), .B(n11225), .Z(n11227) );
  NAND U13522 ( .A(n11228), .B(n11227), .Z(n11230) );
  XOR U13523 ( .A(n11231), .B(n11230), .Z(n11229) );
  XNOR U13524 ( .A(n11232), .B(n11229), .Z(N238) );
  NANDN U13525 ( .A(n11234), .B(n11233), .Z(n11238) );
  NANDN U13526 ( .A(n11236), .B(n11235), .Z(n11237) );
  NAND U13527 ( .A(n11238), .B(n11237), .Z(n11383) );
  NAND U13528 ( .A(n11240), .B(n11239), .Z(n11244) );
  NAND U13529 ( .A(n11242), .B(n11241), .Z(n11243) );
  NAND U13530 ( .A(n11244), .B(n11243), .Z(n11378) );
  NAND U13531 ( .A(n11246), .B(n11245), .Z(n11250) );
  NAND U13532 ( .A(n11248), .B(n11247), .Z(n11249) );
  NAND U13533 ( .A(n11250), .B(n11249), .Z(n11377) );
  XOR U13534 ( .A(n11378), .B(n11377), .Z(n11380) );
  NAND U13535 ( .A(n11252), .B(n11251), .Z(n11256) );
  NAND U13536 ( .A(n11254), .B(n11253), .Z(n11255) );
  NAND U13537 ( .A(n11256), .B(n11255), .Z(n11303) );
  AND U13538 ( .A(y[7781]), .B(x[491]), .Z(n11421) );
  NAND U13539 ( .A(n11421), .B(n11261), .Z(n11264) );
  NANDN U13540 ( .A(n11262), .B(n12111), .Z(n11263) );
  AND U13541 ( .A(n11264), .B(n11263), .Z(n11335) );
  AND U13542 ( .A(x[487]), .B(y[7788]), .Z(n11834) );
  NAND U13543 ( .A(n11834), .B(n11265), .Z(n11269) );
  NANDN U13544 ( .A(n11267), .B(n11266), .Z(n11268) );
  NAND U13545 ( .A(n11269), .B(n11268), .Z(n11334) );
  XNOR U13546 ( .A(n11335), .B(n11334), .Z(n11337) );
  AND U13547 ( .A(x[484]), .B(y[7786]), .Z(n11735) );
  AND U13548 ( .A(y[7787]), .B(x[483]), .Z(n11271) );
  NAND U13549 ( .A(y[7782]), .B(x[488]), .Z(n11270) );
  XOR U13550 ( .A(n11271), .B(n11270), .Z(n11319) );
  XOR U13551 ( .A(n11628), .B(n11319), .Z(n11328) );
  XNOR U13552 ( .A(n11735), .B(n11328), .Z(n11330) );
  AND U13553 ( .A(x[489]), .B(y[7781]), .Z(n11943) );
  AND U13554 ( .A(x[482]), .B(y[7788]), .Z(n11272) );
  AND U13555 ( .A(y[7780]), .B(x[490]), .Z(n11961) );
  XNOR U13556 ( .A(n11272), .B(n11961), .Z(n11362) );
  XNOR U13557 ( .A(n11943), .B(n11362), .Z(n11329) );
  XOR U13558 ( .A(n11330), .B(n11329), .Z(n11336) );
  XOR U13559 ( .A(n11337), .B(n11336), .Z(n11308) );
  XOR U13560 ( .A(n11308), .B(n11307), .Z(n11310) );
  XOR U13561 ( .A(n11309), .B(n11310), .Z(n11302) );
  AND U13562 ( .A(x[485]), .B(y[7786]), .Z(n11408) );
  NAND U13563 ( .A(n12099), .B(n11408), .Z(n11280) );
  NANDN U13564 ( .A(n11278), .B(n11277), .Z(n11279) );
  AND U13565 ( .A(n11280), .B(n11279), .Z(n11341) );
  AND U13566 ( .A(x[493]), .B(y[7789]), .Z(n12847) );
  NAND U13567 ( .A(y[7779]), .B(x[491]), .Z(n11283) );
  XNOR U13568 ( .A(n11284), .B(n11283), .Z(n11366) );
  NAND U13569 ( .A(x[481]), .B(y[7789]), .Z(n11367) );
  XNOR U13570 ( .A(n11339), .B(n11338), .Z(n11340) );
  XOR U13571 ( .A(n11341), .B(n11340), .Z(n11372) );
  AND U13572 ( .A(x[489]), .B(y[7787]), .Z(n11285) );
  NAND U13573 ( .A(n11285), .B(n11361), .Z(n11288) );
  NAND U13574 ( .A(n12275), .B(n11286), .Z(n11287) );
  AND U13575 ( .A(n11288), .B(n11287), .Z(n11348) );
  AND U13576 ( .A(y[7776]), .B(x[494]), .Z(n11290) );
  NAND U13577 ( .A(y[7790]), .B(x[480]), .Z(n11289) );
  XNOR U13578 ( .A(n11290), .B(n11289), .Z(n11314) );
  AND U13579 ( .A(o[109]), .B(n11291), .Z(n11313) );
  XOR U13580 ( .A(n11314), .B(n11313), .Z(n11345) );
  NAND U13581 ( .A(y[7778]), .B(x[492]), .Z(n11292) );
  XNOR U13582 ( .A(n11293), .B(n11292), .Z(n11353) );
  NAND U13583 ( .A(x[493]), .B(y[7777]), .Z(n11360) );
  XOR U13584 ( .A(n11353), .B(n11352), .Z(n11344) );
  XOR U13585 ( .A(n11345), .B(n11344), .Z(n11347) );
  XOR U13586 ( .A(n11348), .B(n11347), .Z(n11371) );
  XOR U13587 ( .A(n11372), .B(n11371), .Z(n11374) );
  NAND U13588 ( .A(n11295), .B(n11294), .Z(n11299) );
  NAND U13589 ( .A(n11297), .B(n11296), .Z(n11298) );
  AND U13590 ( .A(n11299), .B(n11298), .Z(n11373) );
  XNOR U13591 ( .A(n11374), .B(n11373), .Z(n11301) );
  XOR U13592 ( .A(n11302), .B(n11301), .Z(n11304) );
  XOR U13593 ( .A(n11303), .B(n11304), .Z(n11379) );
  XOR U13594 ( .A(n11380), .B(n11379), .Z(n11385) );
  XOR U13595 ( .A(n11383), .B(n11385), .Z(n11300) );
  XOR U13596 ( .A(n11384), .B(n11300), .Z(N239) );
  NAND U13597 ( .A(n11302), .B(n11301), .Z(n11306) );
  NAND U13598 ( .A(n11304), .B(n11303), .Z(n11305) );
  NAND U13599 ( .A(n11306), .B(n11305), .Z(n11471) );
  NANDN U13600 ( .A(n11308), .B(n11307), .Z(n11312) );
  NANDN U13601 ( .A(n11310), .B(n11309), .Z(n11311) );
  NAND U13602 ( .A(n11312), .B(n11311), .Z(n11389) );
  AND U13603 ( .A(x[494]), .B(y[7790]), .Z(n13096) );
  NAND U13604 ( .A(n11395), .B(n13096), .Z(n11316) );
  NAND U13605 ( .A(n11314), .B(n11313), .Z(n11315) );
  AND U13606 ( .A(n11316), .B(n11315), .Z(n11423) );
  AND U13607 ( .A(x[488]), .B(y[7787]), .Z(n11317) );
  NANDN U13608 ( .A(n11318), .B(n11317), .Z(n11321) );
  NANDN U13609 ( .A(n11319), .B(n11628), .Z(n11320) );
  NAND U13610 ( .A(n11321), .B(n11320), .Z(n11422) );
  AND U13611 ( .A(y[7781]), .B(x[490]), .Z(n11323) );
  NAND U13612 ( .A(y[7787]), .B(x[484]), .Z(n11322) );
  XNOR U13613 ( .A(n11323), .B(n11322), .Z(n11403) );
  AND U13614 ( .A(x[487]), .B(y[7784]), .Z(n11402) );
  XOR U13615 ( .A(n11403), .B(n11402), .Z(n11410) );
  NAND U13616 ( .A(x[486]), .B(y[7785]), .Z(n11541) );
  XNOR U13617 ( .A(n11541), .B(n11408), .Z(n11409) );
  AND U13618 ( .A(y[7789]), .B(x[482]), .Z(n11325) );
  NAND U13619 ( .A(y[7782]), .B(x[489]), .Z(n11324) );
  XNOR U13620 ( .A(n11325), .B(n11324), .Z(n11413) );
  NAND U13621 ( .A(x[483]), .B(y[7788]), .Z(n11414) );
  AND U13622 ( .A(y[7790]), .B(x[481]), .Z(n11327) );
  NAND U13623 ( .A(y[7783]), .B(x[488]), .Z(n11326) );
  XNOR U13624 ( .A(n11327), .B(n11326), .Z(n11392) );
  NAND U13625 ( .A(x[494]), .B(y[7777]), .Z(n11419) );
  XOR U13626 ( .A(n11392), .B(n11391), .Z(n11442) );
  XOR U13627 ( .A(n11443), .B(n11442), .Z(n11445) );
  XOR U13628 ( .A(n11444), .B(n11445), .Z(n11424) );
  XOR U13629 ( .A(n11425), .B(n11424), .Z(n11461) );
  NANDN U13630 ( .A(n11328), .B(n11735), .Z(n11333) );
  IV U13631 ( .A(n11329), .Z(n11331) );
  NANDN U13632 ( .A(n11331), .B(n11330), .Z(n11332) );
  AND U13633 ( .A(n11333), .B(n11332), .Z(n11460) );
  NANDN U13634 ( .A(n11339), .B(n11338), .Z(n11343) );
  NANDN U13635 ( .A(n11341), .B(n11340), .Z(n11342) );
  AND U13636 ( .A(n11343), .B(n11342), .Z(n11451) );
  IV U13637 ( .A(n11344), .Z(n11346) );
  NANDN U13638 ( .A(n11346), .B(n11345), .Z(n11350) );
  NANDN U13639 ( .A(n11348), .B(n11347), .Z(n11349) );
  AND U13640 ( .A(n11350), .B(n11349), .Z(n11449) );
  AND U13641 ( .A(x[492]), .B(y[7783]), .Z(n11826) );
  NAND U13642 ( .A(n11826), .B(n11351), .Z(n11355) );
  NAND U13643 ( .A(n11353), .B(n11352), .Z(n11354) );
  AND U13644 ( .A(n11355), .B(n11354), .Z(n11431) );
  AND U13645 ( .A(y[7780]), .B(x[491]), .Z(n11357) );
  NAND U13646 ( .A(y[7778]), .B(x[493]), .Z(n11356) );
  XNOR U13647 ( .A(n11357), .B(n11356), .Z(n11435) );
  AND U13648 ( .A(x[492]), .B(y[7779]), .Z(n11434) );
  XOR U13649 ( .A(n11435), .B(n11434), .Z(n11429) );
  AND U13650 ( .A(y[7776]), .B(x[495]), .Z(n11359) );
  NAND U13651 ( .A(y[7791]), .B(x[480]), .Z(n11358) );
  XNOR U13652 ( .A(n11359), .B(n11358), .Z(n11397) );
  ANDN U13653 ( .B(o[110]), .A(n11360), .Z(n11396) );
  XNOR U13654 ( .A(n11397), .B(n11396), .Z(n11428) );
  XOR U13655 ( .A(n11431), .B(n11430), .Z(n11457) );
  NAND U13656 ( .A(x[490]), .B(y[7788]), .Z(n12277) );
  NANDN U13657 ( .A(n12277), .B(n11361), .Z(n11364) );
  NANDN U13658 ( .A(n11362), .B(n11943), .Z(n11363) );
  AND U13659 ( .A(n11364), .B(n11363), .Z(n11455) );
  AND U13660 ( .A(x[491]), .B(y[7784]), .Z(n11734) );
  NAND U13661 ( .A(n11734), .B(n11365), .Z(n11369) );
  NANDN U13662 ( .A(n11367), .B(n11366), .Z(n11368) );
  NAND U13663 ( .A(n11369), .B(n11368), .Z(n11454) );
  XNOR U13664 ( .A(n11388), .B(n11387), .Z(n11370) );
  XNOR U13665 ( .A(n11389), .B(n11370), .Z(n11470) );
  NAND U13666 ( .A(n11372), .B(n11371), .Z(n11376) );
  NAND U13667 ( .A(n11374), .B(n11373), .Z(n11375) );
  AND U13668 ( .A(n11376), .B(n11375), .Z(n11469) );
  XOR U13669 ( .A(n11470), .B(n11469), .Z(n11472) );
  XNOR U13670 ( .A(n11471), .B(n11472), .Z(n11468) );
  NAND U13671 ( .A(n11378), .B(n11377), .Z(n11382) );
  NAND U13672 ( .A(n11380), .B(n11379), .Z(n11381) );
  NAND U13673 ( .A(n11382), .B(n11381), .Z(n11467) );
  XOR U13674 ( .A(n11467), .B(n11466), .Z(n11386) );
  XNOR U13675 ( .A(n11468), .B(n11386), .Z(N240) );
  AND U13676 ( .A(x[488]), .B(y[7790]), .Z(n11736) );
  NAND U13677 ( .A(n11736), .B(n11390), .Z(n11394) );
  NAND U13678 ( .A(n11392), .B(n11391), .Z(n11393) );
  AND U13679 ( .A(n11394), .B(n11393), .Z(n11489) );
  AND U13680 ( .A(x[495]), .B(y[7791]), .Z(n13449) );
  NAND U13681 ( .A(n13449), .B(n11395), .Z(n11399) );
  NAND U13682 ( .A(n11397), .B(n11396), .Z(n11398) );
  NAND U13683 ( .A(n11399), .B(n11398), .Z(n11488) );
  AND U13684 ( .A(x[490]), .B(y[7787]), .Z(n11401) );
  NAND U13685 ( .A(n11401), .B(n11400), .Z(n11405) );
  NAND U13686 ( .A(n11403), .B(n11402), .Z(n11404) );
  NAND U13687 ( .A(n11405), .B(n11404), .Z(n11527) );
  AND U13688 ( .A(x[480]), .B(y[7792]), .Z(n11550) );
  NAND U13689 ( .A(x[496]), .B(y[7776]), .Z(n11551) );
  NAND U13690 ( .A(x[495]), .B(y[7777]), .Z(n11537) );
  XOR U13691 ( .A(n11553), .B(n11552), .Z(n11526) );
  NAND U13692 ( .A(y[7785]), .B(x[487]), .Z(n11406) );
  XNOR U13693 ( .A(n11407), .B(n11406), .Z(n11543) );
  AND U13694 ( .A(x[490]), .B(y[7782]), .Z(n11542) );
  XOR U13695 ( .A(n11543), .B(n11542), .Z(n11525) );
  XOR U13696 ( .A(n11526), .B(n11525), .Z(n11528) );
  XOR U13697 ( .A(n11527), .B(n11528), .Z(n11490) );
  XOR U13698 ( .A(n11491), .B(n11490), .Z(n11522) );
  NANDN U13699 ( .A(n11408), .B(n11541), .Z(n11412) );
  NANDN U13700 ( .A(n11410), .B(n11409), .Z(n11411) );
  AND U13701 ( .A(n11412), .B(n11411), .Z(n11520) );
  NAND U13702 ( .A(x[489]), .B(y[7789]), .Z(n12258) );
  NANDN U13703 ( .A(n12258), .B(n11824), .Z(n11416) );
  NANDN U13704 ( .A(n11414), .B(n11413), .Z(n11415) );
  AND U13705 ( .A(n11416), .B(n11415), .Z(n11561) );
  AND U13706 ( .A(y[7791]), .B(x[481]), .Z(n11418) );
  NAND U13707 ( .A(y[7784]), .B(x[488]), .Z(n11417) );
  XNOR U13708 ( .A(n11418), .B(n11417), .Z(n11547) );
  ANDN U13709 ( .B(o[111]), .A(n11419), .Z(n11546) );
  XOR U13710 ( .A(n11547), .B(n11546), .Z(n11559) );
  NAND U13711 ( .A(y[7778]), .B(x[494]), .Z(n11420) );
  XNOR U13712 ( .A(n11421), .B(n11420), .Z(n11500) );
  NAND U13713 ( .A(x[484]), .B(y[7788]), .Z(n11501) );
  XOR U13714 ( .A(n11559), .B(n11558), .Z(n11560) );
  XOR U13715 ( .A(n11561), .B(n11560), .Z(n11519) );
  NANDN U13716 ( .A(n11423), .B(n11422), .Z(n11427) );
  NAND U13717 ( .A(n11425), .B(n11424), .Z(n11426) );
  NAND U13718 ( .A(n11427), .B(n11426), .Z(n11483) );
  NANDN U13719 ( .A(n11429), .B(n11428), .Z(n11433) );
  NAND U13720 ( .A(n11431), .B(n11430), .Z(n11432) );
  AND U13721 ( .A(n11433), .B(n11432), .Z(n11516) );
  AND U13722 ( .A(y[7780]), .B(x[493]), .Z(n11512) );
  NAND U13723 ( .A(n12072), .B(n11512), .Z(n11437) );
  NAND U13724 ( .A(n11435), .B(n11434), .Z(n11436) );
  AND U13725 ( .A(n11437), .B(n11436), .Z(n11497) );
  AND U13726 ( .A(y[7790]), .B(x[482]), .Z(n11439) );
  NAND U13727 ( .A(y[7783]), .B(x[489]), .Z(n11438) );
  XNOR U13728 ( .A(n11439), .B(n11438), .Z(n11505) );
  NAND U13729 ( .A(x[483]), .B(y[7789]), .Z(n11506) );
  AND U13730 ( .A(x[492]), .B(y[7780]), .Z(n12246) );
  AND U13731 ( .A(y[7787]), .B(x[485]), .Z(n11441) );
  NAND U13732 ( .A(y[7779]), .B(x[493]), .Z(n11440) );
  XOR U13733 ( .A(n11441), .B(n11440), .Z(n11532) );
  XOR U13734 ( .A(n11495), .B(n11494), .Z(n11496) );
  NAND U13735 ( .A(n11443), .B(n11442), .Z(n11447) );
  NAND U13736 ( .A(n11445), .B(n11444), .Z(n11446) );
  AND U13737 ( .A(n11447), .B(n11446), .Z(n11514) );
  XOR U13738 ( .A(n11513), .B(n11514), .Z(n11515) );
  XNOR U13739 ( .A(n11485), .B(n11484), .Z(n11564) );
  XNOR U13740 ( .A(n11565), .B(n11564), .Z(n11567) );
  NANDN U13741 ( .A(n11449), .B(n11448), .Z(n11453) );
  NANDN U13742 ( .A(n11451), .B(n11450), .Z(n11452) );
  AND U13743 ( .A(n11453), .B(n11452), .Z(n11479) );
  NANDN U13744 ( .A(n11455), .B(n11454), .Z(n11459) );
  NANDN U13745 ( .A(n11457), .B(n11456), .Z(n11458) );
  AND U13746 ( .A(n11459), .B(n11458), .Z(n11477) );
  NANDN U13747 ( .A(n11461), .B(n11460), .Z(n11465) );
  NANDN U13748 ( .A(n11463), .B(n11462), .Z(n11464) );
  AND U13749 ( .A(n11465), .B(n11464), .Z(n11476) );
  XNOR U13750 ( .A(n11567), .B(n11566), .Z(n11572) );
  NAND U13751 ( .A(n11470), .B(n11469), .Z(n11474) );
  NAND U13752 ( .A(n11472), .B(n11471), .Z(n11473) );
  NAND U13753 ( .A(n11474), .B(n11473), .Z(n11570) );
  XNOR U13754 ( .A(n11571), .B(n11570), .Z(n11475) );
  XNOR U13755 ( .A(n11572), .B(n11475), .Z(N241) );
  NANDN U13756 ( .A(n11477), .B(n11476), .Z(n11481) );
  NANDN U13757 ( .A(n11479), .B(n11478), .Z(n11480) );
  AND U13758 ( .A(n11481), .B(n11480), .Z(n11674) );
  NANDN U13759 ( .A(n11483), .B(n11482), .Z(n11487) );
  NAND U13760 ( .A(n11485), .B(n11484), .Z(n11486) );
  AND U13761 ( .A(n11487), .B(n11486), .Z(n11577) );
  NANDN U13762 ( .A(n11489), .B(n11488), .Z(n11493) );
  NAND U13763 ( .A(n11491), .B(n11490), .Z(n11492) );
  AND U13764 ( .A(n11493), .B(n11492), .Z(n11659) );
  NAND U13765 ( .A(n11495), .B(n11494), .Z(n11499) );
  NANDN U13766 ( .A(n11497), .B(n11496), .Z(n11498) );
  AND U13767 ( .A(n11499), .B(n11498), .Z(n11657) );
  AND U13768 ( .A(x[494]), .B(y[7781]), .Z(n11870) );
  NAND U13769 ( .A(n11870), .B(n12072), .Z(n11503) );
  NANDN U13770 ( .A(n11501), .B(n11500), .Z(n11502) );
  AND U13771 ( .A(n11503), .B(n11502), .Z(n11651) );
  AND U13772 ( .A(x[489]), .B(y[7790]), .Z(n12496) );
  NANDN U13773 ( .A(n11504), .B(n12496), .Z(n11508) );
  NANDN U13774 ( .A(n11506), .B(n11505), .Z(n11507) );
  NAND U13775 ( .A(n11508), .B(n11507), .Z(n11650) );
  AND U13776 ( .A(x[485]), .B(y[7788]), .Z(n11696) );
  NAND U13777 ( .A(y[7785]), .B(x[488]), .Z(n11509) );
  XNOR U13778 ( .A(n11696), .B(n11509), .Z(n11629) );
  XOR U13779 ( .A(n11629), .B(n11510), .Z(n11644) );
  NAND U13780 ( .A(x[487]), .B(y[7786]), .Z(n11645) );
  IV U13781 ( .A(n11645), .Z(n11540) );
  XOR U13782 ( .A(n11644), .B(n11540), .Z(n11647) );
  NAND U13783 ( .A(y[7789]), .B(x[484]), .Z(n11511) );
  XNOR U13784 ( .A(n11512), .B(n11511), .Z(n11591) );
  NAND U13785 ( .A(x[491]), .B(y[7782]), .Z(n11592) );
  XOR U13786 ( .A(n11647), .B(n11646), .Z(n11652) );
  XOR U13787 ( .A(n11653), .B(n11652), .Z(n11656) );
  NAND U13788 ( .A(n11514), .B(n11513), .Z(n11518) );
  NANDN U13789 ( .A(n11516), .B(n11515), .Z(n11517) );
  NAND U13790 ( .A(n11518), .B(n11517), .Z(n11574) );
  XOR U13791 ( .A(n11575), .B(n11574), .Z(n11576) );
  NANDN U13792 ( .A(n11520), .B(n11519), .Z(n11524) );
  NANDN U13793 ( .A(n11522), .B(n11521), .Z(n11523) );
  AND U13794 ( .A(n11524), .B(n11523), .Z(n11583) );
  NAND U13795 ( .A(n11526), .B(n11525), .Z(n11530) );
  NAND U13796 ( .A(n11528), .B(n11527), .Z(n11529) );
  AND U13797 ( .A(n11530), .B(n11529), .Z(n11665) );
  AND U13798 ( .A(x[493]), .B(y[7787]), .Z(n12513) );
  NAND U13799 ( .A(n12513), .B(n11531), .Z(n11534) );
  NANDN U13800 ( .A(n11532), .B(n12246), .Z(n11533) );
  AND U13801 ( .A(n11534), .B(n11533), .Z(n11613) );
  AND U13802 ( .A(y[7792]), .B(x[481]), .Z(n11536) );
  NAND U13803 ( .A(y[7784]), .B(x[489]), .Z(n11535) );
  XNOR U13804 ( .A(n11536), .B(n11535), .Z(n11634) );
  ANDN U13805 ( .B(o[112]), .A(n11537), .Z(n11633) );
  XOR U13806 ( .A(n11634), .B(n11633), .Z(n11611) );
  AND U13807 ( .A(y[7778]), .B(x[495]), .Z(n11539) );
  NAND U13808 ( .A(y[7781]), .B(x[492]), .Z(n11538) );
  XNOR U13809 ( .A(n11539), .B(n11538), .Z(n11587) );
  AND U13810 ( .A(x[494]), .B(y[7779]), .Z(n11586) );
  XOR U13811 ( .A(n11587), .B(n11586), .Z(n11610) );
  XOR U13812 ( .A(n11611), .B(n11610), .Z(n11612) );
  NANDN U13813 ( .A(n11541), .B(n11540), .Z(n11545) );
  NAND U13814 ( .A(n11543), .B(n11542), .Z(n11544) );
  AND U13815 ( .A(n11545), .B(n11544), .Z(n11623) );
  NAND U13816 ( .A(x[488]), .B(y[7791]), .Z(n12400) );
  AND U13817 ( .A(x[481]), .B(y[7784]), .Z(n11714) );
  NANDN U13818 ( .A(n12400), .B(n11714), .Z(n11549) );
  NAND U13819 ( .A(n11547), .B(n11546), .Z(n11548) );
  NAND U13820 ( .A(n11549), .B(n11548), .Z(n11622) );
  NANDN U13821 ( .A(n11551), .B(n11550), .Z(n11555) );
  NAND U13822 ( .A(n11553), .B(n11552), .Z(n11554) );
  AND U13823 ( .A(n11555), .B(n11554), .Z(n11619) );
  AND U13824 ( .A(x[480]), .B(y[7793]), .Z(n11601) );
  AND U13825 ( .A(x[497]), .B(y[7776]), .Z(n11600) );
  XOR U13826 ( .A(n11601), .B(n11600), .Z(n11603) );
  AND U13827 ( .A(x[496]), .B(y[7777]), .Z(n11597) );
  XOR U13828 ( .A(n11597), .B(o[113]), .Z(n11602) );
  XOR U13829 ( .A(n11603), .B(n11602), .Z(n11617) );
  AND U13830 ( .A(y[7791]), .B(x[482]), .Z(n11557) );
  NAND U13831 ( .A(y[7783]), .B(x[490]), .Z(n11556) );
  XNOR U13832 ( .A(n11557), .B(n11556), .Z(n11638) );
  NAND U13833 ( .A(x[483]), .B(y[7790]), .Z(n11639) );
  XOR U13834 ( .A(n11617), .B(n11616), .Z(n11618) );
  XOR U13835 ( .A(n11625), .B(n11624), .Z(n11662) );
  XOR U13836 ( .A(n11663), .B(n11662), .Z(n11664) );
  NAND U13837 ( .A(n11559), .B(n11558), .Z(n11563) );
  NANDN U13838 ( .A(n11561), .B(n11560), .Z(n11562) );
  AND U13839 ( .A(n11563), .B(n11562), .Z(n11581) );
  XOR U13840 ( .A(n11580), .B(n11581), .Z(n11582) );
  XOR U13841 ( .A(n11583), .B(n11582), .Z(n11671) );
  XOR U13842 ( .A(n11672), .B(n11671), .Z(n11673) );
  XOR U13843 ( .A(n11674), .B(n11673), .Z(n11669) );
  NANDN U13844 ( .A(n11565), .B(n11564), .Z(n11569) );
  NAND U13845 ( .A(n11567), .B(n11566), .Z(n11568) );
  AND U13846 ( .A(n11569), .B(n11568), .Z(n11670) );
  XOR U13847 ( .A(n11670), .B(n11668), .Z(n11573) );
  XNOR U13848 ( .A(n11669), .B(n11573), .Z(N242) );
  NAND U13849 ( .A(n11575), .B(n11574), .Z(n11579) );
  NANDN U13850 ( .A(n11577), .B(n11576), .Z(n11578) );
  AND U13851 ( .A(n11579), .B(n11578), .Z(n11790) );
  NAND U13852 ( .A(n11581), .B(n11580), .Z(n11585) );
  NANDN U13853 ( .A(n11583), .B(n11582), .Z(n11584) );
  AND U13854 ( .A(n11585), .B(n11584), .Z(n11788) );
  AND U13855 ( .A(x[492]), .B(y[7778]), .Z(n11933) );
  AND U13856 ( .A(x[495]), .B(y[7781]), .Z(n11832) );
  NAND U13857 ( .A(n11933), .B(n11832), .Z(n11589) );
  NAND U13858 ( .A(n11587), .B(n11586), .Z(n11588) );
  NAND U13859 ( .A(n11589), .B(n11588), .Z(n11762) );
  NAND U13860 ( .A(n12847), .B(n11590), .Z(n11594) );
  NANDN U13861 ( .A(n11592), .B(n11591), .Z(n11593) );
  AND U13862 ( .A(n11594), .B(n11593), .Z(n11753) );
  AND U13863 ( .A(y[7793]), .B(x[481]), .Z(n11596) );
  NAND U13864 ( .A(y[7784]), .B(x[490]), .Z(n11595) );
  XNOR U13865 ( .A(n11596), .B(n11595), .Z(n11715) );
  NAND U13866 ( .A(n11597), .B(o[113]), .Z(n11716) );
  AND U13867 ( .A(y[7779]), .B(x[495]), .Z(n11599) );
  NAND U13868 ( .A(y[7785]), .B(x[489]), .Z(n11598) );
  XNOR U13869 ( .A(n11599), .B(n11598), .Z(n11706) );
  NAND U13870 ( .A(x[494]), .B(y[7780]), .Z(n11707) );
  XOR U13871 ( .A(n11751), .B(n11750), .Z(n11752) );
  XOR U13872 ( .A(n11762), .B(n11763), .Z(n11765) );
  NAND U13873 ( .A(n11601), .B(n11600), .Z(n11605) );
  NAND U13874 ( .A(n11603), .B(n11602), .Z(n11604) );
  NAND U13875 ( .A(n11605), .B(n11604), .Z(n11774) );
  AND U13876 ( .A(y[7778]), .B(x[496]), .Z(n11607) );
  NAND U13877 ( .A(y[7783]), .B(x[491]), .Z(n11606) );
  XNOR U13878 ( .A(n11607), .B(n11606), .Z(n11702) );
  NAND U13879 ( .A(x[482]), .B(y[7792]), .Z(n11703) );
  XOR U13880 ( .A(n11774), .B(n11775), .Z(n11777) );
  AND U13881 ( .A(y[7789]), .B(x[485]), .Z(n11852) );
  NAND U13882 ( .A(y[7788]), .B(x[486]), .Z(n11608) );
  XNOR U13883 ( .A(n11852), .B(n11608), .Z(n11699) );
  NAND U13884 ( .A(y[7790]), .B(x[484]), .Z(n11609) );
  XNOR U13885 ( .A(n12501), .B(n11609), .Z(n11737) );
  NAND U13886 ( .A(x[487]), .B(y[7787]), .Z(n11738) );
  XOR U13887 ( .A(n11699), .B(n11698), .Z(n11776) );
  XOR U13888 ( .A(n11777), .B(n11776), .Z(n11764) );
  XOR U13889 ( .A(n11765), .B(n11764), .Z(n11685) );
  NAND U13890 ( .A(n11611), .B(n11610), .Z(n11615) );
  NANDN U13891 ( .A(n11613), .B(n11612), .Z(n11614) );
  AND U13892 ( .A(n11615), .B(n11614), .Z(n11757) );
  NAND U13893 ( .A(n11617), .B(n11616), .Z(n11621) );
  NANDN U13894 ( .A(n11619), .B(n11618), .Z(n11620) );
  AND U13895 ( .A(n11621), .B(n11620), .Z(n11756) );
  XOR U13896 ( .A(n11757), .B(n11756), .Z(n11759) );
  NANDN U13897 ( .A(n11623), .B(n11622), .Z(n11627) );
  NAND U13898 ( .A(n11625), .B(n11624), .Z(n11626) );
  AND U13899 ( .A(n11627), .B(n11626), .Z(n11758) );
  XOR U13900 ( .A(n11759), .B(n11758), .Z(n11684) );
  AND U13901 ( .A(x[488]), .B(y[7788]), .Z(n11967) );
  NAND U13902 ( .A(n11967), .B(n11628), .Z(n11632) );
  NANDN U13903 ( .A(n11630), .B(n11629), .Z(n11631) );
  NAND U13904 ( .A(n11632), .B(n11631), .Z(n11769) );
  NAND U13905 ( .A(x[489]), .B(y[7792]), .Z(n12617) );
  NANDN U13906 ( .A(n12617), .B(n11714), .Z(n11636) );
  NAND U13907 ( .A(n11634), .B(n11633), .Z(n11635) );
  NAND U13908 ( .A(n11636), .B(n11635), .Z(n11768) );
  XOR U13909 ( .A(n11769), .B(n11768), .Z(n11771) );
  NAND U13910 ( .A(x[490]), .B(y[7791]), .Z(n12618) );
  NANDN U13911 ( .A(n12618), .B(n11637), .Z(n11641) );
  NANDN U13912 ( .A(n11639), .B(n11638), .Z(n11640) );
  AND U13913 ( .A(n11641), .B(n11640), .Z(n11747) );
  AND U13914 ( .A(y[7781]), .B(x[493]), .Z(n11643) );
  NAND U13915 ( .A(y[7791]), .B(x[483]), .Z(n11642) );
  XNOR U13916 ( .A(n11643), .B(n11642), .Z(n11727) );
  NAND U13917 ( .A(x[492]), .B(y[7782]), .Z(n11728) );
  AND U13918 ( .A(x[480]), .B(y[7794]), .Z(n11719) );
  NAND U13919 ( .A(x[498]), .B(y[7776]), .Z(n11720) );
  AND U13920 ( .A(x[497]), .B(y[7777]), .Z(n11741) );
  XOR U13921 ( .A(o[114]), .B(n11741), .Z(n11721) );
  XOR U13922 ( .A(n11722), .B(n11721), .Z(n11744) );
  XOR U13923 ( .A(n11745), .B(n11744), .Z(n11746) );
  XOR U13924 ( .A(n11771), .B(n11770), .Z(n11691) );
  NANDN U13925 ( .A(n11645), .B(n11644), .Z(n11649) );
  NAND U13926 ( .A(n11647), .B(n11646), .Z(n11648) );
  AND U13927 ( .A(n11649), .B(n11648), .Z(n11690) );
  NANDN U13928 ( .A(n11651), .B(n11650), .Z(n11655) );
  NAND U13929 ( .A(n11653), .B(n11652), .Z(n11654) );
  NAND U13930 ( .A(n11655), .B(n11654), .Z(n11693) );
  XOR U13931 ( .A(n11687), .B(n11686), .Z(n11681) );
  NANDN U13932 ( .A(n11657), .B(n11656), .Z(n11661) );
  NANDN U13933 ( .A(n11659), .B(n11658), .Z(n11660) );
  AND U13934 ( .A(n11661), .B(n11660), .Z(n11679) );
  NAND U13935 ( .A(n11663), .B(n11662), .Z(n11667) );
  NANDN U13936 ( .A(n11665), .B(n11664), .Z(n11666) );
  NAND U13937 ( .A(n11667), .B(n11666), .Z(n11678) );
  XOR U13938 ( .A(n11788), .B(n11787), .Z(n11789) );
  XNOR U13939 ( .A(n11790), .B(n11789), .Z(n11783) );
  NAND U13940 ( .A(n11672), .B(n11671), .Z(n11676) );
  NANDN U13941 ( .A(n11674), .B(n11673), .Z(n11675) );
  NAND U13942 ( .A(n11676), .B(n11675), .Z(n11781) );
  IV U13943 ( .A(n11781), .Z(n11780) );
  XOR U13944 ( .A(n11782), .B(n11780), .Z(n11677) );
  XNOR U13945 ( .A(n11783), .B(n11677), .Z(N243) );
  NANDN U13946 ( .A(n11679), .B(n11678), .Z(n11683) );
  NANDN U13947 ( .A(n11681), .B(n11680), .Z(n11682) );
  AND U13948 ( .A(n11683), .B(n11682), .Z(n11797) );
  NANDN U13949 ( .A(n11685), .B(n11684), .Z(n11689) );
  NAND U13950 ( .A(n11687), .B(n11686), .Z(n11688) );
  AND U13951 ( .A(n11689), .B(n11688), .Z(n11795) );
  NANDN U13952 ( .A(n11691), .B(n11690), .Z(n11695) );
  NANDN U13953 ( .A(n11693), .B(n11692), .Z(n11694) );
  AND U13954 ( .A(n11695), .B(n11694), .Z(n11899) );
  AND U13955 ( .A(x[486]), .B(y[7789]), .Z(n11697) );
  NAND U13956 ( .A(n11697), .B(n11696), .Z(n11701) );
  NAND U13957 ( .A(n11699), .B(n11698), .Z(n11700) );
  AND U13958 ( .A(n11701), .B(n11700), .Z(n11893) );
  AND U13959 ( .A(x[496]), .B(y[7783]), .Z(n12262) );
  NAND U13960 ( .A(n12262), .B(n12072), .Z(n11705) );
  NANDN U13961 ( .A(n11703), .B(n11702), .Z(n11704) );
  AND U13962 ( .A(n11705), .B(n11704), .Z(n11891) );
  AND U13963 ( .A(x[495]), .B(y[7785]), .Z(n12524) );
  NAND U13964 ( .A(n12524), .B(n11819), .Z(n11709) );
  NANDN U13965 ( .A(n11707), .B(n11706), .Z(n11708) );
  AND U13966 ( .A(n11709), .B(n11708), .Z(n11810) );
  AND U13967 ( .A(y[7794]), .B(x[481]), .Z(n11711) );
  NAND U13968 ( .A(y[7787]), .B(x[488]), .Z(n11710) );
  XNOR U13969 ( .A(n11711), .B(n11710), .Z(n11869) );
  XOR U13970 ( .A(n11869), .B(n11870), .Z(n11808) );
  AND U13971 ( .A(y[7782]), .B(x[493]), .Z(n11713) );
  NAND U13972 ( .A(y[7793]), .B(x[482]), .Z(n11712) );
  XNOR U13973 ( .A(n11713), .B(n11712), .Z(n11825) );
  XOR U13974 ( .A(n11825), .B(n11826), .Z(n11807) );
  XOR U13975 ( .A(n11808), .B(n11807), .Z(n11809) );
  NAND U13976 ( .A(x[490]), .B(y[7793]), .Z(n12912) );
  NANDN U13977 ( .A(n12912), .B(n11714), .Z(n11718) );
  NANDN U13978 ( .A(n11716), .B(n11715), .Z(n11717) );
  AND U13979 ( .A(n11718), .B(n11717), .Z(n11849) );
  NANDN U13980 ( .A(n11720), .B(n11719), .Z(n11724) );
  NAND U13981 ( .A(n11722), .B(n11721), .Z(n11723) );
  AND U13982 ( .A(n11724), .B(n11723), .Z(n11847) );
  AND U13983 ( .A(y[7779]), .B(x[496]), .Z(n12472) );
  NAND U13984 ( .A(y[7786]), .B(x[489]), .Z(n11725) );
  XNOR U13985 ( .A(n12472), .B(n11725), .Z(n11820) );
  AND U13986 ( .A(x[495]), .B(y[7780]), .Z(n11821) );
  XOR U13987 ( .A(n11820), .B(n11821), .Z(n11846) );
  AND U13988 ( .A(x[493]), .B(y[7791]), .Z(n13126) );
  NANDN U13989 ( .A(n11726), .B(n13126), .Z(n11730) );
  NANDN U13990 ( .A(n11728), .B(n11727), .Z(n11729) );
  AND U13991 ( .A(n11730), .B(n11729), .Z(n11843) );
  AND U13992 ( .A(y[7785]), .B(x[490]), .Z(n11732) );
  NAND U13993 ( .A(y[7778]), .B(x[497]), .Z(n11731) );
  XNOR U13994 ( .A(n11732), .B(n11731), .Z(n11875) );
  AND U13995 ( .A(x[498]), .B(y[7777]), .Z(n11839) );
  XOR U13996 ( .A(o[115]), .B(n11839), .Z(n11874) );
  XOR U13997 ( .A(n11875), .B(n11874), .Z(n11841) );
  NAND U13998 ( .A(y[7792]), .B(x[483]), .Z(n11733) );
  XNOR U13999 ( .A(n11734), .B(n11733), .Z(n11833) );
  XOR U14000 ( .A(n11833), .B(n11834), .Z(n11840) );
  XOR U14001 ( .A(n11841), .B(n11840), .Z(n11842) );
  NAND U14002 ( .A(n11736), .B(n11735), .Z(n11740) );
  NANDN U14003 ( .A(n11738), .B(n11737), .Z(n11739) );
  AND U14004 ( .A(n11740), .B(n11739), .Z(n11816) );
  AND U14005 ( .A(x[480]), .B(y[7795]), .Z(n11856) );
  AND U14006 ( .A(x[499]), .B(y[7776]), .Z(n11857) );
  XOR U14007 ( .A(n11856), .B(n11857), .Z(n11859) );
  AND U14008 ( .A(o[114]), .B(n11741), .Z(n11858) );
  XOR U14009 ( .A(n11859), .B(n11858), .Z(n11814) );
  AND U14010 ( .A(x[484]), .B(y[7791]), .Z(n11981) );
  AND U14011 ( .A(y[7790]), .B(x[485]), .Z(n11743) );
  NAND U14012 ( .A(y[7789]), .B(x[486]), .Z(n11742) );
  XNOR U14013 ( .A(n11743), .B(n11742), .Z(n11853) );
  XOR U14014 ( .A(n11981), .B(n11853), .Z(n11813) );
  XOR U14015 ( .A(n11814), .B(n11813), .Z(n11815) );
  XOR U14016 ( .A(n11816), .B(n11815), .Z(n11884) );
  XOR U14017 ( .A(n11885), .B(n11884), .Z(n11887) );
  XNOR U14018 ( .A(n11886), .B(n11887), .Z(n11880) );
  NAND U14019 ( .A(n11745), .B(n11744), .Z(n11749) );
  NANDN U14020 ( .A(n11747), .B(n11746), .Z(n11748) );
  AND U14021 ( .A(n11749), .B(n11748), .Z(n11879) );
  NAND U14022 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U14023 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U14024 ( .A(n11755), .B(n11754), .Z(n11878) );
  XNOR U14025 ( .A(n11880), .B(n11881), .Z(n11896) );
  XOR U14026 ( .A(n11897), .B(n11896), .Z(n11898) );
  NAND U14027 ( .A(n11757), .B(n11756), .Z(n11761) );
  NAND U14028 ( .A(n11759), .B(n11758), .Z(n11760) );
  AND U14029 ( .A(n11761), .B(n11760), .Z(n11908) );
  NAND U14030 ( .A(n11763), .B(n11762), .Z(n11767) );
  NAND U14031 ( .A(n11765), .B(n11764), .Z(n11766) );
  NAND U14032 ( .A(n11767), .B(n11766), .Z(n11904) );
  NAND U14033 ( .A(n11769), .B(n11768), .Z(n11773) );
  NAND U14034 ( .A(n11771), .B(n11770), .Z(n11772) );
  NAND U14035 ( .A(n11773), .B(n11772), .Z(n11903) );
  NAND U14036 ( .A(n11775), .B(n11774), .Z(n11779) );
  NAND U14037 ( .A(n11777), .B(n11776), .Z(n11778) );
  NAND U14038 ( .A(n11779), .B(n11778), .Z(n11902) );
  XNOR U14039 ( .A(n11903), .B(n11902), .Z(n11905) );
  XNOR U14040 ( .A(n11908), .B(n11909), .Z(n11910) );
  XOR U14041 ( .A(n11795), .B(n11794), .Z(n11796) );
  XOR U14042 ( .A(n11797), .B(n11796), .Z(n11803) );
  OR U14043 ( .A(n11782), .B(n11780), .Z(n11786) );
  ANDN U14044 ( .B(n11782), .A(n11781), .Z(n11784) );
  OR U14045 ( .A(n11784), .B(n11783), .Z(n11785) );
  AND U14046 ( .A(n11786), .B(n11785), .Z(n11802) );
  NAND U14047 ( .A(n11788), .B(n11787), .Z(n11792) );
  NAND U14048 ( .A(n11790), .B(n11789), .Z(n11791) );
  NAND U14049 ( .A(n11792), .B(n11791), .Z(n11801) );
  IV U14050 ( .A(n11801), .Z(n11800) );
  XOR U14051 ( .A(n11802), .B(n11800), .Z(n11793) );
  XNOR U14052 ( .A(n11803), .B(n11793), .Z(N244) );
  NAND U14053 ( .A(n11795), .B(n11794), .Z(n11799) );
  NANDN U14054 ( .A(n11797), .B(n11796), .Z(n11798) );
  NAND U14055 ( .A(n11799), .B(n11798), .Z(n12029) );
  IV U14056 ( .A(n12029), .Z(n12028) );
  OR U14057 ( .A(n11802), .B(n11800), .Z(n11806) );
  ANDN U14058 ( .B(n11802), .A(n11801), .Z(n11804) );
  OR U14059 ( .A(n11804), .B(n11803), .Z(n11805) );
  AND U14060 ( .A(n11806), .B(n11805), .Z(n12030) );
  NAND U14061 ( .A(n11808), .B(n11807), .Z(n11812) );
  NANDN U14062 ( .A(n11810), .B(n11809), .Z(n11811) );
  AND U14063 ( .A(n11812), .B(n11811), .Z(n11916) );
  NAND U14064 ( .A(n11814), .B(n11813), .Z(n11818) );
  NANDN U14065 ( .A(n11816), .B(n11815), .Z(n11817) );
  NAND U14066 ( .A(n11818), .B(n11817), .Z(n11915) );
  AND U14067 ( .A(x[496]), .B(y[7786]), .Z(n12763) );
  NAND U14068 ( .A(n12763), .B(n11819), .Z(n11823) );
  NAND U14069 ( .A(n11821), .B(n11820), .Z(n11822) );
  NAND U14070 ( .A(n11823), .B(n11822), .Z(n11956) );
  AND U14071 ( .A(x[493]), .B(y[7793]), .Z(n13365) );
  NAND U14072 ( .A(n13365), .B(n11824), .Z(n11828) );
  NAND U14073 ( .A(n11826), .B(n11825), .Z(n11827) );
  NAND U14074 ( .A(n11828), .B(n11827), .Z(n12001) );
  AND U14075 ( .A(y[7780]), .B(x[496]), .Z(n11830) );
  NAND U14076 ( .A(y[7786]), .B(x[490]), .Z(n11829) );
  XNOR U14077 ( .A(n11830), .B(n11829), .Z(n11962) );
  AND U14078 ( .A(x[482]), .B(y[7794]), .Z(n11963) );
  XOR U14079 ( .A(n11962), .B(n11963), .Z(n11999) );
  NAND U14080 ( .A(y[7787]), .B(x[489]), .Z(n11831) );
  XNOR U14081 ( .A(n11832), .B(n11831), .Z(n11944) );
  AND U14082 ( .A(x[494]), .B(y[7782]), .Z(n11945) );
  XOR U14083 ( .A(n11944), .B(n11945), .Z(n11998) );
  XOR U14084 ( .A(n11999), .B(n11998), .Z(n12000) );
  XOR U14085 ( .A(n12001), .B(n12000), .Z(n11955) );
  XOR U14086 ( .A(n11956), .B(n11955), .Z(n11958) );
  NAND U14087 ( .A(x[491]), .B(y[7792]), .Z(n12914) );
  NANDN U14088 ( .A(n12914), .B(n12099), .Z(n11836) );
  NAND U14089 ( .A(n11834), .B(n11833), .Z(n11835) );
  NAND U14090 ( .A(n11836), .B(n11835), .Z(n12007) );
  AND U14091 ( .A(y[7785]), .B(x[491]), .Z(n11838) );
  NAND U14092 ( .A(y[7795]), .B(x[481]), .Z(n11837) );
  XNOR U14093 ( .A(n11838), .B(n11837), .Z(n11940) );
  AND U14094 ( .A(x[499]), .B(y[7777]), .Z(n11948) );
  XOR U14095 ( .A(o[116]), .B(n11948), .Z(n11939) );
  XOR U14096 ( .A(n11940), .B(n11939), .Z(n12005) );
  AND U14097 ( .A(x[480]), .B(y[7796]), .Z(n11986) );
  AND U14098 ( .A(x[500]), .B(y[7776]), .Z(n11987) );
  XOR U14099 ( .A(n11986), .B(n11987), .Z(n11989) );
  AND U14100 ( .A(o[115]), .B(n11839), .Z(n11988) );
  XOR U14101 ( .A(n11989), .B(n11988), .Z(n12004) );
  XOR U14102 ( .A(n12005), .B(n12004), .Z(n12006) );
  XOR U14103 ( .A(n12007), .B(n12006), .Z(n11957) );
  XOR U14104 ( .A(n11958), .B(n11957), .Z(n11917) );
  XOR U14105 ( .A(n11918), .B(n11917), .Z(n12013) );
  NAND U14106 ( .A(n11841), .B(n11840), .Z(n11845) );
  NANDN U14107 ( .A(n11843), .B(n11842), .Z(n11844) );
  AND U14108 ( .A(n11845), .B(n11844), .Z(n12011) );
  NANDN U14109 ( .A(n11847), .B(n11846), .Z(n11851) );
  NANDN U14110 ( .A(n11849), .B(n11848), .Z(n11850) );
  AND U14111 ( .A(n11851), .B(n11850), .Z(n11924) );
  NAND U14112 ( .A(x[486]), .B(y[7790]), .Z(n11950) );
  NANDN U14113 ( .A(n11950), .B(n11852), .Z(n11855) );
  NAND U14114 ( .A(n11853), .B(n11981), .Z(n11854) );
  NAND U14115 ( .A(n11855), .B(n11854), .Z(n11930) );
  NAND U14116 ( .A(n11857), .B(n11856), .Z(n11861) );
  NAND U14117 ( .A(n11859), .B(n11858), .Z(n11860) );
  NAND U14118 ( .A(n11861), .B(n11860), .Z(n11928) );
  AND U14119 ( .A(y[7778]), .B(x[498]), .Z(n11863) );
  NAND U14120 ( .A(y[7784]), .B(x[492]), .Z(n11862) );
  XNOR U14121 ( .A(n11863), .B(n11862), .Z(n11934) );
  AND U14122 ( .A(x[497]), .B(y[7779]), .Z(n11935) );
  XOR U14123 ( .A(n11934), .B(n11935), .Z(n11927) );
  XOR U14124 ( .A(n11928), .B(n11927), .Z(n11929) );
  XNOR U14125 ( .A(n11930), .B(n11929), .Z(n11922) );
  AND U14126 ( .A(y[7783]), .B(x[493]), .Z(n11865) );
  NAND U14127 ( .A(y[7793]), .B(x[483]), .Z(n11864) );
  XNOR U14128 ( .A(n11865), .B(n11864), .Z(n11968) );
  XNOR U14129 ( .A(n11968), .B(n11967), .Z(n11952) );
  AND U14130 ( .A(y[7791]), .B(x[485]), .Z(n11867) );
  NAND U14131 ( .A(y[7792]), .B(x[484]), .Z(n11866) );
  XNOR U14132 ( .A(n11867), .B(n11866), .Z(n11983) );
  AND U14133 ( .A(x[487]), .B(y[7789]), .Z(n11982) );
  XNOR U14134 ( .A(n11983), .B(n11982), .Z(n11949) );
  XOR U14135 ( .A(n11950), .B(n11949), .Z(n11951) );
  XNOR U14136 ( .A(n11952), .B(n11951), .Z(n11994) );
  AND U14137 ( .A(x[488]), .B(y[7794]), .Z(n13076) );
  AND U14138 ( .A(x[481]), .B(y[7787]), .Z(n11868) );
  NAND U14139 ( .A(n13076), .B(n11868), .Z(n11872) );
  NAND U14140 ( .A(n11870), .B(n11869), .Z(n11871) );
  NAND U14141 ( .A(n11872), .B(n11871), .Z(n11993) );
  AND U14142 ( .A(x[497]), .B(y[7785]), .Z(n12770) );
  NAND U14143 ( .A(n12770), .B(n11873), .Z(n11877) );
  NAND U14144 ( .A(n11875), .B(n11874), .Z(n11876) );
  NAND U14145 ( .A(n11877), .B(n11876), .Z(n11992) );
  XOR U14146 ( .A(n11993), .B(n11992), .Z(n11995) );
  XNOR U14147 ( .A(n11994), .B(n11995), .Z(n11921) );
  XOR U14148 ( .A(n11922), .B(n11921), .Z(n11923) );
  XOR U14149 ( .A(n11924), .B(n11923), .Z(n12010) );
  XOR U14150 ( .A(n12011), .B(n12010), .Z(n12012) );
  NANDN U14151 ( .A(n11879), .B(n11878), .Z(n11883) );
  NAND U14152 ( .A(n11881), .B(n11880), .Z(n11882) );
  AND U14153 ( .A(n11883), .B(n11882), .Z(n12025) );
  NAND U14154 ( .A(n11885), .B(n11884), .Z(n11889) );
  NAND U14155 ( .A(n11887), .B(n11886), .Z(n11888) );
  AND U14156 ( .A(n11889), .B(n11888), .Z(n12023) );
  NANDN U14157 ( .A(n11891), .B(n11890), .Z(n11895) );
  NANDN U14158 ( .A(n11893), .B(n11892), .Z(n11894) );
  AND U14159 ( .A(n11895), .B(n11894), .Z(n12022) );
  XNOR U14160 ( .A(n12025), .B(n12024), .Z(n12016) );
  XOR U14161 ( .A(n12017), .B(n12016), .Z(n12018) );
  NAND U14162 ( .A(n11897), .B(n11896), .Z(n11901) );
  NANDN U14163 ( .A(n11899), .B(n11898), .Z(n11900) );
  NAND U14164 ( .A(n11901), .B(n11900), .Z(n12019) );
  NAND U14165 ( .A(n11903), .B(n11902), .Z(n11907) );
  NANDN U14166 ( .A(n11905), .B(n11904), .Z(n11906) );
  AND U14167 ( .A(n11907), .B(n11906), .Z(n12036) );
  NANDN U14168 ( .A(n11909), .B(n11908), .Z(n11913) );
  NANDN U14169 ( .A(n11911), .B(n11910), .Z(n11912) );
  AND U14170 ( .A(n11913), .B(n11912), .Z(n12035) );
  XOR U14171 ( .A(n12036), .B(n12035), .Z(n12037) );
  XNOR U14172 ( .A(n12030), .B(n12031), .Z(n11914) );
  XOR U14173 ( .A(n12028), .B(n11914), .Z(N245) );
  NANDN U14174 ( .A(n11916), .B(n11915), .Z(n11920) );
  NAND U14175 ( .A(n11918), .B(n11917), .Z(n11919) );
  AND U14176 ( .A(n11920), .B(n11919), .Z(n12051) );
  NAND U14177 ( .A(n11922), .B(n11921), .Z(n11926) );
  NAND U14178 ( .A(n11924), .B(n11923), .Z(n11925) );
  AND U14179 ( .A(n11926), .B(n11925), .Z(n12049) );
  NAND U14180 ( .A(n11928), .B(n11927), .Z(n11932) );
  NAND U14181 ( .A(n11930), .B(n11929), .Z(n11931) );
  NAND U14182 ( .A(n11932), .B(n11931), .Z(n12142) );
  AND U14183 ( .A(x[498]), .B(y[7784]), .Z(n12769) );
  NAND U14184 ( .A(n12769), .B(n11933), .Z(n11937) );
  NAND U14185 ( .A(n11935), .B(n11934), .Z(n11936) );
  NAND U14186 ( .A(n11937), .B(n11936), .Z(n12122) );
  AND U14187 ( .A(x[491]), .B(y[7795]), .Z(n13487) );
  AND U14188 ( .A(x[481]), .B(y[7785]), .Z(n11938) );
  NAND U14189 ( .A(n13487), .B(n11938), .Z(n11942) );
  NAND U14190 ( .A(n11940), .B(n11939), .Z(n11941) );
  NAND U14191 ( .A(n11942), .B(n11941), .Z(n12121) );
  XOR U14192 ( .A(n12122), .B(n12121), .Z(n12124) );
  AND U14193 ( .A(x[495]), .B(y[7787]), .Z(n12757) );
  NAND U14194 ( .A(n12757), .B(n11943), .Z(n11947) );
  NAND U14195 ( .A(n11945), .B(n11944), .Z(n11946) );
  NAND U14196 ( .A(n11947), .B(n11946), .Z(n12086) );
  AND U14197 ( .A(o[116]), .B(n11948), .Z(n12108) );
  AND U14198 ( .A(x[480]), .B(y[7797]), .Z(n12105) );
  AND U14199 ( .A(x[501]), .B(y[7776]), .Z(n12106) );
  XOR U14200 ( .A(n12105), .B(n12106), .Z(n12107) );
  XOR U14201 ( .A(n12108), .B(n12107), .Z(n12084) );
  AND U14202 ( .A(x[485]), .B(y[7792]), .Z(n12092) );
  AND U14203 ( .A(x[496]), .B(y[7781]), .Z(n12091) );
  XOR U14204 ( .A(n12092), .B(n12091), .Z(n12090) );
  AND U14205 ( .A(x[495]), .B(y[7782]), .Z(n12089) );
  XOR U14206 ( .A(n12090), .B(n12089), .Z(n12083) );
  XOR U14207 ( .A(n12084), .B(n12083), .Z(n12085) );
  XOR U14208 ( .A(n12086), .B(n12085), .Z(n12123) );
  XOR U14209 ( .A(n12124), .B(n12123), .Z(n12139) );
  NAND U14210 ( .A(n11950), .B(n11949), .Z(n11954) );
  NAND U14211 ( .A(n11952), .B(n11951), .Z(n11953) );
  AND U14212 ( .A(n11954), .B(n11953), .Z(n12140) );
  XOR U14213 ( .A(n12139), .B(n12140), .Z(n12141) );
  XOR U14214 ( .A(n12142), .B(n12141), .Z(n12048) );
  XOR U14215 ( .A(n12049), .B(n12048), .Z(n12050) );
  NAND U14216 ( .A(n11956), .B(n11955), .Z(n11960) );
  NAND U14217 ( .A(n11958), .B(n11957), .Z(n11959) );
  NAND U14218 ( .A(n11960), .B(n11959), .Z(n12148) );
  NAND U14219 ( .A(n12763), .B(n11961), .Z(n11965) );
  NAND U14220 ( .A(n11963), .B(n11962), .Z(n11964) );
  NAND U14221 ( .A(n11965), .B(n11964), .Z(n12055) );
  NAND U14222 ( .A(n11966), .B(n13365), .Z(n11970) );
  NAND U14223 ( .A(n11968), .B(n11967), .Z(n11969) );
  NAND U14224 ( .A(n11970), .B(n11969), .Z(n12136) );
  AND U14225 ( .A(y[7778]), .B(x[499]), .Z(n11972) );
  NAND U14226 ( .A(y[7786]), .B(x[491]), .Z(n11971) );
  XNOR U14227 ( .A(n11972), .B(n11971), .Z(n12074) );
  AND U14228 ( .A(x[500]), .B(y[7777]), .Z(n12104) );
  XOR U14229 ( .A(o[117]), .B(n12104), .Z(n12073) );
  XOR U14230 ( .A(n12074), .B(n12073), .Z(n12134) );
  AND U14231 ( .A(y[7779]), .B(x[498]), .Z(n11974) );
  NAND U14232 ( .A(y[7787]), .B(x[490]), .Z(n11973) );
  XNOR U14233 ( .A(n11974), .B(n11973), .Z(n12112) );
  AND U14234 ( .A(x[481]), .B(y[7796]), .Z(n12113) );
  XOR U14235 ( .A(n12112), .B(n12113), .Z(n12133) );
  XOR U14236 ( .A(n12134), .B(n12133), .Z(n12135) );
  XOR U14237 ( .A(n12136), .B(n12135), .Z(n12054) );
  XOR U14238 ( .A(n12055), .B(n12054), .Z(n12057) );
  AND U14239 ( .A(x[487]), .B(y[7790]), .Z(n12398) );
  AND U14240 ( .A(y[7791]), .B(x[486]), .Z(n11976) );
  NAND U14241 ( .A(y[7783]), .B(x[494]), .Z(n11975) );
  XNOR U14242 ( .A(n11976), .B(n11975), .Z(n12116) );
  XNOR U14243 ( .A(n12398), .B(n12116), .Z(n12063) );
  NAND U14244 ( .A(x[489]), .B(y[7788]), .Z(n12061) );
  NAND U14245 ( .A(x[488]), .B(y[7789]), .Z(n12060) );
  XOR U14246 ( .A(n12061), .B(n12060), .Z(n12062) );
  XNOR U14247 ( .A(n12063), .B(n12062), .Z(n12079) );
  AND U14248 ( .A(y[7785]), .B(x[492]), .Z(n11978) );
  NAND U14249 ( .A(y[7780]), .B(x[497]), .Z(n11977) );
  XNOR U14250 ( .A(n11978), .B(n11977), .Z(n12066) );
  AND U14251 ( .A(x[482]), .B(y[7795]), .Z(n12067) );
  XOR U14252 ( .A(n12066), .B(n12067), .Z(n12078) );
  AND U14253 ( .A(y[7784]), .B(x[493]), .Z(n11980) );
  NAND U14254 ( .A(y[7794]), .B(x[483]), .Z(n11979) );
  XNOR U14255 ( .A(n11980), .B(n11979), .Z(n12100) );
  AND U14256 ( .A(x[484]), .B(y[7793]), .Z(n12101) );
  XOR U14257 ( .A(n12100), .B(n12101), .Z(n12077) );
  XOR U14258 ( .A(n12078), .B(n12077), .Z(n12080) );
  XOR U14259 ( .A(n12079), .B(n12080), .Z(n12130) );
  NAND U14260 ( .A(n12092), .B(n11981), .Z(n11985) );
  NAND U14261 ( .A(n11983), .B(n11982), .Z(n11984) );
  NAND U14262 ( .A(n11985), .B(n11984), .Z(n12128) );
  NAND U14263 ( .A(n11987), .B(n11986), .Z(n11991) );
  NAND U14264 ( .A(n11989), .B(n11988), .Z(n11990) );
  NAND U14265 ( .A(n11991), .B(n11990), .Z(n12127) );
  XOR U14266 ( .A(n12128), .B(n12127), .Z(n12129) );
  XOR U14267 ( .A(n12130), .B(n12129), .Z(n12056) );
  XOR U14268 ( .A(n12057), .B(n12056), .Z(n12146) );
  NAND U14269 ( .A(n11993), .B(n11992), .Z(n11997) );
  NAND U14270 ( .A(n11995), .B(n11994), .Z(n11996) );
  NAND U14271 ( .A(n11997), .B(n11996), .Z(n12153) );
  NAND U14272 ( .A(n11999), .B(n11998), .Z(n12003) );
  NAND U14273 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U14274 ( .A(n12003), .B(n12002), .Z(n12152) );
  NAND U14275 ( .A(n12005), .B(n12004), .Z(n12009) );
  NAND U14276 ( .A(n12007), .B(n12006), .Z(n12008) );
  NAND U14277 ( .A(n12009), .B(n12008), .Z(n12151) );
  XOR U14278 ( .A(n12152), .B(n12151), .Z(n12154) );
  XOR U14279 ( .A(n12153), .B(n12154), .Z(n12145) );
  XOR U14280 ( .A(n12146), .B(n12145), .Z(n12147) );
  XNOR U14281 ( .A(n12148), .B(n12147), .Z(n12043) );
  NAND U14282 ( .A(n12011), .B(n12010), .Z(n12015) );
  NANDN U14283 ( .A(n12013), .B(n12012), .Z(n12014) );
  NAND U14284 ( .A(n12015), .B(n12014), .Z(n12042) );
  XOR U14285 ( .A(n12043), .B(n12042), .Z(n12045) );
  XNOR U14286 ( .A(n12044), .B(n12045), .Z(n12166) );
  NAND U14287 ( .A(n12017), .B(n12016), .Z(n12021) );
  NANDN U14288 ( .A(n12019), .B(n12018), .Z(n12020) );
  AND U14289 ( .A(n12021), .B(n12020), .Z(n12165) );
  NANDN U14290 ( .A(n12023), .B(n12022), .Z(n12027) );
  NAND U14291 ( .A(n12025), .B(n12024), .Z(n12026) );
  AND U14292 ( .A(n12027), .B(n12026), .Z(n12164) );
  XNOR U14293 ( .A(n12166), .B(n12167), .Z(n12160) );
  OR U14294 ( .A(n12030), .B(n12028), .Z(n12034) );
  ANDN U14295 ( .B(n12030), .A(n12029), .Z(n12032) );
  OR U14296 ( .A(n12032), .B(n12031), .Z(n12033) );
  AND U14297 ( .A(n12034), .B(n12033), .Z(n12159) );
  NAND U14298 ( .A(n12036), .B(n12035), .Z(n12040) );
  NANDN U14299 ( .A(n12038), .B(n12037), .Z(n12039) );
  AND U14300 ( .A(n12040), .B(n12039), .Z(n12158) );
  IV U14301 ( .A(n12158), .Z(n12157) );
  XOR U14302 ( .A(n12159), .B(n12157), .Z(n12041) );
  XNOR U14303 ( .A(n12160), .B(n12041), .Z(N246) );
  NAND U14304 ( .A(n12043), .B(n12042), .Z(n12047) );
  NAND U14305 ( .A(n12045), .B(n12044), .Z(n12046) );
  AND U14306 ( .A(n12047), .B(n12046), .Z(n12174) );
  NAND U14307 ( .A(n12049), .B(n12048), .Z(n12053) );
  NANDN U14308 ( .A(n12051), .B(n12050), .Z(n12052) );
  AND U14309 ( .A(n12053), .B(n12052), .Z(n12172) );
  NAND U14310 ( .A(n12055), .B(n12054), .Z(n12059) );
  NAND U14311 ( .A(n12057), .B(n12056), .Z(n12058) );
  AND U14312 ( .A(n12059), .B(n12058), .Z(n12301) );
  NAND U14313 ( .A(n12061), .B(n12060), .Z(n12065) );
  NAND U14314 ( .A(n12063), .B(n12062), .Z(n12064) );
  NAND U14315 ( .A(n12065), .B(n12064), .Z(n12295) );
  NAND U14316 ( .A(n12770), .B(n12246), .Z(n12069) );
  NAND U14317 ( .A(n12067), .B(n12066), .Z(n12068) );
  NAND U14318 ( .A(n12069), .B(n12068), .Z(n12222) );
  AND U14319 ( .A(x[485]), .B(y[7793]), .Z(n12268) );
  AND U14320 ( .A(x[497]), .B(y[7781]), .Z(n12269) );
  XOR U14321 ( .A(n12268), .B(n12269), .Z(n12270) );
  AND U14322 ( .A(x[496]), .B(y[7782]), .Z(n12271) );
  XOR U14323 ( .A(n12270), .B(n12271), .Z(n12221) );
  AND U14324 ( .A(y[7780]), .B(x[498]), .Z(n12071) );
  NAND U14325 ( .A(y[7786]), .B(x[492]), .Z(n12070) );
  XNOR U14326 ( .A(n12071), .B(n12070), .Z(n12247) );
  AND U14327 ( .A(x[484]), .B(y[7794]), .Z(n12248) );
  XOR U14328 ( .A(n12247), .B(n12248), .Z(n12220) );
  XOR U14329 ( .A(n12221), .B(n12220), .Z(n12223) );
  XNOR U14330 ( .A(n12222), .B(n12223), .Z(n12292) );
  AND U14331 ( .A(x[499]), .B(y[7786]), .Z(n13256) );
  NAND U14332 ( .A(n13256), .B(n12072), .Z(n12076) );
  NAND U14333 ( .A(n12074), .B(n12073), .Z(n12075) );
  AND U14334 ( .A(n12076), .B(n12075), .Z(n12293) );
  XOR U14335 ( .A(n12292), .B(n12293), .Z(n12294) );
  XNOR U14336 ( .A(n12295), .B(n12294), .Z(n12298) );
  NAND U14337 ( .A(n12078), .B(n12077), .Z(n12082) );
  NAND U14338 ( .A(n12080), .B(n12079), .Z(n12081) );
  NAND U14339 ( .A(n12082), .B(n12081), .Z(n12281) );
  NAND U14340 ( .A(n12084), .B(n12083), .Z(n12088) );
  NAND U14341 ( .A(n12086), .B(n12085), .Z(n12087) );
  NAND U14342 ( .A(n12088), .B(n12087), .Z(n12280) );
  XOR U14343 ( .A(n12281), .B(n12280), .Z(n12283) );
  AND U14344 ( .A(n12090), .B(n12089), .Z(n12094) );
  NAND U14345 ( .A(n12092), .B(n12091), .Z(n12093) );
  NANDN U14346 ( .A(n12094), .B(n12093), .Z(n12243) );
  AND U14347 ( .A(y[7785]), .B(x[493]), .Z(n12096) );
  NAND U14348 ( .A(y[7778]), .B(x[500]), .Z(n12095) );
  XNOR U14349 ( .A(n12096), .B(n12095), .Z(n12264) );
  AND U14350 ( .A(x[482]), .B(y[7796]), .Z(n12265) );
  XOR U14351 ( .A(n12264), .B(n12265), .Z(n12241) );
  AND U14352 ( .A(y[7792]), .B(x[486]), .Z(n12098) );
  NAND U14353 ( .A(y[7783]), .B(x[495]), .Z(n12097) );
  XNOR U14354 ( .A(n12098), .B(n12097), .Z(n12276) );
  XOR U14355 ( .A(n12241), .B(n12240), .Z(n12242) );
  XOR U14356 ( .A(n12243), .B(n12242), .Z(n12287) );
  AND U14357 ( .A(x[493]), .B(y[7794]), .Z(n13527) );
  NAND U14358 ( .A(n12099), .B(n13527), .Z(n12103) );
  NAND U14359 ( .A(n12101), .B(n12100), .Z(n12102) );
  NAND U14360 ( .A(n12103), .B(n12102), .Z(n12211) );
  AND U14361 ( .A(x[481]), .B(y[7797]), .Z(n12234) );
  XOR U14362 ( .A(n12235), .B(n12234), .Z(n12233) );
  AND U14363 ( .A(o[117]), .B(n12104), .Z(n12232) );
  XOR U14364 ( .A(n12233), .B(n12232), .Z(n12209) );
  AND U14365 ( .A(x[494]), .B(y[7784]), .Z(n12226) );
  AND U14366 ( .A(x[483]), .B(y[7795]), .Z(n12227) );
  XOR U14367 ( .A(n12226), .B(n12227), .Z(n12228) );
  AND U14368 ( .A(x[499]), .B(y[7779]), .Z(n12229) );
  XOR U14369 ( .A(n12228), .B(n12229), .Z(n12208) );
  XOR U14370 ( .A(n12209), .B(n12208), .Z(n12210) );
  XOR U14371 ( .A(n12211), .B(n12210), .Z(n12286) );
  XOR U14372 ( .A(n12287), .B(n12286), .Z(n12289) );
  NAND U14373 ( .A(n12106), .B(n12105), .Z(n12110) );
  NAND U14374 ( .A(n12108), .B(n12107), .Z(n12109) );
  NAND U14375 ( .A(n12110), .B(n12109), .Z(n12203) );
  AND U14376 ( .A(x[498]), .B(y[7787]), .Z(n13258) );
  NAND U14377 ( .A(n13258), .B(n12111), .Z(n12115) );
  NAND U14378 ( .A(n12113), .B(n12112), .Z(n12114) );
  NAND U14379 ( .A(n12115), .B(n12114), .Z(n12202) );
  XOR U14380 ( .A(n12203), .B(n12202), .Z(n12205) );
  AND U14381 ( .A(x[494]), .B(y[7791]), .Z(n13268) );
  NAND U14382 ( .A(n12275), .B(n13268), .Z(n12118) );
  NAND U14383 ( .A(n12398), .B(n12116), .Z(n12117) );
  NAND U14384 ( .A(n12118), .B(n12117), .Z(n12217) );
  AND U14385 ( .A(x[480]), .B(y[7798]), .Z(n12251) );
  AND U14386 ( .A(x[502]), .B(y[7776]), .Z(n12252) );
  XOR U14387 ( .A(n12251), .B(n12252), .Z(n12254) );
  AND U14388 ( .A(x[501]), .B(y[7777]), .Z(n12274) );
  XOR U14389 ( .A(o[118]), .B(n12274), .Z(n12253) );
  XOR U14390 ( .A(n12254), .B(n12253), .Z(n12215) );
  AND U14391 ( .A(y[7791]), .B(x[487]), .Z(n12120) );
  NAND U14392 ( .A(y[7790]), .B(x[488]), .Z(n12119) );
  XNOR U14393 ( .A(n12120), .B(n12119), .Z(n12257) );
  XOR U14394 ( .A(n12215), .B(n12214), .Z(n12216) );
  XOR U14395 ( .A(n12217), .B(n12216), .Z(n12204) );
  XOR U14396 ( .A(n12205), .B(n12204), .Z(n12288) );
  XOR U14397 ( .A(n12289), .B(n12288), .Z(n12282) );
  XOR U14398 ( .A(n12283), .B(n12282), .Z(n12299) );
  XOR U14399 ( .A(n12298), .B(n12299), .Z(n12300) );
  NAND U14400 ( .A(n12122), .B(n12121), .Z(n12126) );
  NAND U14401 ( .A(n12124), .B(n12123), .Z(n12125) );
  NAND U14402 ( .A(n12126), .B(n12125), .Z(n12199) );
  NAND U14403 ( .A(n12128), .B(n12127), .Z(n12132) );
  NAND U14404 ( .A(n12130), .B(n12129), .Z(n12131) );
  NAND U14405 ( .A(n12132), .B(n12131), .Z(n12197) );
  NAND U14406 ( .A(n12134), .B(n12133), .Z(n12138) );
  NAND U14407 ( .A(n12136), .B(n12135), .Z(n12137) );
  NAND U14408 ( .A(n12138), .B(n12137), .Z(n12196) );
  XOR U14409 ( .A(n12197), .B(n12196), .Z(n12198) );
  XNOR U14410 ( .A(n12199), .B(n12198), .Z(n12190) );
  NAND U14411 ( .A(n12140), .B(n12139), .Z(n12144) );
  NAND U14412 ( .A(n12142), .B(n12141), .Z(n12143) );
  AND U14413 ( .A(n12144), .B(n12143), .Z(n12191) );
  XOR U14414 ( .A(n12190), .B(n12191), .Z(n12193) );
  XNOR U14415 ( .A(n12192), .B(n12193), .Z(n12186) );
  NAND U14416 ( .A(n12146), .B(n12145), .Z(n12150) );
  NAND U14417 ( .A(n12148), .B(n12147), .Z(n12149) );
  NAND U14418 ( .A(n12150), .B(n12149), .Z(n12185) );
  NAND U14419 ( .A(n12152), .B(n12151), .Z(n12156) );
  NAND U14420 ( .A(n12154), .B(n12153), .Z(n12155) );
  NAND U14421 ( .A(n12156), .B(n12155), .Z(n12184) );
  XOR U14422 ( .A(n12185), .B(n12184), .Z(n12187) );
  XOR U14423 ( .A(n12186), .B(n12187), .Z(n12171) );
  XNOR U14424 ( .A(n12174), .B(n12173), .Z(n12180) );
  OR U14425 ( .A(n12159), .B(n12157), .Z(n12163) );
  ANDN U14426 ( .B(n12159), .A(n12158), .Z(n12161) );
  OR U14427 ( .A(n12161), .B(n12160), .Z(n12162) );
  AND U14428 ( .A(n12163), .B(n12162), .Z(n12179) );
  NANDN U14429 ( .A(n12165), .B(n12164), .Z(n12169) );
  NAND U14430 ( .A(n12167), .B(n12166), .Z(n12168) );
  NAND U14431 ( .A(n12169), .B(n12168), .Z(n12178) );
  IV U14432 ( .A(n12178), .Z(n12177) );
  XOR U14433 ( .A(n12179), .B(n12177), .Z(n12170) );
  XNOR U14434 ( .A(n12180), .B(n12170), .Z(N247) );
  NANDN U14435 ( .A(n12172), .B(n12171), .Z(n12176) );
  NAND U14436 ( .A(n12174), .B(n12173), .Z(n12175) );
  NAND U14437 ( .A(n12176), .B(n12175), .Z(n12312) );
  IV U14438 ( .A(n12312), .Z(n12311) );
  OR U14439 ( .A(n12179), .B(n12177), .Z(n12183) );
  ANDN U14440 ( .B(n12179), .A(n12178), .Z(n12181) );
  OR U14441 ( .A(n12181), .B(n12180), .Z(n12182) );
  AND U14442 ( .A(n12183), .B(n12182), .Z(n12313) );
  NAND U14443 ( .A(n12185), .B(n12184), .Z(n12189) );
  NAND U14444 ( .A(n12187), .B(n12186), .Z(n12188) );
  AND U14445 ( .A(n12189), .B(n12188), .Z(n12308) );
  NAND U14446 ( .A(n12191), .B(n12190), .Z(n12195) );
  NAND U14447 ( .A(n12193), .B(n12192), .Z(n12194) );
  NAND U14448 ( .A(n12195), .B(n12194), .Z(n12306) );
  NAND U14449 ( .A(n12197), .B(n12196), .Z(n12201) );
  NAND U14450 ( .A(n12199), .B(n12198), .Z(n12200) );
  NAND U14451 ( .A(n12201), .B(n12200), .Z(n12434) );
  NAND U14452 ( .A(n12203), .B(n12202), .Z(n12207) );
  NAND U14453 ( .A(n12205), .B(n12204), .Z(n12206) );
  NAND U14454 ( .A(n12207), .B(n12206), .Z(n12381) );
  NAND U14455 ( .A(n12209), .B(n12208), .Z(n12213) );
  NAND U14456 ( .A(n12211), .B(n12210), .Z(n12212) );
  NAND U14457 ( .A(n12213), .B(n12212), .Z(n12379) );
  NAND U14458 ( .A(n12215), .B(n12214), .Z(n12219) );
  NAND U14459 ( .A(n12217), .B(n12216), .Z(n12218) );
  NAND U14460 ( .A(n12219), .B(n12218), .Z(n12378) );
  XOR U14461 ( .A(n12379), .B(n12378), .Z(n12380) );
  XOR U14462 ( .A(n12381), .B(n12380), .Z(n12446) );
  NAND U14463 ( .A(n12221), .B(n12220), .Z(n12225) );
  NAND U14464 ( .A(n12223), .B(n12222), .Z(n12224) );
  NAND U14465 ( .A(n12225), .B(n12224), .Z(n12444) );
  NAND U14466 ( .A(n12227), .B(n12226), .Z(n12231) );
  NAND U14467 ( .A(n12229), .B(n12228), .Z(n12230) );
  NAND U14468 ( .A(n12231), .B(n12230), .Z(n12325) );
  AND U14469 ( .A(n12233), .B(n12232), .Z(n12237) );
  NAND U14470 ( .A(n12235), .B(n12234), .Z(n12236) );
  NANDN U14471 ( .A(n12237), .B(n12236), .Z(n12324) );
  XOR U14472 ( .A(n12325), .B(n12324), .Z(n12327) );
  AND U14473 ( .A(y[7792]), .B(x[487]), .Z(n12239) );
  NAND U14474 ( .A(y[7790]), .B(x[489]), .Z(n12238) );
  XNOR U14475 ( .A(n12239), .B(n12238), .Z(n12399) );
  AND U14476 ( .A(x[490]), .B(y[7789]), .Z(n12330) );
  XOR U14477 ( .A(n12331), .B(n12330), .Z(n12333) );
  AND U14478 ( .A(x[486]), .B(y[7793]), .Z(n12390) );
  NAND U14479 ( .A(x[495]), .B(y[7784]), .Z(n12391) );
  XNOR U14480 ( .A(n12390), .B(n12391), .Z(n12393) );
  AND U14481 ( .A(x[491]), .B(y[7788]), .Z(n12392) );
  XOR U14482 ( .A(n12393), .B(n12392), .Z(n12332) );
  XOR U14483 ( .A(n12333), .B(n12332), .Z(n12326) );
  XOR U14484 ( .A(n12327), .B(n12326), .Z(n12443) );
  XOR U14485 ( .A(n12444), .B(n12443), .Z(n12445) );
  XOR U14486 ( .A(n12446), .B(n12445), .Z(n12432) );
  NAND U14487 ( .A(n12241), .B(n12240), .Z(n12245) );
  NAND U14488 ( .A(n12243), .B(n12242), .Z(n12244) );
  NAND U14489 ( .A(n12245), .B(n12244), .Z(n12426) );
  AND U14490 ( .A(x[498]), .B(y[7786]), .Z(n13114) );
  NAND U14491 ( .A(n13114), .B(n12246), .Z(n12250) );
  NAND U14492 ( .A(n12248), .B(n12247), .Z(n12249) );
  NAND U14493 ( .A(n12250), .B(n12249), .Z(n12355) );
  NAND U14494 ( .A(n12252), .B(n12251), .Z(n12256) );
  NAND U14495 ( .A(n12254), .B(n12253), .Z(n12255) );
  NAND U14496 ( .A(n12256), .B(n12255), .Z(n12354) );
  XOR U14497 ( .A(n12355), .B(n12354), .Z(n12357) );
  NANDN U14498 ( .A(n12400), .B(n12398), .Z(n12260) );
  NANDN U14499 ( .A(n12258), .B(n12257), .Z(n12259) );
  AND U14500 ( .A(n12260), .B(n12259), .Z(n12369) );
  AND U14501 ( .A(x[480]), .B(y[7799]), .Z(n12410) );
  AND U14502 ( .A(x[503]), .B(y[7776]), .Z(n12409) );
  XOR U14503 ( .A(n12410), .B(n12409), .Z(n12412) );
  AND U14504 ( .A(x[502]), .B(y[7777]), .Z(n12389) );
  XOR U14505 ( .A(n12389), .B(o[119]), .Z(n12411) );
  XOR U14506 ( .A(n12412), .B(n12411), .Z(n12366) );
  NAND U14507 ( .A(y[7779]), .B(x[500]), .Z(n12261) );
  XNOR U14508 ( .A(n12262), .B(n12261), .Z(n12385) );
  NAND U14509 ( .A(x[499]), .B(y[7780]), .Z(n12386) );
  XOR U14510 ( .A(n12385), .B(n12386), .Z(n12367) );
  XOR U14511 ( .A(n12357), .B(n12356), .Z(n12425) );
  XOR U14512 ( .A(n12426), .B(n12425), .Z(n12428) );
  AND U14513 ( .A(x[500]), .B(y[7785]), .Z(n13280) );
  AND U14514 ( .A(x[493]), .B(y[7778]), .Z(n12263) );
  NAND U14515 ( .A(n13280), .B(n12263), .Z(n12267) );
  NAND U14516 ( .A(n12265), .B(n12264), .Z(n12266) );
  NAND U14517 ( .A(n12267), .B(n12266), .Z(n12420) );
  NAND U14518 ( .A(n12269), .B(n12268), .Z(n12273) );
  NAND U14519 ( .A(n12271), .B(n12270), .Z(n12272) );
  NAND U14520 ( .A(n12273), .B(n12272), .Z(n12375) );
  AND U14521 ( .A(x[493]), .B(y[7786]), .Z(n12348) );
  AND U14522 ( .A(x[482]), .B(y[7797]), .Z(n12349) );
  XOR U14523 ( .A(n12348), .B(n12349), .Z(n12350) );
  AND U14524 ( .A(x[501]), .B(y[7778]), .Z(n12351) );
  XOR U14525 ( .A(n12350), .B(n12351), .Z(n12373) );
  AND U14526 ( .A(x[492]), .B(y[7787]), .Z(n12403) );
  AND U14527 ( .A(x[481]), .B(y[7798]), .Z(n12404) );
  XOR U14528 ( .A(n12403), .B(n12404), .Z(n12406) );
  AND U14529 ( .A(o[118]), .B(n12274), .Z(n12405) );
  XOR U14530 ( .A(n12406), .B(n12405), .Z(n12372) );
  XOR U14531 ( .A(n12373), .B(n12372), .Z(n12374) );
  XOR U14532 ( .A(n12375), .B(n12374), .Z(n12419) );
  XOR U14533 ( .A(n12420), .B(n12419), .Z(n12422) );
  AND U14534 ( .A(x[495]), .B(y[7792]), .Z(n13528) );
  NAND U14535 ( .A(n13528), .B(n12275), .Z(n12279) );
  NANDN U14536 ( .A(n12277), .B(n12276), .Z(n12278) );
  NAND U14537 ( .A(n12279), .B(n12278), .Z(n12363) );
  AND U14538 ( .A(x[494]), .B(y[7785]), .Z(n12342) );
  AND U14539 ( .A(x[483]), .B(y[7796]), .Z(n12343) );
  XOR U14540 ( .A(n12342), .B(n12343), .Z(n12344) );
  AND U14541 ( .A(x[484]), .B(y[7795]), .Z(n12345) );
  XOR U14542 ( .A(n12344), .B(n12345), .Z(n12360) );
  AND U14543 ( .A(x[485]), .B(y[7794]), .Z(n12336) );
  NAND U14544 ( .A(x[498]), .B(y[7781]), .Z(n12337) );
  XNOR U14545 ( .A(n12336), .B(n12337), .Z(n12338) );
  NAND U14546 ( .A(x[497]), .B(y[7782]), .Z(n12339) );
  XNOR U14547 ( .A(n12338), .B(n12339), .Z(n12361) );
  XOR U14548 ( .A(n12360), .B(n12361), .Z(n12362) );
  XOR U14549 ( .A(n12363), .B(n12362), .Z(n12421) );
  XOR U14550 ( .A(n12422), .B(n12421), .Z(n12427) );
  XOR U14551 ( .A(n12428), .B(n12427), .Z(n12431) );
  XOR U14552 ( .A(n12432), .B(n12431), .Z(n12433) );
  XOR U14553 ( .A(n12434), .B(n12433), .Z(n12321) );
  NAND U14554 ( .A(n12281), .B(n12280), .Z(n12285) );
  NAND U14555 ( .A(n12283), .B(n12282), .Z(n12284) );
  NAND U14556 ( .A(n12285), .B(n12284), .Z(n12440) );
  NAND U14557 ( .A(n12287), .B(n12286), .Z(n12291) );
  NAND U14558 ( .A(n12289), .B(n12288), .Z(n12290) );
  NAND U14559 ( .A(n12291), .B(n12290), .Z(n12438) );
  NAND U14560 ( .A(n12293), .B(n12292), .Z(n12297) );
  NAND U14561 ( .A(n12295), .B(n12294), .Z(n12296) );
  AND U14562 ( .A(n12297), .B(n12296), .Z(n12437) );
  XOR U14563 ( .A(n12438), .B(n12437), .Z(n12439) );
  XOR U14564 ( .A(n12440), .B(n12439), .Z(n12319) );
  NAND U14565 ( .A(n12299), .B(n12298), .Z(n12303) );
  NANDN U14566 ( .A(n12301), .B(n12300), .Z(n12302) );
  AND U14567 ( .A(n12303), .B(n12302), .Z(n12318) );
  XOR U14568 ( .A(n12306), .B(n12305), .Z(n12307) );
  XOR U14569 ( .A(n12308), .B(n12307), .Z(n12314) );
  XNOR U14570 ( .A(n12313), .B(n12314), .Z(n12304) );
  XOR U14571 ( .A(n12311), .B(n12304), .Z(N248) );
  NAND U14572 ( .A(n12306), .B(n12305), .Z(n12310) );
  NAND U14573 ( .A(n12308), .B(n12307), .Z(n12309) );
  NAND U14574 ( .A(n12310), .B(n12309), .Z(n12569) );
  IV U14575 ( .A(n12569), .Z(n12567) );
  OR U14576 ( .A(n12313), .B(n12311), .Z(n12317) );
  ANDN U14577 ( .B(n12313), .A(n12312), .Z(n12315) );
  OR U14578 ( .A(n12315), .B(n12314), .Z(n12316) );
  AND U14579 ( .A(n12317), .B(n12316), .Z(n12568) );
  NANDN U14580 ( .A(n12319), .B(n12318), .Z(n12323) );
  NANDN U14581 ( .A(n12321), .B(n12320), .Z(n12322) );
  AND U14582 ( .A(n12323), .B(n12322), .Z(n12576) );
  NAND U14583 ( .A(n12325), .B(n12324), .Z(n12329) );
  NAND U14584 ( .A(n12327), .B(n12326), .Z(n12328) );
  NAND U14585 ( .A(n12329), .B(n12328), .Z(n12545) );
  NAND U14586 ( .A(n12331), .B(n12330), .Z(n12335) );
  NAND U14587 ( .A(n12333), .B(n12332), .Z(n12334) );
  NAND U14588 ( .A(n12335), .B(n12334), .Z(n12543) );
  NANDN U14589 ( .A(n12337), .B(n12336), .Z(n12341) );
  NANDN U14590 ( .A(n12339), .B(n12338), .Z(n12340) );
  NAND U14591 ( .A(n12341), .B(n12340), .Z(n12470) );
  AND U14592 ( .A(x[480]), .B(y[7800]), .Z(n12528) );
  AND U14593 ( .A(x[504]), .B(y[7776]), .Z(n12527) );
  XOR U14594 ( .A(n12528), .B(n12527), .Z(n12530) );
  AND U14595 ( .A(x[503]), .B(y[7777]), .Z(n12522) );
  XOR U14596 ( .A(n12522), .B(o[120]), .Z(n12529) );
  XOR U14597 ( .A(n12530), .B(n12529), .Z(n12469) );
  AND U14598 ( .A(x[487]), .B(y[7793]), .Z(n12516) );
  NAND U14599 ( .A(x[498]), .B(y[7782]), .Z(n12517) );
  XNOR U14600 ( .A(n12516), .B(n12517), .Z(n12519) );
  AND U14601 ( .A(x[497]), .B(y[7783]), .Z(n12518) );
  XOR U14602 ( .A(n12519), .B(n12518), .Z(n12468) );
  XOR U14603 ( .A(n12469), .B(n12468), .Z(n12471) );
  XOR U14604 ( .A(n12470), .B(n12471), .Z(n12459) );
  NAND U14605 ( .A(n12343), .B(n12342), .Z(n12347) );
  NAND U14606 ( .A(n12345), .B(n12344), .Z(n12346) );
  NAND U14607 ( .A(n12347), .B(n12346), .Z(n12457) );
  NAND U14608 ( .A(n12349), .B(n12348), .Z(n12353) );
  NAND U14609 ( .A(n12351), .B(n12350), .Z(n12352) );
  NAND U14610 ( .A(n12353), .B(n12352), .Z(n12456) );
  XOR U14611 ( .A(n12457), .B(n12456), .Z(n12458) );
  XOR U14612 ( .A(n12459), .B(n12458), .Z(n12544) );
  XOR U14613 ( .A(n12543), .B(n12544), .Z(n12546) );
  XNOR U14614 ( .A(n12545), .B(n12546), .Z(n12452) );
  NAND U14615 ( .A(n12355), .B(n12354), .Z(n12359) );
  NAND U14616 ( .A(n12357), .B(n12356), .Z(n12358) );
  AND U14617 ( .A(n12359), .B(n12358), .Z(n12493) );
  NAND U14618 ( .A(n12361), .B(n12360), .Z(n12365) );
  NAND U14619 ( .A(n12363), .B(n12362), .Z(n12364) );
  AND U14620 ( .A(n12365), .B(n12364), .Z(n12490) );
  NANDN U14621 ( .A(n12367), .B(n12366), .Z(n12371) );
  NANDN U14622 ( .A(n12369), .B(n12368), .Z(n12370) );
  NAND U14623 ( .A(n12371), .B(n12370), .Z(n12491) );
  XOR U14624 ( .A(n12493), .B(n12492), .Z(n12450) );
  NAND U14625 ( .A(n12373), .B(n12372), .Z(n12377) );
  NAND U14626 ( .A(n12375), .B(n12374), .Z(n12376) );
  AND U14627 ( .A(n12377), .B(n12376), .Z(n12451) );
  XOR U14628 ( .A(n12450), .B(n12451), .Z(n12453) );
  XOR U14629 ( .A(n12452), .B(n12453), .Z(n12555) );
  NAND U14630 ( .A(n12379), .B(n12378), .Z(n12383) );
  NAND U14631 ( .A(n12381), .B(n12380), .Z(n12382) );
  AND U14632 ( .A(n12383), .B(n12382), .Z(n12556) );
  XOR U14633 ( .A(n12555), .B(n12556), .Z(n12558) );
  AND U14634 ( .A(x[500]), .B(y[7783]), .Z(n12384) );
  NAND U14635 ( .A(n12472), .B(n12384), .Z(n12388) );
  NANDN U14636 ( .A(n12386), .B(n12385), .Z(n12387) );
  AND U14637 ( .A(n12388), .B(n12387), .Z(n12489) );
  AND U14638 ( .A(x[502]), .B(y[7778]), .Z(n12506) );
  XOR U14639 ( .A(n12507), .B(n12506), .Z(n12504) );
  NAND U14640 ( .A(x[482]), .B(y[7798]), .Z(n12505) );
  XNOR U14641 ( .A(n12504), .B(n12505), .Z(n12487) );
  AND U14642 ( .A(x[481]), .B(y[7799]), .Z(n12512) );
  XOR U14643 ( .A(n12513), .B(n12512), .Z(n12511) );
  NAND U14644 ( .A(n12389), .B(o[119]), .Z(n12510) );
  XNOR U14645 ( .A(n12511), .B(n12510), .Z(n12486) );
  XOR U14646 ( .A(n12487), .B(n12486), .Z(n12488) );
  XNOR U14647 ( .A(n12489), .B(n12488), .Z(n12538) );
  NANDN U14648 ( .A(n12391), .B(n12390), .Z(n12395) );
  NAND U14649 ( .A(n12393), .B(n12392), .Z(n12394) );
  NAND U14650 ( .A(n12395), .B(n12394), .Z(n12484) );
  AND U14651 ( .A(y[7784]), .B(x[496]), .Z(n12397) );
  NAND U14652 ( .A(y[7779]), .B(x[501]), .Z(n12396) );
  XNOR U14653 ( .A(n12397), .B(n12396), .Z(n12474) );
  AND U14654 ( .A(x[485]), .B(y[7795]), .Z(n12473) );
  XOR U14655 ( .A(n12474), .B(n12473), .Z(n12483) );
  AND U14656 ( .A(x[500]), .B(y[7780]), .Z(n12686) );
  AND U14657 ( .A(x[486]), .B(y[7794]), .Z(n12477) );
  XOR U14658 ( .A(n12686), .B(n12477), .Z(n12479) );
  AND U14659 ( .A(x[499]), .B(y[7781]), .Z(n12478) );
  XOR U14660 ( .A(n12479), .B(n12478), .Z(n12482) );
  XOR U14661 ( .A(n12483), .B(n12482), .Z(n12485) );
  XOR U14662 ( .A(n12484), .B(n12485), .Z(n12465) );
  NANDN U14663 ( .A(n12617), .B(n12398), .Z(n12402) );
  NANDN U14664 ( .A(n12400), .B(n12399), .Z(n12401) );
  NAND U14665 ( .A(n12402), .B(n12401), .Z(n12463) );
  NAND U14666 ( .A(n12404), .B(n12403), .Z(n12408) );
  NAND U14667 ( .A(n12406), .B(n12405), .Z(n12407) );
  NAND U14668 ( .A(n12408), .B(n12407), .Z(n12462) );
  XOR U14669 ( .A(n12463), .B(n12462), .Z(n12464) );
  XOR U14670 ( .A(n12465), .B(n12464), .Z(n12537) );
  XOR U14671 ( .A(n12538), .B(n12537), .Z(n12540) );
  NAND U14672 ( .A(n12410), .B(n12409), .Z(n12414) );
  NAND U14673 ( .A(n12412), .B(n12411), .Z(n12413) );
  NAND U14674 ( .A(n12414), .B(n12413), .Z(n12531) );
  AND U14675 ( .A(x[483]), .B(y[7797]), .Z(n12523) );
  XOR U14676 ( .A(n12524), .B(n12523), .Z(n12526) );
  AND U14677 ( .A(x[484]), .B(y[7796]), .Z(n12525) );
  XOR U14678 ( .A(n12526), .B(n12525), .Z(n12532) );
  XOR U14679 ( .A(n12531), .B(n12532), .Z(n12534) );
  AND U14680 ( .A(y[7791]), .B(x[489]), .Z(n12416) );
  NAND U14681 ( .A(y[7790]), .B(x[490]), .Z(n12415) );
  XNOR U14682 ( .A(n12416), .B(n12415), .Z(n12498) );
  AND U14683 ( .A(y[7786]), .B(x[494]), .Z(n12418) );
  NAND U14684 ( .A(y[7792]), .B(x[488]), .Z(n12417) );
  XNOR U14685 ( .A(n12418), .B(n12417), .Z(n12503) );
  AND U14686 ( .A(x[491]), .B(y[7789]), .Z(n12502) );
  XOR U14687 ( .A(n12503), .B(n12502), .Z(n12497) );
  XOR U14688 ( .A(n12498), .B(n12497), .Z(n12533) );
  XOR U14689 ( .A(n12534), .B(n12533), .Z(n12539) );
  XNOR U14690 ( .A(n12540), .B(n12539), .Z(n12550) );
  NAND U14691 ( .A(n12420), .B(n12419), .Z(n12424) );
  NAND U14692 ( .A(n12422), .B(n12421), .Z(n12423) );
  AND U14693 ( .A(n12424), .B(n12423), .Z(n12549) );
  XOR U14694 ( .A(n12550), .B(n12549), .Z(n12551) );
  NAND U14695 ( .A(n12426), .B(n12425), .Z(n12430) );
  NAND U14696 ( .A(n12428), .B(n12427), .Z(n12429) );
  AND U14697 ( .A(n12430), .B(n12429), .Z(n12552) );
  XOR U14698 ( .A(n12551), .B(n12552), .Z(n12557) );
  XNOR U14699 ( .A(n12558), .B(n12557), .Z(n12574) );
  NAND U14700 ( .A(n12432), .B(n12431), .Z(n12436) );
  NAND U14701 ( .A(n12434), .B(n12433), .Z(n12435) );
  NAND U14702 ( .A(n12436), .B(n12435), .Z(n12564) );
  NAND U14703 ( .A(n12438), .B(n12437), .Z(n12442) );
  NAND U14704 ( .A(n12440), .B(n12439), .Z(n12441) );
  NAND U14705 ( .A(n12442), .B(n12441), .Z(n12562) );
  NAND U14706 ( .A(n12444), .B(n12443), .Z(n12448) );
  NAND U14707 ( .A(n12446), .B(n12445), .Z(n12447) );
  NAND U14708 ( .A(n12448), .B(n12447), .Z(n12561) );
  XOR U14709 ( .A(n12562), .B(n12561), .Z(n12563) );
  XNOR U14710 ( .A(n12564), .B(n12563), .Z(n12575) );
  XOR U14711 ( .A(n12574), .B(n12575), .Z(n12577) );
  XNOR U14712 ( .A(n12576), .B(n12577), .Z(n12570) );
  XNOR U14713 ( .A(n12568), .B(n12570), .Z(n12449) );
  XOR U14714 ( .A(n12567), .B(n12449), .Z(N249) );
  NAND U14715 ( .A(n12451), .B(n12450), .Z(n12455) );
  NAND U14716 ( .A(n12453), .B(n12452), .Z(n12454) );
  AND U14717 ( .A(n12455), .B(n12454), .Z(n12590) );
  NAND U14718 ( .A(n12457), .B(n12456), .Z(n12461) );
  NAND U14719 ( .A(n12459), .B(n12458), .Z(n12460) );
  NAND U14720 ( .A(n12461), .B(n12460), .Z(n12606) );
  NAND U14721 ( .A(n12463), .B(n12462), .Z(n12467) );
  NAND U14722 ( .A(n12465), .B(n12464), .Z(n12466) );
  NAND U14723 ( .A(n12467), .B(n12466), .Z(n12605) );
  XOR U14724 ( .A(n12606), .B(n12605), .Z(n12608) );
  AND U14725 ( .A(x[501]), .B(y[7784]), .Z(n13429) );
  NAND U14726 ( .A(x[502]), .B(y[7779]), .Z(n12675) );
  NAND U14727 ( .A(x[485]), .B(y[7796]), .Z(n12674) );
  NAND U14728 ( .A(x[497]), .B(y[7784]), .Z(n12673) );
  XOR U14729 ( .A(n12674), .B(n12673), .Z(n12676) );
  XOR U14730 ( .A(n12675), .B(n12676), .Z(n12702) );
  AND U14731 ( .A(y[7781]), .B(x[500]), .Z(n12476) );
  NAND U14732 ( .A(y[7780]), .B(x[501]), .Z(n12475) );
  XNOR U14733 ( .A(n12476), .B(n12475), .Z(n12688) );
  AND U14734 ( .A(x[499]), .B(y[7782]), .Z(n12687) );
  XOR U14735 ( .A(n12688), .B(n12687), .Z(n12701) );
  XNOR U14736 ( .A(n12702), .B(n12701), .Z(n12704) );
  XOR U14737 ( .A(n12703), .B(n12704), .Z(n12634) );
  IV U14738 ( .A(n12477), .Z(n12859) );
  NANDN U14739 ( .A(n12859), .B(n12686), .Z(n12481) );
  NAND U14740 ( .A(n12479), .B(n12478), .Z(n12480) );
  NAND U14741 ( .A(n12481), .B(n12480), .Z(n12707) );
  NAND U14742 ( .A(x[495]), .B(y[7786]), .Z(n12693) );
  NAND U14743 ( .A(x[498]), .B(y[7783]), .Z(n12692) );
  NAND U14744 ( .A(x[486]), .B(y[7795]), .Z(n12691) );
  XOR U14745 ( .A(n12692), .B(n12691), .Z(n12694) );
  XOR U14746 ( .A(n12693), .B(n12694), .Z(n12706) );
  NAND U14747 ( .A(x[503]), .B(y[7778]), .Z(n12669) );
  NAND U14748 ( .A(x[484]), .B(y[7797]), .Z(n12668) );
  NAND U14749 ( .A(x[496]), .B(y[7785]), .Z(n12667) );
  XNOR U14750 ( .A(n12668), .B(n12667), .Z(n12670) );
  XOR U14751 ( .A(n12669), .B(n12670), .Z(n12705) );
  XNOR U14752 ( .A(n12706), .B(n12705), .Z(n12708) );
  XOR U14753 ( .A(n12707), .B(n12708), .Z(n12633) );
  XNOR U14754 ( .A(n12634), .B(n12633), .Z(n12636) );
  XNOR U14755 ( .A(n12635), .B(n12636), .Z(n12646) );
  XOR U14756 ( .A(n12643), .B(n12644), .Z(n12645) );
  XNOR U14757 ( .A(n12646), .B(n12645), .Z(n12607) );
  XOR U14758 ( .A(n12608), .B(n12607), .Z(n12588) );
  NANDN U14759 ( .A(n12491), .B(n12490), .Z(n12495) );
  NAND U14760 ( .A(n12493), .B(n12492), .Z(n12494) );
  NAND U14761 ( .A(n12495), .B(n12494), .Z(n12587) );
  NANDN U14762 ( .A(n12618), .B(n12496), .Z(n12500) );
  NAND U14763 ( .A(n12498), .B(n12497), .Z(n12499) );
  NAND U14764 ( .A(n12500), .B(n12499), .Z(n12639) );
  AND U14765 ( .A(x[494]), .B(y[7792]), .Z(n13505) );
  NAND U14766 ( .A(x[491]), .B(y[7790]), .Z(n12682) );
  NAND U14767 ( .A(x[492]), .B(y[7789]), .Z(n12681) );
  NAND U14768 ( .A(x[487]), .B(y[7794]), .Z(n12680) );
  XOR U14769 ( .A(n12681), .B(n12680), .Z(n12683) );
  XNOR U14770 ( .A(n12682), .B(n12683), .Z(n12662) );
  AND U14771 ( .A(x[504]), .B(y[7777]), .Z(n12679) );
  XOR U14772 ( .A(o[121]), .B(n12679), .Z(n12650) );
  AND U14773 ( .A(x[481]), .B(y[7800]), .Z(n12649) );
  XOR U14774 ( .A(n12650), .B(n12649), .Z(n12652) );
  AND U14775 ( .A(x[493]), .B(y[7788]), .Z(n12651) );
  XOR U14776 ( .A(n12652), .B(n12651), .Z(n12661) );
  XOR U14777 ( .A(n12662), .B(n12661), .Z(n12664) );
  XOR U14778 ( .A(n12663), .B(n12664), .Z(n12640) );
  XOR U14779 ( .A(n12639), .B(n12640), .Z(n12642) );
  NANDN U14780 ( .A(n12505), .B(n12504), .Z(n12509) );
  AND U14781 ( .A(n12507), .B(n12506), .Z(n12508) );
  ANDN U14782 ( .B(n12509), .A(n12508), .Z(n12628) );
  ANDN U14783 ( .B(n12511), .A(n12510), .Z(n12515) );
  NAND U14784 ( .A(n12513), .B(n12512), .Z(n12514) );
  NANDN U14785 ( .A(n12515), .B(n12514), .Z(n12627) );
  XNOR U14786 ( .A(n12628), .B(n12627), .Z(n12630) );
  NANDN U14787 ( .A(n12517), .B(n12516), .Z(n12521) );
  NAND U14788 ( .A(n12519), .B(n12518), .Z(n12520) );
  AND U14789 ( .A(n12521), .B(n12520), .Z(n12624) );
  NAND U14790 ( .A(x[488]), .B(y[7793]), .Z(n12619) );
  XOR U14791 ( .A(n12617), .B(n12618), .Z(n12620) );
  XOR U14792 ( .A(n12619), .B(n12620), .Z(n12622) );
  NAND U14793 ( .A(n12522), .B(o[120]), .Z(n12613) );
  NAND U14794 ( .A(x[505]), .B(y[7776]), .Z(n12612) );
  NAND U14795 ( .A(x[480]), .B(y[7801]), .Z(n12611) );
  XNOR U14796 ( .A(n12612), .B(n12611), .Z(n12614) );
  XOR U14797 ( .A(n12613), .B(n12614), .Z(n12621) );
  XNOR U14798 ( .A(n12622), .B(n12621), .Z(n12623) );
  XNOR U14799 ( .A(n12624), .B(n12623), .Z(n12629) );
  XOR U14800 ( .A(n12630), .B(n12629), .Z(n12641) );
  XNOR U14801 ( .A(n12642), .B(n12641), .Z(n12596) );
  AND U14802 ( .A(x[494]), .B(y[7787]), .Z(n12656) );
  AND U14803 ( .A(x[482]), .B(y[7799]), .Z(n12655) );
  XOR U14804 ( .A(n12656), .B(n12655), .Z(n12658) );
  AND U14805 ( .A(x[483]), .B(y[7798]), .Z(n12657) );
  XOR U14806 ( .A(n12658), .B(n12657), .Z(n12698) );
  XOR U14807 ( .A(n12697), .B(n12698), .Z(n12700) );
  XNOR U14808 ( .A(n12699), .B(n12700), .Z(n12594) );
  NAND U14809 ( .A(n12532), .B(n12531), .Z(n12536) );
  NAND U14810 ( .A(n12534), .B(n12533), .Z(n12535) );
  AND U14811 ( .A(n12536), .B(n12535), .Z(n12593) );
  XOR U14812 ( .A(n12594), .B(n12593), .Z(n12595) );
  XOR U14813 ( .A(n12596), .B(n12595), .Z(n12600) );
  NAND U14814 ( .A(n12538), .B(n12537), .Z(n12542) );
  NAND U14815 ( .A(n12540), .B(n12539), .Z(n12541) );
  AND U14816 ( .A(n12542), .B(n12541), .Z(n12599) );
  XOR U14817 ( .A(n12600), .B(n12599), .Z(n12602) );
  NAND U14818 ( .A(n12544), .B(n12543), .Z(n12548) );
  NAND U14819 ( .A(n12546), .B(n12545), .Z(n12547) );
  AND U14820 ( .A(n12548), .B(n12547), .Z(n12601) );
  XOR U14821 ( .A(n12602), .B(n12601), .Z(n12582) );
  NAND U14822 ( .A(n12550), .B(n12549), .Z(n12554) );
  NAND U14823 ( .A(n12552), .B(n12551), .Z(n12553) );
  AND U14824 ( .A(n12554), .B(n12553), .Z(n12581) );
  XNOR U14825 ( .A(n12583), .B(n12584), .Z(n12713) );
  NAND U14826 ( .A(n12556), .B(n12555), .Z(n12560) );
  NAND U14827 ( .A(n12558), .B(n12557), .Z(n12559) );
  NAND U14828 ( .A(n12560), .B(n12559), .Z(n12712) );
  XOR U14829 ( .A(n12713), .B(n12712), .Z(n12715) );
  NAND U14830 ( .A(n12562), .B(n12561), .Z(n12566) );
  NAND U14831 ( .A(n12564), .B(n12563), .Z(n12565) );
  AND U14832 ( .A(n12566), .B(n12565), .Z(n12714) );
  XNOR U14833 ( .A(n12715), .B(n12714), .Z(n12711) );
  NANDN U14834 ( .A(n12567), .B(n12568), .Z(n12573) );
  NOR U14835 ( .A(n12569), .B(n12568), .Z(n12571) );
  OR U14836 ( .A(n12571), .B(n12570), .Z(n12572) );
  AND U14837 ( .A(n12573), .B(n12572), .Z(n12710) );
  NANDN U14838 ( .A(n12575), .B(n12574), .Z(n12579) );
  NANDN U14839 ( .A(n12577), .B(n12576), .Z(n12578) );
  AND U14840 ( .A(n12579), .B(n12578), .Z(n12709) );
  XOR U14841 ( .A(n12710), .B(n12709), .Z(n12580) );
  XNOR U14842 ( .A(n12711), .B(n12580), .Z(N250) );
  NANDN U14843 ( .A(n12582), .B(n12581), .Z(n12586) );
  NAND U14844 ( .A(n12584), .B(n12583), .Z(n12585) );
  AND U14845 ( .A(n12586), .B(n12585), .Z(n12720) );
  NANDN U14846 ( .A(n12588), .B(n12587), .Z(n12592) );
  NANDN U14847 ( .A(n12590), .B(n12589), .Z(n12591) );
  AND U14848 ( .A(n12592), .B(n12591), .Z(n12719) );
  NAND U14849 ( .A(n12594), .B(n12593), .Z(n12598) );
  NAND U14850 ( .A(n12596), .B(n12595), .Z(n12597) );
  AND U14851 ( .A(n12598), .B(n12597), .Z(n12729) );
  NAND U14852 ( .A(n12600), .B(n12599), .Z(n12604) );
  NAND U14853 ( .A(n12602), .B(n12601), .Z(n12603) );
  AND U14854 ( .A(n12604), .B(n12603), .Z(n12728) );
  XOR U14855 ( .A(n12729), .B(n12728), .Z(n12730) );
  NAND U14856 ( .A(n12606), .B(n12605), .Z(n12610) );
  NAND U14857 ( .A(n12608), .B(n12607), .Z(n12609) );
  NAND U14858 ( .A(n12610), .B(n12609), .Z(n12736) );
  AND U14859 ( .A(x[482]), .B(y[7800]), .Z(n12756) );
  XOR U14860 ( .A(n12757), .B(n12756), .Z(n12759) );
  AND U14861 ( .A(x[504]), .B(y[7778]), .Z(n12758) );
  XOR U14862 ( .A(n12759), .B(n12758), .Z(n12793) );
  NAND U14863 ( .A(n12612), .B(n12611), .Z(n12616) );
  NANDN U14864 ( .A(n12614), .B(n12613), .Z(n12615) );
  AND U14865 ( .A(n12616), .B(n12615), .Z(n12792) );
  XOR U14866 ( .A(n12793), .B(n12792), .Z(n12795) );
  XOR U14867 ( .A(n12795), .B(n12794), .Z(n12828) );
  NANDN U14868 ( .A(n12622), .B(n12621), .Z(n12626) );
  NANDN U14869 ( .A(n12624), .B(n12623), .Z(n12625) );
  AND U14870 ( .A(n12626), .B(n12625), .Z(n12827) );
  XNOR U14871 ( .A(n12828), .B(n12827), .Z(n12829) );
  NANDN U14872 ( .A(n12628), .B(n12627), .Z(n12632) );
  NAND U14873 ( .A(n12630), .B(n12629), .Z(n12631) );
  NAND U14874 ( .A(n12632), .B(n12631), .Z(n12830) );
  XNOR U14875 ( .A(n12829), .B(n12830), .Z(n12825) );
  OR U14876 ( .A(n12634), .B(n12633), .Z(n12638) );
  NANDN U14877 ( .A(n12636), .B(n12635), .Z(n12637) );
  NAND U14878 ( .A(n12638), .B(n12637), .Z(n12824) );
  XNOR U14879 ( .A(n12824), .B(n12823), .Z(n12826) );
  XOR U14880 ( .A(n12825), .B(n12826), .Z(n12734) );
  AND U14881 ( .A(x[492]), .B(y[7790]), .Z(n12922) );
  AND U14882 ( .A(x[485]), .B(y[7797]), .Z(n12806) );
  XOR U14883 ( .A(n12922), .B(n12806), .Z(n12808) );
  AND U14884 ( .A(x[490]), .B(y[7792]), .Z(n12807) );
  XOR U14885 ( .A(n12808), .B(n12807), .Z(n12835) );
  AND U14886 ( .A(y[7796]), .B(x[486]), .Z(n12648) );
  NAND U14887 ( .A(y[7794]), .B(x[488]), .Z(n12647) );
  XNOR U14888 ( .A(n12648), .B(n12647), .Z(n12861) );
  AND U14889 ( .A(x[489]), .B(y[7793]), .Z(n12860) );
  XOR U14890 ( .A(n12861), .B(n12860), .Z(n12834) );
  AND U14891 ( .A(x[487]), .B(y[7795]), .Z(n12833) );
  XNOR U14892 ( .A(n12834), .B(n12833), .Z(n12836) );
  XNOR U14893 ( .A(n12835), .B(n12836), .Z(n12782) );
  NAND U14894 ( .A(n12650), .B(n12649), .Z(n12654) );
  NAND U14895 ( .A(n12652), .B(n12651), .Z(n12653) );
  NAND U14896 ( .A(n12654), .B(n12653), .Z(n12781) );
  NAND U14897 ( .A(n12656), .B(n12655), .Z(n12660) );
  NAND U14898 ( .A(n12658), .B(n12657), .Z(n12659) );
  NAND U14899 ( .A(n12660), .B(n12659), .Z(n12780) );
  XOR U14900 ( .A(n12781), .B(n12780), .Z(n12783) );
  XNOR U14901 ( .A(n12782), .B(n12783), .Z(n12818) );
  NAND U14902 ( .A(n12662), .B(n12661), .Z(n12666) );
  NAND U14903 ( .A(n12664), .B(n12663), .Z(n12665) );
  AND U14904 ( .A(n12666), .B(n12665), .Z(n12817) );
  XOR U14905 ( .A(n12818), .B(n12817), .Z(n12819) );
  NAND U14906 ( .A(n12668), .B(n12667), .Z(n12672) );
  NANDN U14907 ( .A(n12670), .B(n12669), .Z(n12671) );
  AND U14908 ( .A(n12672), .B(n12671), .Z(n12745) );
  NAND U14909 ( .A(n12674), .B(n12673), .Z(n12678) );
  NAND U14910 ( .A(n12676), .B(n12675), .Z(n12677) );
  AND U14911 ( .A(n12678), .B(n12677), .Z(n12744) );
  XOR U14912 ( .A(n12745), .B(n12744), .Z(n12747) );
  NAND U14913 ( .A(x[494]), .B(y[7788]), .Z(n12854) );
  XNOR U14914 ( .A(n12853), .B(n12854), .Z(n12855) );
  NAND U14915 ( .A(x[481]), .B(y[7801]), .Z(n12856) );
  XNOR U14916 ( .A(n12855), .B(n12856), .Z(n12799) );
  NAND U14917 ( .A(x[505]), .B(y[7777]), .Z(n12864) );
  XNOR U14918 ( .A(o[122]), .B(n12864), .Z(n12812) );
  AND U14919 ( .A(x[506]), .B(y[7776]), .Z(n12811) );
  XOR U14920 ( .A(n12812), .B(n12811), .Z(n12814) );
  AND U14921 ( .A(x[480]), .B(y[7802]), .Z(n12813) );
  XOR U14922 ( .A(n12814), .B(n12813), .Z(n12798) );
  XOR U14923 ( .A(n12799), .B(n12798), .Z(n12801) );
  NAND U14924 ( .A(n12681), .B(n12680), .Z(n12685) );
  NAND U14925 ( .A(n12683), .B(n12682), .Z(n12684) );
  AND U14926 ( .A(n12685), .B(n12684), .Z(n12800) );
  XOR U14927 ( .A(n12801), .B(n12800), .Z(n12746) );
  XNOR U14928 ( .A(n12747), .B(n12746), .Z(n12788) );
  AND U14929 ( .A(x[501]), .B(y[7781]), .Z(n12848) );
  NAND U14930 ( .A(n12848), .B(n12686), .Z(n12690) );
  NAND U14931 ( .A(n12688), .B(n12687), .Z(n12689) );
  NAND U14932 ( .A(n12690), .B(n12689), .Z(n12776) );
  XOR U14933 ( .A(n12848), .B(n12847), .Z(n12849) );
  NAND U14934 ( .A(x[500]), .B(y[7782]), .Z(n12850) );
  XNOR U14935 ( .A(n12849), .B(n12850), .Z(n12775) );
  AND U14936 ( .A(x[503]), .B(y[7779]), .Z(n12762) );
  XOR U14937 ( .A(n12763), .B(n12762), .Z(n12765) );
  AND U14938 ( .A(x[502]), .B(y[7780]), .Z(n12764) );
  XOR U14939 ( .A(n12765), .B(n12764), .Z(n12774) );
  XOR U14940 ( .A(n12775), .B(n12774), .Z(n12777) );
  XNOR U14941 ( .A(n12776), .B(n12777), .Z(n12787) );
  AND U14942 ( .A(x[484]), .B(y[7798]), .Z(n12768) );
  XOR U14943 ( .A(n12769), .B(n12768), .Z(n12771) );
  XOR U14944 ( .A(n12771), .B(n12770), .Z(n12751) );
  AND U14945 ( .A(x[491]), .B(y[7791]), .Z(n12839) );
  NAND U14946 ( .A(x[483]), .B(y[7799]), .Z(n12840) );
  XNOR U14947 ( .A(n12839), .B(n12840), .Z(n12842) );
  AND U14948 ( .A(x[499]), .B(y[7783]), .Z(n12841) );
  XOR U14949 ( .A(n12842), .B(n12841), .Z(n12750) );
  XOR U14950 ( .A(n12751), .B(n12750), .Z(n12753) );
  NAND U14951 ( .A(n12692), .B(n12691), .Z(n12696) );
  NAND U14952 ( .A(n12694), .B(n12693), .Z(n12695) );
  AND U14953 ( .A(n12696), .B(n12695), .Z(n12752) );
  XNOR U14954 ( .A(n12753), .B(n12752), .Z(n12786) );
  XNOR U14955 ( .A(n12787), .B(n12786), .Z(n12789) );
  XOR U14956 ( .A(n12788), .B(n12789), .Z(n12820) );
  XNOR U14957 ( .A(n12819), .B(n12820), .Z(n12740) );
  XOR U14958 ( .A(n12866), .B(n12865), .Z(n12868) );
  XOR U14959 ( .A(n12867), .B(n12868), .Z(n12741) );
  XOR U14960 ( .A(n12740), .B(n12741), .Z(n12742) );
  XNOR U14961 ( .A(n12743), .B(n12742), .Z(n12735) );
  XOR U14962 ( .A(n12734), .B(n12735), .Z(n12737) );
  XOR U14963 ( .A(n12736), .B(n12737), .Z(n12731) );
  XNOR U14964 ( .A(n12730), .B(n12731), .Z(n12721) );
  XNOR U14965 ( .A(n12722), .B(n12721), .Z(n12727) );
  NAND U14966 ( .A(n12713), .B(n12712), .Z(n12717) );
  NAND U14967 ( .A(n12715), .B(n12714), .Z(n12716) );
  AND U14968 ( .A(n12717), .B(n12716), .Z(n12726) );
  XOR U14969 ( .A(n12725), .B(n12726), .Z(n12718) );
  XNOR U14970 ( .A(n12727), .B(n12718), .Z(N251) );
  NANDN U14971 ( .A(n12720), .B(n12719), .Z(n12724) );
  NAND U14972 ( .A(n12722), .B(n12721), .Z(n12723) );
  NAND U14973 ( .A(n12724), .B(n12723), .Z(n13026) );
  IV U14974 ( .A(n13026), .Z(n13025) );
  NAND U14975 ( .A(n12729), .B(n12728), .Z(n12733) );
  NANDN U14976 ( .A(n12731), .B(n12730), .Z(n12732) );
  AND U14977 ( .A(n12733), .B(n12732), .Z(n13022) );
  NANDN U14978 ( .A(n12735), .B(n12734), .Z(n12739) );
  NANDN U14979 ( .A(n12737), .B(n12736), .Z(n12738) );
  AND U14980 ( .A(n12739), .B(n12738), .Z(n13020) );
  NAND U14981 ( .A(n12745), .B(n12744), .Z(n12749) );
  NAND U14982 ( .A(n12747), .B(n12746), .Z(n12748) );
  NAND U14983 ( .A(n12749), .B(n12748), .Z(n12997) );
  NAND U14984 ( .A(n12751), .B(n12750), .Z(n12755) );
  NAND U14985 ( .A(n12753), .B(n12752), .Z(n12754) );
  NAND U14986 ( .A(n12755), .B(n12754), .Z(n12995) );
  AND U14987 ( .A(n12757), .B(n12756), .Z(n12761) );
  NAND U14988 ( .A(n12759), .B(n12758), .Z(n12760) );
  NANDN U14989 ( .A(n12761), .B(n12760), .Z(n12895) );
  NAND U14990 ( .A(n12763), .B(n12762), .Z(n12767) );
  NAND U14991 ( .A(n12765), .B(n12764), .Z(n12766) );
  NAND U14992 ( .A(n12767), .B(n12766), .Z(n12894) );
  XOR U14993 ( .A(n12895), .B(n12894), .Z(n12896) );
  AND U14994 ( .A(n12769), .B(n12768), .Z(n12773) );
  NAND U14995 ( .A(n12771), .B(n12770), .Z(n12772) );
  NANDN U14996 ( .A(n12773), .B(n12772), .Z(n12908) );
  AND U14997 ( .A(x[480]), .B(y[7803]), .Z(n12984) );
  AND U14998 ( .A(x[507]), .B(y[7776]), .Z(n12983) );
  XOR U14999 ( .A(n12984), .B(n12983), .Z(n12986) );
  AND U15000 ( .A(x[506]), .B(y[7777]), .Z(n12968) );
  XOR U15001 ( .A(n12968), .B(o[123]), .Z(n12985) );
  XOR U15002 ( .A(n12986), .B(n12985), .Z(n12907) );
  AND U15003 ( .A(x[489]), .B(y[7794]), .Z(n12972) );
  AND U15004 ( .A(x[501]), .B(y[7782]), .Z(n12971) );
  XOR U15005 ( .A(n12972), .B(n12971), .Z(n12974) );
  AND U15006 ( .A(x[498]), .B(y[7785]), .Z(n12973) );
  XOR U15007 ( .A(n12974), .B(n12973), .Z(n12906) );
  XOR U15008 ( .A(n12907), .B(n12906), .Z(n12909) );
  XNOR U15009 ( .A(n12908), .B(n12909), .Z(n12897) );
  XOR U15010 ( .A(n12995), .B(n12996), .Z(n12998) );
  XOR U15011 ( .A(n12997), .B(n12998), .Z(n13016) );
  NAND U15012 ( .A(n12775), .B(n12774), .Z(n12779) );
  NAND U15013 ( .A(n12777), .B(n12776), .Z(n12778) );
  AND U15014 ( .A(n12779), .B(n12778), .Z(n13014) );
  NAND U15015 ( .A(n12781), .B(n12780), .Z(n12785) );
  NAND U15016 ( .A(n12783), .B(n12782), .Z(n12784) );
  AND U15017 ( .A(n12785), .B(n12784), .Z(n13013) );
  XOR U15018 ( .A(n13014), .B(n13013), .Z(n13015) );
  NAND U15019 ( .A(n12787), .B(n12786), .Z(n12791) );
  NANDN U15020 ( .A(n12789), .B(n12788), .Z(n12790) );
  AND U15021 ( .A(n12791), .B(n12790), .Z(n13001) );
  NAND U15022 ( .A(n12793), .B(n12792), .Z(n12797) );
  NAND U15023 ( .A(n12795), .B(n12794), .Z(n12796) );
  NAND U15024 ( .A(n12797), .B(n12796), .Z(n12991) );
  NAND U15025 ( .A(n12799), .B(n12798), .Z(n12803) );
  NAND U15026 ( .A(n12801), .B(n12800), .Z(n12802) );
  NAND U15027 ( .A(n12803), .B(n12802), .Z(n12989) );
  AND U15028 ( .A(x[495]), .B(y[7788]), .Z(n12928) );
  AND U15029 ( .A(x[482]), .B(y[7801]), .Z(n12927) );
  XOR U15030 ( .A(n12928), .B(n12927), .Z(n12930) );
  AND U15031 ( .A(x[483]), .B(y[7800]), .Z(n12929) );
  XOR U15032 ( .A(n12930), .B(n12929), .Z(n12952) );
  AND U15033 ( .A(x[499]), .B(y[7784]), .Z(n12963) );
  AND U15034 ( .A(x[505]), .B(y[7778]), .Z(n12962) );
  XOR U15035 ( .A(n12963), .B(n12962), .Z(n12965) );
  AND U15036 ( .A(x[486]), .B(y[7797]), .Z(n12964) );
  XOR U15037 ( .A(n12965), .B(n12964), .Z(n12951) );
  XOR U15038 ( .A(n12952), .B(n12951), .Z(n12953) );
  NAND U15039 ( .A(x[496]), .B(y[7787]), .Z(n12913) );
  XOR U15040 ( .A(n12913), .B(n12912), .Z(n12915) );
  XOR U15041 ( .A(n12914), .B(n12915), .Z(n12924) );
  AND U15042 ( .A(y[7790]), .B(x[493]), .Z(n12805) );
  AND U15043 ( .A(y[7791]), .B(x[492]), .Z(n12804) );
  XOR U15044 ( .A(n12805), .B(n12804), .Z(n12923) );
  XNOR U15045 ( .A(n12953), .B(n12954), .Z(n12891) );
  AND U15046 ( .A(n12922), .B(n12806), .Z(n12810) );
  NAND U15047 ( .A(n12808), .B(n12807), .Z(n12809) );
  NANDN U15048 ( .A(n12810), .B(n12809), .Z(n12889) );
  NAND U15049 ( .A(n12812), .B(n12811), .Z(n12816) );
  NAND U15050 ( .A(n12814), .B(n12813), .Z(n12815) );
  NAND U15051 ( .A(n12816), .B(n12815), .Z(n12888) );
  XOR U15052 ( .A(n12889), .B(n12888), .Z(n12890) );
  XOR U15053 ( .A(n12891), .B(n12890), .Z(n12990) );
  XNOR U15054 ( .A(n12989), .B(n12990), .Z(n12992) );
  XNOR U15055 ( .A(n13001), .B(n13002), .Z(n13004) );
  NAND U15056 ( .A(n12818), .B(n12817), .Z(n12822) );
  NANDN U15057 ( .A(n12820), .B(n12819), .Z(n12821) );
  AND U15058 ( .A(n12822), .B(n12821), .Z(n13003) );
  XOR U15059 ( .A(n13004), .B(n13003), .Z(n12872) );
  XOR U15060 ( .A(n12873), .B(n12872), .Z(n12875) );
  XOR U15061 ( .A(n12874), .B(n12875), .Z(n12881) );
  NANDN U15062 ( .A(n12828), .B(n12827), .Z(n12832) );
  NANDN U15063 ( .A(n12830), .B(n12829), .Z(n12831) );
  NAND U15064 ( .A(n12832), .B(n12831), .Z(n12882) );
  NAND U15065 ( .A(n12834), .B(n12833), .Z(n12838) );
  NANDN U15066 ( .A(n12836), .B(n12835), .Z(n12837) );
  AND U15067 ( .A(n12838), .B(n12837), .Z(n13009) );
  NANDN U15068 ( .A(n12840), .B(n12839), .Z(n12844) );
  NAND U15069 ( .A(n12842), .B(n12841), .Z(n12843) );
  NAND U15070 ( .A(n12844), .B(n12843), .Z(n12947) );
  AND U15071 ( .A(y[7779]), .B(x[504]), .Z(n12846) );
  NAND U15072 ( .A(y[7783]), .B(x[500]), .Z(n12845) );
  XNOR U15073 ( .A(n12846), .B(n12845), .Z(n12959) );
  AND U15074 ( .A(x[487]), .B(y[7796]), .Z(n12958) );
  XOR U15075 ( .A(n12959), .B(n12958), .Z(n12946) );
  AND U15076 ( .A(x[488]), .B(y[7795]), .Z(n12917) );
  AND U15077 ( .A(x[503]), .B(y[7780]), .Z(n12916) );
  XOR U15078 ( .A(n12917), .B(n12916), .Z(n12919) );
  AND U15079 ( .A(x[502]), .B(y[7781]), .Z(n12918) );
  XOR U15080 ( .A(n12919), .B(n12918), .Z(n12945) );
  XOR U15081 ( .A(n12946), .B(n12945), .Z(n12948) );
  XOR U15082 ( .A(n12947), .B(n12948), .Z(n13008) );
  AND U15083 ( .A(n12848), .B(n12847), .Z(n12852) );
  NANDN U15084 ( .A(n12850), .B(n12849), .Z(n12851) );
  NANDN U15085 ( .A(n12852), .B(n12851), .Z(n12940) );
  NANDN U15086 ( .A(n12854), .B(n12853), .Z(n12858) );
  NANDN U15087 ( .A(n12856), .B(n12855), .Z(n12857) );
  NAND U15088 ( .A(n12858), .B(n12857), .Z(n12939) );
  XOR U15089 ( .A(n12940), .B(n12939), .Z(n12941) );
  AND U15090 ( .A(y[7796]), .B(x[488]), .Z(n12970) );
  NANDN U15091 ( .A(n12859), .B(n12970), .Z(n12863) );
  NAND U15092 ( .A(n12861), .B(n12860), .Z(n12862) );
  NAND U15093 ( .A(n12863), .B(n12862), .Z(n12902) );
  ANDN U15094 ( .B(o[122]), .A(n12864), .Z(n12936) );
  AND U15095 ( .A(x[494]), .B(y[7789]), .Z(n12934) );
  AND U15096 ( .A(x[481]), .B(y[7802]), .Z(n12933) );
  XOR U15097 ( .A(n12934), .B(n12933), .Z(n12935) );
  XOR U15098 ( .A(n12936), .B(n12935), .Z(n12901) );
  AND U15099 ( .A(x[497]), .B(y[7786]), .Z(n12978) );
  AND U15100 ( .A(x[484]), .B(y[7799]), .Z(n12977) );
  XOR U15101 ( .A(n12978), .B(n12977), .Z(n12980) );
  AND U15102 ( .A(x[485]), .B(y[7798]), .Z(n12979) );
  XOR U15103 ( .A(n12980), .B(n12979), .Z(n12900) );
  XOR U15104 ( .A(n12901), .B(n12900), .Z(n12903) );
  XOR U15105 ( .A(n12902), .B(n12903), .Z(n12942) );
  XNOR U15106 ( .A(n12941), .B(n12942), .Z(n13007) );
  XNOR U15107 ( .A(n13009), .B(n13010), .Z(n12883) );
  XOR U15108 ( .A(n12882), .B(n12883), .Z(n12885) );
  NANDN U15109 ( .A(n12866), .B(n12865), .Z(n12870) );
  NANDN U15110 ( .A(n12868), .B(n12867), .Z(n12869) );
  AND U15111 ( .A(n12870), .B(n12869), .Z(n12884) );
  XOR U15112 ( .A(n12885), .B(n12884), .Z(n12879) );
  XOR U15113 ( .A(n12878), .B(n12879), .Z(n12880) );
  XNOR U15114 ( .A(n12881), .B(n12880), .Z(n13019) );
  XOR U15115 ( .A(n13020), .B(n13019), .Z(n13021) );
  XOR U15116 ( .A(n13022), .B(n13021), .Z(n13028) );
  XNOR U15117 ( .A(n13027), .B(n13028), .Z(n12871) );
  XOR U15118 ( .A(n13025), .B(n12871), .Z(N252) );
  NAND U15119 ( .A(n12873), .B(n12872), .Z(n12877) );
  NAND U15120 ( .A(n12875), .B(n12874), .Z(n12876) );
  NAND U15121 ( .A(n12877), .B(n12876), .Z(n13033) );
  XOR U15122 ( .A(n13033), .B(n13034), .Z(n13036) );
  NAND U15123 ( .A(n12883), .B(n12882), .Z(n12887) );
  NAND U15124 ( .A(n12885), .B(n12884), .Z(n12886) );
  AND U15125 ( .A(n12887), .B(n12886), .Z(n13040) );
  NAND U15126 ( .A(n12889), .B(n12888), .Z(n12893) );
  NAND U15127 ( .A(n12891), .B(n12890), .Z(n12892) );
  NAND U15128 ( .A(n12893), .B(n12892), .Z(n13052) );
  NAND U15129 ( .A(n12895), .B(n12894), .Z(n12899) );
  NANDN U15130 ( .A(n12897), .B(n12896), .Z(n12898) );
  NAND U15131 ( .A(n12899), .B(n12898), .Z(n13157) );
  NAND U15132 ( .A(n12901), .B(n12900), .Z(n12905) );
  NAND U15133 ( .A(n12903), .B(n12902), .Z(n12904) );
  NAND U15134 ( .A(n12905), .B(n12904), .Z(n13156) );
  NAND U15135 ( .A(n12907), .B(n12906), .Z(n12911) );
  NAND U15136 ( .A(n12909), .B(n12908), .Z(n12910) );
  NAND U15137 ( .A(n12911), .B(n12910), .Z(n13155) );
  XOR U15138 ( .A(n13156), .B(n13155), .Z(n13158) );
  XOR U15139 ( .A(n13157), .B(n13158), .Z(n13053) );
  XOR U15140 ( .A(n13052), .B(n13053), .Z(n13055) );
  AND U15141 ( .A(x[487]), .B(y[7797]), .Z(n13100) );
  AND U15142 ( .A(x[492]), .B(y[7792]), .Z(n13099) );
  XOR U15143 ( .A(n13100), .B(n13099), .Z(n13102) );
  AND U15144 ( .A(x[491]), .B(y[7793]), .Z(n13101) );
  XOR U15145 ( .A(n13102), .B(n13101), .Z(n13132) );
  AND U15146 ( .A(x[507]), .B(y[7777]), .Z(n13111) );
  XOR U15147 ( .A(o[124]), .B(n13111), .Z(n13120) );
  AND U15148 ( .A(x[506]), .B(y[7778]), .Z(n13119) );
  XOR U15149 ( .A(n13120), .B(n13119), .Z(n13122) );
  AND U15150 ( .A(x[495]), .B(y[7789]), .Z(n13121) );
  XNOR U15151 ( .A(n13122), .B(n13121), .Z(n13131) );
  XOR U15152 ( .A(n13133), .B(n13134), .Z(n13162) );
  NAND U15153 ( .A(n12917), .B(n12916), .Z(n12921) );
  NAND U15154 ( .A(n12919), .B(n12918), .Z(n12920) );
  NAND U15155 ( .A(n12921), .B(n12920), .Z(n13139) );
  AND U15156 ( .A(x[497]), .B(y[7787]), .Z(n13065) );
  AND U15157 ( .A(x[502]), .B(y[7782]), .Z(n13064) );
  XOR U15158 ( .A(n13065), .B(n13064), .Z(n13067) );
  AND U15159 ( .A(x[484]), .B(y[7800]), .Z(n13066) );
  XOR U15160 ( .A(n13067), .B(n13066), .Z(n13138) );
  AND U15161 ( .A(x[486]), .B(y[7798]), .Z(n13286) );
  AND U15162 ( .A(x[499]), .B(y[7785]), .Z(n13112) );
  XOR U15163 ( .A(n13286), .B(n13112), .Z(n13113) );
  XOR U15164 ( .A(n13114), .B(n13113), .Z(n13137) );
  XOR U15165 ( .A(n13138), .B(n13137), .Z(n13140) );
  XOR U15166 ( .A(n13139), .B(n13140), .Z(n13161) );
  NAND U15167 ( .A(n12922), .B(n13126), .Z(n12926) );
  NANDN U15168 ( .A(n12924), .B(n12923), .Z(n12925) );
  NAND U15169 ( .A(n12926), .B(n12925), .Z(n13060) );
  NAND U15170 ( .A(n12928), .B(n12927), .Z(n12932) );
  NAND U15171 ( .A(n12930), .B(n12929), .Z(n12931) );
  NAND U15172 ( .A(n12932), .B(n12931), .Z(n13059) );
  NAND U15173 ( .A(n12934), .B(n12933), .Z(n12938) );
  NAND U15174 ( .A(n12936), .B(n12935), .Z(n12937) );
  NAND U15175 ( .A(n12938), .B(n12937), .Z(n13058) );
  XOR U15176 ( .A(n13059), .B(n13058), .Z(n13061) );
  XOR U15177 ( .A(n13060), .B(n13061), .Z(n13163) );
  XOR U15178 ( .A(n13164), .B(n13163), .Z(n13054) );
  XNOR U15179 ( .A(n13055), .B(n13054), .Z(n13194) );
  NAND U15180 ( .A(n12940), .B(n12939), .Z(n12944) );
  NAND U15181 ( .A(n12942), .B(n12941), .Z(n12943) );
  NAND U15182 ( .A(n12944), .B(n12943), .Z(n13145) );
  NAND U15183 ( .A(n12946), .B(n12945), .Z(n12950) );
  NAND U15184 ( .A(n12948), .B(n12947), .Z(n12949) );
  NAND U15185 ( .A(n12950), .B(n12949), .Z(n13144) );
  NAND U15186 ( .A(n12952), .B(n12951), .Z(n12956) );
  NANDN U15187 ( .A(n12954), .B(n12953), .Z(n12955) );
  NAND U15188 ( .A(n12956), .B(n12955), .Z(n13143) );
  XOR U15189 ( .A(n13144), .B(n13143), .Z(n13146) );
  XOR U15190 ( .A(n13145), .B(n13146), .Z(n13192) );
  AND U15191 ( .A(x[500]), .B(y[7779]), .Z(n12957) );
  AND U15192 ( .A(x[504]), .B(y[7783]), .Z(n13522) );
  NAND U15193 ( .A(n12957), .B(n13522), .Z(n12961) );
  NAND U15194 ( .A(n12959), .B(n12958), .Z(n12960) );
  NAND U15195 ( .A(n12961), .B(n12960), .Z(n13181) );
  AND U15196 ( .A(x[505]), .B(y[7779]), .Z(n13095) );
  XOR U15197 ( .A(n13096), .B(n13095), .Z(n13094) );
  AND U15198 ( .A(x[481]), .B(y[7803]), .Z(n13093) );
  XOR U15199 ( .A(n13094), .B(n13093), .Z(n13180) );
  AND U15200 ( .A(x[496]), .B(y[7788]), .Z(n13088) );
  AND U15201 ( .A(x[504]), .B(y[7780]), .Z(n13087) );
  XOR U15202 ( .A(n13088), .B(n13087), .Z(n13090) );
  AND U15203 ( .A(x[482]), .B(y[7802]), .Z(n13089) );
  XOR U15204 ( .A(n13090), .B(n13089), .Z(n13179) );
  XOR U15205 ( .A(n13180), .B(n13179), .Z(n13182) );
  XOR U15206 ( .A(n13181), .B(n13182), .Z(n13152) );
  NAND U15207 ( .A(n12963), .B(n12962), .Z(n12967) );
  NAND U15208 ( .A(n12965), .B(n12964), .Z(n12966) );
  NAND U15209 ( .A(n12967), .B(n12966), .Z(n13175) );
  AND U15210 ( .A(x[483]), .B(y[7801]), .Z(n13125) );
  XOR U15211 ( .A(n13126), .B(n13125), .Z(n13128) );
  AND U15212 ( .A(x[503]), .B(y[7781]), .Z(n13127) );
  XOR U15213 ( .A(n13128), .B(n13127), .Z(n13174) );
  AND U15214 ( .A(x[485]), .B(y[7799]), .Z(n13106) );
  AND U15215 ( .A(x[501]), .B(y[7783]), .Z(n13105) );
  XOR U15216 ( .A(n13106), .B(n13105), .Z(n13108) );
  AND U15217 ( .A(x[500]), .B(y[7784]), .Z(n13107) );
  XOR U15218 ( .A(n13108), .B(n13107), .Z(n13173) );
  XOR U15219 ( .A(n13174), .B(n13173), .Z(n13176) );
  XOR U15220 ( .A(n13175), .B(n13176), .Z(n13150) );
  AND U15221 ( .A(n12968), .B(o[123]), .Z(n13073) );
  AND U15222 ( .A(x[480]), .B(y[7804]), .Z(n13071) );
  AND U15223 ( .A(x[508]), .B(y[7776]), .Z(n13070) );
  XOR U15224 ( .A(n13071), .B(n13070), .Z(n13072) );
  XOR U15225 ( .A(n13073), .B(n13072), .Z(n13082) );
  NAND U15226 ( .A(y[7794]), .B(x[490]), .Z(n12969) );
  XNOR U15227 ( .A(n12970), .B(n12969), .Z(n13078) );
  AND U15228 ( .A(x[489]), .B(y[7795]), .Z(n13077) );
  XOR U15229 ( .A(n13078), .B(n13077), .Z(n13081) );
  XOR U15230 ( .A(n13082), .B(n13081), .Z(n13084) );
  NAND U15231 ( .A(n12972), .B(n12971), .Z(n12976) );
  NAND U15232 ( .A(n12974), .B(n12973), .Z(n12975) );
  NAND U15233 ( .A(n12976), .B(n12975), .Z(n13083) );
  XOR U15234 ( .A(n13084), .B(n13083), .Z(n13170) );
  NAND U15235 ( .A(n12978), .B(n12977), .Z(n12982) );
  NAND U15236 ( .A(n12980), .B(n12979), .Z(n12981) );
  NAND U15237 ( .A(n12982), .B(n12981), .Z(n13168) );
  NAND U15238 ( .A(n12984), .B(n12983), .Z(n12988) );
  NAND U15239 ( .A(n12986), .B(n12985), .Z(n12987) );
  NAND U15240 ( .A(n12988), .B(n12987), .Z(n13167) );
  XOR U15241 ( .A(n13168), .B(n13167), .Z(n13169) );
  XNOR U15242 ( .A(n13170), .B(n13169), .Z(n13149) );
  XNOR U15243 ( .A(n13194), .B(n13193), .Z(n13187) );
  NAND U15244 ( .A(n12990), .B(n12989), .Z(n12994) );
  NANDN U15245 ( .A(n12992), .B(n12991), .Z(n12993) );
  NAND U15246 ( .A(n12994), .B(n12993), .Z(n13186) );
  NAND U15247 ( .A(n12996), .B(n12995), .Z(n13000) );
  NAND U15248 ( .A(n12998), .B(n12997), .Z(n12999) );
  NAND U15249 ( .A(n13000), .B(n12999), .Z(n13185) );
  XNOR U15250 ( .A(n13186), .B(n13185), .Z(n13188) );
  XNOR U15251 ( .A(n13040), .B(n13041), .Z(n13042) );
  NANDN U15252 ( .A(n13002), .B(n13001), .Z(n13006) );
  NAND U15253 ( .A(n13004), .B(n13003), .Z(n13005) );
  NAND U15254 ( .A(n13006), .B(n13005), .Z(n13048) );
  NANDN U15255 ( .A(n13008), .B(n13007), .Z(n13012) );
  NANDN U15256 ( .A(n13010), .B(n13009), .Z(n13011) );
  AND U15257 ( .A(n13012), .B(n13011), .Z(n13047) );
  NAND U15258 ( .A(n13014), .B(n13013), .Z(n13018) );
  NANDN U15259 ( .A(n13016), .B(n13015), .Z(n13017) );
  AND U15260 ( .A(n13018), .B(n13017), .Z(n13046) );
  XOR U15261 ( .A(n13047), .B(n13046), .Z(n13049) );
  XNOR U15262 ( .A(n13048), .B(n13049), .Z(n13043) );
  XNOR U15263 ( .A(n13036), .B(n13035), .Z(n13039) );
  NAND U15264 ( .A(n13020), .B(n13019), .Z(n13024) );
  NAND U15265 ( .A(n13022), .B(n13021), .Z(n13023) );
  AND U15266 ( .A(n13024), .B(n13023), .Z(n13037) );
  OR U15267 ( .A(n13027), .B(n13025), .Z(n13031) );
  ANDN U15268 ( .B(n13027), .A(n13026), .Z(n13029) );
  OR U15269 ( .A(n13029), .B(n13028), .Z(n13030) );
  AND U15270 ( .A(n13031), .B(n13030), .Z(n13038) );
  XNOR U15271 ( .A(n13037), .B(n13038), .Z(n13032) );
  XNOR U15272 ( .A(n13039), .B(n13032), .Z(N253) );
  NANDN U15273 ( .A(n13041), .B(n13040), .Z(n13045) );
  NANDN U15274 ( .A(n13043), .B(n13042), .Z(n13044) );
  NAND U15275 ( .A(n13045), .B(n13044), .Z(n13203) );
  NAND U15276 ( .A(n13047), .B(n13046), .Z(n13051) );
  NAND U15277 ( .A(n13049), .B(n13048), .Z(n13050) );
  NAND U15278 ( .A(n13051), .B(n13050), .Z(n13201) );
  NAND U15279 ( .A(n13053), .B(n13052), .Z(n13057) );
  NAND U15280 ( .A(n13055), .B(n13054), .Z(n13056) );
  NAND U15281 ( .A(n13057), .B(n13056), .Z(n13225) );
  NAND U15282 ( .A(n13059), .B(n13058), .Z(n13063) );
  NAND U15283 ( .A(n13061), .B(n13060), .Z(n13062) );
  AND U15284 ( .A(n13063), .B(n13062), .Z(n13330) );
  NAND U15285 ( .A(n13065), .B(n13064), .Z(n13069) );
  NAND U15286 ( .A(n13067), .B(n13066), .Z(n13068) );
  NAND U15287 ( .A(n13069), .B(n13068), .Z(n13353) );
  NAND U15288 ( .A(n13071), .B(n13070), .Z(n13075) );
  NAND U15289 ( .A(n13073), .B(n13072), .Z(n13074) );
  NAND U15290 ( .A(n13075), .B(n13074), .Z(n13352) );
  XOR U15291 ( .A(n13353), .B(n13352), .Z(n13354) );
  AND U15292 ( .A(y[7796]), .B(x[490]), .Z(n13366) );
  NAND U15293 ( .A(n13076), .B(n13366), .Z(n13080) );
  NAND U15294 ( .A(n13078), .B(n13077), .Z(n13079) );
  NAND U15295 ( .A(n13080), .B(n13079), .Z(n13342) );
  AND U15296 ( .A(x[502]), .B(y[7783]), .Z(n13275) );
  AND U15297 ( .A(x[492]), .B(y[7793]), .Z(n13485) );
  AND U15298 ( .A(x[481]), .B(y[7804]), .Z(n13273) );
  XOR U15299 ( .A(n13485), .B(n13273), .Z(n13274) );
  XOR U15300 ( .A(n13275), .B(n13274), .Z(n13341) );
  AND U15301 ( .A(x[495]), .B(y[7790]), .Z(n13278) );
  XOR U15302 ( .A(n13429), .B(n13278), .Z(n13279) );
  XOR U15303 ( .A(n13280), .B(n13279), .Z(n13340) );
  XOR U15304 ( .A(n13341), .B(n13340), .Z(n13343) );
  XNOR U15305 ( .A(n13342), .B(n13343), .Z(n13355) );
  NAND U15306 ( .A(n13082), .B(n13081), .Z(n13086) );
  NAND U15307 ( .A(n13084), .B(n13083), .Z(n13085) );
  AND U15308 ( .A(n13086), .B(n13085), .Z(n13328) );
  XNOR U15309 ( .A(n13330), .B(n13331), .Z(n13325) );
  NAND U15310 ( .A(n13088), .B(n13087), .Z(n13092) );
  NAND U15311 ( .A(n13090), .B(n13089), .Z(n13091) );
  NAND U15312 ( .A(n13092), .B(n13091), .Z(n13347) );
  AND U15313 ( .A(n13094), .B(n13093), .Z(n13098) );
  NAND U15314 ( .A(n13096), .B(n13095), .Z(n13097) );
  NANDN U15315 ( .A(n13098), .B(n13097), .Z(n13346) );
  XOR U15316 ( .A(n13347), .B(n13346), .Z(n13348) );
  NAND U15317 ( .A(n13100), .B(n13099), .Z(n13104) );
  NAND U15318 ( .A(n13102), .B(n13101), .Z(n13103) );
  NAND U15319 ( .A(n13104), .B(n13103), .Z(n13239) );
  AND U15320 ( .A(x[491]), .B(y[7794]), .Z(n13296) );
  AND U15321 ( .A(x[483]), .B(y[7802]), .Z(n13294) );
  AND U15322 ( .A(x[497]), .B(y[7788]), .Z(n13293) );
  XOR U15323 ( .A(n13294), .B(n13293), .Z(n13295) );
  XOR U15324 ( .A(n13296), .B(n13295), .Z(n13238) );
  AND U15325 ( .A(x[503]), .B(y[7782]), .Z(n13301) );
  AND U15326 ( .A(x[493]), .B(y[7792]), .Z(n13299) );
  AND U15327 ( .A(x[504]), .B(y[7781]), .Z(n13456) );
  XOR U15328 ( .A(n13299), .B(n13456), .Z(n13300) );
  XOR U15329 ( .A(n13301), .B(n13300), .Z(n13237) );
  XOR U15330 ( .A(n13238), .B(n13237), .Z(n13240) );
  XNOR U15331 ( .A(n13239), .B(n13240), .Z(n13349) );
  NAND U15332 ( .A(n13106), .B(n13105), .Z(n13110) );
  NAND U15333 ( .A(n13108), .B(n13107), .Z(n13109) );
  NAND U15334 ( .A(n13110), .B(n13109), .Z(n13306) );
  AND U15335 ( .A(n13111), .B(o[124]), .Z(n13246) );
  AND U15336 ( .A(x[496]), .B(y[7789]), .Z(n13244) );
  AND U15337 ( .A(x[507]), .B(y[7778]), .Z(n13243) );
  XOR U15338 ( .A(n13244), .B(n13243), .Z(n13245) );
  XOR U15339 ( .A(n13246), .B(n13245), .Z(n13305) );
  AND U15340 ( .A(x[482]), .B(y[7803]), .Z(n13255) );
  XOR U15341 ( .A(n13256), .B(n13255), .Z(n13257) );
  XOR U15342 ( .A(n13258), .B(n13257), .Z(n13304) );
  XOR U15343 ( .A(n13305), .B(n13304), .Z(n13307) );
  XOR U15344 ( .A(n13306), .B(n13307), .Z(n13311) );
  NAND U15345 ( .A(n13286), .B(n13112), .Z(n13116) );
  NAND U15346 ( .A(n13114), .B(n13113), .Z(n13115) );
  AND U15347 ( .A(n13116), .B(n13115), .Z(n13336) );
  AND U15348 ( .A(x[505]), .B(y[7780]), .Z(n13270) );
  AND U15349 ( .A(x[506]), .B(y[7779]), .Z(n13267) );
  XOR U15350 ( .A(n13268), .B(n13267), .Z(n13269) );
  XOR U15351 ( .A(n13270), .B(n13269), .Z(n13335) );
  AND U15352 ( .A(x[508]), .B(y[7777]), .Z(n13285) );
  XOR U15353 ( .A(o[125]), .B(n13285), .Z(n13361) );
  AND U15354 ( .A(x[480]), .B(y[7805]), .Z(n13359) );
  AND U15355 ( .A(x[509]), .B(y[7776]), .Z(n13358) );
  XOR U15356 ( .A(n13359), .B(n13358), .Z(n13360) );
  XNOR U15357 ( .A(n13361), .B(n13360), .Z(n13334) );
  XNOR U15358 ( .A(n13336), .B(n13337), .Z(n13310) );
  AND U15359 ( .A(y[7799]), .B(x[486]), .Z(n13118) );
  NAND U15360 ( .A(y[7798]), .B(x[487]), .Z(n13117) );
  XNOR U15361 ( .A(n13118), .B(n13117), .Z(n13288) );
  AND U15362 ( .A(x[488]), .B(y[7797]), .Z(n13287) );
  XOR U15363 ( .A(n13288), .B(n13287), .Z(n13368) );
  AND U15364 ( .A(x[489]), .B(y[7796]), .Z(n13518) );
  XOR U15365 ( .A(n13368), .B(n13518), .Z(n13370) );
  AND U15366 ( .A(x[484]), .B(y[7801]), .Z(n13250) );
  AND U15367 ( .A(x[490]), .B(y[7795]), .Z(n13249) );
  XOR U15368 ( .A(n13250), .B(n13249), .Z(n13252) );
  AND U15369 ( .A(x[485]), .B(y[7800]), .Z(n13251) );
  XOR U15370 ( .A(n13252), .B(n13251), .Z(n13369) );
  XOR U15371 ( .A(n13370), .B(n13369), .Z(n13263) );
  NAND U15372 ( .A(n13120), .B(n13119), .Z(n13124) );
  NAND U15373 ( .A(n13122), .B(n13121), .Z(n13123) );
  NAND U15374 ( .A(n13124), .B(n13123), .Z(n13262) );
  NAND U15375 ( .A(n13126), .B(n13125), .Z(n13130) );
  NAND U15376 ( .A(n13128), .B(n13127), .Z(n13129) );
  NAND U15377 ( .A(n13130), .B(n13129), .Z(n13261) );
  XNOR U15378 ( .A(n13262), .B(n13261), .Z(n13264) );
  NANDN U15379 ( .A(n13132), .B(n13131), .Z(n13136) );
  NAND U15380 ( .A(n13134), .B(n13133), .Z(n13135) );
  NAND U15381 ( .A(n13136), .B(n13135), .Z(n13231) );
  XNOR U15382 ( .A(n13233), .B(n13234), .Z(n13323) );
  NAND U15383 ( .A(n13138), .B(n13137), .Z(n13142) );
  NAND U15384 ( .A(n13140), .B(n13139), .Z(n13141) );
  NAND U15385 ( .A(n13142), .B(n13141), .Z(n13322) );
  XOR U15386 ( .A(n13225), .B(n13226), .Z(n13228) );
  NAND U15387 ( .A(n13144), .B(n13143), .Z(n13148) );
  NAND U15388 ( .A(n13146), .B(n13145), .Z(n13147) );
  NAND U15389 ( .A(n13148), .B(n13147), .Z(n13219) );
  NANDN U15390 ( .A(n13150), .B(n13149), .Z(n13154) );
  NANDN U15391 ( .A(n13152), .B(n13151), .Z(n13153) );
  AND U15392 ( .A(n13154), .B(n13153), .Z(n13220) );
  XOR U15393 ( .A(n13219), .B(n13220), .Z(n13222) );
  NAND U15394 ( .A(n13156), .B(n13155), .Z(n13160) );
  NAND U15395 ( .A(n13158), .B(n13157), .Z(n13159) );
  NAND U15396 ( .A(n13160), .B(n13159), .Z(n13215) );
  NANDN U15397 ( .A(n13162), .B(n13161), .Z(n13166) );
  NAND U15398 ( .A(n13164), .B(n13163), .Z(n13165) );
  NAND U15399 ( .A(n13166), .B(n13165), .Z(n13213) );
  NAND U15400 ( .A(n13168), .B(n13167), .Z(n13172) );
  NAND U15401 ( .A(n13170), .B(n13169), .Z(n13171) );
  NAND U15402 ( .A(n13172), .B(n13171), .Z(n13318) );
  NAND U15403 ( .A(n13174), .B(n13173), .Z(n13178) );
  NAND U15404 ( .A(n13176), .B(n13175), .Z(n13177) );
  NAND U15405 ( .A(n13178), .B(n13177), .Z(n13317) );
  NAND U15406 ( .A(n13180), .B(n13179), .Z(n13184) );
  NAND U15407 ( .A(n13182), .B(n13181), .Z(n13183) );
  NAND U15408 ( .A(n13184), .B(n13183), .Z(n13316) );
  XOR U15409 ( .A(n13317), .B(n13316), .Z(n13319) );
  XOR U15410 ( .A(n13318), .B(n13319), .Z(n13214) );
  XOR U15411 ( .A(n13213), .B(n13214), .Z(n13216) );
  XOR U15412 ( .A(n13215), .B(n13216), .Z(n13221) );
  XOR U15413 ( .A(n13222), .B(n13221), .Z(n13227) );
  XOR U15414 ( .A(n13228), .B(n13227), .Z(n13209) );
  NAND U15415 ( .A(n13186), .B(n13185), .Z(n13190) );
  NANDN U15416 ( .A(n13188), .B(n13187), .Z(n13189) );
  NAND U15417 ( .A(n13190), .B(n13189), .Z(n13207) );
  NANDN U15418 ( .A(n13192), .B(n13191), .Z(n13196) );
  NAND U15419 ( .A(n13194), .B(n13193), .Z(n13195) );
  AND U15420 ( .A(n13196), .B(n13195), .Z(n13208) );
  XNOR U15421 ( .A(n13207), .B(n13208), .Z(n13210) );
  XOR U15422 ( .A(n13201), .B(n13202), .Z(n13204) );
  XOR U15423 ( .A(n13203), .B(n13204), .Z(n13200) );
  XOR U15424 ( .A(n13198), .B(n13200), .Z(n13197) );
  XOR U15425 ( .A(n13199), .B(n13197), .Z(N254) );
  NAND U15426 ( .A(n13202), .B(n13201), .Z(n13206) );
  NAND U15427 ( .A(n13204), .B(n13203), .Z(n13205) );
  AND U15428 ( .A(n13206), .B(n13205), .Z(n13375) );
  XNOR U15429 ( .A(n13376), .B(n13375), .Z(n13374) );
  NAND U15430 ( .A(n13208), .B(n13207), .Z(n13212) );
  NANDN U15431 ( .A(n13210), .B(n13209), .Z(n13211) );
  NAND U15432 ( .A(n13212), .B(n13211), .Z(n13657) );
  NAND U15433 ( .A(n13214), .B(n13213), .Z(n13218) );
  NAND U15434 ( .A(n13216), .B(n13215), .Z(n13217) );
  AND U15435 ( .A(n13218), .B(n13217), .Z(n13664) );
  NAND U15436 ( .A(n13220), .B(n13219), .Z(n13224) );
  NAND U15437 ( .A(n13222), .B(n13221), .Z(n13223) );
  AND U15438 ( .A(n13224), .B(n13223), .Z(n13666) );
  NAND U15439 ( .A(n13226), .B(n13225), .Z(n13230) );
  NAND U15440 ( .A(n13228), .B(n13227), .Z(n13229) );
  AND U15441 ( .A(n13230), .B(n13229), .Z(n13665) );
  XOR U15442 ( .A(n13666), .B(n13665), .Z(n13663) );
  XNOR U15443 ( .A(n13664), .B(n13663), .Z(n13659) );
  NANDN U15444 ( .A(n13232), .B(n13231), .Z(n13236) );
  NANDN U15445 ( .A(n13234), .B(n13233), .Z(n13235) );
  AND U15446 ( .A(n13236), .B(n13235), .Z(n13645) );
  NAND U15447 ( .A(n13238), .B(n13237), .Z(n13242) );
  NAND U15448 ( .A(n13240), .B(n13239), .Z(n13241) );
  AND U15449 ( .A(n13242), .B(n13241), .Z(n13629) );
  NAND U15450 ( .A(n13244), .B(n13243), .Z(n13248) );
  NAND U15451 ( .A(n13246), .B(n13245), .Z(n13247) );
  NAND U15452 ( .A(n13248), .B(n13247), .Z(n13587) );
  NAND U15453 ( .A(n13250), .B(n13249), .Z(n13254) );
  NAND U15454 ( .A(n13252), .B(n13251), .Z(n13253) );
  NAND U15455 ( .A(n13254), .B(n13253), .Z(n13590) );
  AND U15456 ( .A(x[486]), .B(y[7800]), .Z(n13437) );
  AND U15457 ( .A(x[485]), .B(y[7801]), .Z(n13435) );
  AND U15458 ( .A(x[499]), .B(y[7787]), .Z(n13434) );
  XOR U15459 ( .A(n13435), .B(n13434), .Z(n13436) );
  XNOR U15460 ( .A(n13437), .B(n13436), .Z(n13417) );
  AND U15461 ( .A(x[484]), .B(y[7802]), .Z(n13480) );
  AND U15462 ( .A(x[483]), .B(y[7803]), .Z(n13482) );
  AND U15463 ( .A(x[498]), .B(y[7788]), .Z(n13481) );
  XOR U15464 ( .A(n13482), .B(n13481), .Z(n13479) );
  XOR U15465 ( .A(n13480), .B(n13479), .Z(n13420) );
  NAND U15466 ( .A(n13256), .B(n13255), .Z(n13260) );
  NAND U15467 ( .A(n13258), .B(n13257), .Z(n13259) );
  AND U15468 ( .A(n13260), .B(n13259), .Z(n13419) );
  XOR U15469 ( .A(n13417), .B(n13418), .Z(n13589) );
  XOR U15470 ( .A(n13590), .B(n13589), .Z(n13588) );
  XOR U15471 ( .A(n13587), .B(n13588), .Z(n13630) );
  NAND U15472 ( .A(n13262), .B(n13261), .Z(n13266) );
  NANDN U15473 ( .A(n13264), .B(n13263), .Z(n13265) );
  AND U15474 ( .A(n13266), .B(n13265), .Z(n13627) );
  XOR U15475 ( .A(n13628), .B(n13627), .Z(n13648) );
  AND U15476 ( .A(n13268), .B(n13267), .Z(n13272) );
  NAND U15477 ( .A(n13270), .B(n13269), .Z(n13271) );
  NANDN U15478 ( .A(n13272), .B(n13271), .Z(n13581) );
  AND U15479 ( .A(n13485), .B(n13273), .Z(n13277) );
  NAND U15480 ( .A(n13275), .B(n13274), .Z(n13276) );
  NANDN U15481 ( .A(n13277), .B(n13276), .Z(n13584) );
  NAND U15482 ( .A(n13429), .B(n13278), .Z(n13282) );
  NAND U15483 ( .A(n13280), .B(n13279), .Z(n13281) );
  AND U15484 ( .A(n13282), .B(n13281), .Z(n13398) );
  AND U15485 ( .A(x[503]), .B(y[7783]), .Z(n13455) );
  AND U15486 ( .A(x[504]), .B(y[7782]), .Z(n13284) );
  AND U15487 ( .A(y[7781]), .B(x[505]), .Z(n13283) );
  XOR U15488 ( .A(n13284), .B(n13283), .Z(n13454) );
  XOR U15489 ( .A(n13455), .B(n13454), .Z(n13400) );
  AND U15490 ( .A(n13285), .B(o[125]), .Z(n13443) );
  AND U15491 ( .A(x[508]), .B(y[7778]), .Z(n13445) );
  AND U15492 ( .A(x[496]), .B(y[7790]), .Z(n13444) );
  XOR U15493 ( .A(n13445), .B(n13444), .Z(n13442) );
  XNOR U15494 ( .A(n13443), .B(n13442), .Z(n13399) );
  XNOR U15495 ( .A(n13398), .B(n13397), .Z(n13583) );
  XOR U15496 ( .A(n13584), .B(n13583), .Z(n13582) );
  XOR U15497 ( .A(n13581), .B(n13582), .Z(n13622) );
  AND U15498 ( .A(x[487]), .B(y[7799]), .Z(n13431) );
  NAND U15499 ( .A(n13286), .B(n13431), .Z(n13290) );
  NAND U15500 ( .A(n13288), .B(n13287), .Z(n13289) );
  AND U15501 ( .A(n13290), .B(n13289), .Z(n13409) );
  AND U15502 ( .A(y[7785]), .B(x[501]), .Z(n13292) );
  AND U15503 ( .A(y[7784]), .B(x[502]), .Z(n13291) );
  XOR U15504 ( .A(n13292), .B(n13291), .Z(n13430) );
  XOR U15505 ( .A(n13431), .B(n13430), .Z(n13412) );
  AND U15506 ( .A(x[497]), .B(y[7789]), .Z(n13509) );
  AND U15507 ( .A(x[482]), .B(y[7804]), .Z(n13511) );
  AND U15508 ( .A(x[506]), .B(y[7780]), .Z(n13510) );
  XOR U15509 ( .A(n13511), .B(n13510), .Z(n13508) );
  XNOR U15510 ( .A(n13509), .B(n13508), .Z(n13411) );
  XNOR U15511 ( .A(n13409), .B(n13410), .Z(n13610) );
  NAND U15512 ( .A(n13294), .B(n13293), .Z(n13298) );
  NAND U15513 ( .A(n13296), .B(n13295), .Z(n13297) );
  AND U15514 ( .A(n13298), .B(n13297), .Z(n13423) );
  AND U15515 ( .A(x[480]), .B(y[7806]), .Z(n13497) );
  AND U15516 ( .A(x[509]), .B(y[7777]), .Z(n13521) );
  XOR U15517 ( .A(o[126]), .B(n13521), .Z(n13499) );
  AND U15518 ( .A(x[510]), .B(y[7776]), .Z(n13498) );
  XOR U15519 ( .A(n13499), .B(n13498), .Z(n13496) );
  XOR U15520 ( .A(n13497), .B(n13496), .Z(n13426) );
  AND U15521 ( .A(x[500]), .B(y[7786]), .Z(n13504) );
  XOR U15522 ( .A(n13505), .B(n13504), .Z(n13503) );
  AND U15523 ( .A(x[488]), .B(y[7798]), .Z(n13502) );
  XNOR U15524 ( .A(n13503), .B(n13502), .Z(n13425) );
  XNOR U15525 ( .A(n13423), .B(n13424), .Z(n13612) );
  NAND U15526 ( .A(n13299), .B(n13456), .Z(n13303) );
  NAND U15527 ( .A(n13301), .B(n13300), .Z(n13302) );
  NAND U15528 ( .A(n13303), .B(n13302), .Z(n13611) );
  NAND U15529 ( .A(n13305), .B(n13304), .Z(n13309) );
  NAND U15530 ( .A(n13307), .B(n13306), .Z(n13308) );
  NAND U15531 ( .A(n13309), .B(n13308), .Z(n13623) );
  XOR U15532 ( .A(n13624), .B(n13623), .Z(n13621) );
  XOR U15533 ( .A(n13622), .B(n13621), .Z(n13647) );
  XOR U15534 ( .A(n13645), .B(n13646), .Z(n13640) );
  NANDN U15535 ( .A(n13311), .B(n13310), .Z(n13315) );
  NANDN U15536 ( .A(n13313), .B(n13312), .Z(n13314) );
  NAND U15537 ( .A(n13315), .B(n13314), .Z(n13641) );
  NAND U15538 ( .A(n13317), .B(n13316), .Z(n13321) );
  NAND U15539 ( .A(n13319), .B(n13318), .Z(n13320) );
  AND U15540 ( .A(n13321), .B(n13320), .Z(n13642) );
  XOR U15541 ( .A(n13641), .B(n13642), .Z(n13639) );
  XNOR U15542 ( .A(n13640), .B(n13639), .Z(n13379) );
  NANDN U15543 ( .A(n13323), .B(n13322), .Z(n13327) );
  NANDN U15544 ( .A(n13325), .B(n13324), .Z(n13326) );
  NAND U15545 ( .A(n13327), .B(n13326), .Z(n13381) );
  NANDN U15546 ( .A(n13329), .B(n13328), .Z(n13333) );
  NANDN U15547 ( .A(n13331), .B(n13330), .Z(n13332) );
  AND U15548 ( .A(n13333), .B(n13332), .Z(n13386) );
  NANDN U15549 ( .A(n13335), .B(n13334), .Z(n13339) );
  NANDN U15550 ( .A(n13337), .B(n13336), .Z(n13338) );
  NAND U15551 ( .A(n13339), .B(n13338), .Z(n13603) );
  NAND U15552 ( .A(n13341), .B(n13340), .Z(n13345) );
  NAND U15553 ( .A(n13343), .B(n13342), .Z(n13344) );
  AND U15554 ( .A(n13345), .B(n13344), .Z(n13606) );
  NAND U15555 ( .A(n13347), .B(n13346), .Z(n13351) );
  NANDN U15556 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U15557 ( .A(n13351), .B(n13350), .Z(n13605) );
  XOR U15558 ( .A(n13606), .B(n13605), .Z(n13604) );
  XOR U15559 ( .A(n13603), .B(n13604), .Z(n13388) );
  NAND U15560 ( .A(n13353), .B(n13352), .Z(n13357) );
  NANDN U15561 ( .A(n13355), .B(n13354), .Z(n13356) );
  AND U15562 ( .A(n13357), .B(n13356), .Z(n13392) );
  NAND U15563 ( .A(n13359), .B(n13358), .Z(n13363) );
  NAND U15564 ( .A(n13361), .B(n13360), .Z(n13362) );
  NAND U15565 ( .A(n13363), .B(n13362), .Z(n13403) );
  AND U15566 ( .A(y[7794]), .B(x[492]), .Z(n13364) );
  XOR U15567 ( .A(n13365), .B(n13364), .Z(n13486) );
  XOR U15568 ( .A(n13487), .B(n13486), .Z(n13517) );
  AND U15569 ( .A(y[7797]), .B(x[489]), .Z(n13367) );
  XOR U15570 ( .A(n13367), .B(n13366), .Z(n13516) );
  XOR U15571 ( .A(n13517), .B(n13516), .Z(n13406) );
  AND U15572 ( .A(x[507]), .B(y[7779]), .Z(n13451) );
  AND U15573 ( .A(x[481]), .B(y[7805]), .Z(n13450) );
  XOR U15574 ( .A(n13451), .B(n13450), .Z(n13448) );
  XOR U15575 ( .A(n13449), .B(n13448), .Z(n13405) );
  XOR U15576 ( .A(n13406), .B(n13405), .Z(n13404) );
  XOR U15577 ( .A(n13403), .B(n13404), .Z(n13394) );
  NAND U15578 ( .A(n13368), .B(n13518), .Z(n13372) );
  NAND U15579 ( .A(n13370), .B(n13369), .Z(n13371) );
  AND U15580 ( .A(n13372), .B(n13371), .Z(n13393) );
  XNOR U15581 ( .A(n13392), .B(n13391), .Z(n13387) );
  XOR U15582 ( .A(n13386), .B(n13385), .Z(n13382) );
  XNOR U15583 ( .A(n13381), .B(n13382), .Z(n13380) );
  XOR U15584 ( .A(n13659), .B(n13660), .Z(n13658) );
  XOR U15585 ( .A(n13657), .B(n13658), .Z(n13373) );
  XNOR U15586 ( .A(n13374), .B(n13373), .Z(N255) );
  NAND U15587 ( .A(n13374), .B(n13373), .Z(n13378) );
  NANDN U15588 ( .A(n13376), .B(n13375), .Z(n13377) );
  AND U15589 ( .A(n13378), .B(n13377), .Z(n13674) );
  NANDN U15590 ( .A(n13380), .B(n13379), .Z(n13384) );
  NAND U15591 ( .A(n13382), .B(n13381), .Z(n13383) );
  AND U15592 ( .A(n13384), .B(n13383), .Z(n13656) );
  NAND U15593 ( .A(n13386), .B(n13385), .Z(n13390) );
  NANDN U15594 ( .A(n13388), .B(n13387), .Z(n13389) );
  AND U15595 ( .A(n13390), .B(n13389), .Z(n13638) );
  NAND U15596 ( .A(n13392), .B(n13391), .Z(n13396) );
  NANDN U15597 ( .A(n13394), .B(n13393), .Z(n13395) );
  AND U15598 ( .A(n13396), .B(n13395), .Z(n13620) );
  NAND U15599 ( .A(n13398), .B(n13397), .Z(n13402) );
  NANDN U15600 ( .A(n13400), .B(n13399), .Z(n13401) );
  AND U15601 ( .A(n13402), .B(n13401), .Z(n13602) );
  NAND U15602 ( .A(n13404), .B(n13403), .Z(n13408) );
  NAND U15603 ( .A(n13406), .B(n13405), .Z(n13407) );
  AND U15604 ( .A(n13408), .B(n13407), .Z(n13416) );
  NANDN U15605 ( .A(n13410), .B(n13409), .Z(n13414) );
  NANDN U15606 ( .A(n13412), .B(n13411), .Z(n13413) );
  NAND U15607 ( .A(n13414), .B(n13413), .Z(n13415) );
  XNOR U15608 ( .A(n13416), .B(n13415), .Z(n13600) );
  NANDN U15609 ( .A(n13418), .B(n13417), .Z(n13422) );
  NANDN U15610 ( .A(n13420), .B(n13419), .Z(n13421) );
  AND U15611 ( .A(n13422), .B(n13421), .Z(n13598) );
  NANDN U15612 ( .A(n13424), .B(n13423), .Z(n13428) );
  NANDN U15613 ( .A(n13426), .B(n13425), .Z(n13427) );
  AND U15614 ( .A(n13428), .B(n13427), .Z(n13580) );
  AND U15615 ( .A(x[502]), .B(y[7785]), .Z(n13541) );
  AND U15616 ( .A(n13429), .B(n13541), .Z(n13433) );
  AND U15617 ( .A(n13431), .B(n13430), .Z(n13432) );
  NOR U15618 ( .A(n13433), .B(n13432), .Z(n13441) );
  NAND U15619 ( .A(n13435), .B(n13434), .Z(n13439) );
  NAND U15620 ( .A(n13437), .B(n13436), .Z(n13438) );
  AND U15621 ( .A(n13439), .B(n13438), .Z(n13440) );
  XNOR U15622 ( .A(n13441), .B(n13440), .Z(n13495) );
  NAND U15623 ( .A(n13443), .B(n13442), .Z(n13447) );
  NAND U15624 ( .A(n13445), .B(n13444), .Z(n13446) );
  AND U15625 ( .A(n13447), .B(n13446), .Z(n13478) );
  NAND U15626 ( .A(n13449), .B(n13448), .Z(n13453) );
  NAND U15627 ( .A(n13451), .B(n13450), .Z(n13452) );
  AND U15628 ( .A(n13453), .B(n13452), .Z(n13460) );
  NAND U15629 ( .A(n13455), .B(n13454), .Z(n13458) );
  AND U15630 ( .A(x[505]), .B(y[7782]), .Z(n13542) );
  NAND U15631 ( .A(n13456), .B(n13542), .Z(n13457) );
  NAND U15632 ( .A(n13458), .B(n13457), .Z(n13459) );
  XNOR U15633 ( .A(n13460), .B(n13459), .Z(n13476) );
  AND U15634 ( .A(y[7784]), .B(x[503]), .Z(n13462) );
  NAND U15635 ( .A(y[7805]), .B(x[482]), .Z(n13461) );
  XNOR U15636 ( .A(n13462), .B(n13461), .Z(n13466) );
  AND U15637 ( .A(y[7801]), .B(x[486]), .Z(n13464) );
  NAND U15638 ( .A(y[7804]), .B(x[483]), .Z(n13463) );
  XNOR U15639 ( .A(n13464), .B(n13463), .Z(n13465) );
  XOR U15640 ( .A(n13466), .B(n13465), .Z(n13474) );
  AND U15641 ( .A(y[7800]), .B(x[487]), .Z(n13468) );
  NAND U15642 ( .A(y[7790]), .B(x[497]), .Z(n13467) );
  XNOR U15643 ( .A(n13468), .B(n13467), .Z(n13472) );
  AND U15644 ( .A(y[7802]), .B(x[485]), .Z(n13470) );
  NAND U15645 ( .A(y[7803]), .B(x[484]), .Z(n13469) );
  XNOR U15646 ( .A(n13470), .B(n13469), .Z(n13471) );
  XNOR U15647 ( .A(n13472), .B(n13471), .Z(n13473) );
  XNOR U15648 ( .A(n13474), .B(n13473), .Z(n13475) );
  XNOR U15649 ( .A(n13476), .B(n13475), .Z(n13477) );
  XNOR U15650 ( .A(n13478), .B(n13477), .Z(n13493) );
  NAND U15651 ( .A(n13480), .B(n13479), .Z(n13484) );
  NAND U15652 ( .A(n13482), .B(n13481), .Z(n13483) );
  AND U15653 ( .A(n13484), .B(n13483), .Z(n13491) );
  NAND U15654 ( .A(n13527), .B(n13485), .Z(n13489) );
  NAND U15655 ( .A(n13487), .B(n13486), .Z(n13488) );
  AND U15656 ( .A(n13489), .B(n13488), .Z(n13490) );
  XNOR U15657 ( .A(n13491), .B(n13490), .Z(n13492) );
  XNOR U15658 ( .A(n13493), .B(n13492), .Z(n13494) );
  XNOR U15659 ( .A(n13495), .B(n13494), .Z(n13578) );
  NAND U15660 ( .A(n13497), .B(n13496), .Z(n13501) );
  NAND U15661 ( .A(n13499), .B(n13498), .Z(n13500) );
  AND U15662 ( .A(n13501), .B(n13500), .Z(n13576) );
  NAND U15663 ( .A(n13503), .B(n13502), .Z(n13507) );
  NAND U15664 ( .A(n13505), .B(n13504), .Z(n13506) );
  AND U15665 ( .A(n13507), .B(n13506), .Z(n13515) );
  NAND U15666 ( .A(n13509), .B(n13508), .Z(n13513) );
  NAND U15667 ( .A(n13511), .B(n13510), .Z(n13512) );
  NAND U15668 ( .A(n13513), .B(n13512), .Z(n13514) );
  XNOR U15669 ( .A(n13515), .B(n13514), .Z(n13574) );
  NAND U15670 ( .A(n13517), .B(n13516), .Z(n13520) );
  AND U15671 ( .A(x[490]), .B(y[7797]), .Z(n13536) );
  NAND U15672 ( .A(n13518), .B(n13536), .Z(n13519) );
  AND U15673 ( .A(n13520), .B(n13519), .Z(n13572) );
  AND U15674 ( .A(n13521), .B(o[126]), .Z(n13526) );
  AND U15675 ( .A(y[7788]), .B(x[499]), .Z(n13524) );
  XNOR U15676 ( .A(n13522), .B(o[127]), .Z(n13523) );
  XNOR U15677 ( .A(n13524), .B(n13523), .Z(n13525) );
  XOR U15678 ( .A(n13526), .B(n13525), .Z(n13530) );
  XNOR U15679 ( .A(n13528), .B(n13527), .Z(n13529) );
  XNOR U15680 ( .A(n13530), .B(n13529), .Z(n13570) );
  AND U15681 ( .A(y[7795]), .B(x[492]), .Z(n13532) );
  NAND U15682 ( .A(y[7781]), .B(x[506]), .Z(n13531) );
  XNOR U15683 ( .A(n13532), .B(n13531), .Z(n13540) );
  AND U15684 ( .A(y[7796]), .B(x[491]), .Z(n13538) );
  AND U15685 ( .A(y[7806]), .B(x[481]), .Z(n13534) );
  NAND U15686 ( .A(y[7779]), .B(x[508]), .Z(n13533) );
  XNOR U15687 ( .A(n13534), .B(n13533), .Z(n13535) );
  XNOR U15688 ( .A(n13536), .B(n13535), .Z(n13537) );
  XNOR U15689 ( .A(n13538), .B(n13537), .Z(n13539) );
  XOR U15690 ( .A(n13540), .B(n13539), .Z(n13544) );
  XNOR U15691 ( .A(n13542), .B(n13541), .Z(n13543) );
  XNOR U15692 ( .A(n13544), .B(n13543), .Z(n13560) );
  AND U15693 ( .A(y[7777]), .B(x[510]), .Z(n13546) );
  NAND U15694 ( .A(y[7791]), .B(x[496]), .Z(n13545) );
  XNOR U15695 ( .A(n13546), .B(n13545), .Z(n13550) );
  AND U15696 ( .A(y[7789]), .B(x[498]), .Z(n13548) );
  NAND U15697 ( .A(y[7787]), .B(x[500]), .Z(n13547) );
  XNOR U15698 ( .A(n13548), .B(n13547), .Z(n13549) );
  XOR U15699 ( .A(n13550), .B(n13549), .Z(n13558) );
  AND U15700 ( .A(y[7798]), .B(x[489]), .Z(n13552) );
  NAND U15701 ( .A(y[7807]), .B(x[480]), .Z(n13551) );
  XNOR U15702 ( .A(n13552), .B(n13551), .Z(n13556) );
  AND U15703 ( .A(y[7778]), .B(x[509]), .Z(n13554) );
  NAND U15704 ( .A(y[7793]), .B(x[494]), .Z(n13553) );
  XNOR U15705 ( .A(n13554), .B(n13553), .Z(n13555) );
  XNOR U15706 ( .A(n13556), .B(n13555), .Z(n13557) );
  XNOR U15707 ( .A(n13558), .B(n13557), .Z(n13559) );
  XOR U15708 ( .A(n13560), .B(n13559), .Z(n13568) );
  AND U15709 ( .A(y[7786]), .B(x[501]), .Z(n13562) );
  NAND U15710 ( .A(y[7799]), .B(x[488]), .Z(n13561) );
  XNOR U15711 ( .A(n13562), .B(n13561), .Z(n13566) );
  AND U15712 ( .A(y[7776]), .B(x[511]), .Z(n13564) );
  NAND U15713 ( .A(y[7780]), .B(x[507]), .Z(n13563) );
  XNOR U15714 ( .A(n13564), .B(n13563), .Z(n13565) );
  XNOR U15715 ( .A(n13566), .B(n13565), .Z(n13567) );
  XNOR U15716 ( .A(n13568), .B(n13567), .Z(n13569) );
  XNOR U15717 ( .A(n13570), .B(n13569), .Z(n13571) );
  XNOR U15718 ( .A(n13572), .B(n13571), .Z(n13573) );
  XNOR U15719 ( .A(n13574), .B(n13573), .Z(n13575) );
  XNOR U15720 ( .A(n13576), .B(n13575), .Z(n13577) );
  XNOR U15721 ( .A(n13578), .B(n13577), .Z(n13579) );
  XNOR U15722 ( .A(n13580), .B(n13579), .Z(n13596) );
  NAND U15723 ( .A(n13582), .B(n13581), .Z(n13586) );
  NAND U15724 ( .A(n13584), .B(n13583), .Z(n13585) );
  AND U15725 ( .A(n13586), .B(n13585), .Z(n13594) );
  NAND U15726 ( .A(n13588), .B(n13587), .Z(n13592) );
  NAND U15727 ( .A(n13590), .B(n13589), .Z(n13591) );
  NAND U15728 ( .A(n13592), .B(n13591), .Z(n13593) );
  XNOR U15729 ( .A(n13594), .B(n13593), .Z(n13595) );
  XNOR U15730 ( .A(n13596), .B(n13595), .Z(n13597) );
  XNOR U15731 ( .A(n13598), .B(n13597), .Z(n13599) );
  XNOR U15732 ( .A(n13600), .B(n13599), .Z(n13601) );
  XNOR U15733 ( .A(n13602), .B(n13601), .Z(n13618) );
  NAND U15734 ( .A(n13604), .B(n13603), .Z(n13608) );
  NAND U15735 ( .A(n13606), .B(n13605), .Z(n13607) );
  AND U15736 ( .A(n13608), .B(n13607), .Z(n13616) );
  NANDN U15737 ( .A(n13610), .B(n13609), .Z(n13614) );
  NANDN U15738 ( .A(n13612), .B(n13611), .Z(n13613) );
  NAND U15739 ( .A(n13614), .B(n13613), .Z(n13615) );
  XNOR U15740 ( .A(n13616), .B(n13615), .Z(n13617) );
  XNOR U15741 ( .A(n13618), .B(n13617), .Z(n13619) );
  XNOR U15742 ( .A(n13620), .B(n13619), .Z(n13636) );
  NAND U15743 ( .A(n13622), .B(n13621), .Z(n13626) );
  NAND U15744 ( .A(n13624), .B(n13623), .Z(n13625) );
  AND U15745 ( .A(n13626), .B(n13625), .Z(n13634) );
  NAND U15746 ( .A(n13628), .B(n13627), .Z(n13632) );
  NANDN U15747 ( .A(n13630), .B(n13629), .Z(n13631) );
  NAND U15748 ( .A(n13632), .B(n13631), .Z(n13633) );
  XNOR U15749 ( .A(n13634), .B(n13633), .Z(n13635) );
  XNOR U15750 ( .A(n13636), .B(n13635), .Z(n13637) );
  XNOR U15751 ( .A(n13638), .B(n13637), .Z(n13654) );
  NAND U15752 ( .A(n13640), .B(n13639), .Z(n13644) );
  NAND U15753 ( .A(n13642), .B(n13641), .Z(n13643) );
  AND U15754 ( .A(n13644), .B(n13643), .Z(n13652) );
  NANDN U15755 ( .A(n13646), .B(n13645), .Z(n13650) );
  NANDN U15756 ( .A(n13648), .B(n13647), .Z(n13649) );
  NAND U15757 ( .A(n13650), .B(n13649), .Z(n13651) );
  XNOR U15758 ( .A(n13652), .B(n13651), .Z(n13653) );
  XNOR U15759 ( .A(n13654), .B(n13653), .Z(n13655) );
  XNOR U15760 ( .A(n13656), .B(n13655), .Z(n13672) );
  NANDN U15761 ( .A(n13658), .B(n13657), .Z(n13662) );
  NANDN U15762 ( .A(n13660), .B(n13659), .Z(n13661) );
  AND U15763 ( .A(n13662), .B(n13661), .Z(n13670) );
  NAND U15764 ( .A(n13664), .B(n13663), .Z(n13668) );
  NAND U15765 ( .A(n13666), .B(n13665), .Z(n13667) );
  NAND U15766 ( .A(n13668), .B(n13667), .Z(n13669) );
  XNOR U15767 ( .A(n13670), .B(n13669), .Z(n13671) );
  XNOR U15768 ( .A(n13672), .B(n13671), .Z(n13673) );
  XNOR U15769 ( .A(n13674), .B(n13673), .Z(N256) );
  AND U15770 ( .A(x[480]), .B(y[7808]), .Z(n14320) );
  XOR U15771 ( .A(n14320), .B(o[128]), .Z(N289) );
  NAND U15772 ( .A(x[481]), .B(y[7808]), .Z(n13684) );
  AND U15773 ( .A(x[480]), .B(y[7809]), .Z(n13680) );
  XNOR U15774 ( .A(n13680), .B(o[129]), .Z(n13675) );
  XOR U15775 ( .A(n13684), .B(n13675), .Z(n13677) );
  NAND U15776 ( .A(n14320), .B(o[128]), .Z(n13676) );
  XNOR U15777 ( .A(n13677), .B(n13676), .Z(N290) );
  AND U15778 ( .A(x[480]), .B(y[7810]), .Z(n13683) );
  XNOR U15779 ( .A(n13683), .B(o[130]), .Z(n13689) );
  XNOR U15780 ( .A(n13690), .B(n13689), .Z(n13692) );
  AND U15781 ( .A(y[7808]), .B(x[482]), .Z(n13679) );
  NAND U15782 ( .A(y[7809]), .B(x[481]), .Z(n13678) );
  XNOR U15783 ( .A(n13679), .B(n13678), .Z(n13686) );
  AND U15784 ( .A(n13680), .B(o[129]), .Z(n13685) );
  XNOR U15785 ( .A(n13686), .B(n13685), .Z(n13691) );
  XNOR U15786 ( .A(n13692), .B(n13691), .Z(N291) );
  AND U15787 ( .A(x[481]), .B(y[7810]), .Z(n13803) );
  AND U15788 ( .A(x[482]), .B(y[7809]), .Z(n13700) );
  XOR U15789 ( .A(n13700), .B(o[131]), .Z(n13704) );
  XOR U15790 ( .A(n13803), .B(n13704), .Z(n13706) );
  AND U15791 ( .A(y[7808]), .B(x[483]), .Z(n13682) );
  NAND U15792 ( .A(y[7811]), .B(x[480]), .Z(n13681) );
  XNOR U15793 ( .A(n13682), .B(n13681), .Z(n13697) );
  AND U15794 ( .A(n13683), .B(o[130]), .Z(n13696) );
  XOR U15795 ( .A(n13697), .B(n13696), .Z(n13705) );
  XNOR U15796 ( .A(n13706), .B(n13705), .Z(n13711) );
  NANDN U15797 ( .A(n13684), .B(n13700), .Z(n13688) );
  NAND U15798 ( .A(n13686), .B(n13685), .Z(n13687) );
  NAND U15799 ( .A(n13688), .B(n13687), .Z(n13709) );
  NANDN U15800 ( .A(n13690), .B(n13689), .Z(n13694) );
  NAND U15801 ( .A(n13692), .B(n13691), .Z(n13693) );
  AND U15802 ( .A(n13694), .B(n13693), .Z(n13710) );
  XOR U15803 ( .A(n13709), .B(n13710), .Z(n13695) );
  XNOR U15804 ( .A(n13711), .B(n13695), .Z(N292) );
  AND U15805 ( .A(x[483]), .B(y[7811]), .Z(n13760) );
  NAND U15806 ( .A(n14320), .B(n13760), .Z(n13699) );
  NAND U15807 ( .A(n13697), .B(n13696), .Z(n13698) );
  NAND U15808 ( .A(n13699), .B(n13698), .Z(n13732) );
  AND U15809 ( .A(n13700), .B(o[131]), .Z(n13724) );
  AND U15810 ( .A(y[7812]), .B(x[480]), .Z(n13702) );
  AND U15811 ( .A(y[7808]), .B(x[484]), .Z(n13701) );
  XOR U15812 ( .A(n13702), .B(n13701), .Z(n13723) );
  XOR U15813 ( .A(n13724), .B(n13723), .Z(n13731) );
  AND U15814 ( .A(y[7810]), .B(x[482]), .Z(n13851) );
  NAND U15815 ( .A(y[7811]), .B(x[481]), .Z(n13703) );
  XNOR U15816 ( .A(n13851), .B(n13703), .Z(n13720) );
  AND U15817 ( .A(x[483]), .B(y[7809]), .Z(n13715) );
  XOR U15818 ( .A(o[132]), .B(n13715), .Z(n13719) );
  XOR U15819 ( .A(n13720), .B(n13719), .Z(n13730) );
  XOR U15820 ( .A(n13731), .B(n13730), .Z(n13733) );
  XOR U15821 ( .A(n13732), .B(n13733), .Z(n13729) );
  NAND U15822 ( .A(n13803), .B(n13704), .Z(n13708) );
  NAND U15823 ( .A(n13706), .B(n13705), .Z(n13707) );
  AND U15824 ( .A(n13708), .B(n13707), .Z(n13728) );
  XNOR U15825 ( .A(n13728), .B(n13727), .Z(n13712) );
  XNOR U15826 ( .A(n13729), .B(n13712), .Z(N293) );
  AND U15827 ( .A(y[7808]), .B(x[485]), .Z(n13714) );
  NAND U15828 ( .A(y[7813]), .B(x[480]), .Z(n13713) );
  XNOR U15829 ( .A(n13714), .B(n13713), .Z(n13753) );
  AND U15830 ( .A(o[132]), .B(n13715), .Z(n13752) );
  XOR U15831 ( .A(n13753), .B(n13752), .Z(n13751) );
  NAND U15832 ( .A(x[482]), .B(y[7811]), .Z(n13811) );
  AND U15833 ( .A(y[7810]), .B(x[483]), .Z(n13717) );
  NAND U15834 ( .A(y[7812]), .B(x[481]), .Z(n13716) );
  XNOR U15835 ( .A(n13717), .B(n13716), .Z(n13747) );
  AND U15836 ( .A(x[484]), .B(y[7809]), .Z(n13758) );
  XOR U15837 ( .A(n13758), .B(o[133]), .Z(n13746) );
  XOR U15838 ( .A(n13747), .B(n13746), .Z(n13750) );
  XOR U15839 ( .A(n13811), .B(n13750), .Z(n13718) );
  XNOR U15840 ( .A(n13751), .B(n13718), .Z(n13739) );
  NANDN U15841 ( .A(n13811), .B(n13803), .Z(n13722) );
  NAND U15842 ( .A(n13720), .B(n13719), .Z(n13721) );
  NAND U15843 ( .A(n13722), .B(n13721), .Z(n13738) );
  AND U15844 ( .A(x[484]), .B(y[7812]), .Z(n14502) );
  NAND U15845 ( .A(n14502), .B(n14320), .Z(n13726) );
  NAND U15846 ( .A(n13724), .B(n13723), .Z(n13725) );
  NAND U15847 ( .A(n13726), .B(n13725), .Z(n13737) );
  XNOR U15848 ( .A(n13738), .B(n13737), .Z(n13740) );
  NAND U15849 ( .A(n13731), .B(n13730), .Z(n13735) );
  NAND U15850 ( .A(n13733), .B(n13732), .Z(n13734) );
  AND U15851 ( .A(n13735), .B(n13734), .Z(n13743) );
  XOR U15852 ( .A(n13744), .B(n13743), .Z(n13736) );
  XNOR U15853 ( .A(n13745), .B(n13736), .Z(N294) );
  NAND U15854 ( .A(n13738), .B(n13737), .Z(n13742) );
  NANDN U15855 ( .A(n13740), .B(n13739), .Z(n13741) );
  AND U15856 ( .A(n13742), .B(n13741), .Z(n13793) );
  AND U15857 ( .A(x[483]), .B(y[7812]), .Z(n13812) );
  NAND U15858 ( .A(n13812), .B(n13803), .Z(n13749) );
  NAND U15859 ( .A(n13747), .B(n13746), .Z(n13748) );
  NAND U15860 ( .A(n13749), .B(n13748), .Z(n13788) );
  XOR U15861 ( .A(n13788), .B(n13787), .Z(n13790) );
  AND U15862 ( .A(x[485]), .B(y[7813]), .Z(n13983) );
  NAND U15863 ( .A(n14320), .B(n13983), .Z(n13755) );
  NAND U15864 ( .A(n13753), .B(n13752), .Z(n13754) );
  NAND U15865 ( .A(n13755), .B(n13754), .Z(n13763) );
  AND U15866 ( .A(y[7808]), .B(x[486]), .Z(n13757) );
  NAND U15867 ( .A(y[7814]), .B(x[480]), .Z(n13756) );
  XNOR U15868 ( .A(n13757), .B(n13756), .Z(n13770) );
  AND U15869 ( .A(n13758), .B(o[133]), .Z(n13771) );
  XOR U15870 ( .A(n13770), .B(n13771), .Z(n13764) );
  XOR U15871 ( .A(n13763), .B(n13764), .Z(n13766) );
  NAND U15872 ( .A(y[7812]), .B(x[482]), .Z(n13759) );
  XNOR U15873 ( .A(n13760), .B(n13759), .Z(n13775) );
  AND U15874 ( .A(y[7813]), .B(x[481]), .Z(n14016) );
  NAND U15875 ( .A(y[7810]), .B(x[484]), .Z(n13761) );
  XNOR U15876 ( .A(n14016), .B(n13761), .Z(n13779) );
  AND U15877 ( .A(x[485]), .B(y[7809]), .Z(n13786) );
  XOR U15878 ( .A(n13786), .B(o[134]), .Z(n13778) );
  XOR U15879 ( .A(n13779), .B(n13778), .Z(n13774) );
  XOR U15880 ( .A(n13775), .B(n13774), .Z(n13765) );
  XOR U15881 ( .A(n13766), .B(n13765), .Z(n13789) );
  XOR U15882 ( .A(n13790), .B(n13789), .Z(n13795) );
  XNOR U15883 ( .A(n13794), .B(n13795), .Z(n13762) );
  XOR U15884 ( .A(n13793), .B(n13762), .Z(N295) );
  NAND U15885 ( .A(n13764), .B(n13763), .Z(n13768) );
  NAND U15886 ( .A(n13766), .B(n13765), .Z(n13767) );
  AND U15887 ( .A(n13768), .B(n13767), .Z(n13834) );
  AND U15888 ( .A(y[7810]), .B(x[485]), .Z(n13905) );
  NAND U15889 ( .A(y[7814]), .B(x[481]), .Z(n13769) );
  XNOR U15890 ( .A(n13905), .B(n13769), .Z(n13805) );
  NAND U15891 ( .A(x[486]), .B(y[7809]), .Z(n13808) );
  XNOR U15892 ( .A(o[135]), .B(n13808), .Z(n13804) );
  XNOR U15893 ( .A(n13805), .B(n13804), .Z(n13823) );
  AND U15894 ( .A(x[486]), .B(y[7814]), .Z(n14036) );
  NAND U15895 ( .A(n14320), .B(n14036), .Z(n13773) );
  NAND U15896 ( .A(n13771), .B(n13770), .Z(n13772) );
  AND U15897 ( .A(n13773), .B(n13772), .Z(n13822) );
  XOR U15898 ( .A(n13823), .B(n13822), .Z(n13824) );
  NANDN U15899 ( .A(n13811), .B(n13812), .Z(n13777) );
  NAND U15900 ( .A(n13775), .B(n13774), .Z(n13776) );
  AND U15901 ( .A(n13777), .B(n13776), .Z(n13825) );
  XOR U15902 ( .A(n13824), .B(n13825), .Z(n13832) );
  AND U15903 ( .A(x[484]), .B(y[7813]), .Z(n14325) );
  NAND U15904 ( .A(n14325), .B(n13803), .Z(n13781) );
  NAND U15905 ( .A(n13779), .B(n13778), .Z(n13780) );
  AND U15906 ( .A(n13781), .B(n13780), .Z(n13800) );
  AND U15907 ( .A(y[7813]), .B(x[482]), .Z(n13783) );
  NAND U15908 ( .A(y[7811]), .B(x[484]), .Z(n13782) );
  XNOR U15909 ( .A(n13783), .B(n13782), .Z(n13813) );
  XNOR U15910 ( .A(n13813), .B(n13812), .Z(n13798) );
  AND U15911 ( .A(y[7808]), .B(x[487]), .Z(n13785) );
  NAND U15912 ( .A(y[7815]), .B(x[480]), .Z(n13784) );
  XNOR U15913 ( .A(n13785), .B(n13784), .Z(n13817) );
  AND U15914 ( .A(n13786), .B(o[134]), .Z(n13816) );
  XNOR U15915 ( .A(n13817), .B(n13816), .Z(n13797) );
  XOR U15916 ( .A(n13798), .B(n13797), .Z(n13799) );
  XOR U15917 ( .A(n13800), .B(n13799), .Z(n13831) );
  XOR U15918 ( .A(n13832), .B(n13831), .Z(n13833) );
  XOR U15919 ( .A(n13834), .B(n13833), .Z(n13830) );
  NAND U15920 ( .A(n13788), .B(n13787), .Z(n13792) );
  NAND U15921 ( .A(n13790), .B(n13789), .Z(n13791) );
  NAND U15922 ( .A(n13792), .B(n13791), .Z(n13829) );
  XOR U15923 ( .A(n13829), .B(n13828), .Z(n13796) );
  XNOR U15924 ( .A(n13830), .B(n13796), .Z(N296) );
  NAND U15925 ( .A(n13798), .B(n13797), .Z(n13802) );
  NAND U15926 ( .A(n13800), .B(n13799), .Z(n13801) );
  AND U15927 ( .A(n13802), .B(n13801), .Z(n13884) );
  AND U15928 ( .A(x[485]), .B(y[7814]), .Z(n13975) );
  NAND U15929 ( .A(n13975), .B(n13803), .Z(n13807) );
  NAND U15930 ( .A(n13805), .B(n13804), .Z(n13806) );
  NAND U15931 ( .A(n13807), .B(n13806), .Z(n13882) );
  ANDN U15932 ( .B(o[135]), .A(n13808), .Z(n13871) );
  AND U15933 ( .A(y[7811]), .B(x[485]), .Z(n14408) );
  NAND U15934 ( .A(y[7815]), .B(x[481]), .Z(n13809) );
  XOR U15935 ( .A(n14408), .B(n13809), .Z(n13872) );
  XOR U15936 ( .A(n13871), .B(n13872), .Z(n13856) );
  NAND U15937 ( .A(x[483]), .B(y[7813]), .Z(n14638) );
  AND U15938 ( .A(x[486]), .B(y[7810]), .Z(n13810) );
  AND U15939 ( .A(y[7814]), .B(x[482]), .Z(n14725) );
  XOR U15940 ( .A(n13810), .B(n14725), .Z(n13852) );
  XOR U15941 ( .A(n14502), .B(n13852), .Z(n13855) );
  XOR U15942 ( .A(n14638), .B(n13855), .Z(n13857) );
  XOR U15943 ( .A(n13856), .B(n13857), .Z(n13881) );
  XOR U15944 ( .A(n13882), .B(n13881), .Z(n13883) );
  XNOR U15945 ( .A(n13884), .B(n13883), .Z(n13841) );
  NANDN U15946 ( .A(n13811), .B(n14325), .Z(n13815) );
  NAND U15947 ( .A(n13813), .B(n13812), .Z(n13814) );
  NAND U15948 ( .A(n13815), .B(n13814), .Z(n13877) );
  AND U15949 ( .A(x[487]), .B(y[7815]), .Z(n14193) );
  NAND U15950 ( .A(n14320), .B(n14193), .Z(n13819) );
  NAND U15951 ( .A(n13817), .B(n13816), .Z(n13818) );
  NAND U15952 ( .A(n13819), .B(n13818), .Z(n13875) );
  AND U15953 ( .A(y[7808]), .B(x[488]), .Z(n13821) );
  NAND U15954 ( .A(y[7816]), .B(x[480]), .Z(n13820) );
  XNOR U15955 ( .A(n13821), .B(n13820), .Z(n13862) );
  NAND U15956 ( .A(x[487]), .B(y[7809]), .Z(n13865) );
  XNOR U15957 ( .A(o[136]), .B(n13865), .Z(n13861) );
  XOR U15958 ( .A(n13862), .B(n13861), .Z(n13876) );
  XOR U15959 ( .A(n13875), .B(n13876), .Z(n13878) );
  XNOR U15960 ( .A(n13877), .B(n13878), .Z(n13839) );
  NAND U15961 ( .A(n13823), .B(n13822), .Z(n13827) );
  NAND U15962 ( .A(n13825), .B(n13824), .Z(n13826) );
  NAND U15963 ( .A(n13827), .B(n13826), .Z(n13838) );
  XOR U15964 ( .A(n13839), .B(n13838), .Z(n13840) );
  XOR U15965 ( .A(n13841), .B(n13840), .Z(n13847) );
  NAND U15966 ( .A(n13832), .B(n13831), .Z(n13836) );
  NAND U15967 ( .A(n13834), .B(n13833), .Z(n13835) );
  AND U15968 ( .A(n13836), .B(n13835), .Z(n13845) );
  IV U15969 ( .A(n13845), .Z(n13844) );
  XOR U15970 ( .A(n13846), .B(n13844), .Z(n13837) );
  XNOR U15971 ( .A(n13847), .B(n13837), .Z(N297) );
  NAND U15972 ( .A(n13839), .B(n13838), .Z(n13843) );
  NAND U15973 ( .A(n13841), .B(n13840), .Z(n13842) );
  NAND U15974 ( .A(n13843), .B(n13842), .Z(n13896) );
  IV U15975 ( .A(n13896), .Z(n13894) );
  OR U15976 ( .A(n13846), .B(n13844), .Z(n13850) );
  ANDN U15977 ( .B(n13846), .A(n13845), .Z(n13848) );
  OR U15978 ( .A(n13848), .B(n13847), .Z(n13849) );
  AND U15979 ( .A(n13850), .B(n13849), .Z(n13895) );
  NAND U15980 ( .A(n14036), .B(n13851), .Z(n13854) );
  NAND U15981 ( .A(n14502), .B(n13852), .Z(n13853) );
  NAND U15982 ( .A(n13854), .B(n13853), .Z(n13901) );
  NANDN U15983 ( .A(n13855), .B(n14638), .Z(n13859) );
  NANDN U15984 ( .A(n13857), .B(n13856), .Z(n13858) );
  AND U15985 ( .A(n13859), .B(n13858), .Z(n13902) );
  XOR U15986 ( .A(n13901), .B(n13902), .Z(n13903) );
  AND U15987 ( .A(x[488]), .B(y[7816]), .Z(n13860) );
  NAND U15988 ( .A(n13860), .B(n14320), .Z(n13864) );
  NAND U15989 ( .A(n13862), .B(n13861), .Z(n13863) );
  AND U15990 ( .A(n13864), .B(n13863), .Z(n13934) );
  ANDN U15991 ( .B(o[136]), .A(n13865), .Z(n13907) );
  AND U15992 ( .A(y[7812]), .B(x[485]), .Z(n13867) );
  NAND U15993 ( .A(y[7810]), .B(x[487]), .Z(n13866) );
  XNOR U15994 ( .A(n13867), .B(n13866), .Z(n13906) );
  XNOR U15995 ( .A(n13907), .B(n13906), .Z(n13932) );
  AND U15996 ( .A(y[7808]), .B(x[489]), .Z(n13869) );
  NAND U15997 ( .A(y[7817]), .B(x[480]), .Z(n13868) );
  XNOR U15998 ( .A(n13869), .B(n13868), .Z(n13914) );
  AND U15999 ( .A(x[488]), .B(y[7809]), .Z(n13923) );
  XOR U16000 ( .A(o[137]), .B(n13923), .Z(n13913) );
  XNOR U16001 ( .A(n13914), .B(n13913), .Z(n13931) );
  XOR U16002 ( .A(n13932), .B(n13931), .Z(n13933) );
  XOR U16003 ( .A(n13934), .B(n13933), .Z(n13928) );
  AND U16004 ( .A(y[7811]), .B(x[486]), .Z(n14274) );
  NAND U16005 ( .A(y[7816]), .B(x[481]), .Z(n13870) );
  XNOR U16006 ( .A(n14274), .B(n13870), .Z(n13918) );
  XNOR U16007 ( .A(n14325), .B(n13918), .Z(n13938) );
  AND U16008 ( .A(x[482]), .B(y[7815]), .Z(n14549) );
  NAND U16009 ( .A(x[483]), .B(y[7814]), .Z(n14280) );
  XNOR U16010 ( .A(n14549), .B(n14280), .Z(n13937) );
  XNOR U16011 ( .A(n13938), .B(n13937), .Z(n13926) );
  NAND U16012 ( .A(x[485]), .B(y[7815]), .Z(n14112) );
  AND U16013 ( .A(x[481]), .B(y[7811]), .Z(n13917) );
  NANDN U16014 ( .A(n14112), .B(n13917), .Z(n13874) );
  NANDN U16015 ( .A(n13872), .B(n13871), .Z(n13873) );
  NAND U16016 ( .A(n13874), .B(n13873), .Z(n13925) );
  XOR U16017 ( .A(n13926), .B(n13925), .Z(n13927) );
  XOR U16018 ( .A(n13928), .B(n13927), .Z(n13904) );
  XNOR U16019 ( .A(n13903), .B(n13904), .Z(n13890) );
  NAND U16020 ( .A(n13876), .B(n13875), .Z(n13880) );
  NAND U16021 ( .A(n13878), .B(n13877), .Z(n13879) );
  NAND U16022 ( .A(n13880), .B(n13879), .Z(n13889) );
  NAND U16023 ( .A(n13882), .B(n13881), .Z(n13886) );
  NAND U16024 ( .A(n13884), .B(n13883), .Z(n13885) );
  NAND U16025 ( .A(n13886), .B(n13885), .Z(n13888) );
  XOR U16026 ( .A(n13889), .B(n13888), .Z(n13891) );
  XOR U16027 ( .A(n13890), .B(n13891), .Z(n13897) );
  XNOR U16028 ( .A(n13895), .B(n13897), .Z(n13887) );
  XOR U16029 ( .A(n13894), .B(n13887), .Z(N298) );
  NAND U16030 ( .A(n13889), .B(n13888), .Z(n13893) );
  NAND U16031 ( .A(n13891), .B(n13890), .Z(n13892) );
  AND U16032 ( .A(n13893), .B(n13892), .Z(n13994) );
  NANDN U16033 ( .A(n13894), .B(n13895), .Z(n13900) );
  NOR U16034 ( .A(n13896), .B(n13895), .Z(n13898) );
  OR U16035 ( .A(n13898), .B(n13897), .Z(n13899) );
  AND U16036 ( .A(n13900), .B(n13899), .Z(n13993) );
  XNOR U16037 ( .A(n13994), .B(n13993), .Z(n13996) );
  AND U16038 ( .A(x[487]), .B(y[7812]), .Z(n13977) );
  NAND U16039 ( .A(n13977), .B(n13905), .Z(n13909) );
  NAND U16040 ( .A(n13907), .B(n13906), .Z(n13908) );
  AND U16041 ( .A(n13909), .B(n13908), .Z(n13990) );
  AND U16042 ( .A(y[7811]), .B(x[487]), .Z(n13911) );
  NAND U16043 ( .A(y[7814]), .B(x[484]), .Z(n13910) );
  XNOR U16044 ( .A(n13911), .B(n13910), .Z(n13961) );
  AND U16045 ( .A(x[486]), .B(y[7812]), .Z(n13960) );
  XNOR U16046 ( .A(n13961), .B(n13960), .Z(n13988) );
  AND U16047 ( .A(x[488]), .B(y[7810]), .Z(n14169) );
  AND U16048 ( .A(x[489]), .B(y[7809]), .Z(n13971) );
  XOR U16049 ( .A(o[138]), .B(n13971), .Z(n13982) );
  XOR U16050 ( .A(n14169), .B(n13982), .Z(n13984) );
  XNOR U16051 ( .A(n13984), .B(n13983), .Z(n13987) );
  XOR U16052 ( .A(n13988), .B(n13987), .Z(n13989) );
  XNOR U16053 ( .A(n13990), .B(n13989), .Z(n13950) );
  AND U16054 ( .A(x[489]), .B(y[7817]), .Z(n13912) );
  NAND U16055 ( .A(n13912), .B(n14320), .Z(n13916) );
  NAND U16056 ( .A(n13914), .B(n13913), .Z(n13915) );
  NAND U16057 ( .A(n13916), .B(n13915), .Z(n13948) );
  AND U16058 ( .A(x[486]), .B(y[7816]), .Z(n14203) );
  NAND U16059 ( .A(n14203), .B(n13917), .Z(n13920) );
  NAND U16060 ( .A(n14325), .B(n13918), .Z(n13919) );
  NAND U16061 ( .A(n13920), .B(n13919), .Z(n13956) );
  AND U16062 ( .A(y[7808]), .B(x[490]), .Z(n13922) );
  NAND U16063 ( .A(y[7818]), .B(x[480]), .Z(n13921) );
  XNOR U16064 ( .A(n13922), .B(n13921), .Z(n13966) );
  AND U16065 ( .A(o[137]), .B(n13923), .Z(n13965) );
  XOR U16066 ( .A(n13966), .B(n13965), .Z(n13954) );
  AND U16067 ( .A(y[7815]), .B(x[483]), .Z(n14867) );
  NAND U16068 ( .A(y[7817]), .B(x[481]), .Z(n13924) );
  XNOR U16069 ( .A(n14867), .B(n13924), .Z(n13978) );
  AND U16070 ( .A(x[482]), .B(y[7816]), .Z(n13979) );
  XOR U16071 ( .A(n13978), .B(n13979), .Z(n13953) );
  XOR U16072 ( .A(n13954), .B(n13953), .Z(n13955) );
  XOR U16073 ( .A(n13956), .B(n13955), .Z(n13947) );
  XOR U16074 ( .A(n13948), .B(n13947), .Z(n13949) );
  XOR U16075 ( .A(n13950), .B(n13949), .Z(n14000) );
  NAND U16076 ( .A(n13926), .B(n13925), .Z(n13930) );
  NANDN U16077 ( .A(n13928), .B(n13927), .Z(n13929) );
  AND U16078 ( .A(n13930), .B(n13929), .Z(n13944) );
  NAND U16079 ( .A(n13932), .B(n13931), .Z(n13936) );
  NAND U16080 ( .A(n13934), .B(n13933), .Z(n13935) );
  AND U16081 ( .A(n13936), .B(n13935), .Z(n13941) );
  NAND U16082 ( .A(n13938), .B(n13937), .Z(n13940) );
  ANDN U16083 ( .B(n14280), .A(n14549), .Z(n13939) );
  ANDN U16084 ( .B(n13940), .A(n13939), .Z(n13942) );
  XOR U16085 ( .A(n13941), .B(n13942), .Z(n13943) );
  XOR U16086 ( .A(n13944), .B(n13943), .Z(n13999) );
  XNOR U16087 ( .A(n14000), .B(n13999), .Z(n14001) );
  XNOR U16088 ( .A(n14002), .B(n14001), .Z(n13995) );
  XOR U16089 ( .A(n13996), .B(n13995), .Z(N299) );
  NAND U16090 ( .A(n13942), .B(n13941), .Z(n13946) );
  NANDN U16091 ( .A(n13944), .B(n13943), .Z(n13945) );
  AND U16092 ( .A(n13946), .B(n13945), .Z(n14067) );
  NAND U16093 ( .A(n13948), .B(n13947), .Z(n13952) );
  NAND U16094 ( .A(n13950), .B(n13949), .Z(n13951) );
  NAND U16095 ( .A(n13952), .B(n13951), .Z(n14065) );
  NAND U16096 ( .A(n13954), .B(n13953), .Z(n13958) );
  NAND U16097 ( .A(n13956), .B(n13955), .Z(n13957) );
  NAND U16098 ( .A(n13958), .B(n13957), .Z(n14058) );
  AND U16099 ( .A(x[487]), .B(y[7814]), .Z(n14107) );
  AND U16100 ( .A(x[484]), .B(y[7811]), .Z(n13959) );
  NAND U16101 ( .A(n14107), .B(n13959), .Z(n13963) );
  NAND U16102 ( .A(n13961), .B(n13960), .Z(n13962) );
  NAND U16103 ( .A(n13963), .B(n13962), .Z(n14056) );
  AND U16104 ( .A(x[490]), .B(y[7818]), .Z(n13964) );
  NAND U16105 ( .A(n13964), .B(n14320), .Z(n13968) );
  NAND U16106 ( .A(n13966), .B(n13965), .Z(n13967) );
  NAND U16107 ( .A(n13968), .B(n13967), .Z(n14052) );
  AND U16108 ( .A(y[7808]), .B(x[491]), .Z(n13970) );
  NAND U16109 ( .A(y[7819]), .B(x[480]), .Z(n13969) );
  XNOR U16110 ( .A(n13970), .B(n13969), .Z(n14027) );
  AND U16111 ( .A(o[138]), .B(n13971), .Z(n14026) );
  XOR U16112 ( .A(n14027), .B(n14026), .Z(n14050) );
  AND U16113 ( .A(y[7813]), .B(x[486]), .Z(n13973) );
  NAND U16114 ( .A(y[7818]), .B(x[481]), .Z(n13972) );
  XNOR U16115 ( .A(n13973), .B(n13972), .Z(n14018) );
  AND U16116 ( .A(x[490]), .B(y[7809]), .Z(n14037) );
  XOR U16117 ( .A(o[139]), .B(n14037), .Z(n14017) );
  XOR U16118 ( .A(n14018), .B(n14017), .Z(n14049) );
  XOR U16119 ( .A(n14050), .B(n14049), .Z(n14051) );
  XOR U16120 ( .A(n14052), .B(n14051), .Z(n14055) );
  XOR U16121 ( .A(n14056), .B(n14055), .Z(n14057) );
  XNOR U16122 ( .A(n14058), .B(n14057), .Z(n14040) );
  AND U16123 ( .A(x[483]), .B(y[7816]), .Z(n15006) );
  NAND U16124 ( .A(y[7817]), .B(x[482]), .Z(n13974) );
  XNOR U16125 ( .A(n13975), .B(n13974), .Z(n14013) );
  AND U16126 ( .A(x[484]), .B(y[7815]), .Z(n14012) );
  XNOR U16127 ( .A(n14013), .B(n14012), .Z(n14044) );
  XNOR U16128 ( .A(n15006), .B(n14044), .Z(n14046) );
  NAND U16129 ( .A(y[7810]), .B(x[489]), .Z(n13976) );
  XNOR U16130 ( .A(n13977), .B(n13976), .Z(n14032) );
  AND U16131 ( .A(x[488]), .B(y[7811]), .Z(n14031) );
  XNOR U16132 ( .A(n14032), .B(n14031), .Z(n14045) );
  XNOR U16133 ( .A(n14046), .B(n14045), .Z(n14009) );
  NAND U16134 ( .A(x[483]), .B(y[7817]), .Z(n14103) );
  AND U16135 ( .A(x[481]), .B(y[7815]), .Z(n14315) );
  NANDN U16136 ( .A(n14103), .B(n14315), .Z(n13981) );
  NAND U16137 ( .A(n13979), .B(n13978), .Z(n13980) );
  NAND U16138 ( .A(n13981), .B(n13980), .Z(n14007) );
  NAND U16139 ( .A(n14169), .B(n13982), .Z(n13986) );
  NAND U16140 ( .A(n13984), .B(n13983), .Z(n13985) );
  NAND U16141 ( .A(n13986), .B(n13985), .Z(n14006) );
  XOR U16142 ( .A(n14007), .B(n14006), .Z(n14008) );
  XNOR U16143 ( .A(n14009), .B(n14008), .Z(n14039) );
  NAND U16144 ( .A(n13988), .B(n13987), .Z(n13992) );
  NAND U16145 ( .A(n13990), .B(n13989), .Z(n13991) );
  NAND U16146 ( .A(n13992), .B(n13991), .Z(n14038) );
  XOR U16147 ( .A(n14039), .B(n14038), .Z(n14041) );
  XNOR U16148 ( .A(n14040), .B(n14041), .Z(n14064) );
  XOR U16149 ( .A(n14065), .B(n14064), .Z(n14066) );
  XOR U16150 ( .A(n14067), .B(n14066), .Z(n14063) );
  NANDN U16151 ( .A(n13994), .B(n13993), .Z(n13998) );
  NAND U16152 ( .A(n13996), .B(n13995), .Z(n13997) );
  NAND U16153 ( .A(n13998), .B(n13997), .Z(n14061) );
  NANDN U16154 ( .A(n14000), .B(n13999), .Z(n14004) );
  NAND U16155 ( .A(n14002), .B(n14001), .Z(n14003) );
  AND U16156 ( .A(n14004), .B(n14003), .Z(n14062) );
  XOR U16157 ( .A(n14061), .B(n14062), .Z(n14005) );
  XNOR U16158 ( .A(n14063), .B(n14005), .Z(N300) );
  NAND U16159 ( .A(n14007), .B(n14006), .Z(n14011) );
  NAND U16160 ( .A(n14009), .B(n14008), .Z(n14010) );
  NAND U16161 ( .A(n14011), .B(n14010), .Z(n14144) );
  AND U16162 ( .A(x[485]), .B(y[7817]), .Z(n14540) );
  NAND U16163 ( .A(n14725), .B(n14540), .Z(n14015) );
  NAND U16164 ( .A(n14013), .B(n14012), .Z(n14014) );
  NAND U16165 ( .A(n14015), .B(n14014), .Z(n14091) );
  AND U16166 ( .A(x[486]), .B(y[7818]), .Z(n14332) );
  NAND U16167 ( .A(n14332), .B(n14016), .Z(n14020) );
  NAND U16168 ( .A(n14018), .B(n14017), .Z(n14019) );
  NAND U16169 ( .A(n14020), .B(n14019), .Z(n14090) );
  XOR U16170 ( .A(n14091), .B(n14090), .Z(n14092) );
  AND U16171 ( .A(x[489]), .B(y[7811]), .Z(n14720) );
  AND U16172 ( .A(x[490]), .B(y[7810]), .Z(n14774) );
  AND U16173 ( .A(y[7816]), .B(x[484]), .Z(n14021) );
  XOR U16174 ( .A(n14774), .B(n14021), .Z(n14134) );
  XOR U16175 ( .A(n14720), .B(n14134), .Z(n14113) );
  NAND U16176 ( .A(x[487]), .B(y[7813]), .Z(n14111) );
  XOR U16177 ( .A(n14112), .B(n14111), .Z(n14114) );
  AND U16178 ( .A(y[7808]), .B(x[492]), .Z(n14023) );
  NAND U16179 ( .A(y[7820]), .B(x[480]), .Z(n14022) );
  XNOR U16180 ( .A(n14023), .B(n14022), .Z(n14127) );
  NAND U16181 ( .A(x[491]), .B(y[7809]), .Z(n14108) );
  XNOR U16182 ( .A(o[140]), .B(n14108), .Z(n14128) );
  XOR U16183 ( .A(n14127), .B(n14128), .Z(n14097) );
  AND U16184 ( .A(y[7818]), .B(x[482]), .Z(n14025) );
  NAND U16185 ( .A(y[7812]), .B(x[488]), .Z(n14024) );
  XNOR U16186 ( .A(n14025), .B(n14024), .Z(n14102) );
  XOR U16187 ( .A(n14097), .B(n14096), .Z(n14098) );
  XNOR U16188 ( .A(n14092), .B(n14093), .Z(n14142) );
  AND U16189 ( .A(x[491]), .B(y[7819]), .Z(n15114) );
  NAND U16190 ( .A(n15114), .B(n14320), .Z(n14029) );
  NAND U16191 ( .A(n14027), .B(n14026), .Z(n14028) );
  NAND U16192 ( .A(n14029), .B(n14028), .Z(n14119) );
  AND U16193 ( .A(x[487]), .B(y[7810]), .Z(n14260) );
  AND U16194 ( .A(x[489]), .B(y[7812]), .Z(n14030) );
  NAND U16195 ( .A(n14260), .B(n14030), .Z(n14034) );
  NAND U16196 ( .A(n14032), .B(n14031), .Z(n14033) );
  NAND U16197 ( .A(n14034), .B(n14033), .Z(n14117) );
  NAND U16198 ( .A(y[7819]), .B(x[481]), .Z(n14035) );
  XNOR U16199 ( .A(n14036), .B(n14035), .Z(n14124) );
  AND U16200 ( .A(o[139]), .B(n14037), .Z(n14123) );
  XOR U16201 ( .A(n14124), .B(n14123), .Z(n14118) );
  XOR U16202 ( .A(n14117), .B(n14118), .Z(n14120) );
  XOR U16203 ( .A(n14119), .B(n14120), .Z(n14141) );
  XOR U16204 ( .A(n14142), .B(n14141), .Z(n14143) );
  XNOR U16205 ( .A(n14144), .B(n14143), .Z(n14072) );
  NAND U16206 ( .A(n14039), .B(n14038), .Z(n14043) );
  NAND U16207 ( .A(n14041), .B(n14040), .Z(n14042) );
  NAND U16208 ( .A(n14043), .B(n14042), .Z(n14071) );
  XOR U16209 ( .A(n14072), .B(n14071), .Z(n14074) );
  NANDN U16210 ( .A(n15006), .B(n14044), .Z(n14048) );
  NAND U16211 ( .A(n14046), .B(n14045), .Z(n14047) );
  NAND U16212 ( .A(n14048), .B(n14047), .Z(n14085) );
  NAND U16213 ( .A(n14050), .B(n14049), .Z(n14054) );
  NAND U16214 ( .A(n14052), .B(n14051), .Z(n14053) );
  AND U16215 ( .A(n14054), .B(n14053), .Z(n14084) );
  XOR U16216 ( .A(n14085), .B(n14084), .Z(n14086) );
  NAND U16217 ( .A(n14056), .B(n14055), .Z(n14060) );
  NAND U16218 ( .A(n14058), .B(n14057), .Z(n14059) );
  AND U16219 ( .A(n14060), .B(n14059), .Z(n14087) );
  XOR U16220 ( .A(n14086), .B(n14087), .Z(n14073) );
  XNOR U16221 ( .A(n14074), .B(n14073), .Z(n14081) );
  NAND U16222 ( .A(n14065), .B(n14064), .Z(n14069) );
  NANDN U16223 ( .A(n14067), .B(n14066), .Z(n14068) );
  AND U16224 ( .A(n14069), .B(n14068), .Z(n14079) );
  IV U16225 ( .A(n14079), .Z(n14077) );
  XOR U16226 ( .A(n14078), .B(n14077), .Z(n14070) );
  XNOR U16227 ( .A(n14081), .B(n14070), .Z(N301) );
  NAND U16228 ( .A(n14072), .B(n14071), .Z(n14076) );
  NAND U16229 ( .A(n14074), .B(n14073), .Z(n14075) );
  AND U16230 ( .A(n14076), .B(n14075), .Z(n14155) );
  NANDN U16231 ( .A(n14077), .B(n14078), .Z(n14083) );
  NOR U16232 ( .A(n14079), .B(n14078), .Z(n14080) );
  OR U16233 ( .A(n14081), .B(n14080), .Z(n14082) );
  AND U16234 ( .A(n14083), .B(n14082), .Z(n14154) );
  NAND U16235 ( .A(n14085), .B(n14084), .Z(n14089) );
  NAND U16236 ( .A(n14087), .B(n14086), .Z(n14088) );
  NAND U16237 ( .A(n14089), .B(n14088), .Z(n14151) );
  NAND U16238 ( .A(n14091), .B(n14090), .Z(n14095) );
  NANDN U16239 ( .A(n14093), .B(n14092), .Z(n14094) );
  NAND U16240 ( .A(n14095), .B(n14094), .Z(n14210) );
  NAND U16241 ( .A(n14097), .B(n14096), .Z(n14101) );
  NANDN U16242 ( .A(n14099), .B(n14098), .Z(n14100) );
  NAND U16243 ( .A(n14101), .B(n14100), .Z(n14218) );
  AND U16244 ( .A(y[7818]), .B(x[488]), .Z(n15393) );
  AND U16245 ( .A(x[482]), .B(y[7812]), .Z(n14270) );
  NAND U16246 ( .A(n15393), .B(n14270), .Z(n14105) );
  NANDN U16247 ( .A(n14103), .B(n14102), .Z(n14104) );
  NAND U16248 ( .A(n14105), .B(n14104), .Z(n14182) );
  NAND U16249 ( .A(y[7820]), .B(x[481]), .Z(n14106) );
  XNOR U16250 ( .A(n14107), .B(n14106), .Z(n14175) );
  ANDN U16251 ( .B(o[140]), .A(n14108), .Z(n14174) );
  XOR U16252 ( .A(n14175), .B(n14174), .Z(n14179) );
  AND U16253 ( .A(x[486]), .B(y[7815]), .Z(n15152) );
  AND U16254 ( .A(y[7819]), .B(x[482]), .Z(n14110) );
  NAND U16255 ( .A(y[7812]), .B(x[489]), .Z(n14109) );
  XOR U16256 ( .A(n14110), .B(n14109), .Z(n14186) );
  XNOR U16257 ( .A(n15152), .B(n14186), .Z(n14180) );
  XOR U16258 ( .A(n14179), .B(n14180), .Z(n14181) );
  XOR U16259 ( .A(n14182), .B(n14181), .Z(n14217) );
  NAND U16260 ( .A(n14112), .B(n14111), .Z(n14116) );
  ANDN U16261 ( .B(n14114), .A(n14113), .Z(n14115) );
  ANDN U16262 ( .B(n14116), .A(n14115), .Z(n14216) );
  XOR U16263 ( .A(n14217), .B(n14216), .Z(n14219) );
  XOR U16264 ( .A(n14218), .B(n14219), .Z(n14211) );
  XOR U16265 ( .A(n14210), .B(n14211), .Z(n14213) );
  NAND U16266 ( .A(n14118), .B(n14117), .Z(n14122) );
  NAND U16267 ( .A(n14120), .B(n14119), .Z(n14121) );
  NAND U16268 ( .A(n14122), .B(n14121), .Z(n14159) );
  NAND U16269 ( .A(x[486]), .B(y[7819]), .Z(n14542) );
  AND U16270 ( .A(x[481]), .B(y[7814]), .Z(n14173) );
  NANDN U16271 ( .A(n14542), .B(n14173), .Z(n14126) );
  NAND U16272 ( .A(n14124), .B(n14123), .Z(n14125) );
  NAND U16273 ( .A(n14126), .B(n14125), .Z(n14166) );
  AND U16274 ( .A(x[492]), .B(y[7820]), .Z(n15399) );
  NAND U16275 ( .A(n15399), .B(n14320), .Z(n14130) );
  NAND U16276 ( .A(n14128), .B(n14127), .Z(n14129) );
  NAND U16277 ( .A(n14130), .B(n14129), .Z(n14164) );
  AND U16278 ( .A(x[490]), .B(y[7811]), .Z(n15018) );
  AND U16279 ( .A(y[7810]), .B(x[491]), .Z(n14979) );
  NAND U16280 ( .A(y[7813]), .B(x[488]), .Z(n14131) );
  XOR U16281 ( .A(n14979), .B(n14131), .Z(n14170) );
  XNOR U16282 ( .A(n15018), .B(n14170), .Z(n14163) );
  XOR U16283 ( .A(n14164), .B(n14163), .Z(n14165) );
  XOR U16284 ( .A(n14166), .B(n14165), .Z(n14157) );
  AND U16285 ( .A(x[490]), .B(y[7816]), .Z(n14133) );
  AND U16286 ( .A(x[484]), .B(y[7810]), .Z(n14132) );
  NAND U16287 ( .A(n14133), .B(n14132), .Z(n14136) );
  NAND U16288 ( .A(n14720), .B(n14134), .Z(n14135) );
  NAND U16289 ( .A(n14136), .B(n14135), .Z(n14206) );
  AND U16290 ( .A(y[7808]), .B(x[493]), .Z(n14138) );
  NAND U16291 ( .A(y[7821]), .B(x[480]), .Z(n14137) );
  XNOR U16292 ( .A(n14138), .B(n14137), .Z(n14198) );
  NAND U16293 ( .A(x[492]), .B(y[7809]), .Z(n14191) );
  XOR U16294 ( .A(o[141]), .B(n14191), .Z(n14199) );
  XNOR U16295 ( .A(n14198), .B(n14199), .Z(n14205) );
  AND U16296 ( .A(y[7816]), .B(x[485]), .Z(n14140) );
  NAND U16297 ( .A(y[7818]), .B(x[483]), .Z(n14139) );
  XNOR U16298 ( .A(n14140), .B(n14139), .Z(n14194) );
  NAND U16299 ( .A(x[484]), .B(y[7817]), .Z(n14195) );
  XNOR U16300 ( .A(n14194), .B(n14195), .Z(n14204) );
  XOR U16301 ( .A(n14205), .B(n14204), .Z(n14207) );
  XNOR U16302 ( .A(n14206), .B(n14207), .Z(n14158) );
  XOR U16303 ( .A(n14159), .B(n14160), .Z(n14212) );
  XNOR U16304 ( .A(n14213), .B(n14212), .Z(n14149) );
  NAND U16305 ( .A(n14142), .B(n14141), .Z(n14146) );
  NAND U16306 ( .A(n14144), .B(n14143), .Z(n14145) );
  AND U16307 ( .A(n14146), .B(n14145), .Z(n14148) );
  XOR U16308 ( .A(n14149), .B(n14148), .Z(n14150) );
  XOR U16309 ( .A(n14151), .B(n14150), .Z(n14156) );
  XNOR U16310 ( .A(n14154), .B(n14156), .Z(n14147) );
  XOR U16311 ( .A(n14155), .B(n14147), .Z(N302) );
  NAND U16312 ( .A(n14149), .B(n14148), .Z(n14153) );
  NAND U16313 ( .A(n14151), .B(n14150), .Z(n14152) );
  NAND U16314 ( .A(n14153), .B(n14152), .Z(n14231) );
  IV U16315 ( .A(n14231), .Z(n14229) );
  NANDN U16316 ( .A(n14158), .B(n14157), .Z(n14162) );
  NAND U16317 ( .A(n14160), .B(n14159), .Z(n14161) );
  NAND U16318 ( .A(n14162), .B(n14161), .Z(n14238) );
  NAND U16319 ( .A(n14164), .B(n14163), .Z(n14168) );
  NAND U16320 ( .A(n14166), .B(n14165), .Z(n14167) );
  AND U16321 ( .A(n14168), .B(n14167), .Z(n14245) );
  AND U16322 ( .A(x[491]), .B(y[7813]), .Z(n14346) );
  NAND U16323 ( .A(n14346), .B(n14169), .Z(n14172) );
  NANDN U16324 ( .A(n14170), .B(n15018), .Z(n14171) );
  AND U16325 ( .A(n14172), .B(n14171), .Z(n14294) );
  AND U16326 ( .A(x[487]), .B(y[7820]), .Z(n14734) );
  XNOR U16327 ( .A(n14294), .B(n14293), .Z(n14296) );
  AND U16328 ( .A(x[484]), .B(y[7818]), .Z(n14647) );
  AND U16329 ( .A(y[7819]), .B(x[483]), .Z(n14177) );
  NAND U16330 ( .A(y[7814]), .B(x[488]), .Z(n14176) );
  XOR U16331 ( .A(n14177), .B(n14176), .Z(n14281) );
  XOR U16332 ( .A(n14540), .B(n14281), .Z(n14290) );
  XNOR U16333 ( .A(n14647), .B(n14290), .Z(n14292) );
  AND U16334 ( .A(x[489]), .B(y[7813]), .Z(n14844) );
  AND U16335 ( .A(x[482]), .B(y[7820]), .Z(n14178) );
  AND U16336 ( .A(y[7812]), .B(x[490]), .Z(n14862) );
  XOR U16337 ( .A(n14178), .B(n14862), .Z(n14271) );
  XOR U16338 ( .A(n14844), .B(n14271), .Z(n14291) );
  XOR U16339 ( .A(n14292), .B(n14291), .Z(n14295) );
  XNOR U16340 ( .A(n14296), .B(n14295), .Z(n14243) );
  NAND U16341 ( .A(n14180), .B(n14179), .Z(n14184) );
  NAND U16342 ( .A(n14182), .B(n14181), .Z(n14183) );
  AND U16343 ( .A(n14184), .B(n14183), .Z(n14242) );
  XOR U16344 ( .A(n14243), .B(n14242), .Z(n14244) );
  XOR U16345 ( .A(n14245), .B(n14244), .Z(n14237) );
  AND U16346 ( .A(x[489]), .B(y[7819]), .Z(n14185) );
  NAND U16347 ( .A(n14185), .B(n14270), .Z(n14188) );
  NANDN U16348 ( .A(n14186), .B(n15152), .Z(n14187) );
  AND U16349 ( .A(n14188), .B(n14187), .Z(n14257) );
  AND U16350 ( .A(y[7808]), .B(x[494]), .Z(n14190) );
  NAND U16351 ( .A(y[7822]), .B(x[480]), .Z(n14189) );
  XNOR U16352 ( .A(n14190), .B(n14189), .Z(n14278) );
  ANDN U16353 ( .B(o[141]), .A(n14191), .Z(n14277) );
  XOR U16354 ( .A(n14278), .B(n14277), .Z(n14254) );
  NAND U16355 ( .A(y[7810]), .B(x[492]), .Z(n14192) );
  XNOR U16356 ( .A(n14193), .B(n14192), .Z(n14261) );
  NAND U16357 ( .A(x[493]), .B(y[7809]), .Z(n14269) );
  XOR U16358 ( .A(o[142]), .B(n14269), .Z(n14262) );
  XOR U16359 ( .A(n14261), .B(n14262), .Z(n14255) );
  XNOR U16360 ( .A(n14254), .B(n14255), .Z(n14256) );
  XOR U16361 ( .A(n14257), .B(n14256), .Z(n14300) );
  AND U16362 ( .A(x[485]), .B(y[7818]), .Z(n14333) );
  NAND U16363 ( .A(n15006), .B(n14333), .Z(n14197) );
  NANDN U16364 ( .A(n14195), .B(n14194), .Z(n14196) );
  AND U16365 ( .A(n14197), .B(n14196), .Z(n14250) );
  AND U16366 ( .A(x[493]), .B(y[7821]), .Z(n15711) );
  NAND U16367 ( .A(n15711), .B(n14320), .Z(n14201) );
  NANDN U16368 ( .A(n14199), .B(n14198), .Z(n14200) );
  AND U16369 ( .A(n14201), .B(n14200), .Z(n14249) );
  NAND U16370 ( .A(y[7811]), .B(x[491]), .Z(n14202) );
  XNOR U16371 ( .A(n14203), .B(n14202), .Z(n14276) );
  AND U16372 ( .A(x[481]), .B(y[7821]), .Z(n14275) );
  XOR U16373 ( .A(n14276), .B(n14275), .Z(n14248) );
  XOR U16374 ( .A(n14249), .B(n14248), .Z(n14251) );
  XNOR U16375 ( .A(n14250), .B(n14251), .Z(n14299) );
  XOR U16376 ( .A(n14300), .B(n14299), .Z(n14302) );
  NAND U16377 ( .A(n14205), .B(n14204), .Z(n14209) );
  NAND U16378 ( .A(n14207), .B(n14206), .Z(n14208) );
  AND U16379 ( .A(n14209), .B(n14208), .Z(n14301) );
  XNOR U16380 ( .A(n14302), .B(n14301), .Z(n14236) );
  XOR U16381 ( .A(n14238), .B(n14239), .Z(n14225) );
  NAND U16382 ( .A(n14211), .B(n14210), .Z(n14215) );
  NAND U16383 ( .A(n14213), .B(n14212), .Z(n14214) );
  NAND U16384 ( .A(n14215), .B(n14214), .Z(n14224) );
  NAND U16385 ( .A(n14217), .B(n14216), .Z(n14221) );
  NAND U16386 ( .A(n14219), .B(n14218), .Z(n14220) );
  NAND U16387 ( .A(n14221), .B(n14220), .Z(n14223) );
  XNOR U16388 ( .A(n14224), .B(n14223), .Z(n14226) );
  XNOR U16389 ( .A(n14230), .B(n14232), .Z(n14222) );
  XOR U16390 ( .A(n14229), .B(n14222), .Z(N303) );
  NAND U16391 ( .A(n14224), .B(n14223), .Z(n14228) );
  NANDN U16392 ( .A(n14226), .B(n14225), .Z(n14227) );
  AND U16393 ( .A(n14228), .B(n14227), .Z(n14312) );
  NANDN U16394 ( .A(n14229), .B(n14230), .Z(n14235) );
  NOR U16395 ( .A(n14231), .B(n14230), .Z(n14233) );
  OR U16396 ( .A(n14233), .B(n14232), .Z(n14234) );
  AND U16397 ( .A(n14235), .B(n14234), .Z(n14313) );
  NANDN U16398 ( .A(n14237), .B(n14236), .Z(n14241) );
  NAND U16399 ( .A(n14239), .B(n14238), .Z(n14240) );
  NAND U16400 ( .A(n14241), .B(n14240), .Z(n14308) );
  NAND U16401 ( .A(n14243), .B(n14242), .Z(n14247) );
  NAND U16402 ( .A(n14245), .B(n14244), .Z(n14246) );
  NAND U16403 ( .A(n14247), .B(n14246), .Z(n14374) );
  NANDN U16404 ( .A(n14249), .B(n14248), .Z(n14253) );
  OR U16405 ( .A(n14251), .B(n14250), .Z(n14252) );
  NAND U16406 ( .A(n14253), .B(n14252), .Z(n14379) );
  NANDN U16407 ( .A(n14255), .B(n14254), .Z(n14259) );
  NANDN U16408 ( .A(n14257), .B(n14256), .Z(n14258) );
  NAND U16409 ( .A(n14259), .B(n14258), .Z(n14377) );
  AND U16410 ( .A(x[492]), .B(y[7815]), .Z(n14726) );
  NAND U16411 ( .A(n14726), .B(n14260), .Z(n14264) );
  NANDN U16412 ( .A(n14262), .B(n14261), .Z(n14263) );
  AND U16413 ( .A(n14264), .B(n14263), .Z(n14353) );
  AND U16414 ( .A(y[7812]), .B(x[491]), .Z(n14266) );
  NAND U16415 ( .A(y[7810]), .B(x[493]), .Z(n14265) );
  XNOR U16416 ( .A(n14266), .B(n14265), .Z(n14358) );
  AND U16417 ( .A(x[492]), .B(y[7811]), .Z(n14357) );
  XOR U16418 ( .A(n14358), .B(n14357), .Z(n14352) );
  AND U16419 ( .A(y[7808]), .B(x[495]), .Z(n14268) );
  NAND U16420 ( .A(y[7823]), .B(x[480]), .Z(n14267) );
  XNOR U16421 ( .A(n14268), .B(n14267), .Z(n14322) );
  ANDN U16422 ( .B(o[142]), .A(n14269), .Z(n14321) );
  XNOR U16423 ( .A(n14322), .B(n14321), .Z(n14351) );
  XOR U16424 ( .A(n14352), .B(n14351), .Z(n14354) );
  XOR U16425 ( .A(n14353), .B(n14354), .Z(n14385) );
  NAND U16426 ( .A(x[490]), .B(y[7820]), .Z(n15154) );
  NANDN U16427 ( .A(n15154), .B(n14270), .Z(n14273) );
  NAND U16428 ( .A(n14844), .B(n14271), .Z(n14272) );
  NAND U16429 ( .A(n14273), .B(n14272), .Z(n14383) );
  AND U16430 ( .A(x[491]), .B(y[7816]), .Z(n14646) );
  XNOR U16431 ( .A(n14383), .B(n14384), .Z(n14386) );
  XOR U16432 ( .A(n14385), .B(n14386), .Z(n14378) );
  XOR U16433 ( .A(n14377), .B(n14378), .Z(n14380) );
  XOR U16434 ( .A(n14379), .B(n14380), .Z(n14371) );
  AND U16435 ( .A(x[494]), .B(y[7822]), .Z(n15946) );
  AND U16436 ( .A(x[488]), .B(y[7819]), .Z(n14279) );
  NANDN U16437 ( .A(n14280), .B(n14279), .Z(n14283) );
  NANDN U16438 ( .A(n14281), .B(n14540), .Z(n14282) );
  NAND U16439 ( .A(n14283), .B(n14282), .Z(n14347) );
  XNOR U16440 ( .A(n14348), .B(n14347), .Z(n14350) );
  AND U16441 ( .A(y[7813]), .B(x[490]), .Z(n14285) );
  NAND U16442 ( .A(y[7819]), .B(x[484]), .Z(n14284) );
  XNOR U16443 ( .A(n14285), .B(n14284), .Z(n14328) );
  AND U16444 ( .A(x[487]), .B(y[7816]), .Z(n14327) );
  XOR U16445 ( .A(n14328), .B(n14327), .Z(n14335) );
  NAND U16446 ( .A(x[486]), .B(y[7817]), .Z(n14417) );
  XNOR U16447 ( .A(n14417), .B(n14333), .Z(n14334) );
  XOR U16448 ( .A(n14335), .B(n14334), .Z(n14367) );
  AND U16449 ( .A(y[7821]), .B(x[482]), .Z(n14287) );
  NAND U16450 ( .A(y[7814]), .B(x[489]), .Z(n14286) );
  XNOR U16451 ( .A(n14287), .B(n14286), .Z(n14338) );
  NAND U16452 ( .A(x[483]), .B(y[7820]), .Z(n14339) );
  XNOR U16453 ( .A(n14338), .B(n14339), .Z(n14365) );
  AND U16454 ( .A(y[7822]), .B(x[481]), .Z(n14289) );
  NAND U16455 ( .A(y[7815]), .B(x[488]), .Z(n14288) );
  XNOR U16456 ( .A(n14289), .B(n14288), .Z(n14316) );
  NAND U16457 ( .A(x[494]), .B(y[7809]), .Z(n14344) );
  XOR U16458 ( .A(o[143]), .B(n14344), .Z(n14317) );
  XNOR U16459 ( .A(n14316), .B(n14317), .Z(n14366) );
  XOR U16460 ( .A(n14365), .B(n14366), .Z(n14368) );
  XOR U16461 ( .A(n14367), .B(n14368), .Z(n14349) );
  XOR U16462 ( .A(n14350), .B(n14349), .Z(n14388) );
  XNOR U16463 ( .A(n14388), .B(n14387), .Z(n14390) );
  NANDN U16464 ( .A(n14294), .B(n14293), .Z(n14298) );
  NAND U16465 ( .A(n14296), .B(n14295), .Z(n14297) );
  AND U16466 ( .A(n14298), .B(n14297), .Z(n14389) );
  XOR U16467 ( .A(n14390), .B(n14389), .Z(n14372) );
  XOR U16468 ( .A(n14371), .B(n14372), .Z(n14373) );
  XOR U16469 ( .A(n14374), .B(n14373), .Z(n14307) );
  NAND U16470 ( .A(n14300), .B(n14299), .Z(n14304) );
  NAND U16471 ( .A(n14302), .B(n14301), .Z(n14303) );
  AND U16472 ( .A(n14304), .B(n14303), .Z(n14306) );
  XOR U16473 ( .A(n14308), .B(n14309), .Z(n14314) );
  XNOR U16474 ( .A(n14313), .B(n14314), .Z(n14305) );
  XOR U16475 ( .A(n14312), .B(n14305), .Z(N304) );
  NANDN U16476 ( .A(n14307), .B(n14306), .Z(n14311) );
  NAND U16477 ( .A(n14309), .B(n14308), .Z(n14310) );
  AND U16478 ( .A(n14311), .B(n14310), .Z(n14482) );
  AND U16479 ( .A(x[488]), .B(y[7822]), .Z(n14648) );
  NAND U16480 ( .A(n14648), .B(n14315), .Z(n14319) );
  NANDN U16481 ( .A(n14317), .B(n14316), .Z(n14318) );
  NAND U16482 ( .A(n14319), .B(n14318), .Z(n14447) );
  AND U16483 ( .A(x[495]), .B(y[7823]), .Z(n16388) );
  NAND U16484 ( .A(n16388), .B(n14320), .Z(n14324) );
  NAND U16485 ( .A(n14322), .B(n14321), .Z(n14323) );
  NAND U16486 ( .A(n14324), .B(n14323), .Z(n14446) );
  XOR U16487 ( .A(n14447), .B(n14446), .Z(n14449) );
  AND U16488 ( .A(x[490]), .B(y[7819]), .Z(n14326) );
  NAND U16489 ( .A(n14326), .B(n14325), .Z(n14330) );
  NAND U16490 ( .A(n14328), .B(n14327), .Z(n14329) );
  NAND U16491 ( .A(n14330), .B(n14329), .Z(n14404) );
  AND U16492 ( .A(x[480]), .B(y[7824]), .Z(n14426) );
  AND U16493 ( .A(x[496]), .B(y[7808]), .Z(n14427) );
  XOR U16494 ( .A(n14426), .B(n14427), .Z(n14429) );
  NAND U16495 ( .A(x[495]), .B(y[7809]), .Z(n14414) );
  XOR U16496 ( .A(n14429), .B(n14428), .Z(n14403) );
  NAND U16497 ( .A(y[7817]), .B(x[487]), .Z(n14331) );
  XNOR U16498 ( .A(n14332), .B(n14331), .Z(n14419) );
  AND U16499 ( .A(x[490]), .B(y[7814]), .Z(n14418) );
  XOR U16500 ( .A(n14419), .B(n14418), .Z(n14402) );
  XOR U16501 ( .A(n14403), .B(n14402), .Z(n14405) );
  XOR U16502 ( .A(n14404), .B(n14405), .Z(n14448) );
  XOR U16503 ( .A(n14449), .B(n14448), .Z(n14399) );
  NANDN U16504 ( .A(n14333), .B(n14417), .Z(n14337) );
  NANDN U16505 ( .A(n14335), .B(n14334), .Z(n14336) );
  AND U16506 ( .A(n14337), .B(n14336), .Z(n14397) );
  NAND U16507 ( .A(x[489]), .B(y[7821]), .Z(n15135) );
  NANDN U16508 ( .A(n15135), .B(n14725), .Z(n14341) );
  NANDN U16509 ( .A(n14339), .B(n14338), .Z(n14340) );
  AND U16510 ( .A(n14341), .B(n14340), .Z(n14437) );
  AND U16511 ( .A(y[7823]), .B(x[481]), .Z(n14343) );
  NAND U16512 ( .A(y[7816]), .B(x[488]), .Z(n14342) );
  XNOR U16513 ( .A(n14343), .B(n14342), .Z(n14423) );
  ANDN U16514 ( .B(o[143]), .A(n14344), .Z(n14422) );
  XOR U16515 ( .A(n14423), .B(n14422), .Z(n14435) );
  NAND U16516 ( .A(y[7810]), .B(x[494]), .Z(n14345) );
  XNOR U16517 ( .A(n14346), .B(n14345), .Z(n14458) );
  AND U16518 ( .A(x[484]), .B(y[7820]), .Z(n14459) );
  XOR U16519 ( .A(n14458), .B(n14459), .Z(n14434) );
  XOR U16520 ( .A(n14435), .B(n14434), .Z(n14436) );
  XOR U16521 ( .A(n14437), .B(n14436), .Z(n14396) );
  XNOR U16522 ( .A(n14397), .B(n14396), .Z(n14398) );
  XNOR U16523 ( .A(n14399), .B(n14398), .Z(n14440) );
  XNOR U16524 ( .A(n14440), .B(n14441), .Z(n14443) );
  NANDN U16525 ( .A(n14352), .B(n14351), .Z(n14356) );
  NANDN U16526 ( .A(n14354), .B(n14353), .Z(n14355) );
  NAND U16527 ( .A(n14356), .B(n14355), .Z(n14473) );
  AND U16528 ( .A(x[493]), .B(y[7812]), .Z(n14469) );
  NAND U16529 ( .A(n14979), .B(n14469), .Z(n14360) );
  NAND U16530 ( .A(n14358), .B(n14357), .Z(n14359) );
  NAND U16531 ( .A(n14360), .B(n14359), .Z(n14455) );
  AND U16532 ( .A(y[7822]), .B(x[482]), .Z(n14362) );
  NAND U16533 ( .A(y[7815]), .B(x[489]), .Z(n14361) );
  XNOR U16534 ( .A(n14362), .B(n14361), .Z(n14462) );
  AND U16535 ( .A(x[483]), .B(y[7821]), .Z(n14463) );
  XOR U16536 ( .A(n14462), .B(n14463), .Z(n14452) );
  AND U16537 ( .A(x[492]), .B(y[7812]), .Z(n15123) );
  AND U16538 ( .A(y[7819]), .B(x[485]), .Z(n14364) );
  NAND U16539 ( .A(y[7811]), .B(x[493]), .Z(n14363) );
  XOR U16540 ( .A(n14364), .B(n14363), .Z(n14409) );
  XNOR U16541 ( .A(n15123), .B(n14409), .Z(n14453) );
  XOR U16542 ( .A(n14452), .B(n14453), .Z(n14454) );
  XNOR U16543 ( .A(n14455), .B(n14454), .Z(n14470) );
  NAND U16544 ( .A(n14366), .B(n14365), .Z(n14370) );
  NAND U16545 ( .A(n14368), .B(n14367), .Z(n14369) );
  AND U16546 ( .A(n14370), .B(n14369), .Z(n14471) );
  XOR U16547 ( .A(n14470), .B(n14471), .Z(n14472) );
  XOR U16548 ( .A(n14473), .B(n14472), .Z(n14442) );
  XNOR U16549 ( .A(n14443), .B(n14442), .Z(n14477) );
  NAND U16550 ( .A(n14372), .B(n14371), .Z(n14376) );
  NAND U16551 ( .A(n14374), .B(n14373), .Z(n14375) );
  AND U16552 ( .A(n14376), .B(n14375), .Z(n14476) );
  XOR U16553 ( .A(n14477), .B(n14476), .Z(n14479) );
  NANDN U16554 ( .A(n14378), .B(n14377), .Z(n14382) );
  NANDN U16555 ( .A(n14380), .B(n14379), .Z(n14381) );
  NAND U16556 ( .A(n14382), .B(n14381), .Z(n14394) );
  XOR U16557 ( .A(n14392), .B(n14393), .Z(n14395) );
  XOR U16558 ( .A(n14394), .B(n14395), .Z(n14478) );
  XOR U16559 ( .A(n14479), .B(n14478), .Z(n14484) );
  XNOR U16560 ( .A(n14483), .B(n14484), .Z(n14391) );
  XOR U16561 ( .A(n14482), .B(n14391), .Z(N305) );
  NANDN U16562 ( .A(n14397), .B(n14396), .Z(n14401) );
  NANDN U16563 ( .A(n14399), .B(n14398), .Z(n14400) );
  NAND U16564 ( .A(n14401), .B(n14400), .Z(n14495) );
  NAND U16565 ( .A(n14403), .B(n14402), .Z(n14407) );
  NAND U16566 ( .A(n14405), .B(n14404), .Z(n14406) );
  NAND U16567 ( .A(n14407), .B(n14406), .Z(n14577) );
  AND U16568 ( .A(x[493]), .B(y[7819]), .Z(n15407) );
  NAND U16569 ( .A(n15407), .B(n14408), .Z(n14411) );
  NANDN U16570 ( .A(n14409), .B(n15123), .Z(n14410) );
  NAND U16571 ( .A(n14411), .B(n14410), .Z(n14525) );
  AND U16572 ( .A(y[7824]), .B(x[481]), .Z(n14413) );
  NAND U16573 ( .A(y[7816]), .B(x[489]), .Z(n14412) );
  XNOR U16574 ( .A(n14413), .B(n14412), .Z(n14546) );
  ANDN U16575 ( .B(o[144]), .A(n14414), .Z(n14545) );
  XOR U16576 ( .A(n14546), .B(n14545), .Z(n14523) );
  AND U16577 ( .A(y[7810]), .B(x[495]), .Z(n14416) );
  NAND U16578 ( .A(y[7813]), .B(x[492]), .Z(n14415) );
  XNOR U16579 ( .A(n14416), .B(n14415), .Z(n14498) );
  NAND U16580 ( .A(x[494]), .B(y[7811]), .Z(n14499) );
  XOR U16581 ( .A(n14523), .B(n14522), .Z(n14524) );
  XOR U16582 ( .A(n14525), .B(n14524), .Z(n14575) );
  NAND U16583 ( .A(x[487]), .B(y[7818]), .Z(n14557) );
  IV U16584 ( .A(n14557), .Z(n14467) );
  NANDN U16585 ( .A(n14417), .B(n14467), .Z(n14421) );
  NAND U16586 ( .A(n14419), .B(n14418), .Z(n14420) );
  NAND U16587 ( .A(n14421), .B(n14420), .Z(n14535) );
  NAND U16588 ( .A(x[488]), .B(y[7823]), .Z(n15210) );
  AND U16589 ( .A(x[481]), .B(y[7816]), .Z(n14626) );
  NANDN U16590 ( .A(n15210), .B(n14626), .Z(n14425) );
  NAND U16591 ( .A(n14423), .B(n14422), .Z(n14424) );
  NAND U16592 ( .A(n14425), .B(n14424), .Z(n14534) );
  XOR U16593 ( .A(n14535), .B(n14534), .Z(n14537) );
  NAND U16594 ( .A(n14427), .B(n14426), .Z(n14431) );
  NAND U16595 ( .A(n14429), .B(n14428), .Z(n14430) );
  NAND U16596 ( .A(n14431), .B(n14430), .Z(n14531) );
  AND U16597 ( .A(x[480]), .B(y[7825]), .Z(n14512) );
  NAND U16598 ( .A(x[497]), .B(y[7808]), .Z(n14513) );
  AND U16599 ( .A(x[496]), .B(y[7809]), .Z(n14509) );
  XOR U16600 ( .A(o[145]), .B(n14509), .Z(n14514) );
  XOR U16601 ( .A(n14515), .B(n14514), .Z(n14529) );
  AND U16602 ( .A(y[7823]), .B(x[482]), .Z(n14433) );
  NAND U16603 ( .A(y[7815]), .B(x[490]), .Z(n14432) );
  XNOR U16604 ( .A(n14433), .B(n14432), .Z(n14550) );
  NAND U16605 ( .A(x[483]), .B(y[7822]), .Z(n14551) );
  XOR U16606 ( .A(n14529), .B(n14528), .Z(n14530) );
  XOR U16607 ( .A(n14531), .B(n14530), .Z(n14536) );
  XOR U16608 ( .A(n14537), .B(n14536), .Z(n14574) );
  XOR U16609 ( .A(n14575), .B(n14574), .Z(n14576) );
  XNOR U16610 ( .A(n14577), .B(n14576), .Z(n14492) );
  NAND U16611 ( .A(n14435), .B(n14434), .Z(n14439) );
  NANDN U16612 ( .A(n14437), .B(n14436), .Z(n14438) );
  AND U16613 ( .A(n14439), .B(n14438), .Z(n14493) );
  XOR U16614 ( .A(n14492), .B(n14493), .Z(n14494) );
  XOR U16615 ( .A(n14495), .B(n14494), .Z(n14584) );
  NANDN U16616 ( .A(n14441), .B(n14440), .Z(n14445) );
  NAND U16617 ( .A(n14443), .B(n14442), .Z(n14444) );
  NAND U16618 ( .A(n14445), .B(n14444), .Z(n14489) );
  NAND U16619 ( .A(n14447), .B(n14446), .Z(n14451) );
  NAND U16620 ( .A(n14449), .B(n14448), .Z(n14450) );
  NAND U16621 ( .A(n14451), .B(n14450), .Z(n14571) );
  NAND U16622 ( .A(n14453), .B(n14452), .Z(n14457) );
  NAND U16623 ( .A(n14455), .B(n14454), .Z(n14456) );
  NAND U16624 ( .A(n14457), .B(n14456), .Z(n14569) );
  NAND U16625 ( .A(x[494]), .B(y[7813]), .Z(n14771) );
  NANDN U16626 ( .A(n14771), .B(n14979), .Z(n14461) );
  NAND U16627 ( .A(n14459), .B(n14458), .Z(n14460) );
  NAND U16628 ( .A(n14461), .B(n14460), .Z(n14563) );
  AND U16629 ( .A(x[489]), .B(y[7822]), .Z(n15388) );
  NAND U16630 ( .A(n14549), .B(n15388), .Z(n14465) );
  NAND U16631 ( .A(n14463), .B(n14462), .Z(n14464) );
  NAND U16632 ( .A(n14465), .B(n14464), .Z(n14562) );
  XOR U16633 ( .A(n14563), .B(n14562), .Z(n14565) );
  AND U16634 ( .A(x[485]), .B(y[7820]), .Z(n14608) );
  NAND U16635 ( .A(y[7817]), .B(x[488]), .Z(n14466) );
  XNOR U16636 ( .A(n14608), .B(n14466), .Z(n14541) );
  XOR U16637 ( .A(n14556), .B(n14467), .Z(n14559) );
  NAND U16638 ( .A(y[7821]), .B(x[484]), .Z(n14468) );
  XNOR U16639 ( .A(n14469), .B(n14468), .Z(n14503) );
  AND U16640 ( .A(x[491]), .B(y[7814]), .Z(n14504) );
  XOR U16641 ( .A(n14503), .B(n14504), .Z(n14558) );
  XOR U16642 ( .A(n14559), .B(n14558), .Z(n14564) );
  XOR U16643 ( .A(n14565), .B(n14564), .Z(n14568) );
  XOR U16644 ( .A(n14569), .B(n14568), .Z(n14570) );
  XNOR U16645 ( .A(n14571), .B(n14570), .Z(n14487) );
  NAND U16646 ( .A(n14471), .B(n14470), .Z(n14475) );
  NAND U16647 ( .A(n14473), .B(n14472), .Z(n14474) );
  NAND U16648 ( .A(n14475), .B(n14474), .Z(n14486) );
  XOR U16649 ( .A(n14487), .B(n14486), .Z(n14488) );
  XOR U16650 ( .A(n14489), .B(n14488), .Z(n14583) );
  XNOR U16651 ( .A(n14584), .B(n14583), .Z(n14586) );
  XOR U16652 ( .A(n14585), .B(n14586), .Z(n14582) );
  NAND U16653 ( .A(n14477), .B(n14476), .Z(n14481) );
  NAND U16654 ( .A(n14479), .B(n14478), .Z(n14480) );
  NAND U16655 ( .A(n14481), .B(n14480), .Z(n14581) );
  XOR U16656 ( .A(n14581), .B(n14580), .Z(n14485) );
  XNOR U16657 ( .A(n14582), .B(n14485), .Z(N306) );
  NAND U16658 ( .A(n14487), .B(n14486), .Z(n14491) );
  NAND U16659 ( .A(n14489), .B(n14488), .Z(n14490) );
  AND U16660 ( .A(n14491), .B(n14490), .Z(n14695) );
  NAND U16661 ( .A(n14493), .B(n14492), .Z(n14497) );
  NAND U16662 ( .A(n14495), .B(n14494), .Z(n14496) );
  AND U16663 ( .A(n14497), .B(n14496), .Z(n14693) );
  AND U16664 ( .A(x[495]), .B(y[7813]), .Z(n14733) );
  AND U16665 ( .A(x[492]), .B(y[7810]), .Z(n14837) );
  NAND U16666 ( .A(n14733), .B(n14837), .Z(n14501) );
  NANDN U16667 ( .A(n14499), .B(n14498), .Z(n14500) );
  NAND U16668 ( .A(n14501), .B(n14500), .Z(n14675) );
  NAND U16669 ( .A(n15711), .B(n14502), .Z(n14506) );
  NAND U16670 ( .A(n14504), .B(n14503), .Z(n14505) );
  NAND U16671 ( .A(n14506), .B(n14505), .Z(n14664) );
  AND U16672 ( .A(y[7825]), .B(x[481]), .Z(n14508) );
  NAND U16673 ( .A(y[7816]), .B(x[490]), .Z(n14507) );
  XNOR U16674 ( .A(n14508), .B(n14507), .Z(n14628) );
  AND U16675 ( .A(n14509), .B(o[145]), .Z(n14627) );
  XOR U16676 ( .A(n14628), .B(n14627), .Z(n14663) );
  AND U16677 ( .A(y[7811]), .B(x[495]), .Z(n14511) );
  NAND U16678 ( .A(y[7817]), .B(x[489]), .Z(n14510) );
  XNOR U16679 ( .A(n14511), .B(n14510), .Z(n14619) );
  AND U16680 ( .A(x[494]), .B(y[7812]), .Z(n14618) );
  XOR U16681 ( .A(n14619), .B(n14618), .Z(n14662) );
  XOR U16682 ( .A(n14663), .B(n14662), .Z(n14665) );
  XOR U16683 ( .A(n14664), .B(n14665), .Z(n14674) );
  XOR U16684 ( .A(n14675), .B(n14674), .Z(n14677) );
  NANDN U16685 ( .A(n14513), .B(n14512), .Z(n14517) );
  NAND U16686 ( .A(n14515), .B(n14514), .Z(n14516) );
  AND U16687 ( .A(n14517), .B(n14516), .Z(n14687) );
  AND U16688 ( .A(y[7810]), .B(x[496]), .Z(n14519) );
  NAND U16689 ( .A(y[7815]), .B(x[491]), .Z(n14518) );
  XNOR U16690 ( .A(n14519), .B(n14518), .Z(n14615) );
  AND U16691 ( .A(x[482]), .B(y[7824]), .Z(n14614) );
  XOR U16692 ( .A(n14615), .B(n14614), .Z(n14686) );
  AND U16693 ( .A(y[7821]), .B(x[485]), .Z(n14753) );
  NAND U16694 ( .A(y[7820]), .B(x[486]), .Z(n14520) );
  XNOR U16695 ( .A(n14753), .B(n14520), .Z(n14611) );
  NAND U16696 ( .A(y[7822]), .B(x[484]), .Z(n14521) );
  XNOR U16697 ( .A(n15393), .B(n14521), .Z(n14650) );
  AND U16698 ( .A(x[487]), .B(y[7819]), .Z(n14649) );
  XOR U16699 ( .A(n14650), .B(n14649), .Z(n14610) );
  XOR U16700 ( .A(n14611), .B(n14610), .Z(n14688) );
  XOR U16701 ( .A(n14689), .B(n14688), .Z(n14676) );
  XNOR U16702 ( .A(n14677), .B(n14676), .Z(n14597) );
  NAND U16703 ( .A(n14523), .B(n14522), .Z(n14527) );
  NAND U16704 ( .A(n14525), .B(n14524), .Z(n14526) );
  AND U16705 ( .A(n14527), .B(n14526), .Z(n14668) );
  NAND U16706 ( .A(n14529), .B(n14528), .Z(n14533) );
  NAND U16707 ( .A(n14531), .B(n14530), .Z(n14532) );
  AND U16708 ( .A(n14533), .B(n14532), .Z(n14669) );
  XOR U16709 ( .A(n14668), .B(n14669), .Z(n14670) );
  NAND U16710 ( .A(n14535), .B(n14534), .Z(n14539) );
  NAND U16711 ( .A(n14537), .B(n14536), .Z(n14538) );
  AND U16712 ( .A(n14539), .B(n14538), .Z(n14671) );
  XOR U16713 ( .A(n14670), .B(n14671), .Z(n14596) );
  XOR U16714 ( .A(n14597), .B(n14596), .Z(n14599) );
  AND U16715 ( .A(x[488]), .B(y[7820]), .Z(n14868) );
  NAND U16716 ( .A(n14868), .B(n14540), .Z(n14544) );
  NANDN U16717 ( .A(n14542), .B(n14541), .Z(n14543) );
  NAND U16718 ( .A(n14544), .B(n14543), .Z(n14681) );
  NAND U16719 ( .A(x[489]), .B(y[7824]), .Z(n15491) );
  NANDN U16720 ( .A(n15491), .B(n14626), .Z(n14548) );
  NAND U16721 ( .A(n14546), .B(n14545), .Z(n14547) );
  NAND U16722 ( .A(n14548), .B(n14547), .Z(n14680) );
  XOR U16723 ( .A(n14681), .B(n14680), .Z(n14683) );
  NAND U16724 ( .A(x[490]), .B(y[7823]), .Z(n15492) );
  NANDN U16725 ( .A(n15492), .B(n14549), .Z(n14553) );
  NANDN U16726 ( .A(n14551), .B(n14550), .Z(n14552) );
  NAND U16727 ( .A(n14553), .B(n14552), .Z(n14658) );
  AND U16728 ( .A(x[480]), .B(y[7826]), .Z(n14632) );
  AND U16729 ( .A(x[498]), .B(y[7808]), .Z(n14631) );
  XOR U16730 ( .A(n14632), .B(n14631), .Z(n14634) );
  AND U16731 ( .A(x[497]), .B(y[7809]), .Z(n14653) );
  XOR U16732 ( .A(n14653), .B(o[146]), .Z(n14633) );
  XOR U16733 ( .A(n14634), .B(n14633), .Z(n14657) );
  AND U16734 ( .A(y[7813]), .B(x[493]), .Z(n14555) );
  NAND U16735 ( .A(y[7823]), .B(x[483]), .Z(n14554) );
  XNOR U16736 ( .A(n14555), .B(n14554), .Z(n14640) );
  AND U16737 ( .A(x[492]), .B(y[7814]), .Z(n14639) );
  XOR U16738 ( .A(n14640), .B(n14639), .Z(n14656) );
  XOR U16739 ( .A(n14657), .B(n14656), .Z(n14659) );
  XOR U16740 ( .A(n14658), .B(n14659), .Z(n14682) );
  XNOR U16741 ( .A(n14683), .B(n14682), .Z(n14603) );
  NANDN U16742 ( .A(n14557), .B(n14556), .Z(n14561) );
  NAND U16743 ( .A(n14559), .B(n14558), .Z(n14560) );
  AND U16744 ( .A(n14561), .B(n14560), .Z(n14602) );
  XOR U16745 ( .A(n14603), .B(n14602), .Z(n14604) );
  NAND U16746 ( .A(n14563), .B(n14562), .Z(n14567) );
  NAND U16747 ( .A(n14565), .B(n14564), .Z(n14566) );
  AND U16748 ( .A(n14567), .B(n14566), .Z(n14605) );
  XOR U16749 ( .A(n14604), .B(n14605), .Z(n14598) );
  XNOR U16750 ( .A(n14599), .B(n14598), .Z(n14593) );
  NAND U16751 ( .A(n14569), .B(n14568), .Z(n14573) );
  NAND U16752 ( .A(n14571), .B(n14570), .Z(n14572) );
  NAND U16753 ( .A(n14573), .B(n14572), .Z(n14591) );
  NAND U16754 ( .A(n14575), .B(n14574), .Z(n14579) );
  NAND U16755 ( .A(n14577), .B(n14576), .Z(n14578) );
  NAND U16756 ( .A(n14579), .B(n14578), .Z(n14590) );
  XOR U16757 ( .A(n14591), .B(n14590), .Z(n14592) );
  XOR U16758 ( .A(n14593), .B(n14592), .Z(n14692) );
  XOR U16759 ( .A(n14693), .B(n14692), .Z(n14694) );
  XOR U16760 ( .A(n14695), .B(n14694), .Z(n14698) );
  OR U16761 ( .A(n14584), .B(n14583), .Z(n14588) );
  NANDN U16762 ( .A(n14586), .B(n14585), .Z(n14587) );
  NAND U16763 ( .A(n14588), .B(n14587), .Z(n14699) );
  XOR U16764 ( .A(n14700), .B(n14699), .Z(n14589) );
  XNOR U16765 ( .A(n14698), .B(n14589), .Z(N307) );
  NAND U16766 ( .A(n14591), .B(n14590), .Z(n14595) );
  NAND U16767 ( .A(n14593), .B(n14592), .Z(n14594) );
  AND U16768 ( .A(n14595), .B(n14594), .Z(n14815) );
  NAND U16769 ( .A(n14597), .B(n14596), .Z(n14601) );
  NAND U16770 ( .A(n14599), .B(n14598), .Z(n14600) );
  AND U16771 ( .A(n14601), .B(n14600), .Z(n14813) );
  NAND U16772 ( .A(n14603), .B(n14602), .Z(n14607) );
  NAND U16773 ( .A(n14605), .B(n14604), .Z(n14606) );
  NAND U16774 ( .A(n14607), .B(n14606), .Z(n14704) );
  AND U16775 ( .A(x[486]), .B(y[7821]), .Z(n14609) );
  NAND U16776 ( .A(n14609), .B(n14608), .Z(n14613) );
  NAND U16777 ( .A(n14611), .B(n14610), .Z(n14612) );
  NAND U16778 ( .A(n14613), .B(n14612), .Z(n14793) );
  AND U16779 ( .A(x[496]), .B(y[7815]), .Z(n15139) );
  NAND U16780 ( .A(n15139), .B(n14979), .Z(n14617) );
  NAND U16781 ( .A(n14615), .B(n14614), .Z(n14616) );
  NAND U16782 ( .A(n14617), .B(n14616), .Z(n14791) );
  AND U16783 ( .A(x[495]), .B(y[7817]), .Z(n15418) );
  NAND U16784 ( .A(n15418), .B(n14720), .Z(n14621) );
  NAND U16785 ( .A(n14619), .B(n14618), .Z(n14620) );
  NAND U16786 ( .A(n14621), .B(n14620), .Z(n14710) );
  AND U16787 ( .A(y[7826]), .B(x[481]), .Z(n14623) );
  NAND U16788 ( .A(y[7819]), .B(x[488]), .Z(n14622) );
  XNOR U16789 ( .A(n14623), .B(n14622), .Z(n14770) );
  XNOR U16790 ( .A(n14770), .B(n14771), .Z(n14709) );
  AND U16791 ( .A(y[7814]), .B(x[493]), .Z(n14625) );
  NAND U16792 ( .A(y[7825]), .B(x[482]), .Z(n14624) );
  XNOR U16793 ( .A(n14625), .B(n14624), .Z(n14727) );
  XOR U16794 ( .A(n14727), .B(n14726), .Z(n14708) );
  XOR U16795 ( .A(n14709), .B(n14708), .Z(n14711) );
  XOR U16796 ( .A(n14710), .B(n14711), .Z(n14792) );
  XOR U16797 ( .A(n14791), .B(n14792), .Z(n14794) );
  XOR U16798 ( .A(n14793), .B(n14794), .Z(n14703) );
  AND U16799 ( .A(x[490]), .B(y[7825]), .Z(n15799) );
  IV U16800 ( .A(n15799), .Z(n15672) );
  NANDN U16801 ( .A(n15672), .B(n14626), .Z(n14630) );
  NAND U16802 ( .A(n14628), .B(n14627), .Z(n14629) );
  NAND U16803 ( .A(n14630), .B(n14629), .Z(n14749) );
  NAND U16804 ( .A(n14632), .B(n14631), .Z(n14636) );
  NAND U16805 ( .A(n14634), .B(n14633), .Z(n14635) );
  NAND U16806 ( .A(n14636), .B(n14635), .Z(n14747) );
  AND U16807 ( .A(y[7811]), .B(x[496]), .Z(n15359) );
  NAND U16808 ( .A(y[7818]), .B(x[489]), .Z(n14637) );
  XNOR U16809 ( .A(n15359), .B(n14637), .Z(n14721) );
  NAND U16810 ( .A(x[495]), .B(y[7812]), .Z(n14722) );
  XNOR U16811 ( .A(n14721), .B(n14722), .Z(n14748) );
  XOR U16812 ( .A(n14747), .B(n14748), .Z(n14750) );
  XOR U16813 ( .A(n14749), .B(n14750), .Z(n14788) );
  AND U16814 ( .A(x[493]), .B(y[7823]), .Z(n15966) );
  NANDN U16815 ( .A(n14638), .B(n15966), .Z(n14642) );
  NAND U16816 ( .A(n14640), .B(n14639), .Z(n14641) );
  NAND U16817 ( .A(n14642), .B(n14641), .Z(n14743) );
  AND U16818 ( .A(y[7817]), .B(x[490]), .Z(n14644) );
  NAND U16819 ( .A(y[7810]), .B(x[497]), .Z(n14643) );
  XNOR U16820 ( .A(n14644), .B(n14643), .Z(n14775) );
  NAND U16821 ( .A(x[498]), .B(y[7809]), .Z(n14740) );
  XOR U16822 ( .A(o[147]), .B(n14740), .Z(n14776) );
  XNOR U16823 ( .A(n14775), .B(n14776), .Z(n14742) );
  NAND U16824 ( .A(y[7824]), .B(x[483]), .Z(n14645) );
  XNOR U16825 ( .A(n14646), .B(n14645), .Z(n14735) );
  XOR U16826 ( .A(n14735), .B(n14734), .Z(n14741) );
  XOR U16827 ( .A(n14742), .B(n14741), .Z(n14744) );
  XOR U16828 ( .A(n14743), .B(n14744), .Z(n14786) );
  NAND U16829 ( .A(n14648), .B(n14647), .Z(n14652) );
  NAND U16830 ( .A(n14650), .B(n14649), .Z(n14651) );
  NAND U16831 ( .A(n14652), .B(n14651), .Z(n14716) );
  AND U16832 ( .A(x[480]), .B(y[7827]), .Z(n14757) );
  NAND U16833 ( .A(x[499]), .B(y[7808]), .Z(n14758) );
  XNOR U16834 ( .A(n14757), .B(n14758), .Z(n14759) );
  NAND U16835 ( .A(n14653), .B(o[146]), .Z(n14760) );
  XNOR U16836 ( .A(n14759), .B(n14760), .Z(n14715) );
  AND U16837 ( .A(x[484]), .B(y[7823]), .Z(n14882) );
  AND U16838 ( .A(y[7822]), .B(x[485]), .Z(n14655) );
  NAND U16839 ( .A(y[7821]), .B(x[486]), .Z(n14654) );
  XOR U16840 ( .A(n14655), .B(n14654), .Z(n14754) );
  XNOR U16841 ( .A(n14882), .B(n14754), .Z(n14714) );
  XOR U16842 ( .A(n14715), .B(n14714), .Z(n14717) );
  XNOR U16843 ( .A(n14716), .B(n14717), .Z(n14785) );
  NAND U16844 ( .A(n14657), .B(n14656), .Z(n14661) );
  NAND U16845 ( .A(n14659), .B(n14658), .Z(n14660) );
  NAND U16846 ( .A(n14661), .B(n14660), .Z(n14780) );
  NAND U16847 ( .A(n14663), .B(n14662), .Z(n14667) );
  NAND U16848 ( .A(n14665), .B(n14664), .Z(n14666) );
  NAND U16849 ( .A(n14667), .B(n14666), .Z(n14779) );
  XOR U16850 ( .A(n14780), .B(n14779), .Z(n14781) );
  XNOR U16851 ( .A(n14782), .B(n14781), .Z(n14702) );
  XOR U16852 ( .A(n14704), .B(n14705), .Z(n14805) );
  NAND U16853 ( .A(n14669), .B(n14668), .Z(n14673) );
  NAND U16854 ( .A(n14671), .B(n14670), .Z(n14672) );
  AND U16855 ( .A(n14673), .B(n14672), .Z(n14804) );
  NAND U16856 ( .A(n14675), .B(n14674), .Z(n14679) );
  NAND U16857 ( .A(n14677), .B(n14676), .Z(n14678) );
  AND U16858 ( .A(n14679), .B(n14678), .Z(n14800) );
  NAND U16859 ( .A(n14681), .B(n14680), .Z(n14685) );
  NAND U16860 ( .A(n14683), .B(n14682), .Z(n14684) );
  AND U16861 ( .A(n14685), .B(n14684), .Z(n14798) );
  NANDN U16862 ( .A(n14687), .B(n14686), .Z(n14691) );
  NAND U16863 ( .A(n14689), .B(n14688), .Z(n14690) );
  NAND U16864 ( .A(n14691), .B(n14690), .Z(n14797) );
  XOR U16865 ( .A(n14804), .B(n14803), .Z(n14806) );
  XOR U16866 ( .A(n14805), .B(n14806), .Z(n14812) );
  XOR U16867 ( .A(n14813), .B(n14812), .Z(n14814) );
  XOR U16868 ( .A(n14815), .B(n14814), .Z(n14811) );
  NAND U16869 ( .A(n14693), .B(n14692), .Z(n14697) );
  NAND U16870 ( .A(n14695), .B(n14694), .Z(n14696) );
  NAND U16871 ( .A(n14697), .B(n14696), .Z(n14810) );
  XOR U16872 ( .A(n14810), .B(n14809), .Z(n14701) );
  XNOR U16873 ( .A(n14811), .B(n14701), .Z(N308) );
  NANDN U16874 ( .A(n14703), .B(n14702), .Z(n14707) );
  NANDN U16875 ( .A(n14705), .B(n14704), .Z(n14706) );
  AND U16876 ( .A(n14707), .B(n14706), .Z(n14916) );
  NAND U16877 ( .A(n14709), .B(n14708), .Z(n14713) );
  NAND U16878 ( .A(n14711), .B(n14710), .Z(n14712) );
  NAND U16879 ( .A(n14713), .B(n14712), .Z(n14820) );
  NAND U16880 ( .A(n14715), .B(n14714), .Z(n14719) );
  NAND U16881 ( .A(n14717), .B(n14716), .Z(n14718) );
  NAND U16882 ( .A(n14719), .B(n14718), .Z(n14819) );
  XOR U16883 ( .A(n14820), .B(n14819), .Z(n14822) );
  AND U16884 ( .A(x[496]), .B(y[7818]), .Z(n15634) );
  NAND U16885 ( .A(n15634), .B(n14720), .Z(n14724) );
  NANDN U16886 ( .A(n14722), .B(n14721), .Z(n14723) );
  AND U16887 ( .A(n14724), .B(n14723), .Z(n14857) );
  AND U16888 ( .A(x[493]), .B(y[7825]), .Z(n16189) );
  NAND U16889 ( .A(n16189), .B(n14725), .Z(n14729) );
  NAND U16890 ( .A(n14727), .B(n14726), .Z(n14728) );
  AND U16891 ( .A(n14729), .B(n14728), .Z(n14900) );
  AND U16892 ( .A(y[7812]), .B(x[496]), .Z(n14731) );
  NAND U16893 ( .A(y[7818]), .B(x[490]), .Z(n14730) );
  XNOR U16894 ( .A(n14731), .B(n14730), .Z(n14863) );
  NAND U16895 ( .A(x[482]), .B(y[7826]), .Z(n14864) );
  XNOR U16896 ( .A(n14863), .B(n14864), .Z(n14897) );
  NAND U16897 ( .A(y[7819]), .B(x[489]), .Z(n14732) );
  XNOR U16898 ( .A(n14733), .B(n14732), .Z(n14845) );
  NAND U16899 ( .A(x[494]), .B(y[7814]), .Z(n14846) );
  XOR U16900 ( .A(n14845), .B(n14846), .Z(n14898) );
  XNOR U16901 ( .A(n14897), .B(n14898), .Z(n14899) );
  XNOR U16902 ( .A(n14900), .B(n14899), .Z(n14856) );
  XNOR U16903 ( .A(n14857), .B(n14856), .Z(n14859) );
  NAND U16904 ( .A(x[491]), .B(y[7824]), .Z(n15800) );
  NANDN U16905 ( .A(n15800), .B(n15006), .Z(n14737) );
  NAND U16906 ( .A(n14735), .B(n14734), .Z(n14736) );
  AND U16907 ( .A(n14737), .B(n14736), .Z(n14906) );
  AND U16908 ( .A(y[7817]), .B(x[491]), .Z(n14739) );
  NAND U16909 ( .A(y[7827]), .B(x[481]), .Z(n14738) );
  XNOR U16910 ( .A(n14739), .B(n14738), .Z(n14843) );
  NAND U16911 ( .A(x[499]), .B(y[7809]), .Z(n14849) );
  XOR U16912 ( .A(n14843), .B(n14842), .Z(n14904) );
  AND U16913 ( .A(x[480]), .B(y[7828]), .Z(n14887) );
  NAND U16914 ( .A(x[500]), .B(y[7808]), .Z(n14888) );
  XNOR U16915 ( .A(n14887), .B(n14888), .Z(n14890) );
  ANDN U16916 ( .B(o[147]), .A(n14740), .Z(n14889) );
  XOR U16917 ( .A(n14890), .B(n14889), .Z(n14903) );
  XOR U16918 ( .A(n14904), .B(n14903), .Z(n14905) );
  XNOR U16919 ( .A(n14906), .B(n14905), .Z(n14858) );
  XOR U16920 ( .A(n14859), .B(n14858), .Z(n14821) );
  XNOR U16921 ( .A(n14822), .B(n14821), .Z(n14910) );
  NAND U16922 ( .A(n14742), .B(n14741), .Z(n14746) );
  NAND U16923 ( .A(n14744), .B(n14743), .Z(n14745) );
  AND U16924 ( .A(n14746), .B(n14745), .Z(n14908) );
  NAND U16925 ( .A(n14748), .B(n14747), .Z(n14752) );
  NAND U16926 ( .A(n14750), .B(n14749), .Z(n14751) );
  AND U16927 ( .A(n14752), .B(n14751), .Z(n14828) );
  AND U16928 ( .A(x[486]), .B(y[7822]), .Z(n14851) );
  NAND U16929 ( .A(n14851), .B(n14753), .Z(n14756) );
  NANDN U16930 ( .A(n14754), .B(n14882), .Z(n14755) );
  AND U16931 ( .A(n14756), .B(n14755), .Z(n14834) );
  NANDN U16932 ( .A(n14758), .B(n14757), .Z(n14762) );
  NANDN U16933 ( .A(n14760), .B(n14759), .Z(n14761) );
  AND U16934 ( .A(n14762), .B(n14761), .Z(n14832) );
  AND U16935 ( .A(y[7810]), .B(x[498]), .Z(n14764) );
  NAND U16936 ( .A(y[7816]), .B(x[492]), .Z(n14763) );
  XNOR U16937 ( .A(n14764), .B(n14763), .Z(n14838) );
  NAND U16938 ( .A(x[497]), .B(y[7811]), .Z(n14839) );
  XNOR U16939 ( .A(n14838), .B(n14839), .Z(n14831) );
  XNOR U16940 ( .A(n14832), .B(n14831), .Z(n14833) );
  XOR U16941 ( .A(n14834), .B(n14833), .Z(n14826) );
  AND U16942 ( .A(y[7815]), .B(x[493]), .Z(n14766) );
  NAND U16943 ( .A(y[7825]), .B(x[483]), .Z(n14765) );
  XNOR U16944 ( .A(n14766), .B(n14765), .Z(n14869) );
  XOR U16945 ( .A(n14869), .B(n14868), .Z(n14852) );
  AND U16946 ( .A(y[7823]), .B(x[485]), .Z(n14768) );
  NAND U16947 ( .A(y[7824]), .B(x[484]), .Z(n14767) );
  XNOR U16948 ( .A(n14768), .B(n14767), .Z(n14884) );
  AND U16949 ( .A(x[487]), .B(y[7821]), .Z(n14883) );
  XNOR U16950 ( .A(n14884), .B(n14883), .Z(n14850) );
  XOR U16951 ( .A(n14851), .B(n14850), .Z(n14853) );
  XOR U16952 ( .A(n14852), .B(n14853), .Z(n14893) );
  AND U16953 ( .A(x[488]), .B(y[7826]), .Z(n15930) );
  AND U16954 ( .A(x[481]), .B(y[7819]), .Z(n14769) );
  NAND U16955 ( .A(n15930), .B(n14769), .Z(n14773) );
  NANDN U16956 ( .A(n14771), .B(n14770), .Z(n14772) );
  AND U16957 ( .A(n14773), .B(n14772), .Z(n14892) );
  NAND U16958 ( .A(x[497]), .B(y[7817]), .Z(n15642) );
  NANDN U16959 ( .A(n15642), .B(n14774), .Z(n14778) );
  NANDN U16960 ( .A(n14776), .B(n14775), .Z(n14777) );
  NAND U16961 ( .A(n14778), .B(n14777), .Z(n14891) );
  XOR U16962 ( .A(n14892), .B(n14891), .Z(n14894) );
  XNOR U16963 ( .A(n14893), .B(n14894), .Z(n14825) );
  XOR U16964 ( .A(n14826), .B(n14825), .Z(n14827) );
  XOR U16965 ( .A(n14828), .B(n14827), .Z(n14907) );
  XOR U16966 ( .A(n14908), .B(n14907), .Z(n14909) );
  XOR U16967 ( .A(n14910), .B(n14909), .Z(n14914) );
  NAND U16968 ( .A(n14780), .B(n14779), .Z(n14784) );
  NAND U16969 ( .A(n14782), .B(n14781), .Z(n14783) );
  AND U16970 ( .A(n14784), .B(n14783), .Z(n14922) );
  NANDN U16971 ( .A(n14786), .B(n14785), .Z(n14790) );
  NANDN U16972 ( .A(n14788), .B(n14787), .Z(n14789) );
  NAND U16973 ( .A(n14790), .B(n14789), .Z(n14919) );
  NAND U16974 ( .A(n14792), .B(n14791), .Z(n14796) );
  NAND U16975 ( .A(n14794), .B(n14793), .Z(n14795) );
  AND U16976 ( .A(n14796), .B(n14795), .Z(n14920) );
  XOR U16977 ( .A(n14919), .B(n14920), .Z(n14921) );
  XNOR U16978 ( .A(n14922), .B(n14921), .Z(n14913) );
  XOR U16979 ( .A(n14916), .B(n14915), .Z(n14935) );
  NANDN U16980 ( .A(n14798), .B(n14797), .Z(n14802) );
  NANDN U16981 ( .A(n14800), .B(n14799), .Z(n14801) );
  AND U16982 ( .A(n14802), .B(n14801), .Z(n14932) );
  NAND U16983 ( .A(n14804), .B(n14803), .Z(n14808) );
  NAND U16984 ( .A(n14806), .B(n14805), .Z(n14807) );
  AND U16985 ( .A(n14808), .B(n14807), .Z(n14933) );
  XOR U16986 ( .A(n14932), .B(n14933), .Z(n14934) );
  XOR U16987 ( .A(n14935), .B(n14934), .Z(n14928) );
  NAND U16988 ( .A(n14813), .B(n14812), .Z(n14817) );
  NANDN U16989 ( .A(n14815), .B(n14814), .Z(n14816) );
  AND U16990 ( .A(n14817), .B(n14816), .Z(n14927) );
  IV U16991 ( .A(n14927), .Z(n14925) );
  XOR U16992 ( .A(n14926), .B(n14925), .Z(n14818) );
  XNOR U16993 ( .A(n14928), .B(n14818), .Z(N309) );
  NAND U16994 ( .A(n14820), .B(n14819), .Z(n14824) );
  NAND U16995 ( .A(n14822), .B(n14821), .Z(n14823) );
  NAND U16996 ( .A(n14824), .B(n14823), .Z(n14947) );
  NAND U16997 ( .A(n14826), .B(n14825), .Z(n14830) );
  NAND U16998 ( .A(n14828), .B(n14827), .Z(n14829) );
  AND U16999 ( .A(n14830), .B(n14829), .Z(n14946) );
  NANDN U17000 ( .A(n14832), .B(n14831), .Z(n14836) );
  NANDN U17001 ( .A(n14834), .B(n14833), .Z(n14835) );
  AND U17002 ( .A(n14836), .B(n14835), .Z(n15030) );
  AND U17003 ( .A(x[498]), .B(y[7816]), .Z(n15641) );
  NAND U17004 ( .A(n15641), .B(n14837), .Z(n14841) );
  NANDN U17005 ( .A(n14839), .B(n14838), .Z(n14840) );
  AND U17006 ( .A(n14841), .B(n14840), .Z(n15035) );
  AND U17007 ( .A(x[491]), .B(y[7827]), .Z(n16334) );
  XNOR U17008 ( .A(n15035), .B(n15034), .Z(n15036) );
  AND U17009 ( .A(x[495]), .B(y[7819]), .Z(n15629) );
  NAND U17010 ( .A(n15629), .B(n14844), .Z(n14848) );
  NANDN U17011 ( .A(n14846), .B(n14845), .Z(n14847) );
  AND U17012 ( .A(n14848), .B(n14847), .Z(n14993) );
  AND U17013 ( .A(x[480]), .B(y[7829]), .Z(n15012) );
  NAND U17014 ( .A(x[501]), .B(y[7808]), .Z(n15013) );
  ANDN U17015 ( .B(o[148]), .A(n14849), .Z(n15014) );
  XOR U17016 ( .A(n15015), .B(n15014), .Z(n14991) );
  AND U17017 ( .A(x[485]), .B(y[7824]), .Z(n14997) );
  AND U17018 ( .A(x[496]), .B(y[7813]), .Z(n14996) );
  XOR U17019 ( .A(n14997), .B(n14996), .Z(n14999) );
  AND U17020 ( .A(x[495]), .B(y[7814]), .Z(n14998) );
  XOR U17021 ( .A(n14999), .B(n14998), .Z(n14990) );
  XOR U17022 ( .A(n14991), .B(n14990), .Z(n14992) );
  XNOR U17023 ( .A(n15036), .B(n15037), .Z(n15028) );
  NANDN U17024 ( .A(n14851), .B(n14850), .Z(n14855) );
  OR U17025 ( .A(n14853), .B(n14852), .Z(n14854) );
  NAND U17026 ( .A(n14855), .B(n14854), .Z(n15029) );
  XOR U17027 ( .A(n15028), .B(n15029), .Z(n15031) );
  XOR U17028 ( .A(n15030), .B(n15031), .Z(n14945) );
  XOR U17029 ( .A(n14946), .B(n14945), .Z(n14948) );
  XNOR U17030 ( .A(n14947), .B(n14948), .Z(n14942) );
  NANDN U17031 ( .A(n14857), .B(n14856), .Z(n14861) );
  NAND U17032 ( .A(n14859), .B(n14858), .Z(n14860) );
  AND U17033 ( .A(n14861), .B(n14860), .Z(n14954) );
  NAND U17034 ( .A(n15634), .B(n14862), .Z(n14866) );
  NANDN U17035 ( .A(n14864), .B(n14863), .Z(n14865) );
  AND U17036 ( .A(n14866), .B(n14865), .Z(n14962) );
  NAND U17037 ( .A(n14867), .B(n16189), .Z(n14871) );
  NAND U17038 ( .A(n14869), .B(n14868), .Z(n14870) );
  AND U17039 ( .A(n14871), .B(n14870), .Z(n15049) );
  AND U17040 ( .A(y[7810]), .B(x[499]), .Z(n14873) );
  NAND U17041 ( .A(y[7818]), .B(x[491]), .Z(n14872) );
  XNOR U17042 ( .A(n14873), .B(n14872), .Z(n14981) );
  AND U17043 ( .A(x[500]), .B(y[7809]), .Z(n15011) );
  XOR U17044 ( .A(o[149]), .B(n15011), .Z(n14980) );
  XOR U17045 ( .A(n14981), .B(n14980), .Z(n15047) );
  AND U17046 ( .A(y[7811]), .B(x[498]), .Z(n14875) );
  NAND U17047 ( .A(y[7819]), .B(x[490]), .Z(n14874) );
  XNOR U17048 ( .A(n14875), .B(n14874), .Z(n15019) );
  NAND U17049 ( .A(x[481]), .B(y[7828]), .Z(n15020) );
  XOR U17050 ( .A(n15047), .B(n15046), .Z(n15048) );
  XNOR U17051 ( .A(n15049), .B(n15048), .Z(n14961) );
  XNOR U17052 ( .A(n14962), .B(n14961), .Z(n14963) );
  AND U17053 ( .A(x[487]), .B(y[7822]), .Z(n15208) );
  AND U17054 ( .A(y[7823]), .B(x[486]), .Z(n14877) );
  NAND U17055 ( .A(y[7815]), .B(x[494]), .Z(n14876) );
  XNOR U17056 ( .A(n14877), .B(n14876), .Z(n15023) );
  XOR U17057 ( .A(n15208), .B(n15023), .Z(n14970) );
  AND U17058 ( .A(x[489]), .B(y[7820]), .Z(n14968) );
  NAND U17059 ( .A(x[488]), .B(y[7821]), .Z(n14967) );
  AND U17060 ( .A(y[7817]), .B(x[492]), .Z(n14879) );
  NAND U17061 ( .A(y[7812]), .B(x[497]), .Z(n14878) );
  XNOR U17062 ( .A(n14879), .B(n14878), .Z(n14973) );
  NAND U17063 ( .A(x[482]), .B(y[7827]), .Z(n14974) );
  AND U17064 ( .A(y[7816]), .B(x[493]), .Z(n14881) );
  NAND U17065 ( .A(y[7826]), .B(x[483]), .Z(n14880) );
  XNOR U17066 ( .A(n14881), .B(n14880), .Z(n15007) );
  NAND U17067 ( .A(x[484]), .B(y[7825]), .Z(n15008) );
  XOR U17068 ( .A(n14985), .B(n14984), .Z(n14987) );
  XOR U17069 ( .A(n14986), .B(n14987), .Z(n15042) );
  NAND U17070 ( .A(n14997), .B(n14882), .Z(n14886) );
  NAND U17071 ( .A(n14884), .B(n14883), .Z(n14885) );
  AND U17072 ( .A(n14886), .B(n14885), .Z(n15041) );
  XOR U17073 ( .A(n15041), .B(n15040), .Z(n15043) );
  XOR U17074 ( .A(n15042), .B(n15043), .Z(n14964) );
  XNOR U17075 ( .A(n14963), .B(n14964), .Z(n14952) );
  NANDN U17076 ( .A(n14892), .B(n14891), .Z(n14896) );
  OR U17077 ( .A(n14894), .B(n14893), .Z(n14895) );
  NAND U17078 ( .A(n14896), .B(n14895), .Z(n14957) );
  NANDN U17079 ( .A(n14898), .B(n14897), .Z(n14902) );
  NANDN U17080 ( .A(n14900), .B(n14899), .Z(n14901) );
  NAND U17081 ( .A(n14902), .B(n14901), .Z(n14956) );
  XOR U17082 ( .A(n14956), .B(n14955), .Z(n14958) );
  XOR U17083 ( .A(n14957), .B(n14958), .Z(n14951) );
  XOR U17084 ( .A(n14952), .B(n14951), .Z(n14953) );
  XOR U17085 ( .A(n14954), .B(n14953), .Z(n14940) );
  NAND U17086 ( .A(n14908), .B(n14907), .Z(n14912) );
  NAND U17087 ( .A(n14910), .B(n14909), .Z(n14911) );
  NAND U17088 ( .A(n14912), .B(n14911), .Z(n14939) );
  XOR U17089 ( .A(n14940), .B(n14939), .Z(n14941) );
  XNOR U17090 ( .A(n14942), .B(n14941), .Z(n15052) );
  NANDN U17091 ( .A(n14914), .B(n14913), .Z(n14918) );
  NAND U17092 ( .A(n14916), .B(n14915), .Z(n14917) );
  NAND U17093 ( .A(n14918), .B(n14917), .Z(n15050) );
  NAND U17094 ( .A(n14920), .B(n14919), .Z(n14924) );
  NAND U17095 ( .A(n14922), .B(n14921), .Z(n14923) );
  AND U17096 ( .A(n14924), .B(n14923), .Z(n15051) );
  XNOR U17097 ( .A(n15050), .B(n15051), .Z(n15053) );
  XOR U17098 ( .A(n15052), .B(n15053), .Z(n15058) );
  NANDN U17099 ( .A(n14925), .B(n14926), .Z(n14931) );
  NOR U17100 ( .A(n14927), .B(n14926), .Z(n14929) );
  OR U17101 ( .A(n14929), .B(n14928), .Z(n14930) );
  AND U17102 ( .A(n14931), .B(n14930), .Z(n15056) );
  NAND U17103 ( .A(n14933), .B(n14932), .Z(n14937) );
  NANDN U17104 ( .A(n14935), .B(n14934), .Z(n14936) );
  AND U17105 ( .A(n14937), .B(n14936), .Z(n15057) );
  XOR U17106 ( .A(n15056), .B(n15057), .Z(n14938) );
  XNOR U17107 ( .A(n15058), .B(n14938), .Z(N310) );
  NAND U17108 ( .A(n14940), .B(n14939), .Z(n14944) );
  NAND U17109 ( .A(n14942), .B(n14941), .Z(n14943) );
  AND U17110 ( .A(n14944), .B(n14943), .Z(n15062) );
  NAND U17111 ( .A(n14946), .B(n14945), .Z(n14950) );
  NAND U17112 ( .A(n14948), .B(n14947), .Z(n14949) );
  NAND U17113 ( .A(n14950), .B(n14949), .Z(n15060) );
  NAND U17114 ( .A(n14956), .B(n14955), .Z(n14960) );
  NAND U17115 ( .A(n14958), .B(n14957), .Z(n14959) );
  NAND U17116 ( .A(n14960), .B(n14959), .Z(n15069) );
  XNOR U17117 ( .A(n15070), .B(n15069), .Z(n15072) );
  NANDN U17118 ( .A(n14962), .B(n14961), .Z(n14966) );
  NANDN U17119 ( .A(n14964), .B(n14963), .Z(n14965) );
  AND U17120 ( .A(n14966), .B(n14965), .Z(n15178) );
  NANDN U17121 ( .A(n14968), .B(n14967), .Z(n14972) );
  NANDN U17122 ( .A(n14970), .B(n14969), .Z(n14971) );
  AND U17123 ( .A(n14972), .B(n14971), .Z(n15172) );
  NANDN U17124 ( .A(n15642), .B(n15123), .Z(n14976) );
  NANDN U17125 ( .A(n14974), .B(n14973), .Z(n14975) );
  NAND U17126 ( .A(n14976), .B(n14975), .Z(n15101) );
  AND U17127 ( .A(x[485]), .B(y[7825]), .Z(n15145) );
  AND U17128 ( .A(x[497]), .B(y[7813]), .Z(n15146) );
  XOR U17129 ( .A(n15145), .B(n15146), .Z(n15147) );
  AND U17130 ( .A(x[496]), .B(y[7814]), .Z(n15148) );
  XOR U17131 ( .A(n15147), .B(n15148), .Z(n15100) );
  AND U17132 ( .A(y[7812]), .B(x[498]), .Z(n14978) );
  NAND U17133 ( .A(y[7818]), .B(x[492]), .Z(n14977) );
  XNOR U17134 ( .A(n14978), .B(n14977), .Z(n15124) );
  AND U17135 ( .A(x[484]), .B(y[7826]), .Z(n15125) );
  XOR U17136 ( .A(n15124), .B(n15125), .Z(n15099) );
  XNOR U17137 ( .A(n15100), .B(n15099), .Z(n15102) );
  XOR U17138 ( .A(n15101), .B(n15102), .Z(n15170) );
  AND U17139 ( .A(x[499]), .B(y[7818]), .Z(n16101) );
  NAND U17140 ( .A(n16101), .B(n14979), .Z(n14983) );
  NAND U17141 ( .A(n14981), .B(n14980), .Z(n14982) );
  AND U17142 ( .A(n14983), .B(n14982), .Z(n15169) );
  XOR U17143 ( .A(n15170), .B(n15169), .Z(n15171) );
  XNOR U17144 ( .A(n15172), .B(n15171), .Z(n15176) );
  NAND U17145 ( .A(n14985), .B(n14984), .Z(n14989) );
  NAND U17146 ( .A(n14987), .B(n14986), .Z(n14988) );
  AND U17147 ( .A(n14989), .B(n14988), .Z(n15158) );
  NAND U17148 ( .A(n14991), .B(n14990), .Z(n14995) );
  NANDN U17149 ( .A(n14993), .B(n14992), .Z(n14994) );
  NAND U17150 ( .A(n14995), .B(n14994), .Z(n15157) );
  XNOR U17151 ( .A(n15158), .B(n15157), .Z(n15159) );
  NAND U17152 ( .A(n14997), .B(n14996), .Z(n15001) );
  AND U17153 ( .A(n14999), .B(n14998), .Z(n15000) );
  ANDN U17154 ( .B(n15001), .A(n15000), .Z(n15122) );
  AND U17155 ( .A(y[7817]), .B(x[493]), .Z(n15003) );
  NAND U17156 ( .A(y[7810]), .B(x[500]), .Z(n15002) );
  XNOR U17157 ( .A(n15003), .B(n15002), .Z(n15141) );
  AND U17158 ( .A(x[482]), .B(y[7828]), .Z(n15142) );
  XOR U17159 ( .A(n15141), .B(n15142), .Z(n15120) );
  AND U17160 ( .A(y[7824]), .B(x[486]), .Z(n15005) );
  NAND U17161 ( .A(y[7815]), .B(x[495]), .Z(n15004) );
  XNOR U17162 ( .A(n15005), .B(n15004), .Z(n15153) );
  XOR U17163 ( .A(n15120), .B(n15119), .Z(n15121) );
  XNOR U17164 ( .A(n15122), .B(n15121), .Z(n15163) );
  AND U17165 ( .A(x[493]), .B(y[7826]), .Z(n16332) );
  NAND U17166 ( .A(n15006), .B(n16332), .Z(n15010) );
  NANDN U17167 ( .A(n15008), .B(n15007), .Z(n15009) );
  AND U17168 ( .A(n15010), .B(n15009), .Z(n15090) );
  AND U17169 ( .A(x[481]), .B(y[7829]), .Z(n15113) );
  XOR U17170 ( .A(n15114), .B(n15113), .Z(n15112) );
  AND U17171 ( .A(o[149]), .B(n15011), .Z(n15111) );
  XOR U17172 ( .A(n15112), .B(n15111), .Z(n15087) );
  AND U17173 ( .A(x[494]), .B(y[7816]), .Z(n15105) );
  AND U17174 ( .A(x[483]), .B(y[7827]), .Z(n15106) );
  XOR U17175 ( .A(n15105), .B(n15106), .Z(n15107) );
  AND U17176 ( .A(x[499]), .B(y[7811]), .Z(n15108) );
  XNOR U17177 ( .A(n15107), .B(n15108), .Z(n15088) );
  XNOR U17178 ( .A(n15087), .B(n15088), .Z(n15089) );
  XOR U17179 ( .A(n15090), .B(n15089), .Z(n15164) );
  NANDN U17180 ( .A(n15013), .B(n15012), .Z(n15017) );
  NAND U17181 ( .A(n15015), .B(n15014), .Z(n15016) );
  AND U17182 ( .A(n15017), .B(n15016), .Z(n15082) );
  AND U17183 ( .A(x[498]), .B(y[7819]), .Z(n16103) );
  NAND U17184 ( .A(n16103), .B(n15018), .Z(n15022) );
  NANDN U17185 ( .A(n15020), .B(n15019), .Z(n15021) );
  NAND U17186 ( .A(n15022), .B(n15021), .Z(n15081) );
  XNOR U17187 ( .A(n15082), .B(n15081), .Z(n15083) );
  AND U17188 ( .A(x[494]), .B(y[7823]), .Z(n16136) );
  NAND U17189 ( .A(n15152), .B(n16136), .Z(n15025) );
  NAND U17190 ( .A(n15208), .B(n15023), .Z(n15024) );
  AND U17191 ( .A(n15025), .B(n15024), .Z(n15096) );
  AND U17192 ( .A(x[480]), .B(y[7830]), .Z(n15128) );
  AND U17193 ( .A(x[502]), .B(y[7808]), .Z(n15129) );
  XOR U17194 ( .A(n15128), .B(n15129), .Z(n15131) );
  AND U17195 ( .A(x[501]), .B(y[7809]), .Z(n15151) );
  XOR U17196 ( .A(o[150]), .B(n15151), .Z(n15130) );
  XOR U17197 ( .A(n15131), .B(n15130), .Z(n15094) );
  AND U17198 ( .A(y[7823]), .B(x[487]), .Z(n15027) );
  NAND U17199 ( .A(y[7822]), .B(x[488]), .Z(n15026) );
  XNOR U17200 ( .A(n15027), .B(n15026), .Z(n15134) );
  XOR U17201 ( .A(n15094), .B(n15093), .Z(n15095) );
  XNOR U17202 ( .A(n15083), .B(n15084), .Z(n15165) );
  XNOR U17203 ( .A(n15166), .B(n15165), .Z(n15160) );
  XNOR U17204 ( .A(n15159), .B(n15160), .Z(n15175) );
  XNOR U17205 ( .A(n15176), .B(n15175), .Z(n15177) );
  XNOR U17206 ( .A(n15178), .B(n15177), .Z(n15183) );
  NANDN U17207 ( .A(n15029), .B(n15028), .Z(n15033) );
  OR U17208 ( .A(n15031), .B(n15030), .Z(n15032) );
  AND U17209 ( .A(n15033), .B(n15032), .Z(n15182) );
  NANDN U17210 ( .A(n15035), .B(n15034), .Z(n15039) );
  NANDN U17211 ( .A(n15037), .B(n15036), .Z(n15038) );
  AND U17212 ( .A(n15039), .B(n15038), .Z(n15078) );
  NANDN U17213 ( .A(n15041), .B(n15040), .Z(n15045) );
  NANDN U17214 ( .A(n15043), .B(n15042), .Z(n15044) );
  AND U17215 ( .A(n15045), .B(n15044), .Z(n15076) );
  XNOR U17216 ( .A(n15076), .B(n15075), .Z(n15077) );
  XNOR U17217 ( .A(n15078), .B(n15077), .Z(n15181) );
  XOR U17218 ( .A(n15182), .B(n15181), .Z(n15184) );
  XNOR U17219 ( .A(n15183), .B(n15184), .Z(n15071) );
  XOR U17220 ( .A(n15072), .B(n15071), .Z(n15061) );
  XOR U17221 ( .A(n15060), .B(n15061), .Z(n15063) );
  XOR U17222 ( .A(n15062), .B(n15063), .Z(n15068) );
  NAND U17223 ( .A(n15051), .B(n15050), .Z(n15055) );
  NANDN U17224 ( .A(n15053), .B(n15052), .Z(n15054) );
  AND U17225 ( .A(n15055), .B(n15054), .Z(n15067) );
  XNOR U17226 ( .A(n15067), .B(n15066), .Z(n15059) );
  XNOR U17227 ( .A(n15068), .B(n15059), .Z(N311) );
  NAND U17228 ( .A(n15061), .B(n15060), .Z(n15065) );
  NAND U17229 ( .A(n15063), .B(n15062), .Z(n15064) );
  NAND U17230 ( .A(n15065), .B(n15064), .Z(n15326) );
  NANDN U17231 ( .A(n15070), .B(n15069), .Z(n15074) );
  NAND U17232 ( .A(n15072), .B(n15071), .Z(n15073) );
  AND U17233 ( .A(n15074), .B(n15073), .Z(n15321) );
  NANDN U17234 ( .A(n15076), .B(n15075), .Z(n15080) );
  NANDN U17235 ( .A(n15078), .B(n15077), .Z(n15079) );
  AND U17236 ( .A(n15080), .B(n15079), .Z(n15304) );
  NANDN U17237 ( .A(n15082), .B(n15081), .Z(n15086) );
  NANDN U17238 ( .A(n15084), .B(n15083), .Z(n15085) );
  AND U17239 ( .A(n15086), .B(n15085), .Z(n15298) );
  NANDN U17240 ( .A(n15088), .B(n15087), .Z(n15092) );
  NANDN U17241 ( .A(n15090), .B(n15089), .Z(n15091) );
  AND U17242 ( .A(n15092), .B(n15091), .Z(n15296) );
  NAND U17243 ( .A(n15094), .B(n15093), .Z(n15098) );
  NANDN U17244 ( .A(n15096), .B(n15095), .Z(n15097) );
  NAND U17245 ( .A(n15098), .B(n15097), .Z(n15295) );
  NAND U17246 ( .A(n15100), .B(n15099), .Z(n15104) );
  NANDN U17247 ( .A(n15102), .B(n15101), .Z(n15103) );
  AND U17248 ( .A(n15104), .B(n15103), .Z(n15314) );
  NAND U17249 ( .A(n15106), .B(n15105), .Z(n15110) );
  NAND U17250 ( .A(n15108), .B(n15107), .Z(n15109) );
  NAND U17251 ( .A(n15110), .B(n15109), .Z(n15242) );
  AND U17252 ( .A(n15112), .B(n15111), .Z(n15116) );
  NAND U17253 ( .A(n15114), .B(n15113), .Z(n15115) );
  NANDN U17254 ( .A(n15116), .B(n15115), .Z(n15241) );
  XOR U17255 ( .A(n15242), .B(n15241), .Z(n15244) );
  AND U17256 ( .A(y[7824]), .B(x[487]), .Z(n15118) );
  NAND U17257 ( .A(y[7822]), .B(x[489]), .Z(n15117) );
  XNOR U17258 ( .A(n15118), .B(n15117), .Z(n15209) );
  AND U17259 ( .A(x[490]), .B(y[7821]), .Z(n15248) );
  XOR U17260 ( .A(n15247), .B(n15248), .Z(n15250) );
  AND U17261 ( .A(x[486]), .B(y[7825]), .Z(n15200) );
  AND U17262 ( .A(x[495]), .B(y[7816]), .Z(n15201) );
  XOR U17263 ( .A(n15200), .B(n15201), .Z(n15202) );
  AND U17264 ( .A(x[491]), .B(y[7820]), .Z(n15203) );
  XOR U17265 ( .A(n15202), .B(n15203), .Z(n15249) );
  XOR U17266 ( .A(n15250), .B(n15249), .Z(n15243) );
  XOR U17267 ( .A(n15244), .B(n15243), .Z(n15313) );
  XOR U17268 ( .A(n15316), .B(n15315), .Z(n15302) );
  AND U17269 ( .A(x[498]), .B(y[7818]), .Z(n15957) );
  NAND U17270 ( .A(n15957), .B(n15123), .Z(n15127) );
  NAND U17271 ( .A(n15125), .B(n15124), .Z(n15126) );
  AND U17272 ( .A(n15127), .B(n15126), .Z(n15272) );
  NAND U17273 ( .A(n15129), .B(n15128), .Z(n15133) );
  NAND U17274 ( .A(n15131), .B(n15130), .Z(n15132) );
  NAND U17275 ( .A(n15133), .B(n15132), .Z(n15271) );
  NANDN U17276 ( .A(n15210), .B(n15208), .Z(n15137) );
  NANDN U17277 ( .A(n15135), .B(n15134), .Z(n15136) );
  AND U17278 ( .A(n15137), .B(n15136), .Z(n15286) );
  AND U17279 ( .A(x[480]), .B(y[7831]), .Z(n15219) );
  AND U17280 ( .A(x[503]), .B(y[7808]), .Z(n15220) );
  XOR U17281 ( .A(n15219), .B(n15220), .Z(n15222) );
  AND U17282 ( .A(x[502]), .B(y[7809]), .Z(n15199) );
  XOR U17283 ( .A(o[151]), .B(n15199), .Z(n15221) );
  XOR U17284 ( .A(n15222), .B(n15221), .Z(n15284) );
  NAND U17285 ( .A(y[7811]), .B(x[500]), .Z(n15138) );
  XNOR U17286 ( .A(n15139), .B(n15138), .Z(n15195) );
  AND U17287 ( .A(x[499]), .B(y[7812]), .Z(n15196) );
  XOR U17288 ( .A(n15195), .B(n15196), .Z(n15283) );
  XOR U17289 ( .A(n15284), .B(n15283), .Z(n15285) );
  XOR U17290 ( .A(n15274), .B(n15273), .Z(n15235) );
  XOR U17291 ( .A(n15236), .B(n15235), .Z(n15238) );
  AND U17292 ( .A(x[500]), .B(y[7817]), .Z(n16141) );
  AND U17293 ( .A(x[493]), .B(y[7810]), .Z(n15140) );
  NAND U17294 ( .A(n16141), .B(n15140), .Z(n15144) );
  NAND U17295 ( .A(n15142), .B(n15141), .Z(n15143) );
  NAND U17296 ( .A(n15144), .B(n15143), .Z(n15230) );
  NAND U17297 ( .A(n15146), .B(n15145), .Z(n15150) );
  NAND U17298 ( .A(n15148), .B(n15147), .Z(n15149) );
  AND U17299 ( .A(n15150), .B(n15149), .Z(n15292) );
  AND U17300 ( .A(x[493]), .B(y[7818]), .Z(n15265) );
  AND U17301 ( .A(x[482]), .B(y[7829]), .Z(n15266) );
  XOR U17302 ( .A(n15265), .B(n15266), .Z(n15267) );
  AND U17303 ( .A(x[501]), .B(y[7810]), .Z(n15268) );
  XOR U17304 ( .A(n15267), .B(n15268), .Z(n15290) );
  AND U17305 ( .A(x[492]), .B(y[7819]), .Z(n15213) );
  AND U17306 ( .A(x[481]), .B(y[7830]), .Z(n15214) );
  XOR U17307 ( .A(n15213), .B(n15214), .Z(n15216) );
  AND U17308 ( .A(o[150]), .B(n15151), .Z(n15215) );
  XOR U17309 ( .A(n15216), .B(n15215), .Z(n15289) );
  XOR U17310 ( .A(n15290), .B(n15289), .Z(n15291) );
  XOR U17311 ( .A(n15230), .B(n15229), .Z(n15232) );
  AND U17312 ( .A(x[495]), .B(y[7824]), .Z(n16271) );
  NAND U17313 ( .A(n16271), .B(n15152), .Z(n15156) );
  NANDN U17314 ( .A(n15154), .B(n15153), .Z(n15155) );
  AND U17315 ( .A(n15156), .B(n15155), .Z(n15280) );
  AND U17316 ( .A(x[494]), .B(y[7817]), .Z(n15259) );
  AND U17317 ( .A(x[483]), .B(y[7828]), .Z(n15260) );
  XOR U17318 ( .A(n15259), .B(n15260), .Z(n15261) );
  AND U17319 ( .A(x[484]), .B(y[7827]), .Z(n15262) );
  XOR U17320 ( .A(n15261), .B(n15262), .Z(n15278) );
  AND U17321 ( .A(x[485]), .B(y[7826]), .Z(n15253) );
  AND U17322 ( .A(x[498]), .B(y[7813]), .Z(n15254) );
  XOR U17323 ( .A(n15253), .B(n15254), .Z(n15255) );
  AND U17324 ( .A(x[497]), .B(y[7814]), .Z(n15256) );
  XOR U17325 ( .A(n15255), .B(n15256), .Z(n15277) );
  XOR U17326 ( .A(n15278), .B(n15277), .Z(n15279) );
  XOR U17327 ( .A(n15232), .B(n15231), .Z(n15237) );
  XOR U17328 ( .A(n15238), .B(n15237), .Z(n15301) );
  XOR U17329 ( .A(n15302), .B(n15301), .Z(n15303) );
  NANDN U17330 ( .A(n15158), .B(n15157), .Z(n15162) );
  NANDN U17331 ( .A(n15160), .B(n15159), .Z(n15161) );
  AND U17332 ( .A(n15162), .B(n15161), .Z(n15310) );
  NANDN U17333 ( .A(n15164), .B(n15163), .Z(n15168) );
  NAND U17334 ( .A(n15166), .B(n15165), .Z(n15167) );
  AND U17335 ( .A(n15168), .B(n15167), .Z(n15308) );
  NAND U17336 ( .A(n15170), .B(n15169), .Z(n15174) );
  NANDN U17337 ( .A(n15172), .B(n15171), .Z(n15173) );
  AND U17338 ( .A(n15174), .B(n15173), .Z(n15307) );
  NANDN U17339 ( .A(n15176), .B(n15175), .Z(n15180) );
  NANDN U17340 ( .A(n15178), .B(n15177), .Z(n15179) );
  AND U17341 ( .A(n15180), .B(n15179), .Z(n15188) );
  NANDN U17342 ( .A(n15182), .B(n15181), .Z(n15186) );
  NANDN U17343 ( .A(n15184), .B(n15183), .Z(n15185) );
  NAND U17344 ( .A(n15186), .B(n15185), .Z(n15320) );
  XOR U17345 ( .A(n15319), .B(n15320), .Z(n15322) );
  XNOR U17346 ( .A(n15321), .B(n15322), .Z(n15327) );
  XOR U17347 ( .A(n15325), .B(n15327), .Z(n15187) );
  XNOR U17348 ( .A(n15326), .B(n15187), .Z(N312) );
  NANDN U17349 ( .A(n15189), .B(n15188), .Z(n15193) );
  NANDN U17350 ( .A(n15191), .B(n15190), .Z(n15192) );
  AND U17351 ( .A(n15193), .B(n15192), .Z(n15464) );
  AND U17352 ( .A(x[500]), .B(y[7815]), .Z(n15194) );
  NAND U17353 ( .A(n15359), .B(n15194), .Z(n15198) );
  NAND U17354 ( .A(n15196), .B(n15195), .Z(n15197) );
  AND U17355 ( .A(n15198), .B(n15197), .Z(n15379) );
  AND U17356 ( .A(x[502]), .B(y[7810]), .Z(n15398) );
  XOR U17357 ( .A(n15399), .B(n15398), .Z(n15401) );
  AND U17358 ( .A(x[482]), .B(y[7830]), .Z(n15400) );
  XOR U17359 ( .A(n15401), .B(n15400), .Z(n15377) );
  AND U17360 ( .A(x[481]), .B(y[7831]), .Z(n15406) );
  XOR U17361 ( .A(n15407), .B(n15406), .Z(n15405) );
  AND U17362 ( .A(o[151]), .B(n15199), .Z(n15404) );
  XOR U17363 ( .A(n15405), .B(n15404), .Z(n15376) );
  XOR U17364 ( .A(n15377), .B(n15376), .Z(n15378) );
  NAND U17365 ( .A(n15201), .B(n15200), .Z(n15205) );
  NAND U17366 ( .A(n15203), .B(n15202), .Z(n15204) );
  AND U17367 ( .A(n15205), .B(n15204), .Z(n15373) );
  AND U17368 ( .A(y[7816]), .B(x[496]), .Z(n15207) );
  NAND U17369 ( .A(y[7811]), .B(x[501]), .Z(n15206) );
  XNOR U17370 ( .A(n15207), .B(n15206), .Z(n15360) );
  NAND U17371 ( .A(x[485]), .B(y[7827]), .Z(n15361) );
  AND U17372 ( .A(x[500]), .B(y[7812]), .Z(n15558) );
  NAND U17373 ( .A(x[486]), .B(y[7826]), .Z(n15722) );
  NAND U17374 ( .A(x[499]), .B(y[7813]), .Z(n15367) );
  XOR U17375 ( .A(n15371), .B(n15370), .Z(n15372) );
  NANDN U17376 ( .A(n15491), .B(n15208), .Z(n15212) );
  NANDN U17377 ( .A(n15210), .B(n15209), .Z(n15211) );
  AND U17378 ( .A(n15212), .B(n15211), .Z(n15348) );
  NAND U17379 ( .A(n15214), .B(n15213), .Z(n15218) );
  NAND U17380 ( .A(n15216), .B(n15215), .Z(n15217) );
  NAND U17381 ( .A(n15218), .B(n15217), .Z(n15347) );
  XOR U17382 ( .A(n15350), .B(n15349), .Z(n15435) );
  XOR U17383 ( .A(n15436), .B(n15435), .Z(n15438) );
  NAND U17384 ( .A(n15220), .B(n15219), .Z(n15224) );
  NAND U17385 ( .A(n15222), .B(n15221), .Z(n15223) );
  NAND U17386 ( .A(n15224), .B(n15223), .Z(n15430) );
  AND U17387 ( .A(x[483]), .B(y[7829]), .Z(n15417) );
  XOR U17388 ( .A(n15418), .B(n15417), .Z(n15420) );
  AND U17389 ( .A(x[484]), .B(y[7828]), .Z(n15419) );
  XOR U17390 ( .A(n15420), .B(n15419), .Z(n15429) );
  XOR U17391 ( .A(n15430), .B(n15429), .Z(n15432) );
  AND U17392 ( .A(y[7823]), .B(x[489]), .Z(n15226) );
  NAND U17393 ( .A(y[7822]), .B(x[490]), .Z(n15225) );
  XNOR U17394 ( .A(n15226), .B(n15225), .Z(n15390) );
  AND U17395 ( .A(y[7818]), .B(x[494]), .Z(n15228) );
  NAND U17396 ( .A(y[7824]), .B(x[488]), .Z(n15227) );
  XNOR U17397 ( .A(n15228), .B(n15227), .Z(n15394) );
  NAND U17398 ( .A(x[491]), .B(y[7821]), .Z(n15395) );
  XOR U17399 ( .A(n15390), .B(n15389), .Z(n15431) );
  XOR U17400 ( .A(n15432), .B(n15431), .Z(n15437) );
  XNOR U17401 ( .A(n15438), .B(n15437), .Z(n15448) );
  NAND U17402 ( .A(n15230), .B(n15229), .Z(n15234) );
  NAND U17403 ( .A(n15232), .B(n15231), .Z(n15233) );
  AND U17404 ( .A(n15234), .B(n15233), .Z(n15447) );
  XOR U17405 ( .A(n15448), .B(n15447), .Z(n15449) );
  NAND U17406 ( .A(n15236), .B(n15235), .Z(n15240) );
  NAND U17407 ( .A(n15238), .B(n15237), .Z(n15239) );
  AND U17408 ( .A(n15240), .B(n15239), .Z(n15450) );
  XOR U17409 ( .A(n15449), .B(n15450), .Z(n15456) );
  NAND U17410 ( .A(n15242), .B(n15241), .Z(n15246) );
  NAND U17411 ( .A(n15244), .B(n15243), .Z(n15245) );
  NAND U17412 ( .A(n15246), .B(n15245), .Z(n15444) );
  NAND U17413 ( .A(n15248), .B(n15247), .Z(n15252) );
  NAND U17414 ( .A(n15250), .B(n15249), .Z(n15251) );
  NAND U17415 ( .A(n15252), .B(n15251), .Z(n15442) );
  NAND U17416 ( .A(n15254), .B(n15253), .Z(n15258) );
  NAND U17417 ( .A(n15256), .B(n15255), .Z(n15257) );
  AND U17418 ( .A(n15258), .B(n15257), .Z(n15356) );
  AND U17419 ( .A(x[480]), .B(y[7832]), .Z(n15423) );
  AND U17420 ( .A(x[504]), .B(y[7808]), .Z(n15424) );
  XOR U17421 ( .A(n15423), .B(n15424), .Z(n15425) );
  NAND U17422 ( .A(x[503]), .B(y[7809]), .Z(n15416) );
  XNOR U17423 ( .A(o[152]), .B(n15416), .Z(n15426) );
  XOR U17424 ( .A(n15425), .B(n15426), .Z(n15354) );
  AND U17425 ( .A(x[487]), .B(y[7825]), .Z(n15410) );
  AND U17426 ( .A(x[498]), .B(y[7814]), .Z(n15411) );
  XOR U17427 ( .A(n15410), .B(n15411), .Z(n15412) );
  AND U17428 ( .A(x[497]), .B(y[7815]), .Z(n15413) );
  XOR U17429 ( .A(n15412), .B(n15413), .Z(n15353) );
  XOR U17430 ( .A(n15354), .B(n15353), .Z(n15355) );
  NAND U17431 ( .A(n15260), .B(n15259), .Z(n15264) );
  NAND U17432 ( .A(n15262), .B(n15261), .Z(n15263) );
  AND U17433 ( .A(n15264), .B(n15263), .Z(n15342) );
  NAND U17434 ( .A(n15266), .B(n15265), .Z(n15270) );
  NAND U17435 ( .A(n15268), .B(n15267), .Z(n15269) );
  NAND U17436 ( .A(n15270), .B(n15269), .Z(n15341) );
  XOR U17437 ( .A(n15344), .B(n15343), .Z(n15441) );
  XOR U17438 ( .A(n15442), .B(n15441), .Z(n15443) );
  XNOR U17439 ( .A(n15444), .B(n15443), .Z(n15384) );
  NANDN U17440 ( .A(n15272), .B(n15271), .Z(n15276) );
  NAND U17441 ( .A(n15274), .B(n15273), .Z(n15275) );
  AND U17442 ( .A(n15276), .B(n15275), .Z(n15338) );
  NAND U17443 ( .A(n15278), .B(n15277), .Z(n15282) );
  NANDN U17444 ( .A(n15280), .B(n15279), .Z(n15281) );
  AND U17445 ( .A(n15282), .B(n15281), .Z(n15335) );
  NAND U17446 ( .A(n15284), .B(n15283), .Z(n15288) );
  NANDN U17447 ( .A(n15286), .B(n15285), .Z(n15287) );
  AND U17448 ( .A(n15288), .B(n15287), .Z(n15336) );
  XOR U17449 ( .A(n15335), .B(n15336), .Z(n15337) );
  XOR U17450 ( .A(n15338), .B(n15337), .Z(n15382) );
  NAND U17451 ( .A(n15290), .B(n15289), .Z(n15294) );
  NANDN U17452 ( .A(n15292), .B(n15291), .Z(n15293) );
  AND U17453 ( .A(n15294), .B(n15293), .Z(n15383) );
  XOR U17454 ( .A(n15382), .B(n15383), .Z(n15385) );
  XOR U17455 ( .A(n15384), .B(n15385), .Z(n15453) );
  NANDN U17456 ( .A(n15296), .B(n15295), .Z(n15300) );
  NANDN U17457 ( .A(n15298), .B(n15297), .Z(n15299) );
  NAND U17458 ( .A(n15300), .B(n15299), .Z(n15454) );
  XNOR U17459 ( .A(n15456), .B(n15455), .Z(n15462) );
  NAND U17460 ( .A(n15302), .B(n15301), .Z(n15306) );
  NANDN U17461 ( .A(n15304), .B(n15303), .Z(n15305) );
  AND U17462 ( .A(n15306), .B(n15305), .Z(n15332) );
  NANDN U17463 ( .A(n15308), .B(n15307), .Z(n15312) );
  NANDN U17464 ( .A(n15310), .B(n15309), .Z(n15311) );
  AND U17465 ( .A(n15312), .B(n15311), .Z(n15330) );
  NANDN U17466 ( .A(n15314), .B(n15313), .Z(n15318) );
  NAND U17467 ( .A(n15316), .B(n15315), .Z(n15317) );
  NAND U17468 ( .A(n15318), .B(n15317), .Z(n15329) );
  XOR U17469 ( .A(n15462), .B(n15463), .Z(n15465) );
  XNOR U17470 ( .A(n15464), .B(n15465), .Z(n15461) );
  NANDN U17471 ( .A(n15320), .B(n15319), .Z(n15324) );
  NANDN U17472 ( .A(n15322), .B(n15321), .Z(n15323) );
  AND U17473 ( .A(n15324), .B(n15323), .Z(n15460) );
  XOR U17474 ( .A(n15460), .B(n15459), .Z(n15328) );
  XNOR U17475 ( .A(n15461), .B(n15328), .Z(N313) );
  NANDN U17476 ( .A(n15330), .B(n15329), .Z(n15334) );
  NANDN U17477 ( .A(n15332), .B(n15331), .Z(n15333) );
  AND U17478 ( .A(n15334), .B(n15333), .Z(n15601) );
  NAND U17479 ( .A(n15336), .B(n15335), .Z(n15340) );
  NAND U17480 ( .A(n15338), .B(n15337), .Z(n15339) );
  AND U17481 ( .A(n15340), .B(n15339), .Z(n15476) );
  NANDN U17482 ( .A(n15342), .B(n15341), .Z(n15346) );
  NAND U17483 ( .A(n15344), .B(n15343), .Z(n15345) );
  AND U17484 ( .A(n15346), .B(n15345), .Z(n15482) );
  NANDN U17485 ( .A(n15348), .B(n15347), .Z(n15352) );
  NAND U17486 ( .A(n15350), .B(n15349), .Z(n15351) );
  NAND U17487 ( .A(n15352), .B(n15351), .Z(n15481) );
  NAND U17488 ( .A(n15354), .B(n15353), .Z(n15358) );
  NANDN U17489 ( .A(n15356), .B(n15355), .Z(n15357) );
  AND U17490 ( .A(n15358), .B(n15357), .Z(n15510) );
  AND U17491 ( .A(x[501]), .B(y[7816]), .Z(n16249) );
  NAND U17492 ( .A(n16249), .B(n15359), .Z(n15363) );
  NANDN U17493 ( .A(n15361), .B(n15360), .Z(n15362) );
  AND U17494 ( .A(n15363), .B(n15362), .Z(n15577) );
  NAND U17495 ( .A(x[502]), .B(y[7811]), .Z(n15551) );
  NAND U17496 ( .A(x[485]), .B(y[7828]), .Z(n15549) );
  NAND U17497 ( .A(x[497]), .B(y[7816]), .Z(n15550) );
  XNOR U17498 ( .A(n15549), .B(n15550), .Z(n15552) );
  XOR U17499 ( .A(n15551), .B(n15552), .Z(n15574) );
  AND U17500 ( .A(y[7813]), .B(x[500]), .Z(n15365) );
  NAND U17501 ( .A(y[7812]), .B(x[501]), .Z(n15364) );
  XNOR U17502 ( .A(n15365), .B(n15364), .Z(n15560) );
  AND U17503 ( .A(x[499]), .B(y[7814]), .Z(n15559) );
  XOR U17504 ( .A(n15560), .B(n15559), .Z(n15575) );
  XOR U17505 ( .A(n15574), .B(n15575), .Z(n15576) );
  NANDN U17506 ( .A(n15722), .B(n15558), .Z(n15369) );
  NANDN U17507 ( .A(n15367), .B(n15366), .Z(n15368) );
  AND U17508 ( .A(n15369), .B(n15368), .Z(n15583) );
  NAND U17509 ( .A(x[495]), .B(y[7818]), .Z(n15565) );
  NAND U17510 ( .A(x[498]), .B(y[7815]), .Z(n15563) );
  NAND U17511 ( .A(x[486]), .B(y[7827]), .Z(n15564) );
  XNOR U17512 ( .A(n15563), .B(n15564), .Z(n15566) );
  XOR U17513 ( .A(n15565), .B(n15566), .Z(n15581) );
  NAND U17514 ( .A(x[503]), .B(y[7810]), .Z(n15547) );
  NAND U17515 ( .A(x[484]), .B(y[7829]), .Z(n15545) );
  NAND U17516 ( .A(x[496]), .B(y[7817]), .Z(n15546) );
  XNOR U17517 ( .A(n15545), .B(n15546), .Z(n15548) );
  XOR U17518 ( .A(n15547), .B(n15548), .Z(n15580) );
  XOR U17519 ( .A(n15581), .B(n15580), .Z(n15582) );
  XOR U17520 ( .A(n15583), .B(n15582), .Z(n15507) );
  XOR U17521 ( .A(n15508), .B(n15507), .Z(n15509) );
  XOR U17522 ( .A(n15510), .B(n15509), .Z(n15522) );
  NAND U17523 ( .A(n15371), .B(n15370), .Z(n15375) );
  NANDN U17524 ( .A(n15373), .B(n15372), .Z(n15374) );
  AND U17525 ( .A(n15375), .B(n15374), .Z(n15520) );
  NAND U17526 ( .A(n15377), .B(n15376), .Z(n15381) );
  NANDN U17527 ( .A(n15379), .B(n15378), .Z(n15380) );
  NAND U17528 ( .A(n15381), .B(n15380), .Z(n15519) );
  XNOR U17529 ( .A(n15484), .B(n15483), .Z(n15475) );
  NAND U17530 ( .A(n15383), .B(n15382), .Z(n15387) );
  NAND U17531 ( .A(n15385), .B(n15384), .Z(n15386) );
  NAND U17532 ( .A(n15387), .B(n15386), .Z(n15477) );
  XNOR U17533 ( .A(n15478), .B(n15477), .Z(n15472) );
  NANDN U17534 ( .A(n15492), .B(n15388), .Z(n15392) );
  NAND U17535 ( .A(n15390), .B(n15389), .Z(n15391) );
  AND U17536 ( .A(n15392), .B(n15391), .Z(n15514) );
  AND U17537 ( .A(x[494]), .B(y[7824]), .Z(n16382) );
  NAND U17538 ( .A(n16382), .B(n15393), .Z(n15397) );
  NANDN U17539 ( .A(n15395), .B(n15394), .Z(n15396) );
  NAND U17540 ( .A(n15397), .B(n15396), .Z(n15541) );
  NAND U17541 ( .A(x[491]), .B(y[7822]), .Z(n15556) );
  NAND U17542 ( .A(x[492]), .B(y[7821]), .Z(n15554) );
  NAND U17543 ( .A(x[487]), .B(y[7826]), .Z(n15555) );
  XOR U17544 ( .A(n15554), .B(n15555), .Z(n15557) );
  XOR U17545 ( .A(n15556), .B(n15557), .Z(n15540) );
  NAND U17546 ( .A(x[504]), .B(y[7809]), .Z(n15553) );
  XNOR U17547 ( .A(o[153]), .B(n15553), .Z(n15528) );
  AND U17548 ( .A(x[481]), .B(y[7832]), .Z(n15527) );
  XOR U17549 ( .A(n15528), .B(n15527), .Z(n15530) );
  AND U17550 ( .A(x[493]), .B(y[7820]), .Z(n15529) );
  XOR U17551 ( .A(n15530), .B(n15529), .Z(n15539) );
  XOR U17552 ( .A(n15541), .B(n15542), .Z(n15513) );
  NAND U17553 ( .A(n15399), .B(n15398), .Z(n15403) );
  AND U17554 ( .A(n15401), .B(n15400), .Z(n15402) );
  ANDN U17555 ( .B(n15403), .A(n15402), .Z(n15502) );
  AND U17556 ( .A(n15405), .B(n15404), .Z(n15409) );
  NAND U17557 ( .A(n15407), .B(n15406), .Z(n15408) );
  NANDN U17558 ( .A(n15409), .B(n15408), .Z(n15501) );
  NAND U17559 ( .A(n15411), .B(n15410), .Z(n15415) );
  NAND U17560 ( .A(n15413), .B(n15412), .Z(n15414) );
  AND U17561 ( .A(n15415), .B(n15414), .Z(n15498) );
  NAND U17562 ( .A(x[488]), .B(y[7825]), .Z(n15493) );
  XNOR U17563 ( .A(n15491), .B(n15492), .Z(n15494) );
  XOR U17564 ( .A(n15493), .B(n15494), .Z(n15496) );
  ANDN U17565 ( .B(o[152]), .A(n15416), .Z(n15489) );
  NAND U17566 ( .A(x[505]), .B(y[7808]), .Z(n15487) );
  NAND U17567 ( .A(x[480]), .B(y[7833]), .Z(n15488) );
  XNOR U17568 ( .A(n15487), .B(n15488), .Z(n15490) );
  XNOR U17569 ( .A(n15489), .B(n15490), .Z(n15495) );
  XOR U17570 ( .A(n15496), .B(n15495), .Z(n15497) );
  XOR U17571 ( .A(n15504), .B(n15503), .Z(n15515) );
  XOR U17572 ( .A(n15516), .B(n15515), .Z(n15595) );
  NAND U17573 ( .A(n15418), .B(n15417), .Z(n15422) );
  AND U17574 ( .A(n15420), .B(n15419), .Z(n15421) );
  ANDN U17575 ( .B(n15422), .A(n15421), .Z(n15571) );
  NAND U17576 ( .A(n15424), .B(n15423), .Z(n15428) );
  NAND U17577 ( .A(n15426), .B(n15425), .Z(n15427) );
  AND U17578 ( .A(n15428), .B(n15427), .Z(n15569) );
  AND U17579 ( .A(x[494]), .B(y[7819]), .Z(n15534) );
  AND U17580 ( .A(x[482]), .B(y[7831]), .Z(n15533) );
  XOR U17581 ( .A(n15534), .B(n15533), .Z(n15536) );
  AND U17582 ( .A(x[483]), .B(y[7830]), .Z(n15535) );
  XOR U17583 ( .A(n15536), .B(n15535), .Z(n15568) );
  NAND U17584 ( .A(n15430), .B(n15429), .Z(n15434) );
  NAND U17585 ( .A(n15432), .B(n15431), .Z(n15433) );
  AND U17586 ( .A(n15434), .B(n15433), .Z(n15592) );
  NAND U17587 ( .A(n15436), .B(n15435), .Z(n15440) );
  NAND U17588 ( .A(n15438), .B(n15437), .Z(n15439) );
  NAND U17589 ( .A(n15440), .B(n15439), .Z(n15587) );
  NAND U17590 ( .A(n15442), .B(n15441), .Z(n15446) );
  NAND U17591 ( .A(n15444), .B(n15443), .Z(n15445) );
  AND U17592 ( .A(n15446), .B(n15445), .Z(n15588) );
  XNOR U17593 ( .A(n15589), .B(n15588), .Z(n15470) );
  NAND U17594 ( .A(n15448), .B(n15447), .Z(n15452) );
  NAND U17595 ( .A(n15450), .B(n15449), .Z(n15451) );
  AND U17596 ( .A(n15452), .B(n15451), .Z(n15469) );
  XOR U17597 ( .A(n15470), .B(n15469), .Z(n15471) );
  XNOR U17598 ( .A(n15472), .B(n15471), .Z(n15599) );
  NANDN U17599 ( .A(n15454), .B(n15453), .Z(n15458) );
  NAND U17600 ( .A(n15456), .B(n15455), .Z(n15457) );
  NAND U17601 ( .A(n15458), .B(n15457), .Z(n15598) );
  XOR U17602 ( .A(n15599), .B(n15598), .Z(n15600) );
  XNOR U17603 ( .A(n15601), .B(n15600), .Z(n15606) );
  NANDN U17604 ( .A(n15463), .B(n15462), .Z(n15467) );
  NANDN U17605 ( .A(n15465), .B(n15464), .Z(n15466) );
  AND U17606 ( .A(n15467), .B(n15466), .Z(n15604) );
  XOR U17607 ( .A(n15605), .B(n15604), .Z(n15468) );
  XNOR U17608 ( .A(n15606), .B(n15468), .Z(N314) );
  NAND U17609 ( .A(n15470), .B(n15469), .Z(n15474) );
  NAND U17610 ( .A(n15472), .B(n15471), .Z(n15473) );
  NAND U17611 ( .A(n15474), .B(n15473), .Z(n15749) );
  NANDN U17612 ( .A(n15476), .B(n15475), .Z(n15480) );
  NAND U17613 ( .A(n15478), .B(n15477), .Z(n15479) );
  AND U17614 ( .A(n15480), .B(n15479), .Z(n15748) );
  XOR U17615 ( .A(n15749), .B(n15748), .Z(n15751) );
  NANDN U17616 ( .A(n15482), .B(n15481), .Z(n15486) );
  NAND U17617 ( .A(n15484), .B(n15483), .Z(n15485) );
  AND U17618 ( .A(n15486), .B(n15485), .Z(n15745) );
  AND U17619 ( .A(x[482]), .B(y[7832]), .Z(n15628) );
  XOR U17620 ( .A(n15629), .B(n15628), .Z(n15631) );
  NAND U17621 ( .A(x[504]), .B(y[7810]), .Z(n15630) );
  XNOR U17622 ( .A(n15631), .B(n15630), .Z(n15665) );
  XOR U17623 ( .A(n15665), .B(n15664), .Z(n15667) );
  XOR U17624 ( .A(n15667), .B(n15666), .Z(n15699) );
  NAND U17625 ( .A(n15496), .B(n15495), .Z(n15500) );
  NANDN U17626 ( .A(n15498), .B(n15497), .Z(n15499) );
  AND U17627 ( .A(n15500), .B(n15499), .Z(n15698) );
  NANDN U17628 ( .A(n15502), .B(n15501), .Z(n15506) );
  NAND U17629 ( .A(n15504), .B(n15503), .Z(n15505) );
  NAND U17630 ( .A(n15506), .B(n15505), .Z(n15701) );
  NAND U17631 ( .A(n15508), .B(n15507), .Z(n15512) );
  NAND U17632 ( .A(n15510), .B(n15509), .Z(n15511) );
  AND U17633 ( .A(n15512), .B(n15511), .Z(n15693) );
  NANDN U17634 ( .A(n15514), .B(n15513), .Z(n15518) );
  NAND U17635 ( .A(n15516), .B(n15515), .Z(n15517) );
  AND U17636 ( .A(n15518), .B(n15517), .Z(n15692) );
  XOR U17637 ( .A(n15695), .B(n15694), .Z(n15743) );
  NANDN U17638 ( .A(n15520), .B(n15519), .Z(n15524) );
  NANDN U17639 ( .A(n15522), .B(n15521), .Z(n15523) );
  AND U17640 ( .A(n15524), .B(n15523), .Z(n15617) );
  AND U17641 ( .A(x[492]), .B(y[7822]), .Z(n15806) );
  AND U17642 ( .A(x[485]), .B(y[7829]), .Z(n15675) );
  XOR U17643 ( .A(n15806), .B(n15675), .Z(n15677) );
  NAND U17644 ( .A(x[490]), .B(y[7824]), .Z(n15676) );
  XNOR U17645 ( .A(n15677), .B(n15676), .Z(n15707) );
  AND U17646 ( .A(x[487]), .B(y[7827]), .Z(n15704) );
  AND U17647 ( .A(y[7828]), .B(x[486]), .Z(n15526) );
  NAND U17648 ( .A(y[7826]), .B(x[488]), .Z(n15525) );
  XNOR U17649 ( .A(n15526), .B(n15525), .Z(n15723) );
  NAND U17650 ( .A(x[489]), .B(y[7825]), .Z(n15724) );
  XOR U17651 ( .A(n15723), .B(n15724), .Z(n15705) );
  XOR U17652 ( .A(n15707), .B(n15706), .Z(n15654) );
  NAND U17653 ( .A(n15528), .B(n15527), .Z(n15532) );
  NAND U17654 ( .A(n15530), .B(n15529), .Z(n15531) );
  NAND U17655 ( .A(n15532), .B(n15531), .Z(n15653) );
  NAND U17656 ( .A(n15534), .B(n15533), .Z(n15538) );
  NAND U17657 ( .A(n15536), .B(n15535), .Z(n15537) );
  NAND U17658 ( .A(n15538), .B(n15537), .Z(n15652) );
  XNOR U17659 ( .A(n15653), .B(n15652), .Z(n15655) );
  NANDN U17660 ( .A(n15540), .B(n15539), .Z(n15544) );
  NAND U17661 ( .A(n15542), .B(n15541), .Z(n15543) );
  AND U17662 ( .A(n15544), .B(n15543), .Z(n15686) );
  XOR U17663 ( .A(n15621), .B(n15620), .Z(n15623) );
  ANDN U17664 ( .B(o[153]), .A(n15553), .Z(n15716) );
  NAND U17665 ( .A(x[494]), .B(y[7820]), .Z(n15717) );
  XNOR U17666 ( .A(n15716), .B(n15717), .Z(n15718) );
  NAND U17667 ( .A(x[481]), .B(y[7833]), .Z(n15719) );
  XNOR U17668 ( .A(n15718), .B(n15719), .Z(n15669) );
  NAND U17669 ( .A(x[505]), .B(y[7809]), .Z(n15727) );
  XNOR U17670 ( .A(o[154]), .B(n15727), .Z(n15680) );
  NAND U17671 ( .A(x[506]), .B(y[7808]), .Z(n15681) );
  XNOR U17672 ( .A(n15680), .B(n15681), .Z(n15683) );
  AND U17673 ( .A(x[480]), .B(y[7834]), .Z(n15682) );
  XOR U17674 ( .A(n15683), .B(n15682), .Z(n15668) );
  XOR U17675 ( .A(n15669), .B(n15668), .Z(n15671) );
  XOR U17676 ( .A(n15671), .B(n15670), .Z(n15622) );
  XOR U17677 ( .A(n15623), .B(n15622), .Z(n15661) );
  AND U17678 ( .A(x[501]), .B(y[7813]), .Z(n15710) );
  NAND U17679 ( .A(n15710), .B(n15558), .Z(n15562) );
  NAND U17680 ( .A(n15560), .B(n15559), .Z(n15561) );
  NAND U17681 ( .A(n15562), .B(n15561), .Z(n15648) );
  XOR U17682 ( .A(n15711), .B(n15710), .Z(n15713) );
  NAND U17683 ( .A(x[500]), .B(y[7814]), .Z(n15712) );
  XNOR U17684 ( .A(n15713), .B(n15712), .Z(n15647) );
  NAND U17685 ( .A(x[503]), .B(y[7811]), .Z(n15635) );
  XNOR U17686 ( .A(n15634), .B(n15635), .Z(n15637) );
  AND U17687 ( .A(x[502]), .B(y[7812]), .Z(n15636) );
  XOR U17688 ( .A(n15637), .B(n15636), .Z(n15646) );
  XOR U17689 ( .A(n15647), .B(n15646), .Z(n15649) );
  XOR U17690 ( .A(n15648), .B(n15649), .Z(n15659) );
  IV U17691 ( .A(n15659), .Z(n15567) );
  AND U17692 ( .A(x[484]), .B(y[7830]), .Z(n15640) );
  XOR U17693 ( .A(n15641), .B(n15640), .Z(n15643) );
  AND U17694 ( .A(x[499]), .B(y[7815]), .Z(n15728) );
  NAND U17695 ( .A(x[483]), .B(y[7831]), .Z(n15729) );
  XNOR U17696 ( .A(n15728), .B(n15729), .Z(n15731) );
  AND U17697 ( .A(x[491]), .B(y[7823]), .Z(n15730) );
  XOR U17698 ( .A(n15731), .B(n15730), .Z(n15624) );
  XOR U17699 ( .A(n15625), .B(n15624), .Z(n15627) );
  XNOR U17700 ( .A(n15627), .B(n15626), .Z(n15658) );
  XOR U17701 ( .A(n15567), .B(n15658), .Z(n15660) );
  XOR U17702 ( .A(n15689), .B(n15688), .Z(n15615) );
  NANDN U17703 ( .A(n15569), .B(n15568), .Z(n15573) );
  NANDN U17704 ( .A(n15571), .B(n15570), .Z(n15572) );
  AND U17705 ( .A(n15573), .B(n15572), .Z(n15739) );
  NAND U17706 ( .A(n15575), .B(n15574), .Z(n15579) );
  NANDN U17707 ( .A(n15577), .B(n15576), .Z(n15578) );
  AND U17708 ( .A(n15579), .B(n15578), .Z(n15737) );
  NAND U17709 ( .A(n15581), .B(n15580), .Z(n15585) );
  NANDN U17710 ( .A(n15583), .B(n15582), .Z(n15584) );
  NAND U17711 ( .A(n15585), .B(n15584), .Z(n15736) );
  NANDN U17712 ( .A(n15587), .B(n15586), .Z(n15591) );
  NAND U17713 ( .A(n15589), .B(n15588), .Z(n15590) );
  AND U17714 ( .A(n15591), .B(n15590), .Z(n15608) );
  NANDN U17715 ( .A(n15593), .B(n15592), .Z(n15597) );
  NANDN U17716 ( .A(n15595), .B(n15594), .Z(n15596) );
  NAND U17717 ( .A(n15597), .B(n15596), .Z(n15609) );
  XOR U17718 ( .A(n15611), .B(n15610), .Z(n15750) );
  XOR U17719 ( .A(n15751), .B(n15750), .Z(n15756) );
  NAND U17720 ( .A(n15599), .B(n15598), .Z(n15603) );
  NAND U17721 ( .A(n15601), .B(n15600), .Z(n15602) );
  NAND U17722 ( .A(n15603), .B(n15602), .Z(n15754) );
  XOR U17723 ( .A(n15754), .B(n15755), .Z(n15607) );
  XNOR U17724 ( .A(n15756), .B(n15607), .Z(N315) );
  NANDN U17725 ( .A(n15609), .B(n15608), .Z(n15613) );
  NAND U17726 ( .A(n15611), .B(n15610), .Z(n15612) );
  AND U17727 ( .A(n15613), .B(n15612), .Z(n15897) );
  NANDN U17728 ( .A(n15615), .B(n15614), .Z(n15619) );
  NANDN U17729 ( .A(n15617), .B(n15616), .Z(n15618) );
  NAND U17730 ( .A(n15619), .B(n15618), .Z(n15760) );
  NAND U17731 ( .A(n15629), .B(n15628), .Z(n15633) );
  ANDN U17732 ( .B(n15631), .A(n15630), .Z(n15632) );
  ANDN U17733 ( .B(n15633), .A(n15632), .Z(n15783) );
  NANDN U17734 ( .A(n15635), .B(n15634), .Z(n15639) );
  NAND U17735 ( .A(n15637), .B(n15636), .Z(n15638) );
  NAND U17736 ( .A(n15639), .B(n15638), .Z(n15782) );
  XNOR U17737 ( .A(n15783), .B(n15782), .Z(n15784) );
  NAND U17738 ( .A(n15641), .B(n15640), .Z(n15645) );
  ANDN U17739 ( .B(n15643), .A(n15642), .Z(n15644) );
  ANDN U17740 ( .B(n15645), .A(n15644), .Z(n15795) );
  AND U17741 ( .A(x[480]), .B(y[7835]), .Z(n15859) );
  NAND U17742 ( .A(x[507]), .B(y[7808]), .Z(n15860) );
  XNOR U17743 ( .A(n15859), .B(n15860), .Z(n15861) );
  NAND U17744 ( .A(x[506]), .B(y[7809]), .Z(n15850) );
  XOR U17745 ( .A(o[155]), .B(n15850), .Z(n15862) );
  XNOR U17746 ( .A(n15861), .B(n15862), .Z(n15792) );
  AND U17747 ( .A(x[489]), .B(y[7826]), .Z(n15844) );
  NAND U17748 ( .A(x[501]), .B(y[7814]), .Z(n15845) );
  XNOR U17749 ( .A(n15844), .B(n15845), .Z(n15846) );
  NAND U17750 ( .A(x[498]), .B(y[7817]), .Z(n15847) );
  XOR U17751 ( .A(n15846), .B(n15847), .Z(n15793) );
  XNOR U17752 ( .A(n15792), .B(n15793), .Z(n15794) );
  XOR U17753 ( .A(n15795), .B(n15794), .Z(n15785) );
  XNOR U17754 ( .A(n15784), .B(n15785), .Z(n15870) );
  XOR U17755 ( .A(n15869), .B(n15870), .Z(n15872) );
  XOR U17756 ( .A(n15871), .B(n15872), .Z(n15888) );
  NAND U17757 ( .A(n15647), .B(n15646), .Z(n15651) );
  NAND U17758 ( .A(n15649), .B(n15648), .Z(n15650) );
  AND U17759 ( .A(n15651), .B(n15650), .Z(n15886) );
  NAND U17760 ( .A(n15653), .B(n15652), .Z(n15657) );
  NANDN U17761 ( .A(n15655), .B(n15654), .Z(n15656) );
  AND U17762 ( .A(n15657), .B(n15656), .Z(n15885) );
  XOR U17763 ( .A(n15886), .B(n15885), .Z(n15887) );
  NANDN U17764 ( .A(n15659), .B(n15658), .Z(n15663) );
  NANDN U17765 ( .A(n15661), .B(n15660), .Z(n15662) );
  AND U17766 ( .A(n15663), .B(n15662), .Z(n15873) );
  AND U17767 ( .A(x[495]), .B(y[7820]), .Z(n15812) );
  AND U17768 ( .A(x[482]), .B(y[7833]), .Z(n15811) );
  XOR U17769 ( .A(n15812), .B(n15811), .Z(n15814) );
  AND U17770 ( .A(x[483]), .B(y[7832]), .Z(n15813) );
  XOR U17771 ( .A(n15814), .B(n15813), .Z(n15827) );
  AND U17772 ( .A(x[499]), .B(y[7816]), .Z(n15838) );
  NAND U17773 ( .A(x[505]), .B(y[7810]), .Z(n15839) );
  XNOR U17774 ( .A(n15838), .B(n15839), .Z(n15840) );
  NAND U17775 ( .A(x[486]), .B(y[7829]), .Z(n15841) );
  XOR U17776 ( .A(n15840), .B(n15841), .Z(n15828) );
  XNOR U17777 ( .A(n15827), .B(n15828), .Z(n15829) );
  NAND U17778 ( .A(x[496]), .B(y[7819]), .Z(n15798) );
  XOR U17779 ( .A(n15798), .B(n15672), .Z(n15801) );
  XOR U17780 ( .A(n15800), .B(n15801), .Z(n15808) );
  AND U17781 ( .A(y[7822]), .B(x[493]), .Z(n15674) );
  NAND U17782 ( .A(y[7823]), .B(x[492]), .Z(n15673) );
  XNOR U17783 ( .A(n15674), .B(n15673), .Z(n15807) );
  XOR U17784 ( .A(n15808), .B(n15807), .Z(n15830) );
  XNOR U17785 ( .A(n15829), .B(n15830), .Z(n15779) );
  NAND U17786 ( .A(n15806), .B(n15675), .Z(n15679) );
  ANDN U17787 ( .B(n15677), .A(n15676), .Z(n15678) );
  ANDN U17788 ( .B(n15679), .A(n15678), .Z(n15777) );
  NANDN U17789 ( .A(n15681), .B(n15680), .Z(n15685) );
  NAND U17790 ( .A(n15683), .B(n15682), .Z(n15684) );
  NAND U17791 ( .A(n15685), .B(n15684), .Z(n15776) );
  XNOR U17792 ( .A(n15777), .B(n15776), .Z(n15778) );
  XOR U17793 ( .A(n15779), .B(n15778), .Z(n15865) );
  XNOR U17794 ( .A(n15866), .B(n15865), .Z(n15868) );
  XOR U17795 ( .A(n15867), .B(n15868), .Z(n15874) );
  NANDN U17796 ( .A(n15687), .B(n15686), .Z(n15691) );
  NAND U17797 ( .A(n15689), .B(n15688), .Z(n15690) );
  AND U17798 ( .A(n15691), .B(n15690), .Z(n15875) );
  XOR U17799 ( .A(n15876), .B(n15875), .Z(n15758) );
  XOR U17800 ( .A(n15760), .B(n15761), .Z(n15766) );
  NANDN U17801 ( .A(n15693), .B(n15692), .Z(n15697) );
  NAND U17802 ( .A(n15695), .B(n15694), .Z(n15696) );
  AND U17803 ( .A(n15697), .B(n15696), .Z(n15765) );
  NANDN U17804 ( .A(n15699), .B(n15698), .Z(n15703) );
  NANDN U17805 ( .A(n15701), .B(n15700), .Z(n15702) );
  NAND U17806 ( .A(n15703), .B(n15702), .Z(n15771) );
  NANDN U17807 ( .A(n15705), .B(n15704), .Z(n15709) );
  NAND U17808 ( .A(n15707), .B(n15706), .Z(n15708) );
  NAND U17809 ( .A(n15709), .B(n15708), .Z(n15881) );
  NAND U17810 ( .A(n15711), .B(n15710), .Z(n15715) );
  ANDN U17811 ( .B(n15713), .A(n15712), .Z(n15714) );
  ANDN U17812 ( .B(n15715), .A(n15714), .Z(n15820) );
  NANDN U17813 ( .A(n15717), .B(n15716), .Z(n15721) );
  NANDN U17814 ( .A(n15719), .B(n15718), .Z(n15720) );
  NAND U17815 ( .A(n15721), .B(n15720), .Z(n15819) );
  XNOR U17816 ( .A(n15820), .B(n15819), .Z(n15822) );
  AND U17817 ( .A(x[488]), .B(y[7828]), .Z(n15852) );
  NANDN U17818 ( .A(n15722), .B(n15852), .Z(n15726) );
  NANDN U17819 ( .A(n15724), .B(n15723), .Z(n15725) );
  NAND U17820 ( .A(n15726), .B(n15725), .Z(n15790) );
  ANDN U17821 ( .B(o[154]), .A(n15727), .Z(n15818) );
  AND U17822 ( .A(x[494]), .B(y[7821]), .Z(n15816) );
  AND U17823 ( .A(x[481]), .B(y[7834]), .Z(n15815) );
  XOR U17824 ( .A(n15816), .B(n15815), .Z(n15817) );
  XOR U17825 ( .A(n15818), .B(n15817), .Z(n15789) );
  AND U17826 ( .A(x[497]), .B(y[7818]), .Z(n15853) );
  NAND U17827 ( .A(x[484]), .B(y[7831]), .Z(n15854) );
  XNOR U17828 ( .A(n15853), .B(n15854), .Z(n15856) );
  AND U17829 ( .A(x[485]), .B(y[7830]), .Z(n15855) );
  XOR U17830 ( .A(n15856), .B(n15855), .Z(n15788) );
  XOR U17831 ( .A(n15789), .B(n15788), .Z(n15791) );
  XOR U17832 ( .A(n15790), .B(n15791), .Z(n15821) );
  XOR U17833 ( .A(n15822), .B(n15821), .Z(n15880) );
  NANDN U17834 ( .A(n15729), .B(n15728), .Z(n15733) );
  NAND U17835 ( .A(n15731), .B(n15730), .Z(n15732) );
  AND U17836 ( .A(n15733), .B(n15732), .Z(n15826) );
  AND U17837 ( .A(y[7811]), .B(x[504]), .Z(n15735) );
  NAND U17838 ( .A(y[7815]), .B(x[500]), .Z(n15734) );
  XNOR U17839 ( .A(n15735), .B(n15734), .Z(n15834) );
  NAND U17840 ( .A(x[487]), .B(y[7828]), .Z(n15835) );
  XNOR U17841 ( .A(n15834), .B(n15835), .Z(n15824) );
  AND U17842 ( .A(x[488]), .B(y[7827]), .Z(n15803) );
  AND U17843 ( .A(x[503]), .B(y[7812]), .Z(n15802) );
  XOR U17844 ( .A(n15803), .B(n15802), .Z(n15805) );
  AND U17845 ( .A(x[502]), .B(y[7813]), .Z(n15804) );
  XOR U17846 ( .A(n15805), .B(n15804), .Z(n15823) );
  XOR U17847 ( .A(n15824), .B(n15823), .Z(n15825) );
  XNOR U17848 ( .A(n15826), .B(n15825), .Z(n15879) );
  XOR U17849 ( .A(n15880), .B(n15879), .Z(n15882) );
  XNOR U17850 ( .A(n15881), .B(n15882), .Z(n15770) );
  XOR U17851 ( .A(n15771), .B(n15770), .Z(n15773) );
  NANDN U17852 ( .A(n15737), .B(n15736), .Z(n15741) );
  NANDN U17853 ( .A(n15739), .B(n15738), .Z(n15740) );
  AND U17854 ( .A(n15741), .B(n15740), .Z(n15772) );
  XOR U17855 ( .A(n15773), .B(n15772), .Z(n15764) );
  XNOR U17856 ( .A(n15766), .B(n15767), .Z(n15895) );
  NANDN U17857 ( .A(n15743), .B(n15742), .Z(n15747) );
  NANDN U17858 ( .A(n15745), .B(n15744), .Z(n15746) );
  NAND U17859 ( .A(n15747), .B(n15746), .Z(n15894) );
  XOR U17860 ( .A(n15895), .B(n15894), .Z(n15896) );
  XOR U17861 ( .A(n15897), .B(n15896), .Z(n15893) );
  NAND U17862 ( .A(n15749), .B(n15748), .Z(n15753) );
  NAND U17863 ( .A(n15751), .B(n15750), .Z(n15752) );
  NAND U17864 ( .A(n15753), .B(n15752), .Z(n15892) );
  XOR U17865 ( .A(n15892), .B(n15891), .Z(n15757) );
  XNOR U17866 ( .A(n15893), .B(n15757), .Z(N316) );
  NANDN U17867 ( .A(n15759), .B(n15758), .Z(n15763) );
  NANDN U17868 ( .A(n15761), .B(n15760), .Z(n15762) );
  AND U17869 ( .A(n15763), .B(n15762), .Z(n16029) );
  NANDN U17870 ( .A(n15765), .B(n15764), .Z(n15769) );
  NAND U17871 ( .A(n15767), .B(n15766), .Z(n15768) );
  AND U17872 ( .A(n15769), .B(n15768), .Z(n16028) );
  NAND U17873 ( .A(n15771), .B(n15770), .Z(n15775) );
  NAND U17874 ( .A(n15773), .B(n15772), .Z(n15774) );
  AND U17875 ( .A(n15775), .B(n15774), .Z(n15901) );
  NANDN U17876 ( .A(n15777), .B(n15776), .Z(n15781) );
  NAND U17877 ( .A(n15779), .B(n15778), .Z(n15780) );
  AND U17878 ( .A(n15781), .B(n15780), .Z(n15914) );
  NANDN U17879 ( .A(n15783), .B(n15782), .Z(n15787) );
  NANDN U17880 ( .A(n15785), .B(n15784), .Z(n15786) );
  AND U17881 ( .A(n15787), .B(n15786), .Z(n15992) );
  NANDN U17882 ( .A(n15793), .B(n15792), .Z(n15797) );
  NANDN U17883 ( .A(n15795), .B(n15794), .Z(n15796) );
  NAND U17884 ( .A(n15797), .B(n15796), .Z(n15989) );
  XNOR U17885 ( .A(n15990), .B(n15989), .Z(n15991) );
  XNOR U17886 ( .A(n15992), .B(n15991), .Z(n15913) );
  XNOR U17887 ( .A(n15914), .B(n15913), .Z(n15916) );
  AND U17888 ( .A(x[487]), .B(y[7829]), .Z(n15948) );
  AND U17889 ( .A(x[492]), .B(y[7824]), .Z(n15947) );
  XOR U17890 ( .A(n15948), .B(n15947), .Z(n15950) );
  AND U17891 ( .A(x[491]), .B(y[7825]), .Z(n15949) );
  XOR U17892 ( .A(n15950), .B(n15949), .Z(n15970) );
  AND U17893 ( .A(x[507]), .B(y[7809]), .Z(n15955) );
  XOR U17894 ( .A(o[156]), .B(n15955), .Z(n15962) );
  AND U17895 ( .A(x[506]), .B(y[7810]), .Z(n15961) );
  XOR U17896 ( .A(n15962), .B(n15961), .Z(n15964) );
  AND U17897 ( .A(x[495]), .B(y[7821]), .Z(n15963) );
  XOR U17898 ( .A(n15964), .B(n15963), .Z(n15969) );
  XOR U17899 ( .A(n15970), .B(n15969), .Z(n15971) );
  XNOR U17900 ( .A(n15972), .B(n15971), .Z(n15996) );
  AND U17901 ( .A(x[497]), .B(y[7819]), .Z(n15922) );
  AND U17902 ( .A(x[502]), .B(y[7814]), .Z(n15921) );
  XOR U17903 ( .A(n15922), .B(n15921), .Z(n15924) );
  AND U17904 ( .A(x[484]), .B(y[7832]), .Z(n15923) );
  XOR U17905 ( .A(n15924), .B(n15923), .Z(n15974) );
  AND U17906 ( .A(x[486]), .B(y[7830]), .Z(n16117) );
  AND U17907 ( .A(x[499]), .B(y[7817]), .Z(n15956) );
  XOR U17908 ( .A(n16117), .B(n15956), .Z(n15958) );
  XOR U17909 ( .A(n15958), .B(n15957), .Z(n15973) );
  XOR U17910 ( .A(n15974), .B(n15973), .Z(n15976) );
  XOR U17911 ( .A(n15975), .B(n15976), .Z(n15995) );
  XOR U17912 ( .A(n15996), .B(n15995), .Z(n15998) );
  NAND U17913 ( .A(n15806), .B(n15966), .Z(n15810) );
  NANDN U17914 ( .A(n15808), .B(n15807), .Z(n15809) );
  NAND U17915 ( .A(n15810), .B(n15809), .Z(n15919) );
  XOR U17916 ( .A(n15917), .B(n15918), .Z(n15920) );
  XOR U17917 ( .A(n15919), .B(n15920), .Z(n15997) );
  XOR U17918 ( .A(n15998), .B(n15997), .Z(n15915) );
  XOR U17919 ( .A(n15916), .B(n15915), .Z(n16018) );
  NANDN U17920 ( .A(n15828), .B(n15827), .Z(n15832) );
  NANDN U17921 ( .A(n15830), .B(n15829), .Z(n15831) );
  NAND U17922 ( .A(n15832), .B(n15831), .Z(n15977) );
  XNOR U17923 ( .A(n15978), .B(n15977), .Z(n15979) );
  XNOR U17924 ( .A(n15980), .B(n15979), .Z(n16016) );
  AND U17925 ( .A(x[500]), .B(y[7811]), .Z(n15833) );
  AND U17926 ( .A(x[504]), .B(y[7815]), .Z(n16266) );
  NAND U17927 ( .A(n15833), .B(n16266), .Z(n15837) );
  NANDN U17928 ( .A(n15835), .B(n15834), .Z(n15836) );
  NAND U17929 ( .A(n15837), .B(n15836), .Z(n16010) );
  AND U17930 ( .A(x[505]), .B(y[7811]), .Z(n15945) );
  XOR U17931 ( .A(n15946), .B(n15945), .Z(n15944) );
  AND U17932 ( .A(x[481]), .B(y[7835]), .Z(n15943) );
  XOR U17933 ( .A(n15944), .B(n15943), .Z(n16008) );
  AND U17934 ( .A(x[496]), .B(y[7820]), .Z(n15940) );
  AND U17935 ( .A(x[504]), .B(y[7812]), .Z(n15939) );
  XOR U17936 ( .A(n15940), .B(n15939), .Z(n15942) );
  AND U17937 ( .A(x[482]), .B(y[7834]), .Z(n15941) );
  XOR U17938 ( .A(n15942), .B(n15941), .Z(n16007) );
  XOR U17939 ( .A(n16008), .B(n16007), .Z(n16009) );
  XNOR U17940 ( .A(n16010), .B(n16009), .Z(n15986) );
  NANDN U17941 ( .A(n15839), .B(n15838), .Z(n15843) );
  NANDN U17942 ( .A(n15841), .B(n15840), .Z(n15842) );
  NAND U17943 ( .A(n15843), .B(n15842), .Z(n16006) );
  AND U17944 ( .A(x[483]), .B(y[7833]), .Z(n15965) );
  XOR U17945 ( .A(n15966), .B(n15965), .Z(n15968) );
  AND U17946 ( .A(x[503]), .B(y[7813]), .Z(n15967) );
  XOR U17947 ( .A(n15968), .B(n15967), .Z(n16004) );
  AND U17948 ( .A(x[485]), .B(y[7831]), .Z(n15952) );
  AND U17949 ( .A(x[501]), .B(y[7815]), .Z(n15951) );
  XOR U17950 ( .A(n15952), .B(n15951), .Z(n15954) );
  AND U17951 ( .A(x[500]), .B(y[7816]), .Z(n15953) );
  XOR U17952 ( .A(n15954), .B(n15953), .Z(n16003) );
  XOR U17953 ( .A(n16004), .B(n16003), .Z(n16005) );
  XNOR U17954 ( .A(n16006), .B(n16005), .Z(n15984) );
  NANDN U17955 ( .A(n15845), .B(n15844), .Z(n15849) );
  NANDN U17956 ( .A(n15847), .B(n15846), .Z(n15848) );
  NAND U17957 ( .A(n15849), .B(n15848), .Z(n15937) );
  ANDN U17958 ( .B(o[155]), .A(n15850), .Z(n15928) );
  AND U17959 ( .A(x[480]), .B(y[7836]), .Z(n15926) );
  AND U17960 ( .A(x[508]), .B(y[7808]), .Z(n15925) );
  XOR U17961 ( .A(n15926), .B(n15925), .Z(n15927) );
  XOR U17962 ( .A(n15928), .B(n15927), .Z(n15936) );
  NAND U17963 ( .A(y[7826]), .B(x[490]), .Z(n15851) );
  XNOR U17964 ( .A(n15852), .B(n15851), .Z(n15932) );
  AND U17965 ( .A(x[489]), .B(y[7827]), .Z(n15931) );
  XOR U17966 ( .A(n15932), .B(n15931), .Z(n15935) );
  XOR U17967 ( .A(n15936), .B(n15935), .Z(n15938) );
  XOR U17968 ( .A(n15937), .B(n15938), .Z(n16002) );
  NANDN U17969 ( .A(n15854), .B(n15853), .Z(n15858) );
  NAND U17970 ( .A(n15856), .B(n15855), .Z(n15857) );
  NAND U17971 ( .A(n15858), .B(n15857), .Z(n15999) );
  NANDN U17972 ( .A(n15860), .B(n15859), .Z(n15864) );
  NANDN U17973 ( .A(n15862), .B(n15861), .Z(n15863) );
  NAND U17974 ( .A(n15864), .B(n15863), .Z(n16000) );
  XOR U17975 ( .A(n15999), .B(n16000), .Z(n16001) );
  XNOR U17976 ( .A(n16002), .B(n16001), .Z(n15983) );
  XOR U17977 ( .A(n15984), .B(n15983), .Z(n15985) );
  XOR U17978 ( .A(n15986), .B(n15985), .Z(n16015) );
  XNOR U17979 ( .A(n16016), .B(n16015), .Z(n16017) );
  XOR U17980 ( .A(n16018), .B(n16017), .Z(n16013) );
  XNOR U17981 ( .A(n16011), .B(n16012), .Z(n16014) );
  XOR U17982 ( .A(n16013), .B(n16014), .Z(n15902) );
  NANDN U17983 ( .A(n15874), .B(n15873), .Z(n15878) );
  NAND U17984 ( .A(n15876), .B(n15875), .Z(n15877) );
  NAND U17985 ( .A(n15878), .B(n15877), .Z(n15909) );
  NAND U17986 ( .A(n15880), .B(n15879), .Z(n15884) );
  NAND U17987 ( .A(n15882), .B(n15881), .Z(n15883) );
  NAND U17988 ( .A(n15884), .B(n15883), .Z(n15907) );
  NAND U17989 ( .A(n15886), .B(n15885), .Z(n15890) );
  NANDN U17990 ( .A(n15888), .B(n15887), .Z(n15889) );
  AND U17991 ( .A(n15890), .B(n15889), .Z(n15908) );
  XNOR U17992 ( .A(n15907), .B(n15908), .Z(n15910) );
  XNOR U17993 ( .A(n15903), .B(n15904), .Z(n16030) );
  XNOR U17994 ( .A(n16031), .B(n16030), .Z(n16024) );
  NAND U17995 ( .A(n15895), .B(n15894), .Z(n15899) );
  NANDN U17996 ( .A(n15897), .B(n15896), .Z(n15898) );
  NAND U17997 ( .A(n15899), .B(n15898), .Z(n16022) );
  IV U17998 ( .A(n16022), .Z(n16021) );
  XOR U17999 ( .A(n16023), .B(n16021), .Z(n15900) );
  XNOR U18000 ( .A(n16024), .B(n15900), .Z(N317) );
  NANDN U18001 ( .A(n15902), .B(n15901), .Z(n15906) );
  NANDN U18002 ( .A(n15904), .B(n15903), .Z(n15905) );
  NAND U18003 ( .A(n15906), .B(n15905), .Z(n16044) );
  NAND U18004 ( .A(n15908), .B(n15907), .Z(n15912) );
  NANDN U18005 ( .A(n15910), .B(n15909), .Z(n15911) );
  NAND U18006 ( .A(n15912), .B(n15911), .Z(n16042) );
  XOR U18007 ( .A(n16180), .B(n16181), .Z(n16182) );
  AND U18008 ( .A(x[490]), .B(y[7828]), .Z(n15929) );
  NAND U18009 ( .A(n15930), .B(n15929), .Z(n15934) );
  NAND U18010 ( .A(n15932), .B(n15931), .Z(n15933) );
  NAND U18011 ( .A(n15934), .B(n15933), .Z(n16172) );
  AND U18012 ( .A(x[502]), .B(y[7815]), .Z(n16147) );
  AND U18013 ( .A(x[492]), .B(y[7825]), .Z(n16331) );
  AND U18014 ( .A(x[481]), .B(y[7836]), .Z(n16145) );
  XOR U18015 ( .A(n16331), .B(n16145), .Z(n16146) );
  XOR U18016 ( .A(n16147), .B(n16146), .Z(n16171) );
  AND U18017 ( .A(x[495]), .B(y[7822]), .Z(n16139) );
  XOR U18018 ( .A(n16249), .B(n16139), .Z(n16140) );
  XOR U18019 ( .A(n16141), .B(n16140), .Z(n16170) );
  XOR U18020 ( .A(n16171), .B(n16170), .Z(n16173) );
  XNOR U18021 ( .A(n16172), .B(n16173), .Z(n16183) );
  XOR U18022 ( .A(n16182), .B(n16183), .Z(n16161) );
  XNOR U18023 ( .A(n16161), .B(n16160), .Z(n16163) );
  XOR U18024 ( .A(n16162), .B(n16163), .Z(n16155) );
  XOR U18025 ( .A(n16176), .B(n16177), .Z(n16178) );
  AND U18026 ( .A(x[483]), .B(y[7834]), .Z(n16125) );
  AND U18027 ( .A(x[497]), .B(y[7820]), .Z(n16124) );
  XOR U18028 ( .A(n16125), .B(n16124), .Z(n16127) );
  AND U18029 ( .A(x[491]), .B(y[7826]), .Z(n16126) );
  XOR U18030 ( .A(n16127), .B(n16126), .Z(n16109) );
  AND U18031 ( .A(x[493]), .B(y[7824]), .Z(n16130) );
  AND U18032 ( .A(x[504]), .B(y[7813]), .Z(n16396) );
  XOR U18033 ( .A(n16130), .B(n16396), .Z(n16132) );
  AND U18034 ( .A(x[503]), .B(y[7814]), .Z(n16131) );
  XOR U18035 ( .A(n16132), .B(n16131), .Z(n16108) );
  XOR U18036 ( .A(n16109), .B(n16108), .Z(n16110) );
  XNOR U18037 ( .A(n16111), .B(n16110), .Z(n16179) );
  XNOR U18038 ( .A(n16178), .B(n16179), .Z(n16078) );
  AND U18039 ( .A(x[482]), .B(y[7835]), .Z(n16100) );
  XOR U18040 ( .A(n16101), .B(n16100), .Z(n16102) );
  XOR U18041 ( .A(n16103), .B(n16102), .Z(n16114) );
  AND U18042 ( .A(n15955), .B(o[156]), .Z(n16107) );
  AND U18043 ( .A(x[496]), .B(y[7821]), .Z(n16105) );
  AND U18044 ( .A(x[507]), .B(y[7810]), .Z(n16104) );
  XOR U18045 ( .A(n16105), .B(n16104), .Z(n16106) );
  XOR U18046 ( .A(n16107), .B(n16106), .Z(n16113) );
  XOR U18047 ( .A(n16114), .B(n16113), .Z(n16116) );
  XOR U18048 ( .A(n16115), .B(n16116), .Z(n16076) );
  AND U18049 ( .A(x[505]), .B(y[7812]), .Z(n16138) );
  AND U18050 ( .A(x[506]), .B(y[7811]), .Z(n16135) );
  XOR U18051 ( .A(n16136), .B(n16135), .Z(n16137) );
  XOR U18052 ( .A(n16138), .B(n16137), .Z(n16165) );
  AND U18053 ( .A(x[508]), .B(y[7809]), .Z(n16144) );
  XOR U18054 ( .A(o[157]), .B(n16144), .Z(n16187) );
  AND U18055 ( .A(x[480]), .B(y[7837]), .Z(n16185) );
  AND U18056 ( .A(x[509]), .B(y[7808]), .Z(n16184) );
  XOR U18057 ( .A(n16185), .B(n16184), .Z(n16186) );
  XOR U18058 ( .A(n16187), .B(n16186), .Z(n16164) );
  XOR U18059 ( .A(n16165), .B(n16164), .Z(n16166) );
  XOR U18060 ( .A(n16167), .B(n16166), .Z(n16075) );
  XNOR U18061 ( .A(n16076), .B(n16075), .Z(n16077) );
  XNOR U18062 ( .A(n16078), .B(n16077), .Z(n16083) );
  AND U18063 ( .A(x[485]), .B(y[7832]), .Z(n16097) );
  AND U18064 ( .A(x[484]), .B(y[7833]), .Z(n16095) );
  AND U18065 ( .A(x[490]), .B(y[7827]), .Z(n16094) );
  XOR U18066 ( .A(n16095), .B(n16094), .Z(n16096) );
  XOR U18067 ( .A(n16097), .B(n16096), .Z(n16194) );
  AND U18068 ( .A(x[488]), .B(y[7829]), .Z(n16119) );
  AND U18069 ( .A(y[7831]), .B(x[486]), .Z(n15960) );
  AND U18070 ( .A(y[7830]), .B(x[487]), .Z(n15959) );
  XOR U18071 ( .A(n15960), .B(n15959), .Z(n16118) );
  XOR U18072 ( .A(n16119), .B(n16118), .Z(n16192) );
  AND U18073 ( .A(x[489]), .B(y[7828]), .Z(n16262) );
  XOR U18074 ( .A(n16192), .B(n16262), .Z(n16193) );
  XOR U18075 ( .A(n16194), .B(n16193), .Z(n16090) );
  XNOR U18076 ( .A(n16087), .B(n16088), .Z(n16091) );
  XNOR U18077 ( .A(n16090), .B(n16091), .Z(n16082) );
  XOR U18078 ( .A(n16082), .B(n16081), .Z(n16084) );
  XOR U18079 ( .A(n16083), .B(n16084), .Z(n16152) );
  XOR U18080 ( .A(n16152), .B(n16153), .Z(n16156) );
  XOR U18081 ( .A(n16155), .B(n16156), .Z(n16067) );
  XNOR U18082 ( .A(n16068), .B(n16067), .Z(n16070) );
  NANDN U18083 ( .A(n15978), .B(n15977), .Z(n15982) );
  NANDN U18084 ( .A(n15980), .B(n15979), .Z(n15981) );
  AND U18085 ( .A(n15982), .B(n15981), .Z(n16061) );
  NAND U18086 ( .A(n15984), .B(n15983), .Z(n15988) );
  NAND U18087 ( .A(n15986), .B(n15985), .Z(n15987) );
  AND U18088 ( .A(n15988), .B(n15987), .Z(n16060) );
  XNOR U18089 ( .A(n16061), .B(n16060), .Z(n16063) );
  NANDN U18090 ( .A(n15990), .B(n15989), .Z(n15994) );
  NANDN U18091 ( .A(n15992), .B(n15991), .Z(n15993) );
  NAND U18092 ( .A(n15994), .B(n15993), .Z(n16055) );
  XOR U18093 ( .A(n16148), .B(n16149), .Z(n16151) );
  XOR U18094 ( .A(n16150), .B(n16151), .Z(n16053) );
  XOR U18095 ( .A(n16052), .B(n16053), .Z(n16056) );
  XOR U18096 ( .A(n16055), .B(n16056), .Z(n16062) );
  XOR U18097 ( .A(n16063), .B(n16062), .Z(n16069) );
  XOR U18098 ( .A(n16070), .B(n16069), .Z(n16051) );
  NANDN U18099 ( .A(n16016), .B(n16015), .Z(n16020) );
  NANDN U18100 ( .A(n16018), .B(n16017), .Z(n16019) );
  AND U18101 ( .A(n16020), .B(n16019), .Z(n16049) );
  XOR U18102 ( .A(n16048), .B(n16049), .Z(n16050) );
  XOR U18103 ( .A(n16051), .B(n16050), .Z(n16043) );
  XNOR U18104 ( .A(n16042), .B(n16043), .Z(n16045) );
  XOR U18105 ( .A(n16044), .B(n16045), .Z(n16038) );
  OR U18106 ( .A(n16023), .B(n16021), .Z(n16027) );
  ANDN U18107 ( .B(n16023), .A(n16022), .Z(n16025) );
  OR U18108 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U18109 ( .A(n16027), .B(n16026), .Z(n16037) );
  NANDN U18110 ( .A(n16029), .B(n16028), .Z(n16033) );
  NAND U18111 ( .A(n16031), .B(n16030), .Z(n16032) );
  NAND U18112 ( .A(n16033), .B(n16032), .Z(n16036) );
  IV U18113 ( .A(n16036), .Z(n16035) );
  XOR U18114 ( .A(n16037), .B(n16035), .Z(n16034) );
  XNOR U18115 ( .A(n16038), .B(n16034), .Z(N318) );
  OR U18116 ( .A(n16037), .B(n16035), .Z(n16041) );
  ANDN U18117 ( .B(n16037), .A(n16036), .Z(n16039) );
  OR U18118 ( .A(n16039), .B(n16038), .Z(n16040) );
  AND U18119 ( .A(n16041), .B(n16040), .Z(n16486) );
  NAND U18120 ( .A(n16043), .B(n16042), .Z(n16047) );
  NANDN U18121 ( .A(n16045), .B(n16044), .Z(n16046) );
  NAND U18122 ( .A(n16047), .B(n16046), .Z(n16487) );
  IV U18123 ( .A(n16052), .Z(n16054) );
  NANDN U18124 ( .A(n16054), .B(n16053), .Z(n16059) );
  IV U18125 ( .A(n16055), .Z(n16057) );
  NANDN U18126 ( .A(n16057), .B(n16056), .Z(n16058) );
  AND U18127 ( .A(n16059), .B(n16058), .Z(n16471) );
  NANDN U18128 ( .A(n16061), .B(n16060), .Z(n16066) );
  IV U18129 ( .A(n16062), .Z(n16064) );
  NANDN U18130 ( .A(n16064), .B(n16063), .Z(n16065) );
  AND U18131 ( .A(n16066), .B(n16065), .Z(n16472) );
  NANDN U18132 ( .A(n16068), .B(n16067), .Z(n16073) );
  IV U18133 ( .A(n16069), .Z(n16071) );
  NANDN U18134 ( .A(n16071), .B(n16070), .Z(n16072) );
  NAND U18135 ( .A(n16073), .B(n16072), .Z(n16473) );
  IV U18136 ( .A(n16473), .Z(n16074) );
  XOR U18137 ( .A(n16472), .B(n16074), .Z(n16470) );
  XOR U18138 ( .A(n16471), .B(n16470), .Z(n16481) );
  NANDN U18139 ( .A(n16076), .B(n16075), .Z(n16080) );
  NANDN U18140 ( .A(n16078), .B(n16077), .Z(n16079) );
  AND U18141 ( .A(n16080), .B(n16079), .Z(n16462) );
  NANDN U18142 ( .A(n16082), .B(n16081), .Z(n16086) );
  NANDN U18143 ( .A(n16084), .B(n16083), .Z(n16085) );
  AND U18144 ( .A(n16086), .B(n16085), .Z(n16455) );
  IV U18145 ( .A(n16087), .Z(n16089) );
  NANDN U18146 ( .A(n16089), .B(n16088), .Z(n16093) );
  NANDN U18147 ( .A(n16091), .B(n16090), .Z(n16092) );
  AND U18148 ( .A(n16093), .B(n16092), .Z(n16197) );
  NAND U18149 ( .A(n16095), .B(n16094), .Z(n16099) );
  NAND U18150 ( .A(n16097), .B(n16096), .Z(n16098) );
  NAND U18151 ( .A(n16099), .B(n16098), .Z(n16212) );
  AND U18152 ( .A(x[486]), .B(y[7832]), .Z(n16326) );
  AND U18153 ( .A(x[485]), .B(y[7833]), .Z(n16328) );
  AND U18154 ( .A(x[499]), .B(y[7819]), .Z(n16327) );
  XOR U18155 ( .A(n16328), .B(n16327), .Z(n16325) );
  XNOR U18156 ( .A(n16326), .B(n16325), .Z(n16363) );
  AND U18157 ( .A(x[484]), .B(y[7834]), .Z(n16253) );
  AND U18158 ( .A(x[483]), .B(y[7835]), .Z(n16255) );
  AND U18159 ( .A(x[498]), .B(y[7820]), .Z(n16254) );
  XOR U18160 ( .A(n16255), .B(n16254), .Z(n16252) );
  XOR U18161 ( .A(n16253), .B(n16252), .Z(n16366) );
  XOR U18162 ( .A(n16363), .B(n16364), .Z(n16211) );
  XOR U18163 ( .A(n16212), .B(n16211), .Z(n16210) );
  XOR U18164 ( .A(n16210), .B(n16209), .Z(n16200) );
  IV U18165 ( .A(n16200), .Z(n16112) );
  XNOR U18166 ( .A(n16112), .B(n16199), .Z(n16198) );
  XOR U18167 ( .A(n16197), .B(n16198), .Z(n16456) );
  AND U18168 ( .A(x[487]), .B(y[7831]), .Z(n16248) );
  NAND U18169 ( .A(n16117), .B(n16248), .Z(n16121) );
  NAND U18170 ( .A(n16119), .B(n16118), .Z(n16120) );
  AND U18171 ( .A(n16121), .B(n16120), .Z(n16215) );
  AND U18172 ( .A(x[501]), .B(y[7817]), .Z(n16123) );
  AND U18173 ( .A(y[7816]), .B(x[502]), .Z(n16122) );
  XOR U18174 ( .A(n16123), .B(n16122), .Z(n16247) );
  XOR U18175 ( .A(n16248), .B(n16247), .Z(n16218) );
  AND U18176 ( .A(x[497]), .B(y[7821]), .Z(n16322) );
  AND U18177 ( .A(x[482]), .B(y[7836]), .Z(n16320) );
  AND U18178 ( .A(x[506]), .B(y[7812]), .Z(n16319) );
  XOR U18179 ( .A(n16320), .B(n16319), .Z(n16321) );
  XNOR U18180 ( .A(n16322), .B(n16321), .Z(n16217) );
  XNOR U18181 ( .A(n16215), .B(n16216), .Z(n16204) );
  NAND U18182 ( .A(n16125), .B(n16124), .Z(n16129) );
  NAND U18183 ( .A(n16127), .B(n16126), .Z(n16128) );
  AND U18184 ( .A(n16129), .B(n16128), .Z(n16227) );
  AND U18185 ( .A(x[480]), .B(y[7838]), .Z(n16242) );
  AND U18186 ( .A(x[509]), .B(y[7809]), .Z(n16265) );
  XOR U18187 ( .A(o[158]), .B(n16265), .Z(n16244) );
  AND U18188 ( .A(x[510]), .B(y[7808]), .Z(n16243) );
  XOR U18189 ( .A(n16244), .B(n16243), .Z(n16241) );
  XOR U18190 ( .A(n16242), .B(n16241), .Z(n16230) );
  AND U18191 ( .A(x[500]), .B(y[7818]), .Z(n16381) );
  XOR U18192 ( .A(n16382), .B(n16381), .Z(n16380) );
  AND U18193 ( .A(x[488]), .B(y[7830]), .Z(n16379) );
  XNOR U18194 ( .A(n16380), .B(n16379), .Z(n16229) );
  XNOR U18195 ( .A(n16227), .B(n16228), .Z(n16206) );
  NAND U18196 ( .A(n16130), .B(n16396), .Z(n16134) );
  NAND U18197 ( .A(n16132), .B(n16131), .Z(n16133) );
  NAND U18198 ( .A(n16134), .B(n16133), .Z(n16205) );
  XNOR U18199 ( .A(n16204), .B(n16203), .Z(n16441) );
  XOR U18200 ( .A(n16440), .B(n16441), .Z(n16438) );
  AND U18201 ( .A(x[503]), .B(y[7815]), .Z(n16394) );
  AND U18202 ( .A(x[504]), .B(y[7814]), .Z(n16143) );
  AND U18203 ( .A(y[7813]), .B(x[505]), .Z(n16142) );
  XOR U18204 ( .A(n16143), .B(n16142), .Z(n16393) );
  XOR U18205 ( .A(n16394), .B(n16393), .Z(n16224) );
  AND U18206 ( .A(x[508]), .B(y[7810]), .Z(n16376) );
  AND U18207 ( .A(x[496]), .B(y[7822]), .Z(n16375) );
  XOR U18208 ( .A(n16376), .B(n16375), .Z(n16373) );
  XNOR U18209 ( .A(n16374), .B(n16373), .Z(n16223) );
  XOR U18210 ( .A(n16221), .B(n16222), .Z(n16238) );
  XNOR U18211 ( .A(n16238), .B(n16237), .Z(n16236) );
  XOR U18212 ( .A(n16235), .B(n16236), .Z(n16439) );
  XNOR U18213 ( .A(n16438), .B(n16439), .Z(n16457) );
  XOR U18214 ( .A(n16456), .B(n16457), .Z(n16454) );
  XOR U18215 ( .A(n16455), .B(n16454), .Z(n16464) );
  IV U18216 ( .A(n16152), .Z(n16154) );
  NANDN U18217 ( .A(n16154), .B(n16153), .Z(n16159) );
  IV U18218 ( .A(n16155), .Z(n16157) );
  NANDN U18219 ( .A(n16157), .B(n16156), .Z(n16158) );
  AND U18220 ( .A(n16159), .B(n16158), .Z(n16453) );
  NAND U18221 ( .A(n16165), .B(n16164), .Z(n16169) );
  NANDN U18222 ( .A(n16167), .B(n16166), .Z(n16168) );
  AND U18223 ( .A(n16169), .B(n16168), .Z(n16420) );
  NAND U18224 ( .A(n16171), .B(n16170), .Z(n16175) );
  NAND U18225 ( .A(n16173), .B(n16172), .Z(n16174) );
  AND U18226 ( .A(n16175), .B(n16174), .Z(n16421) );
  XOR U18227 ( .A(n16420), .B(n16419), .Z(n16435) );
  AND U18228 ( .A(y[7826]), .B(x[492]), .Z(n16188) );
  XOR U18229 ( .A(n16189), .B(n16188), .Z(n16333) );
  XOR U18230 ( .A(n16334), .B(n16333), .Z(n16260) );
  AND U18231 ( .A(y[7829]), .B(x[489]), .Z(n16191) );
  NAND U18232 ( .A(y[7828]), .B(x[490]), .Z(n16190) );
  XOR U18233 ( .A(n16191), .B(n16190), .Z(n16261) );
  XNOR U18234 ( .A(n16260), .B(n16261), .Z(n16360) );
  AND U18235 ( .A(x[507]), .B(y[7811]), .Z(n16389) );
  NAND U18236 ( .A(x[481]), .B(y[7837]), .Z(n16390) );
  XOR U18237 ( .A(n16388), .B(n16387), .Z(n16359) );
  XOR U18238 ( .A(n16360), .B(n16359), .Z(n16357) );
  XOR U18239 ( .A(n16358), .B(n16357), .Z(n16415) );
  NAND U18240 ( .A(n16192), .B(n16262), .Z(n16196) );
  NAND U18241 ( .A(n16194), .B(n16193), .Z(n16195) );
  AND U18242 ( .A(n16196), .B(n16195), .Z(n16416) );
  XOR U18243 ( .A(n16415), .B(n16416), .Z(n16413) );
  XNOR U18244 ( .A(n16414), .B(n16413), .Z(n16434) );
  XOR U18245 ( .A(n16432), .B(n16431), .Z(n16452) );
  XOR U18246 ( .A(n16451), .B(n16450), .Z(n16480) );
  XOR U18247 ( .A(n16479), .B(n16478), .Z(n16484) );
  XNOR U18248 ( .A(n16485), .B(n16484), .Z(N319) );
  NANDN U18249 ( .A(n16198), .B(n16197), .Z(n16202) );
  NANDN U18250 ( .A(n16200), .B(n16199), .Z(n16201) );
  AND U18251 ( .A(n16202), .B(n16201), .Z(n16461) );
  NANDN U18252 ( .A(n16204), .B(n16203), .Z(n16208) );
  NANDN U18253 ( .A(n16206), .B(n16205), .Z(n16207) );
  AND U18254 ( .A(n16208), .B(n16207), .Z(n16449) );
  NAND U18255 ( .A(n16210), .B(n16209), .Z(n16214) );
  NAND U18256 ( .A(n16212), .B(n16211), .Z(n16213) );
  AND U18257 ( .A(n16214), .B(n16213), .Z(n16430) );
  NANDN U18258 ( .A(n16216), .B(n16215), .Z(n16220) );
  NANDN U18259 ( .A(n16218), .B(n16217), .Z(n16219) );
  AND U18260 ( .A(n16220), .B(n16219), .Z(n16412) );
  NANDN U18261 ( .A(n16222), .B(n16221), .Z(n16226) );
  NANDN U18262 ( .A(n16224), .B(n16223), .Z(n16225) );
  AND U18263 ( .A(n16226), .B(n16225), .Z(n16234) );
  NANDN U18264 ( .A(n16228), .B(n16227), .Z(n16232) );
  NANDN U18265 ( .A(n16230), .B(n16229), .Z(n16231) );
  NAND U18266 ( .A(n16232), .B(n16231), .Z(n16233) );
  XNOR U18267 ( .A(n16234), .B(n16233), .Z(n16410) );
  NANDN U18268 ( .A(n16236), .B(n16235), .Z(n16240) );
  NAND U18269 ( .A(n16238), .B(n16237), .Z(n16239) );
  AND U18270 ( .A(n16240), .B(n16239), .Z(n16408) );
  NAND U18271 ( .A(n16242), .B(n16241), .Z(n16246) );
  NAND U18272 ( .A(n16244), .B(n16243), .Z(n16245) );
  AND U18273 ( .A(n16246), .B(n16245), .Z(n16318) );
  NAND U18274 ( .A(n16248), .B(n16247), .Z(n16251) );
  AND U18275 ( .A(x[502]), .B(y[7817]), .Z(n16284) );
  NAND U18276 ( .A(n16249), .B(n16284), .Z(n16250) );
  AND U18277 ( .A(n16251), .B(n16250), .Z(n16259) );
  NAND U18278 ( .A(n16253), .B(n16252), .Z(n16257) );
  NAND U18279 ( .A(n16255), .B(n16254), .Z(n16256) );
  NAND U18280 ( .A(n16257), .B(n16256), .Z(n16258) );
  XNOR U18281 ( .A(n16259), .B(n16258), .Z(n16316) );
  NANDN U18282 ( .A(n16261), .B(n16260), .Z(n16264) );
  AND U18283 ( .A(x[490]), .B(y[7829]), .Z(n16279) );
  NAND U18284 ( .A(n16262), .B(n16279), .Z(n16263) );
  AND U18285 ( .A(n16264), .B(n16263), .Z(n16314) );
  AND U18286 ( .A(n16265), .B(o[158]), .Z(n16270) );
  AND U18287 ( .A(y[7808]), .B(x[511]), .Z(n16268) );
  XNOR U18288 ( .A(n16266), .B(o[159]), .Z(n16267) );
  XNOR U18289 ( .A(n16268), .B(n16267), .Z(n16269) );
  XOR U18290 ( .A(n16270), .B(n16269), .Z(n16273) );
  XNOR U18291 ( .A(n16271), .B(n16332), .Z(n16272) );
  XNOR U18292 ( .A(n16273), .B(n16272), .Z(n16312) );
  AND U18293 ( .A(y[7836]), .B(x[483]), .Z(n16275) );
  NAND U18294 ( .A(y[7813]), .B(x[506]), .Z(n16274) );
  XNOR U18295 ( .A(n16275), .B(n16274), .Z(n16283) );
  AND U18296 ( .A(y[7821]), .B(x[498]), .Z(n16281) );
  AND U18297 ( .A(y[7828]), .B(x[491]), .Z(n16277) );
  NAND U18298 ( .A(y[7827]), .B(x[492]), .Z(n16276) );
  XNOR U18299 ( .A(n16277), .B(n16276), .Z(n16278) );
  XNOR U18300 ( .A(n16279), .B(n16278), .Z(n16280) );
  XNOR U18301 ( .A(n16281), .B(n16280), .Z(n16282) );
  XOR U18302 ( .A(n16283), .B(n16282), .Z(n16286) );
  AND U18303 ( .A(x[505]), .B(y[7814]), .Z(n16395) );
  XNOR U18304 ( .A(n16284), .B(n16395), .Z(n16285) );
  XNOR U18305 ( .A(n16286), .B(n16285), .Z(n16302) );
  AND U18306 ( .A(y[7810]), .B(x[509]), .Z(n16288) );
  NAND U18307 ( .A(y[7819]), .B(x[500]), .Z(n16287) );
  XNOR U18308 ( .A(n16288), .B(n16287), .Z(n16292) );
  AND U18309 ( .A(y[7809]), .B(x[510]), .Z(n16290) );
  NAND U18310 ( .A(y[7825]), .B(x[494]), .Z(n16289) );
  XNOR U18311 ( .A(n16290), .B(n16289), .Z(n16291) );
  XOR U18312 ( .A(n16292), .B(n16291), .Z(n16300) );
  AND U18313 ( .A(y[7811]), .B(x[508]), .Z(n16294) );
  NAND U18314 ( .A(y[7839]), .B(x[480]), .Z(n16293) );
  XNOR U18315 ( .A(n16294), .B(n16293), .Z(n16298) );
  AND U18316 ( .A(y[7823]), .B(x[496]), .Z(n16296) );
  NAND U18317 ( .A(y[7838]), .B(x[481]), .Z(n16295) );
  XNOR U18318 ( .A(n16296), .B(n16295), .Z(n16297) );
  XNOR U18319 ( .A(n16298), .B(n16297), .Z(n16299) );
  XNOR U18320 ( .A(n16300), .B(n16299), .Z(n16301) );
  XOR U18321 ( .A(n16302), .B(n16301), .Z(n16310) );
  AND U18322 ( .A(y[7833]), .B(x[486]), .Z(n16304) );
  NAND U18323 ( .A(y[7835]), .B(x[484]), .Z(n16303) );
  XNOR U18324 ( .A(n16304), .B(n16303), .Z(n16308) );
  AND U18325 ( .A(y[7837]), .B(x[482]), .Z(n16306) );
  NAND U18326 ( .A(y[7822]), .B(x[497]), .Z(n16305) );
  XNOR U18327 ( .A(n16306), .B(n16305), .Z(n16307) );
  XNOR U18328 ( .A(n16308), .B(n16307), .Z(n16309) );
  XNOR U18329 ( .A(n16310), .B(n16309), .Z(n16311) );
  XNOR U18330 ( .A(n16312), .B(n16311), .Z(n16313) );
  XNOR U18331 ( .A(n16314), .B(n16313), .Z(n16315) );
  XNOR U18332 ( .A(n16316), .B(n16315), .Z(n16317) );
  XNOR U18333 ( .A(n16318), .B(n16317), .Z(n16406) );
  AND U18334 ( .A(n16320), .B(n16319), .Z(n16324) );
  AND U18335 ( .A(n16322), .B(n16321), .Z(n16323) );
  NOR U18336 ( .A(n16324), .B(n16323), .Z(n16356) );
  NAND U18337 ( .A(n16326), .B(n16325), .Z(n16330) );
  NAND U18338 ( .A(n16328), .B(n16327), .Z(n16329) );
  AND U18339 ( .A(n16330), .B(n16329), .Z(n16338) );
  NAND U18340 ( .A(n16332), .B(n16331), .Z(n16336) );
  NAND U18341 ( .A(n16334), .B(n16333), .Z(n16335) );
  AND U18342 ( .A(n16336), .B(n16335), .Z(n16337) );
  XNOR U18343 ( .A(n16338), .B(n16337), .Z(n16354) );
  AND U18344 ( .A(y[7820]), .B(x[499]), .Z(n16340) );
  NAND U18345 ( .A(y[7831]), .B(x[488]), .Z(n16339) );
  XNOR U18346 ( .A(n16340), .B(n16339), .Z(n16344) );
  AND U18347 ( .A(y[7818]), .B(x[501]), .Z(n16342) );
  NAND U18348 ( .A(y[7830]), .B(x[489]), .Z(n16341) );
  XNOR U18349 ( .A(n16342), .B(n16341), .Z(n16343) );
  XOR U18350 ( .A(n16344), .B(n16343), .Z(n16352) );
  AND U18351 ( .A(y[7812]), .B(x[507]), .Z(n16346) );
  NAND U18352 ( .A(y[7816]), .B(x[503]), .Z(n16345) );
  XNOR U18353 ( .A(n16346), .B(n16345), .Z(n16350) );
  AND U18354 ( .A(y[7834]), .B(x[485]), .Z(n16348) );
  NAND U18355 ( .A(y[7832]), .B(x[487]), .Z(n16347) );
  XNOR U18356 ( .A(n16348), .B(n16347), .Z(n16349) );
  XNOR U18357 ( .A(n16350), .B(n16349), .Z(n16351) );
  XNOR U18358 ( .A(n16352), .B(n16351), .Z(n16353) );
  XOR U18359 ( .A(n16354), .B(n16353), .Z(n16355) );
  XNOR U18360 ( .A(n16356), .B(n16355), .Z(n16372) );
  NANDN U18361 ( .A(n16358), .B(n16357), .Z(n16362) );
  NAND U18362 ( .A(n16360), .B(n16359), .Z(n16361) );
  AND U18363 ( .A(n16362), .B(n16361), .Z(n16370) );
  NANDN U18364 ( .A(n16364), .B(n16363), .Z(n16368) );
  NANDN U18365 ( .A(n16366), .B(n16365), .Z(n16367) );
  NAND U18366 ( .A(n16368), .B(n16367), .Z(n16369) );
  XNOR U18367 ( .A(n16370), .B(n16369), .Z(n16371) );
  XOR U18368 ( .A(n16372), .B(n16371), .Z(n16404) );
  NAND U18369 ( .A(n16374), .B(n16373), .Z(n16378) );
  NAND U18370 ( .A(n16376), .B(n16375), .Z(n16377) );
  AND U18371 ( .A(n16378), .B(n16377), .Z(n16386) );
  NAND U18372 ( .A(n16380), .B(n16379), .Z(n16384) );
  NAND U18373 ( .A(n16382), .B(n16381), .Z(n16383) );
  NAND U18374 ( .A(n16384), .B(n16383), .Z(n16385) );
  XNOR U18375 ( .A(n16386), .B(n16385), .Z(n16402) );
  NAND U18376 ( .A(n16388), .B(n16387), .Z(n16392) );
  NANDN U18377 ( .A(n16390), .B(n16389), .Z(n16391) );
  AND U18378 ( .A(n16392), .B(n16391), .Z(n16400) );
  NAND U18379 ( .A(n16394), .B(n16393), .Z(n16398) );
  NAND U18380 ( .A(n16396), .B(n16395), .Z(n16397) );
  NAND U18381 ( .A(n16398), .B(n16397), .Z(n16399) );
  XNOR U18382 ( .A(n16400), .B(n16399), .Z(n16401) );
  XNOR U18383 ( .A(n16402), .B(n16401), .Z(n16403) );
  XNOR U18384 ( .A(n16404), .B(n16403), .Z(n16405) );
  XNOR U18385 ( .A(n16406), .B(n16405), .Z(n16407) );
  XNOR U18386 ( .A(n16408), .B(n16407), .Z(n16409) );
  XNOR U18387 ( .A(n16410), .B(n16409), .Z(n16411) );
  XNOR U18388 ( .A(n16412), .B(n16411), .Z(n16428) );
  NAND U18389 ( .A(n16414), .B(n16413), .Z(n16418) );
  NAND U18390 ( .A(n16416), .B(n16415), .Z(n16417) );
  AND U18391 ( .A(n16418), .B(n16417), .Z(n16426) );
  NAND U18392 ( .A(n16420), .B(n16419), .Z(n16424) );
  NANDN U18393 ( .A(n16422), .B(n16421), .Z(n16423) );
  NAND U18394 ( .A(n16424), .B(n16423), .Z(n16425) );
  XNOR U18395 ( .A(n16426), .B(n16425), .Z(n16427) );
  XNOR U18396 ( .A(n16428), .B(n16427), .Z(n16429) );
  XNOR U18397 ( .A(n16430), .B(n16429), .Z(n16447) );
  IV U18398 ( .A(n16431), .Z(n16433) );
  NANDN U18399 ( .A(n16433), .B(n16432), .Z(n16437) );
  NANDN U18400 ( .A(n16435), .B(n16434), .Z(n16436) );
  AND U18401 ( .A(n16437), .B(n16436), .Z(n16445) );
  NANDN U18402 ( .A(n16439), .B(n16438), .Z(n16443) );
  NAND U18403 ( .A(n16441), .B(n16440), .Z(n16442) );
  NAND U18404 ( .A(n16443), .B(n16442), .Z(n16444) );
  XNOR U18405 ( .A(n16445), .B(n16444), .Z(n16446) );
  XNOR U18406 ( .A(n16447), .B(n16446), .Z(n16448) );
  XNOR U18407 ( .A(n16449), .B(n16448), .Z(n16459) );
  XNOR U18408 ( .A(n16459), .B(n16458), .Z(n16460) );
  XNOR U18409 ( .A(n16461), .B(n16460), .Z(n16469) );
  NANDN U18410 ( .A(n16463), .B(n16462), .Z(n16467) );
  ANDN U18411 ( .B(n16463), .A(n16462), .Z(n16465) );
  NANDN U18412 ( .A(n16465), .B(n16464), .Z(n16466) );
  NAND U18413 ( .A(n16467), .B(n16466), .Z(n16468) );
  XNOR U18414 ( .A(n16469), .B(n16468), .Z(n16477) );
  NAND U18415 ( .A(n16471), .B(n16470), .Z(n16475) );
  NANDN U18416 ( .A(n16473), .B(n16472), .Z(n16474) );
  NAND U18417 ( .A(n16475), .B(n16474), .Z(n16476) );
  XNOR U18418 ( .A(n16477), .B(n16476), .Z(n16493) );
  NANDN U18419 ( .A(n16479), .B(n16478), .Z(n16483) );
  NANDN U18420 ( .A(n16481), .B(n16480), .Z(n16482) );
  AND U18421 ( .A(n16483), .B(n16482), .Z(n16491) );
  NAND U18422 ( .A(n16485), .B(n16484), .Z(n16489) );
  NANDN U18423 ( .A(n16487), .B(n16486), .Z(n16488) );
  NAND U18424 ( .A(n16489), .B(n16488), .Z(n16490) );
  XNOR U18425 ( .A(n16491), .B(n16490), .Z(n16492) );
  XNOR U18426 ( .A(n16493), .B(n16492), .Z(N320) );
  AND U18427 ( .A(x[480]), .B(y[7840]), .Z(n17140) );
  XOR U18428 ( .A(n17140), .B(o[160]), .Z(N353) );
  AND U18429 ( .A(x[481]), .B(y[7840]), .Z(n16502) );
  AND U18430 ( .A(x[480]), .B(y[7841]), .Z(n16501) );
  XNOR U18431 ( .A(n16501), .B(o[161]), .Z(n16494) );
  XNOR U18432 ( .A(n16502), .B(n16494), .Z(n16496) );
  NAND U18433 ( .A(n17140), .B(o[160]), .Z(n16495) );
  XNOR U18434 ( .A(n16496), .B(n16495), .Z(N354) );
  NANDN U18435 ( .A(n16502), .B(n16494), .Z(n16498) );
  NAND U18436 ( .A(n16496), .B(n16495), .Z(n16497) );
  AND U18437 ( .A(n16498), .B(n16497), .Z(n16508) );
  AND U18438 ( .A(x[480]), .B(y[7842]), .Z(n16516) );
  XNOR U18439 ( .A(n16516), .B(o[162]), .Z(n16507) );
  XNOR U18440 ( .A(n16508), .B(n16507), .Z(n16510) );
  AND U18441 ( .A(y[7840]), .B(x[482]), .Z(n16500) );
  NAND U18442 ( .A(y[7841]), .B(x[481]), .Z(n16499) );
  XNOR U18443 ( .A(n16500), .B(n16499), .Z(n16504) );
  AND U18444 ( .A(n16501), .B(o[161]), .Z(n16503) );
  XNOR U18445 ( .A(n16504), .B(n16503), .Z(n16509) );
  XNOR U18446 ( .A(n16510), .B(n16509), .Z(N355) );
  AND U18447 ( .A(x[482]), .B(y[7841]), .Z(n16513) );
  IV U18448 ( .A(n16513), .Z(n16521) );
  NANDN U18449 ( .A(n16521), .B(n16502), .Z(n16506) );
  NAND U18450 ( .A(n16504), .B(n16503), .Z(n16505) );
  AND U18451 ( .A(n16506), .B(n16505), .Z(n16529) );
  NANDN U18452 ( .A(n16508), .B(n16507), .Z(n16512) );
  NAND U18453 ( .A(n16510), .B(n16509), .Z(n16511) );
  AND U18454 ( .A(n16512), .B(n16511), .Z(n16528) );
  XNOR U18455 ( .A(n16529), .B(n16528), .Z(n16531) );
  AND U18456 ( .A(x[481]), .B(y[7842]), .Z(n16619) );
  XOR U18457 ( .A(o[163]), .B(n16513), .Z(n16525) );
  XOR U18458 ( .A(n16619), .B(n16525), .Z(n16527) );
  AND U18459 ( .A(y[7840]), .B(x[483]), .Z(n16515) );
  NAND U18460 ( .A(y[7843]), .B(x[480]), .Z(n16514) );
  XNOR U18461 ( .A(n16515), .B(n16514), .Z(n16518) );
  AND U18462 ( .A(n16516), .B(o[162]), .Z(n16517) );
  XOR U18463 ( .A(n16518), .B(n16517), .Z(n16526) );
  XOR U18464 ( .A(n16527), .B(n16526), .Z(n16530) );
  XOR U18465 ( .A(n16531), .B(n16530), .Z(N356) );
  AND U18466 ( .A(x[483]), .B(y[7843]), .Z(n16576) );
  NAND U18467 ( .A(n17140), .B(n16576), .Z(n16520) );
  NAND U18468 ( .A(n16518), .B(n16517), .Z(n16519) );
  NAND U18469 ( .A(n16520), .B(n16519), .Z(n16550) );
  ANDN U18470 ( .B(o[163]), .A(n16521), .Z(n16544) );
  AND U18471 ( .A(x[480]), .B(y[7844]), .Z(n16523) );
  AND U18472 ( .A(y[7840]), .B(x[484]), .Z(n16522) );
  XOR U18473 ( .A(n16523), .B(n16522), .Z(n16543) );
  XOR U18474 ( .A(n16544), .B(n16543), .Z(n16549) );
  AND U18475 ( .A(y[7842]), .B(x[482]), .Z(n16655) );
  NAND U18476 ( .A(y[7843]), .B(x[481]), .Z(n16524) );
  XNOR U18477 ( .A(n16655), .B(n16524), .Z(n16542) );
  AND U18478 ( .A(x[483]), .B(y[7841]), .Z(n16537) );
  XOR U18479 ( .A(n16537), .B(o[164]), .Z(n16541) );
  XOR U18480 ( .A(n16542), .B(n16541), .Z(n16548) );
  XOR U18481 ( .A(n16549), .B(n16548), .Z(n16551) );
  XNOR U18482 ( .A(n16550), .B(n16551), .Z(n16547) );
  NANDN U18483 ( .A(n16529), .B(n16528), .Z(n16533) );
  NAND U18484 ( .A(n16531), .B(n16530), .Z(n16532) );
  NAND U18485 ( .A(n16533), .B(n16532), .Z(n16546) );
  XOR U18486 ( .A(n16545), .B(n16546), .Z(n16534) );
  XNOR U18487 ( .A(n16547), .B(n16534), .Z(N357) );
  AND U18488 ( .A(y[7840]), .B(x[485]), .Z(n16536) );
  NAND U18489 ( .A(y[7845]), .B(x[480]), .Z(n16535) );
  XNOR U18490 ( .A(n16536), .B(n16535), .Z(n16569) );
  AND U18491 ( .A(n16537), .B(o[164]), .Z(n16568) );
  XOR U18492 ( .A(n16569), .B(n16568), .Z(n16567) );
  NAND U18493 ( .A(x[482]), .B(y[7843]), .Z(n16628) );
  AND U18494 ( .A(y[7842]), .B(x[483]), .Z(n16539) );
  NAND U18495 ( .A(y[7844]), .B(x[481]), .Z(n16538) );
  XNOR U18496 ( .A(n16539), .B(n16538), .Z(n16563) );
  AND U18497 ( .A(x[484]), .B(y[7841]), .Z(n16572) );
  XOR U18498 ( .A(n16572), .B(o[165]), .Z(n16562) );
  XOR U18499 ( .A(n16563), .B(n16562), .Z(n16566) );
  XOR U18500 ( .A(n16628), .B(n16566), .Z(n16540) );
  XNOR U18501 ( .A(n16567), .B(n16540), .Z(n16558) );
  AND U18502 ( .A(x[484]), .B(y[7844]), .Z(n17340) );
  XOR U18503 ( .A(n16555), .B(n16556), .Z(n16557) );
  XNOR U18504 ( .A(n16558), .B(n16557), .Z(n16561) );
  NAND U18505 ( .A(n16549), .B(n16548), .Z(n16553) );
  NAND U18506 ( .A(n16551), .B(n16550), .Z(n16552) );
  NAND U18507 ( .A(n16553), .B(n16552), .Z(n16559) );
  XNOR U18508 ( .A(n16560), .B(n16559), .Z(n16554) );
  XNOR U18509 ( .A(n16561), .B(n16554), .Z(N358) );
  AND U18510 ( .A(x[483]), .B(y[7844]), .Z(n16630) );
  NAND U18511 ( .A(n16630), .B(n16619), .Z(n16565) );
  NAND U18512 ( .A(n16563), .B(n16562), .Z(n16564) );
  NAND U18513 ( .A(n16565), .B(n16564), .Z(n16604) );
  XOR U18514 ( .A(n16604), .B(n16603), .Z(n16606) );
  AND U18515 ( .A(x[485]), .B(y[7845]), .Z(n16803) );
  NAND U18516 ( .A(n17140), .B(n16803), .Z(n16571) );
  NAND U18517 ( .A(n16569), .B(n16568), .Z(n16570) );
  NAND U18518 ( .A(n16571), .B(n16570), .Z(n16579) );
  AND U18519 ( .A(n16572), .B(o[165]), .Z(n16587) );
  AND U18520 ( .A(y[7840]), .B(x[486]), .Z(n16574) );
  AND U18521 ( .A(y[7846]), .B(x[480]), .Z(n16573) );
  XOR U18522 ( .A(n16574), .B(n16573), .Z(n16586) );
  XOR U18523 ( .A(n16587), .B(n16586), .Z(n16580) );
  XOR U18524 ( .A(n16579), .B(n16580), .Z(n16582) );
  NAND U18525 ( .A(y[7844]), .B(x[482]), .Z(n16575) );
  XNOR U18526 ( .A(n16576), .B(n16575), .Z(n16591) );
  AND U18527 ( .A(x[481]), .B(y[7845]), .Z(n16854) );
  NAND U18528 ( .A(y[7842]), .B(x[484]), .Z(n16577) );
  XNOR U18529 ( .A(n16854), .B(n16577), .Z(n16595) );
  AND U18530 ( .A(x[485]), .B(y[7841]), .Z(n16600) );
  XOR U18531 ( .A(o[166]), .B(n16600), .Z(n16594) );
  XOR U18532 ( .A(n16595), .B(n16594), .Z(n16590) );
  XOR U18533 ( .A(n16591), .B(n16590), .Z(n16581) );
  XOR U18534 ( .A(n16582), .B(n16581), .Z(n16605) );
  XOR U18535 ( .A(n16606), .B(n16605), .Z(n16611) );
  XOR U18536 ( .A(n16609), .B(n16611), .Z(n16578) );
  XOR U18537 ( .A(n16610), .B(n16578), .Z(N359) );
  NAND U18538 ( .A(n16580), .B(n16579), .Z(n16584) );
  NAND U18539 ( .A(n16582), .B(n16581), .Z(n16583) );
  AND U18540 ( .A(n16584), .B(n16583), .Z(n16651) );
  AND U18541 ( .A(y[7842]), .B(x[485]), .Z(n16711) );
  NAND U18542 ( .A(y[7846]), .B(x[481]), .Z(n16585) );
  XNOR U18543 ( .A(n16711), .B(n16585), .Z(n16621) );
  AND U18544 ( .A(x[486]), .B(y[7841]), .Z(n16625) );
  XOR U18545 ( .A(o[167]), .B(n16625), .Z(n16620) );
  XOR U18546 ( .A(n16621), .B(n16620), .Z(n16640) );
  AND U18547 ( .A(x[486]), .B(y[7846]), .Z(n16874) );
  NAND U18548 ( .A(n17140), .B(n16874), .Z(n16589) );
  NAND U18549 ( .A(n16587), .B(n16586), .Z(n16588) );
  AND U18550 ( .A(n16589), .B(n16588), .Z(n16639) );
  NANDN U18551 ( .A(n16628), .B(n16630), .Z(n16593) );
  NAND U18552 ( .A(n16591), .B(n16590), .Z(n16592) );
  AND U18553 ( .A(n16593), .B(n16592), .Z(n16641) );
  XOR U18554 ( .A(n16642), .B(n16641), .Z(n16649) );
  AND U18555 ( .A(x[484]), .B(y[7845]), .Z(n17145) );
  NAND U18556 ( .A(n17145), .B(n16619), .Z(n16597) );
  NAND U18557 ( .A(n16595), .B(n16594), .Z(n16596) );
  AND U18558 ( .A(n16597), .B(n16596), .Z(n16616) );
  AND U18559 ( .A(y[7845]), .B(x[482]), .Z(n16599) );
  NAND U18560 ( .A(y[7843]), .B(x[484]), .Z(n16598) );
  XNOR U18561 ( .A(n16599), .B(n16598), .Z(n16629) );
  XNOR U18562 ( .A(n16630), .B(n16629), .Z(n16614) );
  AND U18563 ( .A(o[166]), .B(n16600), .Z(n16634) );
  AND U18564 ( .A(y[7840]), .B(x[487]), .Z(n16602) );
  NAND U18565 ( .A(y[7847]), .B(x[480]), .Z(n16601) );
  XNOR U18566 ( .A(n16602), .B(n16601), .Z(n16633) );
  XNOR U18567 ( .A(n16634), .B(n16633), .Z(n16613) );
  XOR U18568 ( .A(n16614), .B(n16613), .Z(n16615) );
  XOR U18569 ( .A(n16616), .B(n16615), .Z(n16648) );
  XOR U18570 ( .A(n16649), .B(n16648), .Z(n16650) );
  XOR U18571 ( .A(n16651), .B(n16650), .Z(n16647) );
  NAND U18572 ( .A(n16604), .B(n16603), .Z(n16608) );
  NAND U18573 ( .A(n16606), .B(n16605), .Z(n16607) );
  NAND U18574 ( .A(n16608), .B(n16607), .Z(n16646) );
  XOR U18575 ( .A(n16646), .B(n16645), .Z(n16612) );
  XNOR U18576 ( .A(n16647), .B(n16612), .Z(N360) );
  NAND U18577 ( .A(n16614), .B(n16613), .Z(n16618) );
  NAND U18578 ( .A(n16616), .B(n16615), .Z(n16617) );
  AND U18579 ( .A(n16618), .B(n16617), .Z(n16688) );
  AND U18580 ( .A(x[485]), .B(y[7846]), .Z(n16795) );
  NAND U18581 ( .A(n16795), .B(n16619), .Z(n16623) );
  NAND U18582 ( .A(n16621), .B(n16620), .Z(n16622) );
  NAND U18583 ( .A(n16623), .B(n16622), .Z(n16686) );
  AND U18584 ( .A(y[7843]), .B(x[485]), .Z(n17250) );
  NAND U18585 ( .A(y[7847]), .B(x[481]), .Z(n16624) );
  XNOR U18586 ( .A(n17250), .B(n16624), .Z(n16676) );
  AND U18587 ( .A(o[167]), .B(n16625), .Z(n16675) );
  XOR U18588 ( .A(n16676), .B(n16675), .Z(n16661) );
  NAND U18589 ( .A(x[483]), .B(y[7845]), .Z(n17458) );
  AND U18590 ( .A(y[7842]), .B(x[486]), .Z(n16627) );
  NAND U18591 ( .A(y[7846]), .B(x[482]), .Z(n16626) );
  XNOR U18592 ( .A(n16627), .B(n16626), .Z(n16656) );
  XNOR U18593 ( .A(n17340), .B(n16656), .Z(n16659) );
  XOR U18594 ( .A(n17458), .B(n16659), .Z(n16660) );
  XOR U18595 ( .A(n16661), .B(n16660), .Z(n16685) );
  XOR U18596 ( .A(n16686), .B(n16685), .Z(n16687) );
  XOR U18597 ( .A(n16688), .B(n16687), .Z(n16701) );
  NANDN U18598 ( .A(n16628), .B(n17145), .Z(n16632) );
  NAND U18599 ( .A(n16630), .B(n16629), .Z(n16631) );
  NAND U18600 ( .A(n16632), .B(n16631), .Z(n16682) );
  AND U18601 ( .A(x[487]), .B(y[7847]), .Z(n17013) );
  NAND U18602 ( .A(n17140), .B(n17013), .Z(n16636) );
  NAND U18603 ( .A(n16634), .B(n16633), .Z(n16635) );
  NAND U18604 ( .A(n16636), .B(n16635), .Z(n16680) );
  AND U18605 ( .A(y[7840]), .B(x[488]), .Z(n16638) );
  NAND U18606 ( .A(y[7848]), .B(x[480]), .Z(n16637) );
  XNOR U18607 ( .A(n16638), .B(n16637), .Z(n16666) );
  AND U18608 ( .A(x[487]), .B(y[7841]), .Z(n16671) );
  XOR U18609 ( .A(o[168]), .B(n16671), .Z(n16665) );
  XOR U18610 ( .A(n16666), .B(n16665), .Z(n16679) );
  XOR U18611 ( .A(n16680), .B(n16679), .Z(n16681) );
  XOR U18612 ( .A(n16682), .B(n16681), .Z(n16699) );
  NANDN U18613 ( .A(n16640), .B(n16639), .Z(n16644) );
  NAND U18614 ( .A(n16642), .B(n16641), .Z(n16643) );
  NAND U18615 ( .A(n16644), .B(n16643), .Z(n16698) );
  NAND U18616 ( .A(n16649), .B(n16648), .Z(n16653) );
  NAND U18617 ( .A(n16651), .B(n16650), .Z(n16652) );
  AND U18618 ( .A(n16653), .B(n16652), .Z(n16692) );
  IV U18619 ( .A(n16692), .Z(n16691) );
  XOR U18620 ( .A(n16693), .B(n16691), .Z(n16654) );
  XNOR U18621 ( .A(n16694), .B(n16654), .Z(N361) );
  NAND U18622 ( .A(n16874), .B(n16655), .Z(n16658) );
  NAND U18623 ( .A(n17340), .B(n16656), .Z(n16657) );
  AND U18624 ( .A(n16658), .B(n16657), .Z(n16706) );
  NAND U18625 ( .A(n17458), .B(n16659), .Z(n16663) );
  NANDN U18626 ( .A(n16661), .B(n16660), .Z(n16662) );
  AND U18627 ( .A(n16663), .B(n16662), .Z(n16705) );
  AND U18628 ( .A(x[488]), .B(y[7848]), .Z(n16664) );
  NAND U18629 ( .A(n16664), .B(n17140), .Z(n16668) );
  NAND U18630 ( .A(n16666), .B(n16665), .Z(n16667) );
  AND U18631 ( .A(n16668), .B(n16667), .Z(n16740) );
  AND U18632 ( .A(y[7844]), .B(x[485]), .Z(n16670) );
  NAND U18633 ( .A(y[7842]), .B(x[487]), .Z(n16669) );
  XNOR U18634 ( .A(n16670), .B(n16669), .Z(n16713) );
  AND U18635 ( .A(o[168]), .B(n16671), .Z(n16712) );
  XNOR U18636 ( .A(n16713), .B(n16712), .Z(n16738) );
  AND U18637 ( .A(y[7840]), .B(x[489]), .Z(n16673) );
  NAND U18638 ( .A(y[7849]), .B(x[480]), .Z(n16672) );
  XNOR U18639 ( .A(n16673), .B(n16672), .Z(n16720) );
  NAND U18640 ( .A(x[488]), .B(y[7841]), .Z(n16727) );
  XNOR U18641 ( .A(n16720), .B(n16719), .Z(n16737) );
  XOR U18642 ( .A(n16738), .B(n16737), .Z(n16739) );
  XNOR U18643 ( .A(n16740), .B(n16739), .Z(n16734) );
  AND U18644 ( .A(y[7843]), .B(x[486]), .Z(n17084) );
  NAND U18645 ( .A(y[7848]), .B(x[481]), .Z(n16674) );
  XNOR U18646 ( .A(n17084), .B(n16674), .Z(n16724) );
  XNOR U18647 ( .A(n17145), .B(n16724), .Z(n16744) );
  NAND U18648 ( .A(x[482]), .B(y[7847]), .Z(n17381) );
  AND U18649 ( .A(x[483]), .B(y[7846]), .Z(n17094) );
  XNOR U18650 ( .A(n17381), .B(n17094), .Z(n16743) );
  XNOR U18651 ( .A(n16744), .B(n16743), .Z(n16732) );
  NAND U18652 ( .A(x[485]), .B(y[7847]), .Z(n16920) );
  AND U18653 ( .A(x[481]), .B(y[7843]), .Z(n16723) );
  NANDN U18654 ( .A(n16920), .B(n16723), .Z(n16678) );
  NAND U18655 ( .A(n16676), .B(n16675), .Z(n16677) );
  NAND U18656 ( .A(n16678), .B(n16677), .Z(n16731) );
  XOR U18657 ( .A(n16732), .B(n16731), .Z(n16733) );
  XOR U18658 ( .A(n16734), .B(n16733), .Z(n16707) );
  XOR U18659 ( .A(n16708), .B(n16707), .Z(n16757) );
  NAND U18660 ( .A(n16680), .B(n16679), .Z(n16684) );
  NAND U18661 ( .A(n16682), .B(n16681), .Z(n16683) );
  NAND U18662 ( .A(n16684), .B(n16683), .Z(n16755) );
  NAND U18663 ( .A(n16686), .B(n16685), .Z(n16690) );
  NAND U18664 ( .A(n16688), .B(n16687), .Z(n16689) );
  NAND U18665 ( .A(n16690), .B(n16689), .Z(n16754) );
  XOR U18666 ( .A(n16755), .B(n16754), .Z(n16756) );
  XNOR U18667 ( .A(n16757), .B(n16756), .Z(n16750) );
  OR U18668 ( .A(n16693), .B(n16691), .Z(n16697) );
  ANDN U18669 ( .B(n16693), .A(n16692), .Z(n16695) );
  OR U18670 ( .A(n16695), .B(n16694), .Z(n16696) );
  AND U18671 ( .A(n16697), .B(n16696), .Z(n16749) );
  NANDN U18672 ( .A(n16699), .B(n16698), .Z(n16703) );
  NANDN U18673 ( .A(n16701), .B(n16700), .Z(n16702) );
  AND U18674 ( .A(n16703), .B(n16702), .Z(n16748) );
  IV U18675 ( .A(n16748), .Z(n16747) );
  XOR U18676 ( .A(n16749), .B(n16747), .Z(n16704) );
  XNOR U18677 ( .A(n16750), .B(n16704), .Z(N362) );
  NANDN U18678 ( .A(n16706), .B(n16705), .Z(n16710) );
  NAND U18679 ( .A(n16708), .B(n16707), .Z(n16709) );
  AND U18680 ( .A(n16710), .B(n16709), .Z(n16816) );
  AND U18681 ( .A(x[487]), .B(y[7844]), .Z(n16797) );
  NAND U18682 ( .A(n16797), .B(n16711), .Z(n16715) );
  NAND U18683 ( .A(n16713), .B(n16712), .Z(n16714) );
  AND U18684 ( .A(n16715), .B(n16714), .Z(n16810) );
  AND U18685 ( .A(y[7843]), .B(x[487]), .Z(n16717) );
  NAND U18686 ( .A(y[7846]), .B(x[484]), .Z(n16716) );
  XNOR U18687 ( .A(n16717), .B(n16716), .Z(n16781) );
  AND U18688 ( .A(x[486]), .B(y[7844]), .Z(n16780) );
  XOR U18689 ( .A(n16781), .B(n16780), .Z(n16808) );
  AND U18690 ( .A(x[488]), .B(y[7842]), .Z(n16977) );
  AND U18691 ( .A(x[489]), .B(y[7841]), .Z(n16791) );
  XOR U18692 ( .A(n16791), .B(o[170]), .Z(n16802) );
  XOR U18693 ( .A(n16977), .B(n16802), .Z(n16804) );
  XNOR U18694 ( .A(n16804), .B(n16803), .Z(n16807) );
  XNOR U18695 ( .A(n16810), .B(n16809), .Z(n16770) );
  AND U18696 ( .A(x[489]), .B(y[7849]), .Z(n16718) );
  NAND U18697 ( .A(n17140), .B(n16718), .Z(n16722) );
  NAND U18698 ( .A(n16720), .B(n16719), .Z(n16721) );
  NAND U18699 ( .A(n16722), .B(n16721), .Z(n16768) );
  AND U18700 ( .A(x[486]), .B(y[7848]), .Z(n17004) );
  NAND U18701 ( .A(n17004), .B(n16723), .Z(n16726) );
  NAND U18702 ( .A(n17145), .B(n16724), .Z(n16725) );
  NAND U18703 ( .A(n16726), .B(n16725), .Z(n16775) );
  ANDN U18704 ( .B(o[169]), .A(n16727), .Z(n16786) );
  AND U18705 ( .A(y[7840]), .B(x[490]), .Z(n16729) );
  AND U18706 ( .A(y[7850]), .B(x[480]), .Z(n16728) );
  XOR U18707 ( .A(n16729), .B(n16728), .Z(n16785) );
  XOR U18708 ( .A(n16786), .B(n16785), .Z(n16774) );
  AND U18709 ( .A(y[7847]), .B(x[483]), .Z(n17697) );
  NAND U18710 ( .A(y[7849]), .B(x[481]), .Z(n16730) );
  XNOR U18711 ( .A(n17697), .B(n16730), .Z(n16799) );
  AND U18712 ( .A(x[482]), .B(y[7848]), .Z(n16798) );
  XOR U18713 ( .A(n16799), .B(n16798), .Z(n16773) );
  XOR U18714 ( .A(n16774), .B(n16773), .Z(n16776) );
  XOR U18715 ( .A(n16775), .B(n16776), .Z(n16767) );
  XOR U18716 ( .A(n16768), .B(n16767), .Z(n16769) );
  XNOR U18717 ( .A(n16770), .B(n16769), .Z(n16814) );
  NAND U18718 ( .A(n16732), .B(n16731), .Z(n16736) );
  NAND U18719 ( .A(n16734), .B(n16733), .Z(n16735) );
  AND U18720 ( .A(n16736), .B(n16735), .Z(n16764) );
  NAND U18721 ( .A(n16738), .B(n16737), .Z(n16742) );
  NAND U18722 ( .A(n16740), .B(n16739), .Z(n16741) );
  AND U18723 ( .A(n16742), .B(n16741), .Z(n16761) );
  NAND U18724 ( .A(n16744), .B(n16743), .Z(n16746) );
  ANDN U18725 ( .B(n17381), .A(n17094), .Z(n16745) );
  ANDN U18726 ( .B(n16746), .A(n16745), .Z(n16762) );
  XOR U18727 ( .A(n16761), .B(n16762), .Z(n16763) );
  XOR U18728 ( .A(n16764), .B(n16763), .Z(n16813) );
  XOR U18729 ( .A(n16814), .B(n16813), .Z(n16815) );
  XNOR U18730 ( .A(n16816), .B(n16815), .Z(n16822) );
  OR U18731 ( .A(n16749), .B(n16747), .Z(n16753) );
  ANDN U18732 ( .B(n16749), .A(n16748), .Z(n16751) );
  OR U18733 ( .A(n16751), .B(n16750), .Z(n16752) );
  AND U18734 ( .A(n16753), .B(n16752), .Z(n16820) );
  NAND U18735 ( .A(n16755), .B(n16754), .Z(n16759) );
  NAND U18736 ( .A(n16757), .B(n16756), .Z(n16758) );
  AND U18737 ( .A(n16759), .B(n16758), .Z(n16821) );
  IV U18738 ( .A(n16821), .Z(n16819) );
  XOR U18739 ( .A(n16820), .B(n16819), .Z(n16760) );
  XNOR U18740 ( .A(n16822), .B(n16760), .Z(N363) );
  NAND U18741 ( .A(n16762), .B(n16761), .Z(n16766) );
  NANDN U18742 ( .A(n16764), .B(n16763), .Z(n16765) );
  NAND U18743 ( .A(n16766), .B(n16765), .Z(n16885) );
  NAND U18744 ( .A(n16768), .B(n16767), .Z(n16772) );
  NAND U18745 ( .A(n16770), .B(n16769), .Z(n16771) );
  NAND U18746 ( .A(n16772), .B(n16771), .Z(n16883) );
  NAND U18747 ( .A(n16774), .B(n16773), .Z(n16778) );
  NAND U18748 ( .A(n16776), .B(n16775), .Z(n16777) );
  NAND U18749 ( .A(n16778), .B(n16777), .Z(n16840) );
  AND U18750 ( .A(x[487]), .B(y[7846]), .Z(n16915) );
  AND U18751 ( .A(x[484]), .B(y[7843]), .Z(n16779) );
  NAND U18752 ( .A(n16915), .B(n16779), .Z(n16783) );
  NAND U18753 ( .A(n16781), .B(n16780), .Z(n16782) );
  NAND U18754 ( .A(n16783), .B(n16782), .Z(n16838) );
  AND U18755 ( .A(x[490]), .B(y[7850]), .Z(n16784) );
  NAND U18756 ( .A(n16784), .B(n17140), .Z(n16788) );
  NAND U18757 ( .A(n16786), .B(n16785), .Z(n16787) );
  NAND U18758 ( .A(n16788), .B(n16787), .Z(n16834) );
  AND U18759 ( .A(y[7840]), .B(x[491]), .Z(n16790) );
  NAND U18760 ( .A(y[7851]), .B(x[480]), .Z(n16789) );
  XNOR U18761 ( .A(n16790), .B(n16789), .Z(n16864) );
  AND U18762 ( .A(n16791), .B(o[170]), .Z(n16865) );
  XOR U18763 ( .A(n16864), .B(n16865), .Z(n16833) );
  AND U18764 ( .A(y[7845]), .B(x[486]), .Z(n16793) );
  NAND U18765 ( .A(y[7850]), .B(x[481]), .Z(n16792) );
  XNOR U18766 ( .A(n16793), .B(n16792), .Z(n16856) );
  AND U18767 ( .A(x[490]), .B(y[7841]), .Z(n16875) );
  XOR U18768 ( .A(o[171]), .B(n16875), .Z(n16855) );
  XOR U18769 ( .A(n16856), .B(n16855), .Z(n16832) );
  XOR U18770 ( .A(n16833), .B(n16832), .Z(n16835) );
  XOR U18771 ( .A(n16834), .B(n16835), .Z(n16839) );
  XOR U18772 ( .A(n16838), .B(n16839), .Z(n16841) );
  XNOR U18773 ( .A(n16840), .B(n16841), .Z(n16878) );
  AND U18774 ( .A(x[483]), .B(y[7848]), .Z(n17820) );
  NAND U18775 ( .A(y[7849]), .B(x[482]), .Z(n16794) );
  XNOR U18776 ( .A(n16795), .B(n16794), .Z(n16851) );
  AND U18777 ( .A(x[484]), .B(y[7847]), .Z(n16850) );
  XNOR U18778 ( .A(n16851), .B(n16850), .Z(n16827) );
  XNOR U18779 ( .A(n17820), .B(n16827), .Z(n16828) );
  NAND U18780 ( .A(y[7842]), .B(x[489]), .Z(n16796) );
  XNOR U18781 ( .A(n16797), .B(n16796), .Z(n16869) );
  AND U18782 ( .A(x[488]), .B(y[7843]), .Z(n16870) );
  XOR U18783 ( .A(n16869), .B(n16870), .Z(n16829) );
  AND U18784 ( .A(x[483]), .B(y[7849]), .Z(n16911) );
  AND U18785 ( .A(x[481]), .B(y[7847]), .Z(n17135) );
  NAND U18786 ( .A(n16911), .B(n17135), .Z(n16801) );
  NAND U18787 ( .A(n16799), .B(n16798), .Z(n16800) );
  NAND U18788 ( .A(n16801), .B(n16800), .Z(n16845) );
  NAND U18789 ( .A(n16977), .B(n16802), .Z(n16806) );
  NAND U18790 ( .A(n16804), .B(n16803), .Z(n16805) );
  NAND U18791 ( .A(n16806), .B(n16805), .Z(n16844) );
  XOR U18792 ( .A(n16845), .B(n16844), .Z(n16846) );
  NANDN U18793 ( .A(n16808), .B(n16807), .Z(n16812) );
  NAND U18794 ( .A(n16810), .B(n16809), .Z(n16811) );
  NAND U18795 ( .A(n16812), .B(n16811), .Z(n16876) );
  XOR U18796 ( .A(n16878), .B(n16879), .Z(n16882) );
  XOR U18797 ( .A(n16883), .B(n16882), .Z(n16884) );
  XOR U18798 ( .A(n16885), .B(n16884), .Z(n16890) );
  NAND U18799 ( .A(n16814), .B(n16813), .Z(n16818) );
  NAND U18800 ( .A(n16816), .B(n16815), .Z(n16817) );
  NAND U18801 ( .A(n16818), .B(n16817), .Z(n16888) );
  NANDN U18802 ( .A(n16819), .B(n16820), .Z(n16825) );
  NOR U18803 ( .A(n16821), .B(n16820), .Z(n16823) );
  OR U18804 ( .A(n16823), .B(n16822), .Z(n16824) );
  AND U18805 ( .A(n16825), .B(n16824), .Z(n16889) );
  XOR U18806 ( .A(n16888), .B(n16889), .Z(n16826) );
  XNOR U18807 ( .A(n16890), .B(n16826), .Z(N364) );
  NANDN U18808 ( .A(n17820), .B(n16827), .Z(n16831) );
  NANDN U18809 ( .A(n16829), .B(n16828), .Z(n16830) );
  NAND U18810 ( .A(n16831), .B(n16830), .Z(n16892) );
  NAND U18811 ( .A(n16833), .B(n16832), .Z(n16837) );
  NAND U18812 ( .A(n16835), .B(n16834), .Z(n16836) );
  AND U18813 ( .A(n16837), .B(n16836), .Z(n16893) );
  XOR U18814 ( .A(n16892), .B(n16893), .Z(n16895) );
  NAND U18815 ( .A(n16839), .B(n16838), .Z(n16843) );
  NAND U18816 ( .A(n16841), .B(n16840), .Z(n16842) );
  AND U18817 ( .A(n16843), .B(n16842), .Z(n16894) );
  XOR U18818 ( .A(n16895), .B(n16894), .Z(n16960) );
  NAND U18819 ( .A(n16845), .B(n16844), .Z(n16849) );
  NANDN U18820 ( .A(n16847), .B(n16846), .Z(n16848) );
  NAND U18821 ( .A(n16849), .B(n16848), .Z(n16951) );
  AND U18822 ( .A(x[482]), .B(y[7846]), .Z(n17558) );
  AND U18823 ( .A(x[485]), .B(y[7849]), .Z(n17372) );
  NAND U18824 ( .A(n17558), .B(n17372), .Z(n16853) );
  NAND U18825 ( .A(n16851), .B(n16850), .Z(n16852) );
  AND U18826 ( .A(n16853), .B(n16852), .Z(n16899) );
  AND U18827 ( .A(x[486]), .B(y[7850]), .Z(n17152) );
  NAND U18828 ( .A(n17152), .B(n16854), .Z(n16858) );
  NAND U18829 ( .A(n16856), .B(n16855), .Z(n16857) );
  NAND U18830 ( .A(n16858), .B(n16857), .Z(n16898) );
  AND U18831 ( .A(x[489]), .B(y[7843]), .Z(n17553) );
  AND U18832 ( .A(x[490]), .B(y[7842]), .Z(n17596) );
  NAND U18833 ( .A(y[7848]), .B(x[484]), .Z(n16859) );
  XNOR U18834 ( .A(n17596), .B(n16859), .Z(n16942) );
  XOR U18835 ( .A(n17553), .B(n16942), .Z(n16921) );
  NAND U18836 ( .A(x[487]), .B(y[7845]), .Z(n16919) );
  XOR U18837 ( .A(n16920), .B(n16919), .Z(n16922) );
  AND U18838 ( .A(y[7840]), .B(x[492]), .Z(n16861) );
  NAND U18839 ( .A(y[7852]), .B(x[480]), .Z(n16860) );
  XNOR U18840 ( .A(n16861), .B(n16860), .Z(n16936) );
  AND U18841 ( .A(x[491]), .B(y[7841]), .Z(n16916) );
  XOR U18842 ( .A(o[172]), .B(n16916), .Z(n16935) );
  XOR U18843 ( .A(n16936), .B(n16935), .Z(n16905) );
  AND U18844 ( .A(y[7850]), .B(x[482]), .Z(n16863) );
  NAND U18845 ( .A(y[7844]), .B(x[488]), .Z(n16862) );
  XNOR U18846 ( .A(n16863), .B(n16862), .Z(n16910) );
  XOR U18847 ( .A(n16910), .B(n16911), .Z(n16904) );
  XOR U18848 ( .A(n16905), .B(n16904), .Z(n16907) );
  XOR U18849 ( .A(n16906), .B(n16907), .Z(n16900) );
  XOR U18850 ( .A(n16901), .B(n16900), .Z(n16949) );
  AND U18851 ( .A(x[491]), .B(y[7851]), .Z(n17918) );
  NAND U18852 ( .A(n17918), .B(n17140), .Z(n16867) );
  NAND U18853 ( .A(n16865), .B(n16864), .Z(n16866) );
  NAND U18854 ( .A(n16867), .B(n16866), .Z(n16928) );
  AND U18855 ( .A(x[487]), .B(y[7842]), .Z(n17070) );
  AND U18856 ( .A(x[489]), .B(y[7844]), .Z(n16868) );
  NAND U18857 ( .A(n17070), .B(n16868), .Z(n16872) );
  NAND U18858 ( .A(n16870), .B(n16869), .Z(n16871) );
  NAND U18859 ( .A(n16872), .B(n16871), .Z(n16926) );
  NAND U18860 ( .A(y[7851]), .B(x[481]), .Z(n16873) );
  XNOR U18861 ( .A(n16874), .B(n16873), .Z(n16932) );
  AND U18862 ( .A(o[171]), .B(n16875), .Z(n16931) );
  XOR U18863 ( .A(n16932), .B(n16931), .Z(n16925) );
  XOR U18864 ( .A(n16926), .B(n16925), .Z(n16927) );
  XNOR U18865 ( .A(n16928), .B(n16927), .Z(n16950) );
  XNOR U18866 ( .A(n16949), .B(n16950), .Z(n16952) );
  XOR U18867 ( .A(n16951), .B(n16952), .Z(n16959) );
  NANDN U18868 ( .A(n16877), .B(n16876), .Z(n16881) );
  NANDN U18869 ( .A(n16879), .B(n16878), .Z(n16880) );
  NAND U18870 ( .A(n16881), .B(n16880), .Z(n16958) );
  XNOR U18871 ( .A(n16960), .B(n16961), .Z(n16957) );
  NAND U18872 ( .A(n16883), .B(n16882), .Z(n16887) );
  NAND U18873 ( .A(n16885), .B(n16884), .Z(n16886) );
  NAND U18874 ( .A(n16887), .B(n16886), .Z(n16956) );
  XOR U18875 ( .A(n16956), .B(n16955), .Z(n16891) );
  XNOR U18876 ( .A(n16957), .B(n16891), .Z(N365) );
  NAND U18877 ( .A(n16893), .B(n16892), .Z(n16897) );
  NAND U18878 ( .A(n16895), .B(n16894), .Z(n16896) );
  NAND U18879 ( .A(n16897), .B(n16896), .Z(n17041) );
  NANDN U18880 ( .A(n16899), .B(n16898), .Z(n16903) );
  NAND U18881 ( .A(n16901), .B(n16900), .Z(n16902) );
  AND U18882 ( .A(n16903), .B(n16902), .Z(n17021) );
  NAND U18883 ( .A(n16905), .B(n16904), .Z(n16909) );
  NAND U18884 ( .A(n16907), .B(n16906), .Z(n16908) );
  NAND U18885 ( .A(n16909), .B(n16908), .Z(n17028) );
  AND U18886 ( .A(y[7850]), .B(x[488]), .Z(n18188) );
  AND U18887 ( .A(x[482]), .B(y[7844]), .Z(n17080) );
  NAND U18888 ( .A(n18188), .B(n17080), .Z(n16913) );
  NAND U18889 ( .A(n16911), .B(n16910), .Z(n16912) );
  NAND U18890 ( .A(n16913), .B(n16912), .Z(n16992) );
  NAND U18891 ( .A(y[7852]), .B(x[481]), .Z(n16914) );
  XNOR U18892 ( .A(n16915), .B(n16914), .Z(n16983) );
  AND U18893 ( .A(o[172]), .B(n16916), .Z(n16982) );
  XOR U18894 ( .A(n16983), .B(n16982), .Z(n16990) );
  AND U18895 ( .A(x[486]), .B(y[7847]), .Z(n17956) );
  AND U18896 ( .A(y[7851]), .B(x[482]), .Z(n16918) );
  NAND U18897 ( .A(y[7844]), .B(x[489]), .Z(n16917) );
  XNOR U18898 ( .A(n16918), .B(n16917), .Z(n17006) );
  XOR U18899 ( .A(n17956), .B(n17006), .Z(n16989) );
  XOR U18900 ( .A(n16990), .B(n16989), .Z(n16991) );
  XOR U18901 ( .A(n16992), .B(n16991), .Z(n17027) );
  NAND U18902 ( .A(n16920), .B(n16919), .Z(n16924) );
  ANDN U18903 ( .B(n16922), .A(n16921), .Z(n16923) );
  ANDN U18904 ( .B(n16924), .A(n16923), .Z(n17026) );
  XOR U18905 ( .A(n17027), .B(n17026), .Z(n17029) );
  XOR U18906 ( .A(n17028), .B(n17029), .Z(n17020) );
  NAND U18907 ( .A(n16926), .B(n16925), .Z(n16930) );
  NAND U18908 ( .A(n16928), .B(n16927), .Z(n16929) );
  NAND U18909 ( .A(n16930), .B(n16929), .Z(n16968) );
  AND U18910 ( .A(x[486]), .B(y[7851]), .Z(n17301) );
  IV U18911 ( .A(n17301), .Z(n17374) );
  AND U18912 ( .A(x[481]), .B(y[7846]), .Z(n16981) );
  NANDN U18913 ( .A(n17374), .B(n16981), .Z(n16934) );
  NAND U18914 ( .A(n16932), .B(n16931), .Z(n16933) );
  NAND U18915 ( .A(n16934), .B(n16933), .Z(n16974) );
  AND U18916 ( .A(x[492]), .B(y[7852]), .Z(n18194) );
  NAND U18917 ( .A(n18194), .B(n17140), .Z(n16938) );
  NAND U18918 ( .A(n16936), .B(n16935), .Z(n16937) );
  NAND U18919 ( .A(n16938), .B(n16937), .Z(n16972) );
  AND U18920 ( .A(x[490]), .B(y[7843]), .Z(n17830) );
  AND U18921 ( .A(y[7842]), .B(x[491]), .Z(n17793) );
  NAND U18922 ( .A(y[7845]), .B(x[488]), .Z(n16939) );
  XNOR U18923 ( .A(n17793), .B(n16939), .Z(n16978) );
  XOR U18924 ( .A(n17830), .B(n16978), .Z(n16971) );
  XOR U18925 ( .A(n16972), .B(n16971), .Z(n16973) );
  XOR U18926 ( .A(n16974), .B(n16973), .Z(n16966) );
  AND U18927 ( .A(x[484]), .B(y[7842]), .Z(n16941) );
  AND U18928 ( .A(x[490]), .B(y[7848]), .Z(n16940) );
  NAND U18929 ( .A(n16941), .B(n16940), .Z(n16944) );
  NAND U18930 ( .A(n16942), .B(n17553), .Z(n16943) );
  NAND U18931 ( .A(n16944), .B(n16943), .Z(n17017) );
  AND U18932 ( .A(y[7840]), .B(x[493]), .Z(n16946) );
  NAND U18933 ( .A(y[7853]), .B(x[480]), .Z(n16945) );
  XNOR U18934 ( .A(n16946), .B(n16945), .Z(n17000) );
  AND U18935 ( .A(x[492]), .B(y[7841]), .Z(n17011) );
  XOR U18936 ( .A(o[173]), .B(n17011), .Z(n16999) );
  XOR U18937 ( .A(n17000), .B(n16999), .Z(n17015) );
  AND U18938 ( .A(y[7848]), .B(x[485]), .Z(n16948) );
  NAND U18939 ( .A(y[7850]), .B(x[483]), .Z(n16947) );
  XNOR U18940 ( .A(n16948), .B(n16947), .Z(n16995) );
  AND U18941 ( .A(x[484]), .B(y[7849]), .Z(n16996) );
  XOR U18942 ( .A(n16995), .B(n16996), .Z(n17014) );
  XOR U18943 ( .A(n17015), .B(n17014), .Z(n17016) );
  XOR U18944 ( .A(n17017), .B(n17016), .Z(n16965) );
  XOR U18945 ( .A(n16966), .B(n16965), .Z(n16967) );
  XOR U18946 ( .A(n16968), .B(n16967), .Z(n17022) );
  XOR U18947 ( .A(n17023), .B(n17022), .Z(n17040) );
  NANDN U18948 ( .A(n16950), .B(n16949), .Z(n16954) );
  NAND U18949 ( .A(n16952), .B(n16951), .Z(n16953) );
  AND U18950 ( .A(n16954), .B(n16953), .Z(n17039) );
  XOR U18951 ( .A(n17041), .B(n17042), .Z(n17035) );
  NANDN U18952 ( .A(n16959), .B(n16958), .Z(n16963) );
  NANDN U18953 ( .A(n16961), .B(n16960), .Z(n16962) );
  AND U18954 ( .A(n16963), .B(n16962), .Z(n17033) );
  IV U18955 ( .A(n17033), .Z(n17032) );
  XOR U18956 ( .A(n17034), .B(n17032), .Z(n16964) );
  XNOR U18957 ( .A(n17035), .B(n16964), .Z(N366) );
  NAND U18958 ( .A(n16966), .B(n16965), .Z(n16970) );
  NAND U18959 ( .A(n16968), .B(n16967), .Z(n16969) );
  NAND U18960 ( .A(n16970), .B(n16969), .Z(n17049) );
  NAND U18961 ( .A(n16972), .B(n16971), .Z(n16976) );
  NAND U18962 ( .A(n16974), .B(n16973), .Z(n16975) );
  AND U18963 ( .A(n16976), .B(n16975), .Z(n17055) );
  AND U18964 ( .A(x[491]), .B(y[7845]), .Z(n17167) );
  NAND U18965 ( .A(n17167), .B(n16977), .Z(n16980) );
  NAND U18966 ( .A(n16978), .B(n17830), .Z(n16979) );
  NAND U18967 ( .A(n16980), .B(n16979), .Z(n17110) );
  AND U18968 ( .A(x[487]), .B(y[7852]), .Z(n17567) );
  NAND U18969 ( .A(n17567), .B(n16981), .Z(n16985) );
  NAND U18970 ( .A(n16983), .B(n16982), .Z(n16984) );
  NAND U18971 ( .A(n16985), .B(n16984), .Z(n17109) );
  XOR U18972 ( .A(n17110), .B(n17109), .Z(n17112) );
  AND U18973 ( .A(x[484]), .B(y[7850]), .Z(n17467) );
  AND U18974 ( .A(y[7851]), .B(x[483]), .Z(n16987) );
  NAND U18975 ( .A(y[7846]), .B(x[488]), .Z(n16986) );
  XNOR U18976 ( .A(n16987), .B(n16986), .Z(n17095) );
  XOR U18977 ( .A(n17372), .B(n17095), .Z(n17104) );
  XOR U18978 ( .A(n17467), .B(n17104), .Z(n17106) );
  AND U18979 ( .A(x[489]), .B(y[7845]), .Z(n17670) );
  AND U18980 ( .A(y[7852]), .B(x[482]), .Z(n16988) );
  AND U18981 ( .A(y[7844]), .B(x[490]), .Z(n17694) );
  XOR U18982 ( .A(n16988), .B(n17694), .Z(n17081) );
  XOR U18983 ( .A(n17670), .B(n17081), .Z(n17105) );
  XOR U18984 ( .A(n17106), .B(n17105), .Z(n17111) );
  XNOR U18985 ( .A(n17112), .B(n17111), .Z(n17053) );
  NAND U18986 ( .A(n16990), .B(n16989), .Z(n16994) );
  NAND U18987 ( .A(n16992), .B(n16991), .Z(n16993) );
  AND U18988 ( .A(n16994), .B(n16993), .Z(n17052) );
  XOR U18989 ( .A(n17053), .B(n17052), .Z(n17054) );
  XNOR U18990 ( .A(n17055), .B(n17054), .Z(n17047) );
  NAND U18991 ( .A(x[485]), .B(y[7850]), .Z(n17153) );
  NANDN U18992 ( .A(n17153), .B(n17820), .Z(n16998) );
  NAND U18993 ( .A(n16996), .B(n16995), .Z(n16997) );
  NAND U18994 ( .A(n16998), .B(n16997), .Z(n17061) );
  AND U18995 ( .A(x[493]), .B(y[7853]), .Z(n18527) );
  NAND U18996 ( .A(n18527), .B(n17140), .Z(n17002) );
  NAND U18997 ( .A(n17000), .B(n16999), .Z(n17001) );
  NAND U18998 ( .A(n17002), .B(n17001), .Z(n17059) );
  NAND U18999 ( .A(y[7843]), .B(x[491]), .Z(n17003) );
  XNOR U19000 ( .A(n17004), .B(n17003), .Z(n17085) );
  NAND U19001 ( .A(x[481]), .B(y[7853]), .Z(n17086) );
  XOR U19002 ( .A(n17059), .B(n17058), .Z(n17060) );
  XNOR U19003 ( .A(n17061), .B(n17060), .Z(n17116) );
  AND U19004 ( .A(x[489]), .B(y[7851]), .Z(n17005) );
  NAND U19005 ( .A(n17005), .B(n17080), .Z(n17008) );
  NAND U19006 ( .A(n17006), .B(n17956), .Z(n17007) );
  AND U19007 ( .A(n17008), .B(n17007), .Z(n17067) );
  AND U19008 ( .A(y[7840]), .B(x[494]), .Z(n17010) );
  NAND U19009 ( .A(y[7854]), .B(x[480]), .Z(n17009) );
  XNOR U19010 ( .A(n17010), .B(n17009), .Z(n17090) );
  AND U19011 ( .A(o[173]), .B(n17011), .Z(n17089) );
  XOR U19012 ( .A(n17090), .B(n17089), .Z(n17065) );
  NAND U19013 ( .A(y[7842]), .B(x[492]), .Z(n17012) );
  XNOR U19014 ( .A(n17013), .B(n17012), .Z(n17071) );
  NAND U19015 ( .A(x[493]), .B(y[7841]), .Z(n17079) );
  XNOR U19016 ( .A(o[174]), .B(n17079), .Z(n17072) );
  XOR U19017 ( .A(n17071), .B(n17072), .Z(n17064) );
  XOR U19018 ( .A(n17065), .B(n17064), .Z(n17066) );
  XOR U19019 ( .A(n17067), .B(n17066), .Z(n17115) );
  XOR U19020 ( .A(n17116), .B(n17115), .Z(n17118) );
  NAND U19021 ( .A(n17015), .B(n17014), .Z(n17019) );
  NAND U19022 ( .A(n17017), .B(n17016), .Z(n17018) );
  AND U19023 ( .A(n17019), .B(n17018), .Z(n17117) );
  XNOR U19024 ( .A(n17118), .B(n17117), .Z(n17046) );
  XOR U19025 ( .A(n17047), .B(n17046), .Z(n17048) );
  XOR U19026 ( .A(n17049), .B(n17048), .Z(n17131) );
  NANDN U19027 ( .A(n17021), .B(n17020), .Z(n17025) );
  NAND U19028 ( .A(n17023), .B(n17022), .Z(n17024) );
  AND U19029 ( .A(n17025), .B(n17024), .Z(n17129) );
  NAND U19030 ( .A(n17027), .B(n17026), .Z(n17031) );
  NAND U19031 ( .A(n17029), .B(n17028), .Z(n17030) );
  NAND U19032 ( .A(n17031), .B(n17030), .Z(n17128) );
  XNOR U19033 ( .A(n17131), .B(n17130), .Z(n17124) );
  OR U19034 ( .A(n17034), .B(n17032), .Z(n17038) );
  ANDN U19035 ( .B(n17034), .A(n17033), .Z(n17036) );
  OR U19036 ( .A(n17036), .B(n17035), .Z(n17037) );
  AND U19037 ( .A(n17038), .B(n17037), .Z(n17123) );
  NANDN U19038 ( .A(n17040), .B(n17039), .Z(n17044) );
  NAND U19039 ( .A(n17042), .B(n17041), .Z(n17043) );
  AND U19040 ( .A(n17044), .B(n17043), .Z(n17122) );
  IV U19041 ( .A(n17122), .Z(n17121) );
  XOR U19042 ( .A(n17123), .B(n17121), .Z(n17045) );
  XNOR U19043 ( .A(n17124), .B(n17045), .Z(N367) );
  NAND U19044 ( .A(n17047), .B(n17046), .Z(n17051) );
  NAND U19045 ( .A(n17049), .B(n17048), .Z(n17050) );
  AND U19046 ( .A(n17051), .B(n17050), .Z(n17228) );
  NAND U19047 ( .A(n17053), .B(n17052), .Z(n17057) );
  NAND U19048 ( .A(n17055), .B(n17054), .Z(n17056) );
  NAND U19049 ( .A(n17057), .B(n17056), .Z(n17197) );
  NAND U19050 ( .A(n17059), .B(n17058), .Z(n17063) );
  NAND U19051 ( .A(n17061), .B(n17060), .Z(n17062) );
  AND U19052 ( .A(n17063), .B(n17062), .Z(n17203) );
  NAND U19053 ( .A(n17065), .B(n17064), .Z(n17069) );
  NANDN U19054 ( .A(n17067), .B(n17066), .Z(n17068) );
  AND U19055 ( .A(n17069), .B(n17068), .Z(n17201) );
  AND U19056 ( .A(x[492]), .B(y[7847]), .Z(n17559) );
  NAND U19057 ( .A(n17559), .B(n17070), .Z(n17074) );
  NAND U19058 ( .A(n17072), .B(n17071), .Z(n17073) );
  AND U19059 ( .A(n17074), .B(n17073), .Z(n17177) );
  AND U19060 ( .A(y[7844]), .B(x[491]), .Z(n17076) );
  NAND U19061 ( .A(y[7842]), .B(x[493]), .Z(n17075) );
  XNOR U19062 ( .A(n17076), .B(n17075), .Z(n17181) );
  AND U19063 ( .A(x[492]), .B(y[7843]), .Z(n17180) );
  XNOR U19064 ( .A(n17181), .B(n17180), .Z(n17175) );
  AND U19065 ( .A(y[7840]), .B(x[495]), .Z(n17078) );
  NAND U19066 ( .A(y[7855]), .B(x[480]), .Z(n17077) );
  XNOR U19067 ( .A(n17078), .B(n17077), .Z(n17142) );
  ANDN U19068 ( .B(o[174]), .A(n17079), .Z(n17141) );
  XNOR U19069 ( .A(n17142), .B(n17141), .Z(n17174) );
  XOR U19070 ( .A(n17175), .B(n17174), .Z(n17176) );
  XOR U19071 ( .A(n17177), .B(n17176), .Z(n17209) );
  AND U19072 ( .A(x[490]), .B(y[7852]), .Z(n17957) );
  NAND U19073 ( .A(n17957), .B(n17080), .Z(n17083) );
  NAND U19074 ( .A(n17670), .B(n17081), .Z(n17082) );
  AND U19075 ( .A(n17083), .B(n17082), .Z(n17207) );
  AND U19076 ( .A(x[491]), .B(y[7848]), .Z(n17466) );
  NAND U19077 ( .A(n17466), .B(n17084), .Z(n17088) );
  NANDN U19078 ( .A(n17086), .B(n17085), .Z(n17087) );
  NAND U19079 ( .A(n17088), .B(n17087), .Z(n17206) );
  AND U19080 ( .A(x[494]), .B(y[7854]), .Z(n18809) );
  NAND U19081 ( .A(n18809), .B(n17140), .Z(n17092) );
  NAND U19082 ( .A(n17090), .B(n17089), .Z(n17091) );
  NAND U19083 ( .A(n17092), .B(n17091), .Z(n17169) );
  AND U19084 ( .A(x[488]), .B(y[7851]), .Z(n17093) );
  NAND U19085 ( .A(n17094), .B(n17093), .Z(n17097) );
  NAND U19086 ( .A(n17095), .B(n17372), .Z(n17096) );
  NAND U19087 ( .A(n17097), .B(n17096), .Z(n17168) );
  XOR U19088 ( .A(n17169), .B(n17168), .Z(n17171) );
  AND U19089 ( .A(y[7845]), .B(x[490]), .Z(n17099) );
  NAND U19090 ( .A(y[7851]), .B(x[484]), .Z(n17098) );
  XNOR U19091 ( .A(n17099), .B(n17098), .Z(n17148) );
  AND U19092 ( .A(x[487]), .B(y[7848]), .Z(n17147) );
  XNOR U19093 ( .A(n17148), .B(n17147), .Z(n17156) );
  AND U19094 ( .A(x[486]), .B(y[7849]), .Z(n17154) );
  IV U19095 ( .A(n17154), .Z(n17259) );
  XOR U19096 ( .A(n17259), .B(n17153), .Z(n17155) );
  XNOR U19097 ( .A(n17156), .B(n17155), .Z(n17191) );
  AND U19098 ( .A(y[7853]), .B(x[482]), .Z(n17101) );
  NAND U19099 ( .A(y[7846]), .B(x[489]), .Z(n17100) );
  XNOR U19100 ( .A(n17101), .B(n17100), .Z(n17159) );
  AND U19101 ( .A(x[483]), .B(y[7852]), .Z(n17160) );
  XOR U19102 ( .A(n17159), .B(n17160), .Z(n17189) );
  AND U19103 ( .A(y[7854]), .B(x[481]), .Z(n17103) );
  NAND U19104 ( .A(y[7847]), .B(x[488]), .Z(n17102) );
  XNOR U19105 ( .A(n17103), .B(n17102), .Z(n17137) );
  NAND U19106 ( .A(x[494]), .B(y[7841]), .Z(n17165) );
  XNOR U19107 ( .A(o[175]), .B(n17165), .Z(n17136) );
  XOR U19108 ( .A(n17137), .B(n17136), .Z(n17188) );
  XOR U19109 ( .A(n17189), .B(n17188), .Z(n17190) );
  XOR U19110 ( .A(n17191), .B(n17190), .Z(n17170) );
  XOR U19111 ( .A(n17171), .B(n17170), .Z(n17213) );
  NAND U19112 ( .A(n17467), .B(n17104), .Z(n17108) );
  NAND U19113 ( .A(n17106), .B(n17105), .Z(n17107) );
  AND U19114 ( .A(n17108), .B(n17107), .Z(n17212) );
  NAND U19115 ( .A(n17110), .B(n17109), .Z(n17114) );
  NAND U19116 ( .A(n17112), .B(n17111), .Z(n17113) );
  NAND U19117 ( .A(n17114), .B(n17113), .Z(n17215) );
  XOR U19118 ( .A(n17194), .B(n17195), .Z(n17196) );
  XNOR U19119 ( .A(n17197), .B(n17196), .Z(n17225) );
  NAND U19120 ( .A(n17116), .B(n17115), .Z(n17120) );
  NAND U19121 ( .A(n17118), .B(n17117), .Z(n17119) );
  AND U19122 ( .A(n17120), .B(n17119), .Z(n17226) );
  XOR U19123 ( .A(n17225), .B(n17226), .Z(n17227) );
  XOR U19124 ( .A(n17228), .B(n17227), .Z(n17221) );
  OR U19125 ( .A(n17123), .B(n17121), .Z(n17127) );
  ANDN U19126 ( .B(n17123), .A(n17122), .Z(n17125) );
  OR U19127 ( .A(n17125), .B(n17124), .Z(n17126) );
  AND U19128 ( .A(n17127), .B(n17126), .Z(n17220) );
  NANDN U19129 ( .A(n17129), .B(n17128), .Z(n17133) );
  NAND U19130 ( .A(n17131), .B(n17130), .Z(n17132) );
  NAND U19131 ( .A(n17133), .B(n17132), .Z(n17219) );
  IV U19132 ( .A(n17219), .Z(n17218) );
  XOR U19133 ( .A(n17220), .B(n17218), .Z(n17134) );
  XNOR U19134 ( .A(n17221), .B(n17134), .Z(N368) );
  AND U19135 ( .A(x[488]), .B(y[7854]), .Z(n17468) );
  NAND U19136 ( .A(n17468), .B(n17135), .Z(n17139) );
  NAND U19137 ( .A(n17137), .B(n17136), .Z(n17138) );
  NAND U19138 ( .A(n17139), .B(n17138), .Z(n17284) );
  AND U19139 ( .A(x[495]), .B(y[7855]), .Z(n19160) );
  NAND U19140 ( .A(n19160), .B(n17140), .Z(n17144) );
  NAND U19141 ( .A(n17142), .B(n17141), .Z(n17143) );
  NAND U19142 ( .A(n17144), .B(n17143), .Z(n17285) );
  XOR U19143 ( .A(n17284), .B(n17285), .Z(n17287) );
  AND U19144 ( .A(x[490]), .B(y[7851]), .Z(n17146) );
  NAND U19145 ( .A(n17146), .B(n17145), .Z(n17150) );
  NAND U19146 ( .A(n17148), .B(n17147), .Z(n17149) );
  NAND U19147 ( .A(n17150), .B(n17149), .Z(n17246) );
  AND U19148 ( .A(x[480]), .B(y[7856]), .Z(n17267) );
  AND U19149 ( .A(x[496]), .B(y[7840]), .Z(n17266) );
  XOR U19150 ( .A(n17267), .B(n17266), .Z(n17269) );
  AND U19151 ( .A(x[495]), .B(y[7841]), .Z(n17254) );
  XOR U19152 ( .A(n17254), .B(o[176]), .Z(n17268) );
  XOR U19153 ( .A(n17269), .B(n17268), .Z(n17245) );
  NAND U19154 ( .A(y[7849]), .B(x[487]), .Z(n17151) );
  XNOR U19155 ( .A(n17152), .B(n17151), .Z(n17261) );
  AND U19156 ( .A(x[490]), .B(y[7846]), .Z(n17260) );
  XOR U19157 ( .A(n17261), .B(n17260), .Z(n17244) );
  XOR U19158 ( .A(n17245), .B(n17244), .Z(n17247) );
  XOR U19159 ( .A(n17246), .B(n17247), .Z(n17286) );
  XNOR U19160 ( .A(n17287), .B(n17286), .Z(n17241) );
  NANDN U19161 ( .A(n17154), .B(n17153), .Z(n17158) );
  NAND U19162 ( .A(n17156), .B(n17155), .Z(n17157) );
  NAND U19163 ( .A(n17158), .B(n17157), .Z(n17239) );
  NAND U19164 ( .A(x[489]), .B(y[7853]), .Z(n17939) );
  NANDN U19165 ( .A(n17939), .B(n17558), .Z(n17162) );
  NAND U19166 ( .A(n17160), .B(n17159), .Z(n17161) );
  NAND U19167 ( .A(n17162), .B(n17161), .Z(n17274) );
  AND U19168 ( .A(y[7855]), .B(x[481]), .Z(n17164) );
  NAND U19169 ( .A(y[7848]), .B(x[488]), .Z(n17163) );
  XNOR U19170 ( .A(n17164), .B(n17163), .Z(n17265) );
  ANDN U19171 ( .B(o[175]), .A(n17165), .Z(n17264) );
  XOR U19172 ( .A(n17265), .B(n17264), .Z(n17273) );
  NAND U19173 ( .A(y[7842]), .B(x[494]), .Z(n17166) );
  XNOR U19174 ( .A(n17167), .B(n17166), .Z(n17292) );
  NAND U19175 ( .A(x[484]), .B(y[7852]), .Z(n17293) );
  XNOR U19176 ( .A(n17292), .B(n17293), .Z(n17272) );
  XOR U19177 ( .A(n17273), .B(n17272), .Z(n17275) );
  XNOR U19178 ( .A(n17274), .B(n17275), .Z(n17238) );
  XOR U19179 ( .A(n17239), .B(n17238), .Z(n17240) );
  XOR U19180 ( .A(n17241), .B(n17240), .Z(n17278) );
  NAND U19181 ( .A(n17169), .B(n17168), .Z(n17173) );
  NAND U19182 ( .A(n17171), .B(n17170), .Z(n17172) );
  AND U19183 ( .A(n17173), .B(n17172), .Z(n17279) );
  XOR U19184 ( .A(n17278), .B(n17279), .Z(n17281) );
  NAND U19185 ( .A(n17175), .B(n17174), .Z(n17179) );
  NAND U19186 ( .A(n17177), .B(n17176), .Z(n17178) );
  NAND U19187 ( .A(n17179), .B(n17178), .Z(n17306) );
  AND U19188 ( .A(x[493]), .B(y[7844]), .Z(n17303) );
  NAND U19189 ( .A(n17793), .B(n17303), .Z(n17183) );
  NAND U19190 ( .A(n17181), .B(n17180), .Z(n17182) );
  NAND U19191 ( .A(n17183), .B(n17182), .Z(n17290) );
  AND U19192 ( .A(y[7854]), .B(x[482]), .Z(n17185) );
  NAND U19193 ( .A(y[7847]), .B(x[489]), .Z(n17184) );
  XNOR U19194 ( .A(n17185), .B(n17184), .Z(n17296) );
  NAND U19195 ( .A(x[483]), .B(y[7853]), .Z(n17297) );
  XNOR U19196 ( .A(n17296), .B(n17297), .Z(n17289) );
  AND U19197 ( .A(x[492]), .B(y[7844]), .Z(n17927) );
  AND U19198 ( .A(y[7851]), .B(x[485]), .Z(n17187) );
  NAND U19199 ( .A(y[7843]), .B(x[493]), .Z(n17186) );
  XNOR U19200 ( .A(n17187), .B(n17186), .Z(n17251) );
  XOR U19201 ( .A(n17927), .B(n17251), .Z(n17288) );
  XOR U19202 ( .A(n17289), .B(n17288), .Z(n17291) );
  XNOR U19203 ( .A(n17290), .B(n17291), .Z(n17305) );
  NAND U19204 ( .A(n17189), .B(n17188), .Z(n17193) );
  NAND U19205 ( .A(n17191), .B(n17190), .Z(n17192) );
  AND U19206 ( .A(n17193), .B(n17192), .Z(n17304) );
  XOR U19207 ( .A(n17305), .B(n17304), .Z(n17307) );
  XOR U19208 ( .A(n17306), .B(n17307), .Z(n17280) );
  XNOR U19209 ( .A(n17281), .B(n17280), .Z(n17311) );
  NAND U19210 ( .A(n17195), .B(n17194), .Z(n17199) );
  NAND U19211 ( .A(n17197), .B(n17196), .Z(n17198) );
  AND U19212 ( .A(n17199), .B(n17198), .Z(n17310) );
  XOR U19213 ( .A(n17311), .B(n17310), .Z(n17313) );
  NANDN U19214 ( .A(n17201), .B(n17200), .Z(n17205) );
  NANDN U19215 ( .A(n17203), .B(n17202), .Z(n17204) );
  AND U19216 ( .A(n17205), .B(n17204), .Z(n17235) );
  NANDN U19217 ( .A(n17207), .B(n17206), .Z(n17211) );
  NANDN U19218 ( .A(n17209), .B(n17208), .Z(n17210) );
  AND U19219 ( .A(n17211), .B(n17210), .Z(n17233) );
  NANDN U19220 ( .A(n17213), .B(n17212), .Z(n17217) );
  NANDN U19221 ( .A(n17215), .B(n17214), .Z(n17216) );
  AND U19222 ( .A(n17217), .B(n17216), .Z(n17232) );
  XOR U19223 ( .A(n17313), .B(n17312), .Z(n17319) );
  OR U19224 ( .A(n17220), .B(n17218), .Z(n17224) );
  ANDN U19225 ( .B(n17220), .A(n17219), .Z(n17222) );
  OR U19226 ( .A(n17222), .B(n17221), .Z(n17223) );
  AND U19227 ( .A(n17224), .B(n17223), .Z(n17317) );
  NAND U19228 ( .A(n17226), .B(n17225), .Z(n17230) );
  NANDN U19229 ( .A(n17228), .B(n17227), .Z(n17229) );
  AND U19230 ( .A(n17230), .B(n17229), .Z(n17318) );
  IV U19231 ( .A(n17318), .Z(n17316) );
  XOR U19232 ( .A(n17317), .B(n17316), .Z(n17231) );
  XNOR U19233 ( .A(n17319), .B(n17231), .Z(N369) );
  NANDN U19234 ( .A(n17233), .B(n17232), .Z(n17237) );
  NANDN U19235 ( .A(n17235), .B(n17234), .Z(n17236) );
  AND U19236 ( .A(n17237), .B(n17236), .Z(n17410) );
  NAND U19237 ( .A(n17239), .B(n17238), .Z(n17243) );
  NAND U19238 ( .A(n17241), .B(n17240), .Z(n17242) );
  NAND U19239 ( .A(n17243), .B(n17242), .Z(n17332) );
  NAND U19240 ( .A(n17245), .B(n17244), .Z(n17249) );
  NAND U19241 ( .A(n17247), .B(n17246), .Z(n17248) );
  NAND U19242 ( .A(n17249), .B(n17248), .Z(n17402) );
  AND U19243 ( .A(x[493]), .B(y[7851]), .Z(n18202) );
  NAND U19244 ( .A(n18202), .B(n17250), .Z(n17253) );
  NAND U19245 ( .A(n17927), .B(n17251), .Z(n17252) );
  NAND U19246 ( .A(n17253), .B(n17252), .Z(n17362) );
  AND U19247 ( .A(n17254), .B(o[176]), .Z(n17377) );
  AND U19248 ( .A(y[7856]), .B(x[481]), .Z(n17256) );
  NAND U19249 ( .A(y[7848]), .B(x[489]), .Z(n17255) );
  XOR U19250 ( .A(n17256), .B(n17255), .Z(n17378) );
  AND U19251 ( .A(y[7842]), .B(x[495]), .Z(n17258) );
  NAND U19252 ( .A(y[7845]), .B(x[492]), .Z(n17257) );
  XNOR U19253 ( .A(n17258), .B(n17257), .Z(n17337) );
  AND U19254 ( .A(x[494]), .B(y[7843]), .Z(n17336) );
  XOR U19255 ( .A(n17337), .B(n17336), .Z(n17360) );
  XOR U19256 ( .A(n17361), .B(n17360), .Z(n17363) );
  XOR U19257 ( .A(n17362), .B(n17363), .Z(n17401) );
  AND U19258 ( .A(x[487]), .B(y[7850]), .Z(n17387) );
  NANDN U19259 ( .A(n17259), .B(n17387), .Z(n17263) );
  NAND U19260 ( .A(n17261), .B(n17260), .Z(n17262) );
  NAND U19261 ( .A(n17263), .B(n17262), .Z(n17368) );
  NAND U19262 ( .A(x[488]), .B(y[7855]), .Z(n18015) );
  AND U19263 ( .A(x[481]), .B(y[7848]), .Z(n17446) );
  XOR U19264 ( .A(n17368), .B(n17369), .Z(n17371) );
  AND U19265 ( .A(x[480]), .B(y[7857]), .Z(n17351) );
  AND U19266 ( .A(x[497]), .B(y[7840]), .Z(n17350) );
  XOR U19267 ( .A(n17351), .B(n17350), .Z(n17353) );
  AND U19268 ( .A(x[496]), .B(y[7841]), .Z(n17345) );
  XOR U19269 ( .A(n17345), .B(o[177]), .Z(n17352) );
  XOR U19270 ( .A(n17353), .B(n17352), .Z(n17365) );
  AND U19271 ( .A(y[7855]), .B(x[482]), .Z(n17271) );
  NAND U19272 ( .A(y[7847]), .B(x[490]), .Z(n17270) );
  XNOR U19273 ( .A(n17271), .B(n17270), .Z(n17383) );
  AND U19274 ( .A(x[483]), .B(y[7854]), .Z(n17382) );
  XOR U19275 ( .A(n17383), .B(n17382), .Z(n17364) );
  XOR U19276 ( .A(n17365), .B(n17364), .Z(n17367) );
  XOR U19277 ( .A(n17366), .B(n17367), .Z(n17370) );
  XOR U19278 ( .A(n17371), .B(n17370), .Z(n17400) );
  XOR U19279 ( .A(n17401), .B(n17400), .Z(n17403) );
  XNOR U19280 ( .A(n17402), .B(n17403), .Z(n17331) );
  NAND U19281 ( .A(n17273), .B(n17272), .Z(n17277) );
  NAND U19282 ( .A(n17275), .B(n17274), .Z(n17276) );
  AND U19283 ( .A(n17277), .B(n17276), .Z(n17330) );
  XNOR U19284 ( .A(n17331), .B(n17330), .Z(n17333) );
  XOR U19285 ( .A(n17332), .B(n17333), .Z(n17408) );
  NAND U19286 ( .A(n17279), .B(n17278), .Z(n17283) );
  NAND U19287 ( .A(n17281), .B(n17280), .Z(n17282) );
  NAND U19288 ( .A(n17283), .B(n17282), .Z(n17326) );
  AND U19289 ( .A(x[494]), .B(y[7845]), .Z(n17443) );
  IV U19290 ( .A(n17443), .Z(n17593) );
  NANDN U19291 ( .A(n17593), .B(n17793), .Z(n17295) );
  NANDN U19292 ( .A(n17293), .B(n17292), .Z(n17294) );
  AND U19293 ( .A(n17295), .B(n17294), .Z(n17391) );
  AND U19294 ( .A(x[489]), .B(y[7854]), .Z(n18183) );
  NANDN U19295 ( .A(n17381), .B(n18183), .Z(n17299) );
  NANDN U19296 ( .A(n17297), .B(n17296), .Z(n17298) );
  NAND U19297 ( .A(n17299), .B(n17298), .Z(n17390) );
  XNOR U19298 ( .A(n17391), .B(n17390), .Z(n17392) );
  AND U19299 ( .A(x[485]), .B(y[7852]), .Z(n17428) );
  NAND U19300 ( .A(y[7849]), .B(x[488]), .Z(n17300) );
  XNOR U19301 ( .A(n17428), .B(n17300), .Z(n17373) );
  XOR U19302 ( .A(n17373), .B(n17301), .Z(n17386) );
  XOR U19303 ( .A(n17387), .B(n17386), .Z(n17388) );
  NAND U19304 ( .A(y[7853]), .B(x[484]), .Z(n17302) );
  XNOR U19305 ( .A(n17303), .B(n17302), .Z(n17341) );
  NAND U19306 ( .A(x[491]), .B(y[7846]), .Z(n17342) );
  XOR U19307 ( .A(n17341), .B(n17342), .Z(n17389) );
  XOR U19308 ( .A(n17388), .B(n17389), .Z(n17393) );
  XNOR U19309 ( .A(n17392), .B(n17393), .Z(n17397) );
  XOR U19310 ( .A(n17396), .B(n17397), .Z(n17399) );
  XNOR U19311 ( .A(n17398), .B(n17399), .Z(n17325) );
  NAND U19312 ( .A(n17305), .B(n17304), .Z(n17309) );
  NAND U19313 ( .A(n17307), .B(n17306), .Z(n17308) );
  NAND U19314 ( .A(n17309), .B(n17308), .Z(n17324) );
  XNOR U19315 ( .A(n17325), .B(n17324), .Z(n17327) );
  XOR U19316 ( .A(n17326), .B(n17327), .Z(n17407) );
  XOR U19317 ( .A(n17408), .B(n17407), .Z(n17409) );
  XOR U19318 ( .A(n17410), .B(n17409), .Z(n17406) );
  NAND U19319 ( .A(n17311), .B(n17310), .Z(n17315) );
  NAND U19320 ( .A(n17313), .B(n17312), .Z(n17314) );
  NAND U19321 ( .A(n17315), .B(n17314), .Z(n17405) );
  NANDN U19322 ( .A(n17316), .B(n17317), .Z(n17322) );
  NOR U19323 ( .A(n17318), .B(n17317), .Z(n17320) );
  OR U19324 ( .A(n17320), .B(n17319), .Z(n17321) );
  AND U19325 ( .A(n17322), .B(n17321), .Z(n17404) );
  XOR U19326 ( .A(n17405), .B(n17404), .Z(n17323) );
  XNOR U19327 ( .A(n17406), .B(n17323), .Z(N370) );
  NAND U19328 ( .A(n17325), .B(n17324), .Z(n17329) );
  NANDN U19329 ( .A(n17327), .B(n17326), .Z(n17328) );
  AND U19330 ( .A(n17329), .B(n17328), .Z(n17522) );
  NAND U19331 ( .A(n17331), .B(n17330), .Z(n17335) );
  NANDN U19332 ( .A(n17333), .B(n17332), .Z(n17334) );
  AND U19333 ( .A(n17335), .B(n17334), .Z(n17520) );
  AND U19334 ( .A(x[492]), .B(y[7842]), .Z(n17665) );
  AND U19335 ( .A(x[495]), .B(y[7845]), .Z(n17566) );
  NAND U19336 ( .A(n17665), .B(n17566), .Z(n17339) );
  NAND U19337 ( .A(n17337), .B(n17336), .Z(n17338) );
  NAND U19338 ( .A(n17339), .B(n17338), .Z(n17494) );
  NAND U19339 ( .A(n18527), .B(n17340), .Z(n17344) );
  NANDN U19340 ( .A(n17342), .B(n17341), .Z(n17343) );
  AND U19341 ( .A(n17344), .B(n17343), .Z(n17485) );
  AND U19342 ( .A(n17345), .B(o[177]), .Z(n17447) );
  AND U19343 ( .A(y[7857]), .B(x[481]), .Z(n17347) );
  NAND U19344 ( .A(y[7848]), .B(x[490]), .Z(n17346) );
  XOR U19345 ( .A(n17347), .B(n17346), .Z(n17448) );
  AND U19346 ( .A(y[7843]), .B(x[495]), .Z(n17349) );
  NAND U19347 ( .A(y[7849]), .B(x[489]), .Z(n17348) );
  XNOR U19348 ( .A(n17349), .B(n17348), .Z(n17437) );
  NAND U19349 ( .A(x[494]), .B(y[7844]), .Z(n17438) );
  XOR U19350 ( .A(n17483), .B(n17482), .Z(n17484) );
  XOR U19351 ( .A(n17494), .B(n17495), .Z(n17497) );
  NAND U19352 ( .A(n17351), .B(n17350), .Z(n17355) );
  NAND U19353 ( .A(n17353), .B(n17352), .Z(n17354) );
  NAND U19354 ( .A(n17355), .B(n17354), .Z(n17506) );
  AND U19355 ( .A(y[7842]), .B(x[496]), .Z(n17357) );
  NAND U19356 ( .A(y[7847]), .B(x[491]), .Z(n17356) );
  XNOR U19357 ( .A(n17357), .B(n17356), .Z(n17433) );
  NAND U19358 ( .A(x[482]), .B(y[7856]), .Z(n17434) );
  XOR U19359 ( .A(n17506), .B(n17507), .Z(n17509) );
  AND U19360 ( .A(x[485]), .B(y[7853]), .Z(n17574) );
  NAND U19361 ( .A(y[7852]), .B(x[486]), .Z(n17358) );
  XNOR U19362 ( .A(n17574), .B(n17358), .Z(n17430) );
  NAND U19363 ( .A(y[7854]), .B(x[484]), .Z(n17359) );
  XNOR U19364 ( .A(n18188), .B(n17359), .Z(n17470) );
  AND U19365 ( .A(x[487]), .B(y[7851]), .Z(n17469) );
  XOR U19366 ( .A(n17470), .B(n17469), .Z(n17429) );
  XOR U19367 ( .A(n17430), .B(n17429), .Z(n17508) );
  XOR U19368 ( .A(n17509), .B(n17508), .Z(n17496) );
  XOR U19369 ( .A(n17497), .B(n17496), .Z(n17419) );
  XOR U19370 ( .A(n17489), .B(n17488), .Z(n17491) );
  XOR U19371 ( .A(n17491), .B(n17490), .Z(n17418) );
  XNOR U19372 ( .A(n17419), .B(n17418), .Z(n17421) );
  AND U19373 ( .A(x[488]), .B(y[7852]), .Z(n17588) );
  IV U19374 ( .A(n17588), .Z(n17699) );
  NANDN U19375 ( .A(n17699), .B(n17372), .Z(n17376) );
  NANDN U19376 ( .A(n17374), .B(n17373), .Z(n17375) );
  NAND U19377 ( .A(n17376), .B(n17375), .Z(n17501) );
  NAND U19378 ( .A(x[489]), .B(y[7856]), .Z(n18295) );
  NANDN U19379 ( .A(n18295), .B(n17446), .Z(n17380) );
  NANDN U19380 ( .A(n17378), .B(n17377), .Z(n17379) );
  NAND U19381 ( .A(n17380), .B(n17379), .Z(n17500) );
  XOR U19382 ( .A(n17501), .B(n17500), .Z(n17503) );
  NAND U19383 ( .A(x[490]), .B(y[7855]), .Z(n18294) );
  AND U19384 ( .A(x[480]), .B(y[7858]), .Z(n17451) );
  NAND U19385 ( .A(x[498]), .B(y[7840]), .Z(n17452) );
  NAND U19386 ( .A(x[497]), .B(y[7841]), .Z(n17473) );
  XOR U19387 ( .A(n17454), .B(n17453), .Z(n17477) );
  AND U19388 ( .A(y[7845]), .B(x[493]), .Z(n17385) );
  NAND U19389 ( .A(y[7855]), .B(x[483]), .Z(n17384) );
  XNOR U19390 ( .A(n17385), .B(n17384), .Z(n17459) );
  NAND U19391 ( .A(x[492]), .B(y[7846]), .Z(n17460) );
  XOR U19392 ( .A(n17477), .B(n17476), .Z(n17478) );
  XOR U19393 ( .A(n17503), .B(n17502), .Z(n17423) );
  NANDN U19394 ( .A(n17391), .B(n17390), .Z(n17395) );
  NANDN U19395 ( .A(n17393), .B(n17392), .Z(n17394) );
  AND U19396 ( .A(n17395), .B(n17394), .Z(n17424) );
  XOR U19397 ( .A(n17425), .B(n17424), .Z(n17420) );
  XOR U19398 ( .A(n17421), .B(n17420), .Z(n17416) );
  XNOR U19399 ( .A(n17414), .B(n17415), .Z(n17417) );
  XOR U19400 ( .A(n17416), .B(n17417), .Z(n17519) );
  XOR U19401 ( .A(n17520), .B(n17519), .Z(n17521) );
  XNOR U19402 ( .A(n17522), .B(n17521), .Z(n17515) );
  NAND U19403 ( .A(n17408), .B(n17407), .Z(n17412) );
  NANDN U19404 ( .A(n17410), .B(n17409), .Z(n17411) );
  NAND U19405 ( .A(n17412), .B(n17411), .Z(n17513) );
  IV U19406 ( .A(n17513), .Z(n17512) );
  XOR U19407 ( .A(n17514), .B(n17512), .Z(n17413) );
  XNOR U19408 ( .A(n17515), .B(n17413), .Z(N371) );
  NANDN U19409 ( .A(n17423), .B(n17422), .Z(n17427) );
  NAND U19410 ( .A(n17425), .B(n17424), .Z(n17426) );
  AND U19411 ( .A(n17427), .B(n17426), .Z(n17538) );
  AND U19412 ( .A(y[7853]), .B(x[486]), .Z(n17474) );
  NAND U19413 ( .A(n17474), .B(n17428), .Z(n17432) );
  NAND U19414 ( .A(n17430), .B(n17429), .Z(n17431) );
  AND U19415 ( .A(n17432), .B(n17431), .Z(n17628) );
  AND U19416 ( .A(x[496]), .B(y[7847]), .Z(n17943) );
  NAND U19417 ( .A(n17943), .B(n17793), .Z(n17436) );
  NANDN U19418 ( .A(n17434), .B(n17433), .Z(n17435) );
  AND U19419 ( .A(n17436), .B(n17435), .Z(n17626) );
  AND U19420 ( .A(x[495]), .B(y[7849]), .Z(n18215) );
  NAND U19421 ( .A(n18215), .B(n17553), .Z(n17440) );
  NANDN U19422 ( .A(n17438), .B(n17437), .Z(n17439) );
  NAND U19423 ( .A(n17440), .B(n17439), .Z(n17543) );
  AND U19424 ( .A(y[7858]), .B(x[481]), .Z(n17442) );
  NAND U19425 ( .A(y[7851]), .B(x[488]), .Z(n17441) );
  XNOR U19426 ( .A(n17442), .B(n17441), .Z(n17592) );
  XOR U19427 ( .A(n17592), .B(n17443), .Z(n17542) );
  AND U19428 ( .A(y[7846]), .B(x[493]), .Z(n17445) );
  NAND U19429 ( .A(y[7857]), .B(x[482]), .Z(n17444) );
  XNOR U19430 ( .A(n17445), .B(n17444), .Z(n17560) );
  XOR U19431 ( .A(n17560), .B(n17559), .Z(n17541) );
  XOR U19432 ( .A(n17542), .B(n17541), .Z(n17544) );
  XOR U19433 ( .A(n17543), .B(n17544), .Z(n17625) );
  AND U19434 ( .A(x[490]), .B(y[7857]), .Z(n18623) );
  IV U19435 ( .A(n18623), .Z(n18488) );
  NANDN U19436 ( .A(n18488), .B(n17446), .Z(n17450) );
  NANDN U19437 ( .A(n17448), .B(n17447), .Z(n17449) );
  NAND U19438 ( .A(n17450), .B(n17449), .Z(n17603) );
  NANDN U19439 ( .A(n17452), .B(n17451), .Z(n17456) );
  NAND U19440 ( .A(n17454), .B(n17453), .Z(n17455) );
  NAND U19441 ( .A(n17456), .B(n17455), .Z(n17601) );
  AND U19442 ( .A(y[7843]), .B(x[496]), .Z(n18154) );
  NAND U19443 ( .A(y[7850]), .B(x[489]), .Z(n17457) );
  XNOR U19444 ( .A(n18154), .B(n17457), .Z(n17555) );
  AND U19445 ( .A(x[495]), .B(y[7844]), .Z(n17554) );
  XOR U19446 ( .A(n17555), .B(n17554), .Z(n17602) );
  XNOR U19447 ( .A(n17601), .B(n17602), .Z(n17604) );
  AND U19448 ( .A(x[493]), .B(y[7855]), .Z(n18838) );
  NANDN U19449 ( .A(n17458), .B(n18838), .Z(n17462) );
  NANDN U19450 ( .A(n17460), .B(n17459), .Z(n17461) );
  NAND U19451 ( .A(n17462), .B(n17461), .Z(n17609) );
  AND U19452 ( .A(y[7849]), .B(x[490]), .Z(n17464) );
  NAND U19453 ( .A(y[7842]), .B(x[497]), .Z(n17463) );
  XNOR U19454 ( .A(n17464), .B(n17463), .Z(n17598) );
  AND U19455 ( .A(x[498]), .B(y[7841]), .Z(n17573) );
  XOR U19456 ( .A(n17573), .B(o[179]), .Z(n17597) );
  XOR U19457 ( .A(n17598), .B(n17597), .Z(n17608) );
  NAND U19458 ( .A(y[7856]), .B(x[483]), .Z(n17465) );
  XNOR U19459 ( .A(n17466), .B(n17465), .Z(n17568) );
  XOR U19460 ( .A(n17568), .B(n17567), .Z(n17607) );
  XOR U19461 ( .A(n17608), .B(n17607), .Z(n17610) );
  XNOR U19462 ( .A(n17609), .B(n17610), .Z(n17620) );
  NAND U19463 ( .A(n17468), .B(n17467), .Z(n17472) );
  NAND U19464 ( .A(n17470), .B(n17469), .Z(n17471) );
  NAND U19465 ( .A(n17472), .B(n17471), .Z(n17549) );
  AND U19466 ( .A(x[480]), .B(y[7859]), .Z(n17579) );
  AND U19467 ( .A(x[499]), .B(y[7840]), .Z(n17578) );
  XOR U19468 ( .A(n17579), .B(n17578), .Z(n17581) );
  ANDN U19469 ( .B(o[178]), .A(n17473), .Z(n17580) );
  XOR U19470 ( .A(n17581), .B(n17580), .Z(n17548) );
  AND U19471 ( .A(x[484]), .B(y[7855]), .Z(n17712) );
  AND U19472 ( .A(x[485]), .B(y[7854]), .Z(n17475) );
  XOR U19473 ( .A(n17475), .B(n17474), .Z(n17575) );
  XOR U19474 ( .A(n17712), .B(n17575), .Z(n17547) );
  XOR U19475 ( .A(n17548), .B(n17547), .Z(n17550) );
  XNOR U19476 ( .A(n17549), .B(n17550), .Z(n17619) );
  XOR U19477 ( .A(n17620), .B(n17619), .Z(n17622) );
  XNOR U19478 ( .A(n17621), .B(n17622), .Z(n17615) );
  NAND U19479 ( .A(n17477), .B(n17476), .Z(n17481) );
  NANDN U19480 ( .A(n17479), .B(n17478), .Z(n17480) );
  AND U19481 ( .A(n17481), .B(n17480), .Z(n17614) );
  NAND U19482 ( .A(n17483), .B(n17482), .Z(n17487) );
  NANDN U19483 ( .A(n17485), .B(n17484), .Z(n17486) );
  NAND U19484 ( .A(n17487), .B(n17486), .Z(n17613) );
  XNOR U19485 ( .A(n17615), .B(n17616), .Z(n17535) );
  XOR U19486 ( .A(n17536), .B(n17535), .Z(n17537) );
  NAND U19487 ( .A(n17489), .B(n17488), .Z(n17493) );
  NAND U19488 ( .A(n17491), .B(n17490), .Z(n17492) );
  AND U19489 ( .A(n17493), .B(n17492), .Z(n17631) );
  NAND U19490 ( .A(n17495), .B(n17494), .Z(n17499) );
  NAND U19491 ( .A(n17497), .B(n17496), .Z(n17498) );
  NAND U19492 ( .A(n17499), .B(n17498), .Z(n17639) );
  NAND U19493 ( .A(n17501), .B(n17500), .Z(n17505) );
  NAND U19494 ( .A(n17503), .B(n17502), .Z(n17504) );
  NAND U19495 ( .A(n17505), .B(n17504), .Z(n17638) );
  NAND U19496 ( .A(n17507), .B(n17506), .Z(n17511) );
  NAND U19497 ( .A(n17509), .B(n17508), .Z(n17510) );
  NAND U19498 ( .A(n17511), .B(n17510), .Z(n17637) );
  XNOR U19499 ( .A(n17638), .B(n17637), .Z(n17640) );
  XNOR U19500 ( .A(n17631), .B(n17632), .Z(n17633) );
  XNOR U19501 ( .A(n17527), .B(n17526), .Z(n17529) );
  XOR U19502 ( .A(n17528), .B(n17529), .Z(n17534) );
  OR U19503 ( .A(n17514), .B(n17512), .Z(n17518) );
  ANDN U19504 ( .B(n17514), .A(n17513), .Z(n17516) );
  OR U19505 ( .A(n17516), .B(n17515), .Z(n17517) );
  AND U19506 ( .A(n17518), .B(n17517), .Z(n17533) );
  NAND U19507 ( .A(n17520), .B(n17519), .Z(n17524) );
  NAND U19508 ( .A(n17522), .B(n17521), .Z(n17523) );
  NAND U19509 ( .A(n17524), .B(n17523), .Z(n17532) );
  XNOR U19510 ( .A(n17533), .B(n17532), .Z(n17525) );
  XNOR U19511 ( .A(n17534), .B(n17525), .Z(N372) );
  NAND U19512 ( .A(n17527), .B(n17526), .Z(n17531) );
  NANDN U19513 ( .A(n17529), .B(n17528), .Z(n17530) );
  AND U19514 ( .A(n17531), .B(n17530), .Z(n17651) );
  NAND U19515 ( .A(n17536), .B(n17535), .Z(n17540) );
  NANDN U19516 ( .A(n17538), .B(n17537), .Z(n17539) );
  AND U19517 ( .A(n17540), .B(n17539), .Z(n17748) );
  NAND U19518 ( .A(n17542), .B(n17541), .Z(n17546) );
  NAND U19519 ( .A(n17544), .B(n17543), .Z(n17545) );
  NAND U19520 ( .A(n17546), .B(n17545), .Z(n17654) );
  NAND U19521 ( .A(n17548), .B(n17547), .Z(n17552) );
  NAND U19522 ( .A(n17550), .B(n17549), .Z(n17551) );
  NAND U19523 ( .A(n17552), .B(n17551), .Z(n17653) );
  XOR U19524 ( .A(n17654), .B(n17653), .Z(n17656) );
  AND U19525 ( .A(x[496]), .B(y[7850]), .Z(n18446) );
  NAND U19526 ( .A(n18446), .B(n17553), .Z(n17557) );
  NAND U19527 ( .A(n17555), .B(n17554), .Z(n17556) );
  NAND U19528 ( .A(n17557), .B(n17556), .Z(n17688) );
  AND U19529 ( .A(y[7857]), .B(x[493]), .Z(n19075) );
  NAND U19530 ( .A(n19075), .B(n17558), .Z(n17562) );
  NAND U19531 ( .A(n17560), .B(n17559), .Z(n17561) );
  NAND U19532 ( .A(n17562), .B(n17561), .Z(n17729) );
  AND U19533 ( .A(y[7844]), .B(x[496]), .Z(n17564) );
  NAND U19534 ( .A(y[7850]), .B(x[490]), .Z(n17563) );
  XNOR U19535 ( .A(n17564), .B(n17563), .Z(n17696) );
  AND U19536 ( .A(x[482]), .B(y[7858]), .Z(n17695) );
  XOR U19537 ( .A(n17696), .B(n17695), .Z(n17728) );
  NAND U19538 ( .A(y[7851]), .B(x[489]), .Z(n17565) );
  XNOR U19539 ( .A(n17566), .B(n17565), .Z(n17672) );
  AND U19540 ( .A(x[494]), .B(y[7846]), .Z(n17671) );
  XOR U19541 ( .A(n17672), .B(n17671), .Z(n17727) );
  XOR U19542 ( .A(n17728), .B(n17727), .Z(n17730) );
  XOR U19543 ( .A(n17729), .B(n17730), .Z(n17689) );
  XOR U19544 ( .A(n17688), .B(n17689), .Z(n17691) );
  NAND U19545 ( .A(x[491]), .B(y[7856]), .Z(n18624) );
  NANDN U19546 ( .A(n18624), .B(n17820), .Z(n17570) );
  NAND U19547 ( .A(n17568), .B(n17567), .Z(n17569) );
  NAND U19548 ( .A(n17570), .B(n17569), .Z(n17735) );
  AND U19549 ( .A(y[7849]), .B(x[491]), .Z(n17572) );
  NAND U19550 ( .A(y[7859]), .B(x[481]), .Z(n17571) );
  XNOR U19551 ( .A(n17572), .B(n17571), .Z(n17669) );
  AND U19552 ( .A(x[499]), .B(y[7841]), .Z(n17675) );
  XOR U19553 ( .A(n17675), .B(o[180]), .Z(n17668) );
  XOR U19554 ( .A(n17669), .B(n17668), .Z(n17734) );
  AND U19555 ( .A(x[480]), .B(y[7860]), .Z(n17718) );
  AND U19556 ( .A(x[500]), .B(y[7840]), .Z(n17717) );
  XOR U19557 ( .A(n17718), .B(n17717), .Z(n17720) );
  AND U19558 ( .A(n17573), .B(o[179]), .Z(n17719) );
  XOR U19559 ( .A(n17720), .B(n17719), .Z(n17733) );
  XOR U19560 ( .A(n17734), .B(n17733), .Z(n17736) );
  XOR U19561 ( .A(n17735), .B(n17736), .Z(n17690) );
  XOR U19562 ( .A(n17691), .B(n17690), .Z(n17655) );
  XOR U19563 ( .A(n17656), .B(n17655), .Z(n17742) );
  NAND U19564 ( .A(x[486]), .B(y[7854]), .Z(n17660) );
  NANDN U19565 ( .A(n17660), .B(n17574), .Z(n17577) );
  NAND U19566 ( .A(n17712), .B(n17575), .Z(n17576) );
  NAND U19567 ( .A(n17577), .B(n17576), .Z(n17678) );
  NAND U19568 ( .A(n17579), .B(n17578), .Z(n17583) );
  NAND U19569 ( .A(n17581), .B(n17580), .Z(n17582) );
  NAND U19570 ( .A(n17583), .B(n17582), .Z(n17676) );
  AND U19571 ( .A(y[7842]), .B(x[498]), .Z(n17585) );
  NAND U19572 ( .A(y[7848]), .B(x[492]), .Z(n17584) );
  XNOR U19573 ( .A(n17585), .B(n17584), .Z(n17667) );
  AND U19574 ( .A(x[497]), .B(y[7843]), .Z(n17666) );
  XOR U19575 ( .A(n17667), .B(n17666), .Z(n17677) );
  XOR U19576 ( .A(n17676), .B(n17677), .Z(n17679) );
  XOR U19577 ( .A(n17678), .B(n17679), .Z(n17683) );
  AND U19578 ( .A(y[7847]), .B(x[493]), .Z(n17587) );
  NAND U19579 ( .A(y[7857]), .B(x[483]), .Z(n17586) );
  XNOR U19580 ( .A(n17587), .B(n17586), .Z(n17698) );
  XNOR U19581 ( .A(n17698), .B(n17588), .Z(n17662) );
  AND U19582 ( .A(y[7855]), .B(x[485]), .Z(n17590) );
  NAND U19583 ( .A(y[7856]), .B(x[484]), .Z(n17589) );
  XNOR U19584 ( .A(n17590), .B(n17589), .Z(n17714) );
  AND U19585 ( .A(x[487]), .B(y[7853]), .Z(n17713) );
  XNOR U19586 ( .A(n17714), .B(n17713), .Z(n17659) );
  XOR U19587 ( .A(n17660), .B(n17659), .Z(n17661) );
  XNOR U19588 ( .A(n17662), .B(n17661), .Z(n17723) );
  AND U19589 ( .A(x[488]), .B(y[7858]), .Z(n18789) );
  AND U19590 ( .A(x[481]), .B(y[7851]), .Z(n17591) );
  NAND U19591 ( .A(n18789), .B(n17591), .Z(n17595) );
  NANDN U19592 ( .A(n17593), .B(n17592), .Z(n17594) );
  NAND U19593 ( .A(n17595), .B(n17594), .Z(n17722) );
  NAND U19594 ( .A(x[497]), .B(y[7849]), .Z(n18455) );
  NANDN U19595 ( .A(n18455), .B(n17596), .Z(n17600) );
  NAND U19596 ( .A(n17598), .B(n17597), .Z(n17599) );
  NAND U19597 ( .A(n17600), .B(n17599), .Z(n17721) );
  XNOR U19598 ( .A(n17722), .B(n17721), .Z(n17724) );
  XOR U19599 ( .A(n17723), .B(n17724), .Z(n17682) );
  NAND U19600 ( .A(n17602), .B(n17601), .Z(n17606) );
  NANDN U19601 ( .A(n17604), .B(n17603), .Z(n17605) );
  AND U19602 ( .A(n17606), .B(n17605), .Z(n17684) );
  XOR U19603 ( .A(n17685), .B(n17684), .Z(n17740) );
  NAND U19604 ( .A(n17608), .B(n17607), .Z(n17612) );
  NAND U19605 ( .A(n17610), .B(n17609), .Z(n17611) );
  AND U19606 ( .A(n17612), .B(n17611), .Z(n17739) );
  XOR U19607 ( .A(n17740), .B(n17739), .Z(n17741) );
  NANDN U19608 ( .A(n17614), .B(n17613), .Z(n17618) );
  NAND U19609 ( .A(n17616), .B(n17615), .Z(n17617) );
  AND U19610 ( .A(n17618), .B(n17617), .Z(n17754) );
  NAND U19611 ( .A(n17620), .B(n17619), .Z(n17624) );
  NAND U19612 ( .A(n17622), .B(n17621), .Z(n17623) );
  AND U19613 ( .A(n17624), .B(n17623), .Z(n17752) );
  NANDN U19614 ( .A(n17626), .B(n17625), .Z(n17630) );
  NANDN U19615 ( .A(n17628), .B(n17627), .Z(n17629) );
  AND U19616 ( .A(n17630), .B(n17629), .Z(n17751) );
  XNOR U19617 ( .A(n17754), .B(n17753), .Z(n17745) );
  XOR U19618 ( .A(n17746), .B(n17745), .Z(n17747) );
  XOR U19619 ( .A(n17748), .B(n17747), .Z(n17646) );
  NANDN U19620 ( .A(n17632), .B(n17631), .Z(n17636) );
  NANDN U19621 ( .A(n17634), .B(n17633), .Z(n17635) );
  NAND U19622 ( .A(n17636), .B(n17635), .Z(n17645) );
  NAND U19623 ( .A(n17638), .B(n17637), .Z(n17642) );
  NANDN U19624 ( .A(n17640), .B(n17639), .Z(n17641) );
  NAND U19625 ( .A(n17642), .B(n17641), .Z(n17644) );
  XNOR U19626 ( .A(n17645), .B(n17644), .Z(n17647) );
  XOR U19627 ( .A(n17650), .B(n17652), .Z(n17643) );
  XOR U19628 ( .A(n17651), .B(n17643), .Z(N373) );
  NAND U19629 ( .A(n17645), .B(n17644), .Z(n17649) );
  NANDN U19630 ( .A(n17647), .B(n17646), .Z(n17648) );
  AND U19631 ( .A(n17649), .B(n17648), .Z(n17764) );
  NAND U19632 ( .A(n17654), .B(n17653), .Z(n17658) );
  NAND U19633 ( .A(n17656), .B(n17655), .Z(n17657) );
  NAND U19634 ( .A(n17658), .B(n17657), .Z(n17775) );
  NAND U19635 ( .A(n17660), .B(n17659), .Z(n17664) );
  NAND U19636 ( .A(n17662), .B(n17661), .Z(n17663) );
  NAND U19637 ( .A(n17664), .B(n17663), .Z(n17855) );
  AND U19638 ( .A(x[498]), .B(y[7848]), .Z(n18453) );
  NAND U19639 ( .A(x[491]), .B(y[7859]), .Z(n19135) );
  XOR U19640 ( .A(n17838), .B(n17839), .Z(n17841) );
  AND U19641 ( .A(x[495]), .B(y[7851]), .Z(n18441) );
  NAND U19642 ( .A(n18441), .B(n17670), .Z(n17674) );
  NAND U19643 ( .A(n17672), .B(n17671), .Z(n17673) );
  NAND U19644 ( .A(n17674), .B(n17673), .Z(n17806) );
  AND U19645 ( .A(n17675), .B(o[180]), .Z(n17829) );
  AND U19646 ( .A(x[480]), .B(y[7861]), .Z(n17827) );
  AND U19647 ( .A(x[501]), .B(y[7840]), .Z(n17826) );
  XOR U19648 ( .A(n17827), .B(n17826), .Z(n17828) );
  XOR U19649 ( .A(n17829), .B(n17828), .Z(n17805) );
  AND U19650 ( .A(x[485]), .B(y[7856]), .Z(n17811) );
  AND U19651 ( .A(x[496]), .B(y[7845]), .Z(n17810) );
  XOR U19652 ( .A(n17811), .B(n17810), .Z(n17813) );
  AND U19653 ( .A(x[495]), .B(y[7846]), .Z(n17812) );
  XOR U19654 ( .A(n17813), .B(n17812), .Z(n17804) );
  XOR U19655 ( .A(n17805), .B(n17804), .Z(n17807) );
  XOR U19656 ( .A(n17806), .B(n17807), .Z(n17840) );
  XNOR U19657 ( .A(n17841), .B(n17840), .Z(n17854) );
  XOR U19658 ( .A(n17855), .B(n17854), .Z(n17857) );
  NAND U19659 ( .A(n17677), .B(n17676), .Z(n17681) );
  NAND U19660 ( .A(n17679), .B(n17678), .Z(n17680) );
  AND U19661 ( .A(n17681), .B(n17680), .Z(n17856) );
  XOR U19662 ( .A(n17857), .B(n17856), .Z(n17774) );
  NANDN U19663 ( .A(n17683), .B(n17682), .Z(n17687) );
  NAND U19664 ( .A(n17685), .B(n17684), .Z(n17686) );
  AND U19665 ( .A(n17687), .B(n17686), .Z(n17773) );
  XNOR U19666 ( .A(n17775), .B(n17776), .Z(n17769) );
  NAND U19667 ( .A(n17689), .B(n17688), .Z(n17693) );
  NAND U19668 ( .A(n17691), .B(n17690), .Z(n17692) );
  NAND U19669 ( .A(n17693), .B(n17692), .Z(n17862) );
  NAND U19670 ( .A(n19075), .B(n17697), .Z(n17701) );
  NANDN U19671 ( .A(n17699), .B(n17698), .Z(n17700) );
  NAND U19672 ( .A(n17701), .B(n17700), .Z(n17849) );
  AND U19673 ( .A(y[7842]), .B(x[499]), .Z(n17703) );
  NAND U19674 ( .A(y[7850]), .B(x[491]), .Z(n17702) );
  XNOR U19675 ( .A(n17703), .B(n17702), .Z(n17795) );
  AND U19676 ( .A(x[500]), .B(y[7841]), .Z(n17825) );
  XOR U19677 ( .A(n17825), .B(o[181]), .Z(n17794) );
  XOR U19678 ( .A(n17795), .B(n17794), .Z(n17847) );
  AND U19679 ( .A(y[7843]), .B(x[498]), .Z(n17705) );
  NAND U19680 ( .A(y[7851]), .B(x[490]), .Z(n17704) );
  XNOR U19681 ( .A(n17705), .B(n17704), .Z(n17832) );
  AND U19682 ( .A(x[481]), .B(y[7860]), .Z(n17831) );
  XOR U19683 ( .A(n17832), .B(n17831), .Z(n17846) );
  XOR U19684 ( .A(n17847), .B(n17846), .Z(n17850) );
  XOR U19685 ( .A(n17849), .B(n17850), .Z(n17780) );
  XOR U19686 ( .A(n17779), .B(n17780), .Z(n17782) );
  AND U19687 ( .A(x[487]), .B(y[7854]), .Z(n18013) );
  AND U19688 ( .A(y[7855]), .B(x[486]), .Z(n17707) );
  AND U19689 ( .A(y[7847]), .B(x[494]), .Z(n17706) );
  XOR U19690 ( .A(n17707), .B(n17706), .Z(n17835) );
  XNOR U19691 ( .A(n18013), .B(n17835), .Z(n17786) );
  NAND U19692 ( .A(x[489]), .B(y[7852]), .Z(n17784) );
  NAND U19693 ( .A(x[488]), .B(y[7853]), .Z(n17783) );
  XOR U19694 ( .A(n17784), .B(n17783), .Z(n17785) );
  XNOR U19695 ( .A(n17786), .B(n17785), .Z(n17801) );
  AND U19696 ( .A(y[7849]), .B(x[492]), .Z(n17709) );
  NAND U19697 ( .A(y[7844]), .B(x[497]), .Z(n17708) );
  XNOR U19698 ( .A(n17709), .B(n17708), .Z(n17790) );
  AND U19699 ( .A(x[482]), .B(y[7859]), .Z(n17789) );
  XOR U19700 ( .A(n17790), .B(n17789), .Z(n17799) );
  AND U19701 ( .A(y[7848]), .B(x[493]), .Z(n17711) );
  NAND U19702 ( .A(y[7858]), .B(x[483]), .Z(n17710) );
  XNOR U19703 ( .A(n17711), .B(n17710), .Z(n17822) );
  AND U19704 ( .A(x[484]), .B(y[7857]), .Z(n17821) );
  XOR U19705 ( .A(n17822), .B(n17821), .Z(n17798) );
  XOR U19706 ( .A(n17799), .B(n17798), .Z(n17800) );
  XOR U19707 ( .A(n17801), .B(n17800), .Z(n17845) );
  NAND U19708 ( .A(n17811), .B(n17712), .Z(n17716) );
  NAND U19709 ( .A(n17714), .B(n17713), .Z(n17715) );
  NAND U19710 ( .A(n17716), .B(n17715), .Z(n17842) );
  XOR U19711 ( .A(n17842), .B(n17843), .Z(n17844) );
  XOR U19712 ( .A(n17845), .B(n17844), .Z(n17781) );
  XOR U19713 ( .A(n17782), .B(n17781), .Z(n17860) );
  NAND U19714 ( .A(n17722), .B(n17721), .Z(n17726) );
  NANDN U19715 ( .A(n17724), .B(n17723), .Z(n17725) );
  NAND U19716 ( .A(n17726), .B(n17725), .Z(n17868) );
  NAND U19717 ( .A(n17728), .B(n17727), .Z(n17732) );
  NAND U19718 ( .A(n17730), .B(n17729), .Z(n17731) );
  NAND U19719 ( .A(n17732), .B(n17731), .Z(n17867) );
  NAND U19720 ( .A(n17734), .B(n17733), .Z(n17738) );
  NAND U19721 ( .A(n17736), .B(n17735), .Z(n17737) );
  NAND U19722 ( .A(n17738), .B(n17737), .Z(n17866) );
  XNOR U19723 ( .A(n17867), .B(n17866), .Z(n17869) );
  XNOR U19724 ( .A(n17860), .B(n17861), .Z(n17863) );
  XOR U19725 ( .A(n17862), .B(n17863), .Z(n17768) );
  NAND U19726 ( .A(n17740), .B(n17739), .Z(n17744) );
  NANDN U19727 ( .A(n17742), .B(n17741), .Z(n17743) );
  NAND U19728 ( .A(n17744), .B(n17743), .Z(n17767) );
  XOR U19729 ( .A(n17769), .B(n17770), .Z(n17760) );
  NAND U19730 ( .A(n17746), .B(n17745), .Z(n17750) );
  NAND U19731 ( .A(n17748), .B(n17747), .Z(n17749) );
  AND U19732 ( .A(n17750), .B(n17749), .Z(n17759) );
  NANDN U19733 ( .A(n17752), .B(n17751), .Z(n17756) );
  NAND U19734 ( .A(n17754), .B(n17753), .Z(n17755) );
  AND U19735 ( .A(n17756), .B(n17755), .Z(n17758) );
  XOR U19736 ( .A(n17760), .B(n17761), .Z(n17766) );
  XNOR U19737 ( .A(n17765), .B(n17766), .Z(n17757) );
  XOR U19738 ( .A(n17764), .B(n17757), .Z(N374) );
  NANDN U19739 ( .A(n17759), .B(n17758), .Z(n17763) );
  NAND U19740 ( .A(n17761), .B(n17760), .Z(n17762) );
  NAND U19741 ( .A(n17763), .B(n17762), .Z(n17983) );
  IV U19742 ( .A(n17983), .Z(n17979) );
  NANDN U19743 ( .A(n17768), .B(n17767), .Z(n17772) );
  NANDN U19744 ( .A(n17770), .B(n17769), .Z(n17771) );
  AND U19745 ( .A(n17772), .B(n17771), .Z(n17988) );
  NANDN U19746 ( .A(n17774), .B(n17773), .Z(n17778) );
  NAND U19747 ( .A(n17776), .B(n17775), .Z(n17777) );
  NAND U19748 ( .A(n17778), .B(n17777), .Z(n17986) );
  NAND U19749 ( .A(n17784), .B(n17783), .Z(n17788) );
  NAND U19750 ( .A(n17786), .B(n17785), .Z(n17787) );
  NAND U19751 ( .A(n17788), .B(n17787), .Z(n17973) );
  AND U19752 ( .A(x[485]), .B(y[7857]), .Z(n17950) );
  AND U19753 ( .A(x[497]), .B(y[7845]), .Z(n17949) );
  XOR U19754 ( .A(n17950), .B(n17949), .Z(n17952) );
  AND U19755 ( .A(x[496]), .B(y[7846]), .Z(n17951) );
  XOR U19756 ( .A(n17952), .B(n17951), .Z(n17903) );
  AND U19757 ( .A(y[7844]), .B(x[498]), .Z(n17792) );
  NAND U19758 ( .A(y[7850]), .B(x[492]), .Z(n17791) );
  XNOR U19759 ( .A(n17792), .B(n17791), .Z(n17929) );
  AND U19760 ( .A(x[484]), .B(y[7858]), .Z(n17928) );
  XNOR U19761 ( .A(n17929), .B(n17928), .Z(n17904) );
  XNOR U19762 ( .A(n17903), .B(n17904), .Z(n17905) );
  XNOR U19763 ( .A(n17906), .B(n17905), .Z(n17972) );
  NAND U19764 ( .A(x[499]), .B(y[7850]), .Z(n18973) );
  NANDN U19765 ( .A(n18973), .B(n17793), .Z(n17797) );
  NAND U19766 ( .A(n17795), .B(n17794), .Z(n17796) );
  AND U19767 ( .A(n17797), .B(n17796), .Z(n17971) );
  XNOR U19768 ( .A(n17972), .B(n17971), .Z(n17974) );
  XOR U19769 ( .A(n17973), .B(n17974), .Z(n17976) );
  NAND U19770 ( .A(n17799), .B(n17798), .Z(n17803) );
  NAND U19771 ( .A(n17801), .B(n17800), .Z(n17802) );
  NAND U19772 ( .A(n17803), .B(n17802), .Z(n17961) );
  NAND U19773 ( .A(n17805), .B(n17804), .Z(n17809) );
  NAND U19774 ( .A(n17807), .B(n17806), .Z(n17808) );
  NAND U19775 ( .A(n17809), .B(n17808), .Z(n17962) );
  XOR U19776 ( .A(n17961), .B(n17962), .Z(n17964) );
  AND U19777 ( .A(n17811), .B(n17810), .Z(n17815) );
  NAND U19778 ( .A(n17813), .B(n17812), .Z(n17814) );
  NANDN U19779 ( .A(n17815), .B(n17814), .Z(n17925) );
  AND U19780 ( .A(y[7849]), .B(x[493]), .Z(n17817) );
  NAND U19781 ( .A(y[7842]), .B(x[500]), .Z(n17816) );
  XNOR U19782 ( .A(n17817), .B(n17816), .Z(n17946) );
  AND U19783 ( .A(x[482]), .B(y[7860]), .Z(n17945) );
  XOR U19784 ( .A(n17946), .B(n17945), .Z(n17924) );
  AND U19785 ( .A(y[7856]), .B(x[486]), .Z(n17819) );
  NAND U19786 ( .A(y[7847]), .B(x[495]), .Z(n17818) );
  XNOR U19787 ( .A(n17819), .B(n17818), .Z(n17958) );
  XOR U19788 ( .A(n17958), .B(n17957), .Z(n17923) );
  XOR U19789 ( .A(n17924), .B(n17923), .Z(n17926) );
  XOR U19790 ( .A(n17925), .B(n17926), .Z(n17965) );
  AND U19791 ( .A(x[493]), .B(y[7858]), .Z(n19251) );
  NAND U19792 ( .A(n17820), .B(n19251), .Z(n17824) );
  NAND U19793 ( .A(n17822), .B(n17821), .Z(n17823) );
  NAND U19794 ( .A(n17824), .B(n17823), .Z(n17896) );
  AND U19795 ( .A(x[481]), .B(y[7861]), .Z(n17917) );
  XOR U19796 ( .A(n17918), .B(n17917), .Z(n17916) );
  AND U19797 ( .A(n17825), .B(o[181]), .Z(n17915) );
  XOR U19798 ( .A(n17916), .B(n17915), .Z(n17894) );
  AND U19799 ( .A(x[494]), .B(y[7848]), .Z(n17909) );
  AND U19800 ( .A(x[483]), .B(y[7859]), .Z(n17910) );
  XOR U19801 ( .A(n17909), .B(n17910), .Z(n17911) );
  AND U19802 ( .A(x[499]), .B(y[7843]), .Z(n17912) );
  XOR U19803 ( .A(n17911), .B(n17912), .Z(n17893) );
  XOR U19804 ( .A(n17894), .B(n17893), .Z(n17895) );
  XNOR U19805 ( .A(n17896), .B(n17895), .Z(n17966) );
  XNOR U19806 ( .A(n17965), .B(n17966), .Z(n17968) );
  AND U19807 ( .A(x[498]), .B(y[7851]), .Z(n18975) );
  NAND U19808 ( .A(n18975), .B(n17830), .Z(n17834) );
  NAND U19809 ( .A(n17832), .B(n17831), .Z(n17833) );
  NAND U19810 ( .A(n17834), .B(n17833), .Z(n17890) );
  XOR U19811 ( .A(n17889), .B(n17890), .Z(n17891) );
  AND U19812 ( .A(x[494]), .B(y[7855]), .Z(n18985) );
  AND U19813 ( .A(x[480]), .B(y[7862]), .Z(n17933) );
  AND U19814 ( .A(x[502]), .B(y[7840]), .Z(n17932) );
  XOR U19815 ( .A(n17933), .B(n17932), .Z(n17935) );
  AND U19816 ( .A(x[501]), .B(y[7841]), .Z(n17955) );
  XOR U19817 ( .A(n17955), .B(o[182]), .Z(n17934) );
  XOR U19818 ( .A(n17935), .B(n17934), .Z(n17898) );
  AND U19819 ( .A(y[7855]), .B(x[487]), .Z(n17837) );
  NAND U19820 ( .A(y[7854]), .B(x[488]), .Z(n17836) );
  XNOR U19821 ( .A(n17837), .B(n17836), .Z(n17938) );
  XOR U19822 ( .A(n17898), .B(n17897), .Z(n17900) );
  XNOR U19823 ( .A(n17899), .B(n17900), .Z(n17892) );
  XNOR U19824 ( .A(n17891), .B(n17892), .Z(n17967) );
  XOR U19825 ( .A(n17968), .B(n17967), .Z(n17963) );
  XOR U19826 ( .A(n17964), .B(n17963), .Z(n17975) );
  XNOR U19827 ( .A(n17976), .B(n17975), .Z(n17978) );
  XNOR U19828 ( .A(n17977), .B(n17978), .Z(n17882) );
  IV U19829 ( .A(n17846), .Z(n17848) );
  NANDN U19830 ( .A(n17848), .B(n17847), .Z(n17853) );
  IV U19831 ( .A(n17849), .Z(n17851) );
  NANDN U19832 ( .A(n17851), .B(n17850), .Z(n17852) );
  NAND U19833 ( .A(n17853), .B(n17852), .Z(n17886) );
  XOR U19834 ( .A(n17885), .B(n17886), .Z(n17888) );
  XOR U19835 ( .A(n17887), .B(n17888), .Z(n17880) );
  NAND U19836 ( .A(n17855), .B(n17854), .Z(n17859) );
  NAND U19837 ( .A(n17857), .B(n17856), .Z(n17858) );
  NAND U19838 ( .A(n17859), .B(n17858), .Z(n17879) );
  XNOR U19839 ( .A(n17882), .B(n17881), .Z(n17875) );
  NANDN U19840 ( .A(n17861), .B(n17860), .Z(n17865) );
  NAND U19841 ( .A(n17863), .B(n17862), .Z(n17864) );
  NAND U19842 ( .A(n17865), .B(n17864), .Z(n17874) );
  NAND U19843 ( .A(n17867), .B(n17866), .Z(n17871) );
  NANDN U19844 ( .A(n17869), .B(n17868), .Z(n17870) );
  NAND U19845 ( .A(n17871), .B(n17870), .Z(n17873) );
  XNOR U19846 ( .A(n17874), .B(n17873), .Z(n17876) );
  XOR U19847 ( .A(n17986), .B(n17987), .Z(n17989) );
  XNOR U19848 ( .A(n17988), .B(n17989), .Z(n17980) );
  XNOR U19849 ( .A(n17982), .B(n17980), .Z(n17872) );
  XOR U19850 ( .A(n17979), .B(n17872), .Z(N375) );
  NAND U19851 ( .A(n17874), .B(n17873), .Z(n17878) );
  NANDN U19852 ( .A(n17876), .B(n17875), .Z(n17877) );
  AND U19853 ( .A(n17878), .B(n17877), .Z(n18126) );
  NANDN U19854 ( .A(n17880), .B(n17879), .Z(n17884) );
  NAND U19855 ( .A(n17882), .B(n17881), .Z(n17883) );
  NAND U19856 ( .A(n17884), .B(n17883), .Z(n18123) );
  NAND U19857 ( .A(n17898), .B(n17897), .Z(n17902) );
  NAND U19858 ( .A(n17900), .B(n17899), .Z(n17901) );
  NAND U19859 ( .A(n17902), .B(n17901), .Z(n18100) );
  XOR U19860 ( .A(n18101), .B(n18100), .Z(n18103) );
  XOR U19861 ( .A(n18102), .B(n18103), .Z(n18116) );
  NANDN U19862 ( .A(n17904), .B(n17903), .Z(n17908) );
  NANDN U19863 ( .A(n17906), .B(n17905), .Z(n17907) );
  NAND U19864 ( .A(n17908), .B(n17907), .Z(n18114) );
  NAND U19865 ( .A(n17910), .B(n17909), .Z(n17914) );
  NAND U19866 ( .A(n17912), .B(n17911), .Z(n17913) );
  NAND U19867 ( .A(n17914), .B(n17913), .Z(n18047) );
  AND U19868 ( .A(n17916), .B(n17915), .Z(n17920) );
  NAND U19869 ( .A(n17918), .B(n17917), .Z(n17919) );
  NANDN U19870 ( .A(n17920), .B(n17919), .Z(n18046) );
  XOR U19871 ( .A(n18047), .B(n18046), .Z(n18049) );
  AND U19872 ( .A(y[7856]), .B(x[487]), .Z(n17922) );
  NAND U19873 ( .A(y[7854]), .B(x[489]), .Z(n17921) );
  XNOR U19874 ( .A(n17922), .B(n17921), .Z(n18014) );
  NAND U19875 ( .A(x[490]), .B(y[7853]), .Z(n18053) );
  AND U19876 ( .A(x[486]), .B(y[7857]), .Z(n18005) );
  AND U19877 ( .A(x[495]), .B(y[7848]), .Z(n18006) );
  XOR U19878 ( .A(n18005), .B(n18006), .Z(n18007) );
  AND U19879 ( .A(x[491]), .B(y[7852]), .Z(n18008) );
  XOR U19880 ( .A(n18007), .B(n18008), .Z(n18054) );
  XOR U19881 ( .A(n18055), .B(n18054), .Z(n18048) );
  XOR U19882 ( .A(n18049), .B(n18048), .Z(n18115) );
  XOR U19883 ( .A(n18114), .B(n18115), .Z(n18117) );
  XOR U19884 ( .A(n18116), .B(n18117), .Z(n18107) );
  AND U19885 ( .A(x[498]), .B(y[7850]), .Z(n18820) );
  NAND U19886 ( .A(n18820), .B(n17927), .Z(n17931) );
  NAND U19887 ( .A(n17929), .B(n17928), .Z(n17930) );
  NAND U19888 ( .A(n17931), .B(n17930), .Z(n18077) );
  NAND U19889 ( .A(n17933), .B(n17932), .Z(n17937) );
  NAND U19890 ( .A(n17935), .B(n17934), .Z(n17936) );
  NAND U19891 ( .A(n17937), .B(n17936), .Z(n18076) );
  XOR U19892 ( .A(n18077), .B(n18076), .Z(n18078) );
  NANDN U19893 ( .A(n18015), .B(n18013), .Z(n17941) );
  NANDN U19894 ( .A(n17939), .B(n17938), .Z(n17940) );
  NAND U19895 ( .A(n17941), .B(n17940), .Z(n18090) );
  AND U19896 ( .A(x[480]), .B(y[7863]), .Z(n18024) );
  NAND U19897 ( .A(x[503]), .B(y[7840]), .Z(n18025) );
  AND U19898 ( .A(x[502]), .B(y[7841]), .Z(n18004) );
  XOR U19899 ( .A(o[183]), .B(n18004), .Z(n18026) );
  XOR U19900 ( .A(n18027), .B(n18026), .Z(n18089) );
  NAND U19901 ( .A(y[7843]), .B(x[500]), .Z(n17942) );
  XNOR U19902 ( .A(n17943), .B(n17942), .Z(n18000) );
  AND U19903 ( .A(x[499]), .B(y[7844]), .Z(n18001) );
  XOR U19904 ( .A(n18000), .B(n18001), .Z(n18088) );
  XOR U19905 ( .A(n18089), .B(n18088), .Z(n18091) );
  XOR U19906 ( .A(n18090), .B(n18091), .Z(n18079) );
  XOR U19907 ( .A(n18078), .B(n18079), .Z(n18041) );
  XOR U19908 ( .A(n18040), .B(n18041), .Z(n18043) );
  NAND U19909 ( .A(x[500]), .B(y[7849]), .Z(n18997) );
  AND U19910 ( .A(x[493]), .B(y[7842]), .Z(n17944) );
  NANDN U19911 ( .A(n18997), .B(n17944), .Z(n17948) );
  NAND U19912 ( .A(n17946), .B(n17945), .Z(n17947) );
  NAND U19913 ( .A(n17948), .B(n17947), .Z(n18034) );
  NAND U19914 ( .A(n17950), .B(n17949), .Z(n17954) );
  NAND U19915 ( .A(n17952), .B(n17951), .Z(n17953) );
  NAND U19916 ( .A(n17954), .B(n17953), .Z(n18096) );
  AND U19917 ( .A(x[493]), .B(y[7850]), .Z(n18070) );
  NAND U19918 ( .A(x[482]), .B(y[7861]), .Z(n18071) );
  NAND U19919 ( .A(x[501]), .B(y[7842]), .Z(n18073) );
  AND U19920 ( .A(x[492]), .B(y[7851]), .Z(n18018) );
  NAND U19921 ( .A(x[481]), .B(y[7862]), .Z(n18019) );
  AND U19922 ( .A(n17955), .B(o[182]), .Z(n18020) );
  XOR U19923 ( .A(n18021), .B(n18020), .Z(n18094) );
  XOR U19924 ( .A(n18095), .B(n18094), .Z(n18097) );
  XOR U19925 ( .A(n18096), .B(n18097), .Z(n18035) );
  XOR U19926 ( .A(n18034), .B(n18035), .Z(n18036) );
  AND U19927 ( .A(x[495]), .B(y[7856]), .Z(n19239) );
  NAND U19928 ( .A(n17956), .B(n19239), .Z(n17960) );
  NAND U19929 ( .A(n17958), .B(n17957), .Z(n17959) );
  NAND U19930 ( .A(n17960), .B(n17959), .Z(n18084) );
  AND U19931 ( .A(x[494]), .B(y[7849]), .Z(n18064) );
  NAND U19932 ( .A(x[483]), .B(y[7860]), .Z(n18065) );
  NAND U19933 ( .A(x[484]), .B(y[7859]), .Z(n18067) );
  AND U19934 ( .A(x[485]), .B(y[7858]), .Z(n18058) );
  AND U19935 ( .A(x[498]), .B(y[7845]), .Z(n18059) );
  XOR U19936 ( .A(n18058), .B(n18059), .Z(n18060) );
  AND U19937 ( .A(x[497]), .B(y[7846]), .Z(n18061) );
  XOR U19938 ( .A(n18060), .B(n18061), .Z(n18082) );
  XOR U19939 ( .A(n18083), .B(n18082), .Z(n18085) );
  XOR U19940 ( .A(n18084), .B(n18085), .Z(n18037) );
  XOR U19941 ( .A(n18036), .B(n18037), .Z(n18042) );
  XOR U19942 ( .A(n18043), .B(n18042), .Z(n18106) );
  XOR U19943 ( .A(n18107), .B(n18106), .Z(n18109) );
  XOR U19944 ( .A(n18108), .B(n18109), .Z(n17996) );
  NANDN U19945 ( .A(n17966), .B(n17965), .Z(n17970) );
  NAND U19946 ( .A(n17968), .B(n17967), .Z(n17969) );
  NAND U19947 ( .A(n17970), .B(n17969), .Z(n18110) );
  XOR U19948 ( .A(n18110), .B(n18111), .Z(n18113) );
  XOR U19949 ( .A(n18112), .B(n18113), .Z(n17994) );
  XNOR U19950 ( .A(n17994), .B(n17993), .Z(n17995) );
  XNOR U19951 ( .A(n17996), .B(n17995), .Z(n18124) );
  XOR U19952 ( .A(n18123), .B(n18124), .Z(n18125) );
  XNOR U19953 ( .A(n18126), .B(n18125), .Z(n18122) );
  ANDN U19954 ( .B(n17982), .A(n17979), .Z(n17981) );
  OR U19955 ( .A(n17981), .B(n17980), .Z(n17985) );
  NOR U19956 ( .A(n17983), .B(n17982), .Z(n17984) );
  ANDN U19957 ( .B(n17985), .A(n17984), .Z(n18121) );
  NANDN U19958 ( .A(n17987), .B(n17986), .Z(n17991) );
  NANDN U19959 ( .A(n17989), .B(n17988), .Z(n17990) );
  AND U19960 ( .A(n17991), .B(n17990), .Z(n18120) );
  XOR U19961 ( .A(n18121), .B(n18120), .Z(n17992) );
  XNOR U19962 ( .A(n18122), .B(n17992), .Z(N376) );
  NANDN U19963 ( .A(n17994), .B(n17993), .Z(n17998) );
  NANDN U19964 ( .A(n17996), .B(n17995), .Z(n17997) );
  AND U19965 ( .A(n17998), .B(n17997), .Z(n18266) );
  AND U19966 ( .A(x[500]), .B(y[7847]), .Z(n17999) );
  NAND U19967 ( .A(n17999), .B(n18154), .Z(n18003) );
  NAND U19968 ( .A(n18001), .B(n18000), .Z(n18002) );
  NAND U19969 ( .A(n18003), .B(n18002), .Z(n18174) );
  AND U19970 ( .A(x[502]), .B(y[7842]), .Z(n18193) );
  XOR U19971 ( .A(n18194), .B(n18193), .Z(n18195) );
  AND U19972 ( .A(x[482]), .B(y[7862]), .Z(n18196) );
  XOR U19973 ( .A(n18195), .B(n18196), .Z(n18172) );
  AND U19974 ( .A(x[481]), .B(y[7863]), .Z(n18201) );
  XOR U19975 ( .A(n18202), .B(n18201), .Z(n18200) );
  AND U19976 ( .A(o[183]), .B(n18004), .Z(n18199) );
  XOR U19977 ( .A(n18200), .B(n18199), .Z(n18171) );
  XOR U19978 ( .A(n18172), .B(n18171), .Z(n18173) );
  XOR U19979 ( .A(n18174), .B(n18173), .Z(n18231) );
  NAND U19980 ( .A(n18006), .B(n18005), .Z(n18010) );
  NAND U19981 ( .A(n18008), .B(n18007), .Z(n18009) );
  NAND U19982 ( .A(n18010), .B(n18009), .Z(n18168) );
  AND U19983 ( .A(y[7848]), .B(x[496]), .Z(n18012) );
  NAND U19984 ( .A(y[7843]), .B(x[501]), .Z(n18011) );
  XNOR U19985 ( .A(n18012), .B(n18011), .Z(n18155) );
  AND U19986 ( .A(x[485]), .B(y[7859]), .Z(n18156) );
  XOR U19987 ( .A(n18155), .B(n18156), .Z(n18166) );
  AND U19988 ( .A(x[486]), .B(y[7858]), .Z(n18538) );
  AND U19989 ( .A(x[500]), .B(y[7844]), .Z(n18369) );
  XOR U19990 ( .A(n18538), .B(n18369), .Z(n18161) );
  AND U19991 ( .A(x[499]), .B(y[7845]), .Z(n18162) );
  XOR U19992 ( .A(n18161), .B(n18162), .Z(n18165) );
  XOR U19993 ( .A(n18166), .B(n18165), .Z(n18167) );
  XOR U19994 ( .A(n18168), .B(n18167), .Z(n18145) );
  NANDN U19995 ( .A(n18295), .B(n18013), .Z(n18017) );
  NANDN U19996 ( .A(n18015), .B(n18014), .Z(n18016) );
  NAND U19997 ( .A(n18017), .B(n18016), .Z(n18143) );
  NANDN U19998 ( .A(n18019), .B(n18018), .Z(n18023) );
  NAND U19999 ( .A(n18021), .B(n18020), .Z(n18022) );
  NAND U20000 ( .A(n18023), .B(n18022), .Z(n18142) );
  XOR U20001 ( .A(n18143), .B(n18142), .Z(n18144) );
  XOR U20002 ( .A(n18145), .B(n18144), .Z(n18230) );
  XOR U20003 ( .A(n18231), .B(n18230), .Z(n18233) );
  NANDN U20004 ( .A(n18025), .B(n18024), .Z(n18029) );
  NAND U20005 ( .A(n18027), .B(n18026), .Z(n18028) );
  NAND U20006 ( .A(n18029), .B(n18028), .Z(n18225) );
  AND U20007 ( .A(x[483]), .B(y[7861]), .Z(n18214) );
  XOR U20008 ( .A(n18215), .B(n18214), .Z(n18213) );
  AND U20009 ( .A(x[484]), .B(y[7860]), .Z(n18212) );
  XOR U20010 ( .A(n18213), .B(n18212), .Z(n18224) );
  XOR U20011 ( .A(n18225), .B(n18224), .Z(n18227) );
  AND U20012 ( .A(y[7855]), .B(x[489]), .Z(n18031) );
  NAND U20013 ( .A(y[7854]), .B(x[490]), .Z(n18030) );
  XNOR U20014 ( .A(n18031), .B(n18030), .Z(n18185) );
  AND U20015 ( .A(y[7850]), .B(x[494]), .Z(n18033) );
  NAND U20016 ( .A(y[7856]), .B(x[488]), .Z(n18032) );
  XNOR U20017 ( .A(n18033), .B(n18032), .Z(n18189) );
  NAND U20018 ( .A(x[491]), .B(y[7853]), .Z(n18190) );
  XOR U20019 ( .A(n18185), .B(n18184), .Z(n18226) );
  XOR U20020 ( .A(n18227), .B(n18226), .Z(n18232) );
  XNOR U20021 ( .A(n18233), .B(n18232), .Z(n18243) );
  NAND U20022 ( .A(n18035), .B(n18034), .Z(n18039) );
  NAND U20023 ( .A(n18037), .B(n18036), .Z(n18038) );
  AND U20024 ( .A(n18039), .B(n18038), .Z(n18242) );
  XOR U20025 ( .A(n18243), .B(n18242), .Z(n18245) );
  NAND U20026 ( .A(n18041), .B(n18040), .Z(n18045) );
  NAND U20027 ( .A(n18043), .B(n18042), .Z(n18044) );
  AND U20028 ( .A(n18045), .B(n18044), .Z(n18244) );
  XOR U20029 ( .A(n18245), .B(n18244), .Z(n18251) );
  NAND U20030 ( .A(n18047), .B(n18046), .Z(n18051) );
  NAND U20031 ( .A(n18049), .B(n18048), .Z(n18050) );
  AND U20032 ( .A(n18051), .B(n18050), .Z(n18239) );
  NANDN U20033 ( .A(n18053), .B(n18052), .Z(n18057) );
  NAND U20034 ( .A(n18055), .B(n18054), .Z(n18056) );
  AND U20035 ( .A(n18057), .B(n18056), .Z(n18237) );
  NAND U20036 ( .A(n18059), .B(n18058), .Z(n18063) );
  NAND U20037 ( .A(n18061), .B(n18060), .Z(n18062) );
  NAND U20038 ( .A(n18063), .B(n18062), .Z(n18151) );
  AND U20039 ( .A(x[480]), .B(y[7864]), .Z(n18219) );
  AND U20040 ( .A(x[504]), .B(y[7840]), .Z(n18218) );
  XOR U20041 ( .A(n18219), .B(n18218), .Z(n18221) );
  AND U20042 ( .A(x[503]), .B(y[7841]), .Z(n18211) );
  XOR U20043 ( .A(n18211), .B(o[184]), .Z(n18220) );
  XOR U20044 ( .A(n18221), .B(n18220), .Z(n18149) );
  AND U20045 ( .A(x[487]), .B(y[7857]), .Z(n18205) );
  AND U20046 ( .A(x[498]), .B(y[7846]), .Z(n18206) );
  XOR U20047 ( .A(n18205), .B(n18206), .Z(n18207) );
  AND U20048 ( .A(x[497]), .B(y[7847]), .Z(n18208) );
  XOR U20049 ( .A(n18207), .B(n18208), .Z(n18148) );
  XOR U20050 ( .A(n18149), .B(n18148), .Z(n18150) );
  XOR U20051 ( .A(n18151), .B(n18150), .Z(n18139) );
  NANDN U20052 ( .A(n18065), .B(n18064), .Z(n18069) );
  NANDN U20053 ( .A(n18067), .B(n18066), .Z(n18068) );
  AND U20054 ( .A(n18069), .B(n18068), .Z(n18137) );
  NANDN U20055 ( .A(n18071), .B(n18070), .Z(n18075) );
  NANDN U20056 ( .A(n18073), .B(n18072), .Z(n18074) );
  NAND U20057 ( .A(n18075), .B(n18074), .Z(n18136) );
  XOR U20058 ( .A(n18139), .B(n18138), .Z(n18236) );
  NAND U20059 ( .A(n18077), .B(n18076), .Z(n18081) );
  NAND U20060 ( .A(n18079), .B(n18078), .Z(n18080) );
  AND U20061 ( .A(n18081), .B(n18080), .Z(n18180) );
  NAND U20062 ( .A(n18083), .B(n18082), .Z(n18087) );
  NAND U20063 ( .A(n18085), .B(n18084), .Z(n18086) );
  AND U20064 ( .A(n18087), .B(n18086), .Z(n18178) );
  NAND U20065 ( .A(n18089), .B(n18088), .Z(n18093) );
  NAND U20066 ( .A(n18091), .B(n18090), .Z(n18092) );
  AND U20067 ( .A(n18093), .B(n18092), .Z(n18177) );
  XOR U20068 ( .A(n18178), .B(n18177), .Z(n18179) );
  XOR U20069 ( .A(n18180), .B(n18179), .Z(n18131) );
  NAND U20070 ( .A(n18095), .B(n18094), .Z(n18099) );
  NAND U20071 ( .A(n18097), .B(n18096), .Z(n18098) );
  AND U20072 ( .A(n18099), .B(n18098), .Z(n18130) );
  XOR U20073 ( .A(n18131), .B(n18130), .Z(n18132) );
  XOR U20074 ( .A(n18133), .B(n18132), .Z(n18249) );
  NAND U20075 ( .A(n18101), .B(n18100), .Z(n18105) );
  NAND U20076 ( .A(n18103), .B(n18102), .Z(n18104) );
  AND U20077 ( .A(n18105), .B(n18104), .Z(n18248) );
  XOR U20078 ( .A(n18249), .B(n18248), .Z(n18250) );
  XOR U20079 ( .A(n18251), .B(n18250), .Z(n18264) );
  NAND U20080 ( .A(n18115), .B(n18114), .Z(n18119) );
  NAND U20081 ( .A(n18117), .B(n18116), .Z(n18118) );
  NAND U20082 ( .A(n18119), .B(n18118), .Z(n18254) );
  XOR U20083 ( .A(n18255), .B(n18254), .Z(n18257) );
  XOR U20084 ( .A(n18256), .B(n18257), .Z(n18263) );
  XNOR U20085 ( .A(n18264), .B(n18263), .Z(n18265) );
  XNOR U20086 ( .A(n18266), .B(n18265), .Z(n18262) );
  NAND U20087 ( .A(n18124), .B(n18123), .Z(n18128) );
  NAND U20088 ( .A(n18126), .B(n18125), .Z(n18127) );
  AND U20089 ( .A(n18128), .B(n18127), .Z(n18260) );
  XOR U20090 ( .A(n18261), .B(n18260), .Z(n18129) );
  XNOR U20091 ( .A(n18262), .B(n18129), .Z(N377) );
  NAND U20092 ( .A(n18131), .B(n18130), .Z(n18135) );
  NAND U20093 ( .A(n18133), .B(n18132), .Z(n18134) );
  NAND U20094 ( .A(n18135), .B(n18134), .Z(n18278) );
  NANDN U20095 ( .A(n18137), .B(n18136), .Z(n18141) );
  NAND U20096 ( .A(n18139), .B(n18138), .Z(n18140) );
  AND U20097 ( .A(n18141), .B(n18140), .Z(n18283) );
  NAND U20098 ( .A(n18143), .B(n18142), .Z(n18147) );
  NAND U20099 ( .A(n18145), .B(n18144), .Z(n18146) );
  NAND U20100 ( .A(n18147), .B(n18146), .Z(n18282) );
  NAND U20101 ( .A(n18149), .B(n18148), .Z(n18153) );
  NAND U20102 ( .A(n18151), .B(n18150), .Z(n18152) );
  AND U20103 ( .A(n18153), .B(n18152), .Z(n18315) );
  NAND U20104 ( .A(x[501]), .B(y[7848]), .Z(n19139) );
  NANDN U20105 ( .A(n19139), .B(n18154), .Z(n18158) );
  NAND U20106 ( .A(n18156), .B(n18155), .Z(n18157) );
  NAND U20107 ( .A(n18158), .B(n18157), .Z(n18389) );
  NAND U20108 ( .A(x[502]), .B(y[7843]), .Z(n18358) );
  NAND U20109 ( .A(x[485]), .B(y[7860]), .Z(n18357) );
  NAND U20110 ( .A(x[497]), .B(y[7848]), .Z(n18356) );
  XOR U20111 ( .A(n18357), .B(n18356), .Z(n18359) );
  XNOR U20112 ( .A(n18358), .B(n18359), .Z(n18388) );
  AND U20113 ( .A(y[7845]), .B(x[500]), .Z(n18160) );
  NAND U20114 ( .A(y[7844]), .B(x[501]), .Z(n18159) );
  XNOR U20115 ( .A(n18160), .B(n18159), .Z(n18371) );
  AND U20116 ( .A(x[499]), .B(y[7846]), .Z(n18370) );
  XOR U20117 ( .A(n18371), .B(n18370), .Z(n18387) );
  XNOR U20118 ( .A(n18388), .B(n18387), .Z(n18390) );
  XOR U20119 ( .A(n18389), .B(n18390), .Z(n18313) );
  NAND U20120 ( .A(n18369), .B(n18538), .Z(n18164) );
  NAND U20121 ( .A(n18162), .B(n18161), .Z(n18163) );
  NAND U20122 ( .A(n18164), .B(n18163), .Z(n18395) );
  NAND U20123 ( .A(x[495]), .B(y[7850]), .Z(n18377) );
  NAND U20124 ( .A(x[498]), .B(y[7847]), .Z(n18376) );
  NAND U20125 ( .A(x[486]), .B(y[7859]), .Z(n18375) );
  XOR U20126 ( .A(n18376), .B(n18375), .Z(n18378) );
  XNOR U20127 ( .A(n18377), .B(n18378), .Z(n18394) );
  NAND U20128 ( .A(x[503]), .B(y[7842]), .Z(n18352) );
  NAND U20129 ( .A(x[484]), .B(y[7861]), .Z(n18351) );
  NAND U20130 ( .A(x[496]), .B(y[7849]), .Z(n18350) );
  XOR U20131 ( .A(n18351), .B(n18350), .Z(n18353) );
  XNOR U20132 ( .A(n18352), .B(n18353), .Z(n18393) );
  XNOR U20133 ( .A(n18394), .B(n18393), .Z(n18396) );
  XOR U20134 ( .A(n18395), .B(n18396), .Z(n18312) );
  XOR U20135 ( .A(n18313), .B(n18312), .Z(n18314) );
  XNOR U20136 ( .A(n18315), .B(n18314), .Z(n18327) );
  NAND U20137 ( .A(n18166), .B(n18165), .Z(n18170) );
  NAND U20138 ( .A(n18168), .B(n18167), .Z(n18169) );
  NAND U20139 ( .A(n18170), .B(n18169), .Z(n18325) );
  NAND U20140 ( .A(n18172), .B(n18171), .Z(n18176) );
  NAND U20141 ( .A(n18174), .B(n18173), .Z(n18175) );
  NAND U20142 ( .A(n18176), .B(n18175), .Z(n18324) );
  XOR U20143 ( .A(n18325), .B(n18324), .Z(n18326) );
  XOR U20144 ( .A(n18327), .B(n18326), .Z(n18284) );
  XOR U20145 ( .A(n18285), .B(n18284), .Z(n18277) );
  NAND U20146 ( .A(n18178), .B(n18177), .Z(n18182) );
  NAND U20147 ( .A(n18180), .B(n18179), .Z(n18181) );
  NAND U20148 ( .A(n18182), .B(n18181), .Z(n18276) );
  XOR U20149 ( .A(n18278), .B(n18279), .Z(n18273) );
  NANDN U20150 ( .A(n18294), .B(n18183), .Z(n18187) );
  NAND U20151 ( .A(n18185), .B(n18184), .Z(n18186) );
  NAND U20152 ( .A(n18187), .B(n18186), .Z(n18319) );
  NAND U20153 ( .A(x[494]), .B(y[7856]), .Z(n19209) );
  NANDN U20154 ( .A(n19209), .B(n18188), .Z(n18192) );
  NANDN U20155 ( .A(n18190), .B(n18189), .Z(n18191) );
  NAND U20156 ( .A(n18192), .B(n18191), .Z(n18346) );
  NAND U20157 ( .A(x[491]), .B(y[7854]), .Z(n18365) );
  NAND U20158 ( .A(x[492]), .B(y[7853]), .Z(n18364) );
  NAND U20159 ( .A(x[487]), .B(y[7858]), .Z(n18363) );
  XOR U20160 ( .A(n18364), .B(n18363), .Z(n18366) );
  XOR U20161 ( .A(n18365), .B(n18366), .Z(n18345) );
  AND U20162 ( .A(x[504]), .B(y[7841]), .Z(n18362) );
  XOR U20163 ( .A(o[185]), .B(n18362), .Z(n18333) );
  AND U20164 ( .A(x[481]), .B(y[7864]), .Z(n18332) );
  XOR U20165 ( .A(n18333), .B(n18332), .Z(n18335) );
  AND U20166 ( .A(x[493]), .B(y[7852]), .Z(n18334) );
  XOR U20167 ( .A(n18335), .B(n18334), .Z(n18344) );
  XOR U20168 ( .A(n18346), .B(n18347), .Z(n18318) );
  XOR U20169 ( .A(n18319), .B(n18318), .Z(n18321) );
  AND U20170 ( .A(n18194), .B(n18193), .Z(n18198) );
  NAND U20171 ( .A(n18196), .B(n18195), .Z(n18197) );
  NANDN U20172 ( .A(n18198), .B(n18197), .Z(n18307) );
  AND U20173 ( .A(n18200), .B(n18199), .Z(n18204) );
  NAND U20174 ( .A(n18202), .B(n18201), .Z(n18203) );
  NANDN U20175 ( .A(n18204), .B(n18203), .Z(n18306) );
  XOR U20176 ( .A(n18307), .B(n18306), .Z(n18308) );
  NAND U20177 ( .A(n18206), .B(n18205), .Z(n18210) );
  NAND U20178 ( .A(n18208), .B(n18207), .Z(n18209) );
  NAND U20179 ( .A(n18210), .B(n18209), .Z(n18302) );
  NAND U20180 ( .A(x[488]), .B(y[7857]), .Z(n18296) );
  XOR U20181 ( .A(n18295), .B(n18294), .Z(n18297) );
  XNOR U20182 ( .A(n18296), .B(n18297), .Z(n18301) );
  NAND U20183 ( .A(n18211), .B(o[184]), .Z(n18290) );
  NAND U20184 ( .A(x[505]), .B(y[7840]), .Z(n18289) );
  NAND U20185 ( .A(x[480]), .B(y[7865]), .Z(n18288) );
  XOR U20186 ( .A(n18289), .B(n18288), .Z(n18291) );
  XNOR U20187 ( .A(n18290), .B(n18291), .Z(n18300) );
  XNOR U20188 ( .A(n18301), .B(n18300), .Z(n18303) );
  XOR U20189 ( .A(n18302), .B(n18303), .Z(n18309) );
  XNOR U20190 ( .A(n18308), .B(n18309), .Z(n18320) );
  XOR U20191 ( .A(n18321), .B(n18320), .Z(n18402) );
  AND U20192 ( .A(n18213), .B(n18212), .Z(n18217) );
  NAND U20193 ( .A(n18215), .B(n18214), .Z(n18216) );
  NANDN U20194 ( .A(n18217), .B(n18216), .Z(n18384) );
  NAND U20195 ( .A(n18219), .B(n18218), .Z(n18223) );
  NAND U20196 ( .A(n18221), .B(n18220), .Z(n18222) );
  NAND U20197 ( .A(n18223), .B(n18222), .Z(n18382) );
  AND U20198 ( .A(x[494]), .B(y[7851]), .Z(n18339) );
  AND U20199 ( .A(x[482]), .B(y[7863]), .Z(n18338) );
  XOR U20200 ( .A(n18339), .B(n18338), .Z(n18341) );
  AND U20201 ( .A(x[483]), .B(y[7862]), .Z(n18340) );
  XOR U20202 ( .A(n18341), .B(n18340), .Z(n18381) );
  XOR U20203 ( .A(n18382), .B(n18381), .Z(n18383) );
  XNOR U20204 ( .A(n18384), .B(n18383), .Z(n18399) );
  NAND U20205 ( .A(n18225), .B(n18224), .Z(n18229) );
  NAND U20206 ( .A(n18227), .B(n18226), .Z(n18228) );
  AND U20207 ( .A(n18229), .B(n18228), .Z(n18400) );
  XOR U20208 ( .A(n18399), .B(n18400), .Z(n18401) );
  NAND U20209 ( .A(n18231), .B(n18230), .Z(n18235) );
  NAND U20210 ( .A(n18233), .B(n18232), .Z(n18234) );
  NAND U20211 ( .A(n18235), .B(n18234), .Z(n18406) );
  NANDN U20212 ( .A(n18237), .B(n18236), .Z(n18241) );
  NANDN U20213 ( .A(n18239), .B(n18238), .Z(n18240) );
  NAND U20214 ( .A(n18241), .B(n18240), .Z(n18408) );
  NAND U20215 ( .A(n18243), .B(n18242), .Z(n18247) );
  NAND U20216 ( .A(n18245), .B(n18244), .Z(n18246) );
  AND U20217 ( .A(n18247), .B(n18246), .Z(n18270) );
  NAND U20218 ( .A(n18249), .B(n18248), .Z(n18253) );
  NAND U20219 ( .A(n18251), .B(n18250), .Z(n18252) );
  NAND U20220 ( .A(n18253), .B(n18252), .Z(n18415) );
  XOR U20221 ( .A(n18416), .B(n18415), .Z(n18418) );
  NAND U20222 ( .A(n18255), .B(n18254), .Z(n18259) );
  NAND U20223 ( .A(n18257), .B(n18256), .Z(n18258) );
  AND U20224 ( .A(n18259), .B(n18258), .Z(n18417) );
  XNOR U20225 ( .A(n18418), .B(n18417), .Z(n18414) );
  NANDN U20226 ( .A(n18264), .B(n18263), .Z(n18268) );
  NAND U20227 ( .A(n18266), .B(n18265), .Z(n18267) );
  AND U20228 ( .A(n18268), .B(n18267), .Z(n18413) );
  IV U20229 ( .A(n18413), .Z(n18411) );
  XOR U20230 ( .A(n18412), .B(n18411), .Z(n18269) );
  XNOR U20231 ( .A(n18414), .B(n18269), .Z(N378) );
  NANDN U20232 ( .A(n18271), .B(n18270), .Z(n18275) );
  NANDN U20233 ( .A(n18273), .B(n18272), .Z(n18274) );
  NAND U20234 ( .A(n18275), .B(n18274), .Z(n18573) );
  NANDN U20235 ( .A(n18277), .B(n18276), .Z(n18281) );
  NAND U20236 ( .A(n18279), .B(n18278), .Z(n18280) );
  AND U20237 ( .A(n18281), .B(n18280), .Z(n18574) );
  XOR U20238 ( .A(n18573), .B(n18574), .Z(n18576) );
  NANDN U20239 ( .A(n18283), .B(n18282), .Z(n18287) );
  NAND U20240 ( .A(n18285), .B(n18284), .Z(n18286) );
  AND U20241 ( .A(n18287), .B(n18286), .Z(n18567) );
  AND U20242 ( .A(x[482]), .B(y[7864]), .Z(n18440) );
  XOR U20243 ( .A(n18441), .B(n18440), .Z(n18443) );
  AND U20244 ( .A(x[504]), .B(y[7842]), .Z(n18442) );
  XOR U20245 ( .A(n18443), .B(n18442), .Z(n18477) );
  NAND U20246 ( .A(n18289), .B(n18288), .Z(n18293) );
  NAND U20247 ( .A(n18291), .B(n18290), .Z(n18292) );
  AND U20248 ( .A(n18293), .B(n18292), .Z(n18476) );
  XOR U20249 ( .A(n18477), .B(n18476), .Z(n18479) );
  NAND U20250 ( .A(n18295), .B(n18294), .Z(n18299) );
  NAND U20251 ( .A(n18297), .B(n18296), .Z(n18298) );
  AND U20252 ( .A(n18299), .B(n18298), .Z(n18478) );
  XNOR U20253 ( .A(n18479), .B(n18478), .Z(n18515) );
  NAND U20254 ( .A(n18301), .B(n18300), .Z(n18305) );
  NANDN U20255 ( .A(n18303), .B(n18302), .Z(n18304) );
  AND U20256 ( .A(n18305), .B(n18304), .Z(n18514) );
  XOR U20257 ( .A(n18515), .B(n18514), .Z(n18517) );
  NAND U20258 ( .A(n18307), .B(n18306), .Z(n18311) );
  NANDN U20259 ( .A(n18309), .B(n18308), .Z(n18310) );
  AND U20260 ( .A(n18311), .B(n18310), .Z(n18516) );
  XOR U20261 ( .A(n18517), .B(n18516), .Z(n18561) );
  NAND U20262 ( .A(n18313), .B(n18312), .Z(n18317) );
  NAND U20263 ( .A(n18315), .B(n18314), .Z(n18316) );
  NAND U20264 ( .A(n18317), .B(n18316), .Z(n18559) );
  NAND U20265 ( .A(n18319), .B(n18318), .Z(n18323) );
  NAND U20266 ( .A(n18321), .B(n18320), .Z(n18322) );
  AND U20267 ( .A(n18323), .B(n18322), .Z(n18558) );
  XOR U20268 ( .A(n18559), .B(n18558), .Z(n18560) );
  XOR U20269 ( .A(n18561), .B(n18560), .Z(n18565) );
  NAND U20270 ( .A(n18325), .B(n18324), .Z(n18329) );
  NAND U20271 ( .A(n18327), .B(n18326), .Z(n18328) );
  NAND U20272 ( .A(n18329), .B(n18328), .Z(n18511) );
  AND U20273 ( .A(y[7860]), .B(x[486]), .Z(n18331) );
  NAND U20274 ( .A(y[7858]), .B(x[488]), .Z(n18330) );
  XNOR U20275 ( .A(n18331), .B(n18330), .Z(n18540) );
  AND U20276 ( .A(x[489]), .B(y[7857]), .Z(n18539) );
  XOR U20277 ( .A(n18540), .B(n18539), .Z(n18520) );
  AND U20278 ( .A(x[487]), .B(y[7859]), .Z(n18521) );
  XOR U20279 ( .A(n18520), .B(n18521), .Z(n18523) );
  AND U20280 ( .A(x[492]), .B(y[7854]), .Z(n18634) );
  AND U20281 ( .A(x[485]), .B(y[7861]), .Z(n18491) );
  XOR U20282 ( .A(n18634), .B(n18491), .Z(n18493) );
  AND U20283 ( .A(x[490]), .B(y[7856]), .Z(n18492) );
  XOR U20284 ( .A(n18493), .B(n18492), .Z(n18522) );
  XOR U20285 ( .A(n18523), .B(n18522), .Z(n18467) );
  NAND U20286 ( .A(n18333), .B(n18332), .Z(n18337) );
  NAND U20287 ( .A(n18335), .B(n18334), .Z(n18336) );
  NAND U20288 ( .A(n18337), .B(n18336), .Z(n18465) );
  NAND U20289 ( .A(n18339), .B(n18338), .Z(n18343) );
  NAND U20290 ( .A(n18341), .B(n18340), .Z(n18342) );
  NAND U20291 ( .A(n18343), .B(n18342), .Z(n18464) );
  XOR U20292 ( .A(n18465), .B(n18464), .Z(n18466) );
  XNOR U20293 ( .A(n18467), .B(n18466), .Z(n18503) );
  NANDN U20294 ( .A(n18345), .B(n18344), .Z(n18349) );
  NAND U20295 ( .A(n18347), .B(n18346), .Z(n18348) );
  AND U20296 ( .A(n18349), .B(n18348), .Z(n18502) );
  XOR U20297 ( .A(n18503), .B(n18502), .Z(n18505) );
  NAND U20298 ( .A(n18351), .B(n18350), .Z(n18355) );
  NAND U20299 ( .A(n18353), .B(n18352), .Z(n18354) );
  AND U20300 ( .A(n18355), .B(n18354), .Z(n18428) );
  NAND U20301 ( .A(n18357), .B(n18356), .Z(n18361) );
  NAND U20302 ( .A(n18359), .B(n18358), .Z(n18360) );
  AND U20303 ( .A(n18361), .B(n18360), .Z(n18429) );
  XOR U20304 ( .A(n18428), .B(n18429), .Z(n18431) );
  AND U20305 ( .A(n18362), .B(o[185]), .Z(n18532) );
  AND U20306 ( .A(x[494]), .B(y[7852]), .Z(n18533) );
  XOR U20307 ( .A(n18532), .B(n18533), .Z(n18534) );
  AND U20308 ( .A(x[481]), .B(y[7865]), .Z(n18535) );
  XOR U20309 ( .A(n18534), .B(n18535), .Z(n18483) );
  AND U20310 ( .A(x[505]), .B(y[7841]), .Z(n18543) );
  XOR U20311 ( .A(o[186]), .B(n18543), .Z(n18497) );
  AND U20312 ( .A(x[506]), .B(y[7840]), .Z(n18496) );
  XOR U20313 ( .A(n18497), .B(n18496), .Z(n18499) );
  AND U20314 ( .A(x[480]), .B(y[7866]), .Z(n18498) );
  XOR U20315 ( .A(n18499), .B(n18498), .Z(n18482) );
  XOR U20316 ( .A(n18483), .B(n18482), .Z(n18485) );
  NAND U20317 ( .A(n18364), .B(n18363), .Z(n18368) );
  NAND U20318 ( .A(n18366), .B(n18365), .Z(n18367) );
  AND U20319 ( .A(n18368), .B(n18367), .Z(n18484) );
  XOR U20320 ( .A(n18485), .B(n18484), .Z(n18430) );
  XNOR U20321 ( .A(n18431), .B(n18430), .Z(n18473) );
  AND U20322 ( .A(x[501]), .B(y[7845]), .Z(n18374) );
  IV U20323 ( .A(n18374), .Z(n18526) );
  NANDN U20324 ( .A(n18526), .B(n18369), .Z(n18373) );
  NAND U20325 ( .A(n18371), .B(n18370), .Z(n18372) );
  NAND U20326 ( .A(n18373), .B(n18372), .Z(n18461) );
  XOR U20327 ( .A(n18527), .B(n18374), .Z(n18528) );
  AND U20328 ( .A(x[500]), .B(y[7846]), .Z(n18529) );
  XOR U20329 ( .A(n18528), .B(n18529), .Z(n18459) );
  AND U20330 ( .A(x[503]), .B(y[7843]), .Z(n18447) );
  XOR U20331 ( .A(n18446), .B(n18447), .Z(n18448) );
  AND U20332 ( .A(x[502]), .B(y[7844]), .Z(n18449) );
  XOR U20333 ( .A(n18448), .B(n18449), .Z(n18458) );
  XOR U20334 ( .A(n18459), .B(n18458), .Z(n18460) );
  XNOR U20335 ( .A(n18461), .B(n18460), .Z(n18471) );
  AND U20336 ( .A(x[484]), .B(y[7862]), .Z(n18452) );
  XOR U20337 ( .A(n18453), .B(n18452), .Z(n18454) );
  XNOR U20338 ( .A(n18454), .B(n18455), .Z(n18435) );
  AND U20339 ( .A(x[483]), .B(y[7863]), .Z(n18544) );
  AND U20340 ( .A(x[499]), .B(y[7847]), .Z(n18545) );
  XOR U20341 ( .A(n18544), .B(n18545), .Z(n18546) );
  AND U20342 ( .A(x[491]), .B(y[7855]), .Z(n18547) );
  XOR U20343 ( .A(n18546), .B(n18547), .Z(n18434) );
  XOR U20344 ( .A(n18435), .B(n18434), .Z(n18437) );
  NAND U20345 ( .A(n18376), .B(n18375), .Z(n18380) );
  NAND U20346 ( .A(n18378), .B(n18377), .Z(n18379) );
  AND U20347 ( .A(n18380), .B(n18379), .Z(n18436) );
  XNOR U20348 ( .A(n18437), .B(n18436), .Z(n18470) );
  XOR U20349 ( .A(n18471), .B(n18470), .Z(n18472) );
  XOR U20350 ( .A(n18473), .B(n18472), .Z(n18504) );
  XNOR U20351 ( .A(n18505), .B(n18504), .Z(n18509) );
  NAND U20352 ( .A(n18382), .B(n18381), .Z(n18386) );
  NAND U20353 ( .A(n18384), .B(n18383), .Z(n18385) );
  NAND U20354 ( .A(n18386), .B(n18385), .Z(n18555) );
  NAND U20355 ( .A(n18388), .B(n18387), .Z(n18392) );
  NANDN U20356 ( .A(n18390), .B(n18389), .Z(n18391) );
  NAND U20357 ( .A(n18392), .B(n18391), .Z(n18553) );
  NAND U20358 ( .A(n18394), .B(n18393), .Z(n18398) );
  NANDN U20359 ( .A(n18396), .B(n18395), .Z(n18397) );
  NAND U20360 ( .A(n18398), .B(n18397), .Z(n18552) );
  XOR U20361 ( .A(n18553), .B(n18552), .Z(n18554) );
  XOR U20362 ( .A(n18555), .B(n18554), .Z(n18508) );
  XOR U20363 ( .A(n18509), .B(n18508), .Z(n18510) );
  XOR U20364 ( .A(n18511), .B(n18510), .Z(n18564) );
  NAND U20365 ( .A(n18400), .B(n18399), .Z(n18404) );
  NANDN U20366 ( .A(n18402), .B(n18401), .Z(n18403) );
  AND U20367 ( .A(n18404), .B(n18403), .Z(n18422) );
  NANDN U20368 ( .A(n18406), .B(n18405), .Z(n18410) );
  NANDN U20369 ( .A(n18408), .B(n18407), .Z(n18409) );
  NAND U20370 ( .A(n18410), .B(n18409), .Z(n18423) );
  XOR U20371 ( .A(n18425), .B(n18424), .Z(n18575) );
  XOR U20372 ( .A(n18576), .B(n18575), .Z(n18572) );
  NAND U20373 ( .A(n18416), .B(n18415), .Z(n18420) );
  NAND U20374 ( .A(n18418), .B(n18417), .Z(n18419) );
  NAND U20375 ( .A(n18420), .B(n18419), .Z(n18570) );
  XOR U20376 ( .A(n18571), .B(n18570), .Z(n18421) );
  XNOR U20377 ( .A(n18572), .B(n18421), .Z(N379) );
  NANDN U20378 ( .A(n18423), .B(n18422), .Z(n18427) );
  NAND U20379 ( .A(n18425), .B(n18424), .Z(n18426) );
  AND U20380 ( .A(n18427), .B(n18426), .Z(n18734) );
  NAND U20381 ( .A(n18429), .B(n18428), .Z(n18433) );
  NAND U20382 ( .A(n18431), .B(n18430), .Z(n18432) );
  NAND U20383 ( .A(n18433), .B(n18432), .Z(n18709) );
  NAND U20384 ( .A(n18435), .B(n18434), .Z(n18439) );
  NAND U20385 ( .A(n18437), .B(n18436), .Z(n18438) );
  NAND U20386 ( .A(n18439), .B(n18438), .Z(n18707) );
  AND U20387 ( .A(n18441), .B(n18440), .Z(n18445) );
  NAND U20388 ( .A(n18443), .B(n18442), .Z(n18444) );
  NANDN U20389 ( .A(n18445), .B(n18444), .Z(n18605) );
  NAND U20390 ( .A(n18447), .B(n18446), .Z(n18451) );
  NAND U20391 ( .A(n18449), .B(n18448), .Z(n18450) );
  NAND U20392 ( .A(n18451), .B(n18450), .Z(n18604) );
  XOR U20393 ( .A(n18605), .B(n18604), .Z(n18606) );
  AND U20394 ( .A(n18453), .B(n18452), .Z(n18457) );
  NANDN U20395 ( .A(n18455), .B(n18454), .Z(n18456) );
  NANDN U20396 ( .A(n18457), .B(n18456), .Z(n18618) );
  AND U20397 ( .A(x[480]), .B(y[7867]), .Z(n18696) );
  AND U20398 ( .A(x[507]), .B(y[7840]), .Z(n18695) );
  XOR U20399 ( .A(n18696), .B(n18695), .Z(n18698) );
  AND U20400 ( .A(x[506]), .B(y[7841]), .Z(n18686) );
  XOR U20401 ( .A(n18686), .B(o[187]), .Z(n18697) );
  XOR U20402 ( .A(n18698), .B(n18697), .Z(n18617) );
  AND U20403 ( .A(x[489]), .B(y[7858]), .Z(n18681) );
  AND U20404 ( .A(x[501]), .B(y[7846]), .Z(n18680) );
  XOR U20405 ( .A(n18681), .B(n18680), .Z(n18683) );
  AND U20406 ( .A(x[498]), .B(y[7849]), .Z(n18682) );
  XOR U20407 ( .A(n18683), .B(n18682), .Z(n18616) );
  XOR U20408 ( .A(n18617), .B(n18616), .Z(n18619) );
  XNOR U20409 ( .A(n18618), .B(n18619), .Z(n18607) );
  XOR U20410 ( .A(n18707), .B(n18708), .Z(n18710) );
  XOR U20411 ( .A(n18709), .B(n18710), .Z(n18728) );
  NAND U20412 ( .A(n18459), .B(n18458), .Z(n18463) );
  NAND U20413 ( .A(n18461), .B(n18460), .Z(n18462) );
  AND U20414 ( .A(n18463), .B(n18462), .Z(n18726) );
  NAND U20415 ( .A(n18465), .B(n18464), .Z(n18469) );
  NAND U20416 ( .A(n18467), .B(n18466), .Z(n18468) );
  AND U20417 ( .A(n18469), .B(n18468), .Z(n18725) );
  XOR U20418 ( .A(n18726), .B(n18725), .Z(n18727) );
  NAND U20419 ( .A(n18471), .B(n18470), .Z(n18475) );
  NAND U20420 ( .A(n18473), .B(n18472), .Z(n18474) );
  AND U20421 ( .A(n18475), .B(n18474), .Z(n18713) );
  NAND U20422 ( .A(n18477), .B(n18476), .Z(n18481) );
  NAND U20423 ( .A(n18479), .B(n18478), .Z(n18480) );
  NAND U20424 ( .A(n18481), .B(n18480), .Z(n18703) );
  NAND U20425 ( .A(n18483), .B(n18482), .Z(n18487) );
  NAND U20426 ( .A(n18485), .B(n18484), .Z(n18486) );
  NAND U20427 ( .A(n18487), .B(n18486), .Z(n18701) );
  AND U20428 ( .A(x[499]), .B(y[7848]), .Z(n18675) );
  AND U20429 ( .A(x[505]), .B(y[7842]), .Z(n18674) );
  XOR U20430 ( .A(n18675), .B(n18674), .Z(n18677) );
  AND U20431 ( .A(x[486]), .B(y[7861]), .Z(n18676) );
  XOR U20432 ( .A(n18677), .B(n18676), .Z(n18664) );
  AND U20433 ( .A(x[495]), .B(y[7852]), .Z(n18640) );
  AND U20434 ( .A(x[482]), .B(y[7865]), .Z(n18639) );
  XOR U20435 ( .A(n18640), .B(n18639), .Z(n18642) );
  AND U20436 ( .A(x[483]), .B(y[7864]), .Z(n18641) );
  XOR U20437 ( .A(n18642), .B(n18641), .Z(n18663) );
  XOR U20438 ( .A(n18664), .B(n18663), .Z(n18665) );
  NAND U20439 ( .A(x[496]), .B(y[7851]), .Z(n18622) );
  XOR U20440 ( .A(n18622), .B(n18488), .Z(n18625) );
  XOR U20441 ( .A(n18624), .B(n18625), .Z(n18636) );
  AND U20442 ( .A(y[7854]), .B(x[493]), .Z(n18490) );
  AND U20443 ( .A(y[7855]), .B(x[492]), .Z(n18489) );
  XOR U20444 ( .A(n18490), .B(n18489), .Z(n18635) );
  XNOR U20445 ( .A(n18665), .B(n18666), .Z(n18601) );
  AND U20446 ( .A(n18634), .B(n18491), .Z(n18495) );
  NAND U20447 ( .A(n18493), .B(n18492), .Z(n18494) );
  NANDN U20448 ( .A(n18495), .B(n18494), .Z(n18599) );
  NAND U20449 ( .A(n18497), .B(n18496), .Z(n18501) );
  NAND U20450 ( .A(n18499), .B(n18498), .Z(n18500) );
  NAND U20451 ( .A(n18501), .B(n18500), .Z(n18598) );
  XOR U20452 ( .A(n18599), .B(n18598), .Z(n18600) );
  XOR U20453 ( .A(n18601), .B(n18600), .Z(n18702) );
  XNOR U20454 ( .A(n18701), .B(n18702), .Z(n18704) );
  XNOR U20455 ( .A(n18713), .B(n18714), .Z(n18716) );
  NAND U20456 ( .A(n18503), .B(n18502), .Z(n18507) );
  NAND U20457 ( .A(n18505), .B(n18504), .Z(n18506) );
  AND U20458 ( .A(n18507), .B(n18506), .Z(n18715) );
  XOR U20459 ( .A(n18716), .B(n18715), .Z(n18586) );
  NAND U20460 ( .A(n18509), .B(n18508), .Z(n18513) );
  NAND U20461 ( .A(n18511), .B(n18510), .Z(n18512) );
  NAND U20462 ( .A(n18513), .B(n18512), .Z(n18588) );
  XOR U20463 ( .A(n18589), .B(n18588), .Z(n18583) );
  NAND U20464 ( .A(n18515), .B(n18514), .Z(n18519) );
  NAND U20465 ( .A(n18517), .B(n18516), .Z(n18518) );
  NAND U20466 ( .A(n18519), .B(n18518), .Z(n18593) );
  NAND U20467 ( .A(n18521), .B(n18520), .Z(n18525) );
  NAND U20468 ( .A(n18523), .B(n18522), .Z(n18524) );
  NAND U20469 ( .A(n18525), .B(n18524), .Z(n18721) );
  ANDN U20470 ( .B(n18527), .A(n18526), .Z(n18531) );
  NAND U20471 ( .A(n18529), .B(n18528), .Z(n18530) );
  NANDN U20472 ( .A(n18531), .B(n18530), .Z(n18652) );
  NAND U20473 ( .A(n18533), .B(n18532), .Z(n18537) );
  NAND U20474 ( .A(n18535), .B(n18534), .Z(n18536) );
  NAND U20475 ( .A(n18537), .B(n18536), .Z(n18651) );
  XOR U20476 ( .A(n18652), .B(n18651), .Z(n18653) );
  AND U20477 ( .A(y[7860]), .B(x[488]), .Z(n18688) );
  NAND U20478 ( .A(n18538), .B(n18688), .Z(n18542) );
  NAND U20479 ( .A(n18540), .B(n18539), .Z(n18541) );
  NAND U20480 ( .A(n18542), .B(n18541), .Z(n18612) );
  AND U20481 ( .A(x[494]), .B(y[7853]), .Z(n18646) );
  AND U20482 ( .A(x[481]), .B(y[7866]), .Z(n18645) );
  XOR U20483 ( .A(n18646), .B(n18645), .Z(n18648) );
  AND U20484 ( .A(o[186]), .B(n18543), .Z(n18647) );
  XOR U20485 ( .A(n18648), .B(n18647), .Z(n18611) );
  AND U20486 ( .A(x[497]), .B(y[7850]), .Z(n18690) );
  AND U20487 ( .A(x[484]), .B(y[7863]), .Z(n18689) );
  XOR U20488 ( .A(n18690), .B(n18689), .Z(n18692) );
  AND U20489 ( .A(x[485]), .B(y[7862]), .Z(n18691) );
  XOR U20490 ( .A(n18692), .B(n18691), .Z(n18610) );
  XOR U20491 ( .A(n18611), .B(n18610), .Z(n18613) );
  XNOR U20492 ( .A(n18612), .B(n18613), .Z(n18654) );
  NAND U20493 ( .A(n18545), .B(n18544), .Z(n18549) );
  NAND U20494 ( .A(n18547), .B(n18546), .Z(n18548) );
  NAND U20495 ( .A(n18549), .B(n18548), .Z(n18659) );
  AND U20496 ( .A(y[7843]), .B(x[504]), .Z(n18551) );
  NAND U20497 ( .A(y[7847]), .B(x[500]), .Z(n18550) );
  XNOR U20498 ( .A(n18551), .B(n18550), .Z(n18671) );
  AND U20499 ( .A(x[487]), .B(y[7860]), .Z(n18670) );
  XOR U20500 ( .A(n18671), .B(n18670), .Z(n18658) );
  AND U20501 ( .A(x[488]), .B(y[7859]), .Z(n18629) );
  AND U20502 ( .A(x[503]), .B(y[7844]), .Z(n18628) );
  XOR U20503 ( .A(n18629), .B(n18628), .Z(n18631) );
  AND U20504 ( .A(x[502]), .B(y[7845]), .Z(n18630) );
  XOR U20505 ( .A(n18631), .B(n18630), .Z(n18657) );
  XOR U20506 ( .A(n18658), .B(n18657), .Z(n18660) );
  XOR U20507 ( .A(n18659), .B(n18660), .Z(n18719) );
  XOR U20508 ( .A(n18720), .B(n18719), .Z(n18722) );
  XNOR U20509 ( .A(n18721), .B(n18722), .Z(n18592) );
  XOR U20510 ( .A(n18593), .B(n18592), .Z(n18595) );
  NAND U20511 ( .A(n18553), .B(n18552), .Z(n18557) );
  NAND U20512 ( .A(n18555), .B(n18554), .Z(n18556) );
  AND U20513 ( .A(n18557), .B(n18556), .Z(n18594) );
  XNOR U20514 ( .A(n18595), .B(n18594), .Z(n18581) );
  NAND U20515 ( .A(n18559), .B(n18558), .Z(n18563) );
  NAND U20516 ( .A(n18561), .B(n18560), .Z(n18562) );
  AND U20517 ( .A(n18563), .B(n18562), .Z(n18580) );
  XOR U20518 ( .A(n18581), .B(n18580), .Z(n18582) );
  XOR U20519 ( .A(n18583), .B(n18582), .Z(n18732) );
  NANDN U20520 ( .A(n18565), .B(n18564), .Z(n18569) );
  NANDN U20521 ( .A(n18567), .B(n18566), .Z(n18568) );
  AND U20522 ( .A(n18569), .B(n18568), .Z(n18731) );
  XNOR U20523 ( .A(n18734), .B(n18733), .Z(n18739) );
  NAND U20524 ( .A(n18574), .B(n18573), .Z(n18578) );
  NAND U20525 ( .A(n18576), .B(n18575), .Z(n18577) );
  AND U20526 ( .A(n18578), .B(n18577), .Z(n18737) );
  XOR U20527 ( .A(n18738), .B(n18737), .Z(n18579) );
  XNOR U20528 ( .A(n18739), .B(n18579), .Z(N380) );
  NAND U20529 ( .A(n18581), .B(n18580), .Z(n18585) );
  NAND U20530 ( .A(n18583), .B(n18582), .Z(n18584) );
  NAND U20531 ( .A(n18585), .B(n18584), .Z(n18900) );
  NANDN U20532 ( .A(n18587), .B(n18586), .Z(n18591) );
  NAND U20533 ( .A(n18589), .B(n18588), .Z(n18590) );
  NAND U20534 ( .A(n18591), .B(n18590), .Z(n18899) );
  XOR U20535 ( .A(n18900), .B(n18899), .Z(n18902) );
  NAND U20536 ( .A(n18593), .B(n18592), .Z(n18597) );
  NAND U20537 ( .A(n18595), .B(n18594), .Z(n18596) );
  AND U20538 ( .A(n18597), .B(n18596), .Z(n18741) );
  NAND U20539 ( .A(n18599), .B(n18598), .Z(n18603) );
  NAND U20540 ( .A(n18601), .B(n18600), .Z(n18602) );
  NAND U20541 ( .A(n18603), .B(n18602), .Z(n18765) );
  NAND U20542 ( .A(n18605), .B(n18604), .Z(n18609) );
  NANDN U20543 ( .A(n18607), .B(n18606), .Z(n18608) );
  NAND U20544 ( .A(n18609), .B(n18608), .Z(n18871) );
  NAND U20545 ( .A(n18611), .B(n18610), .Z(n18615) );
  NAND U20546 ( .A(n18613), .B(n18612), .Z(n18614) );
  NAND U20547 ( .A(n18615), .B(n18614), .Z(n18870) );
  NAND U20548 ( .A(n18617), .B(n18616), .Z(n18621) );
  NAND U20549 ( .A(n18619), .B(n18618), .Z(n18620) );
  NAND U20550 ( .A(n18621), .B(n18620), .Z(n18869) );
  XOR U20551 ( .A(n18870), .B(n18869), .Z(n18872) );
  XOR U20552 ( .A(n18871), .B(n18872), .Z(n18766) );
  XOR U20553 ( .A(n18765), .B(n18766), .Z(n18768) );
  NANDN U20554 ( .A(n18623), .B(n18622), .Z(n18627) );
  NAND U20555 ( .A(n18625), .B(n18624), .Z(n18626) );
  NAND U20556 ( .A(n18627), .B(n18626), .Z(n18833) );
  AND U20557 ( .A(x[487]), .B(y[7861]), .Z(n18813) );
  AND U20558 ( .A(x[492]), .B(y[7856]), .Z(n18812) );
  XOR U20559 ( .A(n18813), .B(n18812), .Z(n18815) );
  AND U20560 ( .A(x[491]), .B(y[7857]), .Z(n18814) );
  XOR U20561 ( .A(n18815), .B(n18814), .Z(n18832) );
  AND U20562 ( .A(x[507]), .B(y[7841]), .Z(n18830) );
  XOR U20563 ( .A(o[188]), .B(n18830), .Z(n18844) );
  AND U20564 ( .A(x[506]), .B(y[7842]), .Z(n18843) );
  XOR U20565 ( .A(n18844), .B(n18843), .Z(n18846) );
  AND U20566 ( .A(x[495]), .B(y[7853]), .Z(n18845) );
  XNOR U20567 ( .A(n18846), .B(n18845), .Z(n18831) );
  XOR U20568 ( .A(n18833), .B(n18834), .Z(n18876) );
  NAND U20569 ( .A(n18629), .B(n18628), .Z(n18633) );
  NAND U20570 ( .A(n18631), .B(n18630), .Z(n18632) );
  NAND U20571 ( .A(n18633), .B(n18632), .Z(n18853) );
  AND U20572 ( .A(x[497]), .B(y[7851]), .Z(n18778) );
  AND U20573 ( .A(x[502]), .B(y[7846]), .Z(n18777) );
  XOR U20574 ( .A(n18778), .B(n18777), .Z(n18780) );
  AND U20575 ( .A(x[484]), .B(y[7864]), .Z(n18779) );
  XOR U20576 ( .A(n18780), .B(n18779), .Z(n18852) );
  AND U20577 ( .A(x[486]), .B(y[7862]), .Z(n19014) );
  AND U20578 ( .A(x[499]), .B(y[7849]), .Z(n18819) );
  XOR U20579 ( .A(n19014), .B(n18819), .Z(n18821) );
  XOR U20580 ( .A(n18821), .B(n18820), .Z(n18851) );
  XOR U20581 ( .A(n18852), .B(n18851), .Z(n18854) );
  XOR U20582 ( .A(n18853), .B(n18854), .Z(n18875) );
  NAND U20583 ( .A(n18838), .B(n18634), .Z(n18638) );
  NANDN U20584 ( .A(n18636), .B(n18635), .Z(n18637) );
  NAND U20585 ( .A(n18638), .B(n18637), .Z(n18773) );
  NAND U20586 ( .A(n18640), .B(n18639), .Z(n18644) );
  NAND U20587 ( .A(n18642), .B(n18641), .Z(n18643) );
  NAND U20588 ( .A(n18644), .B(n18643), .Z(n18772) );
  NAND U20589 ( .A(n18646), .B(n18645), .Z(n18650) );
  NAND U20590 ( .A(n18648), .B(n18647), .Z(n18649) );
  NAND U20591 ( .A(n18650), .B(n18649), .Z(n18771) );
  XOR U20592 ( .A(n18772), .B(n18771), .Z(n18774) );
  XOR U20593 ( .A(n18773), .B(n18774), .Z(n18877) );
  XOR U20594 ( .A(n18878), .B(n18877), .Z(n18767) );
  XNOR U20595 ( .A(n18768), .B(n18767), .Z(n18762) );
  NAND U20596 ( .A(n18652), .B(n18651), .Z(n18656) );
  NANDN U20597 ( .A(n18654), .B(n18653), .Z(n18655) );
  NAND U20598 ( .A(n18656), .B(n18655), .Z(n18859) );
  NAND U20599 ( .A(n18658), .B(n18657), .Z(n18662) );
  NAND U20600 ( .A(n18660), .B(n18659), .Z(n18661) );
  NAND U20601 ( .A(n18662), .B(n18661), .Z(n18858) );
  NAND U20602 ( .A(n18664), .B(n18663), .Z(n18668) );
  NANDN U20603 ( .A(n18666), .B(n18665), .Z(n18667) );
  NAND U20604 ( .A(n18668), .B(n18667), .Z(n18857) );
  XOR U20605 ( .A(n18858), .B(n18857), .Z(n18860) );
  XOR U20606 ( .A(n18859), .B(n18860), .Z(n18760) );
  AND U20607 ( .A(x[504]), .B(y[7847]), .Z(n19229) );
  AND U20608 ( .A(x[500]), .B(y[7843]), .Z(n18669) );
  NAND U20609 ( .A(n19229), .B(n18669), .Z(n18673) );
  NAND U20610 ( .A(n18671), .B(n18670), .Z(n18672) );
  NAND U20611 ( .A(n18673), .B(n18672), .Z(n18895) );
  AND U20612 ( .A(x[505]), .B(y[7843]), .Z(n18808) );
  XOR U20613 ( .A(n18809), .B(n18808), .Z(n18807) );
  AND U20614 ( .A(x[481]), .B(y[7867]), .Z(n18806) );
  XOR U20615 ( .A(n18807), .B(n18806), .Z(n18894) );
  AND U20616 ( .A(x[496]), .B(y[7852]), .Z(n18801) );
  AND U20617 ( .A(x[504]), .B(y[7844]), .Z(n18800) );
  XOR U20618 ( .A(n18801), .B(n18800), .Z(n18803) );
  AND U20619 ( .A(x[482]), .B(y[7866]), .Z(n18802) );
  XOR U20620 ( .A(n18803), .B(n18802), .Z(n18893) );
  XOR U20621 ( .A(n18894), .B(n18893), .Z(n18896) );
  XOR U20622 ( .A(n18895), .B(n18896), .Z(n18866) );
  NAND U20623 ( .A(n18675), .B(n18674), .Z(n18679) );
  NAND U20624 ( .A(n18677), .B(n18676), .Z(n18678) );
  NAND U20625 ( .A(n18679), .B(n18678), .Z(n18889) );
  AND U20626 ( .A(x[483]), .B(y[7865]), .Z(n18837) );
  XOR U20627 ( .A(n18838), .B(n18837), .Z(n18840) );
  AND U20628 ( .A(x[503]), .B(y[7845]), .Z(n18839) );
  XOR U20629 ( .A(n18840), .B(n18839), .Z(n18888) );
  AND U20630 ( .A(x[485]), .B(y[7863]), .Z(n18825) );
  AND U20631 ( .A(x[501]), .B(y[7847]), .Z(n18824) );
  XOR U20632 ( .A(n18825), .B(n18824), .Z(n18827) );
  AND U20633 ( .A(x[500]), .B(y[7848]), .Z(n18826) );
  XOR U20634 ( .A(n18827), .B(n18826), .Z(n18887) );
  XOR U20635 ( .A(n18888), .B(n18887), .Z(n18890) );
  XOR U20636 ( .A(n18889), .B(n18890), .Z(n18864) );
  NAND U20637 ( .A(n18681), .B(n18680), .Z(n18685) );
  NAND U20638 ( .A(n18683), .B(n18682), .Z(n18684) );
  NAND U20639 ( .A(n18685), .B(n18684), .Z(n18796) );
  AND U20640 ( .A(x[480]), .B(y[7868]), .Z(n18784) );
  AND U20641 ( .A(x[508]), .B(y[7840]), .Z(n18783) );
  XOR U20642 ( .A(n18784), .B(n18783), .Z(n18786) );
  AND U20643 ( .A(n18686), .B(o[187]), .Z(n18785) );
  XOR U20644 ( .A(n18786), .B(n18785), .Z(n18795) );
  NAND U20645 ( .A(y[7858]), .B(x[490]), .Z(n18687) );
  XNOR U20646 ( .A(n18688), .B(n18687), .Z(n18791) );
  AND U20647 ( .A(x[489]), .B(y[7859]), .Z(n18790) );
  XOR U20648 ( .A(n18791), .B(n18790), .Z(n18794) );
  XOR U20649 ( .A(n18795), .B(n18794), .Z(n18797) );
  XOR U20650 ( .A(n18796), .B(n18797), .Z(n18884) );
  NAND U20651 ( .A(n18690), .B(n18689), .Z(n18694) );
  NAND U20652 ( .A(n18692), .B(n18691), .Z(n18693) );
  NAND U20653 ( .A(n18694), .B(n18693), .Z(n18882) );
  NAND U20654 ( .A(n18696), .B(n18695), .Z(n18700) );
  NAND U20655 ( .A(n18698), .B(n18697), .Z(n18699) );
  NAND U20656 ( .A(n18700), .B(n18699), .Z(n18881) );
  XOR U20657 ( .A(n18882), .B(n18881), .Z(n18883) );
  XNOR U20658 ( .A(n18884), .B(n18883), .Z(n18863) );
  XNOR U20659 ( .A(n18762), .B(n18761), .Z(n18755) );
  NAND U20660 ( .A(n18702), .B(n18701), .Z(n18706) );
  NANDN U20661 ( .A(n18704), .B(n18703), .Z(n18705) );
  NAND U20662 ( .A(n18706), .B(n18705), .Z(n18754) );
  NAND U20663 ( .A(n18708), .B(n18707), .Z(n18712) );
  NAND U20664 ( .A(n18710), .B(n18709), .Z(n18711) );
  NAND U20665 ( .A(n18712), .B(n18711), .Z(n18753) );
  XNOR U20666 ( .A(n18754), .B(n18753), .Z(n18756) );
  XNOR U20667 ( .A(n18741), .B(n18742), .Z(n18743) );
  NANDN U20668 ( .A(n18714), .B(n18713), .Z(n18718) );
  NAND U20669 ( .A(n18716), .B(n18715), .Z(n18717) );
  NAND U20670 ( .A(n18718), .B(n18717), .Z(n18749) );
  NAND U20671 ( .A(n18720), .B(n18719), .Z(n18724) );
  NAND U20672 ( .A(n18722), .B(n18721), .Z(n18723) );
  NAND U20673 ( .A(n18724), .B(n18723), .Z(n18747) );
  NAND U20674 ( .A(n18726), .B(n18725), .Z(n18730) );
  NANDN U20675 ( .A(n18728), .B(n18727), .Z(n18729) );
  AND U20676 ( .A(n18730), .B(n18729), .Z(n18748) );
  XNOR U20677 ( .A(n18747), .B(n18748), .Z(n18750) );
  XNOR U20678 ( .A(n18743), .B(n18744), .Z(n18901) );
  XOR U20679 ( .A(n18902), .B(n18901), .Z(n18907) );
  NANDN U20680 ( .A(n18732), .B(n18731), .Z(n18736) );
  NAND U20681 ( .A(n18734), .B(n18733), .Z(n18735) );
  NAND U20682 ( .A(n18736), .B(n18735), .Z(n18905) );
  XOR U20683 ( .A(n18905), .B(n18906), .Z(n18740) );
  XNOR U20684 ( .A(n18907), .B(n18740), .Z(N381) );
  NANDN U20685 ( .A(n18742), .B(n18741), .Z(n18746) );
  NANDN U20686 ( .A(n18744), .B(n18743), .Z(n18745) );
  NAND U20687 ( .A(n18746), .B(n18745), .Z(n18914) );
  NAND U20688 ( .A(n18748), .B(n18747), .Z(n18752) );
  NANDN U20689 ( .A(n18750), .B(n18749), .Z(n18751) );
  NAND U20690 ( .A(n18752), .B(n18751), .Z(n18912) );
  NAND U20691 ( .A(n18754), .B(n18753), .Z(n18758) );
  NANDN U20692 ( .A(n18756), .B(n18755), .Z(n18757) );
  NAND U20693 ( .A(n18758), .B(n18757), .Z(n18918) );
  NANDN U20694 ( .A(n18760), .B(n18759), .Z(n18764) );
  NAND U20695 ( .A(n18762), .B(n18761), .Z(n18763) );
  AND U20696 ( .A(n18764), .B(n18763), .Z(n18919) );
  XOR U20697 ( .A(n18918), .B(n18919), .Z(n18921) );
  NAND U20698 ( .A(n18766), .B(n18765), .Z(n18770) );
  NAND U20699 ( .A(n18768), .B(n18767), .Z(n18769) );
  NAND U20700 ( .A(n18770), .B(n18769), .Z(n18930) );
  NAND U20701 ( .A(n18772), .B(n18771), .Z(n18776) );
  NAND U20702 ( .A(n18774), .B(n18773), .Z(n18775) );
  AND U20703 ( .A(n18776), .B(n18775), .Z(n19041) );
  NAND U20704 ( .A(n18778), .B(n18777), .Z(n18782) );
  NAND U20705 ( .A(n18780), .B(n18779), .Z(n18781) );
  NAND U20706 ( .A(n18782), .B(n18781), .Z(n19079) );
  NAND U20707 ( .A(n18784), .B(n18783), .Z(n18788) );
  NAND U20708 ( .A(n18786), .B(n18785), .Z(n18787) );
  NAND U20709 ( .A(n18788), .B(n18787), .Z(n19078) );
  XOR U20710 ( .A(n19079), .B(n19078), .Z(n19080) );
  AND U20711 ( .A(y[7860]), .B(x[490]), .Z(n19076) );
  NAND U20712 ( .A(n18789), .B(n19076), .Z(n18793) );
  NAND U20713 ( .A(n18791), .B(n18790), .Z(n18792) );
  NAND U20714 ( .A(n18793), .B(n18792), .Z(n19047) );
  AND U20715 ( .A(x[502]), .B(y[7847]), .Z(n18992) );
  AND U20716 ( .A(x[492]), .B(y[7857]), .Z(n19134) );
  AND U20717 ( .A(x[481]), .B(y[7868]), .Z(n18990) );
  XOR U20718 ( .A(n19134), .B(n18990), .Z(n18991) );
  XOR U20719 ( .A(n18992), .B(n18991), .Z(n19046) );
  AND U20720 ( .A(x[495]), .B(y[7854]), .Z(n18995) );
  XOR U20721 ( .A(n19046), .B(n19045), .Z(n19048) );
  XNOR U20722 ( .A(n19047), .B(n19048), .Z(n19081) );
  NAND U20723 ( .A(n18795), .B(n18794), .Z(n18799) );
  NAND U20724 ( .A(n18797), .B(n18796), .Z(n18798) );
  AND U20725 ( .A(n18799), .B(n18798), .Z(n19039) );
  XNOR U20726 ( .A(n19041), .B(n19042), .Z(n19036) );
  NAND U20727 ( .A(n18801), .B(n18800), .Z(n18805) );
  NAND U20728 ( .A(n18803), .B(n18802), .Z(n18804) );
  NAND U20729 ( .A(n18805), .B(n18804), .Z(n19052) );
  AND U20730 ( .A(n18807), .B(n18806), .Z(n18811) );
  NAND U20731 ( .A(n18809), .B(n18808), .Z(n18810) );
  NANDN U20732 ( .A(n18811), .B(n18810), .Z(n19051) );
  XOR U20733 ( .A(n19052), .B(n19051), .Z(n19053) );
  NAND U20734 ( .A(n18813), .B(n18812), .Z(n18817) );
  NAND U20735 ( .A(n18815), .B(n18814), .Z(n18816) );
  NAND U20736 ( .A(n18817), .B(n18816), .Z(n18956) );
  AND U20737 ( .A(x[491]), .B(y[7858]), .Z(n19011) );
  AND U20738 ( .A(x[483]), .B(y[7866]), .Z(n19009) );
  AND U20739 ( .A(x[497]), .B(y[7852]), .Z(n19008) );
  XOR U20740 ( .A(n19009), .B(n19008), .Z(n19010) );
  XOR U20741 ( .A(n19011), .B(n19010), .Z(n18955) );
  AND U20742 ( .A(x[503]), .B(y[7846]), .Z(n19005) );
  AND U20743 ( .A(x[493]), .B(y[7856]), .Z(n19003) );
  AND U20744 ( .A(x[504]), .B(y[7845]), .Z(n19174) );
  XOR U20745 ( .A(n19003), .B(n19174), .Z(n19004) );
  XOR U20746 ( .A(n19005), .B(n19004), .Z(n18954) );
  XOR U20747 ( .A(n18955), .B(n18954), .Z(n18957) );
  XNOR U20748 ( .A(n18956), .B(n18957), .Z(n19054) );
  IV U20749 ( .A(n19054), .Z(n18818) );
  XOR U20750 ( .A(n19053), .B(n18818), .Z(n18945) );
  NAND U20751 ( .A(n19014), .B(n18819), .Z(n18823) );
  NAND U20752 ( .A(n18821), .B(n18820), .Z(n18822) );
  AND U20753 ( .A(n18823), .B(n18822), .Z(n19059) );
  AND U20754 ( .A(x[505]), .B(y[7844]), .Z(n18987) );
  AND U20755 ( .A(x[506]), .B(y[7843]), .Z(n18984) );
  XOR U20756 ( .A(n18985), .B(n18984), .Z(n18986) );
  XOR U20757 ( .A(n18987), .B(n18986), .Z(n19058) );
  AND U20758 ( .A(x[508]), .B(y[7841]), .Z(n19002) );
  XOR U20759 ( .A(o[189]), .B(n19002), .Z(n19071) );
  AND U20760 ( .A(x[480]), .B(y[7869]), .Z(n19069) );
  AND U20761 ( .A(x[509]), .B(y[7840]), .Z(n19068) );
  XOR U20762 ( .A(n19069), .B(n19068), .Z(n19070) );
  XNOR U20763 ( .A(n19071), .B(n19070), .Z(n19057) );
  XNOR U20764 ( .A(n19059), .B(n19060), .Z(n18942) );
  NAND U20765 ( .A(n18825), .B(n18824), .Z(n18829) );
  NAND U20766 ( .A(n18827), .B(n18826), .Z(n18828) );
  NAND U20767 ( .A(n18829), .B(n18828), .Z(n19023) );
  AND U20768 ( .A(o[188]), .B(n18830), .Z(n18963) );
  AND U20769 ( .A(x[496]), .B(y[7853]), .Z(n18961) );
  AND U20770 ( .A(x[507]), .B(y[7842]), .Z(n18960) );
  XOR U20771 ( .A(n18961), .B(n18960), .Z(n18962) );
  XOR U20772 ( .A(n18963), .B(n18962), .Z(n19022) );
  AND U20773 ( .A(x[482]), .B(y[7867]), .Z(n18972) );
  XOR U20774 ( .A(n18975), .B(n18974), .Z(n19021) );
  XOR U20775 ( .A(n19022), .B(n19021), .Z(n19024) );
  XOR U20776 ( .A(n19023), .B(n19024), .Z(n18943) );
  NANDN U20777 ( .A(n18832), .B(n18831), .Z(n18836) );
  NAND U20778 ( .A(n18834), .B(n18833), .Z(n18835) );
  NAND U20779 ( .A(n18836), .B(n18835), .Z(n18948) );
  NAND U20780 ( .A(n18838), .B(n18837), .Z(n18842) );
  NAND U20781 ( .A(n18840), .B(n18839), .Z(n18841) );
  NAND U20782 ( .A(n18842), .B(n18841), .Z(n18979) );
  NAND U20783 ( .A(n18844), .B(n18843), .Z(n18848) );
  NAND U20784 ( .A(n18846), .B(n18845), .Z(n18847) );
  NAND U20785 ( .A(n18848), .B(n18847), .Z(n18978) );
  XOR U20786 ( .A(n18979), .B(n18978), .Z(n18981) );
  AND U20787 ( .A(x[489]), .B(y[7860]), .Z(n19203) );
  AND U20788 ( .A(x[488]), .B(y[7861]), .Z(n19016) );
  AND U20789 ( .A(y[7863]), .B(x[486]), .Z(n18850) );
  NAND U20790 ( .A(y[7862]), .B(x[487]), .Z(n18849) );
  XNOR U20791 ( .A(n18850), .B(n18849), .Z(n19015) );
  XOR U20792 ( .A(n19016), .B(n19015), .Z(n19063) );
  XOR U20793 ( .A(n19203), .B(n19063), .Z(n19065) );
  AND U20794 ( .A(x[485]), .B(y[7864]), .Z(n18969) );
  AND U20795 ( .A(x[484]), .B(y[7865]), .Z(n18967) );
  AND U20796 ( .A(x[490]), .B(y[7859]), .Z(n18966) );
  XOR U20797 ( .A(n18967), .B(n18966), .Z(n18968) );
  XOR U20798 ( .A(n18969), .B(n18968), .Z(n19064) );
  XOR U20799 ( .A(n19065), .B(n19064), .Z(n18980) );
  XOR U20800 ( .A(n18981), .B(n18980), .Z(n18949) );
  XNOR U20801 ( .A(n18950), .B(n18951), .Z(n19034) );
  NAND U20802 ( .A(n18852), .B(n18851), .Z(n18856) );
  NAND U20803 ( .A(n18854), .B(n18853), .Z(n18855) );
  NAND U20804 ( .A(n18856), .B(n18855), .Z(n19033) );
  XOR U20805 ( .A(n18930), .B(n18931), .Z(n18933) );
  NAND U20806 ( .A(n18858), .B(n18857), .Z(n18862) );
  NAND U20807 ( .A(n18860), .B(n18859), .Z(n18861) );
  NAND U20808 ( .A(n18862), .B(n18861), .Z(n18924) );
  NANDN U20809 ( .A(n18864), .B(n18863), .Z(n18868) );
  NANDN U20810 ( .A(n18866), .B(n18865), .Z(n18867) );
  AND U20811 ( .A(n18868), .B(n18867), .Z(n18925) );
  XOR U20812 ( .A(n18924), .B(n18925), .Z(n18927) );
  NAND U20813 ( .A(n18870), .B(n18869), .Z(n18874) );
  NAND U20814 ( .A(n18872), .B(n18871), .Z(n18873) );
  NAND U20815 ( .A(n18874), .B(n18873), .Z(n18938) );
  NANDN U20816 ( .A(n18876), .B(n18875), .Z(n18880) );
  NAND U20817 ( .A(n18878), .B(n18877), .Z(n18879) );
  NAND U20818 ( .A(n18880), .B(n18879), .Z(n18936) );
  NAND U20819 ( .A(n18882), .B(n18881), .Z(n18886) );
  NAND U20820 ( .A(n18884), .B(n18883), .Z(n18885) );
  NAND U20821 ( .A(n18886), .B(n18885), .Z(n19029) );
  NAND U20822 ( .A(n18888), .B(n18887), .Z(n18892) );
  NAND U20823 ( .A(n18890), .B(n18889), .Z(n18891) );
  NAND U20824 ( .A(n18892), .B(n18891), .Z(n19028) );
  NAND U20825 ( .A(n18894), .B(n18893), .Z(n18898) );
  NAND U20826 ( .A(n18896), .B(n18895), .Z(n18897) );
  NAND U20827 ( .A(n18898), .B(n18897), .Z(n19027) );
  XOR U20828 ( .A(n19028), .B(n19027), .Z(n19030) );
  XOR U20829 ( .A(n19029), .B(n19030), .Z(n18937) );
  XOR U20830 ( .A(n18936), .B(n18937), .Z(n18939) );
  XOR U20831 ( .A(n18938), .B(n18939), .Z(n18926) );
  XOR U20832 ( .A(n18927), .B(n18926), .Z(n18932) );
  XOR U20833 ( .A(n18933), .B(n18932), .Z(n18920) );
  XOR U20834 ( .A(n18921), .B(n18920), .Z(n18913) );
  XNOR U20835 ( .A(n18912), .B(n18913), .Z(n18915) );
  XOR U20836 ( .A(n18914), .B(n18915), .Z(n18911) );
  NAND U20837 ( .A(n18900), .B(n18899), .Z(n18904) );
  NAND U20838 ( .A(n18902), .B(n18901), .Z(n18903) );
  NAND U20839 ( .A(n18904), .B(n18903), .Z(n18910) );
  XOR U20840 ( .A(n18910), .B(n18909), .Z(n18908) );
  XNOR U20841 ( .A(n18911), .B(n18908), .Z(N382) );
  NAND U20842 ( .A(n18913), .B(n18912), .Z(n18917) );
  NANDN U20843 ( .A(n18915), .B(n18914), .Z(n18916) );
  NAND U20844 ( .A(n18917), .B(n18916), .Z(n19087) );
  NAND U20845 ( .A(n18919), .B(n18918), .Z(n18923) );
  NAND U20846 ( .A(n18921), .B(n18920), .Z(n18922) );
  NAND U20847 ( .A(n18923), .B(n18922), .Z(n19370) );
  NAND U20848 ( .A(n18925), .B(n18924), .Z(n18929) );
  NAND U20849 ( .A(n18927), .B(n18926), .Z(n18928) );
  AND U20850 ( .A(n18929), .B(n18928), .Z(n19377) );
  NAND U20851 ( .A(n18931), .B(n18930), .Z(n18935) );
  NAND U20852 ( .A(n18933), .B(n18932), .Z(n18934) );
  AND U20853 ( .A(n18935), .B(n18934), .Z(n19376) );
  XOR U20854 ( .A(n19377), .B(n19376), .Z(n19379) );
  NAND U20855 ( .A(n18937), .B(n18936), .Z(n18941) );
  NAND U20856 ( .A(n18939), .B(n18938), .Z(n18940) );
  AND U20857 ( .A(n18941), .B(n18940), .Z(n19378) );
  XOR U20858 ( .A(n19379), .B(n19378), .Z(n19372) );
  NANDN U20859 ( .A(n18943), .B(n18942), .Z(n18947) );
  NANDN U20860 ( .A(n18945), .B(n18944), .Z(n18946) );
  AND U20861 ( .A(n18947), .B(n18946), .Z(n19358) );
  NANDN U20862 ( .A(n18949), .B(n18948), .Z(n18953) );
  NANDN U20863 ( .A(n18951), .B(n18950), .Z(n18952) );
  AND U20864 ( .A(n18953), .B(n18952), .Z(n19350) );
  NAND U20865 ( .A(n18955), .B(n18954), .Z(n18959) );
  NAND U20866 ( .A(n18957), .B(n18956), .Z(n18958) );
  AND U20867 ( .A(n18959), .B(n18958), .Z(n19334) );
  NAND U20868 ( .A(n18961), .B(n18960), .Z(n18965) );
  NAND U20869 ( .A(n18963), .B(n18962), .Z(n18964) );
  NAND U20870 ( .A(n18965), .B(n18964), .Z(n19292) );
  NAND U20871 ( .A(n18967), .B(n18966), .Z(n18971) );
  NAND U20872 ( .A(n18969), .B(n18968), .Z(n18970) );
  NAND U20873 ( .A(n18971), .B(n18970), .Z(n19295) );
  AND U20874 ( .A(x[486]), .B(y[7864]), .Z(n19153) );
  AND U20875 ( .A(x[485]), .B(y[7865]), .Z(n19155) );
  AND U20876 ( .A(x[499]), .B(y[7851]), .Z(n19154) );
  XOR U20877 ( .A(n19155), .B(n19154), .Z(n19152) );
  XNOR U20878 ( .A(n19153), .B(n19152), .Z(n19102) );
  AND U20879 ( .A(x[484]), .B(y[7866]), .Z(n19147) );
  AND U20880 ( .A(x[483]), .B(y[7867]), .Z(n19149) );
  AND U20881 ( .A(x[498]), .B(y[7852]), .Z(n19148) );
  XOR U20882 ( .A(n19149), .B(n19148), .Z(n19146) );
  XOR U20883 ( .A(n19147), .B(n19146), .Z(n19105) );
  NANDN U20884 ( .A(n18973), .B(n18972), .Z(n18977) );
  NAND U20885 ( .A(n18975), .B(n18974), .Z(n18976) );
  AND U20886 ( .A(n18977), .B(n18976), .Z(n19104) );
  XOR U20887 ( .A(n19102), .B(n19103), .Z(n19294) );
  XOR U20888 ( .A(n19295), .B(n19294), .Z(n19293) );
  XOR U20889 ( .A(n19292), .B(n19293), .Z(n19335) );
  NAND U20890 ( .A(n18979), .B(n18978), .Z(n18983) );
  NAND U20891 ( .A(n18981), .B(n18980), .Z(n18982) );
  AND U20892 ( .A(n18983), .B(n18982), .Z(n19332) );
  XOR U20893 ( .A(n19333), .B(n19332), .Z(n19353) );
  AND U20894 ( .A(n18985), .B(n18984), .Z(n18989) );
  NAND U20895 ( .A(n18987), .B(n18986), .Z(n18988) );
  NANDN U20896 ( .A(n18989), .B(n18988), .Z(n19286) );
  AND U20897 ( .A(n19134), .B(n18990), .Z(n18994) );
  NAND U20898 ( .A(n18992), .B(n18991), .Z(n18993) );
  NANDN U20899 ( .A(n18994), .B(n18993), .Z(n19289) );
  NANDN U20900 ( .A(n19139), .B(n18995), .Z(n18999) );
  NANDN U20901 ( .A(n18997), .B(n18996), .Z(n18998) );
  AND U20902 ( .A(n18999), .B(n18998), .Z(n19123) );
  AND U20903 ( .A(x[503]), .B(y[7847]), .Z(n19173) );
  AND U20904 ( .A(y[7846]), .B(x[504]), .Z(n19001) );
  AND U20905 ( .A(y[7845]), .B(x[505]), .Z(n19000) );
  XOR U20906 ( .A(n19001), .B(n19000), .Z(n19172) );
  XOR U20907 ( .A(n19173), .B(n19172), .Z(n19125) );
  AND U20908 ( .A(n19002), .B(o[189]), .Z(n19213) );
  AND U20909 ( .A(x[508]), .B(y[7842]), .Z(n19215) );
  AND U20910 ( .A(x[496]), .B(y[7854]), .Z(n19214) );
  XOR U20911 ( .A(n19215), .B(n19214), .Z(n19212) );
  XNOR U20912 ( .A(n19213), .B(n19212), .Z(n19124) );
  XNOR U20913 ( .A(n19123), .B(n19122), .Z(n19288) );
  XOR U20914 ( .A(n19289), .B(n19288), .Z(n19287) );
  XOR U20915 ( .A(n19286), .B(n19287), .Z(n19091) );
  NAND U20916 ( .A(n19003), .B(n19174), .Z(n19007) );
  NAND U20917 ( .A(n19005), .B(n19004), .Z(n19006) );
  NAND U20918 ( .A(n19007), .B(n19006), .Z(n19317) );
  NAND U20919 ( .A(n19009), .B(n19008), .Z(n19013) );
  NAND U20920 ( .A(n19011), .B(n19010), .Z(n19012) );
  AND U20921 ( .A(n19013), .B(n19012), .Z(n19129) );
  AND U20922 ( .A(x[480]), .B(y[7870]), .Z(n19221) );
  AND U20923 ( .A(x[509]), .B(y[7841]), .Z(n19226) );
  XOR U20924 ( .A(o[190]), .B(n19226), .Z(n19223) );
  AND U20925 ( .A(x[510]), .B(y[7840]), .Z(n19222) );
  XOR U20926 ( .A(n19223), .B(n19222), .Z(n19220) );
  XOR U20927 ( .A(n19221), .B(n19220), .Z(n19131) );
  AND U20928 ( .A(x[500]), .B(y[7850]), .Z(n19208) );
  AND U20929 ( .A(x[488]), .B(y[7862]), .Z(n19206) );
  XNOR U20930 ( .A(n19207), .B(n19206), .Z(n19130) );
  XNOR U20931 ( .A(n19129), .B(n19128), .Z(n19316) );
  XOR U20932 ( .A(n19317), .B(n19316), .Z(n19314) );
  AND U20933 ( .A(x[487]), .B(y[7863]), .Z(n19141) );
  NAND U20934 ( .A(n19014), .B(n19141), .Z(n19018) );
  NAND U20935 ( .A(n19016), .B(n19015), .Z(n19017) );
  AND U20936 ( .A(n19018), .B(n19017), .Z(n19114) );
  AND U20937 ( .A(y[7849]), .B(x[501]), .Z(n19020) );
  AND U20938 ( .A(y[7848]), .B(x[502]), .Z(n19019) );
  XOR U20939 ( .A(n19020), .B(n19019), .Z(n19140) );
  XOR U20940 ( .A(n19141), .B(n19140), .Z(n19117) );
  AND U20941 ( .A(x[497]), .B(y[7853]), .Z(n19167) );
  AND U20942 ( .A(x[482]), .B(y[7868]), .Z(n19169) );
  AND U20943 ( .A(x[506]), .B(y[7844]), .Z(n19168) );
  XOR U20944 ( .A(n19169), .B(n19168), .Z(n19166) );
  XNOR U20945 ( .A(n19167), .B(n19166), .Z(n19116) );
  XNOR U20946 ( .A(n19114), .B(n19115), .Z(n19315) );
  NAND U20947 ( .A(n19022), .B(n19021), .Z(n19026) );
  NAND U20948 ( .A(n19024), .B(n19023), .Z(n19025) );
  NAND U20949 ( .A(n19026), .B(n19025), .Z(n19092) );
  XOR U20950 ( .A(n19093), .B(n19092), .Z(n19090) );
  XOR U20951 ( .A(n19091), .B(n19090), .Z(n19352) );
  XNOR U20952 ( .A(n19350), .B(n19351), .Z(n19360) );
  NAND U20953 ( .A(n19028), .B(n19027), .Z(n19032) );
  NAND U20954 ( .A(n19030), .B(n19029), .Z(n19031) );
  AND U20955 ( .A(n19032), .B(n19031), .Z(n19359) );
  NANDN U20956 ( .A(n19034), .B(n19033), .Z(n19038) );
  NANDN U20957 ( .A(n19036), .B(n19035), .Z(n19037) );
  NAND U20958 ( .A(n19038), .B(n19037), .Z(n19346) );
  NANDN U20959 ( .A(n19040), .B(n19039), .Z(n19044) );
  NANDN U20960 ( .A(n19042), .B(n19041), .Z(n19043) );
  AND U20961 ( .A(n19044), .B(n19043), .Z(n19326) );
  NAND U20962 ( .A(n19046), .B(n19045), .Z(n19050) );
  NAND U20963 ( .A(n19048), .B(n19047), .Z(n19049) );
  AND U20964 ( .A(n19050), .B(n19049), .Z(n19311) );
  NAND U20965 ( .A(n19052), .B(n19051), .Z(n19056) );
  NANDN U20966 ( .A(n19054), .B(n19053), .Z(n19055) );
  AND U20967 ( .A(n19056), .B(n19055), .Z(n19310) );
  XOR U20968 ( .A(n19311), .B(n19310), .Z(n19309) );
  NANDN U20969 ( .A(n19058), .B(n19057), .Z(n19062) );
  NANDN U20970 ( .A(n19060), .B(n19059), .Z(n19061) );
  NAND U20971 ( .A(n19062), .B(n19061), .Z(n19308) );
  XOR U20972 ( .A(n19309), .B(n19308), .Z(n19329) );
  NAND U20973 ( .A(n19203), .B(n19063), .Z(n19067) );
  NAND U20974 ( .A(n19065), .B(n19064), .Z(n19066) );
  AND U20975 ( .A(n19067), .B(n19066), .Z(n19098) );
  NAND U20976 ( .A(n19069), .B(n19068), .Z(n19073) );
  NAND U20977 ( .A(n19071), .B(n19070), .Z(n19072) );
  NAND U20978 ( .A(n19073), .B(n19072), .Z(n19108) );
  NAND U20979 ( .A(y[7858]), .B(x[492]), .Z(n19074) );
  XNOR U20980 ( .A(n19075), .B(n19074), .Z(n19136) );
  AND U20981 ( .A(y[7861]), .B(x[489]), .Z(n19077) );
  XOR U20982 ( .A(n19077), .B(n19076), .Z(n19201) );
  XOR U20983 ( .A(n19202), .B(n19201), .Z(n19111) );
  AND U20984 ( .A(x[507]), .B(y[7843]), .Z(n19163) );
  AND U20985 ( .A(x[481]), .B(y[7869]), .Z(n19162) );
  XOR U20986 ( .A(n19163), .B(n19162), .Z(n19161) );
  XOR U20987 ( .A(n19161), .B(n19160), .Z(n19110) );
  XOR U20988 ( .A(n19111), .B(n19110), .Z(n19109) );
  XOR U20989 ( .A(n19108), .B(n19109), .Z(n19099) );
  NAND U20990 ( .A(n19079), .B(n19078), .Z(n19083) );
  NANDN U20991 ( .A(n19081), .B(n19080), .Z(n19082) );
  AND U20992 ( .A(n19083), .B(n19082), .Z(n19096) );
  XNOR U20993 ( .A(n19097), .B(n19096), .Z(n19328) );
  XNOR U20994 ( .A(n19326), .B(n19327), .Z(n19347) );
  XOR U20995 ( .A(n19346), .B(n19347), .Z(n19344) );
  XOR U20996 ( .A(n19345), .B(n19344), .Z(n19373) );
  XOR U20997 ( .A(n19370), .B(n19371), .Z(n19084) );
  XNOR U20998 ( .A(n19085), .B(n19084), .Z(N383) );
  NAND U20999 ( .A(n19085), .B(n19084), .Z(n19089) );
  NANDN U21000 ( .A(n19087), .B(n19086), .Z(n19088) );
  AND U21001 ( .A(n19089), .B(n19088), .Z(n19369) );
  NAND U21002 ( .A(n19091), .B(n19090), .Z(n19095) );
  NAND U21003 ( .A(n19093), .B(n19092), .Z(n19094) );
  AND U21004 ( .A(n19095), .B(n19094), .Z(n19343) );
  NAND U21005 ( .A(n19097), .B(n19096), .Z(n19101) );
  NANDN U21006 ( .A(n19099), .B(n19098), .Z(n19100) );
  AND U21007 ( .A(n19101), .B(n19100), .Z(n19325) );
  NANDN U21008 ( .A(n19103), .B(n19102), .Z(n19107) );
  NANDN U21009 ( .A(n19105), .B(n19104), .Z(n19106) );
  AND U21010 ( .A(n19107), .B(n19106), .Z(n19307) );
  NAND U21011 ( .A(n19109), .B(n19108), .Z(n19113) );
  NAND U21012 ( .A(n19111), .B(n19110), .Z(n19112) );
  AND U21013 ( .A(n19113), .B(n19112), .Z(n19121) );
  NANDN U21014 ( .A(n19115), .B(n19114), .Z(n19119) );
  NANDN U21015 ( .A(n19117), .B(n19116), .Z(n19118) );
  NAND U21016 ( .A(n19119), .B(n19118), .Z(n19120) );
  XNOR U21017 ( .A(n19121), .B(n19120), .Z(n19305) );
  NAND U21018 ( .A(n19123), .B(n19122), .Z(n19127) );
  NANDN U21019 ( .A(n19125), .B(n19124), .Z(n19126) );
  AND U21020 ( .A(n19127), .B(n19126), .Z(n19303) );
  NAND U21021 ( .A(n19129), .B(n19128), .Z(n19133) );
  NANDN U21022 ( .A(n19131), .B(n19130), .Z(n19132) );
  AND U21023 ( .A(n19133), .B(n19132), .Z(n19285) );
  AND U21024 ( .A(n19134), .B(n19251), .Z(n19138) );
  ANDN U21025 ( .B(n19136), .A(n19135), .Z(n19137) );
  NOR U21026 ( .A(n19138), .B(n19137), .Z(n19145) );
  AND U21027 ( .A(x[502]), .B(y[7849]), .Z(n19227) );
  NANDN U21028 ( .A(n19139), .B(n19227), .Z(n19143) );
  NAND U21029 ( .A(n19141), .B(n19140), .Z(n19142) );
  AND U21030 ( .A(n19143), .B(n19142), .Z(n19144) );
  XNOR U21031 ( .A(n19145), .B(n19144), .Z(n19200) );
  NAND U21032 ( .A(n19147), .B(n19146), .Z(n19151) );
  NAND U21033 ( .A(n19149), .B(n19148), .Z(n19150) );
  AND U21034 ( .A(n19151), .B(n19150), .Z(n19159) );
  NAND U21035 ( .A(n19153), .B(n19152), .Z(n19157) );
  NAND U21036 ( .A(n19155), .B(n19154), .Z(n19156) );
  NAND U21037 ( .A(n19157), .B(n19156), .Z(n19158) );
  XNOR U21038 ( .A(n19159), .B(n19158), .Z(n19198) );
  NAND U21039 ( .A(n19161), .B(n19160), .Z(n19165) );
  NAND U21040 ( .A(n19163), .B(n19162), .Z(n19164) );
  AND U21041 ( .A(n19165), .B(n19164), .Z(n19196) );
  NAND U21042 ( .A(n19167), .B(n19166), .Z(n19171) );
  NAND U21043 ( .A(n19169), .B(n19168), .Z(n19170) );
  AND U21044 ( .A(n19171), .B(n19170), .Z(n19178) );
  NAND U21045 ( .A(n19173), .B(n19172), .Z(n19176) );
  AND U21046 ( .A(x[505]), .B(y[7846]), .Z(n19228) );
  NAND U21047 ( .A(n19174), .B(n19228), .Z(n19175) );
  NAND U21048 ( .A(n19176), .B(n19175), .Z(n19177) );
  XNOR U21049 ( .A(n19178), .B(n19177), .Z(n19194) );
  AND U21050 ( .A(y[7844]), .B(x[507]), .Z(n19180) );
  NAND U21051 ( .A(y[7848]), .B(x[503]), .Z(n19179) );
  XNOR U21052 ( .A(n19180), .B(n19179), .Z(n19184) );
  AND U21053 ( .A(y[7869]), .B(x[482]), .Z(n19182) );
  NAND U21054 ( .A(y[7854]), .B(x[497]), .Z(n19181) );
  XNOR U21055 ( .A(n19182), .B(n19181), .Z(n19183) );
  XOR U21056 ( .A(n19184), .B(n19183), .Z(n19192) );
  AND U21057 ( .A(y[7865]), .B(x[486]), .Z(n19186) );
  NAND U21058 ( .A(y[7864]), .B(x[487]), .Z(n19185) );
  XNOR U21059 ( .A(n19186), .B(n19185), .Z(n19190) );
  AND U21060 ( .A(y[7866]), .B(x[485]), .Z(n19188) );
  NAND U21061 ( .A(y[7867]), .B(x[484]), .Z(n19187) );
  XNOR U21062 ( .A(n19188), .B(n19187), .Z(n19189) );
  XNOR U21063 ( .A(n19190), .B(n19189), .Z(n19191) );
  XNOR U21064 ( .A(n19192), .B(n19191), .Z(n19193) );
  XNOR U21065 ( .A(n19194), .B(n19193), .Z(n19195) );
  XNOR U21066 ( .A(n19196), .B(n19195), .Z(n19197) );
  XOR U21067 ( .A(n19198), .B(n19197), .Z(n19199) );
  XNOR U21068 ( .A(n19200), .B(n19199), .Z(n19283) );
  NAND U21069 ( .A(n19202), .B(n19201), .Z(n19205) );
  AND U21070 ( .A(x[490]), .B(y[7861]), .Z(n19250) );
  NAND U21071 ( .A(n19203), .B(n19250), .Z(n19204) );
  AND U21072 ( .A(n19205), .B(n19204), .Z(n19281) );
  NAND U21073 ( .A(n19207), .B(n19206), .Z(n19211) );
  NANDN U21074 ( .A(n19209), .B(n19208), .Z(n19210) );
  AND U21075 ( .A(n19211), .B(n19210), .Z(n19219) );
  NAND U21076 ( .A(n19213), .B(n19212), .Z(n19217) );
  NAND U21077 ( .A(n19215), .B(n19214), .Z(n19216) );
  NAND U21078 ( .A(n19217), .B(n19216), .Z(n19218) );
  XNOR U21079 ( .A(n19219), .B(n19218), .Z(n19279) );
  NAND U21080 ( .A(n19221), .B(n19220), .Z(n19225) );
  NAND U21081 ( .A(n19223), .B(n19222), .Z(n19224) );
  AND U21082 ( .A(n19225), .B(n19224), .Z(n19277) );
  AND U21083 ( .A(y[7850]), .B(x[501]), .Z(n19235) );
  AND U21084 ( .A(n19226), .B(o[190]), .Z(n19233) );
  XOR U21085 ( .A(n19227), .B(o[191]), .Z(n19231) );
  XNOR U21086 ( .A(n19229), .B(n19228), .Z(n19230) );
  XNOR U21087 ( .A(n19231), .B(n19230), .Z(n19232) );
  XNOR U21088 ( .A(n19233), .B(n19232), .Z(n19234) );
  XNOR U21089 ( .A(n19235), .B(n19234), .Z(n19275) );
  AND U21090 ( .A(y[7857]), .B(x[494]), .Z(n19241) );
  AND U21091 ( .A(y[7870]), .B(x[481]), .Z(n19237) );
  NAND U21092 ( .A(y[7843]), .B(x[508]), .Z(n19236) );
  XNOR U21093 ( .A(n19237), .B(n19236), .Z(n19238) );
  XNOR U21094 ( .A(n19239), .B(n19238), .Z(n19240) );
  XNOR U21095 ( .A(n19241), .B(n19240), .Z(n19265) );
  AND U21096 ( .A(y[7842]), .B(x[509]), .Z(n19243) );
  NAND U21097 ( .A(y[7863]), .B(x[488]), .Z(n19242) );
  XNOR U21098 ( .A(n19243), .B(n19242), .Z(n19255) );
  AND U21099 ( .A(y[7841]), .B(x[510]), .Z(n19245) );
  NAND U21100 ( .A(y[7855]), .B(x[496]), .Z(n19244) );
  XNOR U21101 ( .A(n19245), .B(n19244), .Z(n19249) );
  AND U21102 ( .A(y[7860]), .B(x[491]), .Z(n19247) );
  NAND U21103 ( .A(y[7851]), .B(x[500]), .Z(n19246) );
  XNOR U21104 ( .A(n19247), .B(n19246), .Z(n19248) );
  XOR U21105 ( .A(n19249), .B(n19248), .Z(n19253) );
  XNOR U21106 ( .A(n19251), .B(n19250), .Z(n19252) );
  XNOR U21107 ( .A(n19253), .B(n19252), .Z(n19254) );
  XOR U21108 ( .A(n19255), .B(n19254), .Z(n19263) );
  AND U21109 ( .A(y[7852]), .B(x[499]), .Z(n19257) );
  NAND U21110 ( .A(y[7868]), .B(x[483]), .Z(n19256) );
  XNOR U21111 ( .A(n19257), .B(n19256), .Z(n19261) );
  AND U21112 ( .A(y[7840]), .B(x[511]), .Z(n19259) );
  NAND U21113 ( .A(y[7853]), .B(x[498]), .Z(n19258) );
  XNOR U21114 ( .A(n19259), .B(n19258), .Z(n19260) );
  XNOR U21115 ( .A(n19261), .B(n19260), .Z(n19262) );
  XNOR U21116 ( .A(n19263), .B(n19262), .Z(n19264) );
  XOR U21117 ( .A(n19265), .B(n19264), .Z(n19273) );
  AND U21118 ( .A(y[7859]), .B(x[492]), .Z(n19267) );
  NAND U21119 ( .A(y[7845]), .B(x[506]), .Z(n19266) );
  XNOR U21120 ( .A(n19267), .B(n19266), .Z(n19271) );
  AND U21121 ( .A(y[7862]), .B(x[489]), .Z(n19269) );
  NAND U21122 ( .A(y[7871]), .B(x[480]), .Z(n19268) );
  XNOR U21123 ( .A(n19269), .B(n19268), .Z(n19270) );
  XNOR U21124 ( .A(n19271), .B(n19270), .Z(n19272) );
  XNOR U21125 ( .A(n19273), .B(n19272), .Z(n19274) );
  XNOR U21126 ( .A(n19275), .B(n19274), .Z(n19276) );
  XNOR U21127 ( .A(n19277), .B(n19276), .Z(n19278) );
  XNOR U21128 ( .A(n19279), .B(n19278), .Z(n19280) );
  XNOR U21129 ( .A(n19281), .B(n19280), .Z(n19282) );
  XNOR U21130 ( .A(n19283), .B(n19282), .Z(n19284) );
  XNOR U21131 ( .A(n19285), .B(n19284), .Z(n19301) );
  NAND U21132 ( .A(n19287), .B(n19286), .Z(n19291) );
  NAND U21133 ( .A(n19289), .B(n19288), .Z(n19290) );
  AND U21134 ( .A(n19291), .B(n19290), .Z(n19299) );
  NAND U21135 ( .A(n19293), .B(n19292), .Z(n19297) );
  NAND U21136 ( .A(n19295), .B(n19294), .Z(n19296) );
  NAND U21137 ( .A(n19297), .B(n19296), .Z(n19298) );
  XNOR U21138 ( .A(n19299), .B(n19298), .Z(n19300) );
  XNOR U21139 ( .A(n19301), .B(n19300), .Z(n19302) );
  XNOR U21140 ( .A(n19303), .B(n19302), .Z(n19304) );
  XNOR U21141 ( .A(n19305), .B(n19304), .Z(n19306) );
  XNOR U21142 ( .A(n19307), .B(n19306), .Z(n19323) );
  NAND U21143 ( .A(n19309), .B(n19308), .Z(n19313) );
  NAND U21144 ( .A(n19311), .B(n19310), .Z(n19312) );
  AND U21145 ( .A(n19313), .B(n19312), .Z(n19321) );
  NANDN U21146 ( .A(n19315), .B(n19314), .Z(n19319) );
  NAND U21147 ( .A(n19317), .B(n19316), .Z(n19318) );
  NAND U21148 ( .A(n19319), .B(n19318), .Z(n19320) );
  XNOR U21149 ( .A(n19321), .B(n19320), .Z(n19322) );
  XNOR U21150 ( .A(n19323), .B(n19322), .Z(n19324) );
  XNOR U21151 ( .A(n19325), .B(n19324), .Z(n19341) );
  NANDN U21152 ( .A(n19327), .B(n19326), .Z(n19331) );
  NANDN U21153 ( .A(n19329), .B(n19328), .Z(n19330) );
  AND U21154 ( .A(n19331), .B(n19330), .Z(n19339) );
  NAND U21155 ( .A(n19333), .B(n19332), .Z(n19337) );
  NANDN U21156 ( .A(n19335), .B(n19334), .Z(n19336) );
  NAND U21157 ( .A(n19337), .B(n19336), .Z(n19338) );
  XNOR U21158 ( .A(n19339), .B(n19338), .Z(n19340) );
  XNOR U21159 ( .A(n19341), .B(n19340), .Z(n19342) );
  XNOR U21160 ( .A(n19343), .B(n19342), .Z(n19367) );
  NAND U21161 ( .A(n19345), .B(n19344), .Z(n19349) );
  NAND U21162 ( .A(n19347), .B(n19346), .Z(n19348) );
  AND U21163 ( .A(n19349), .B(n19348), .Z(n19357) );
  NANDN U21164 ( .A(n19351), .B(n19350), .Z(n19355) );
  NANDN U21165 ( .A(n19353), .B(n19352), .Z(n19354) );
  NAND U21166 ( .A(n19355), .B(n19354), .Z(n19356) );
  XNOR U21167 ( .A(n19357), .B(n19356), .Z(n19365) );
  ANDN U21168 ( .B(n19359), .A(n19358), .Z(n19361) );
  NANDN U21169 ( .A(n19361), .B(n19360), .Z(n19362) );
  NAND U21170 ( .A(n19363), .B(n19362), .Z(n19364) );
  XNOR U21171 ( .A(n19365), .B(n19364), .Z(n19366) );
  XNOR U21172 ( .A(n19367), .B(n19366), .Z(n19368) );
  XNOR U21173 ( .A(n19369), .B(n19368), .Z(n19385) );
  NANDN U21174 ( .A(n19371), .B(n19370), .Z(n19375) );
  ANDN U21175 ( .B(n19373), .A(n19372), .Z(n19374) );
  ANDN U21176 ( .B(n19375), .A(n19374), .Z(n19383) );
  AND U21177 ( .A(n19377), .B(n19376), .Z(n19381) );
  AND U21178 ( .A(n19379), .B(n19378), .Z(n19380) );
  OR U21179 ( .A(n19381), .B(n19380), .Z(n19382) );
  XNOR U21180 ( .A(n19383), .B(n19382), .Z(n19384) );
  XNOR U21181 ( .A(n19385), .B(n19384), .Z(N384) );
  AND U21182 ( .A(x[480]), .B(y[7872]), .Z(n19997) );
  XOR U21183 ( .A(n19997), .B(o[192]), .Z(N417) );
  AND U21184 ( .A(x[481]), .B(y[7872]), .Z(n19394) );
  AND U21185 ( .A(x[480]), .B(y[7873]), .Z(n19393) );
  XNOR U21186 ( .A(n19393), .B(o[193]), .Z(n19386) );
  XNOR U21187 ( .A(n19394), .B(n19386), .Z(n19388) );
  NAND U21188 ( .A(n19997), .B(o[192]), .Z(n19387) );
  XNOR U21189 ( .A(n19388), .B(n19387), .Z(N418) );
  NANDN U21190 ( .A(n19394), .B(n19386), .Z(n19390) );
  NAND U21191 ( .A(n19388), .B(n19387), .Z(n19389) );
  AND U21192 ( .A(n19390), .B(n19389), .Z(n19400) );
  AND U21193 ( .A(x[480]), .B(y[7874]), .Z(n19405) );
  XNOR U21194 ( .A(n19405), .B(o[194]), .Z(n19399) );
  XNOR U21195 ( .A(n19400), .B(n19399), .Z(n19402) );
  AND U21196 ( .A(y[7872]), .B(x[482]), .Z(n19392) );
  NAND U21197 ( .A(y[7873]), .B(x[481]), .Z(n19391) );
  XNOR U21198 ( .A(n19392), .B(n19391), .Z(n19396) );
  AND U21199 ( .A(n19393), .B(o[193]), .Z(n19395) );
  XNOR U21200 ( .A(n19396), .B(n19395), .Z(n19401) );
  XNOR U21201 ( .A(n19402), .B(n19401), .Z(N419) );
  AND U21202 ( .A(x[482]), .B(y[7873]), .Z(n19412) );
  NAND U21203 ( .A(n19412), .B(n19394), .Z(n19398) );
  NAND U21204 ( .A(n19396), .B(n19395), .Z(n19397) );
  AND U21205 ( .A(n19398), .B(n19397), .Z(n19417) );
  NANDN U21206 ( .A(n19400), .B(n19399), .Z(n19404) );
  NAND U21207 ( .A(n19402), .B(n19401), .Z(n19403) );
  AND U21208 ( .A(n19404), .B(n19403), .Z(n19416) );
  XNOR U21209 ( .A(n19417), .B(n19416), .Z(n19419) );
  AND U21210 ( .A(x[481]), .B(y[7874]), .Z(n19519) );
  XOR U21211 ( .A(n19412), .B(o[195]), .Z(n19422) );
  XOR U21212 ( .A(n19519), .B(n19422), .Z(n19424) );
  AND U21213 ( .A(n19405), .B(o[194]), .Z(n19409) );
  AND U21214 ( .A(y[7872]), .B(x[483]), .Z(n19407) );
  NAND U21215 ( .A(y[7875]), .B(x[480]), .Z(n19406) );
  XNOR U21216 ( .A(n19407), .B(n19406), .Z(n19408) );
  XOR U21217 ( .A(n19409), .B(n19408), .Z(n19423) );
  XOR U21218 ( .A(n19424), .B(n19423), .Z(n19418) );
  XOR U21219 ( .A(n19419), .B(n19418), .Z(N420) );
  AND U21220 ( .A(y[7875]), .B(x[483]), .Z(n19476) );
  NAND U21221 ( .A(n19997), .B(n19476), .Z(n19411) );
  NAND U21222 ( .A(n19409), .B(n19408), .Z(n19410) );
  NAND U21223 ( .A(n19411), .B(n19410), .Z(n19430) );
  AND U21224 ( .A(n19412), .B(o[195]), .Z(n19449) );
  AND U21225 ( .A(y[7876]), .B(x[480]), .Z(n19414) );
  AND U21226 ( .A(y[7872]), .B(x[484]), .Z(n19413) );
  XOR U21227 ( .A(n19414), .B(n19413), .Z(n19448) );
  XOR U21228 ( .A(n19449), .B(n19448), .Z(n19429) );
  AND U21229 ( .A(y[7874]), .B(x[482]), .Z(n19573) );
  NAND U21230 ( .A(y[7875]), .B(x[481]), .Z(n19415) );
  XNOR U21231 ( .A(n19573), .B(n19415), .Z(n19445) );
  NAND U21232 ( .A(x[483]), .B(y[7873]), .Z(n19442) );
  XOR U21233 ( .A(n19445), .B(n19444), .Z(n19428) );
  XOR U21234 ( .A(n19429), .B(n19428), .Z(n19431) );
  XOR U21235 ( .A(n19430), .B(n19431), .Z(n19435) );
  NANDN U21236 ( .A(n19417), .B(n19416), .Z(n19421) );
  NAND U21237 ( .A(n19419), .B(n19418), .Z(n19420) );
  NAND U21238 ( .A(n19421), .B(n19420), .Z(n19436) );
  NAND U21239 ( .A(n19519), .B(n19422), .Z(n19426) );
  NAND U21240 ( .A(n19424), .B(n19423), .Z(n19425) );
  NAND U21241 ( .A(n19426), .B(n19425), .Z(n19437) );
  IV U21242 ( .A(n19437), .Z(n19434) );
  XOR U21243 ( .A(n19436), .B(n19434), .Z(n19427) );
  XNOR U21244 ( .A(n19435), .B(n19427), .Z(N421) );
  NAND U21245 ( .A(n19429), .B(n19428), .Z(n19433) );
  NAND U21246 ( .A(n19431), .B(n19430), .Z(n19432) );
  AND U21247 ( .A(n19433), .B(n19432), .Z(n19459) );
  AND U21248 ( .A(y[7874]), .B(x[483]), .Z(n19439) );
  NAND U21249 ( .A(y[7876]), .B(x[481]), .Z(n19438) );
  XNOR U21250 ( .A(n19439), .B(n19438), .Z(n19463) );
  AND U21251 ( .A(x[484]), .B(y[7873]), .Z(n19474) );
  XOR U21252 ( .A(n19474), .B(o[197]), .Z(n19462) );
  XNOR U21253 ( .A(n19463), .B(n19462), .Z(n19466) );
  NAND U21254 ( .A(x[482]), .B(y[7875]), .Z(n19528) );
  AND U21255 ( .A(y[7872]), .B(x[485]), .Z(n19441) );
  NAND U21256 ( .A(y[7877]), .B(x[480]), .Z(n19440) );
  XNOR U21257 ( .A(n19441), .B(n19440), .Z(n19469) );
  ANDN U21258 ( .B(o[196]), .A(n19442), .Z(n19468) );
  XOR U21259 ( .A(n19469), .B(n19468), .Z(n19467) );
  XOR U21260 ( .A(n19528), .B(n19467), .Z(n19443) );
  XOR U21261 ( .A(n19466), .B(n19443), .Z(n19455) );
  NANDN U21262 ( .A(n19528), .B(n19519), .Z(n19447) );
  NAND U21263 ( .A(n19445), .B(n19444), .Z(n19446) );
  NAND U21264 ( .A(n19447), .B(n19446), .Z(n19454) );
  AND U21265 ( .A(x[484]), .B(y[7876]), .Z(n20201) );
  NAND U21266 ( .A(n20201), .B(n19997), .Z(n19451) );
  NAND U21267 ( .A(n19449), .B(n19448), .Z(n19450) );
  NAND U21268 ( .A(n19451), .B(n19450), .Z(n19453) );
  XNOR U21269 ( .A(n19454), .B(n19453), .Z(n19456) );
  XNOR U21270 ( .A(n19460), .B(n19461), .Z(n19452) );
  XOR U21271 ( .A(n19459), .B(n19452), .Z(N422) );
  NAND U21272 ( .A(n19454), .B(n19453), .Z(n19458) );
  NANDN U21273 ( .A(n19456), .B(n19455), .Z(n19457) );
  AND U21274 ( .A(n19458), .B(n19457), .Z(n19503) );
  AND U21275 ( .A(x[483]), .B(y[7876]), .Z(n19529) );
  NAND U21276 ( .A(n19529), .B(n19519), .Z(n19465) );
  NAND U21277 ( .A(n19463), .B(n19462), .Z(n19464) );
  NAND U21278 ( .A(n19465), .B(n19464), .Z(n19506) );
  XOR U21279 ( .A(n19506), .B(n19507), .Z(n19509) );
  AND U21280 ( .A(x[485]), .B(y[7877]), .Z(n19702) );
  NAND U21281 ( .A(n19997), .B(n19702), .Z(n19471) );
  NAND U21282 ( .A(n19469), .B(n19468), .Z(n19470) );
  AND U21283 ( .A(n19471), .B(n19470), .Z(n19480) );
  AND U21284 ( .A(y[7872]), .B(x[486]), .Z(n19473) );
  NAND U21285 ( .A(y[7878]), .B(x[480]), .Z(n19472) );
  XNOR U21286 ( .A(n19473), .B(n19472), .Z(n19486) );
  NAND U21287 ( .A(n19474), .B(o[197]), .Z(n19487) );
  NAND U21288 ( .A(y[7876]), .B(x[482]), .Z(n19475) );
  XNOR U21289 ( .A(n19476), .B(n19475), .Z(n19491) );
  AND U21290 ( .A(y[7877]), .B(x[481]), .Z(n19723) );
  NAND U21291 ( .A(y[7874]), .B(x[484]), .Z(n19477) );
  XNOR U21292 ( .A(n19723), .B(n19477), .Z(n19495) );
  AND U21293 ( .A(x[485]), .B(y[7873]), .Z(n19502) );
  XOR U21294 ( .A(o[198]), .B(n19502), .Z(n19494) );
  XOR U21295 ( .A(n19495), .B(n19494), .Z(n19490) );
  XOR U21296 ( .A(n19491), .B(n19490), .Z(n19481) );
  XOR U21297 ( .A(n19482), .B(n19481), .Z(n19508) );
  XOR U21298 ( .A(n19509), .B(n19508), .Z(n19505) );
  XNOR U21299 ( .A(n19504), .B(n19505), .Z(n19478) );
  XOR U21300 ( .A(n19503), .B(n19478), .Z(N423) );
  NANDN U21301 ( .A(n19480), .B(n19479), .Z(n19484) );
  NAND U21302 ( .A(n19482), .B(n19481), .Z(n19483) );
  AND U21303 ( .A(n19484), .B(n19483), .Z(n19548) );
  AND U21304 ( .A(y[7874]), .B(x[485]), .Z(n19605) );
  NAND U21305 ( .A(y[7878]), .B(x[481]), .Z(n19485) );
  XNOR U21306 ( .A(n19605), .B(n19485), .Z(n19521) );
  AND U21307 ( .A(x[486]), .B(y[7873]), .Z(n19525) );
  XOR U21308 ( .A(o[199]), .B(n19525), .Z(n19520) );
  XOR U21309 ( .A(n19521), .B(n19520), .Z(n19540) );
  AND U21310 ( .A(x[486]), .B(y[7878]), .Z(n19744) );
  NAND U21311 ( .A(n19997), .B(n19744), .Z(n19489) );
  NANDN U21312 ( .A(n19487), .B(n19486), .Z(n19488) );
  AND U21313 ( .A(n19489), .B(n19488), .Z(n19539) );
  NANDN U21314 ( .A(n19528), .B(n19529), .Z(n19493) );
  NAND U21315 ( .A(n19491), .B(n19490), .Z(n19492) );
  NAND U21316 ( .A(n19493), .B(n19492), .Z(n19542) );
  AND U21317 ( .A(x[484]), .B(y[7877]), .Z(n20002) );
  NAND U21318 ( .A(n20002), .B(n19519), .Z(n19497) );
  NAND U21319 ( .A(n19495), .B(n19494), .Z(n19496) );
  AND U21320 ( .A(n19497), .B(n19496), .Z(n19516) );
  AND U21321 ( .A(y[7877]), .B(x[482]), .Z(n19499) );
  NAND U21322 ( .A(y[7875]), .B(x[484]), .Z(n19498) );
  XNOR U21323 ( .A(n19499), .B(n19498), .Z(n19530) );
  XNOR U21324 ( .A(n19530), .B(n19529), .Z(n19514) );
  AND U21325 ( .A(y[7872]), .B(x[487]), .Z(n19501) );
  NAND U21326 ( .A(y[7879]), .B(x[480]), .Z(n19500) );
  XNOR U21327 ( .A(n19501), .B(n19500), .Z(n19534) );
  AND U21328 ( .A(o[198]), .B(n19502), .Z(n19533) );
  XNOR U21329 ( .A(n19534), .B(n19533), .Z(n19513) );
  XOR U21330 ( .A(n19514), .B(n19513), .Z(n19515) );
  XOR U21331 ( .A(n19516), .B(n19515), .Z(n19545) );
  XOR U21332 ( .A(n19546), .B(n19545), .Z(n19547) );
  XNOR U21333 ( .A(n19548), .B(n19547), .Z(n19553) );
  NAND U21334 ( .A(n19507), .B(n19506), .Z(n19511) );
  NAND U21335 ( .A(n19509), .B(n19508), .Z(n19510) );
  AND U21336 ( .A(n19511), .B(n19510), .Z(n19551) );
  XOR U21337 ( .A(n19552), .B(n19551), .Z(n19512) );
  XNOR U21338 ( .A(n19553), .B(n19512), .Z(N424) );
  NAND U21339 ( .A(n19514), .B(n19513), .Z(n19518) );
  NAND U21340 ( .A(n19516), .B(n19515), .Z(n19517) );
  AND U21341 ( .A(n19518), .B(n19517), .Z(n19586) );
  AND U21342 ( .A(x[485]), .B(y[7878]), .Z(n19694) );
  NAND U21343 ( .A(n19694), .B(n19519), .Z(n19523) );
  NAND U21344 ( .A(n19521), .B(n19520), .Z(n19522) );
  NAND U21345 ( .A(n19523), .B(n19522), .Z(n19584) );
  AND U21346 ( .A(x[485]), .B(y[7875]), .Z(n20143) );
  NAND U21347 ( .A(y[7879]), .B(x[481]), .Z(n19524) );
  XNOR U21348 ( .A(n20143), .B(n19524), .Z(n19567) );
  AND U21349 ( .A(o[199]), .B(n19525), .Z(n19566) );
  XOR U21350 ( .A(n19567), .B(n19566), .Z(n19572) );
  NAND U21351 ( .A(x[483]), .B(y[7877]), .Z(n20337) );
  AND U21352 ( .A(y[7874]), .B(x[486]), .Z(n19527) );
  NAND U21353 ( .A(y[7878]), .B(x[482]), .Z(n19526) );
  XNOR U21354 ( .A(n19527), .B(n19526), .Z(n19574) );
  XNOR U21355 ( .A(n20201), .B(n19574), .Z(n19570) );
  XOR U21356 ( .A(n20337), .B(n19570), .Z(n19571) );
  XOR U21357 ( .A(n19572), .B(n19571), .Z(n19583) );
  XOR U21358 ( .A(n19584), .B(n19583), .Z(n19585) );
  XOR U21359 ( .A(n19586), .B(n19585), .Z(n19592) );
  NANDN U21360 ( .A(n19528), .B(n20002), .Z(n19532) );
  NAND U21361 ( .A(n19530), .B(n19529), .Z(n19531) );
  NAND U21362 ( .A(n19532), .B(n19531), .Z(n19580) );
  AND U21363 ( .A(x[487]), .B(y[7879]), .Z(n19881) );
  NAND U21364 ( .A(n19997), .B(n19881), .Z(n19536) );
  NAND U21365 ( .A(n19534), .B(n19533), .Z(n19535) );
  NAND U21366 ( .A(n19536), .B(n19535), .Z(n19578) );
  AND U21367 ( .A(y[7872]), .B(x[488]), .Z(n19538) );
  NAND U21368 ( .A(y[7880]), .B(x[480]), .Z(n19537) );
  XNOR U21369 ( .A(n19538), .B(n19537), .Z(n19557) );
  AND U21370 ( .A(x[487]), .B(y[7873]), .Z(n19562) );
  XOR U21371 ( .A(o[200]), .B(n19562), .Z(n19556) );
  XOR U21372 ( .A(n19557), .B(n19556), .Z(n19577) );
  XOR U21373 ( .A(n19578), .B(n19577), .Z(n19579) );
  XNOR U21374 ( .A(n19580), .B(n19579), .Z(n19590) );
  NANDN U21375 ( .A(n19540), .B(n19539), .Z(n19544) );
  NANDN U21376 ( .A(n19542), .B(n19541), .Z(n19543) );
  NAND U21377 ( .A(n19544), .B(n19543), .Z(n19589) );
  XOR U21378 ( .A(n19590), .B(n19589), .Z(n19591) );
  XOR U21379 ( .A(n19592), .B(n19591), .Z(n19597) );
  NAND U21380 ( .A(n19546), .B(n19545), .Z(n19550) );
  NAND U21381 ( .A(n19548), .B(n19547), .Z(n19549) );
  NAND U21382 ( .A(n19550), .B(n19549), .Z(n19595) );
  XOR U21383 ( .A(n19595), .B(n19596), .Z(n19554) );
  XNOR U21384 ( .A(n19597), .B(n19554), .Z(N425) );
  AND U21385 ( .A(x[488]), .B(y[7880]), .Z(n19555) );
  NAND U21386 ( .A(n19555), .B(n19997), .Z(n19559) );
  NAND U21387 ( .A(n19557), .B(n19556), .Z(n19558) );
  AND U21388 ( .A(n19559), .B(n19558), .Z(n19634) );
  AND U21389 ( .A(y[7876]), .B(x[485]), .Z(n19561) );
  NAND U21390 ( .A(y[7874]), .B(x[487]), .Z(n19560) );
  XNOR U21391 ( .A(n19561), .B(n19560), .Z(n19607) );
  AND U21392 ( .A(o[200]), .B(n19562), .Z(n19606) );
  XNOR U21393 ( .A(n19607), .B(n19606), .Z(n19632) );
  AND U21394 ( .A(y[7872]), .B(x[489]), .Z(n19564) );
  NAND U21395 ( .A(y[7881]), .B(x[480]), .Z(n19563) );
  XNOR U21396 ( .A(n19564), .B(n19563), .Z(n19614) );
  AND U21397 ( .A(x[488]), .B(y[7873]), .Z(n19623) );
  XOR U21398 ( .A(o[201]), .B(n19623), .Z(n19613) );
  XNOR U21399 ( .A(n19614), .B(n19613), .Z(n19631) );
  XOR U21400 ( .A(n19632), .B(n19631), .Z(n19633) );
  XNOR U21401 ( .A(n19634), .B(n19633), .Z(n19628) );
  AND U21402 ( .A(y[7875]), .B(x[486]), .Z(n19951) );
  NAND U21403 ( .A(y[7880]), .B(x[481]), .Z(n19565) );
  XNOR U21404 ( .A(n19951), .B(n19565), .Z(n19618) );
  XNOR U21405 ( .A(n20002), .B(n19618), .Z(n19637) );
  NAND U21406 ( .A(x[482]), .B(y[7879]), .Z(n20117) );
  NAND U21407 ( .A(x[483]), .B(y[7878]), .Z(n19959) );
  XNOR U21408 ( .A(n20117), .B(n19959), .Z(n19638) );
  XOR U21409 ( .A(n19637), .B(n19638), .Z(n19626) );
  NAND U21410 ( .A(x[485]), .B(y[7879]), .Z(n19810) );
  AND U21411 ( .A(x[481]), .B(y[7875]), .Z(n19617) );
  NANDN U21412 ( .A(n19810), .B(n19617), .Z(n19569) );
  NAND U21413 ( .A(n19567), .B(n19566), .Z(n19568) );
  NAND U21414 ( .A(n19569), .B(n19568), .Z(n19625) );
  XOR U21415 ( .A(n19626), .B(n19625), .Z(n19627) );
  XNOR U21416 ( .A(n19628), .B(n19627), .Z(n19601) );
  NAND U21417 ( .A(n19744), .B(n19573), .Z(n19576) );
  NAND U21418 ( .A(n20201), .B(n19574), .Z(n19575) );
  AND U21419 ( .A(n19576), .B(n19575), .Z(n19599) );
  XOR U21420 ( .A(n19600), .B(n19599), .Z(n19602) );
  XNOR U21421 ( .A(n19601), .B(n19602), .Z(n19643) );
  NAND U21422 ( .A(n19578), .B(n19577), .Z(n19582) );
  NAND U21423 ( .A(n19580), .B(n19579), .Z(n19581) );
  NAND U21424 ( .A(n19582), .B(n19581), .Z(n19642) );
  NAND U21425 ( .A(n19584), .B(n19583), .Z(n19588) );
  NAND U21426 ( .A(n19586), .B(n19585), .Z(n19587) );
  NAND U21427 ( .A(n19588), .B(n19587), .Z(n19641) );
  XOR U21428 ( .A(n19642), .B(n19641), .Z(n19644) );
  XOR U21429 ( .A(n19643), .B(n19644), .Z(n19649) );
  NAND U21430 ( .A(n19590), .B(n19589), .Z(n19594) );
  NANDN U21431 ( .A(n19592), .B(n19591), .Z(n19593) );
  NAND U21432 ( .A(n19594), .B(n19593), .Z(n19647) );
  XOR U21433 ( .A(n19647), .B(n19648), .Z(n19598) );
  XNOR U21434 ( .A(n19649), .B(n19598), .Z(N426) );
  NAND U21435 ( .A(n19600), .B(n19599), .Z(n19604) );
  NAND U21436 ( .A(n19602), .B(n19601), .Z(n19603) );
  NAND U21437 ( .A(n19604), .B(n19603), .Z(n19654) );
  AND U21438 ( .A(x[487]), .B(y[7876]), .Z(n19696) );
  NAND U21439 ( .A(n19696), .B(n19605), .Z(n19609) );
  NAND U21440 ( .A(n19607), .B(n19606), .Z(n19608) );
  AND U21441 ( .A(n19609), .B(n19608), .Z(n19709) );
  AND U21442 ( .A(y[7875]), .B(x[487]), .Z(n19611) );
  NAND U21443 ( .A(y[7878]), .B(x[484]), .Z(n19610) );
  XNOR U21444 ( .A(n19611), .B(n19610), .Z(n19680) );
  AND U21445 ( .A(x[486]), .B(y[7876]), .Z(n19679) );
  XOR U21446 ( .A(n19680), .B(n19679), .Z(n19707) );
  AND U21447 ( .A(x[488]), .B(y[7874]), .Z(n19861) );
  AND U21448 ( .A(x[489]), .B(y[7873]), .Z(n19690) );
  XOR U21449 ( .A(o[202]), .B(n19690), .Z(n19701) );
  XOR U21450 ( .A(n19861), .B(n19701), .Z(n19703) );
  XNOR U21451 ( .A(n19703), .B(n19702), .Z(n19706) );
  XNOR U21452 ( .A(n19709), .B(n19708), .Z(n19668) );
  AND U21453 ( .A(x[489]), .B(y[7881]), .Z(n19612) );
  NAND U21454 ( .A(n19612), .B(n19997), .Z(n19616) );
  NAND U21455 ( .A(n19614), .B(n19613), .Z(n19615) );
  NAND U21456 ( .A(n19616), .B(n19615), .Z(n19666) );
  AND U21457 ( .A(x[486]), .B(y[7880]), .Z(n19887) );
  NAND U21458 ( .A(n19887), .B(n19617), .Z(n19620) );
  NAND U21459 ( .A(n19618), .B(n20002), .Z(n19619) );
  AND U21460 ( .A(n19620), .B(n19619), .Z(n19675) );
  AND U21461 ( .A(y[7872]), .B(x[490]), .Z(n19622) );
  NAND U21462 ( .A(y[7882]), .B(x[480]), .Z(n19621) );
  XNOR U21463 ( .A(n19622), .B(n19621), .Z(n19685) );
  AND U21464 ( .A(o[201]), .B(n19623), .Z(n19684) );
  XOR U21465 ( .A(n19685), .B(n19684), .Z(n19673) );
  AND U21466 ( .A(x[483]), .B(y[7879]), .Z(n20562) );
  NAND U21467 ( .A(y[7881]), .B(x[481]), .Z(n19624) );
  XNOR U21468 ( .A(n20562), .B(n19624), .Z(n19697) );
  NAND U21469 ( .A(x[482]), .B(y[7880]), .Z(n19698) );
  XOR U21470 ( .A(n19673), .B(n19672), .Z(n19674) );
  XOR U21471 ( .A(n19666), .B(n19667), .Z(n19669) );
  XOR U21472 ( .A(n19668), .B(n19669), .Z(n19652) );
  NAND U21473 ( .A(n19626), .B(n19625), .Z(n19630) );
  NAND U21474 ( .A(n19628), .B(n19627), .Z(n19629) );
  NAND U21475 ( .A(n19630), .B(n19629), .Z(n19662) );
  NAND U21476 ( .A(n19632), .B(n19631), .Z(n19636) );
  NAND U21477 ( .A(n19634), .B(n19633), .Z(n19635) );
  AND U21478 ( .A(n19636), .B(n19635), .Z(n19661) );
  NANDN U21479 ( .A(n19638), .B(n19637), .Z(n19640) );
  IV U21480 ( .A(n20117), .Z(n20248) );
  ANDN U21481 ( .B(n19959), .A(n20248), .Z(n19639) );
  ANDN U21482 ( .B(n19640), .A(n19639), .Z(n19660) );
  XOR U21483 ( .A(n19661), .B(n19660), .Z(n19663) );
  XNOR U21484 ( .A(n19662), .B(n19663), .Z(n19651) );
  XOR U21485 ( .A(n19652), .B(n19651), .Z(n19653) );
  XOR U21486 ( .A(n19654), .B(n19653), .Z(n19659) );
  NAND U21487 ( .A(n19642), .B(n19641), .Z(n19646) );
  NAND U21488 ( .A(n19644), .B(n19643), .Z(n19645) );
  NAND U21489 ( .A(n19646), .B(n19645), .Z(n19658) );
  XOR U21490 ( .A(n19658), .B(n19657), .Z(n19650) );
  XNOR U21491 ( .A(n19659), .B(n19650), .Z(N427) );
  NAND U21492 ( .A(n19652), .B(n19651), .Z(n19656) );
  NAND U21493 ( .A(n19654), .B(n19653), .Z(n19655) );
  NAND U21494 ( .A(n19656), .B(n19655), .Z(n19770) );
  IV U21495 ( .A(n19770), .Z(n19768) );
  NAND U21496 ( .A(n19661), .B(n19660), .Z(n19665) );
  NAND U21497 ( .A(n19663), .B(n19662), .Z(n19664) );
  NAND U21498 ( .A(n19665), .B(n19664), .Z(n19777) );
  NANDN U21499 ( .A(n19667), .B(n19666), .Z(n19671) );
  NANDN U21500 ( .A(n19669), .B(n19668), .Z(n19670) );
  NAND U21501 ( .A(n19671), .B(n19670), .Z(n19776) );
  NAND U21502 ( .A(n19673), .B(n19672), .Z(n19677) );
  NANDN U21503 ( .A(n19675), .B(n19674), .Z(n19676) );
  AND U21504 ( .A(n19677), .B(n19676), .Z(n19765) );
  AND U21505 ( .A(x[487]), .B(y[7878]), .Z(n19806) );
  AND U21506 ( .A(x[484]), .B(y[7875]), .Z(n19678) );
  NAND U21507 ( .A(n19806), .B(n19678), .Z(n19682) );
  NAND U21508 ( .A(n19680), .B(n19679), .Z(n19681) );
  AND U21509 ( .A(n19682), .B(n19681), .Z(n19763) );
  AND U21510 ( .A(x[490]), .B(y[7882]), .Z(n19683) );
  NAND U21511 ( .A(n19683), .B(n19997), .Z(n19687) );
  NAND U21512 ( .A(n19685), .B(n19684), .Z(n19686) );
  AND U21513 ( .A(n19687), .B(n19686), .Z(n19759) );
  AND U21514 ( .A(y[7872]), .B(x[491]), .Z(n19689) );
  NAND U21515 ( .A(y[7883]), .B(x[480]), .Z(n19688) );
  XNOR U21516 ( .A(n19689), .B(n19688), .Z(n19735) );
  AND U21517 ( .A(o[202]), .B(n19690), .Z(n19734) );
  XOR U21518 ( .A(n19735), .B(n19734), .Z(n19757) );
  AND U21519 ( .A(y[7877]), .B(x[486]), .Z(n19692) );
  NAND U21520 ( .A(y[7882]), .B(x[481]), .Z(n19691) );
  XNOR U21521 ( .A(n19692), .B(n19691), .Z(n19725) );
  AND U21522 ( .A(x[490]), .B(y[7873]), .Z(n19743) );
  XOR U21523 ( .A(o[203]), .B(n19743), .Z(n19724) );
  XOR U21524 ( .A(n19725), .B(n19724), .Z(n19756) );
  XOR U21525 ( .A(n19757), .B(n19756), .Z(n19758) );
  NAND U21526 ( .A(x[483]), .B(y[7880]), .Z(n20691) );
  NAND U21527 ( .A(y[7881]), .B(x[482]), .Z(n19693) );
  XNOR U21528 ( .A(n19694), .B(n19693), .Z(n19720) );
  AND U21529 ( .A(x[484]), .B(y[7879]), .Z(n19719) );
  XNOR U21530 ( .A(n19720), .B(n19719), .Z(n19751) );
  XOR U21531 ( .A(n20691), .B(n19751), .Z(n19753) );
  NAND U21532 ( .A(y[7874]), .B(x[489]), .Z(n19695) );
  XNOR U21533 ( .A(n19696), .B(n19695), .Z(n19740) );
  AND U21534 ( .A(x[488]), .B(y[7875]), .Z(n19739) );
  XNOR U21535 ( .A(n19740), .B(n19739), .Z(n19752) );
  XOR U21536 ( .A(n19753), .B(n19752), .Z(n19716) );
  AND U21537 ( .A(x[483]), .B(y[7881]), .Z(n19733) );
  IV U21538 ( .A(n19733), .Z(n19801) );
  AND U21539 ( .A(x[481]), .B(y[7879]), .Z(n19992) );
  NANDN U21540 ( .A(n19801), .B(n19992), .Z(n19700) );
  NANDN U21541 ( .A(n19698), .B(n19697), .Z(n19699) );
  AND U21542 ( .A(n19700), .B(n19699), .Z(n19714) );
  NAND U21543 ( .A(n19861), .B(n19701), .Z(n19705) );
  NAND U21544 ( .A(n19703), .B(n19702), .Z(n19704) );
  NAND U21545 ( .A(n19705), .B(n19704), .Z(n19713) );
  NANDN U21546 ( .A(n19707), .B(n19706), .Z(n19711) );
  NAND U21547 ( .A(n19709), .B(n19708), .Z(n19710) );
  NAND U21548 ( .A(n19711), .B(n19710), .Z(n19745) );
  XOR U21549 ( .A(n19746), .B(n19745), .Z(n19748) );
  XNOR U21550 ( .A(n19747), .B(n19748), .Z(n19775) );
  XOR U21551 ( .A(n19776), .B(n19775), .Z(n19778) );
  XOR U21552 ( .A(n19777), .B(n19778), .Z(n19771) );
  XNOR U21553 ( .A(n19769), .B(n19771), .Z(n19712) );
  XOR U21554 ( .A(n19768), .B(n19712), .Z(N428) );
  NANDN U21555 ( .A(n19714), .B(n19713), .Z(n19718) );
  NANDN U21556 ( .A(n19716), .B(n19715), .Z(n19717) );
  AND U21557 ( .A(n19718), .B(n19717), .Z(n19838) );
  AND U21558 ( .A(x[482]), .B(y[7878]), .Z(n20409) );
  AND U21559 ( .A(x[485]), .B(y[7881]), .Z(n20239) );
  NAND U21560 ( .A(n20409), .B(n20239), .Z(n19722) );
  NAND U21561 ( .A(n19720), .B(n19719), .Z(n19721) );
  NAND U21562 ( .A(n19722), .B(n19721), .Z(n19789) );
  AND U21563 ( .A(x[486]), .B(y[7882]), .Z(n20009) );
  NAND U21564 ( .A(n20009), .B(n19723), .Z(n19727) );
  NAND U21565 ( .A(n19725), .B(n19724), .Z(n19726) );
  NAND U21566 ( .A(n19727), .B(n19726), .Z(n19788) );
  XOR U21567 ( .A(n19789), .B(n19788), .Z(n19791) );
  AND U21568 ( .A(x[489]), .B(y[7875]), .Z(n20404) );
  AND U21569 ( .A(x[490]), .B(y[7874]), .Z(n20448) );
  AND U21570 ( .A(y[7880]), .B(x[484]), .Z(n19728) );
  XOR U21571 ( .A(n20448), .B(n19728), .Z(n19828) );
  XOR U21572 ( .A(n20404), .B(n19828), .Z(n19811) );
  NAND U21573 ( .A(x[487]), .B(y[7877]), .Z(n19809) );
  XOR U21574 ( .A(n19810), .B(n19809), .Z(n19812) );
  AND U21575 ( .A(y[7872]), .B(x[492]), .Z(n19730) );
  NAND U21576 ( .A(y[7884]), .B(x[480]), .Z(n19729) );
  XNOR U21577 ( .A(n19730), .B(n19729), .Z(n19824) );
  AND U21578 ( .A(x[491]), .B(y[7873]), .Z(n19804) );
  XOR U21579 ( .A(n19804), .B(o[204]), .Z(n19823) );
  XOR U21580 ( .A(n19824), .B(n19823), .Z(n19795) );
  AND U21581 ( .A(y[7882]), .B(x[482]), .Z(n19732) );
  NAND U21582 ( .A(y[7876]), .B(x[488]), .Z(n19731) );
  XNOR U21583 ( .A(n19732), .B(n19731), .Z(n19800) );
  XOR U21584 ( .A(n19800), .B(n19733), .Z(n19794) );
  XOR U21585 ( .A(n19795), .B(n19794), .Z(n19797) );
  XOR U21586 ( .A(n19796), .B(n19797), .Z(n19790) );
  XOR U21587 ( .A(n19791), .B(n19790), .Z(n19836) );
  AND U21588 ( .A(x[491]), .B(y[7883]), .Z(n20810) );
  NAND U21589 ( .A(n20810), .B(n19997), .Z(n19737) );
  NAND U21590 ( .A(n19735), .B(n19734), .Z(n19736) );
  NAND U21591 ( .A(n19737), .B(n19736), .Z(n19818) );
  AND U21592 ( .A(x[489]), .B(y[7876]), .Z(n19738) );
  AND U21593 ( .A(x[487]), .B(y[7874]), .Z(n19937) );
  NAND U21594 ( .A(n19738), .B(n19937), .Z(n19742) );
  NAND U21595 ( .A(n19740), .B(n19739), .Z(n19741) );
  NAND U21596 ( .A(n19742), .B(n19741), .Z(n19816) );
  AND U21597 ( .A(x[481]), .B(y[7883]), .Z(n20443) );
  XOR U21598 ( .A(n19744), .B(n20443), .Z(n19821) );
  XOR U21599 ( .A(n19822), .B(n19821), .Z(n19815) );
  XOR U21600 ( .A(n19816), .B(n19815), .Z(n19817) );
  XOR U21601 ( .A(n19818), .B(n19817), .Z(n19835) );
  XOR U21602 ( .A(n19836), .B(n19835), .Z(n19837) );
  NAND U21603 ( .A(n19746), .B(n19745), .Z(n19750) );
  NAND U21604 ( .A(n19748), .B(n19747), .Z(n19749) );
  NAND U21605 ( .A(n19750), .B(n19749), .Z(n19841) );
  XOR U21606 ( .A(n19842), .B(n19841), .Z(n19844) );
  IV U21607 ( .A(n20691), .Z(n20418) );
  NANDN U21608 ( .A(n20418), .B(n19751), .Z(n19755) );
  NAND U21609 ( .A(n19753), .B(n19752), .Z(n19754) );
  AND U21610 ( .A(n19755), .B(n19754), .Z(n19783) );
  NAND U21611 ( .A(n19757), .B(n19756), .Z(n19761) );
  NANDN U21612 ( .A(n19759), .B(n19758), .Z(n19760) );
  AND U21613 ( .A(n19761), .B(n19760), .Z(n19782) );
  NANDN U21614 ( .A(n19763), .B(n19762), .Z(n19767) );
  NANDN U21615 ( .A(n19765), .B(n19764), .Z(n19766) );
  NAND U21616 ( .A(n19767), .B(n19766), .Z(n19785) );
  XNOR U21617 ( .A(n19844), .B(n19843), .Z(n19849) );
  NANDN U21618 ( .A(n19768), .B(n19769), .Z(n19774) );
  NOR U21619 ( .A(n19770), .B(n19769), .Z(n19772) );
  OR U21620 ( .A(n19772), .B(n19771), .Z(n19773) );
  AND U21621 ( .A(n19774), .B(n19773), .Z(n19848) );
  NAND U21622 ( .A(n19776), .B(n19775), .Z(n19780) );
  NAND U21623 ( .A(n19778), .B(n19777), .Z(n19779) );
  AND U21624 ( .A(n19780), .B(n19779), .Z(n19847) );
  XOR U21625 ( .A(n19848), .B(n19847), .Z(n19781) );
  XNOR U21626 ( .A(n19849), .B(n19781), .Z(N429) );
  NANDN U21627 ( .A(n19783), .B(n19782), .Z(n19787) );
  NANDN U21628 ( .A(n19785), .B(n19784), .Z(n19786) );
  AND U21629 ( .A(n19787), .B(n19786), .Z(n19909) );
  NAND U21630 ( .A(n19789), .B(n19788), .Z(n19793) );
  NAND U21631 ( .A(n19791), .B(n19790), .Z(n19792) );
  NAND U21632 ( .A(n19793), .B(n19792), .Z(n19895) );
  NAND U21633 ( .A(n19795), .B(n19794), .Z(n19799) );
  NAND U21634 ( .A(n19797), .B(n19796), .Z(n19798) );
  NAND U21635 ( .A(n19799), .B(n19798), .Z(n19902) );
  AND U21636 ( .A(y[7882]), .B(x[488]), .Z(n21094) );
  AND U21637 ( .A(x[482]), .B(y[7876]), .Z(n19947) );
  NAND U21638 ( .A(n21094), .B(n19947), .Z(n19803) );
  NANDN U21639 ( .A(n19801), .B(n19800), .Z(n19802) );
  NAND U21640 ( .A(n19803), .B(n19802), .Z(n19871) );
  AND U21641 ( .A(n19804), .B(o[204]), .Z(n19865) );
  AND U21642 ( .A(y[7884]), .B(x[481]), .Z(n19805) );
  XOR U21643 ( .A(n19806), .B(n19805), .Z(n19864) );
  XOR U21644 ( .A(n19865), .B(n19864), .Z(n19870) );
  AND U21645 ( .A(x[486]), .B(y[7879]), .Z(n20850) );
  AND U21646 ( .A(y[7883]), .B(x[482]), .Z(n19808) );
  NAND U21647 ( .A(y[7876]), .B(x[489]), .Z(n19807) );
  XNOR U21648 ( .A(n19808), .B(n19807), .Z(n19874) );
  XOR U21649 ( .A(n20850), .B(n19874), .Z(n19869) );
  XOR U21650 ( .A(n19870), .B(n19869), .Z(n19872) );
  XOR U21651 ( .A(n19871), .B(n19872), .Z(n19901) );
  NAND U21652 ( .A(n19810), .B(n19809), .Z(n19814) );
  ANDN U21653 ( .B(n19812), .A(n19811), .Z(n19813) );
  ANDN U21654 ( .B(n19814), .A(n19813), .Z(n19900) );
  XOR U21655 ( .A(n19901), .B(n19900), .Z(n19903) );
  XOR U21656 ( .A(n19902), .B(n19903), .Z(n19894) );
  XOR U21657 ( .A(n19895), .B(n19894), .Z(n19897) );
  NAND U21658 ( .A(n19816), .B(n19815), .Z(n19820) );
  NAND U21659 ( .A(n19818), .B(n19817), .Z(n19819) );
  NAND U21660 ( .A(n19820), .B(n19819), .Z(n19853) );
  NAND U21661 ( .A(x[486]), .B(y[7883]), .Z(n20241) );
  AND U21662 ( .A(x[481]), .B(y[7878]), .Z(n19863) );
  AND U21663 ( .A(x[492]), .B(y[7884]), .Z(n21100) );
  AND U21664 ( .A(x[490]), .B(y[7875]), .Z(n20703) );
  AND U21665 ( .A(x[491]), .B(y[7874]), .Z(n20664) );
  AND U21666 ( .A(y[7877]), .B(x[488]), .Z(n19825) );
  XOR U21667 ( .A(n20664), .B(n19825), .Z(n19862) );
  XOR U21668 ( .A(n20703), .B(n19862), .Z(n19858) );
  XOR U21669 ( .A(n19857), .B(n19858), .Z(n19860) );
  XOR U21670 ( .A(n19859), .B(n19860), .Z(n19851) );
  AND U21671 ( .A(x[490]), .B(y[7880]), .Z(n19827) );
  AND U21672 ( .A(x[484]), .B(y[7874]), .Z(n19826) );
  NAND U21673 ( .A(n19827), .B(n19826), .Z(n19830) );
  NAND U21674 ( .A(n20404), .B(n19828), .Z(n19829) );
  NAND U21675 ( .A(n19830), .B(n19829), .Z(n19890) );
  AND U21676 ( .A(y[7872]), .B(x[493]), .Z(n19832) );
  NAND U21677 ( .A(y[7885]), .B(x[480]), .Z(n19831) );
  XNOR U21678 ( .A(n19832), .B(n19831), .Z(n19885) );
  AND U21679 ( .A(x[492]), .B(y[7873]), .Z(n19877) );
  XOR U21680 ( .A(n19877), .B(o[205]), .Z(n19884) );
  XOR U21681 ( .A(n19885), .B(n19884), .Z(n19889) );
  AND U21682 ( .A(y[7880]), .B(x[485]), .Z(n19834) );
  NAND U21683 ( .A(y[7882]), .B(x[483]), .Z(n19833) );
  XNOR U21684 ( .A(n19834), .B(n19833), .Z(n19883) );
  AND U21685 ( .A(x[484]), .B(y[7881]), .Z(n19882) );
  XOR U21686 ( .A(n19883), .B(n19882), .Z(n19888) );
  XOR U21687 ( .A(n19889), .B(n19888), .Z(n19891) );
  XOR U21688 ( .A(n19890), .B(n19891), .Z(n19852) );
  XOR U21689 ( .A(n19851), .B(n19852), .Z(n19854) );
  XOR U21690 ( .A(n19853), .B(n19854), .Z(n19896) );
  XOR U21691 ( .A(n19897), .B(n19896), .Z(n19907) );
  NAND U21692 ( .A(n19836), .B(n19835), .Z(n19840) );
  NANDN U21693 ( .A(n19838), .B(n19837), .Z(n19839) );
  AND U21694 ( .A(n19840), .B(n19839), .Z(n19906) );
  XOR U21695 ( .A(n19909), .B(n19908), .Z(n19915) );
  NAND U21696 ( .A(n19842), .B(n19841), .Z(n19846) );
  NAND U21697 ( .A(n19844), .B(n19843), .Z(n19845) );
  NAND U21698 ( .A(n19846), .B(n19845), .Z(n19913) );
  IV U21699 ( .A(n19914), .Z(n19912) );
  XOR U21700 ( .A(n19913), .B(n19912), .Z(n19850) );
  XNOR U21701 ( .A(n19915), .B(n19850), .Z(N430) );
  NAND U21702 ( .A(n19852), .B(n19851), .Z(n19856) );
  NAND U21703 ( .A(n19854), .B(n19853), .Z(n19855) );
  NAND U21704 ( .A(n19856), .B(n19855), .Z(n19919) );
  AND U21705 ( .A(x[491]), .B(y[7877]), .Z(n20021) );
  NAND U21706 ( .A(x[487]), .B(y[7884]), .Z(n20420) );
  XOR U21707 ( .A(n19972), .B(n19973), .Z(n19975) );
  AND U21708 ( .A(x[484]), .B(y[7882]), .Z(n20346) );
  AND U21709 ( .A(y[7883]), .B(x[483]), .Z(n19867) );
  NAND U21710 ( .A(y[7878]), .B(x[488]), .Z(n19866) );
  XNOR U21711 ( .A(n19867), .B(n19866), .Z(n19960) );
  XOR U21712 ( .A(n20239), .B(n19960), .Z(n19969) );
  XOR U21713 ( .A(n20346), .B(n19969), .Z(n19971) );
  AND U21714 ( .A(x[489]), .B(y[7877]), .Z(n20539) );
  AND U21715 ( .A(x[482]), .B(y[7884]), .Z(n19868) );
  AND U21716 ( .A(x[490]), .B(y[7876]), .Z(n20557) );
  XOR U21717 ( .A(n19868), .B(n20557), .Z(n19948) );
  XOR U21718 ( .A(n20539), .B(n19948), .Z(n19970) );
  XOR U21719 ( .A(n19971), .B(n19970), .Z(n19974) );
  XOR U21720 ( .A(n19975), .B(n19974), .Z(n19924) );
  XOR U21721 ( .A(n19924), .B(n19923), .Z(n19926) );
  XOR U21722 ( .A(n19925), .B(n19926), .Z(n19918) );
  AND U21723 ( .A(x[489]), .B(y[7883]), .Z(n19873) );
  NAND U21724 ( .A(n19873), .B(n19947), .Z(n19876) );
  NAND U21725 ( .A(n20850), .B(n19874), .Z(n19875) );
  NAND U21726 ( .A(n19876), .B(n19875), .Z(n19935) );
  AND U21727 ( .A(n19877), .B(o[205]), .Z(n19957) );
  AND U21728 ( .A(x[494]), .B(y[7872]), .Z(n19879) );
  AND U21729 ( .A(y[7886]), .B(x[480]), .Z(n19878) );
  XOR U21730 ( .A(n19879), .B(n19878), .Z(n19956) );
  XOR U21731 ( .A(n19957), .B(n19956), .Z(n19934) );
  NAND U21732 ( .A(y[7874]), .B(x[492]), .Z(n19880) );
  XNOR U21733 ( .A(n19881), .B(n19880), .Z(n19939) );
  AND U21734 ( .A(x[493]), .B(y[7873]), .Z(n19944) );
  XOR U21735 ( .A(o[206]), .B(n19944), .Z(n19938) );
  XOR U21736 ( .A(n19939), .B(n19938), .Z(n19933) );
  XOR U21737 ( .A(n19934), .B(n19933), .Z(n19936) );
  XNOR U21738 ( .A(n19935), .B(n19936), .Z(n19977) );
  NAND U21739 ( .A(x[485]), .B(y[7882]), .Z(n20010) );
  AND U21740 ( .A(x[493]), .B(y[7885]), .Z(n21407) );
  NAND U21741 ( .A(y[7875]), .B(x[491]), .Z(n19886) );
  XNOR U21742 ( .A(n19887), .B(n19886), .Z(n19953) );
  AND U21743 ( .A(x[481]), .B(y[7885]), .Z(n19952) );
  XOR U21744 ( .A(n19953), .B(n19952), .Z(n19929) );
  XNOR U21745 ( .A(n19930), .B(n19929), .Z(n19932) );
  XOR U21746 ( .A(n19931), .B(n19932), .Z(n19976) );
  XOR U21747 ( .A(n19977), .B(n19976), .Z(n19979) );
  NAND U21748 ( .A(n19889), .B(n19888), .Z(n19893) );
  NAND U21749 ( .A(n19891), .B(n19890), .Z(n19892) );
  AND U21750 ( .A(n19893), .B(n19892), .Z(n19978) );
  XNOR U21751 ( .A(n19979), .B(n19978), .Z(n19917) );
  XOR U21752 ( .A(n19918), .B(n19917), .Z(n19920) );
  XOR U21753 ( .A(n19919), .B(n19920), .Z(n19985) );
  NAND U21754 ( .A(n19895), .B(n19894), .Z(n19899) );
  NAND U21755 ( .A(n19897), .B(n19896), .Z(n19898) );
  NAND U21756 ( .A(n19899), .B(n19898), .Z(n19983) );
  NAND U21757 ( .A(n19901), .B(n19900), .Z(n19905) );
  NAND U21758 ( .A(n19903), .B(n19902), .Z(n19904) );
  NAND U21759 ( .A(n19905), .B(n19904), .Z(n19982) );
  XOR U21760 ( .A(n19983), .B(n19982), .Z(n19984) );
  XOR U21761 ( .A(n19985), .B(n19984), .Z(n19990) );
  NANDN U21762 ( .A(n19907), .B(n19906), .Z(n19911) );
  NANDN U21763 ( .A(n19909), .B(n19908), .Z(n19910) );
  NAND U21764 ( .A(n19911), .B(n19910), .Z(n19988) );
  XOR U21765 ( .A(n19988), .B(n19989), .Z(n19916) );
  XNOR U21766 ( .A(n19990), .B(n19916), .Z(N431) );
  NAND U21767 ( .A(n19918), .B(n19917), .Z(n19922) );
  NAND U21768 ( .A(n19920), .B(n19919), .Z(n19921) );
  NAND U21769 ( .A(n19922), .B(n19921), .Z(n20075) );
  NANDN U21770 ( .A(n19924), .B(n19923), .Z(n19928) );
  NANDN U21771 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U21772 ( .A(n19928), .B(n19927), .Z(n20050) );
  NAND U21773 ( .A(x[492]), .B(y[7879]), .Z(n20411) );
  NANDN U21774 ( .A(n20411), .B(n19937), .Z(n19941) );
  NAND U21775 ( .A(n19939), .B(n19938), .Z(n19940) );
  AND U21776 ( .A(n19941), .B(n19940), .Z(n20030) );
  AND U21777 ( .A(y[7876]), .B(x[491]), .Z(n19943) );
  NAND U21778 ( .A(y[7874]), .B(x[493]), .Z(n19942) );
  XNOR U21779 ( .A(n19943), .B(n19942), .Z(n20035) );
  AND U21780 ( .A(x[492]), .B(y[7875]), .Z(n20034) );
  XNOR U21781 ( .A(n20035), .B(n20034), .Z(n20029) );
  AND U21782 ( .A(n19944), .B(o[206]), .Z(n19999) );
  AND U21783 ( .A(x[495]), .B(y[7872]), .Z(n19946) );
  AND U21784 ( .A(y[7887]), .B(x[480]), .Z(n19945) );
  XOR U21785 ( .A(n19946), .B(n19945), .Z(n19998) );
  XNOR U21786 ( .A(n19999), .B(n19998), .Z(n20028) );
  XNOR U21787 ( .A(n20029), .B(n20028), .Z(n20031) );
  XNOR U21788 ( .A(n20030), .B(n20031), .Z(n20061) );
  NAND U21789 ( .A(x[490]), .B(y[7884]), .Z(n20852) );
  NANDN U21790 ( .A(n20852), .B(n19947), .Z(n19950) );
  NAND U21791 ( .A(n20539), .B(n19948), .Z(n19949) );
  NAND U21792 ( .A(n19950), .B(n19949), .Z(n20059) );
  AND U21793 ( .A(y[7880]), .B(x[491]), .Z(n20345) );
  NAND U21794 ( .A(n20345), .B(n19951), .Z(n19955) );
  NAND U21795 ( .A(n19953), .B(n19952), .Z(n19954) );
  NAND U21796 ( .A(n19955), .B(n19954), .Z(n20058) );
  XOR U21797 ( .A(n20059), .B(n20058), .Z(n20060) );
  XOR U21798 ( .A(n20052), .B(n20053), .Z(n20055) );
  XOR U21799 ( .A(n20054), .B(n20055), .Z(n20049) );
  AND U21800 ( .A(x[494]), .B(y[7886]), .Z(n21647) );
  AND U21801 ( .A(x[488]), .B(y[7883]), .Z(n19958) );
  NANDN U21802 ( .A(n19959), .B(n19958), .Z(n19962) );
  NAND U21803 ( .A(n20239), .B(n19960), .Z(n19961) );
  NAND U21804 ( .A(n19962), .B(n19961), .Z(n20022) );
  XOR U21805 ( .A(n20023), .B(n20022), .Z(n20024) );
  AND U21806 ( .A(y[7877]), .B(x[490]), .Z(n19964) );
  NAND U21807 ( .A(y[7883]), .B(x[484]), .Z(n19963) );
  XNOR U21808 ( .A(n19964), .B(n19963), .Z(n20005) );
  AND U21809 ( .A(x[487]), .B(y[7880]), .Z(n20004) );
  XNOR U21810 ( .A(n20005), .B(n20004), .Z(n20012) );
  NAND U21811 ( .A(x[486]), .B(y[7881]), .Z(n20152) );
  XOR U21812 ( .A(n20152), .B(n20010), .Z(n20011) );
  XOR U21813 ( .A(n20012), .B(n20011), .Z(n20045) );
  AND U21814 ( .A(y[7885]), .B(x[482]), .Z(n19966) );
  NAND U21815 ( .A(y[7878]), .B(x[489]), .Z(n19965) );
  XNOR U21816 ( .A(n19966), .B(n19965), .Z(n20014) );
  AND U21817 ( .A(x[483]), .B(y[7884]), .Z(n20013) );
  XOR U21818 ( .A(n20014), .B(n20013), .Z(n20043) );
  AND U21819 ( .A(y[7886]), .B(x[481]), .Z(n19968) );
  NAND U21820 ( .A(y[7879]), .B(x[488]), .Z(n19967) );
  XNOR U21821 ( .A(n19968), .B(n19967), .Z(n19994) );
  AND U21822 ( .A(x[494]), .B(y[7873]), .Z(n20019) );
  XOR U21823 ( .A(n20019), .B(o[207]), .Z(n19993) );
  XOR U21824 ( .A(n19994), .B(n19993), .Z(n20042) );
  XOR U21825 ( .A(n20043), .B(n20042), .Z(n20044) );
  XNOR U21826 ( .A(n20024), .B(n20025), .Z(n20065) );
  XOR U21827 ( .A(n20067), .B(n20066), .Z(n20048) );
  XNOR U21828 ( .A(n20049), .B(n20048), .Z(n20051) );
  XNOR U21829 ( .A(n20050), .B(n20051), .Z(n20074) );
  NAND U21830 ( .A(n19977), .B(n19976), .Z(n19981) );
  NAND U21831 ( .A(n19979), .B(n19978), .Z(n19980) );
  AND U21832 ( .A(n19981), .B(n19980), .Z(n20073) );
  XNOR U21833 ( .A(n20074), .B(n20073), .Z(n20076) );
  XOR U21834 ( .A(n20075), .B(n20076), .Z(n20072) );
  NAND U21835 ( .A(n19983), .B(n19982), .Z(n19987) );
  NAND U21836 ( .A(n19985), .B(n19984), .Z(n19986) );
  NAND U21837 ( .A(n19987), .B(n19986), .Z(n20071) );
  XOR U21838 ( .A(n20071), .B(n20070), .Z(n19991) );
  XNOR U21839 ( .A(n20072), .B(n19991), .Z(N432) );
  AND U21840 ( .A(x[488]), .B(y[7886]), .Z(n20347) );
  NAND U21841 ( .A(n20347), .B(n19992), .Z(n19996) );
  NAND U21842 ( .A(n19994), .B(n19993), .Z(n19995) );
  NAND U21843 ( .A(n19996), .B(n19995), .Z(n20102) );
  AND U21844 ( .A(x[495]), .B(y[7887]), .Z(n21935) );
  NAND U21845 ( .A(n19997), .B(n21935), .Z(n20001) );
  NAND U21846 ( .A(n19999), .B(n19998), .Z(n20000) );
  NAND U21847 ( .A(n20001), .B(n20000), .Z(n20101) );
  XOR U21848 ( .A(n20102), .B(n20101), .Z(n20103) );
  AND U21849 ( .A(x[490]), .B(y[7883]), .Z(n20003) );
  NAND U21850 ( .A(n20003), .B(n20002), .Z(n20007) );
  NAND U21851 ( .A(n20005), .B(n20004), .Z(n20006) );
  NAND U21852 ( .A(n20007), .B(n20006), .Z(n20139) );
  AND U21853 ( .A(x[480]), .B(y[7888]), .Z(n20161) );
  NAND U21854 ( .A(x[496]), .B(y[7872]), .Z(n20162) );
  NAND U21855 ( .A(x[495]), .B(y[7873]), .Z(n20149) );
  XOR U21856 ( .A(n20164), .B(n20163), .Z(n20138) );
  NAND U21857 ( .A(y[7881]), .B(x[487]), .Z(n20008) );
  XNOR U21858 ( .A(n20009), .B(n20008), .Z(n20153) );
  NAND U21859 ( .A(x[490]), .B(y[7878]), .Z(n20154) );
  XOR U21860 ( .A(n20138), .B(n20137), .Z(n20140) );
  XNOR U21861 ( .A(n20139), .B(n20140), .Z(n20104) );
  AND U21862 ( .A(x[489]), .B(y[7885]), .Z(n20822) );
  NAND U21863 ( .A(n20822), .B(n20409), .Z(n20016) );
  NAND U21864 ( .A(n20014), .B(n20013), .Z(n20015) );
  NAND U21865 ( .A(n20016), .B(n20015), .Z(n20171) );
  AND U21866 ( .A(y[7887]), .B(x[481]), .Z(n20018) );
  NAND U21867 ( .A(y[7880]), .B(x[488]), .Z(n20017) );
  XNOR U21868 ( .A(n20018), .B(n20017), .Z(n20157) );
  NAND U21869 ( .A(n20019), .B(o[207]), .Z(n20158) );
  NAND U21870 ( .A(y[7874]), .B(x[494]), .Z(n20020) );
  XNOR U21871 ( .A(n20021), .B(n20020), .Z(n20113) );
  NAND U21872 ( .A(x[484]), .B(y[7884]), .Z(n20114) );
  XOR U21873 ( .A(n20170), .B(n20169), .Z(n20172) );
  XNOR U21874 ( .A(n20171), .B(n20172), .Z(n20131) );
  XOR U21875 ( .A(n20132), .B(n20131), .Z(n20133) );
  NAND U21876 ( .A(n20023), .B(n20022), .Z(n20027) );
  NANDN U21877 ( .A(n20025), .B(n20024), .Z(n20026) );
  AND U21878 ( .A(n20027), .B(n20026), .Z(n20095) );
  XOR U21879 ( .A(n20096), .B(n20095), .Z(n20097) );
  NAND U21880 ( .A(n20029), .B(n20028), .Z(n20033) );
  NANDN U21881 ( .A(n20031), .B(n20030), .Z(n20032) );
  NAND U21882 ( .A(n20033), .B(n20032), .Z(n20127) );
  AND U21883 ( .A(y[7876]), .B(x[493]), .Z(n20124) );
  NAND U21884 ( .A(n20664), .B(n20124), .Z(n20037) );
  NAND U21885 ( .A(n20035), .B(n20034), .Z(n20036) );
  NAND U21886 ( .A(n20037), .B(n20036), .Z(n20109) );
  AND U21887 ( .A(y[7886]), .B(x[482]), .Z(n20039) );
  NAND U21888 ( .A(y[7879]), .B(x[489]), .Z(n20038) );
  XNOR U21889 ( .A(n20039), .B(n20038), .Z(n20118) );
  NAND U21890 ( .A(x[483]), .B(y[7885]), .Z(n20119) );
  AND U21891 ( .A(x[492]), .B(y[7876]), .Z(n20833) );
  AND U21892 ( .A(y[7883]), .B(x[485]), .Z(n20041) );
  NAND U21893 ( .A(y[7875]), .B(x[493]), .Z(n20040) );
  XNOR U21894 ( .A(n20041), .B(n20040), .Z(n20144) );
  XOR U21895 ( .A(n20833), .B(n20144), .Z(n20107) );
  XOR U21896 ( .A(n20108), .B(n20107), .Z(n20110) );
  XOR U21897 ( .A(n20109), .B(n20110), .Z(n20126) );
  NAND U21898 ( .A(n20043), .B(n20042), .Z(n20047) );
  NANDN U21899 ( .A(n20045), .B(n20044), .Z(n20046) );
  AND U21900 ( .A(n20047), .B(n20046), .Z(n20125) );
  XOR U21901 ( .A(n20127), .B(n20128), .Z(n20098) );
  XNOR U21902 ( .A(n20097), .B(n20098), .Z(n20081) );
  XNOR U21903 ( .A(n20081), .B(n20080), .Z(n20083) );
  NAND U21904 ( .A(n20053), .B(n20052), .Z(n20057) );
  NAND U21905 ( .A(n20055), .B(n20054), .Z(n20056) );
  NAND U21906 ( .A(n20057), .B(n20056), .Z(n20091) );
  NAND U21907 ( .A(n20059), .B(n20058), .Z(n20063) );
  NANDN U21908 ( .A(n20061), .B(n20060), .Z(n20062) );
  NAND U21909 ( .A(n20063), .B(n20062), .Z(n20089) );
  NANDN U21910 ( .A(n20065), .B(n20064), .Z(n20069) );
  NAND U21911 ( .A(n20067), .B(n20066), .Z(n20068) );
  AND U21912 ( .A(n20069), .B(n20068), .Z(n20090) );
  XOR U21913 ( .A(n20089), .B(n20090), .Z(n20092) );
  XOR U21914 ( .A(n20091), .B(n20092), .Z(n20082) );
  XNOR U21915 ( .A(n20083), .B(n20082), .Z(n20088) );
  NAND U21916 ( .A(n20074), .B(n20073), .Z(n20078) );
  NANDN U21917 ( .A(n20076), .B(n20075), .Z(n20077) );
  NAND U21918 ( .A(n20078), .B(n20077), .Z(n20086) );
  XNOR U21919 ( .A(n20087), .B(n20086), .Z(n20079) );
  XNOR U21920 ( .A(n20088), .B(n20079), .Z(N433) );
  NANDN U21921 ( .A(n20081), .B(n20080), .Z(n20085) );
  NAND U21922 ( .A(n20083), .B(n20082), .Z(n20084) );
  AND U21923 ( .A(n20085), .B(n20084), .Z(n20183) );
  NAND U21924 ( .A(n20090), .B(n20089), .Z(n20094) );
  NAND U21925 ( .A(n20092), .B(n20091), .Z(n20093) );
  NAND U21926 ( .A(n20094), .B(n20093), .Z(n20178) );
  NAND U21927 ( .A(n20096), .B(n20095), .Z(n20100) );
  NANDN U21928 ( .A(n20098), .B(n20097), .Z(n20099) );
  NAND U21929 ( .A(n20100), .B(n20099), .Z(n20187) );
  NAND U21930 ( .A(n20102), .B(n20101), .Z(n20106) );
  NANDN U21931 ( .A(n20104), .B(n20103), .Z(n20105) );
  NAND U21932 ( .A(n20106), .B(n20105), .Z(n20269) );
  NAND U21933 ( .A(n20108), .B(n20107), .Z(n20112) );
  NAND U21934 ( .A(n20110), .B(n20109), .Z(n20111) );
  NAND U21935 ( .A(n20112), .B(n20111), .Z(n20267) );
  NAND U21936 ( .A(x[494]), .B(y[7877]), .Z(n20445) );
  NANDN U21937 ( .A(n20445), .B(n20664), .Z(n20116) );
  NANDN U21938 ( .A(n20114), .B(n20113), .Z(n20115) );
  AND U21939 ( .A(n20116), .B(n20115), .Z(n20262) );
  AND U21940 ( .A(x[489]), .B(y[7886]), .Z(n21089) );
  NANDN U21941 ( .A(n20117), .B(n21089), .Z(n20121) );
  NANDN U21942 ( .A(n20119), .B(n20118), .Z(n20120) );
  NAND U21943 ( .A(n20121), .B(n20120), .Z(n20261) );
  AND U21944 ( .A(x[487]), .B(y[7882]), .Z(n20256) );
  AND U21945 ( .A(x[485]), .B(y[7884]), .Z(n20307) );
  NAND U21946 ( .A(y[7881]), .B(x[488]), .Z(n20122) );
  XNOR U21947 ( .A(n20307), .B(n20122), .Z(n20240) );
  XOR U21948 ( .A(n20256), .B(n20255), .Z(n20258) );
  NAND U21949 ( .A(y[7885]), .B(x[484]), .Z(n20123) );
  XNOR U21950 ( .A(n20124), .B(n20123), .Z(n20202) );
  NAND U21951 ( .A(x[491]), .B(y[7878]), .Z(n20203) );
  XOR U21952 ( .A(n20258), .B(n20257), .Z(n20263) );
  XOR U21953 ( .A(n20264), .B(n20263), .Z(n20268) );
  XOR U21954 ( .A(n20267), .B(n20268), .Z(n20270) );
  XOR U21955 ( .A(n20269), .B(n20270), .Z(n20186) );
  NANDN U21956 ( .A(n20126), .B(n20125), .Z(n20130) );
  NANDN U21957 ( .A(n20128), .B(n20127), .Z(n20129) );
  NAND U21958 ( .A(n20130), .B(n20129), .Z(n20185) );
  XOR U21959 ( .A(n20187), .B(n20188), .Z(n20177) );
  NAND U21960 ( .A(n20132), .B(n20131), .Z(n20136) );
  NANDN U21961 ( .A(n20134), .B(n20133), .Z(n20135) );
  NAND U21962 ( .A(n20136), .B(n20135), .Z(n20193) );
  NAND U21963 ( .A(n20138), .B(n20137), .Z(n20142) );
  NAND U21964 ( .A(n20140), .B(n20139), .Z(n20141) );
  NAND U21965 ( .A(n20142), .B(n20141), .Z(n20275) );
  AND U21966 ( .A(x[493]), .B(y[7883]), .Z(n21108) );
  NAND U21967 ( .A(n21108), .B(n20143), .Z(n20146) );
  NAND U21968 ( .A(n20833), .B(n20144), .Z(n20145) );
  AND U21969 ( .A(n20146), .B(n20145), .Z(n20224) );
  AND U21970 ( .A(y[7888]), .B(x[481]), .Z(n20148) );
  NAND U21971 ( .A(y[7880]), .B(x[489]), .Z(n20147) );
  XNOR U21972 ( .A(n20148), .B(n20147), .Z(n20245) );
  ANDN U21973 ( .B(o[208]), .A(n20149), .Z(n20244) );
  XOR U21974 ( .A(n20245), .B(n20244), .Z(n20222) );
  AND U21975 ( .A(y[7874]), .B(x[495]), .Z(n20151) );
  NAND U21976 ( .A(y[7877]), .B(x[492]), .Z(n20150) );
  XNOR U21977 ( .A(n20151), .B(n20150), .Z(n20197) );
  NAND U21978 ( .A(x[494]), .B(y[7875]), .Z(n20198) );
  XOR U21979 ( .A(n20222), .B(n20221), .Z(n20223) );
  NANDN U21980 ( .A(n20152), .B(n20256), .Z(n20156) );
  NANDN U21981 ( .A(n20154), .B(n20153), .Z(n20155) );
  AND U21982 ( .A(n20156), .B(n20155), .Z(n20234) );
  AND U21983 ( .A(x[488]), .B(y[7887]), .Z(n20910) );
  AND U21984 ( .A(x[481]), .B(y[7880]), .Z(n20325) );
  NAND U21985 ( .A(n20910), .B(n20325), .Z(n20160) );
  NANDN U21986 ( .A(n20158), .B(n20157), .Z(n20159) );
  NAND U21987 ( .A(n20160), .B(n20159), .Z(n20233) );
  NANDN U21988 ( .A(n20162), .B(n20161), .Z(n20166) );
  NAND U21989 ( .A(n20164), .B(n20163), .Z(n20165) );
  AND U21990 ( .A(n20166), .B(n20165), .Z(n20230) );
  AND U21991 ( .A(x[480]), .B(y[7889]), .Z(n20211) );
  NAND U21992 ( .A(x[497]), .B(y[7872]), .Z(n20212) );
  NAND U21993 ( .A(x[496]), .B(y[7873]), .Z(n20208) );
  XOR U21994 ( .A(n20214), .B(n20213), .Z(n20228) );
  AND U21995 ( .A(y[7887]), .B(x[482]), .Z(n20168) );
  NAND U21996 ( .A(y[7879]), .B(x[490]), .Z(n20167) );
  XNOR U21997 ( .A(n20168), .B(n20167), .Z(n20249) );
  NAND U21998 ( .A(x[483]), .B(y[7886]), .Z(n20250) );
  XOR U21999 ( .A(n20228), .B(n20227), .Z(n20229) );
  XOR U22000 ( .A(n20236), .B(n20235), .Z(n20273) );
  XOR U22001 ( .A(n20274), .B(n20273), .Z(n20276) );
  XOR U22002 ( .A(n20275), .B(n20276), .Z(n20192) );
  NAND U22003 ( .A(n20170), .B(n20169), .Z(n20174) );
  NAND U22004 ( .A(n20172), .B(n20171), .Z(n20173) );
  AND U22005 ( .A(n20174), .B(n20173), .Z(n20191) );
  XOR U22006 ( .A(n20193), .B(n20194), .Z(n20176) );
  XOR U22007 ( .A(n20178), .B(n20179), .Z(n20184) );
  XOR U22008 ( .A(n20182), .B(n20184), .Z(n20175) );
  XOR U22009 ( .A(n20183), .B(n20175), .Z(N434) );
  NANDN U22010 ( .A(n20177), .B(n20176), .Z(n20181) );
  NAND U22011 ( .A(n20179), .B(n20178), .Z(n20180) );
  AND U22012 ( .A(n20181), .B(n20180), .Z(n20286) );
  NANDN U22013 ( .A(n20186), .B(n20185), .Z(n20190) );
  NAND U22014 ( .A(n20188), .B(n20187), .Z(n20189) );
  AND U22015 ( .A(n20190), .B(n20189), .Z(n20283) );
  NANDN U22016 ( .A(n20192), .B(n20191), .Z(n20196) );
  NANDN U22017 ( .A(n20194), .B(n20193), .Z(n20195) );
  AND U22018 ( .A(n20196), .B(n20195), .Z(n20281) );
  AND U22019 ( .A(y[7877]), .B(x[495]), .Z(n20417) );
  AND U22020 ( .A(x[492]), .B(y[7874]), .Z(n20529) );
  NAND U22021 ( .A(n20417), .B(n20529), .Z(n20200) );
  NANDN U22022 ( .A(n20198), .B(n20197), .Z(n20199) );
  AND U22023 ( .A(n20200), .B(n20199), .Z(n20374) );
  NAND U22024 ( .A(n21407), .B(n20201), .Z(n20205) );
  NANDN U22025 ( .A(n20203), .B(n20202), .Z(n20204) );
  NAND U22026 ( .A(n20205), .B(n20204), .Z(n20363) );
  AND U22027 ( .A(y[7889]), .B(x[481]), .Z(n20207) );
  NAND U22028 ( .A(y[7880]), .B(x[490]), .Z(n20206) );
  XNOR U22029 ( .A(n20207), .B(n20206), .Z(n20327) );
  ANDN U22030 ( .B(o[209]), .A(n20208), .Z(n20326) );
  XOR U22031 ( .A(n20327), .B(n20326), .Z(n20362) );
  AND U22032 ( .A(y[7875]), .B(x[495]), .Z(n20210) );
  NAND U22033 ( .A(y[7881]), .B(x[489]), .Z(n20209) );
  XNOR U22034 ( .A(n20210), .B(n20209), .Z(n20318) );
  AND U22035 ( .A(x[494]), .B(y[7876]), .Z(n20317) );
  XOR U22036 ( .A(n20318), .B(n20317), .Z(n20361) );
  XOR U22037 ( .A(n20362), .B(n20361), .Z(n20364) );
  XOR U22038 ( .A(n20363), .B(n20364), .Z(n20373) );
  NANDN U22039 ( .A(n20212), .B(n20211), .Z(n20216) );
  NAND U22040 ( .A(n20214), .B(n20213), .Z(n20215) );
  AND U22041 ( .A(n20216), .B(n20215), .Z(n20386) );
  AND U22042 ( .A(y[7874]), .B(x[496]), .Z(n20218) );
  NAND U22043 ( .A(y[7879]), .B(x[491]), .Z(n20217) );
  XNOR U22044 ( .A(n20218), .B(n20217), .Z(n20314) );
  AND U22045 ( .A(x[482]), .B(y[7888]), .Z(n20313) );
  XOR U22046 ( .A(n20314), .B(n20313), .Z(n20385) );
  AND U22047 ( .A(x[485]), .B(y[7885]), .Z(n20426) );
  NAND U22048 ( .A(y[7884]), .B(x[486]), .Z(n20219) );
  XNOR U22049 ( .A(n20426), .B(n20219), .Z(n20310) );
  NAND U22050 ( .A(y[7886]), .B(x[484]), .Z(n20220) );
  XNOR U22051 ( .A(n21094), .B(n20220), .Z(n20349) );
  AND U22052 ( .A(x[487]), .B(y[7883]), .Z(n20348) );
  XOR U22053 ( .A(n20349), .B(n20348), .Z(n20309) );
  XOR U22054 ( .A(n20310), .B(n20309), .Z(n20387) );
  XOR U22055 ( .A(n20388), .B(n20387), .Z(n20375) );
  XOR U22056 ( .A(n20376), .B(n20375), .Z(n20296) );
  NAND U22057 ( .A(n20222), .B(n20221), .Z(n20226) );
  NANDN U22058 ( .A(n20224), .B(n20223), .Z(n20225) );
  AND U22059 ( .A(n20226), .B(n20225), .Z(n20367) );
  NAND U22060 ( .A(n20228), .B(n20227), .Z(n20232) );
  NANDN U22061 ( .A(n20230), .B(n20229), .Z(n20231) );
  NAND U22062 ( .A(n20232), .B(n20231), .Z(n20368) );
  NANDN U22063 ( .A(n20234), .B(n20233), .Z(n20238) );
  NAND U22064 ( .A(n20236), .B(n20235), .Z(n20237) );
  NAND U22065 ( .A(n20238), .B(n20237), .Z(n20370) );
  AND U22066 ( .A(x[488]), .B(y[7884]), .Z(n20563) );
  NAND U22067 ( .A(n20563), .B(n20239), .Z(n20243) );
  NANDN U22068 ( .A(n20241), .B(n20240), .Z(n20242) );
  AND U22069 ( .A(n20243), .B(n20242), .Z(n20380) );
  NAND U22070 ( .A(x[489]), .B(y[7888]), .Z(n21217) );
  NANDN U22071 ( .A(n21217), .B(n20325), .Z(n20247) );
  NAND U22072 ( .A(n20245), .B(n20244), .Z(n20246) );
  NAND U22073 ( .A(n20247), .B(n20246), .Z(n20379) );
  NAND U22074 ( .A(x[490]), .B(y[7887]), .Z(n21218) );
  NANDN U22075 ( .A(n21218), .B(n20248), .Z(n20252) );
  NANDN U22076 ( .A(n20250), .B(n20249), .Z(n20251) );
  NAND U22077 ( .A(n20252), .B(n20251), .Z(n20357) );
  AND U22078 ( .A(y[7877]), .B(x[493]), .Z(n20254) );
  NAND U22079 ( .A(y[7887]), .B(x[483]), .Z(n20253) );
  XNOR U22080 ( .A(n20254), .B(n20253), .Z(n20338) );
  NAND U22081 ( .A(x[492]), .B(y[7878]), .Z(n20339) );
  AND U22082 ( .A(x[480]), .B(y[7890]), .Z(n20330) );
  NAND U22083 ( .A(x[498]), .B(y[7872]), .Z(n20331) );
  NAND U22084 ( .A(x[497]), .B(y[7873]), .Z(n20352) );
  XOR U22085 ( .A(n20333), .B(n20332), .Z(n20355) );
  XOR U22086 ( .A(n20356), .B(n20355), .Z(n20358) );
  XOR U22087 ( .A(n20357), .B(n20358), .Z(n20381) );
  XOR U22088 ( .A(n20382), .B(n20381), .Z(n20302) );
  NAND U22089 ( .A(n20256), .B(n20255), .Z(n20260) );
  NAND U22090 ( .A(n20258), .B(n20257), .Z(n20259) );
  AND U22091 ( .A(n20260), .B(n20259), .Z(n20301) );
  NANDN U22092 ( .A(n20262), .B(n20261), .Z(n20266) );
  NAND U22093 ( .A(n20264), .B(n20263), .Z(n20265) );
  AND U22094 ( .A(n20266), .B(n20265), .Z(n20303) );
  XOR U22095 ( .A(n20304), .B(n20303), .Z(n20297) );
  XOR U22096 ( .A(n20298), .B(n20297), .Z(n20292) );
  NAND U22097 ( .A(n20268), .B(n20267), .Z(n20272) );
  NAND U22098 ( .A(n20270), .B(n20269), .Z(n20271) );
  NAND U22099 ( .A(n20272), .B(n20271), .Z(n20290) );
  NAND U22100 ( .A(n20274), .B(n20273), .Z(n20278) );
  NAND U22101 ( .A(n20276), .B(n20275), .Z(n20277) );
  NAND U22102 ( .A(n20278), .B(n20277), .Z(n20289) );
  XOR U22103 ( .A(n20290), .B(n20289), .Z(n20291) );
  XOR U22104 ( .A(n20281), .B(n20280), .Z(n20282) );
  XOR U22105 ( .A(n20283), .B(n20282), .Z(n20288) );
  XNOR U22106 ( .A(n20287), .B(n20288), .Z(n20279) );
  XOR U22107 ( .A(n20286), .B(n20279), .Z(N435) );
  NAND U22108 ( .A(n20281), .B(n20280), .Z(n20285) );
  NAND U22109 ( .A(n20283), .B(n20282), .Z(n20284) );
  AND U22110 ( .A(n20285), .B(n20284), .Z(n20501) );
  NAND U22111 ( .A(n20290), .B(n20289), .Z(n20294) );
  NANDN U22112 ( .A(n20292), .B(n20291), .Z(n20293) );
  NAND U22113 ( .A(n20294), .B(n20293), .Z(n20506) );
  NANDN U22114 ( .A(n20296), .B(n20295), .Z(n20300) );
  NAND U22115 ( .A(n20298), .B(n20297), .Z(n20299) );
  AND U22116 ( .A(n20300), .B(n20299), .Z(n20504) );
  NANDN U22117 ( .A(n20302), .B(n20301), .Z(n20306) );
  NAND U22118 ( .A(n20304), .B(n20303), .Z(n20305) );
  NAND U22119 ( .A(n20306), .B(n20305), .Z(n20485) );
  AND U22120 ( .A(x[486]), .B(y[7885]), .Z(n20308) );
  NAND U22121 ( .A(n20308), .B(n20307), .Z(n20312) );
  NAND U22122 ( .A(n20310), .B(n20309), .Z(n20311) );
  NAND U22123 ( .A(n20312), .B(n20311), .Z(n20479) );
  AND U22124 ( .A(x[496]), .B(y[7879]), .Z(n20826) );
  NAND U22125 ( .A(n20826), .B(n20664), .Z(n20316) );
  NAND U22126 ( .A(n20314), .B(n20313), .Z(n20315) );
  NAND U22127 ( .A(n20316), .B(n20315), .Z(n20477) );
  AND U22128 ( .A(x[495]), .B(y[7881]), .Z(n21121) );
  NAND U22129 ( .A(n21121), .B(n20404), .Z(n20320) );
  NAND U22130 ( .A(n20318), .B(n20317), .Z(n20319) );
  AND U22131 ( .A(n20320), .B(n20319), .Z(n20395) );
  AND U22132 ( .A(y[7890]), .B(x[481]), .Z(n20322) );
  NAND U22133 ( .A(y[7883]), .B(x[488]), .Z(n20321) );
  XNOR U22134 ( .A(n20322), .B(n20321), .Z(n20444) );
  AND U22135 ( .A(y[7878]), .B(x[493]), .Z(n20324) );
  NAND U22136 ( .A(y[7889]), .B(x[482]), .Z(n20323) );
  XNOR U22137 ( .A(n20324), .B(n20323), .Z(n20410) );
  XOR U22138 ( .A(n20393), .B(n20392), .Z(n20394) );
  XOR U22139 ( .A(n20477), .B(n20478), .Z(n20480) );
  XOR U22140 ( .A(n20479), .B(n20480), .Z(n20484) );
  NAND U22141 ( .A(x[490]), .B(y[7889]), .Z(n21496) );
  NANDN U22142 ( .A(n21496), .B(n20325), .Z(n20329) );
  NAND U22143 ( .A(n20327), .B(n20326), .Z(n20328) );
  AND U22144 ( .A(n20329), .B(n20328), .Z(n20456) );
  NANDN U22145 ( .A(n20331), .B(n20330), .Z(n20335) );
  NAND U22146 ( .A(n20333), .B(n20332), .Z(n20334) );
  AND U22147 ( .A(n20335), .B(n20334), .Z(n20454) );
  AND U22148 ( .A(y[7875]), .B(x[496]), .Z(n21054) );
  NAND U22149 ( .A(y[7882]), .B(x[489]), .Z(n20336) );
  XNOR U22150 ( .A(n21054), .B(n20336), .Z(n20405) );
  NAND U22151 ( .A(x[495]), .B(y[7876]), .Z(n20406) );
  AND U22152 ( .A(x[493]), .B(y[7887]), .Z(n21668) );
  NANDN U22153 ( .A(n20337), .B(n21668), .Z(n20341) );
  NANDN U22154 ( .A(n20339), .B(n20338), .Z(n20340) );
  AND U22155 ( .A(n20341), .B(n20340), .Z(n20462) );
  AND U22156 ( .A(y[7881]), .B(x[490]), .Z(n20343) );
  NAND U22157 ( .A(y[7874]), .B(x[497]), .Z(n20342) );
  XNOR U22158 ( .A(n20343), .B(n20342), .Z(n20450) );
  NAND U22159 ( .A(x[498]), .B(y[7873]), .Z(n20425) );
  XOR U22160 ( .A(n20450), .B(n20449), .Z(n20460) );
  NAND U22161 ( .A(y[7888]), .B(x[483]), .Z(n20344) );
  XNOR U22162 ( .A(n20345), .B(n20344), .Z(n20419) );
  XOR U22163 ( .A(n20460), .B(n20459), .Z(n20461) );
  NAND U22164 ( .A(n20347), .B(n20346), .Z(n20351) );
  NAND U22165 ( .A(n20349), .B(n20348), .Z(n20350) );
  AND U22166 ( .A(n20351), .B(n20350), .Z(n20401) );
  AND U22167 ( .A(x[480]), .B(y[7891]), .Z(n20430) );
  NAND U22168 ( .A(x[499]), .B(y[7872]), .Z(n20431) );
  ANDN U22169 ( .B(o[210]), .A(n20352), .Z(n20432) );
  XOR U22170 ( .A(n20433), .B(n20432), .Z(n20399) );
  AND U22171 ( .A(x[484]), .B(y[7887]), .Z(n20577) );
  AND U22172 ( .A(y[7886]), .B(x[485]), .Z(n20354) );
  NAND U22173 ( .A(y[7885]), .B(x[486]), .Z(n20353) );
  XOR U22174 ( .A(n20354), .B(n20353), .Z(n20427) );
  XOR U22175 ( .A(n20399), .B(n20398), .Z(n20400) );
  XOR U22176 ( .A(n20401), .B(n20400), .Z(n20471) );
  NAND U22177 ( .A(n20356), .B(n20355), .Z(n20360) );
  NAND U22178 ( .A(n20358), .B(n20357), .Z(n20359) );
  NAND U22179 ( .A(n20360), .B(n20359), .Z(n20466) );
  NAND U22180 ( .A(n20362), .B(n20361), .Z(n20366) );
  NAND U22181 ( .A(n20364), .B(n20363), .Z(n20365) );
  NAND U22182 ( .A(n20366), .B(n20365), .Z(n20465) );
  XOR U22183 ( .A(n20466), .B(n20465), .Z(n20467) );
  XNOR U22184 ( .A(n20468), .B(n20467), .Z(n20483) );
  XOR U22185 ( .A(n20485), .B(n20486), .Z(n20497) );
  NANDN U22186 ( .A(n20368), .B(n20367), .Z(n20372) );
  NANDN U22187 ( .A(n20370), .B(n20369), .Z(n20371) );
  AND U22188 ( .A(n20372), .B(n20371), .Z(n20496) );
  NANDN U22189 ( .A(n20374), .B(n20373), .Z(n20378) );
  NAND U22190 ( .A(n20376), .B(n20375), .Z(n20377) );
  AND U22191 ( .A(n20378), .B(n20377), .Z(n20492) );
  NANDN U22192 ( .A(n20380), .B(n20379), .Z(n20384) );
  NAND U22193 ( .A(n20382), .B(n20381), .Z(n20383) );
  AND U22194 ( .A(n20384), .B(n20383), .Z(n20490) );
  NANDN U22195 ( .A(n20386), .B(n20385), .Z(n20390) );
  NAND U22196 ( .A(n20388), .B(n20387), .Z(n20389) );
  NAND U22197 ( .A(n20390), .B(n20389), .Z(n20489) );
  XOR U22198 ( .A(n20496), .B(n20495), .Z(n20498) );
  XNOR U22199 ( .A(n20497), .B(n20498), .Z(n20505) );
  XOR U22200 ( .A(n20506), .B(n20507), .Z(n20503) );
  XNOR U22201 ( .A(n20502), .B(n20503), .Z(n20391) );
  XOR U22202 ( .A(n20501), .B(n20391), .Z(N436) );
  NAND U22203 ( .A(n20393), .B(n20392), .Z(n20397) );
  NANDN U22204 ( .A(n20395), .B(n20394), .Z(n20396) );
  AND U22205 ( .A(n20397), .B(n20396), .Z(n20512) );
  NAND U22206 ( .A(n20399), .B(n20398), .Z(n20403) );
  NANDN U22207 ( .A(n20401), .B(n20400), .Z(n20402) );
  NAND U22208 ( .A(n20403), .B(n20402), .Z(n20511) );
  AND U22209 ( .A(x[496]), .B(y[7882]), .Z(n21335) );
  NAND U22210 ( .A(n21335), .B(n20404), .Z(n20408) );
  NANDN U22211 ( .A(n20406), .B(n20405), .Z(n20407) );
  AND U22212 ( .A(n20408), .B(n20407), .Z(n20552) );
  AND U22213 ( .A(x[493]), .B(y[7889]), .Z(n21876) );
  NAND U22214 ( .A(n21876), .B(n20409), .Z(n20413) );
  NANDN U22215 ( .A(n20411), .B(n20410), .Z(n20412) );
  AND U22216 ( .A(n20413), .B(n20412), .Z(n20597) );
  AND U22217 ( .A(y[7876]), .B(x[496]), .Z(n20415) );
  NAND U22218 ( .A(y[7882]), .B(x[490]), .Z(n20414) );
  XNOR U22219 ( .A(n20415), .B(n20414), .Z(n20558) );
  NAND U22220 ( .A(x[482]), .B(y[7890]), .Z(n20559) );
  NAND U22221 ( .A(y[7883]), .B(x[489]), .Z(n20416) );
  XNOR U22222 ( .A(n20417), .B(n20416), .Z(n20540) );
  NAND U22223 ( .A(x[494]), .B(y[7878]), .Z(n20541) );
  XOR U22224 ( .A(n20595), .B(n20594), .Z(n20596) );
  NAND U22225 ( .A(x[491]), .B(y[7888]), .Z(n21497) );
  NANDN U22226 ( .A(n21497), .B(n20418), .Z(n20422) );
  NANDN U22227 ( .A(n20420), .B(n20419), .Z(n20421) );
  AND U22228 ( .A(n20422), .B(n20421), .Z(n20603) );
  AND U22229 ( .A(y[7881]), .B(x[491]), .Z(n20424) );
  NAND U22230 ( .A(y[7891]), .B(x[481]), .Z(n20423) );
  XNOR U22231 ( .A(n20424), .B(n20423), .Z(n20536) );
  NAND U22232 ( .A(x[499]), .B(y[7873]), .Z(n20544) );
  XOR U22233 ( .A(n20536), .B(n20535), .Z(n20601) );
  AND U22234 ( .A(x[480]), .B(y[7892]), .Z(n20582) );
  NAND U22235 ( .A(x[500]), .B(y[7872]), .Z(n20583) );
  ANDN U22236 ( .B(o[211]), .A(n20425), .Z(n20584) );
  XOR U22237 ( .A(n20585), .B(n20584), .Z(n20600) );
  XOR U22238 ( .A(n20601), .B(n20600), .Z(n20602) );
  XOR U22239 ( .A(n20554), .B(n20553), .Z(n20513) );
  XOR U22240 ( .A(n20514), .B(n20513), .Z(n20609) );
  AND U22241 ( .A(x[486]), .B(y[7886]), .Z(n20546) );
  IV U22242 ( .A(n20546), .Z(n20442) );
  NANDN U22243 ( .A(n20442), .B(n20426), .Z(n20429) );
  NANDN U22244 ( .A(n20427), .B(n20577), .Z(n20428) );
  AND U22245 ( .A(n20429), .B(n20428), .Z(n20526) );
  NANDN U22246 ( .A(n20431), .B(n20430), .Z(n20435) );
  NAND U22247 ( .A(n20433), .B(n20432), .Z(n20434) );
  AND U22248 ( .A(n20435), .B(n20434), .Z(n20524) );
  AND U22249 ( .A(y[7874]), .B(x[498]), .Z(n20437) );
  NAND U22250 ( .A(y[7880]), .B(x[492]), .Z(n20436) );
  XNOR U22251 ( .A(n20437), .B(n20436), .Z(n20530) );
  NAND U22252 ( .A(x[497]), .B(y[7875]), .Z(n20531) );
  AND U22253 ( .A(y[7879]), .B(x[493]), .Z(n20439) );
  NAND U22254 ( .A(y[7889]), .B(x[483]), .Z(n20438) );
  XNOR U22255 ( .A(n20439), .B(n20438), .Z(n20564) );
  XOR U22256 ( .A(n20564), .B(n20563), .Z(n20548) );
  AND U22257 ( .A(y[7887]), .B(x[485]), .Z(n20441) );
  NAND U22258 ( .A(y[7888]), .B(x[484]), .Z(n20440) );
  XNOR U22259 ( .A(n20441), .B(n20440), .Z(n20579) );
  AND U22260 ( .A(x[487]), .B(y[7885]), .Z(n20578) );
  XNOR U22261 ( .A(n20579), .B(n20578), .Z(n20545) );
  XOR U22262 ( .A(n20442), .B(n20545), .Z(n20547) );
  AND U22263 ( .A(x[488]), .B(y[7890]), .Z(n21631) );
  NAND U22264 ( .A(n21631), .B(n20443), .Z(n20447) );
  NANDN U22265 ( .A(n20445), .B(n20444), .Z(n20446) );
  AND U22266 ( .A(n20447), .B(n20446), .Z(n20589) );
  AND U22267 ( .A(x[497]), .B(y[7881]), .Z(n21289) );
  IV U22268 ( .A(n21289), .Z(n21344) );
  NANDN U22269 ( .A(n21344), .B(n20448), .Z(n20452) );
  NAND U22270 ( .A(n20450), .B(n20449), .Z(n20451) );
  NAND U22271 ( .A(n20452), .B(n20451), .Z(n20588) );
  XNOR U22272 ( .A(n20590), .B(n20591), .Z(n20517) );
  XOR U22273 ( .A(n20518), .B(n20517), .Z(n20519) );
  NANDN U22274 ( .A(n20454), .B(n20453), .Z(n20458) );
  NANDN U22275 ( .A(n20456), .B(n20455), .Z(n20457) );
  NAND U22276 ( .A(n20458), .B(n20457), .Z(n20520) );
  NAND U22277 ( .A(n20460), .B(n20459), .Z(n20464) );
  NANDN U22278 ( .A(n20462), .B(n20461), .Z(n20463) );
  NAND U22279 ( .A(n20464), .B(n20463), .Z(n20607) );
  NAND U22280 ( .A(n20466), .B(n20465), .Z(n20470) );
  NAND U22281 ( .A(n20468), .B(n20467), .Z(n20469) );
  AND U22282 ( .A(n20470), .B(n20469), .Z(n20621) );
  NANDN U22283 ( .A(n20472), .B(n20471), .Z(n20476) );
  NANDN U22284 ( .A(n20474), .B(n20473), .Z(n20475) );
  NAND U22285 ( .A(n20476), .B(n20475), .Z(n20618) );
  NAND U22286 ( .A(n20478), .B(n20477), .Z(n20482) );
  NAND U22287 ( .A(n20480), .B(n20479), .Z(n20481) );
  AND U22288 ( .A(n20482), .B(n20481), .Z(n20619) );
  XOR U22289 ( .A(n20618), .B(n20619), .Z(n20620) );
  XNOR U22290 ( .A(n20621), .B(n20620), .Z(n20612) );
  NANDN U22291 ( .A(n20484), .B(n20483), .Z(n20488) );
  NANDN U22292 ( .A(n20486), .B(n20485), .Z(n20487) );
  AND U22293 ( .A(n20488), .B(n20487), .Z(n20614) );
  XOR U22294 ( .A(n20615), .B(n20614), .Z(n20627) );
  NANDN U22295 ( .A(n20490), .B(n20489), .Z(n20494) );
  NANDN U22296 ( .A(n20492), .B(n20491), .Z(n20493) );
  AND U22297 ( .A(n20494), .B(n20493), .Z(n20624) );
  NAND U22298 ( .A(n20496), .B(n20495), .Z(n20500) );
  NAND U22299 ( .A(n20498), .B(n20497), .Z(n20499) );
  NAND U22300 ( .A(n20500), .B(n20499), .Z(n20625) );
  XOR U22301 ( .A(n20627), .B(n20626), .Z(n20632) );
  NANDN U22302 ( .A(n20505), .B(n20504), .Z(n20509) );
  NAND U22303 ( .A(n20507), .B(n20506), .Z(n20508) );
  AND U22304 ( .A(n20509), .B(n20508), .Z(n20630) );
  XOR U22305 ( .A(n20631), .B(n20630), .Z(n20510) );
  XNOR U22306 ( .A(n20632), .B(n20510), .Z(N437) );
  NANDN U22307 ( .A(n20512), .B(n20511), .Z(n20516) );
  NAND U22308 ( .A(n20514), .B(n20513), .Z(n20515) );
  AND U22309 ( .A(n20516), .B(n20515), .Z(n20643) );
  NAND U22310 ( .A(n20518), .B(n20517), .Z(n20522) );
  NANDN U22311 ( .A(n20520), .B(n20519), .Z(n20521) );
  AND U22312 ( .A(n20522), .B(n20521), .Z(n20641) );
  NANDN U22313 ( .A(n20524), .B(n20523), .Z(n20528) );
  NANDN U22314 ( .A(n20526), .B(n20525), .Z(n20527) );
  AND U22315 ( .A(n20528), .B(n20527), .Z(n20734) );
  AND U22316 ( .A(x[498]), .B(y[7880]), .Z(n21342) );
  NAND U22317 ( .A(n21342), .B(n20529), .Z(n20533) );
  NANDN U22318 ( .A(n20531), .B(n20530), .Z(n20532) );
  AND U22319 ( .A(n20533), .B(n20532), .Z(n20714) );
  AND U22320 ( .A(x[491]), .B(y[7891]), .Z(n21941) );
  AND U22321 ( .A(x[481]), .B(y[7881]), .Z(n20534) );
  NAND U22322 ( .A(n21941), .B(n20534), .Z(n20538) );
  NAND U22323 ( .A(n20536), .B(n20535), .Z(n20537) );
  NAND U22324 ( .A(n20538), .B(n20537), .Z(n20713) );
  AND U22325 ( .A(x[495]), .B(y[7883]), .Z(n21332) );
  NAND U22326 ( .A(n21332), .B(n20539), .Z(n20543) );
  NANDN U22327 ( .A(n20541), .B(n20540), .Z(n20542) );
  AND U22328 ( .A(n20543), .B(n20542), .Z(n20678) );
  AND U22329 ( .A(x[480]), .B(y[7893]), .Z(n20697) );
  NAND U22330 ( .A(x[501]), .B(y[7872]), .Z(n20698) );
  ANDN U22331 ( .B(o[212]), .A(n20544), .Z(n20699) );
  XOR U22332 ( .A(n20700), .B(n20699), .Z(n20676) );
  AND U22333 ( .A(x[485]), .B(y[7888]), .Z(n20684) );
  AND U22334 ( .A(x[496]), .B(y[7877]), .Z(n20683) );
  XOR U22335 ( .A(n20684), .B(n20683), .Z(n20682) );
  AND U22336 ( .A(x[495]), .B(y[7878]), .Z(n20681) );
  XOR U22337 ( .A(n20682), .B(n20681), .Z(n20675) );
  XOR U22338 ( .A(n20676), .B(n20675), .Z(n20677) );
  XOR U22339 ( .A(n20716), .B(n20715), .Z(n20731) );
  NANDN U22340 ( .A(n20546), .B(n20545), .Z(n20550) );
  NANDN U22341 ( .A(n20548), .B(n20547), .Z(n20549) );
  NAND U22342 ( .A(n20550), .B(n20549), .Z(n20732) );
  XOR U22343 ( .A(n20641), .B(n20640), .Z(n20642) );
  NANDN U22344 ( .A(n20552), .B(n20551), .Z(n20556) );
  NAND U22345 ( .A(n20554), .B(n20553), .Z(n20555) );
  AND U22346 ( .A(n20556), .B(n20555), .Z(n20740) );
  NAND U22347 ( .A(n21335), .B(n20557), .Z(n20561) );
  NANDN U22348 ( .A(n20559), .B(n20558), .Z(n20560) );
  AND U22349 ( .A(n20561), .B(n20560), .Z(n20647) );
  NAND U22350 ( .A(n20562), .B(n21876), .Z(n20566) );
  NAND U22351 ( .A(n20564), .B(n20563), .Z(n20565) );
  AND U22352 ( .A(n20566), .B(n20565), .Z(n20728) );
  AND U22353 ( .A(y[7874]), .B(x[499]), .Z(n20568) );
  NAND U22354 ( .A(y[7882]), .B(x[491]), .Z(n20567) );
  XNOR U22355 ( .A(n20568), .B(n20567), .Z(n20666) );
  AND U22356 ( .A(x[500]), .B(y[7873]), .Z(n20696) );
  XOR U22357 ( .A(o[213]), .B(n20696), .Z(n20665) );
  XOR U22358 ( .A(n20666), .B(n20665), .Z(n20726) );
  AND U22359 ( .A(y[7875]), .B(x[498]), .Z(n20570) );
  NAND U22360 ( .A(y[7883]), .B(x[490]), .Z(n20569) );
  XNOR U22361 ( .A(n20570), .B(n20569), .Z(n20704) );
  NAND U22362 ( .A(x[481]), .B(y[7892]), .Z(n20705) );
  XOR U22363 ( .A(n20726), .B(n20725), .Z(n20727) );
  AND U22364 ( .A(x[487]), .B(y[7886]), .Z(n20909) );
  AND U22365 ( .A(y[7887]), .B(x[486]), .Z(n20572) );
  NAND U22366 ( .A(y[7879]), .B(x[494]), .Z(n20571) );
  XNOR U22367 ( .A(n20572), .B(n20571), .Z(n20708) );
  XOR U22368 ( .A(n20909), .B(n20708), .Z(n20655) );
  AND U22369 ( .A(x[489]), .B(y[7884]), .Z(n20653) );
  NAND U22370 ( .A(x[488]), .B(y[7885]), .Z(n20652) );
  AND U22371 ( .A(y[7880]), .B(x[493]), .Z(n20574) );
  NAND U22372 ( .A(y[7890]), .B(x[483]), .Z(n20573) );
  XNOR U22373 ( .A(n20574), .B(n20573), .Z(n20692) );
  NAND U22374 ( .A(x[484]), .B(y[7889]), .Z(n20693) );
  AND U22375 ( .A(y[7881]), .B(x[492]), .Z(n20576) );
  NAND U22376 ( .A(y[7876]), .B(x[497]), .Z(n20575) );
  XNOR U22377 ( .A(n20576), .B(n20575), .Z(n20658) );
  NAND U22378 ( .A(x[482]), .B(y[7891]), .Z(n20659) );
  XOR U22379 ( .A(n20670), .B(n20669), .Z(n20672) );
  XOR U22380 ( .A(n20671), .B(n20672), .Z(n20722) );
  NAND U22381 ( .A(n20684), .B(n20577), .Z(n20581) );
  NAND U22382 ( .A(n20579), .B(n20578), .Z(n20580) );
  AND U22383 ( .A(n20581), .B(n20580), .Z(n20720) );
  NANDN U22384 ( .A(n20583), .B(n20582), .Z(n20587) );
  NAND U22385 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U22386 ( .A(n20587), .B(n20586), .Z(n20719) );
  XOR U22387 ( .A(n20722), .B(n20721), .Z(n20648) );
  XOR U22388 ( .A(n20649), .B(n20648), .Z(n20738) );
  NANDN U22389 ( .A(n20589), .B(n20588), .Z(n20593) );
  NAND U22390 ( .A(n20591), .B(n20590), .Z(n20592) );
  NAND U22391 ( .A(n20593), .B(n20592), .Z(n20745) );
  NAND U22392 ( .A(n20595), .B(n20594), .Z(n20599) );
  NANDN U22393 ( .A(n20597), .B(n20596), .Z(n20598) );
  NAND U22394 ( .A(n20599), .B(n20598), .Z(n20744) );
  NAND U22395 ( .A(n20601), .B(n20600), .Z(n20605) );
  NANDN U22396 ( .A(n20603), .B(n20602), .Z(n20604) );
  NAND U22397 ( .A(n20605), .B(n20604), .Z(n20743) );
  XOR U22398 ( .A(n20744), .B(n20743), .Z(n20746) );
  XOR U22399 ( .A(n20745), .B(n20746), .Z(n20737) );
  XOR U22400 ( .A(n20738), .B(n20737), .Z(n20739) );
  NANDN U22401 ( .A(n20607), .B(n20606), .Z(n20611) );
  NANDN U22402 ( .A(n20609), .B(n20608), .Z(n20610) );
  NAND U22403 ( .A(n20611), .B(n20610), .Z(n20634) );
  XOR U22404 ( .A(n20635), .B(n20634), .Z(n20637) );
  XOR U22405 ( .A(n20636), .B(n20637), .Z(n20755) );
  NANDN U22406 ( .A(n20613), .B(n20612), .Z(n20617) );
  NAND U22407 ( .A(n20615), .B(n20614), .Z(n20616) );
  NAND U22408 ( .A(n20617), .B(n20616), .Z(n20752) );
  NAND U22409 ( .A(n20619), .B(n20618), .Z(n20623) );
  NAND U22410 ( .A(n20621), .B(n20620), .Z(n20622) );
  AND U22411 ( .A(n20623), .B(n20622), .Z(n20753) );
  XOR U22412 ( .A(n20752), .B(n20753), .Z(n20754) );
  NANDN U22413 ( .A(n20625), .B(n20624), .Z(n20629) );
  NANDN U22414 ( .A(n20627), .B(n20626), .Z(n20628) );
  NAND U22415 ( .A(n20629), .B(n20628), .Z(n20749) );
  XOR U22416 ( .A(n20749), .B(n20750), .Z(n20633) );
  XNOR U22417 ( .A(n20751), .B(n20633), .Z(N438) );
  NAND U22418 ( .A(n20635), .B(n20634), .Z(n20639) );
  NAND U22419 ( .A(n20637), .B(n20636), .Z(n20638) );
  AND U22420 ( .A(n20639), .B(n20638), .Z(n20882) );
  NAND U22421 ( .A(n20641), .B(n20640), .Z(n20645) );
  NANDN U22422 ( .A(n20643), .B(n20642), .Z(n20644) );
  AND U22423 ( .A(n20645), .B(n20644), .Z(n20880) );
  NANDN U22424 ( .A(n20647), .B(n20646), .Z(n20651) );
  NAND U22425 ( .A(n20649), .B(n20648), .Z(n20650) );
  NAND U22426 ( .A(n20651), .B(n20650), .Z(n20875) );
  NANDN U22427 ( .A(n20653), .B(n20652), .Z(n20657) );
  NANDN U22428 ( .A(n20655), .B(n20654), .Z(n20656) );
  AND U22429 ( .A(n20657), .B(n20656), .Z(n20870) );
  NANDN U22430 ( .A(n21344), .B(n20833), .Z(n20661) );
  NANDN U22431 ( .A(n20659), .B(n20658), .Z(n20660) );
  NAND U22432 ( .A(n20661), .B(n20660), .Z(n20797) );
  AND U22433 ( .A(x[485]), .B(y[7889]), .Z(n20843) );
  AND U22434 ( .A(x[497]), .B(y[7877]), .Z(n20844) );
  XOR U22435 ( .A(n20843), .B(n20844), .Z(n20845) );
  AND U22436 ( .A(x[496]), .B(y[7878]), .Z(n20846) );
  XOR U22437 ( .A(n20845), .B(n20846), .Z(n20796) );
  AND U22438 ( .A(y[7876]), .B(x[498]), .Z(n20663) );
  NAND U22439 ( .A(y[7882]), .B(x[492]), .Z(n20662) );
  XNOR U22440 ( .A(n20663), .B(n20662), .Z(n20834) );
  AND U22441 ( .A(x[484]), .B(y[7890]), .Z(n20835) );
  XOR U22442 ( .A(n20834), .B(n20835), .Z(n20795) );
  XOR U22443 ( .A(n20796), .B(n20795), .Z(n20798) );
  XNOR U22444 ( .A(n20797), .B(n20798), .Z(n20867) );
  AND U22445 ( .A(x[499]), .B(y[7882]), .Z(n21775) );
  NAND U22446 ( .A(n21775), .B(n20664), .Z(n20668) );
  NAND U22447 ( .A(n20666), .B(n20665), .Z(n20667) );
  AND U22448 ( .A(n20668), .B(n20667), .Z(n20868) );
  XOR U22449 ( .A(n20867), .B(n20868), .Z(n20869) );
  NAND U22450 ( .A(n20670), .B(n20669), .Z(n20674) );
  NAND U22451 ( .A(n20672), .B(n20671), .Z(n20673) );
  AND U22452 ( .A(n20674), .B(n20673), .Z(n20856) );
  NAND U22453 ( .A(n20676), .B(n20675), .Z(n20680) );
  NANDN U22454 ( .A(n20678), .B(n20677), .Z(n20679) );
  NAND U22455 ( .A(n20680), .B(n20679), .Z(n20855) );
  AND U22456 ( .A(n20682), .B(n20681), .Z(n20686) );
  NAND U22457 ( .A(n20684), .B(n20683), .Z(n20685) );
  NANDN U22458 ( .A(n20686), .B(n20685), .Z(n20818) );
  AND U22459 ( .A(y[7881]), .B(x[493]), .Z(n20688) );
  NAND U22460 ( .A(y[7874]), .B(x[500]), .Z(n20687) );
  XNOR U22461 ( .A(n20688), .B(n20687), .Z(n20839) );
  AND U22462 ( .A(x[482]), .B(y[7892]), .Z(n20840) );
  XOR U22463 ( .A(n20839), .B(n20840), .Z(n20816) );
  AND U22464 ( .A(y[7888]), .B(x[486]), .Z(n20690) );
  NAND U22465 ( .A(y[7879]), .B(x[495]), .Z(n20689) );
  XNOR U22466 ( .A(n20690), .B(n20689), .Z(n20851) );
  XOR U22467 ( .A(n20816), .B(n20815), .Z(n20817) );
  XOR U22468 ( .A(n20818), .B(n20817), .Z(n20862) );
  AND U22469 ( .A(x[493]), .B(y[7890]), .Z(n21959) );
  NANDN U22470 ( .A(n20691), .B(n21959), .Z(n20695) );
  NANDN U22471 ( .A(n20693), .B(n20692), .Z(n20694) );
  AND U22472 ( .A(n20695), .B(n20694), .Z(n20786) );
  AND U22473 ( .A(x[481]), .B(y[7893]), .Z(n20809) );
  XOR U22474 ( .A(n20810), .B(n20809), .Z(n20808) );
  AND U22475 ( .A(o[213]), .B(n20696), .Z(n20807) );
  XOR U22476 ( .A(n20808), .B(n20807), .Z(n20784) );
  AND U22477 ( .A(x[494]), .B(y[7880]), .Z(n20801) );
  AND U22478 ( .A(x[483]), .B(y[7891]), .Z(n20802) );
  XOR U22479 ( .A(n20801), .B(n20802), .Z(n20803) );
  AND U22480 ( .A(x[499]), .B(y[7875]), .Z(n20804) );
  XOR U22481 ( .A(n20803), .B(n20804), .Z(n20783) );
  XOR U22482 ( .A(n20784), .B(n20783), .Z(n20785) );
  XOR U22483 ( .A(n20862), .B(n20861), .Z(n20864) );
  NANDN U22484 ( .A(n20698), .B(n20697), .Z(n20702) );
  NAND U22485 ( .A(n20700), .B(n20699), .Z(n20701) );
  AND U22486 ( .A(n20702), .B(n20701), .Z(n20778) );
  AND U22487 ( .A(x[498]), .B(y[7883]), .Z(n21777) );
  NAND U22488 ( .A(n21777), .B(n20703), .Z(n20707) );
  NANDN U22489 ( .A(n20705), .B(n20704), .Z(n20706) );
  NAND U22490 ( .A(n20707), .B(n20706), .Z(n20777) );
  AND U22491 ( .A(x[494]), .B(y[7887]), .Z(n21787) );
  NAND U22492 ( .A(n20850), .B(n21787), .Z(n20710) );
  NAND U22493 ( .A(n20909), .B(n20708), .Z(n20709) );
  AND U22494 ( .A(n20710), .B(n20709), .Z(n20792) );
  AND U22495 ( .A(x[480]), .B(y[7894]), .Z(n20827) );
  AND U22496 ( .A(x[502]), .B(y[7872]), .Z(n20828) );
  XOR U22497 ( .A(n20827), .B(n20828), .Z(n20830) );
  AND U22498 ( .A(x[501]), .B(y[7873]), .Z(n20849) );
  XOR U22499 ( .A(o[214]), .B(n20849), .Z(n20829) );
  XOR U22500 ( .A(n20830), .B(n20829), .Z(n20790) );
  AND U22501 ( .A(y[7887]), .B(x[487]), .Z(n20712) );
  NAND U22502 ( .A(y[7886]), .B(x[488]), .Z(n20711) );
  XNOR U22503 ( .A(n20712), .B(n20711), .Z(n20821) );
  XOR U22504 ( .A(n20821), .B(n20822), .Z(n20789) );
  XOR U22505 ( .A(n20790), .B(n20789), .Z(n20791) );
  XOR U22506 ( .A(n20780), .B(n20779), .Z(n20863) );
  XOR U22507 ( .A(n20864), .B(n20863), .Z(n20857) );
  XOR U22508 ( .A(n20858), .B(n20857), .Z(n20873) );
  XOR U22509 ( .A(n20875), .B(n20876), .Z(n20768) );
  NANDN U22510 ( .A(n20714), .B(n20713), .Z(n20718) );
  NAND U22511 ( .A(n20716), .B(n20715), .Z(n20717) );
  AND U22512 ( .A(n20718), .B(n20717), .Z(n20774) );
  NANDN U22513 ( .A(n20720), .B(n20719), .Z(n20724) );
  NAND U22514 ( .A(n20722), .B(n20721), .Z(n20723) );
  AND U22515 ( .A(n20724), .B(n20723), .Z(n20772) );
  NAND U22516 ( .A(n20726), .B(n20725), .Z(n20730) );
  NANDN U22517 ( .A(n20728), .B(n20727), .Z(n20729) );
  NAND U22518 ( .A(n20730), .B(n20729), .Z(n20771) );
  NANDN U22519 ( .A(n20732), .B(n20731), .Z(n20736) );
  NANDN U22520 ( .A(n20734), .B(n20733), .Z(n20735) );
  AND U22521 ( .A(n20736), .B(n20735), .Z(n20765) );
  NAND U22522 ( .A(n20738), .B(n20737), .Z(n20742) );
  NANDN U22523 ( .A(n20740), .B(n20739), .Z(n20741) );
  NAND U22524 ( .A(n20742), .B(n20741), .Z(n20760) );
  NAND U22525 ( .A(n20744), .B(n20743), .Z(n20748) );
  NAND U22526 ( .A(n20746), .B(n20745), .Z(n20747) );
  NAND U22527 ( .A(n20748), .B(n20747), .Z(n20759) );
  XOR U22528 ( .A(n20760), .B(n20759), .Z(n20761) );
  XNOR U22529 ( .A(n20882), .B(n20881), .Z(n20887) );
  NAND U22530 ( .A(n20753), .B(n20752), .Z(n20757) );
  NANDN U22531 ( .A(n20755), .B(n20754), .Z(n20756) );
  NAND U22532 ( .A(n20757), .B(n20756), .Z(n20885) );
  XOR U22533 ( .A(n20886), .B(n20885), .Z(n20758) );
  XNOR U22534 ( .A(n20887), .B(n20758), .Z(N439) );
  NAND U22535 ( .A(n20760), .B(n20759), .Z(n20764) );
  NANDN U22536 ( .A(n20762), .B(n20761), .Z(n20763) );
  AND U22537 ( .A(n20764), .B(n20763), .Z(n21025) );
  NANDN U22538 ( .A(n20766), .B(n20765), .Z(n20770) );
  NANDN U22539 ( .A(n20768), .B(n20767), .Z(n20769) );
  NAND U22540 ( .A(n20770), .B(n20769), .Z(n21023) );
  NANDN U22541 ( .A(n20772), .B(n20771), .Z(n20776) );
  NANDN U22542 ( .A(n20774), .B(n20773), .Z(n20775) );
  NAND U22543 ( .A(n20776), .B(n20775), .Z(n21005) );
  NANDN U22544 ( .A(n20778), .B(n20777), .Z(n20782) );
  NAND U22545 ( .A(n20780), .B(n20779), .Z(n20781) );
  AND U22546 ( .A(n20782), .B(n20781), .Z(n20999) );
  NAND U22547 ( .A(n20784), .B(n20783), .Z(n20788) );
  NANDN U22548 ( .A(n20786), .B(n20785), .Z(n20787) );
  AND U22549 ( .A(n20788), .B(n20787), .Z(n20997) );
  NAND U22550 ( .A(n20790), .B(n20789), .Z(n20794) );
  NANDN U22551 ( .A(n20792), .B(n20791), .Z(n20793) );
  NAND U22552 ( .A(n20794), .B(n20793), .Z(n20996) );
  NAND U22553 ( .A(n20796), .B(n20795), .Z(n20800) );
  NAND U22554 ( .A(n20798), .B(n20797), .Z(n20799) );
  AND U22555 ( .A(n20800), .B(n20799), .Z(n21015) );
  NAND U22556 ( .A(n20802), .B(n20801), .Z(n20806) );
  NAND U22557 ( .A(n20804), .B(n20803), .Z(n20805) );
  NAND U22558 ( .A(n20806), .B(n20805), .Z(n20943) );
  AND U22559 ( .A(n20808), .B(n20807), .Z(n20812) );
  NAND U22560 ( .A(n20810), .B(n20809), .Z(n20811) );
  NANDN U22561 ( .A(n20812), .B(n20811), .Z(n20942) );
  XOR U22562 ( .A(n20943), .B(n20942), .Z(n20945) );
  AND U22563 ( .A(y[7888]), .B(x[487]), .Z(n20814) );
  NAND U22564 ( .A(y[7886]), .B(x[489]), .Z(n20813) );
  XNOR U22565 ( .A(n20814), .B(n20813), .Z(n20911) );
  XOR U22566 ( .A(n20910), .B(n20911), .Z(n20949) );
  AND U22567 ( .A(x[490]), .B(y[7885]), .Z(n20948) );
  XOR U22568 ( .A(n20949), .B(n20948), .Z(n20951) );
  AND U22569 ( .A(x[486]), .B(y[7889]), .Z(n20901) );
  AND U22570 ( .A(x[495]), .B(y[7880]), .Z(n20902) );
  XOR U22571 ( .A(n20901), .B(n20902), .Z(n20904) );
  AND U22572 ( .A(x[491]), .B(y[7884]), .Z(n20903) );
  XOR U22573 ( .A(n20904), .B(n20903), .Z(n20950) );
  XOR U22574 ( .A(n20951), .B(n20950), .Z(n20944) );
  XOR U22575 ( .A(n20945), .B(n20944), .Z(n21014) );
  XOR U22576 ( .A(n21017), .B(n21016), .Z(n21003) );
  NAND U22577 ( .A(n20816), .B(n20815), .Z(n20820) );
  NAND U22578 ( .A(n20818), .B(n20817), .Z(n20819) );
  NAND U22579 ( .A(n20820), .B(n20819), .Z(n20937) );
  NAND U22580 ( .A(n20909), .B(n20910), .Z(n20824) );
  NAND U22581 ( .A(n20822), .B(n20821), .Z(n20823) );
  AND U22582 ( .A(n20824), .B(n20823), .Z(n20981) );
  AND U22583 ( .A(x[480]), .B(y[7895]), .Z(n20921) );
  AND U22584 ( .A(x[503]), .B(y[7872]), .Z(n20920) );
  XOR U22585 ( .A(n20921), .B(n20920), .Z(n20923) );
  AND U22586 ( .A(x[502]), .B(y[7873]), .Z(n20900) );
  XOR U22587 ( .A(n20900), .B(o[215]), .Z(n20922) );
  XOR U22588 ( .A(n20923), .B(n20922), .Z(n20979) );
  NAND U22589 ( .A(y[7875]), .B(x[500]), .Z(n20825) );
  XNOR U22590 ( .A(n20826), .B(n20825), .Z(n20896) );
  AND U22591 ( .A(x[499]), .B(y[7876]), .Z(n20897) );
  XOR U22592 ( .A(n20896), .B(n20897), .Z(n20978) );
  XOR U22593 ( .A(n20979), .B(n20978), .Z(n20980) );
  NAND U22594 ( .A(n20828), .B(n20827), .Z(n20832) );
  NAND U22595 ( .A(n20830), .B(n20829), .Z(n20831) );
  AND U22596 ( .A(n20832), .B(n20831), .Z(n20985) );
  AND U22597 ( .A(x[498]), .B(y[7882]), .Z(n21655) );
  NAND U22598 ( .A(n21655), .B(n20833), .Z(n20837) );
  NAND U22599 ( .A(n20835), .B(n20834), .Z(n20836) );
  NAND U22600 ( .A(n20837), .B(n20836), .Z(n20984) );
  XOR U22601 ( .A(n20987), .B(n20986), .Z(n20936) );
  XOR U22602 ( .A(n20937), .B(n20936), .Z(n20939) );
  AND U22603 ( .A(x[500]), .B(y[7881]), .Z(n21797) );
  AND U22604 ( .A(x[493]), .B(y[7874]), .Z(n20838) );
  NAND U22605 ( .A(n21797), .B(n20838), .Z(n20842) );
  NAND U22606 ( .A(n20840), .B(n20839), .Z(n20841) );
  NAND U22607 ( .A(n20842), .B(n20841), .Z(n20931) );
  NAND U22608 ( .A(n20844), .B(n20843), .Z(n20848) );
  NAND U22609 ( .A(n20846), .B(n20845), .Z(n20847) );
  AND U22610 ( .A(n20848), .B(n20847), .Z(n20993) );
  AND U22611 ( .A(x[493]), .B(y[7882]), .Z(n20966) );
  AND U22612 ( .A(x[482]), .B(y[7893]), .Z(n20967) );
  XOR U22613 ( .A(n20966), .B(n20967), .Z(n20968) );
  AND U22614 ( .A(x[501]), .B(y[7874]), .Z(n20969) );
  XOR U22615 ( .A(n20968), .B(n20969), .Z(n20991) );
  AND U22616 ( .A(x[492]), .B(y[7883]), .Z(n20914) );
  AND U22617 ( .A(x[481]), .B(y[7894]), .Z(n20915) );
  XOR U22618 ( .A(n20914), .B(n20915), .Z(n20916) );
  AND U22619 ( .A(n20849), .B(o[214]), .Z(n20917) );
  XOR U22620 ( .A(n20916), .B(n20917), .Z(n20990) );
  XOR U22621 ( .A(n20991), .B(n20990), .Z(n20992) );
  XOR U22622 ( .A(n20931), .B(n20930), .Z(n20933) );
  AND U22623 ( .A(x[495]), .B(y[7888]), .Z(n21960) );
  NAND U22624 ( .A(n21960), .B(n20850), .Z(n20854) );
  NANDN U22625 ( .A(n20852), .B(n20851), .Z(n20853) );
  AND U22626 ( .A(n20854), .B(n20853), .Z(n20975) );
  AND U22627 ( .A(x[494]), .B(y[7881]), .Z(n20961) );
  AND U22628 ( .A(x[483]), .B(y[7892]), .Z(n20960) );
  XOR U22629 ( .A(n20961), .B(n20960), .Z(n20963) );
  AND U22630 ( .A(x[484]), .B(y[7891]), .Z(n20962) );
  XOR U22631 ( .A(n20963), .B(n20962), .Z(n20973) );
  AND U22632 ( .A(x[485]), .B(y[7890]), .Z(n20954) );
  AND U22633 ( .A(x[498]), .B(y[7877]), .Z(n20955) );
  XOR U22634 ( .A(n20954), .B(n20955), .Z(n20956) );
  AND U22635 ( .A(x[497]), .B(y[7878]), .Z(n20957) );
  XOR U22636 ( .A(n20956), .B(n20957), .Z(n20972) );
  XOR U22637 ( .A(n20973), .B(n20972), .Z(n20974) );
  XOR U22638 ( .A(n20933), .B(n20932), .Z(n20938) );
  XOR U22639 ( .A(n20939), .B(n20938), .Z(n21002) );
  XOR U22640 ( .A(n21003), .B(n21002), .Z(n21004) );
  XNOR U22641 ( .A(n21005), .B(n21004), .Z(n20891) );
  NANDN U22642 ( .A(n20856), .B(n20855), .Z(n20860) );
  NAND U22643 ( .A(n20858), .B(n20857), .Z(n20859) );
  AND U22644 ( .A(n20860), .B(n20859), .Z(n21011) );
  NAND U22645 ( .A(n20862), .B(n20861), .Z(n20866) );
  NAND U22646 ( .A(n20864), .B(n20863), .Z(n20865) );
  AND U22647 ( .A(n20866), .B(n20865), .Z(n21009) );
  NAND U22648 ( .A(n20868), .B(n20867), .Z(n20872) );
  NANDN U22649 ( .A(n20870), .B(n20869), .Z(n20871) );
  AND U22650 ( .A(n20872), .B(n20871), .Z(n21008) );
  NANDN U22651 ( .A(n20874), .B(n20873), .Z(n20878) );
  NAND U22652 ( .A(n20876), .B(n20875), .Z(n20877) );
  AND U22653 ( .A(n20878), .B(n20877), .Z(n20889) );
  XOR U22654 ( .A(n20891), .B(n20892), .Z(n21024) );
  XOR U22655 ( .A(n21023), .B(n21024), .Z(n21026) );
  XNOR U22656 ( .A(n21025), .B(n21026), .Z(n21022) );
  NANDN U22657 ( .A(n20880), .B(n20879), .Z(n20884) );
  NAND U22658 ( .A(n20882), .B(n20881), .Z(n20883) );
  NAND U22659 ( .A(n20884), .B(n20883), .Z(n21020) );
  XOR U22660 ( .A(n21020), .B(n21021), .Z(n20888) );
  XNOR U22661 ( .A(n21022), .B(n20888), .Z(N440) );
  NANDN U22662 ( .A(n20890), .B(n20889), .Z(n20894) );
  NANDN U22663 ( .A(n20892), .B(n20891), .Z(n20893) );
  AND U22664 ( .A(n20894), .B(n20893), .Z(n21163) );
  AND U22665 ( .A(x[500]), .B(y[7879]), .Z(n20895) );
  NAND U22666 ( .A(n20895), .B(n21054), .Z(n20899) );
  NAND U22667 ( .A(n20897), .B(n20896), .Z(n20898) );
  NAND U22668 ( .A(n20899), .B(n20898), .Z(n21080) );
  AND U22669 ( .A(x[502]), .B(y[7874]), .Z(n21099) );
  XOR U22670 ( .A(n21100), .B(n21099), .Z(n21101) );
  NAND U22671 ( .A(x[482]), .B(y[7894]), .Z(n21102) );
  AND U22672 ( .A(x[481]), .B(y[7895]), .Z(n21107) );
  XOR U22673 ( .A(n21108), .B(n21107), .Z(n21106) );
  NAND U22674 ( .A(n20900), .B(o[215]), .Z(n21105) );
  XOR U22675 ( .A(n21078), .B(n21077), .Z(n21079) );
  XOR U22676 ( .A(n21080), .B(n21079), .Z(n21137) );
  NAND U22677 ( .A(n20902), .B(n20901), .Z(n20906) );
  NAND U22678 ( .A(n20904), .B(n20903), .Z(n20905) );
  NAND U22679 ( .A(n20906), .B(n20905), .Z(n21074) );
  AND U22680 ( .A(y[7880]), .B(x[496]), .Z(n20908) );
  NAND U22681 ( .A(y[7875]), .B(x[501]), .Z(n20907) );
  XNOR U22682 ( .A(n20908), .B(n20907), .Z(n21055) );
  AND U22683 ( .A(x[485]), .B(y[7891]), .Z(n21056) );
  XOR U22684 ( .A(n21055), .B(n21056), .Z(n21072) );
  AND U22685 ( .A(x[486]), .B(y[7890]), .Z(n21418) );
  AND U22686 ( .A(x[500]), .B(y[7876]), .Z(n21284) );
  XOR U22687 ( .A(n21418), .B(n21284), .Z(n21061) );
  AND U22688 ( .A(x[499]), .B(y[7877]), .Z(n21062) );
  XOR U22689 ( .A(n21061), .B(n21062), .Z(n21071) );
  XOR U22690 ( .A(n21072), .B(n21071), .Z(n21073) );
  XOR U22691 ( .A(n21074), .B(n21073), .Z(n21051) );
  NANDN U22692 ( .A(n21217), .B(n20909), .Z(n20913) );
  NAND U22693 ( .A(n20911), .B(n20910), .Z(n20912) );
  NAND U22694 ( .A(n20913), .B(n20912), .Z(n21049) );
  NAND U22695 ( .A(n20915), .B(n20914), .Z(n20919) );
  NAND U22696 ( .A(n20917), .B(n20916), .Z(n20918) );
  NAND U22697 ( .A(n20919), .B(n20918), .Z(n21048) );
  XOR U22698 ( .A(n21049), .B(n21048), .Z(n21050) );
  XOR U22699 ( .A(n21051), .B(n21050), .Z(n21136) );
  XOR U22700 ( .A(n21137), .B(n21136), .Z(n21139) );
  NAND U22701 ( .A(n20921), .B(n20920), .Z(n20925) );
  NAND U22702 ( .A(n20923), .B(n20922), .Z(n20924) );
  NAND U22703 ( .A(n20925), .B(n20924), .Z(n21130) );
  AND U22704 ( .A(x[483]), .B(y[7893]), .Z(n21120) );
  XOR U22705 ( .A(n21121), .B(n21120), .Z(n21119) );
  AND U22706 ( .A(x[484]), .B(y[7892]), .Z(n21118) );
  XOR U22707 ( .A(n21119), .B(n21118), .Z(n21131) );
  XOR U22708 ( .A(n21130), .B(n21131), .Z(n21133) );
  AND U22709 ( .A(y[7887]), .B(x[489]), .Z(n20927) );
  NAND U22710 ( .A(y[7886]), .B(x[490]), .Z(n20926) );
  XNOR U22711 ( .A(n20927), .B(n20926), .Z(n21091) );
  AND U22712 ( .A(y[7882]), .B(x[494]), .Z(n20929) );
  NAND U22713 ( .A(y[7888]), .B(x[488]), .Z(n20928) );
  XNOR U22714 ( .A(n20929), .B(n20928), .Z(n21095) );
  AND U22715 ( .A(x[491]), .B(y[7885]), .Z(n21096) );
  XOR U22716 ( .A(n21095), .B(n21096), .Z(n21090) );
  XOR U22717 ( .A(n21091), .B(n21090), .Z(n21132) );
  XOR U22718 ( .A(n21133), .B(n21132), .Z(n21138) );
  XNOR U22719 ( .A(n21139), .B(n21138), .Z(n21149) );
  NAND U22720 ( .A(n20931), .B(n20930), .Z(n20935) );
  NAND U22721 ( .A(n20933), .B(n20932), .Z(n20934) );
  AND U22722 ( .A(n20935), .B(n20934), .Z(n21148) );
  XOR U22723 ( .A(n21149), .B(n21148), .Z(n21150) );
  NAND U22724 ( .A(n20937), .B(n20936), .Z(n20941) );
  NAND U22725 ( .A(n20939), .B(n20938), .Z(n20940) );
  AND U22726 ( .A(n20941), .B(n20940), .Z(n21151) );
  XOR U22727 ( .A(n21150), .B(n21151), .Z(n21157) );
  NAND U22728 ( .A(n20943), .B(n20942), .Z(n20947) );
  NAND U22729 ( .A(n20945), .B(n20944), .Z(n20946) );
  NAND U22730 ( .A(n20947), .B(n20946), .Z(n21144) );
  NAND U22731 ( .A(n20949), .B(n20948), .Z(n20953) );
  NAND U22732 ( .A(n20951), .B(n20950), .Z(n20952) );
  NAND U22733 ( .A(n20953), .B(n20952), .Z(n21142) );
  NAND U22734 ( .A(n20955), .B(n20954), .Z(n20959) );
  NAND U22735 ( .A(n20957), .B(n20956), .Z(n20958) );
  NAND U22736 ( .A(n20959), .B(n20958), .Z(n21068) );
  AND U22737 ( .A(x[480]), .B(y[7896]), .Z(n21125) );
  AND U22738 ( .A(x[504]), .B(y[7872]), .Z(n21124) );
  XOR U22739 ( .A(n21125), .B(n21124), .Z(n21127) );
  AND U22740 ( .A(x[503]), .B(y[7873]), .Z(n21117) );
  XOR U22741 ( .A(n21117), .B(o[216]), .Z(n21126) );
  XOR U22742 ( .A(n21127), .B(n21126), .Z(n21066) );
  AND U22743 ( .A(x[487]), .B(y[7889]), .Z(n21111) );
  NAND U22744 ( .A(x[498]), .B(y[7878]), .Z(n21112) );
  NAND U22745 ( .A(x[497]), .B(y[7879]), .Z(n21114) );
  XOR U22746 ( .A(n21066), .B(n21065), .Z(n21067) );
  XOR U22747 ( .A(n21068), .B(n21067), .Z(n21045) );
  NAND U22748 ( .A(n20961), .B(n20960), .Z(n20965) );
  NAND U22749 ( .A(n20963), .B(n20962), .Z(n20964) );
  NAND U22750 ( .A(n20965), .B(n20964), .Z(n21043) );
  NAND U22751 ( .A(n20967), .B(n20966), .Z(n20971) );
  NAND U22752 ( .A(n20969), .B(n20968), .Z(n20970) );
  NAND U22753 ( .A(n20971), .B(n20970), .Z(n21042) );
  XOR U22754 ( .A(n21043), .B(n21042), .Z(n21044) );
  XOR U22755 ( .A(n21045), .B(n21044), .Z(n21143) );
  XOR U22756 ( .A(n21142), .B(n21143), .Z(n21145) );
  XNOR U22757 ( .A(n21144), .B(n21145), .Z(n21085) );
  NAND U22758 ( .A(n20973), .B(n20972), .Z(n20977) );
  NANDN U22759 ( .A(n20975), .B(n20974), .Z(n20976) );
  AND U22760 ( .A(n20977), .B(n20976), .Z(n21036) );
  NAND U22761 ( .A(n20979), .B(n20978), .Z(n20983) );
  NANDN U22762 ( .A(n20981), .B(n20980), .Z(n20982) );
  AND U22763 ( .A(n20983), .B(n20982), .Z(n21037) );
  XOR U22764 ( .A(n21036), .B(n21037), .Z(n21038) );
  NANDN U22765 ( .A(n20985), .B(n20984), .Z(n20989) );
  NAND U22766 ( .A(n20987), .B(n20986), .Z(n20988) );
  AND U22767 ( .A(n20989), .B(n20988), .Z(n21039) );
  XOR U22768 ( .A(n21038), .B(n21039), .Z(n21083) );
  NAND U22769 ( .A(n20991), .B(n20990), .Z(n20995) );
  NANDN U22770 ( .A(n20993), .B(n20992), .Z(n20994) );
  AND U22771 ( .A(n20995), .B(n20994), .Z(n21084) );
  XOR U22772 ( .A(n21083), .B(n21084), .Z(n21086) );
  XOR U22773 ( .A(n21085), .B(n21086), .Z(n21154) );
  NANDN U22774 ( .A(n20997), .B(n20996), .Z(n21001) );
  NANDN U22775 ( .A(n20999), .B(n20998), .Z(n21000) );
  NAND U22776 ( .A(n21001), .B(n21000), .Z(n21155) );
  XOR U22777 ( .A(n21157), .B(n21156), .Z(n21161) );
  NAND U22778 ( .A(n21003), .B(n21002), .Z(n21007) );
  NAND U22779 ( .A(n21005), .B(n21004), .Z(n21006) );
  AND U22780 ( .A(n21007), .B(n21006), .Z(n21033) );
  NANDN U22781 ( .A(n21009), .B(n21008), .Z(n21013) );
  NANDN U22782 ( .A(n21011), .B(n21010), .Z(n21012) );
  AND U22783 ( .A(n21013), .B(n21012), .Z(n21031) );
  NANDN U22784 ( .A(n21015), .B(n21014), .Z(n21019) );
  NAND U22785 ( .A(n21017), .B(n21016), .Z(n21018) );
  NAND U22786 ( .A(n21019), .B(n21018), .Z(n21030) );
  XNOR U22787 ( .A(n21163), .B(n21162), .Z(n21169) );
  NANDN U22788 ( .A(n21024), .B(n21023), .Z(n21028) );
  NANDN U22789 ( .A(n21026), .B(n21025), .Z(n21027) );
  AND U22790 ( .A(n21028), .B(n21027), .Z(n21167) );
  IV U22791 ( .A(n21167), .Z(n21166) );
  XOR U22792 ( .A(n21168), .B(n21166), .Z(n21029) );
  XNOR U22793 ( .A(n21169), .B(n21029), .Z(N441) );
  NANDN U22794 ( .A(n21031), .B(n21030), .Z(n21035) );
  NANDN U22795 ( .A(n21033), .B(n21032), .Z(n21034) );
  AND U22796 ( .A(n21035), .B(n21034), .Z(n21180) );
  NAND U22797 ( .A(n21037), .B(n21036), .Z(n21041) );
  NAND U22798 ( .A(n21039), .B(n21038), .Z(n21040) );
  AND U22799 ( .A(n21041), .B(n21040), .Z(n21190) );
  NAND U22800 ( .A(n21043), .B(n21042), .Z(n21047) );
  NAND U22801 ( .A(n21045), .B(n21044), .Z(n21046) );
  NAND U22802 ( .A(n21047), .B(n21046), .Z(n21208) );
  NAND U22803 ( .A(n21049), .B(n21048), .Z(n21053) );
  NAND U22804 ( .A(n21051), .B(n21050), .Z(n21052) );
  NAND U22805 ( .A(n21053), .B(n21052), .Z(n21207) );
  XOR U22806 ( .A(n21208), .B(n21207), .Z(n21210) );
  AND U22807 ( .A(x[501]), .B(y[7880]), .Z(n22012) );
  NAND U22808 ( .A(n22012), .B(n21054), .Z(n21058) );
  NAND U22809 ( .A(n21056), .B(n21055), .Z(n21057) );
  NAND U22810 ( .A(n21058), .B(n21057), .Z(n21302) );
  NAND U22811 ( .A(x[502]), .B(y[7875]), .Z(n21277) );
  NAND U22812 ( .A(x[485]), .B(y[7892]), .Z(n21275) );
  NAND U22813 ( .A(x[497]), .B(y[7880]), .Z(n21276) );
  XOR U22814 ( .A(n21275), .B(n21276), .Z(n21278) );
  XNOR U22815 ( .A(n21277), .B(n21278), .Z(n21301) );
  AND U22816 ( .A(y[7877]), .B(x[500]), .Z(n21060) );
  NAND U22817 ( .A(y[7876]), .B(x[501]), .Z(n21059) );
  XNOR U22818 ( .A(n21060), .B(n21059), .Z(n21286) );
  AND U22819 ( .A(x[499]), .B(y[7878]), .Z(n21285) );
  XOR U22820 ( .A(n21286), .B(n21285), .Z(n21300) );
  XNOR U22821 ( .A(n21301), .B(n21300), .Z(n21303) );
  XOR U22822 ( .A(n21302), .B(n21303), .Z(n21234) );
  NAND U22823 ( .A(n21284), .B(n21418), .Z(n21064) );
  NAND U22824 ( .A(n21062), .B(n21061), .Z(n21063) );
  NAND U22825 ( .A(n21064), .B(n21063), .Z(n21308) );
  NAND U22826 ( .A(x[495]), .B(y[7882]), .Z(n21292) );
  NAND U22827 ( .A(x[498]), .B(y[7879]), .Z(n21290) );
  NAND U22828 ( .A(x[486]), .B(y[7891]), .Z(n21291) );
  XOR U22829 ( .A(n21290), .B(n21291), .Z(n21293) );
  XNOR U22830 ( .A(n21292), .B(n21293), .Z(n21307) );
  NAND U22831 ( .A(x[503]), .B(y[7874]), .Z(n21274) );
  NAND U22832 ( .A(x[484]), .B(y[7893]), .Z(n21271) );
  NAND U22833 ( .A(x[496]), .B(y[7881]), .Z(n21272) );
  XOR U22834 ( .A(n21271), .B(n21272), .Z(n21273) );
  XNOR U22835 ( .A(n21274), .B(n21273), .Z(n21306) );
  XNOR U22836 ( .A(n21307), .B(n21306), .Z(n21309) );
  XOR U22837 ( .A(n21308), .B(n21309), .Z(n21233) );
  XOR U22838 ( .A(n21234), .B(n21233), .Z(n21236) );
  NAND U22839 ( .A(n21066), .B(n21065), .Z(n21070) );
  NAND U22840 ( .A(n21068), .B(n21067), .Z(n21069) );
  AND U22841 ( .A(n21070), .B(n21069), .Z(n21235) );
  XNOR U22842 ( .A(n21236), .B(n21235), .Z(n21248) );
  NAND U22843 ( .A(n21072), .B(n21071), .Z(n21076) );
  NAND U22844 ( .A(n21074), .B(n21073), .Z(n21075) );
  NAND U22845 ( .A(n21076), .B(n21075), .Z(n21246) );
  NAND U22846 ( .A(n21078), .B(n21077), .Z(n21082) );
  NAND U22847 ( .A(n21080), .B(n21079), .Z(n21081) );
  NAND U22848 ( .A(n21082), .B(n21081), .Z(n21245) );
  XOR U22849 ( .A(n21246), .B(n21245), .Z(n21247) );
  XOR U22850 ( .A(n21248), .B(n21247), .Z(n21209) );
  XNOR U22851 ( .A(n21210), .B(n21209), .Z(n21189) );
  NAND U22852 ( .A(n21084), .B(n21083), .Z(n21088) );
  NAND U22853 ( .A(n21086), .B(n21085), .Z(n21087) );
  NAND U22854 ( .A(n21088), .B(n21087), .Z(n21191) );
  XNOR U22855 ( .A(n21192), .B(n21191), .Z(n21186) );
  NANDN U22856 ( .A(n21218), .B(n21089), .Z(n21093) );
  NAND U22857 ( .A(n21091), .B(n21090), .Z(n21092) );
  NAND U22858 ( .A(n21093), .B(n21092), .Z(n21240) );
  AND U22859 ( .A(x[494]), .B(y[7888]), .Z(n22056) );
  NAND U22860 ( .A(n22056), .B(n21094), .Z(n21098) );
  NAND U22861 ( .A(n21096), .B(n21095), .Z(n21097) );
  NAND U22862 ( .A(n21098), .B(n21097), .Z(n21267) );
  NAND U22863 ( .A(x[491]), .B(y[7886]), .Z(n21282) );
  NAND U22864 ( .A(x[492]), .B(y[7885]), .Z(n21280) );
  NAND U22865 ( .A(x[487]), .B(y[7890]), .Z(n21281) );
  XOR U22866 ( .A(n21280), .B(n21281), .Z(n21283) );
  XNOR U22867 ( .A(n21282), .B(n21283), .Z(n21266) );
  AND U22868 ( .A(x[504]), .B(y[7873]), .Z(n21279) );
  XOR U22869 ( .A(o[217]), .B(n21279), .Z(n21254) );
  AND U22870 ( .A(x[481]), .B(y[7896]), .Z(n21253) );
  XOR U22871 ( .A(n21254), .B(n21253), .Z(n21256) );
  AND U22872 ( .A(x[493]), .B(y[7884]), .Z(n21255) );
  XOR U22873 ( .A(n21256), .B(n21255), .Z(n21265) );
  XOR U22874 ( .A(n21266), .B(n21265), .Z(n21268) );
  XOR U22875 ( .A(n21267), .B(n21268), .Z(n21239) );
  XOR U22876 ( .A(n21240), .B(n21239), .Z(n21242) );
  AND U22877 ( .A(n21100), .B(n21099), .Z(n21104) );
  NANDN U22878 ( .A(n21102), .B(n21101), .Z(n21103) );
  NANDN U22879 ( .A(n21104), .B(n21103), .Z(n21228) );
  ANDN U22880 ( .B(n21106), .A(n21105), .Z(n21110) );
  NAND U22881 ( .A(n21108), .B(n21107), .Z(n21109) );
  NANDN U22882 ( .A(n21110), .B(n21109), .Z(n21227) );
  XOR U22883 ( .A(n21228), .B(n21227), .Z(n21229) );
  NANDN U22884 ( .A(n21112), .B(n21111), .Z(n21116) );
  NANDN U22885 ( .A(n21114), .B(n21113), .Z(n21115) );
  NAND U22886 ( .A(n21116), .B(n21115), .Z(n21223) );
  NAND U22887 ( .A(x[488]), .B(y[7889]), .Z(n21219) );
  XOR U22888 ( .A(n21217), .B(n21218), .Z(n21220) );
  XNOR U22889 ( .A(n21219), .B(n21220), .Z(n21222) );
  NAND U22890 ( .A(n21117), .B(o[216]), .Z(n21216) );
  NAND U22891 ( .A(x[505]), .B(y[7872]), .Z(n21213) );
  NAND U22892 ( .A(x[480]), .B(y[7897]), .Z(n21214) );
  XOR U22893 ( .A(n21213), .B(n21214), .Z(n21215) );
  XNOR U22894 ( .A(n21216), .B(n21215), .Z(n21221) );
  XNOR U22895 ( .A(n21222), .B(n21221), .Z(n21224) );
  XOR U22896 ( .A(n21223), .B(n21224), .Z(n21230) );
  XNOR U22897 ( .A(n21229), .B(n21230), .Z(n21241) );
  XNOR U22898 ( .A(n21242), .B(n21241), .Z(n21198) );
  AND U22899 ( .A(n21119), .B(n21118), .Z(n21123) );
  NAND U22900 ( .A(n21121), .B(n21120), .Z(n21122) );
  NANDN U22901 ( .A(n21123), .B(n21122), .Z(n21297) );
  NAND U22902 ( .A(n21125), .B(n21124), .Z(n21129) );
  NAND U22903 ( .A(n21127), .B(n21126), .Z(n21128) );
  NAND U22904 ( .A(n21129), .B(n21128), .Z(n21295) );
  AND U22905 ( .A(x[494]), .B(y[7883]), .Z(n21260) );
  AND U22906 ( .A(x[482]), .B(y[7895]), .Z(n21259) );
  XOR U22907 ( .A(n21260), .B(n21259), .Z(n21262) );
  AND U22908 ( .A(x[483]), .B(y[7894]), .Z(n21261) );
  XOR U22909 ( .A(n21262), .B(n21261), .Z(n21294) );
  XOR U22910 ( .A(n21295), .B(n21294), .Z(n21296) );
  XNOR U22911 ( .A(n21297), .B(n21296), .Z(n21196) );
  NAND U22912 ( .A(n21131), .B(n21130), .Z(n21135) );
  NAND U22913 ( .A(n21133), .B(n21132), .Z(n21134) );
  AND U22914 ( .A(n21135), .B(n21134), .Z(n21195) );
  XOR U22915 ( .A(n21196), .B(n21195), .Z(n21197) );
  XOR U22916 ( .A(n21198), .B(n21197), .Z(n21202) );
  NAND U22917 ( .A(n21137), .B(n21136), .Z(n21141) );
  NAND U22918 ( .A(n21139), .B(n21138), .Z(n21140) );
  AND U22919 ( .A(n21141), .B(n21140), .Z(n21201) );
  XOR U22920 ( .A(n21202), .B(n21201), .Z(n21204) );
  NAND U22921 ( .A(n21143), .B(n21142), .Z(n21147) );
  NAND U22922 ( .A(n21145), .B(n21144), .Z(n21146) );
  AND U22923 ( .A(n21147), .B(n21146), .Z(n21203) );
  XNOR U22924 ( .A(n21204), .B(n21203), .Z(n21184) );
  NAND U22925 ( .A(n21149), .B(n21148), .Z(n21153) );
  NAND U22926 ( .A(n21151), .B(n21150), .Z(n21152) );
  AND U22927 ( .A(n21153), .B(n21152), .Z(n21183) );
  XOR U22928 ( .A(n21184), .B(n21183), .Z(n21185) );
  XNOR U22929 ( .A(n21186), .B(n21185), .Z(n21178) );
  NANDN U22930 ( .A(n21155), .B(n21154), .Z(n21159) );
  NAND U22931 ( .A(n21157), .B(n21156), .Z(n21158) );
  NAND U22932 ( .A(n21159), .B(n21158), .Z(n21177) );
  XOR U22933 ( .A(n21178), .B(n21177), .Z(n21179) );
  XNOR U22934 ( .A(n21180), .B(n21179), .Z(n21176) );
  NANDN U22935 ( .A(n21161), .B(n21160), .Z(n21165) );
  NAND U22936 ( .A(n21163), .B(n21162), .Z(n21164) );
  AND U22937 ( .A(n21165), .B(n21164), .Z(n21175) );
  OR U22938 ( .A(n21168), .B(n21166), .Z(n21172) );
  ANDN U22939 ( .B(n21168), .A(n21167), .Z(n21170) );
  OR U22940 ( .A(n21170), .B(n21169), .Z(n21171) );
  AND U22941 ( .A(n21172), .B(n21171), .Z(n21174) );
  XNOR U22942 ( .A(n21175), .B(n21174), .Z(n21173) );
  XNOR U22943 ( .A(n21176), .B(n21173), .Z(N442) );
  NAND U22944 ( .A(n21178), .B(n21177), .Z(n21182) );
  NAND U22945 ( .A(n21180), .B(n21179), .Z(n21181) );
  NAND U22946 ( .A(n21182), .B(n21181), .Z(n21454) );
  NAND U22947 ( .A(n21184), .B(n21183), .Z(n21188) );
  NAND U22948 ( .A(n21186), .B(n21185), .Z(n21187) );
  NAND U22949 ( .A(n21188), .B(n21187), .Z(n21449) );
  NANDN U22950 ( .A(n21190), .B(n21189), .Z(n21194) );
  NAND U22951 ( .A(n21192), .B(n21191), .Z(n21193) );
  AND U22952 ( .A(n21194), .B(n21193), .Z(n21448) );
  XOR U22953 ( .A(n21449), .B(n21448), .Z(n21451) );
  NAND U22954 ( .A(n21196), .B(n21195), .Z(n21200) );
  NAND U22955 ( .A(n21198), .B(n21197), .Z(n21199) );
  AND U22956 ( .A(n21200), .B(n21199), .Z(n21314) );
  NAND U22957 ( .A(n21202), .B(n21201), .Z(n21206) );
  NAND U22958 ( .A(n21204), .B(n21203), .Z(n21205) );
  AND U22959 ( .A(n21206), .B(n21205), .Z(n21313) );
  XOR U22960 ( .A(n21314), .B(n21313), .Z(n21315) );
  NAND U22961 ( .A(n21208), .B(n21207), .Z(n21212) );
  NAND U22962 ( .A(n21210), .B(n21209), .Z(n21211) );
  NAND U22963 ( .A(n21212), .B(n21211), .Z(n21444) );
  AND U22964 ( .A(x[482]), .B(y[7896]), .Z(n21331) );
  XOR U22965 ( .A(n21332), .B(n21331), .Z(n21334) );
  AND U22966 ( .A(x[504]), .B(y[7874]), .Z(n21333) );
  XOR U22967 ( .A(n21334), .B(n21333), .Z(n21366) );
  XOR U22968 ( .A(n21366), .B(n21365), .Z(n21368) );
  XNOR U22969 ( .A(n21368), .B(n21367), .Z(n21395) );
  NAND U22970 ( .A(n21222), .B(n21221), .Z(n21226) );
  NANDN U22971 ( .A(n21224), .B(n21223), .Z(n21225) );
  AND U22972 ( .A(n21226), .B(n21225), .Z(n21394) );
  XOR U22973 ( .A(n21395), .B(n21394), .Z(n21397) );
  NAND U22974 ( .A(n21228), .B(n21227), .Z(n21232) );
  NANDN U22975 ( .A(n21230), .B(n21229), .Z(n21231) );
  AND U22976 ( .A(n21232), .B(n21231), .Z(n21396) );
  XOR U22977 ( .A(n21397), .B(n21396), .Z(n21439) );
  NAND U22978 ( .A(n21234), .B(n21233), .Z(n21238) );
  NAND U22979 ( .A(n21236), .B(n21235), .Z(n21237) );
  NAND U22980 ( .A(n21238), .B(n21237), .Z(n21437) );
  NAND U22981 ( .A(n21240), .B(n21239), .Z(n21244) );
  NAND U22982 ( .A(n21242), .B(n21241), .Z(n21243) );
  AND U22983 ( .A(n21244), .B(n21243), .Z(n21436) );
  XOR U22984 ( .A(n21437), .B(n21436), .Z(n21438) );
  XNOR U22985 ( .A(n21439), .B(n21438), .Z(n21442) );
  NAND U22986 ( .A(n21246), .B(n21245), .Z(n21250) );
  NAND U22987 ( .A(n21248), .B(n21247), .Z(n21249) );
  NAND U22988 ( .A(n21250), .B(n21249), .Z(n21391) );
  AND U22989 ( .A(y[7892]), .B(x[486]), .Z(n21252) );
  NAND U22990 ( .A(y[7890]), .B(x[488]), .Z(n21251) );
  XNOR U22991 ( .A(n21252), .B(n21251), .Z(n21420) );
  AND U22992 ( .A(x[489]), .B(y[7889]), .Z(n21419) );
  XOR U22993 ( .A(n21420), .B(n21419), .Z(n21400) );
  NAND U22994 ( .A(x[487]), .B(y[7891]), .Z(n21401) );
  AND U22995 ( .A(x[492]), .B(y[7886]), .Z(n21503) );
  AND U22996 ( .A(x[485]), .B(y[7893]), .Z(n21375) );
  XOR U22997 ( .A(n21503), .B(n21375), .Z(n21377) );
  AND U22998 ( .A(x[490]), .B(y[7888]), .Z(n21376) );
  XOR U22999 ( .A(n21377), .B(n21376), .Z(n21402) );
  XOR U23000 ( .A(n21403), .B(n21402), .Z(n21356) );
  NAND U23001 ( .A(n21254), .B(n21253), .Z(n21258) );
  NAND U23002 ( .A(n21256), .B(n21255), .Z(n21257) );
  NAND U23003 ( .A(n21258), .B(n21257), .Z(n21354) );
  NAND U23004 ( .A(n21260), .B(n21259), .Z(n21264) );
  NAND U23005 ( .A(n21262), .B(n21261), .Z(n21263) );
  NAND U23006 ( .A(n21264), .B(n21263), .Z(n21353) );
  XOR U23007 ( .A(n21354), .B(n21353), .Z(n21355) );
  XNOR U23008 ( .A(n21356), .B(n21355), .Z(n21383) );
  NAND U23009 ( .A(n21266), .B(n21265), .Z(n21270) );
  NAND U23010 ( .A(n21268), .B(n21267), .Z(n21269) );
  AND U23011 ( .A(n21270), .B(n21269), .Z(n21382) );
  XOR U23012 ( .A(n21383), .B(n21382), .Z(n21385) );
  XNOR U23013 ( .A(n21319), .B(n21320), .Z(n21322) );
  NAND U23014 ( .A(x[494]), .B(y[7884]), .Z(n21413) );
  XNOR U23015 ( .A(n21412), .B(n21413), .Z(n21414) );
  NAND U23016 ( .A(x[481]), .B(y[7897]), .Z(n21415) );
  XNOR U23017 ( .A(n21414), .B(n21415), .Z(n21370) );
  NAND U23018 ( .A(x[505]), .B(y[7873]), .Z(n21421) );
  XNOR U23019 ( .A(o[218]), .B(n21421), .Z(n21379) );
  AND U23020 ( .A(x[506]), .B(y[7872]), .Z(n21378) );
  XOR U23021 ( .A(n21379), .B(n21378), .Z(n21381) );
  AND U23022 ( .A(x[480]), .B(y[7898]), .Z(n21380) );
  XOR U23023 ( .A(n21381), .B(n21380), .Z(n21369) );
  XOR U23024 ( .A(n21370), .B(n21369), .Z(n21372) );
  XOR U23025 ( .A(n21372), .B(n21371), .Z(n21321) );
  XNOR U23026 ( .A(n21322), .B(n21321), .Z(n21362) );
  AND U23027 ( .A(x[501]), .B(y[7877]), .Z(n21406) );
  NAND U23028 ( .A(n21284), .B(n21406), .Z(n21288) );
  NAND U23029 ( .A(n21286), .B(n21285), .Z(n21287) );
  NAND U23030 ( .A(n21288), .B(n21287), .Z(n21350) );
  XOR U23031 ( .A(n21407), .B(n21406), .Z(n21408) );
  NAND U23032 ( .A(x[500]), .B(y[7878]), .Z(n21409) );
  XNOR U23033 ( .A(n21408), .B(n21409), .Z(n21347) );
  NAND U23034 ( .A(x[503]), .B(y[7875]), .Z(n21336) );
  XNOR U23035 ( .A(n21335), .B(n21336), .Z(n21337) );
  NAND U23036 ( .A(x[502]), .B(y[7876]), .Z(n21338) );
  XNOR U23037 ( .A(n21337), .B(n21338), .Z(n21348) );
  XOR U23038 ( .A(n21347), .B(n21348), .Z(n21349) );
  XNOR U23039 ( .A(n21350), .B(n21349), .Z(n21360) );
  AND U23040 ( .A(x[484]), .B(y[7894]), .Z(n21341) );
  XOR U23041 ( .A(n21342), .B(n21341), .Z(n21343) );
  XOR U23042 ( .A(n21343), .B(n21289), .Z(n21325) );
  AND U23043 ( .A(x[499]), .B(y[7879]), .Z(n21422) );
  NAND U23044 ( .A(x[483]), .B(y[7895]), .Z(n21423) );
  XNOR U23045 ( .A(n21422), .B(n21423), .Z(n21424) );
  NAND U23046 ( .A(x[491]), .B(y[7887]), .Z(n21425) );
  XOR U23047 ( .A(n21424), .B(n21425), .Z(n21326) );
  XNOR U23048 ( .A(n21325), .B(n21326), .Z(n21328) );
  XNOR U23049 ( .A(n21328), .B(n21327), .Z(n21359) );
  XOR U23050 ( .A(n21360), .B(n21359), .Z(n21361) );
  XOR U23051 ( .A(n21362), .B(n21361), .Z(n21384) );
  XNOR U23052 ( .A(n21385), .B(n21384), .Z(n21389) );
  NAND U23053 ( .A(n21295), .B(n21294), .Z(n21299) );
  NAND U23054 ( .A(n21297), .B(n21296), .Z(n21298) );
  AND U23055 ( .A(n21299), .B(n21298), .Z(n21433) );
  NAND U23056 ( .A(n21301), .B(n21300), .Z(n21305) );
  NANDN U23057 ( .A(n21303), .B(n21302), .Z(n21304) );
  AND U23058 ( .A(n21305), .B(n21304), .Z(n21431) );
  NAND U23059 ( .A(n21307), .B(n21306), .Z(n21311) );
  NANDN U23060 ( .A(n21309), .B(n21308), .Z(n21310) );
  NAND U23061 ( .A(n21311), .B(n21310), .Z(n21430) );
  XOR U23062 ( .A(n21389), .B(n21388), .Z(n21390) );
  XNOR U23063 ( .A(n21391), .B(n21390), .Z(n21443) );
  XOR U23064 ( .A(n21442), .B(n21443), .Z(n21445) );
  XOR U23065 ( .A(n21444), .B(n21445), .Z(n21316) );
  XNOR U23066 ( .A(n21315), .B(n21316), .Z(n21450) );
  XOR U23067 ( .A(n21451), .B(n21450), .Z(n21456) );
  XOR U23068 ( .A(n21454), .B(n21456), .Z(n21312) );
  XOR U23069 ( .A(n21455), .B(n21312), .Z(N443) );
  NAND U23070 ( .A(n21314), .B(n21313), .Z(n21318) );
  NANDN U23071 ( .A(n21316), .B(n21315), .Z(n21317) );
  AND U23072 ( .A(n21318), .B(n21317), .Z(n21585) );
  NANDN U23073 ( .A(n21320), .B(n21319), .Z(n21324) );
  NAND U23074 ( .A(n21322), .B(n21321), .Z(n21323) );
  NAND U23075 ( .A(n21324), .B(n21323), .Z(n21563) );
  NANDN U23076 ( .A(n21326), .B(n21325), .Z(n21330) );
  NAND U23077 ( .A(n21328), .B(n21327), .Z(n21329) );
  NAND U23078 ( .A(n21330), .B(n21329), .Z(n21561) );
  NANDN U23079 ( .A(n21336), .B(n21335), .Z(n21340) );
  NANDN U23080 ( .A(n21338), .B(n21337), .Z(n21339) );
  NAND U23081 ( .A(n21340), .B(n21339), .Z(n21481) );
  XOR U23082 ( .A(n21480), .B(n21481), .Z(n21482) );
  AND U23083 ( .A(n21342), .B(n21341), .Z(n21346) );
  NANDN U23084 ( .A(n21344), .B(n21343), .Z(n21345) );
  NANDN U23085 ( .A(n21346), .B(n21345), .Z(n21491) );
  AND U23086 ( .A(x[480]), .B(y[7899]), .Z(n21543) );
  AND U23087 ( .A(x[507]), .B(y[7872]), .Z(n21542) );
  XOR U23088 ( .A(n21543), .B(n21542), .Z(n21546) );
  AND U23089 ( .A(x[506]), .B(y[7873]), .Z(n21554) );
  XOR U23090 ( .A(n21554), .B(o[219]), .Z(n21545) );
  XOR U23091 ( .A(n21546), .B(n21545), .Z(n21489) );
  AND U23092 ( .A(x[489]), .B(y[7890]), .Z(n21551) );
  AND U23093 ( .A(x[501]), .B(y[7878]), .Z(n21550) );
  XOR U23094 ( .A(n21551), .B(n21550), .Z(n21553) );
  AND U23095 ( .A(x[498]), .B(y[7881]), .Z(n21552) );
  XOR U23096 ( .A(n21553), .B(n21552), .Z(n21488) );
  XOR U23097 ( .A(n21489), .B(n21488), .Z(n21490) );
  XNOR U23098 ( .A(n21491), .B(n21490), .Z(n21483) );
  XNOR U23099 ( .A(n21482), .B(n21483), .Z(n21562) );
  XOR U23100 ( .A(n21561), .B(n21562), .Z(n21564) );
  XOR U23101 ( .A(n21563), .B(n21564), .Z(n21580) );
  NAND U23102 ( .A(n21348), .B(n21347), .Z(n21352) );
  NAND U23103 ( .A(n21350), .B(n21349), .Z(n21351) );
  AND U23104 ( .A(n21352), .B(n21351), .Z(n21578) );
  NAND U23105 ( .A(n21354), .B(n21353), .Z(n21358) );
  NAND U23106 ( .A(n21356), .B(n21355), .Z(n21357) );
  AND U23107 ( .A(n21358), .B(n21357), .Z(n21577) );
  XOR U23108 ( .A(n21578), .B(n21577), .Z(n21579) );
  NAND U23109 ( .A(n21360), .B(n21359), .Z(n21364) );
  NAND U23110 ( .A(n21362), .B(n21361), .Z(n21363) );
  AND U23111 ( .A(n21364), .B(n21363), .Z(n21565) );
  AND U23112 ( .A(x[495]), .B(y[7884]), .Z(n21509) );
  AND U23113 ( .A(x[482]), .B(y[7897]), .Z(n21508) );
  XOR U23114 ( .A(n21509), .B(n21508), .Z(n21511) );
  AND U23115 ( .A(x[483]), .B(y[7896]), .Z(n21510) );
  XOR U23116 ( .A(n21511), .B(n21510), .Z(n21529) );
  AND U23117 ( .A(x[486]), .B(y[7893]), .Z(n21537) );
  AND U23118 ( .A(x[505]), .B(y[7874]), .Z(n21535) );
  AND U23119 ( .A(x[499]), .B(y[7880]), .Z(n21534) );
  XOR U23120 ( .A(n21535), .B(n21534), .Z(n21536) );
  XOR U23121 ( .A(n21537), .B(n21536), .Z(n21528) );
  XOR U23122 ( .A(n21529), .B(n21528), .Z(n21530) );
  NAND U23123 ( .A(x[496]), .B(y[7883]), .Z(n21495) );
  XOR U23124 ( .A(n21495), .B(n21496), .Z(n21498) );
  XOR U23125 ( .A(n21497), .B(n21498), .Z(n21505) );
  AND U23126 ( .A(y[7886]), .B(x[493]), .Z(n21374) );
  AND U23127 ( .A(y[7887]), .B(x[492]), .Z(n21373) );
  XOR U23128 ( .A(n21374), .B(n21373), .Z(n21504) );
  XOR U23129 ( .A(n21505), .B(n21504), .Z(n21531) );
  XNOR U23130 ( .A(n21530), .B(n21531), .Z(n21479) );
  XOR U23131 ( .A(n21476), .B(n21477), .Z(n21478) );
  XOR U23132 ( .A(n21479), .B(n21478), .Z(n21557) );
  XNOR U23133 ( .A(n21558), .B(n21557), .Z(n21560) );
  XOR U23134 ( .A(n21559), .B(n21560), .Z(n21566) );
  NAND U23135 ( .A(n21383), .B(n21382), .Z(n21387) );
  NAND U23136 ( .A(n21385), .B(n21384), .Z(n21386) );
  AND U23137 ( .A(n21387), .B(n21386), .Z(n21567) );
  XOR U23138 ( .A(n21568), .B(n21567), .Z(n21464) );
  NAND U23139 ( .A(n21389), .B(n21388), .Z(n21393) );
  NAND U23140 ( .A(n21391), .B(n21390), .Z(n21392) );
  NAND U23141 ( .A(n21393), .B(n21392), .Z(n21466) );
  XOR U23142 ( .A(n21467), .B(n21466), .Z(n21461) );
  NAND U23143 ( .A(n21395), .B(n21394), .Z(n21399) );
  NAND U23144 ( .A(n21397), .B(n21396), .Z(n21398) );
  NAND U23145 ( .A(n21399), .B(n21398), .Z(n21471) );
  NANDN U23146 ( .A(n21401), .B(n21400), .Z(n21405) );
  NAND U23147 ( .A(n21403), .B(n21402), .Z(n21404) );
  NAND U23148 ( .A(n21405), .B(n21404), .Z(n21573) );
  AND U23149 ( .A(n21407), .B(n21406), .Z(n21411) );
  NANDN U23150 ( .A(n21409), .B(n21408), .Z(n21410) );
  NANDN U23151 ( .A(n21411), .B(n21410), .Z(n21520) );
  NANDN U23152 ( .A(n21413), .B(n21412), .Z(n21417) );
  NANDN U23153 ( .A(n21415), .B(n21414), .Z(n21416) );
  NAND U23154 ( .A(n21417), .B(n21416), .Z(n21521) );
  XOR U23155 ( .A(n21520), .B(n21521), .Z(n21522) );
  AND U23156 ( .A(x[488]), .B(y[7892]), .Z(n21556) );
  AND U23157 ( .A(x[494]), .B(y[7885]), .Z(n21513) );
  AND U23158 ( .A(x[481]), .B(y[7898]), .Z(n21512) );
  XOR U23159 ( .A(n21513), .B(n21512), .Z(n21516) );
  ANDN U23160 ( .B(o[218]), .A(n21421), .Z(n21515) );
  XOR U23161 ( .A(n21516), .B(n21515), .Z(n21485) );
  AND U23162 ( .A(x[497]), .B(y[7882]), .Z(n21539) );
  AND U23163 ( .A(x[484]), .B(y[7895]), .Z(n21538) );
  XOR U23164 ( .A(n21539), .B(n21538), .Z(n21541) );
  AND U23165 ( .A(x[485]), .B(y[7894]), .Z(n21540) );
  XOR U23166 ( .A(n21541), .B(n21540), .Z(n21484) );
  XOR U23167 ( .A(n21485), .B(n21484), .Z(n21486) );
  XNOR U23168 ( .A(n21487), .B(n21486), .Z(n21523) );
  XNOR U23169 ( .A(n21522), .B(n21523), .Z(n21572) );
  NANDN U23170 ( .A(n21423), .B(n21422), .Z(n21427) );
  NANDN U23171 ( .A(n21425), .B(n21424), .Z(n21426) );
  NAND U23172 ( .A(n21427), .B(n21426), .Z(n21526) );
  AND U23173 ( .A(y[7875]), .B(x[504]), .Z(n21429) );
  NAND U23174 ( .A(y[7879]), .B(x[500]), .Z(n21428) );
  XNOR U23175 ( .A(n21429), .B(n21428), .Z(n21533) );
  AND U23176 ( .A(x[487]), .B(y[7892]), .Z(n21532) );
  XOR U23177 ( .A(n21533), .B(n21532), .Z(n21525) );
  AND U23178 ( .A(x[488]), .B(y[7891]), .Z(n21500) );
  AND U23179 ( .A(x[503]), .B(y[7876]), .Z(n21499) );
  XOR U23180 ( .A(n21500), .B(n21499), .Z(n21502) );
  AND U23181 ( .A(x[502]), .B(y[7877]), .Z(n21501) );
  XOR U23182 ( .A(n21502), .B(n21501), .Z(n21524) );
  XOR U23183 ( .A(n21525), .B(n21524), .Z(n21527) );
  XOR U23184 ( .A(n21526), .B(n21527), .Z(n21571) );
  XOR U23185 ( .A(n21572), .B(n21571), .Z(n21574) );
  XNOR U23186 ( .A(n21573), .B(n21574), .Z(n21470) );
  XOR U23187 ( .A(n21471), .B(n21470), .Z(n21473) );
  NANDN U23188 ( .A(n21431), .B(n21430), .Z(n21435) );
  NANDN U23189 ( .A(n21433), .B(n21432), .Z(n21434) );
  AND U23190 ( .A(n21435), .B(n21434), .Z(n21472) );
  XOR U23191 ( .A(n21473), .B(n21472), .Z(n21459) );
  NAND U23192 ( .A(n21437), .B(n21436), .Z(n21441) );
  NAND U23193 ( .A(n21439), .B(n21438), .Z(n21440) );
  AND U23194 ( .A(n21441), .B(n21440), .Z(n21458) );
  XNOR U23195 ( .A(n21461), .B(n21460), .Z(n21584) );
  NANDN U23196 ( .A(n21443), .B(n21442), .Z(n21447) );
  NANDN U23197 ( .A(n21445), .B(n21444), .Z(n21446) );
  AND U23198 ( .A(n21447), .B(n21446), .Z(n21583) );
  XNOR U23199 ( .A(n21584), .B(n21583), .Z(n21586) );
  XNOR U23200 ( .A(n21585), .B(n21586), .Z(n21591) );
  NAND U23201 ( .A(n21449), .B(n21448), .Z(n21453) );
  NAND U23202 ( .A(n21451), .B(n21450), .Z(n21452) );
  NAND U23203 ( .A(n21453), .B(n21452), .Z(n21590) );
  XOR U23204 ( .A(n21590), .B(n21589), .Z(n21457) );
  XNOR U23205 ( .A(n21591), .B(n21457), .Z(N444) );
  NANDN U23206 ( .A(n21459), .B(n21458), .Z(n21463) );
  NAND U23207 ( .A(n21461), .B(n21460), .Z(n21462) );
  AND U23208 ( .A(n21463), .B(n21462), .Z(n21716) );
  NANDN U23209 ( .A(n21465), .B(n21464), .Z(n21469) );
  NAND U23210 ( .A(n21467), .B(n21466), .Z(n21468) );
  NAND U23211 ( .A(n21469), .B(n21468), .Z(n21715) );
  NAND U23212 ( .A(n21471), .B(n21470), .Z(n21475) );
  NAND U23213 ( .A(n21473), .B(n21472), .Z(n21474) );
  AND U23214 ( .A(n21475), .B(n21474), .Z(n21593) );
  NAND U23215 ( .A(n21489), .B(n21488), .Z(n21494) );
  IV U23216 ( .A(n21490), .Z(n21492) );
  NANDN U23217 ( .A(n21492), .B(n21491), .Z(n21493) );
  NAND U23218 ( .A(n21494), .B(n21493), .Z(n21694) );
  XOR U23219 ( .A(n21693), .B(n21694), .Z(n21696) );
  XOR U23220 ( .A(n21695), .B(n21696), .Z(n21616) );
  XOR U23221 ( .A(n21615), .B(n21616), .Z(n21618) );
  AND U23222 ( .A(x[487]), .B(y[7893]), .Z(n21649) );
  AND U23223 ( .A(x[492]), .B(y[7888]), .Z(n21648) );
  XOR U23224 ( .A(n21649), .B(n21648), .Z(n21651) );
  AND U23225 ( .A(x[491]), .B(y[7889]), .Z(n21650) );
  XOR U23226 ( .A(n21651), .B(n21650), .Z(n21664) );
  AND U23227 ( .A(x[507]), .B(y[7873]), .Z(n21662) );
  XOR U23228 ( .A(o[220]), .B(n21662), .Z(n21672) );
  AND U23229 ( .A(x[506]), .B(y[7874]), .Z(n21671) );
  XOR U23230 ( .A(n21672), .B(n21671), .Z(n21674) );
  AND U23231 ( .A(x[495]), .B(y[7885]), .Z(n21673) );
  XNOR U23232 ( .A(n21674), .B(n21673), .Z(n21663) );
  XNOR U23233 ( .A(n21664), .B(n21663), .Z(n21666) );
  XOR U23234 ( .A(n21665), .B(n21666), .Z(n21698) );
  AND U23235 ( .A(x[497]), .B(y[7883]), .Z(n21624) );
  AND U23236 ( .A(x[502]), .B(y[7878]), .Z(n21623) );
  XOR U23237 ( .A(n21624), .B(n21623), .Z(n21626) );
  AND U23238 ( .A(x[484]), .B(y[7896]), .Z(n21625) );
  XOR U23239 ( .A(n21626), .B(n21625), .Z(n21680) );
  AND U23240 ( .A(x[486]), .B(y[7894]), .Z(n21813) );
  AND U23241 ( .A(x[499]), .B(y[7881]), .Z(n21654) );
  XOR U23242 ( .A(n21813), .B(n21654), .Z(n21656) );
  XOR U23243 ( .A(n21656), .B(n21655), .Z(n21679) );
  XOR U23244 ( .A(n21680), .B(n21679), .Z(n21682) );
  XOR U23245 ( .A(n21681), .B(n21682), .Z(n21697) );
  XNOR U23246 ( .A(n21698), .B(n21697), .Z(n21700) );
  NAND U23247 ( .A(n21503), .B(n21668), .Z(n21507) );
  NANDN U23248 ( .A(n21505), .B(n21504), .Z(n21506) );
  NAND U23249 ( .A(n21507), .B(n21506), .Z(n21638) );
  IV U23250 ( .A(n21512), .Z(n21514) );
  NANDN U23251 ( .A(n21514), .B(n21513), .Z(n21519) );
  IV U23252 ( .A(n21515), .Z(n21517) );
  NANDN U23253 ( .A(n21517), .B(n21516), .Z(n21518) );
  NAND U23254 ( .A(n21519), .B(n21518), .Z(n21637) );
  XOR U23255 ( .A(n21636), .B(n21637), .Z(n21639) );
  XOR U23256 ( .A(n21638), .B(n21639), .Z(n21699) );
  XOR U23257 ( .A(n21700), .B(n21699), .Z(n21617) );
  XOR U23258 ( .A(n21618), .B(n21617), .Z(n21612) );
  XOR U23259 ( .A(n21683), .B(n21684), .Z(n21686) );
  XOR U23260 ( .A(n21685), .B(n21686), .Z(n21610) );
  AND U23261 ( .A(x[504]), .B(y[7879]), .Z(n21954) );
  AND U23262 ( .A(x[505]), .B(y[7875]), .Z(n21646) );
  XOR U23263 ( .A(n21647), .B(n21646), .Z(n21645) );
  AND U23264 ( .A(x[481]), .B(y[7899]), .Z(n21644) );
  XOR U23265 ( .A(n21645), .B(n21644), .Z(n21712) );
  AND U23266 ( .A(x[496]), .B(y[7884]), .Z(n21641) );
  AND U23267 ( .A(x[504]), .B(y[7876]), .Z(n21640) );
  XOR U23268 ( .A(n21641), .B(n21640), .Z(n21643) );
  AND U23269 ( .A(x[482]), .B(y[7898]), .Z(n21642) );
  XOR U23270 ( .A(n21643), .B(n21642), .Z(n21711) );
  XOR U23271 ( .A(n21712), .B(n21711), .Z(n21714) );
  XOR U23272 ( .A(n21713), .B(n21714), .Z(n21690) );
  AND U23273 ( .A(x[483]), .B(y[7897]), .Z(n21667) );
  XOR U23274 ( .A(n21668), .B(n21667), .Z(n21670) );
  AND U23275 ( .A(x[503]), .B(y[7877]), .Z(n21669) );
  XOR U23276 ( .A(n21670), .B(n21669), .Z(n21708) );
  AND U23277 ( .A(x[485]), .B(y[7895]), .Z(n21659) );
  AND U23278 ( .A(x[501]), .B(y[7879]), .Z(n21658) );
  XOR U23279 ( .A(n21659), .B(n21658), .Z(n21661) );
  AND U23280 ( .A(x[500]), .B(y[7880]), .Z(n21660) );
  XOR U23281 ( .A(n21661), .B(n21660), .Z(n21707) );
  XOR U23282 ( .A(n21708), .B(n21707), .Z(n21710) );
  XOR U23283 ( .A(n21709), .B(n21710), .Z(n21688) );
  IV U23284 ( .A(n21542), .Z(n21544) );
  NANDN U23285 ( .A(n21544), .B(n21543), .Z(n21549) );
  IV U23286 ( .A(n21545), .Z(n21547) );
  NANDN U23287 ( .A(n21547), .B(n21546), .Z(n21548) );
  NAND U23288 ( .A(n21549), .B(n21548), .Z(n21704) );
  XOR U23289 ( .A(n21703), .B(n21704), .Z(n21706) );
  AND U23290 ( .A(n21554), .B(o[219]), .Z(n21630) );
  AND U23291 ( .A(x[480]), .B(y[7900]), .Z(n21628) );
  AND U23292 ( .A(x[508]), .B(y[7872]), .Z(n21627) );
  XOR U23293 ( .A(n21628), .B(n21627), .Z(n21629) );
  XOR U23294 ( .A(n21630), .B(n21629), .Z(n21620) );
  NAND U23295 ( .A(y[7890]), .B(x[490]), .Z(n21555) );
  XNOR U23296 ( .A(n21556), .B(n21555), .Z(n21633) );
  AND U23297 ( .A(x[489]), .B(y[7891]), .Z(n21632) );
  XOR U23298 ( .A(n21633), .B(n21632), .Z(n21619) );
  XOR U23299 ( .A(n21620), .B(n21619), .Z(n21622) );
  XOR U23300 ( .A(n21621), .B(n21622), .Z(n21705) );
  XNOR U23301 ( .A(n21706), .B(n21705), .Z(n21687) );
  XNOR U23302 ( .A(n21688), .B(n21687), .Z(n21689) );
  XNOR U23303 ( .A(n21690), .B(n21689), .Z(n21609) );
  XNOR U23304 ( .A(n21610), .B(n21609), .Z(n21611) );
  XOR U23305 ( .A(n21612), .B(n21611), .Z(n21607) );
  XNOR U23306 ( .A(n21605), .B(n21606), .Z(n21608) );
  XOR U23307 ( .A(n21607), .B(n21608), .Z(n21594) );
  NANDN U23308 ( .A(n21566), .B(n21565), .Z(n21570) );
  NAND U23309 ( .A(n21568), .B(n21567), .Z(n21569) );
  NAND U23310 ( .A(n21570), .B(n21569), .Z(n21601) );
  NAND U23311 ( .A(n21572), .B(n21571), .Z(n21576) );
  NAND U23312 ( .A(n21574), .B(n21573), .Z(n21575) );
  NAND U23313 ( .A(n21576), .B(n21575), .Z(n21599) );
  NAND U23314 ( .A(n21578), .B(n21577), .Z(n21582) );
  NANDN U23315 ( .A(n21580), .B(n21579), .Z(n21581) );
  AND U23316 ( .A(n21582), .B(n21581), .Z(n21600) );
  XNOR U23317 ( .A(n21599), .B(n21600), .Z(n21602) );
  XNOR U23318 ( .A(n21595), .B(n21596), .Z(n21717) );
  XNOR U23319 ( .A(n21718), .B(n21717), .Z(n21723) );
  NAND U23320 ( .A(n21584), .B(n21583), .Z(n21588) );
  NANDN U23321 ( .A(n21586), .B(n21585), .Z(n21587) );
  AND U23322 ( .A(n21588), .B(n21587), .Z(n21721) );
  XNOR U23323 ( .A(n21721), .B(n21722), .Z(n21592) );
  XNOR U23324 ( .A(n21723), .B(n21592), .Z(N445) );
  NANDN U23325 ( .A(n21594), .B(n21593), .Z(n21598) );
  NANDN U23326 ( .A(n21596), .B(n21595), .Z(n21597) );
  NAND U23327 ( .A(n21598), .B(n21597), .Z(n21730) );
  NAND U23328 ( .A(n21600), .B(n21599), .Z(n21604) );
  NANDN U23329 ( .A(n21602), .B(n21601), .Z(n21603) );
  NAND U23330 ( .A(n21604), .B(n21603), .Z(n21728) );
  NANDN U23331 ( .A(n21610), .B(n21609), .Z(n21614) );
  NANDN U23332 ( .A(n21612), .B(n21611), .Z(n21613) );
  AND U23333 ( .A(n21614), .B(n21613), .Z(n21735) );
  XOR U23334 ( .A(n21734), .B(n21735), .Z(n21737) );
  XOR U23335 ( .A(n21879), .B(n21880), .Z(n21881) );
  AND U23336 ( .A(x[490]), .B(y[7892]), .Z(n21877) );
  NAND U23337 ( .A(n21631), .B(n21877), .Z(n21635) );
  NAND U23338 ( .A(n21633), .B(n21632), .Z(n21634) );
  NAND U23339 ( .A(n21635), .B(n21634), .Z(n21848) );
  AND U23340 ( .A(x[502]), .B(y[7879]), .Z(n21794) );
  AND U23341 ( .A(x[492]), .B(y[7889]), .Z(n21942) );
  AND U23342 ( .A(x[481]), .B(y[7900]), .Z(n21792) );
  XOR U23343 ( .A(n21942), .B(n21792), .Z(n21793) );
  XOR U23344 ( .A(n21794), .B(n21793), .Z(n21847) );
  AND U23345 ( .A(x[495]), .B(y[7886]), .Z(n21795) );
  XOR U23346 ( .A(n22012), .B(n21795), .Z(n21796) );
  XOR U23347 ( .A(n21797), .B(n21796), .Z(n21846) );
  XOR U23348 ( .A(n21847), .B(n21846), .Z(n21849) );
  XNOR U23349 ( .A(n21848), .B(n21849), .Z(n21882) );
  XOR U23350 ( .A(n21881), .B(n21882), .Z(n21842) );
  XOR U23351 ( .A(n21843), .B(n21842), .Z(n21845) );
  XOR U23352 ( .A(n21845), .B(n21844), .Z(n21841) );
  XOR U23353 ( .A(n21853), .B(n21852), .Z(n21854) );
  NAND U23354 ( .A(n21649), .B(n21648), .Z(n21653) );
  NAND U23355 ( .A(n21651), .B(n21650), .Z(n21652) );
  NAND U23356 ( .A(n21653), .B(n21652), .Z(n21758) );
  AND U23357 ( .A(x[491]), .B(y[7890]), .Z(n21810) );
  AND U23358 ( .A(x[483]), .B(y[7898]), .Z(n21808) );
  AND U23359 ( .A(x[497]), .B(y[7884]), .Z(n21807) );
  XOR U23360 ( .A(n21808), .B(n21807), .Z(n21809) );
  XOR U23361 ( .A(n21810), .B(n21809), .Z(n21757) );
  AND U23362 ( .A(x[503]), .B(y[7878]), .Z(n21804) );
  AND U23363 ( .A(x[493]), .B(y[7888]), .Z(n21802) );
  AND U23364 ( .A(x[504]), .B(y[7877]), .Z(n22062) );
  XOR U23365 ( .A(n21802), .B(n22062), .Z(n21803) );
  XOR U23366 ( .A(n21804), .B(n21803), .Z(n21756) );
  XOR U23367 ( .A(n21757), .B(n21756), .Z(n21759) );
  XNOR U23368 ( .A(n21758), .B(n21759), .Z(n21855) );
  AND U23369 ( .A(x[505]), .B(y[7876]), .Z(n21789) );
  AND U23370 ( .A(x[506]), .B(y[7875]), .Z(n21786) );
  XOR U23371 ( .A(n21787), .B(n21786), .Z(n21788) );
  XOR U23372 ( .A(n21789), .B(n21788), .Z(n21859) );
  IV U23373 ( .A(n21859), .Z(n21657) );
  AND U23374 ( .A(x[508]), .B(y[7873]), .Z(n21800) );
  XOR U23375 ( .A(o[221]), .B(n21800), .Z(n21872) );
  AND U23376 ( .A(x[480]), .B(y[7901]), .Z(n21870) );
  AND U23377 ( .A(x[509]), .B(y[7872]), .Z(n21869) );
  XOR U23378 ( .A(n21870), .B(n21869), .Z(n21871) );
  XNOR U23379 ( .A(n21872), .B(n21871), .Z(n21858) );
  XNOR U23380 ( .A(n21657), .B(n21858), .Z(n21860) );
  XOR U23381 ( .A(n21861), .B(n21860), .Z(n21828) );
  AND U23382 ( .A(n21662), .B(o[220]), .Z(n21765) );
  AND U23383 ( .A(x[496]), .B(y[7885]), .Z(n21763) );
  AND U23384 ( .A(x[507]), .B(y[7874]), .Z(n21762) );
  XOR U23385 ( .A(n21763), .B(n21762), .Z(n21764) );
  XOR U23386 ( .A(n21765), .B(n21764), .Z(n21822) );
  AND U23387 ( .A(x[482]), .B(y[7899]), .Z(n21774) );
  XOR U23388 ( .A(n21775), .B(n21774), .Z(n21776) );
  XOR U23389 ( .A(n21777), .B(n21776), .Z(n21821) );
  XOR U23390 ( .A(n21822), .B(n21821), .Z(n21824) );
  XOR U23391 ( .A(n21823), .B(n21824), .Z(n21829) );
  NAND U23392 ( .A(n21672), .B(n21671), .Z(n21676) );
  NAND U23393 ( .A(n21674), .B(n21673), .Z(n21675) );
  NAND U23394 ( .A(n21676), .B(n21675), .Z(n21780) );
  XOR U23395 ( .A(n21781), .B(n21780), .Z(n21783) );
  AND U23396 ( .A(x[488]), .B(y[7893]), .Z(n21815) );
  AND U23397 ( .A(y[7895]), .B(x[486]), .Z(n21678) );
  AND U23398 ( .A(y[7894]), .B(x[487]), .Z(n21677) );
  XOR U23399 ( .A(n21678), .B(n21677), .Z(n21814) );
  XOR U23400 ( .A(n21815), .B(n21814), .Z(n21864) );
  AND U23401 ( .A(x[489]), .B(y[7892]), .Z(n21933) );
  XOR U23402 ( .A(n21864), .B(n21933), .Z(n21866) );
  AND U23403 ( .A(x[485]), .B(y[7896]), .Z(n21771) );
  AND U23404 ( .A(x[484]), .B(y[7897]), .Z(n21769) );
  AND U23405 ( .A(x[490]), .B(y[7891]), .Z(n21768) );
  XOR U23406 ( .A(n21769), .B(n21768), .Z(n21770) );
  XOR U23407 ( .A(n21771), .B(n21770), .Z(n21865) );
  XOR U23408 ( .A(n21866), .B(n21865), .Z(n21782) );
  XOR U23409 ( .A(n21783), .B(n21782), .Z(n21751) );
  XOR U23410 ( .A(n21750), .B(n21751), .Z(n21753) );
  XOR U23411 ( .A(n21752), .B(n21753), .Z(n21838) );
  XOR U23412 ( .A(n21838), .B(n21839), .Z(n21840) );
  XNOR U23413 ( .A(n21841), .B(n21840), .Z(n21747) );
  XOR U23414 ( .A(n21746), .B(n21747), .Z(n21749) );
  NANDN U23415 ( .A(n21688), .B(n21687), .Z(n21692) );
  NANDN U23416 ( .A(n21690), .B(n21689), .Z(n21691) );
  AND U23417 ( .A(n21692), .B(n21691), .Z(n21743) );
  XOR U23418 ( .A(n21742), .B(n21743), .Z(n21745) );
  NANDN U23419 ( .A(n21698), .B(n21697), .Z(n21702) );
  NAND U23420 ( .A(n21700), .B(n21699), .Z(n21701) );
  NAND U23421 ( .A(n21702), .B(n21701), .Z(n21738) );
  XOR U23422 ( .A(n21834), .B(n21835), .Z(n21837) );
  XOR U23423 ( .A(n21836), .B(n21837), .Z(n21739) );
  XOR U23424 ( .A(n21738), .B(n21739), .Z(n21741) );
  XOR U23425 ( .A(n21740), .B(n21741), .Z(n21744) );
  XOR U23426 ( .A(n21745), .B(n21744), .Z(n21748) );
  XOR U23427 ( .A(n21749), .B(n21748), .Z(n21736) );
  XOR U23428 ( .A(n21737), .B(n21736), .Z(n21729) );
  XNOR U23429 ( .A(n21728), .B(n21729), .Z(n21731) );
  XOR U23430 ( .A(n21730), .B(n21731), .Z(n21727) );
  NANDN U23431 ( .A(n21716), .B(n21715), .Z(n21720) );
  NAND U23432 ( .A(n21718), .B(n21717), .Z(n21719) );
  NAND U23433 ( .A(n21720), .B(n21719), .Z(n21725) );
  XOR U23434 ( .A(n21725), .B(n21726), .Z(n21724) );
  XNOR U23435 ( .A(n21727), .B(n21724), .Z(N446) );
  NAND U23436 ( .A(n21729), .B(n21728), .Z(n21733) );
  NANDN U23437 ( .A(n21731), .B(n21730), .Z(n21732) );
  NAND U23438 ( .A(n21733), .B(n21732), .Z(n22160) );
  XOR U23439 ( .A(n22148), .B(n22147), .Z(n22145) );
  XOR U23440 ( .A(n22146), .B(n22145), .Z(n22142) );
  NANDN U23441 ( .A(n21751), .B(n21750), .Z(n21755) );
  NANDN U23442 ( .A(n21753), .B(n21752), .Z(n21754) );
  AND U23443 ( .A(n21755), .B(n21754), .Z(n21883) );
  NAND U23444 ( .A(n21757), .B(n21756), .Z(n21761) );
  NAND U23445 ( .A(n21759), .B(n21758), .Z(n21760) );
  AND U23446 ( .A(n21761), .B(n21760), .Z(n21891) );
  NAND U23447 ( .A(n21763), .B(n21762), .Z(n21767) );
  NAND U23448 ( .A(n21765), .B(n21764), .Z(n21766) );
  NAND U23449 ( .A(n21767), .B(n21766), .Z(n21901) );
  NAND U23450 ( .A(n21769), .B(n21768), .Z(n21773) );
  NAND U23451 ( .A(n21771), .B(n21770), .Z(n21772) );
  NAND U23452 ( .A(n21773), .B(n21772), .Z(n21904) );
  AND U23453 ( .A(x[486]), .B(y[7896]), .Z(n22004) );
  AND U23454 ( .A(x[485]), .B(y[7897]), .Z(n22006) );
  AND U23455 ( .A(x[499]), .B(y[7883]), .Z(n22005) );
  XOR U23456 ( .A(n22006), .B(n22005), .Z(n22003) );
  XNOR U23457 ( .A(n22004), .B(n22003), .Z(n22045) );
  AND U23458 ( .A(x[484]), .B(y[7898]), .Z(n22016) );
  AND U23459 ( .A(x[483]), .B(y[7899]), .Z(n22018) );
  AND U23460 ( .A(x[498]), .B(y[7884]), .Z(n22017) );
  XOR U23461 ( .A(n22018), .B(n22017), .Z(n22015) );
  XOR U23462 ( .A(n22016), .B(n22015), .Z(n22048) );
  NAND U23463 ( .A(n21775), .B(n21774), .Z(n21779) );
  NAND U23464 ( .A(n21777), .B(n21776), .Z(n21778) );
  AND U23465 ( .A(n21779), .B(n21778), .Z(n22047) );
  XOR U23466 ( .A(n22045), .B(n22046), .Z(n21903) );
  XOR U23467 ( .A(n21904), .B(n21903), .Z(n21902) );
  XOR U23468 ( .A(n21901), .B(n21902), .Z(n21892) );
  NAND U23469 ( .A(n21781), .B(n21780), .Z(n21785) );
  NAND U23470 ( .A(n21783), .B(n21782), .Z(n21784) );
  AND U23471 ( .A(n21785), .B(n21784), .Z(n21889) );
  XOR U23472 ( .A(n21890), .B(n21889), .Z(n21886) );
  IV U23473 ( .A(n21886), .Z(n21827) );
  AND U23474 ( .A(n21787), .B(n21786), .Z(n21791) );
  NAND U23475 ( .A(n21789), .B(n21788), .Z(n21790) );
  NANDN U23476 ( .A(n21791), .B(n21790), .Z(n21927) );
  AND U23477 ( .A(x[503]), .B(y[7879]), .Z(n22060) );
  AND U23478 ( .A(x[504]), .B(y[7878]), .Z(n21799) );
  AND U23479 ( .A(y[7877]), .B(x[505]), .Z(n21798) );
  XOR U23480 ( .A(n21799), .B(n21798), .Z(n22059) );
  XOR U23481 ( .A(n22060), .B(n22059), .Z(n21910) );
  IV U23482 ( .A(n21910), .Z(n21801) );
  AND U23483 ( .A(n21800), .B(o[221]), .Z(n22074) );
  AND U23484 ( .A(x[508]), .B(y[7874]), .Z(n22076) );
  AND U23485 ( .A(x[496]), .B(y[7886]), .Z(n22075) );
  XOR U23486 ( .A(n22076), .B(n22075), .Z(n22073) );
  XNOR U23487 ( .A(n22074), .B(n22073), .Z(n21909) );
  XOR U23488 ( .A(n21801), .B(n21909), .Z(n21907) );
  XNOR U23489 ( .A(n21908), .B(n21907), .Z(n21929) );
  XOR U23490 ( .A(n21930), .B(n21929), .Z(n21928) );
  XOR U23491 ( .A(n21927), .B(n21928), .Z(n22110) );
  NAND U23492 ( .A(n21802), .B(n22062), .Z(n21806) );
  NAND U23493 ( .A(n21804), .B(n21803), .Z(n21805) );
  NAND U23494 ( .A(n21806), .B(n21805), .Z(n21898) );
  NAND U23495 ( .A(n21808), .B(n21807), .Z(n21812) );
  NAND U23496 ( .A(n21810), .B(n21809), .Z(n21811) );
  AND U23497 ( .A(n21812), .B(n21811), .Z(n21920) );
  AND U23498 ( .A(x[480]), .B(y[7902]), .Z(n21948) );
  AND U23499 ( .A(x[509]), .B(y[7873]), .Z(n21953) );
  XOR U23500 ( .A(o[222]), .B(n21953), .Z(n21950) );
  AND U23501 ( .A(x[510]), .B(y[7872]), .Z(n21949) );
  XOR U23502 ( .A(n21950), .B(n21949), .Z(n21947) );
  XOR U23503 ( .A(n21948), .B(n21947), .Z(n21922) );
  AND U23504 ( .A(x[500]), .B(y[7882]), .Z(n22055) );
  XOR U23505 ( .A(n22056), .B(n22055), .Z(n22054) );
  AND U23506 ( .A(x[488]), .B(y[7894]), .Z(n22053) );
  XNOR U23507 ( .A(n22054), .B(n22053), .Z(n21921) );
  XNOR U23508 ( .A(n21920), .B(n21919), .Z(n21897) );
  XOR U23509 ( .A(n21898), .B(n21897), .Z(n21895) );
  AND U23510 ( .A(x[487]), .B(y[7895]), .Z(n22010) );
  NAND U23511 ( .A(n21813), .B(n22010), .Z(n21817) );
  NAND U23512 ( .A(n21815), .B(n21814), .Z(n21816) );
  AND U23513 ( .A(n21817), .B(n21816), .Z(n21913) );
  AND U23514 ( .A(y[7881]), .B(x[501]), .Z(n21819) );
  AND U23515 ( .A(y[7880]), .B(x[502]), .Z(n21818) );
  XOR U23516 ( .A(n21819), .B(n21818), .Z(n22009) );
  XOR U23517 ( .A(n22010), .B(n22009), .Z(n21916) );
  AND U23518 ( .A(x[497]), .B(y[7885]), .Z(n22068) );
  AND U23519 ( .A(x[482]), .B(y[7900]), .Z(n22070) );
  AND U23520 ( .A(x[506]), .B(y[7876]), .Z(n22069) );
  XOR U23521 ( .A(n22070), .B(n22069), .Z(n22067) );
  XNOR U23522 ( .A(n22068), .B(n22067), .Z(n21915) );
  XNOR U23523 ( .A(n21913), .B(n21914), .Z(n21896) );
  IV U23524 ( .A(n21896), .Z(n21820) );
  XOR U23525 ( .A(n21895), .B(n21820), .Z(n22112) );
  NAND U23526 ( .A(n21822), .B(n21821), .Z(n21826) );
  NAND U23527 ( .A(n21824), .B(n21823), .Z(n21825) );
  NAND U23528 ( .A(n21826), .B(n21825), .Z(n22111) );
  XOR U23529 ( .A(n22112), .B(n22111), .Z(n22109) );
  XOR U23530 ( .A(n22110), .B(n22109), .Z(n21885) );
  XNOR U23531 ( .A(n21827), .B(n21885), .Z(n21884) );
  XOR U23532 ( .A(n21883), .B(n21884), .Z(n22127) );
  NANDN U23533 ( .A(n21829), .B(n21828), .Z(n21833) );
  NANDN U23534 ( .A(n21831), .B(n21830), .Z(n21832) );
  NAND U23535 ( .A(n21833), .B(n21832), .Z(n22129) );
  XOR U23536 ( .A(n22129), .B(n22130), .Z(n22128) );
  XOR U23537 ( .A(n22127), .B(n22128), .Z(n22121) );
  NAND U23538 ( .A(n21847), .B(n21846), .Z(n21851) );
  NAND U23539 ( .A(n21849), .B(n21848), .Z(n21850) );
  AND U23540 ( .A(n21851), .B(n21850), .Z(n22094) );
  NAND U23541 ( .A(n21853), .B(n21852), .Z(n21857) );
  NANDN U23542 ( .A(n21855), .B(n21854), .Z(n21856) );
  AND U23543 ( .A(n21857), .B(n21856), .Z(n22093) );
  XOR U23544 ( .A(n22094), .B(n22093), .Z(n22092) );
  NANDN U23545 ( .A(n21859), .B(n21858), .Z(n21863) );
  OR U23546 ( .A(n21861), .B(n21860), .Z(n21862) );
  NAND U23547 ( .A(n21863), .B(n21862), .Z(n22091) );
  XOR U23548 ( .A(n22092), .B(n22091), .Z(n22106) );
  NAND U23549 ( .A(n21864), .B(n21933), .Z(n21868) );
  NAND U23550 ( .A(n21866), .B(n21865), .Z(n21867) );
  AND U23551 ( .A(n21868), .B(n21867), .Z(n22087) );
  NAND U23552 ( .A(n21870), .B(n21869), .Z(n21874) );
  NAND U23553 ( .A(n21872), .B(n21871), .Z(n21873) );
  NAND U23554 ( .A(n21874), .B(n21873), .Z(n22041) );
  AND U23555 ( .A(y[7890]), .B(x[492]), .Z(n21875) );
  XOR U23556 ( .A(n21876), .B(n21875), .Z(n21940) );
  XOR U23557 ( .A(n21941), .B(n21940), .Z(n21932) );
  AND U23558 ( .A(y[7893]), .B(x[489]), .Z(n21878) );
  XOR U23559 ( .A(n21878), .B(n21877), .Z(n21931) );
  XOR U23560 ( .A(n21932), .B(n21931), .Z(n22044) );
  AND U23561 ( .A(x[507]), .B(y[7875]), .Z(n21937) );
  AND U23562 ( .A(x[481]), .B(y[7901]), .Z(n21936) );
  XOR U23563 ( .A(n21937), .B(n21936), .Z(n21934) );
  XOR U23564 ( .A(n21935), .B(n21934), .Z(n22043) );
  XOR U23565 ( .A(n22044), .B(n22043), .Z(n22042) );
  XOR U23566 ( .A(n22041), .B(n22042), .Z(n22088) );
  XNOR U23567 ( .A(n22086), .B(n22085), .Z(n22105) );
  XOR U23568 ( .A(n22104), .B(n22103), .Z(n22124) );
  XNOR U23569 ( .A(n22123), .B(n22124), .Z(n22122) );
  XOR U23570 ( .A(n22121), .B(n22122), .Z(n22141) );
  XOR U23571 ( .A(n22139), .B(n22140), .Z(n22157) );
  XNOR U23572 ( .A(n22158), .B(n22157), .Z(N447) );
  NANDN U23573 ( .A(n21884), .B(n21883), .Z(n21888) );
  NANDN U23574 ( .A(n21886), .B(n21885), .Z(n21887) );
  AND U23575 ( .A(n21888), .B(n21887), .Z(n22156) );
  NAND U23576 ( .A(n21890), .B(n21889), .Z(n21894) );
  NANDN U23577 ( .A(n21892), .B(n21891), .Z(n21893) );
  AND U23578 ( .A(n21894), .B(n21893), .Z(n22138) );
  NANDN U23579 ( .A(n21896), .B(n21895), .Z(n21900) );
  NAND U23580 ( .A(n21898), .B(n21897), .Z(n21899) );
  AND U23581 ( .A(n21900), .B(n21899), .Z(n22120) );
  NAND U23582 ( .A(n21902), .B(n21901), .Z(n21906) );
  NAND U23583 ( .A(n21904), .B(n21903), .Z(n21905) );
  AND U23584 ( .A(n21906), .B(n21905), .Z(n22102) );
  NAND U23585 ( .A(n21908), .B(n21907), .Z(n21912) );
  NANDN U23586 ( .A(n21910), .B(n21909), .Z(n21911) );
  AND U23587 ( .A(n21912), .B(n21911), .Z(n22084) );
  NANDN U23588 ( .A(n21914), .B(n21913), .Z(n21918) );
  NANDN U23589 ( .A(n21916), .B(n21915), .Z(n21917) );
  AND U23590 ( .A(n21918), .B(n21917), .Z(n21926) );
  NAND U23591 ( .A(n21920), .B(n21919), .Z(n21924) );
  NANDN U23592 ( .A(n21922), .B(n21921), .Z(n21923) );
  NAND U23593 ( .A(n21924), .B(n21923), .Z(n21925) );
  XNOR U23594 ( .A(n21926), .B(n21925), .Z(n22082) );
  AND U23595 ( .A(x[490]), .B(y[7893]), .Z(n21968) );
  NAND U23596 ( .A(n21935), .B(n21934), .Z(n21939) );
  NAND U23597 ( .A(n21937), .B(n21936), .Z(n21938) );
  AND U23598 ( .A(n21939), .B(n21938), .Z(n21946) );
  NAND U23599 ( .A(n21941), .B(n21940), .Z(n21944) );
  NAND U23600 ( .A(n21959), .B(n21942), .Z(n21943) );
  NAND U23601 ( .A(n21944), .B(n21943), .Z(n21945) );
  NAND U23602 ( .A(n21948), .B(n21947), .Z(n21952) );
  NAND U23603 ( .A(n21950), .B(n21949), .Z(n21951) );
  AND U23604 ( .A(n21952), .B(n21951), .Z(n22002) );
  AND U23605 ( .A(n21953), .B(o[222]), .Z(n21958) );
  AND U23606 ( .A(y[7903]), .B(x[480]), .Z(n21956) );
  XNOR U23607 ( .A(n21954), .B(o[223]), .Z(n21955) );
  XNOR U23608 ( .A(n21956), .B(n21955), .Z(n21957) );
  XOR U23609 ( .A(n21958), .B(n21957), .Z(n21962) );
  XNOR U23610 ( .A(n21960), .B(n21959), .Z(n21961) );
  XNOR U23611 ( .A(n21962), .B(n21961), .Z(n22000) );
  AND U23612 ( .A(y[7884]), .B(x[499]), .Z(n21964) );
  NAND U23613 ( .A(y[7882]), .B(x[501]), .Z(n21963) );
  XNOR U23614 ( .A(n21964), .B(n21963), .Z(n21972) );
  AND U23615 ( .A(y[7895]), .B(x[488]), .Z(n21970) );
  AND U23616 ( .A(y[7892]), .B(x[491]), .Z(n21966) );
  NAND U23617 ( .A(y[7877]), .B(x[506]), .Z(n21965) );
  XNOR U23618 ( .A(n21966), .B(n21965), .Z(n21967) );
  XNOR U23619 ( .A(n21968), .B(n21967), .Z(n21969) );
  XNOR U23620 ( .A(n21970), .B(n21969), .Z(n21971) );
  XOR U23621 ( .A(n21972), .B(n21971), .Z(n21974) );
  AND U23622 ( .A(x[505]), .B(y[7878]), .Z(n22061) );
  AND U23623 ( .A(x[502]), .B(y[7881]), .Z(n22011) );
  XNOR U23624 ( .A(n22061), .B(n22011), .Z(n21973) );
  XNOR U23625 ( .A(n21974), .B(n21973), .Z(n21990) );
  AND U23626 ( .A(y[7876]), .B(x[507]), .Z(n21976) );
  NAND U23627 ( .A(y[7875]), .B(x[508]), .Z(n21975) );
  XNOR U23628 ( .A(n21976), .B(n21975), .Z(n21980) );
  AND U23629 ( .A(y[7896]), .B(x[487]), .Z(n21978) );
  NAND U23630 ( .A(y[7902]), .B(x[481]), .Z(n21977) );
  XNOR U23631 ( .A(n21978), .B(n21977), .Z(n21979) );
  XOR U23632 ( .A(n21980), .B(n21979), .Z(n21988) );
  AND U23633 ( .A(y[7901]), .B(x[482]), .Z(n21982) );
  NAND U23634 ( .A(y[7891]), .B(x[492]), .Z(n21981) );
  XNOR U23635 ( .A(n21982), .B(n21981), .Z(n21986) );
  AND U23636 ( .A(y[7880]), .B(x[503]), .Z(n21984) );
  NAND U23637 ( .A(y[7886]), .B(x[497]), .Z(n21983) );
  XNOR U23638 ( .A(n21984), .B(n21983), .Z(n21985) );
  XNOR U23639 ( .A(n21986), .B(n21985), .Z(n21987) );
  XNOR U23640 ( .A(n21988), .B(n21987), .Z(n21989) );
  XOR U23641 ( .A(n21990), .B(n21989), .Z(n21998) );
  AND U23642 ( .A(y[7887]), .B(x[496]), .Z(n21992) );
  NAND U23643 ( .A(y[7883]), .B(x[500]), .Z(n21991) );
  XNOR U23644 ( .A(n21992), .B(n21991), .Z(n21996) );
  AND U23645 ( .A(y[7873]), .B(x[510]), .Z(n21994) );
  NAND U23646 ( .A(y[7889]), .B(x[494]), .Z(n21993) );
  XNOR U23647 ( .A(n21994), .B(n21993), .Z(n21995) );
  XNOR U23648 ( .A(n21996), .B(n21995), .Z(n21997) );
  XNOR U23649 ( .A(n21998), .B(n21997), .Z(n21999) );
  XNOR U23650 ( .A(n22000), .B(n21999), .Z(n22001) );
  NAND U23651 ( .A(n22004), .B(n22003), .Z(n22008) );
  NAND U23652 ( .A(n22006), .B(n22005), .Z(n22007) );
  AND U23653 ( .A(n22008), .B(n22007), .Z(n22040) );
  NAND U23654 ( .A(n22010), .B(n22009), .Z(n22014) );
  NAND U23655 ( .A(n22012), .B(n22011), .Z(n22013) );
  AND U23656 ( .A(n22014), .B(n22013), .Z(n22022) );
  NAND U23657 ( .A(n22016), .B(n22015), .Z(n22020) );
  NAND U23658 ( .A(n22018), .B(n22017), .Z(n22019) );
  NAND U23659 ( .A(n22020), .B(n22019), .Z(n22021) );
  XNOR U23660 ( .A(n22022), .B(n22021), .Z(n22038) );
  AND U23661 ( .A(y[7872]), .B(x[511]), .Z(n22024) );
  NAND U23662 ( .A(y[7899]), .B(x[484]), .Z(n22023) );
  XNOR U23663 ( .A(n22024), .B(n22023), .Z(n22028) );
  AND U23664 ( .A(y[7898]), .B(x[485]), .Z(n22026) );
  NAND U23665 ( .A(y[7897]), .B(x[486]), .Z(n22025) );
  XNOR U23666 ( .A(n22026), .B(n22025), .Z(n22027) );
  XOR U23667 ( .A(n22028), .B(n22027), .Z(n22036) );
  AND U23668 ( .A(y[7900]), .B(x[483]), .Z(n22030) );
  NAND U23669 ( .A(y[7885]), .B(x[498]), .Z(n22029) );
  XNOR U23670 ( .A(n22030), .B(n22029), .Z(n22034) );
  AND U23671 ( .A(y[7874]), .B(x[509]), .Z(n22032) );
  NAND U23672 ( .A(y[7894]), .B(x[489]), .Z(n22031) );
  XNOR U23673 ( .A(n22032), .B(n22031), .Z(n22033) );
  XNOR U23674 ( .A(n22034), .B(n22033), .Z(n22035) );
  XNOR U23675 ( .A(n22036), .B(n22035), .Z(n22037) );
  XNOR U23676 ( .A(n22038), .B(n22037), .Z(n22039) );
  NANDN U23677 ( .A(n22046), .B(n22045), .Z(n22050) );
  NANDN U23678 ( .A(n22048), .B(n22047), .Z(n22049) );
  NAND U23679 ( .A(n22050), .B(n22049), .Z(n22051) );
  NAND U23680 ( .A(n22054), .B(n22053), .Z(n22058) );
  NAND U23681 ( .A(n22056), .B(n22055), .Z(n22057) );
  AND U23682 ( .A(n22058), .B(n22057), .Z(n22066) );
  NAND U23683 ( .A(n22060), .B(n22059), .Z(n22064) );
  NAND U23684 ( .A(n22062), .B(n22061), .Z(n22063) );
  NAND U23685 ( .A(n22064), .B(n22063), .Z(n22065) );
  NAND U23686 ( .A(n22068), .B(n22067), .Z(n22072) );
  NAND U23687 ( .A(n22070), .B(n22069), .Z(n22071) );
  AND U23688 ( .A(n22072), .B(n22071), .Z(n22080) );
  NAND U23689 ( .A(n22074), .B(n22073), .Z(n22078) );
  NAND U23690 ( .A(n22076), .B(n22075), .Z(n22077) );
  NAND U23691 ( .A(n22078), .B(n22077), .Z(n22079) );
  XNOR U23692 ( .A(n22082), .B(n22081), .Z(n22083) );
  XNOR U23693 ( .A(n22084), .B(n22083), .Z(n22100) );
  NAND U23694 ( .A(n22086), .B(n22085), .Z(n22090) );
  NANDN U23695 ( .A(n22088), .B(n22087), .Z(n22089) );
  AND U23696 ( .A(n22090), .B(n22089), .Z(n22098) );
  NAND U23697 ( .A(n22094), .B(n22093), .Z(n22095) );
  NAND U23698 ( .A(n22096), .B(n22095), .Z(n22097) );
  XNOR U23699 ( .A(n22098), .B(n22097), .Z(n22099) );
  XNOR U23700 ( .A(n22100), .B(n22099), .Z(n22101) );
  XNOR U23701 ( .A(n22102), .B(n22101), .Z(n22118) );
  NAND U23702 ( .A(n22104), .B(n22103), .Z(n22108) );
  NANDN U23703 ( .A(n22106), .B(n22105), .Z(n22107) );
  AND U23704 ( .A(n22108), .B(n22107), .Z(n22116) );
  NAND U23705 ( .A(n22110), .B(n22109), .Z(n22114) );
  NAND U23706 ( .A(n22112), .B(n22111), .Z(n22113) );
  NAND U23707 ( .A(n22114), .B(n22113), .Z(n22115) );
  XNOR U23708 ( .A(n22116), .B(n22115), .Z(n22117) );
  XNOR U23709 ( .A(n22118), .B(n22117), .Z(n22119) );
  XNOR U23710 ( .A(n22120), .B(n22119), .Z(n22136) );
  OR U23711 ( .A(n22122), .B(n22121), .Z(n22126) );
  NAND U23712 ( .A(n22124), .B(n22123), .Z(n22125) );
  AND U23713 ( .A(n22126), .B(n22125), .Z(n22134) );
  NAND U23714 ( .A(n22128), .B(n22127), .Z(n22132) );
  NAND U23715 ( .A(n22130), .B(n22129), .Z(n22131) );
  NAND U23716 ( .A(n22132), .B(n22131), .Z(n22133) );
  XNOR U23717 ( .A(n22134), .B(n22133), .Z(n22135) );
  XNOR U23718 ( .A(n22136), .B(n22135), .Z(n22137) );
  XNOR U23719 ( .A(n22138), .B(n22137), .Z(n22154) );
  NANDN U23720 ( .A(n22140), .B(n22139), .Z(n22144) );
  NANDN U23721 ( .A(n22142), .B(n22141), .Z(n22143) );
  AND U23722 ( .A(n22144), .B(n22143), .Z(n22152) );
  NAND U23723 ( .A(n22146), .B(n22145), .Z(n22150) );
  NAND U23724 ( .A(n22148), .B(n22147), .Z(n22149) );
  NAND U23725 ( .A(n22150), .B(n22149), .Z(n22151) );
  XNOR U23726 ( .A(n22152), .B(n22151), .Z(n22153) );
  XNOR U23727 ( .A(n22154), .B(n22153), .Z(n22155) );
  XNOR U23728 ( .A(n22156), .B(n22155), .Z(n22164) );
  NAND U23729 ( .A(n22158), .B(n22157), .Z(n22162) );
  NANDN U23730 ( .A(n22160), .B(n22159), .Z(n22161) );
  NAND U23731 ( .A(n22162), .B(n22161), .Z(n22163) );
  XNOR U23732 ( .A(n22164), .B(n22163), .Z(N448) );
  AND U23733 ( .A(x[480]), .B(y[7904]), .Z(n22817) );
  XOR U23734 ( .A(n22817), .B(o[224]), .Z(N481) );
  AND U23735 ( .A(x[481]), .B(y[7904]), .Z(n22173) );
  AND U23736 ( .A(x[480]), .B(y[7905]), .Z(n22172) );
  XNOR U23737 ( .A(n22172), .B(o[225]), .Z(n22165) );
  XNOR U23738 ( .A(n22173), .B(n22165), .Z(n22167) );
  NAND U23739 ( .A(n22817), .B(o[224]), .Z(n22166) );
  XNOR U23740 ( .A(n22167), .B(n22166), .Z(N482) );
  NANDN U23741 ( .A(n22173), .B(n22165), .Z(n22169) );
  NAND U23742 ( .A(n22167), .B(n22166), .Z(n22168) );
  AND U23743 ( .A(n22169), .B(n22168), .Z(n22179) );
  AND U23744 ( .A(x[480]), .B(y[7906]), .Z(n22186) );
  XNOR U23745 ( .A(n22186), .B(o[226]), .Z(n22178) );
  XNOR U23746 ( .A(n22179), .B(n22178), .Z(n22181) );
  AND U23747 ( .A(y[7904]), .B(x[482]), .Z(n22171) );
  NAND U23748 ( .A(y[7905]), .B(x[481]), .Z(n22170) );
  XNOR U23749 ( .A(n22171), .B(n22170), .Z(n22175) );
  AND U23750 ( .A(n22172), .B(o[225]), .Z(n22174) );
  XNOR U23751 ( .A(n22175), .B(n22174), .Z(n22180) );
  XNOR U23752 ( .A(n22181), .B(n22180), .Z(N483) );
  AND U23753 ( .A(x[482]), .B(y[7905]), .Z(n22193) );
  NAND U23754 ( .A(n22193), .B(n22173), .Z(n22177) );
  NAND U23755 ( .A(n22175), .B(n22174), .Z(n22176) );
  AND U23756 ( .A(n22177), .B(n22176), .Z(n22196) );
  NANDN U23757 ( .A(n22179), .B(n22178), .Z(n22183) );
  NAND U23758 ( .A(n22181), .B(n22180), .Z(n22182) );
  AND U23759 ( .A(n22183), .B(n22182), .Z(n22195) );
  XNOR U23760 ( .A(n22196), .B(n22195), .Z(n22198) );
  AND U23761 ( .A(x[481]), .B(y[7906]), .Z(n22315) );
  XOR U23762 ( .A(n22193), .B(o[227]), .Z(n22201) );
  XOR U23763 ( .A(n22315), .B(n22201), .Z(n22203) );
  AND U23764 ( .A(y[7904]), .B(x[483]), .Z(n22185) );
  NAND U23765 ( .A(y[7907]), .B(x[480]), .Z(n22184) );
  XNOR U23766 ( .A(n22185), .B(n22184), .Z(n22188) );
  AND U23767 ( .A(n22186), .B(o[226]), .Z(n22187) );
  XOR U23768 ( .A(n22188), .B(n22187), .Z(n22202) );
  XOR U23769 ( .A(n22203), .B(n22202), .Z(n22197) );
  XOR U23770 ( .A(n22198), .B(n22197), .Z(N484) );
  AND U23771 ( .A(x[483]), .B(y[7907]), .Z(n22246) );
  NAND U23772 ( .A(n22817), .B(n22246), .Z(n22190) );
  NAND U23773 ( .A(n22188), .B(n22187), .Z(n22189) );
  NAND U23774 ( .A(n22190), .B(n22189), .Z(n22224) );
  AND U23775 ( .A(y[7908]), .B(x[480]), .Z(n22192) );
  NAND U23776 ( .A(y[7904]), .B(x[484]), .Z(n22191) );
  XNOR U23777 ( .A(n22192), .B(n22191), .Z(n22217) );
  NAND U23778 ( .A(n22193), .B(o[227]), .Z(n22218) );
  AND U23779 ( .A(y[7906]), .B(x[482]), .Z(n22369) );
  NAND U23780 ( .A(y[7907]), .B(x[481]), .Z(n22194) );
  XNOR U23781 ( .A(n22369), .B(n22194), .Z(n22214) );
  AND U23782 ( .A(x[483]), .B(y[7905]), .Z(n22209) );
  XOR U23783 ( .A(o[228]), .B(n22209), .Z(n22213) );
  XOR U23784 ( .A(n22214), .B(n22213), .Z(n22221) );
  XOR U23785 ( .A(n22222), .B(n22221), .Z(n22223) );
  XOR U23786 ( .A(n22224), .B(n22223), .Z(n22228) );
  NANDN U23787 ( .A(n22196), .B(n22195), .Z(n22200) );
  NAND U23788 ( .A(n22198), .B(n22197), .Z(n22199) );
  NAND U23789 ( .A(n22200), .B(n22199), .Z(n22229) );
  NAND U23790 ( .A(n22315), .B(n22201), .Z(n22205) );
  NAND U23791 ( .A(n22203), .B(n22202), .Z(n22204) );
  NAND U23792 ( .A(n22205), .B(n22204), .Z(n22230) );
  IV U23793 ( .A(n22230), .Z(n22227) );
  XOR U23794 ( .A(n22229), .B(n22227), .Z(n22206) );
  XNOR U23795 ( .A(n22228), .B(n22206), .Z(N485) );
  AND U23796 ( .A(y[7906]), .B(x[483]), .Z(n22208) );
  NAND U23797 ( .A(y[7908]), .B(x[481]), .Z(n22207) );
  XNOR U23798 ( .A(n22208), .B(n22207), .Z(n22233) );
  AND U23799 ( .A(x[484]), .B(y[7905]), .Z(n22244) );
  XOR U23800 ( .A(n22244), .B(o[229]), .Z(n22232) );
  XNOR U23801 ( .A(n22233), .B(n22232), .Z(n22236) );
  NAND U23802 ( .A(x[482]), .B(y[7907]), .Z(n22324) );
  AND U23803 ( .A(o[228]), .B(n22209), .Z(n22238) );
  AND U23804 ( .A(y[7904]), .B(x[485]), .Z(n22211) );
  NAND U23805 ( .A(y[7909]), .B(x[480]), .Z(n22210) );
  XNOR U23806 ( .A(n22211), .B(n22210), .Z(n22239) );
  XOR U23807 ( .A(n22238), .B(n22239), .Z(n22237) );
  XOR U23808 ( .A(n22324), .B(n22237), .Z(n22212) );
  XOR U23809 ( .A(n22236), .B(n22212), .Z(n22254) );
  NANDN U23810 ( .A(n22324), .B(n22315), .Z(n22216) );
  NAND U23811 ( .A(n22214), .B(n22213), .Z(n22215) );
  AND U23812 ( .A(n22216), .B(n22215), .Z(n22252) );
  AND U23813 ( .A(x[484]), .B(y[7908]), .Z(n23020) );
  NAND U23814 ( .A(n23020), .B(n22817), .Z(n22220) );
  NANDN U23815 ( .A(n22218), .B(n22217), .Z(n22219) );
  NAND U23816 ( .A(n22220), .B(n22219), .Z(n22251) );
  XNOR U23817 ( .A(n22254), .B(n22253), .Z(n22250) );
  NAND U23818 ( .A(n22222), .B(n22221), .Z(n22226) );
  NAND U23819 ( .A(n22224), .B(n22223), .Z(n22225) );
  NAND U23820 ( .A(n22226), .B(n22225), .Z(n22249) );
  XOR U23821 ( .A(n22249), .B(n22248), .Z(n22231) );
  XNOR U23822 ( .A(n22250), .B(n22231), .Z(N486) );
  AND U23823 ( .A(x[483]), .B(y[7908]), .Z(n22325) );
  NAND U23824 ( .A(n22325), .B(n22315), .Z(n22235) );
  NAND U23825 ( .A(n22233), .B(n22232), .Z(n22234) );
  NAND U23826 ( .A(n22235), .B(n22234), .Z(n22290) );
  XOR U23827 ( .A(n22290), .B(n22289), .Z(n22292) );
  AND U23828 ( .A(x[485]), .B(y[7909]), .Z(n22493) );
  NAND U23829 ( .A(n22817), .B(n22493), .Z(n22241) );
  NAND U23830 ( .A(n22239), .B(n22238), .Z(n22240) );
  NAND U23831 ( .A(n22241), .B(n22240), .Z(n22259) );
  AND U23832 ( .A(y[7904]), .B(x[486]), .Z(n22243) );
  NAND U23833 ( .A(y[7910]), .B(x[480]), .Z(n22242) );
  XNOR U23834 ( .A(n22243), .B(n22242), .Z(n22265) );
  AND U23835 ( .A(n22244), .B(o[229]), .Z(n22266) );
  XOR U23836 ( .A(n22265), .B(n22266), .Z(n22258) );
  XOR U23837 ( .A(n22259), .B(n22258), .Z(n22261) );
  NAND U23838 ( .A(y[7908]), .B(x[482]), .Z(n22245) );
  XNOR U23839 ( .A(n22246), .B(n22245), .Z(n22270) );
  AND U23840 ( .A(y[7909]), .B(x[481]), .Z(n22531) );
  NAND U23841 ( .A(y[7906]), .B(x[484]), .Z(n22247) );
  XNOR U23842 ( .A(n22531), .B(n22247), .Z(n22274) );
  AND U23843 ( .A(x[485]), .B(y[7905]), .Z(n22281) );
  XOR U23844 ( .A(o[230]), .B(n22281), .Z(n22273) );
  XOR U23845 ( .A(n22274), .B(n22273), .Z(n22269) );
  XOR U23846 ( .A(n22270), .B(n22269), .Z(n22260) );
  XOR U23847 ( .A(n22261), .B(n22260), .Z(n22291) );
  XNOR U23848 ( .A(n22292), .B(n22291), .Z(n22285) );
  NANDN U23849 ( .A(n22252), .B(n22251), .Z(n22256) );
  NAND U23850 ( .A(n22254), .B(n22253), .Z(n22255) );
  NAND U23851 ( .A(n22256), .B(n22255), .Z(n22283) );
  IV U23852 ( .A(n22283), .Z(n22282) );
  XOR U23853 ( .A(n22284), .B(n22282), .Z(n22257) );
  XNOR U23854 ( .A(n22285), .B(n22257), .Z(N487) );
  NAND U23855 ( .A(n22259), .B(n22258), .Z(n22263) );
  NAND U23856 ( .A(n22261), .B(n22260), .Z(n22262) );
  AND U23857 ( .A(n22263), .B(n22262), .Z(n22299) );
  AND U23858 ( .A(y[7906]), .B(x[485]), .Z(n22392) );
  NAND U23859 ( .A(y[7910]), .B(x[481]), .Z(n22264) );
  XNOR U23860 ( .A(n22392), .B(n22264), .Z(n22317) );
  AND U23861 ( .A(x[486]), .B(y[7905]), .Z(n22321) );
  XOR U23862 ( .A(o[231]), .B(n22321), .Z(n22316) );
  XNOR U23863 ( .A(n22317), .B(n22316), .Z(n22336) );
  AND U23864 ( .A(x[486]), .B(y[7910]), .Z(n22551) );
  NAND U23865 ( .A(n22817), .B(n22551), .Z(n22268) );
  NAND U23866 ( .A(n22266), .B(n22265), .Z(n22267) );
  AND U23867 ( .A(n22268), .B(n22267), .Z(n22335) );
  XOR U23868 ( .A(n22336), .B(n22335), .Z(n22337) );
  NANDN U23869 ( .A(n22324), .B(n22325), .Z(n22272) );
  NAND U23870 ( .A(n22270), .B(n22269), .Z(n22271) );
  AND U23871 ( .A(n22272), .B(n22271), .Z(n22338) );
  XOR U23872 ( .A(n22337), .B(n22338), .Z(n22297) );
  AND U23873 ( .A(x[484]), .B(y[7909]), .Z(n22822) );
  NAND U23874 ( .A(n22822), .B(n22315), .Z(n22276) );
  NAND U23875 ( .A(n22274), .B(n22273), .Z(n22275) );
  AND U23876 ( .A(n22276), .B(n22275), .Z(n22312) );
  AND U23877 ( .A(y[7909]), .B(x[482]), .Z(n22278) );
  NAND U23878 ( .A(y[7907]), .B(x[484]), .Z(n22277) );
  XNOR U23879 ( .A(n22278), .B(n22277), .Z(n22326) );
  XNOR U23880 ( .A(n22326), .B(n22325), .Z(n22310) );
  AND U23881 ( .A(y[7904]), .B(x[487]), .Z(n22280) );
  NAND U23882 ( .A(y[7911]), .B(x[480]), .Z(n22279) );
  XNOR U23883 ( .A(n22280), .B(n22279), .Z(n22330) );
  AND U23884 ( .A(o[230]), .B(n22281), .Z(n22329) );
  XNOR U23885 ( .A(n22330), .B(n22329), .Z(n22309) );
  XOR U23886 ( .A(n22310), .B(n22309), .Z(n22311) );
  XOR U23887 ( .A(n22312), .B(n22311), .Z(n22296) );
  XOR U23888 ( .A(n22297), .B(n22296), .Z(n22298) );
  XNOR U23889 ( .A(n22299), .B(n22298), .Z(n22305) );
  OR U23890 ( .A(n22284), .B(n22282), .Z(n22288) );
  ANDN U23891 ( .B(n22284), .A(n22283), .Z(n22286) );
  OR U23892 ( .A(n22286), .B(n22285), .Z(n22287) );
  AND U23893 ( .A(n22288), .B(n22287), .Z(n22303) );
  NAND U23894 ( .A(n22290), .B(n22289), .Z(n22294) );
  NAND U23895 ( .A(n22292), .B(n22291), .Z(n22293) );
  AND U23896 ( .A(n22294), .B(n22293), .Z(n22304) );
  IV U23897 ( .A(n22304), .Z(n22302) );
  XOR U23898 ( .A(n22303), .B(n22302), .Z(n22295) );
  XNOR U23899 ( .A(n22305), .B(n22295), .Z(N488) );
  NAND U23900 ( .A(n22297), .B(n22296), .Z(n22301) );
  NAND U23901 ( .A(n22299), .B(n22298), .Z(n22300) );
  AND U23902 ( .A(n22301), .B(n22300), .Z(n22349) );
  NANDN U23903 ( .A(n22302), .B(n22303), .Z(n22308) );
  NOR U23904 ( .A(n22304), .B(n22303), .Z(n22306) );
  OR U23905 ( .A(n22306), .B(n22305), .Z(n22307) );
  AND U23906 ( .A(n22308), .B(n22307), .Z(n22348) );
  NAND U23907 ( .A(n22310), .B(n22309), .Z(n22314) );
  NAND U23908 ( .A(n22312), .B(n22311), .Z(n22313) );
  AND U23909 ( .A(n22314), .B(n22313), .Z(n22382) );
  AND U23910 ( .A(x[485]), .B(y[7910]), .Z(n22485) );
  NAND U23911 ( .A(n22485), .B(n22315), .Z(n22319) );
  NAND U23912 ( .A(n22317), .B(n22316), .Z(n22318) );
  NAND U23913 ( .A(n22319), .B(n22318), .Z(n22380) );
  AND U23914 ( .A(y[7907]), .B(x[485]), .Z(n22926) );
  NAND U23915 ( .A(y[7911]), .B(x[481]), .Z(n22320) );
  XNOR U23916 ( .A(n22926), .B(n22320), .Z(n22363) );
  AND U23917 ( .A(o[231]), .B(n22321), .Z(n22362) );
  XOR U23918 ( .A(n22363), .B(n22362), .Z(n22368) );
  NAND U23919 ( .A(x[483]), .B(y[7909]), .Z(n23156) );
  AND U23920 ( .A(y[7906]), .B(x[486]), .Z(n22323) );
  NAND U23921 ( .A(y[7910]), .B(x[482]), .Z(n22322) );
  XNOR U23922 ( .A(n22323), .B(n22322), .Z(n22370) );
  XNOR U23923 ( .A(n23020), .B(n22370), .Z(n22366) );
  XOR U23924 ( .A(n23156), .B(n22366), .Z(n22367) );
  XOR U23925 ( .A(n22368), .B(n22367), .Z(n22379) );
  XOR U23926 ( .A(n22380), .B(n22379), .Z(n22381) );
  XNOR U23927 ( .A(n22382), .B(n22381), .Z(n22345) );
  NANDN U23928 ( .A(n22324), .B(n22822), .Z(n22328) );
  NAND U23929 ( .A(n22326), .B(n22325), .Z(n22327) );
  NAND U23930 ( .A(n22328), .B(n22327), .Z(n22376) );
  AND U23931 ( .A(x[487]), .B(y[7911]), .Z(n22694) );
  NAND U23932 ( .A(n22817), .B(n22694), .Z(n22332) );
  NAND U23933 ( .A(n22330), .B(n22329), .Z(n22331) );
  NAND U23934 ( .A(n22332), .B(n22331), .Z(n22374) );
  AND U23935 ( .A(y[7904]), .B(x[488]), .Z(n22334) );
  NAND U23936 ( .A(y[7912]), .B(x[480]), .Z(n22333) );
  XNOR U23937 ( .A(n22334), .B(n22333), .Z(n22353) );
  AND U23938 ( .A(x[487]), .B(y[7905]), .Z(n22358) );
  XOR U23939 ( .A(o[232]), .B(n22358), .Z(n22352) );
  XOR U23940 ( .A(n22353), .B(n22352), .Z(n22373) );
  XOR U23941 ( .A(n22374), .B(n22373), .Z(n22375) );
  XNOR U23942 ( .A(n22376), .B(n22375), .Z(n22343) );
  NAND U23943 ( .A(n22336), .B(n22335), .Z(n22340) );
  NAND U23944 ( .A(n22338), .B(n22337), .Z(n22339) );
  NAND U23945 ( .A(n22340), .B(n22339), .Z(n22342) );
  XOR U23946 ( .A(n22343), .B(n22342), .Z(n22344) );
  XOR U23947 ( .A(n22345), .B(n22344), .Z(n22350) );
  XNOR U23948 ( .A(n22348), .B(n22350), .Z(n22341) );
  XOR U23949 ( .A(n22349), .B(n22341), .Z(N489) );
  NAND U23950 ( .A(n22343), .B(n22342), .Z(n22347) );
  NAND U23951 ( .A(n22345), .B(n22344), .Z(n22346) );
  NAND U23952 ( .A(n22347), .B(n22346), .Z(n22436) );
  IV U23953 ( .A(n22436), .Z(n22434) );
  AND U23954 ( .A(x[488]), .B(y[7912]), .Z(n22351) );
  NAND U23955 ( .A(n22351), .B(n22817), .Z(n22355) );
  NAND U23956 ( .A(n22353), .B(n22352), .Z(n22354) );
  AND U23957 ( .A(n22355), .B(n22354), .Z(n22421) );
  AND U23958 ( .A(y[7908]), .B(x[485]), .Z(n22357) );
  NAND U23959 ( .A(y[7906]), .B(x[487]), .Z(n22356) );
  XNOR U23960 ( .A(n22357), .B(n22356), .Z(n22394) );
  AND U23961 ( .A(o[232]), .B(n22358), .Z(n22393) );
  XNOR U23962 ( .A(n22394), .B(n22393), .Z(n22419) );
  AND U23963 ( .A(y[7904]), .B(x[489]), .Z(n22360) );
  NAND U23964 ( .A(y[7913]), .B(x[480]), .Z(n22359) );
  XNOR U23965 ( .A(n22360), .B(n22359), .Z(n22401) );
  AND U23966 ( .A(x[488]), .B(y[7905]), .Z(n22410) );
  XOR U23967 ( .A(o[233]), .B(n22410), .Z(n22400) );
  XNOR U23968 ( .A(n22401), .B(n22400), .Z(n22418) );
  XOR U23969 ( .A(n22419), .B(n22418), .Z(n22420) );
  XNOR U23970 ( .A(n22421), .B(n22420), .Z(n22415) );
  AND U23971 ( .A(y[7907]), .B(x[486]), .Z(n22765) );
  NAND U23972 ( .A(y[7912]), .B(x[481]), .Z(n22361) );
  XNOR U23973 ( .A(n22765), .B(n22361), .Z(n22405) );
  XNOR U23974 ( .A(n22822), .B(n22405), .Z(n22425) );
  NAND U23975 ( .A(x[482]), .B(y[7911]), .Z(n23067) );
  AND U23976 ( .A(x[483]), .B(y[7910]), .Z(n22775) );
  XNOR U23977 ( .A(n23067), .B(n22775), .Z(n22424) );
  XNOR U23978 ( .A(n22425), .B(n22424), .Z(n22413) );
  NAND U23979 ( .A(x[485]), .B(y[7911]), .Z(n22601) );
  AND U23980 ( .A(x[481]), .B(y[7907]), .Z(n22404) );
  NANDN U23981 ( .A(n22601), .B(n22404), .Z(n22365) );
  NAND U23982 ( .A(n22363), .B(n22362), .Z(n22364) );
  NAND U23983 ( .A(n22365), .B(n22364), .Z(n22412) );
  XOR U23984 ( .A(n22413), .B(n22412), .Z(n22414) );
  XNOR U23985 ( .A(n22415), .B(n22414), .Z(n22388) );
  NAND U23986 ( .A(n22551), .B(n22369), .Z(n22372) );
  NAND U23987 ( .A(n23020), .B(n22370), .Z(n22371) );
  AND U23988 ( .A(n22372), .B(n22371), .Z(n22386) );
  XOR U23989 ( .A(n22387), .B(n22386), .Z(n22389) );
  XNOR U23990 ( .A(n22388), .B(n22389), .Z(n22430) );
  NAND U23991 ( .A(n22374), .B(n22373), .Z(n22378) );
  NAND U23992 ( .A(n22376), .B(n22375), .Z(n22377) );
  NAND U23993 ( .A(n22378), .B(n22377), .Z(n22429) );
  NAND U23994 ( .A(n22380), .B(n22379), .Z(n22384) );
  NAND U23995 ( .A(n22382), .B(n22381), .Z(n22383) );
  NAND U23996 ( .A(n22384), .B(n22383), .Z(n22428) );
  XOR U23997 ( .A(n22429), .B(n22428), .Z(n22431) );
  XOR U23998 ( .A(n22430), .B(n22431), .Z(n22437) );
  XNOR U23999 ( .A(n22435), .B(n22437), .Z(n22385) );
  XOR U24000 ( .A(n22434), .B(n22385), .Z(N490) );
  NAND U24001 ( .A(n22387), .B(n22386), .Z(n22391) );
  NAND U24002 ( .A(n22389), .B(n22388), .Z(n22390) );
  NAND U24003 ( .A(n22391), .B(n22390), .Z(n22445) );
  AND U24004 ( .A(x[487]), .B(y[7908]), .Z(n22487) );
  NAND U24005 ( .A(n22487), .B(n22392), .Z(n22396) );
  NAND U24006 ( .A(n22394), .B(n22393), .Z(n22395) );
  AND U24007 ( .A(n22396), .B(n22395), .Z(n22500) );
  AND U24008 ( .A(y[7907]), .B(x[487]), .Z(n22398) );
  NAND U24009 ( .A(y[7910]), .B(x[484]), .Z(n22397) );
  XNOR U24010 ( .A(n22398), .B(n22397), .Z(n22471) );
  AND U24011 ( .A(x[486]), .B(y[7908]), .Z(n22470) );
  XNOR U24012 ( .A(n22471), .B(n22470), .Z(n22498) );
  AND U24013 ( .A(x[488]), .B(y[7906]), .Z(n22658) );
  AND U24014 ( .A(x[489]), .B(y[7905]), .Z(n22481) );
  XOR U24015 ( .A(o[234]), .B(n22481), .Z(n22492) );
  XOR U24016 ( .A(n22658), .B(n22492), .Z(n22494) );
  XNOR U24017 ( .A(n22494), .B(n22493), .Z(n22497) );
  XOR U24018 ( .A(n22498), .B(n22497), .Z(n22499) );
  XNOR U24019 ( .A(n22500), .B(n22499), .Z(n22460) );
  AND U24020 ( .A(x[489]), .B(y[7913]), .Z(n22399) );
  NAND U24021 ( .A(n22399), .B(n22817), .Z(n22403) );
  NAND U24022 ( .A(n22401), .B(n22400), .Z(n22402) );
  NAND U24023 ( .A(n22403), .B(n22402), .Z(n22458) );
  AND U24024 ( .A(x[486]), .B(y[7912]), .Z(n22685) );
  NAND U24025 ( .A(n22685), .B(n22404), .Z(n22407) );
  NAND U24026 ( .A(n22822), .B(n22405), .Z(n22406) );
  NAND U24027 ( .A(n22407), .B(n22406), .Z(n22466) );
  AND U24028 ( .A(y[7904]), .B(x[490]), .Z(n22409) );
  NAND U24029 ( .A(y[7914]), .B(x[480]), .Z(n22408) );
  XNOR U24030 ( .A(n22409), .B(n22408), .Z(n22476) );
  AND U24031 ( .A(o[233]), .B(n22410), .Z(n22475) );
  XOR U24032 ( .A(n22476), .B(n22475), .Z(n22464) );
  AND U24033 ( .A(y[7911]), .B(x[483]), .Z(n23409) );
  NAND U24034 ( .A(y[7913]), .B(x[481]), .Z(n22411) );
  XNOR U24035 ( .A(n23409), .B(n22411), .Z(n22488) );
  AND U24036 ( .A(x[482]), .B(y[7912]), .Z(n22489) );
  XOR U24037 ( .A(n22488), .B(n22489), .Z(n22463) );
  XOR U24038 ( .A(n22464), .B(n22463), .Z(n22465) );
  XOR U24039 ( .A(n22466), .B(n22465), .Z(n22457) );
  XOR U24040 ( .A(n22458), .B(n22457), .Z(n22459) );
  XNOR U24041 ( .A(n22460), .B(n22459), .Z(n22443) );
  NAND U24042 ( .A(n22413), .B(n22412), .Z(n22417) );
  NAND U24043 ( .A(n22415), .B(n22414), .Z(n22416) );
  AND U24044 ( .A(n22417), .B(n22416), .Z(n22454) );
  NAND U24045 ( .A(n22419), .B(n22418), .Z(n22423) );
  NAND U24046 ( .A(n22421), .B(n22420), .Z(n22422) );
  AND U24047 ( .A(n22423), .B(n22422), .Z(n22451) );
  NAND U24048 ( .A(n22425), .B(n22424), .Z(n22427) );
  ANDN U24049 ( .B(n23067), .A(n22775), .Z(n22426) );
  ANDN U24050 ( .B(n22427), .A(n22426), .Z(n22452) );
  XOR U24051 ( .A(n22451), .B(n22452), .Z(n22453) );
  XOR U24052 ( .A(n22454), .B(n22453), .Z(n22442) );
  XOR U24053 ( .A(n22443), .B(n22442), .Z(n22444) );
  XOR U24054 ( .A(n22445), .B(n22444), .Z(n22450) );
  NAND U24055 ( .A(n22429), .B(n22428), .Z(n22433) );
  NAND U24056 ( .A(n22431), .B(n22430), .Z(n22432) );
  NAND U24057 ( .A(n22433), .B(n22432), .Z(n22449) );
  NANDN U24058 ( .A(n22434), .B(n22435), .Z(n22440) );
  NOR U24059 ( .A(n22436), .B(n22435), .Z(n22438) );
  OR U24060 ( .A(n22438), .B(n22437), .Z(n22439) );
  AND U24061 ( .A(n22440), .B(n22439), .Z(n22448) );
  XOR U24062 ( .A(n22449), .B(n22448), .Z(n22441) );
  XNOR U24063 ( .A(n22450), .B(n22441), .Z(N491) );
  NAND U24064 ( .A(n22443), .B(n22442), .Z(n22447) );
  NAND U24065 ( .A(n22445), .B(n22444), .Z(n22446) );
  NAND U24066 ( .A(n22447), .B(n22446), .Z(n22567) );
  IV U24067 ( .A(n22567), .Z(n22565) );
  NAND U24068 ( .A(n22452), .B(n22451), .Z(n22456) );
  NANDN U24069 ( .A(n22454), .B(n22453), .Z(n22455) );
  NAND U24070 ( .A(n22456), .B(n22455), .Z(n22562) );
  NAND U24071 ( .A(n22458), .B(n22457), .Z(n22462) );
  NAND U24072 ( .A(n22460), .B(n22459), .Z(n22461) );
  NAND U24073 ( .A(n22462), .B(n22461), .Z(n22560) );
  NAND U24074 ( .A(n22464), .B(n22463), .Z(n22468) );
  NAND U24075 ( .A(n22466), .B(n22465), .Z(n22467) );
  NAND U24076 ( .A(n22468), .B(n22467), .Z(n22518) );
  AND U24077 ( .A(x[487]), .B(y[7910]), .Z(n22596) );
  AND U24078 ( .A(x[484]), .B(y[7907]), .Z(n22469) );
  NAND U24079 ( .A(n22596), .B(n22469), .Z(n22473) );
  NAND U24080 ( .A(n22471), .B(n22470), .Z(n22472) );
  NAND U24081 ( .A(n22473), .B(n22472), .Z(n22516) );
  AND U24082 ( .A(x[490]), .B(y[7914]), .Z(n22474) );
  NAND U24083 ( .A(n22474), .B(n22817), .Z(n22478) );
  NAND U24084 ( .A(n22476), .B(n22475), .Z(n22477) );
  NAND U24085 ( .A(n22478), .B(n22477), .Z(n22512) );
  AND U24086 ( .A(y[7904]), .B(x[491]), .Z(n22480) );
  NAND U24087 ( .A(y[7915]), .B(x[480]), .Z(n22479) );
  XNOR U24088 ( .A(n22480), .B(n22479), .Z(n22542) );
  AND U24089 ( .A(o[234]), .B(n22481), .Z(n22541) );
  XOR U24090 ( .A(n22542), .B(n22541), .Z(n22510) );
  AND U24091 ( .A(y[7909]), .B(x[486]), .Z(n22483) );
  NAND U24092 ( .A(y[7914]), .B(x[481]), .Z(n22482) );
  XNOR U24093 ( .A(n22483), .B(n22482), .Z(n22533) );
  AND U24094 ( .A(x[490]), .B(y[7905]), .Z(n22552) );
  XOR U24095 ( .A(o[235]), .B(n22552), .Z(n22532) );
  XOR U24096 ( .A(n22533), .B(n22532), .Z(n22509) );
  XOR U24097 ( .A(n22510), .B(n22509), .Z(n22511) );
  XOR U24098 ( .A(n22512), .B(n22511), .Z(n22515) );
  XOR U24099 ( .A(n22516), .B(n22515), .Z(n22517) );
  XNOR U24100 ( .A(n22518), .B(n22517), .Z(n22555) );
  AND U24101 ( .A(x[483]), .B(y[7912]), .Z(n23529) );
  NAND U24102 ( .A(y[7913]), .B(x[482]), .Z(n22484) );
  XNOR U24103 ( .A(n22485), .B(n22484), .Z(n22528) );
  AND U24104 ( .A(x[484]), .B(y[7911]), .Z(n22527) );
  XNOR U24105 ( .A(n22528), .B(n22527), .Z(n22504) );
  XNOR U24106 ( .A(n23529), .B(n22504), .Z(n22506) );
  NAND U24107 ( .A(y[7906]), .B(x[489]), .Z(n22486) );
  XNOR U24108 ( .A(n22487), .B(n22486), .Z(n22547) );
  AND U24109 ( .A(x[488]), .B(y[7907]), .Z(n22546) );
  XNOR U24110 ( .A(n22547), .B(n22546), .Z(n22505) );
  XNOR U24111 ( .A(n22506), .B(n22505), .Z(n22524) );
  NAND U24112 ( .A(x[483]), .B(y[7913]), .Z(n22592) );
  AND U24113 ( .A(x[481]), .B(y[7911]), .Z(n22812) );
  NANDN U24114 ( .A(n22592), .B(n22812), .Z(n22491) );
  NAND U24115 ( .A(n22489), .B(n22488), .Z(n22490) );
  NAND U24116 ( .A(n22491), .B(n22490), .Z(n22522) );
  NAND U24117 ( .A(n22658), .B(n22492), .Z(n22496) );
  NAND U24118 ( .A(n22494), .B(n22493), .Z(n22495) );
  NAND U24119 ( .A(n22496), .B(n22495), .Z(n22521) );
  XOR U24120 ( .A(n22522), .B(n22521), .Z(n22523) );
  XNOR U24121 ( .A(n22524), .B(n22523), .Z(n22554) );
  NAND U24122 ( .A(n22498), .B(n22497), .Z(n22502) );
  NAND U24123 ( .A(n22500), .B(n22499), .Z(n22501) );
  NAND U24124 ( .A(n22502), .B(n22501), .Z(n22553) );
  XOR U24125 ( .A(n22554), .B(n22553), .Z(n22556) );
  XNOR U24126 ( .A(n22555), .B(n22556), .Z(n22559) );
  XOR U24127 ( .A(n22560), .B(n22559), .Z(n22561) );
  XOR U24128 ( .A(n22562), .B(n22561), .Z(n22568) );
  XNOR U24129 ( .A(n22566), .B(n22568), .Z(n22503) );
  XOR U24130 ( .A(n22565), .B(n22503), .Z(N492) );
  NANDN U24131 ( .A(n23529), .B(n22504), .Z(n22508) );
  NAND U24132 ( .A(n22506), .B(n22505), .Z(n22507) );
  NAND U24133 ( .A(n22508), .B(n22507), .Z(n22574) );
  NAND U24134 ( .A(n22510), .B(n22509), .Z(n22514) );
  NAND U24135 ( .A(n22512), .B(n22511), .Z(n22513) );
  AND U24136 ( .A(n22514), .B(n22513), .Z(n22573) );
  XOR U24137 ( .A(n22574), .B(n22573), .Z(n22575) );
  NAND U24138 ( .A(n22516), .B(n22515), .Z(n22520) );
  NAND U24139 ( .A(n22518), .B(n22517), .Z(n22519) );
  AND U24140 ( .A(n22520), .B(n22519), .Z(n22576) );
  XOR U24141 ( .A(n22575), .B(n22576), .Z(n22642) );
  NAND U24142 ( .A(n22522), .B(n22521), .Z(n22526) );
  NAND U24143 ( .A(n22524), .B(n22523), .Z(n22525) );
  NAND U24144 ( .A(n22526), .B(n22525), .Z(n22633) );
  AND U24145 ( .A(x[482]), .B(y[7910]), .Z(n23254) );
  AND U24146 ( .A(x[485]), .B(y[7913]), .Z(n23058) );
  NAND U24147 ( .A(n23254), .B(n23058), .Z(n22530) );
  NAND U24148 ( .A(n22528), .B(n22527), .Z(n22529) );
  NAND U24149 ( .A(n22530), .B(n22529), .Z(n22580) );
  AND U24150 ( .A(x[486]), .B(y[7914]), .Z(n22829) );
  NAND U24151 ( .A(n22829), .B(n22531), .Z(n22535) );
  NAND U24152 ( .A(n22533), .B(n22532), .Z(n22534) );
  NAND U24153 ( .A(n22535), .B(n22534), .Z(n22579) );
  XOR U24154 ( .A(n22580), .B(n22579), .Z(n22582) );
  AND U24155 ( .A(x[489]), .B(y[7907]), .Z(n23249) );
  AND U24156 ( .A(x[490]), .B(y[7906]), .Z(n23291) );
  AND U24157 ( .A(y[7912]), .B(x[484]), .Z(n22536) );
  XOR U24158 ( .A(n23291), .B(n22536), .Z(n22623) );
  XOR U24159 ( .A(n23249), .B(n22623), .Z(n22602) );
  NAND U24160 ( .A(x[487]), .B(y[7909]), .Z(n22600) );
  XOR U24161 ( .A(n22601), .B(n22600), .Z(n22603) );
  AND U24162 ( .A(y[7904]), .B(x[492]), .Z(n22538) );
  NAND U24163 ( .A(y[7916]), .B(x[480]), .Z(n22537) );
  XNOR U24164 ( .A(n22538), .B(n22537), .Z(n22617) );
  AND U24165 ( .A(x[491]), .B(y[7905]), .Z(n22597) );
  XOR U24166 ( .A(o[236]), .B(n22597), .Z(n22616) );
  XOR U24167 ( .A(n22617), .B(n22616), .Z(n22586) );
  AND U24168 ( .A(y[7914]), .B(x[482]), .Z(n22540) );
  NAND U24169 ( .A(y[7908]), .B(x[488]), .Z(n22539) );
  XNOR U24170 ( .A(n22540), .B(n22539), .Z(n22591) );
  XOR U24171 ( .A(n22586), .B(n22585), .Z(n22588) );
  XOR U24172 ( .A(n22587), .B(n22588), .Z(n22581) );
  XOR U24173 ( .A(n22582), .B(n22581), .Z(n22631) );
  AND U24174 ( .A(x[491]), .B(y[7915]), .Z(n23652) );
  NAND U24175 ( .A(n23652), .B(n22817), .Z(n22544) );
  NAND U24176 ( .A(n22542), .B(n22541), .Z(n22543) );
  NAND U24177 ( .A(n22544), .B(n22543), .Z(n22609) );
  AND U24178 ( .A(x[487]), .B(y[7906]), .Z(n22751) );
  AND U24179 ( .A(x[489]), .B(y[7908]), .Z(n22545) );
  NAND U24180 ( .A(n22751), .B(n22545), .Z(n22549) );
  NAND U24181 ( .A(n22547), .B(n22546), .Z(n22548) );
  NAND U24182 ( .A(n22549), .B(n22548), .Z(n22607) );
  NAND U24183 ( .A(y[7915]), .B(x[481]), .Z(n22550) );
  XNOR U24184 ( .A(n22551), .B(n22550), .Z(n22613) );
  AND U24185 ( .A(o[235]), .B(n22552), .Z(n22612) );
  XOR U24186 ( .A(n22613), .B(n22612), .Z(n22606) );
  XOR U24187 ( .A(n22607), .B(n22606), .Z(n22608) );
  XOR U24188 ( .A(n22609), .B(n22608), .Z(n22630) );
  XOR U24189 ( .A(n22631), .B(n22630), .Z(n22632) );
  XNOR U24190 ( .A(n22633), .B(n22632), .Z(n22640) );
  NAND U24191 ( .A(n22554), .B(n22553), .Z(n22558) );
  NAND U24192 ( .A(n22556), .B(n22555), .Z(n22557) );
  NAND U24193 ( .A(n22558), .B(n22557), .Z(n22639) );
  XOR U24194 ( .A(n22640), .B(n22639), .Z(n22641) );
  XOR U24195 ( .A(n22642), .B(n22641), .Z(n22638) );
  NAND U24196 ( .A(n22560), .B(n22559), .Z(n22564) );
  NAND U24197 ( .A(n22562), .B(n22561), .Z(n22563) );
  NAND U24198 ( .A(n22564), .B(n22563), .Z(n22637) );
  NANDN U24199 ( .A(n22565), .B(n22566), .Z(n22571) );
  NOR U24200 ( .A(n22567), .B(n22566), .Z(n22569) );
  OR U24201 ( .A(n22569), .B(n22568), .Z(n22570) );
  AND U24202 ( .A(n22571), .B(n22570), .Z(n22636) );
  XOR U24203 ( .A(n22637), .B(n22636), .Z(n22572) );
  XNOR U24204 ( .A(n22638), .B(n22572), .Z(N493) );
  NAND U24205 ( .A(n22574), .B(n22573), .Z(n22578) );
  NAND U24206 ( .A(n22576), .B(n22575), .Z(n22577) );
  AND U24207 ( .A(n22578), .B(n22577), .Z(n22723) );
  NAND U24208 ( .A(n22580), .B(n22579), .Z(n22584) );
  NAND U24209 ( .A(n22582), .B(n22581), .Z(n22583) );
  AND U24210 ( .A(n22584), .B(n22583), .Z(n22702) );
  NAND U24211 ( .A(n22586), .B(n22585), .Z(n22590) );
  NAND U24212 ( .A(n22588), .B(n22587), .Z(n22589) );
  NAND U24213 ( .A(n22590), .B(n22589), .Z(n22709) );
  AND U24214 ( .A(y[7914]), .B(x[488]), .Z(n23908) );
  AND U24215 ( .A(x[482]), .B(y[7908]), .Z(n22761) );
  NAND U24216 ( .A(n23908), .B(n22761), .Z(n22594) );
  NANDN U24217 ( .A(n22592), .B(n22591), .Z(n22593) );
  NAND U24218 ( .A(n22594), .B(n22593), .Z(n22673) );
  NAND U24219 ( .A(y[7916]), .B(x[481]), .Z(n22595) );
  XNOR U24220 ( .A(n22596), .B(n22595), .Z(n22664) );
  AND U24221 ( .A(o[236]), .B(n22597), .Z(n22663) );
  XOR U24222 ( .A(n22664), .B(n22663), .Z(n22671) );
  AND U24223 ( .A(x[486]), .B(y[7911]), .Z(n23692) );
  AND U24224 ( .A(y[7915]), .B(x[482]), .Z(n22599) );
  NAND U24225 ( .A(y[7908]), .B(x[489]), .Z(n22598) );
  XOR U24226 ( .A(n22599), .B(n22598), .Z(n22687) );
  XOR U24227 ( .A(n22671), .B(n22670), .Z(n22672) );
  XOR U24228 ( .A(n22673), .B(n22672), .Z(n22708) );
  NAND U24229 ( .A(n22601), .B(n22600), .Z(n22605) );
  ANDN U24230 ( .B(n22603), .A(n22602), .Z(n22604) );
  ANDN U24231 ( .B(n22605), .A(n22604), .Z(n22707) );
  XOR U24232 ( .A(n22708), .B(n22707), .Z(n22710) );
  XOR U24233 ( .A(n22709), .B(n22710), .Z(n22701) );
  NAND U24234 ( .A(n22607), .B(n22606), .Z(n22611) );
  NAND U24235 ( .A(n22609), .B(n22608), .Z(n22610) );
  NAND U24236 ( .A(n22611), .B(n22610), .Z(n22648) );
  AND U24237 ( .A(x[486]), .B(y[7915]), .Z(n22985) );
  IV U24238 ( .A(n22985), .Z(n23060) );
  AND U24239 ( .A(x[481]), .B(y[7910]), .Z(n22662) );
  NANDN U24240 ( .A(n23060), .B(n22662), .Z(n22615) );
  NAND U24241 ( .A(n22613), .B(n22612), .Z(n22614) );
  NAND U24242 ( .A(n22615), .B(n22614), .Z(n22655) );
  AND U24243 ( .A(x[492]), .B(y[7916]), .Z(n23914) );
  NAND U24244 ( .A(n23914), .B(n22817), .Z(n22619) );
  NAND U24245 ( .A(n22617), .B(n22616), .Z(n22618) );
  NAND U24246 ( .A(n22619), .B(n22618), .Z(n22653) );
  AND U24247 ( .A(x[490]), .B(y[7907]), .Z(n23541) );
  AND U24248 ( .A(y[7906]), .B(x[491]), .Z(n23502) );
  NAND U24249 ( .A(y[7909]), .B(x[488]), .Z(n22620) );
  XNOR U24250 ( .A(n23502), .B(n22620), .Z(n22659) );
  XOR U24251 ( .A(n23541), .B(n22659), .Z(n22652) );
  XOR U24252 ( .A(n22653), .B(n22652), .Z(n22654) );
  XOR U24253 ( .A(n22655), .B(n22654), .Z(n22646) );
  AND U24254 ( .A(x[490]), .B(y[7912]), .Z(n22622) );
  AND U24255 ( .A(x[484]), .B(y[7906]), .Z(n22621) );
  NAND U24256 ( .A(n22622), .B(n22621), .Z(n22625) );
  NAND U24257 ( .A(n23249), .B(n22623), .Z(n22624) );
  NAND U24258 ( .A(n22625), .B(n22624), .Z(n22697) );
  AND U24259 ( .A(y[7904]), .B(x[493]), .Z(n22627) );
  NAND U24260 ( .A(y[7917]), .B(x[480]), .Z(n22626) );
  XNOR U24261 ( .A(n22627), .B(n22626), .Z(n22681) );
  NAND U24262 ( .A(x[492]), .B(y[7905]), .Z(n22692) );
  XOR U24263 ( .A(n22681), .B(n22680), .Z(n22696) );
  AND U24264 ( .A(y[7912]), .B(x[485]), .Z(n22629) );
  NAND U24265 ( .A(y[7914]), .B(x[483]), .Z(n22628) );
  XNOR U24266 ( .A(n22629), .B(n22628), .Z(n22676) );
  AND U24267 ( .A(x[484]), .B(y[7913]), .Z(n22677) );
  XOR U24268 ( .A(n22676), .B(n22677), .Z(n22695) );
  XOR U24269 ( .A(n22696), .B(n22695), .Z(n22698) );
  XOR U24270 ( .A(n22697), .B(n22698), .Z(n22647) );
  XOR U24271 ( .A(n22646), .B(n22647), .Z(n22649) );
  XOR U24272 ( .A(n22648), .B(n22649), .Z(n22703) );
  XNOR U24273 ( .A(n22704), .B(n22703), .Z(n22721) );
  NAND U24274 ( .A(n22631), .B(n22630), .Z(n22635) );
  NAND U24275 ( .A(n22633), .B(n22632), .Z(n22634) );
  AND U24276 ( .A(n22635), .B(n22634), .Z(n22720) );
  XOR U24277 ( .A(n22721), .B(n22720), .Z(n22722) );
  XOR U24278 ( .A(n22723), .B(n22722), .Z(n22716) );
  NAND U24279 ( .A(n22640), .B(n22639), .Z(n22644) );
  NAND U24280 ( .A(n22642), .B(n22641), .Z(n22643) );
  NAND U24281 ( .A(n22644), .B(n22643), .Z(n22715) );
  IV U24282 ( .A(n22715), .Z(n22713) );
  XOR U24283 ( .A(n22714), .B(n22713), .Z(n22645) );
  XNOR U24284 ( .A(n22716), .B(n22645), .Z(N494) );
  NAND U24285 ( .A(n22647), .B(n22646), .Z(n22651) );
  NAND U24286 ( .A(n22649), .B(n22648), .Z(n22650) );
  NAND U24287 ( .A(n22651), .B(n22650), .Z(n22729) );
  NAND U24288 ( .A(n22653), .B(n22652), .Z(n22657) );
  NAND U24289 ( .A(n22655), .B(n22654), .Z(n22656) );
  AND U24290 ( .A(n22657), .B(n22656), .Z(n22736) );
  AND U24291 ( .A(x[491]), .B(y[7909]), .Z(n22843) );
  NAND U24292 ( .A(n22843), .B(n22658), .Z(n22661) );
  NAND U24293 ( .A(n22659), .B(n23541), .Z(n22660) );
  AND U24294 ( .A(n22661), .B(n22660), .Z(n22791) );
  NAND U24295 ( .A(x[487]), .B(y[7916]), .Z(n23264) );
  NANDN U24296 ( .A(n23264), .B(n22662), .Z(n22666) );
  NAND U24297 ( .A(n22664), .B(n22663), .Z(n22665) );
  NAND U24298 ( .A(n22666), .B(n22665), .Z(n22790) );
  AND U24299 ( .A(x[484]), .B(y[7914]), .Z(n23165) );
  AND U24300 ( .A(y[7915]), .B(x[483]), .Z(n22668) );
  NAND U24301 ( .A(y[7910]), .B(x[488]), .Z(n22667) );
  XOR U24302 ( .A(n22668), .B(n22667), .Z(n22776) );
  XOR U24303 ( .A(n23165), .B(n22785), .Z(n22787) );
  AND U24304 ( .A(x[489]), .B(y[7909]), .Z(n23380) );
  AND U24305 ( .A(y[7916]), .B(x[482]), .Z(n22669) );
  AND U24306 ( .A(y[7908]), .B(x[490]), .Z(n23404) );
  XOR U24307 ( .A(n22669), .B(n23404), .Z(n22762) );
  XOR U24308 ( .A(n23380), .B(n22762), .Z(n22786) );
  XOR U24309 ( .A(n22787), .B(n22786), .Z(n22792) );
  XNOR U24310 ( .A(n22793), .B(n22792), .Z(n22734) );
  NAND U24311 ( .A(n22671), .B(n22670), .Z(n22675) );
  NAND U24312 ( .A(n22673), .B(n22672), .Z(n22674) );
  AND U24313 ( .A(n22675), .B(n22674), .Z(n22733) );
  XOR U24314 ( .A(n22734), .B(n22733), .Z(n22735) );
  XNOR U24315 ( .A(n22736), .B(n22735), .Z(n22728) );
  AND U24316 ( .A(x[485]), .B(y[7914]), .Z(n22830) );
  NAND U24317 ( .A(n23529), .B(n22830), .Z(n22679) );
  NAND U24318 ( .A(n22677), .B(n22676), .Z(n22678) );
  NAND U24319 ( .A(n22679), .B(n22678), .Z(n22742) );
  AND U24320 ( .A(x[493]), .B(y[7917]), .Z(n24216) );
  NAND U24321 ( .A(n24216), .B(n22817), .Z(n22683) );
  NAND U24322 ( .A(n22681), .B(n22680), .Z(n22682) );
  NAND U24323 ( .A(n22683), .B(n22682), .Z(n22740) );
  NAND U24324 ( .A(y[7907]), .B(x[491]), .Z(n22684) );
  XNOR U24325 ( .A(n22685), .B(n22684), .Z(n22766) );
  NAND U24326 ( .A(x[481]), .B(y[7917]), .Z(n22767) );
  XOR U24327 ( .A(n22740), .B(n22739), .Z(n22741) );
  XNOR U24328 ( .A(n22742), .B(n22741), .Z(n22797) );
  AND U24329 ( .A(x[489]), .B(y[7915]), .Z(n22686) );
  NAND U24330 ( .A(n22686), .B(n22761), .Z(n22689) );
  NANDN U24331 ( .A(n22687), .B(n23692), .Z(n22688) );
  AND U24332 ( .A(n22689), .B(n22688), .Z(n22748) );
  AND U24333 ( .A(y[7904]), .B(x[494]), .Z(n22691) );
  NAND U24334 ( .A(y[7918]), .B(x[480]), .Z(n22690) );
  XNOR U24335 ( .A(n22691), .B(n22690), .Z(n22771) );
  ANDN U24336 ( .B(o[237]), .A(n22692), .Z(n22770) );
  XOR U24337 ( .A(n22771), .B(n22770), .Z(n22746) );
  NAND U24338 ( .A(y[7906]), .B(x[492]), .Z(n22693) );
  XNOR U24339 ( .A(n22694), .B(n22693), .Z(n22753) );
  NAND U24340 ( .A(x[493]), .B(y[7905]), .Z(n22760) );
  XOR U24341 ( .A(n22753), .B(n22752), .Z(n22745) );
  XOR U24342 ( .A(n22746), .B(n22745), .Z(n22747) );
  XOR U24343 ( .A(n22748), .B(n22747), .Z(n22796) );
  XOR U24344 ( .A(n22797), .B(n22796), .Z(n22799) );
  NAND U24345 ( .A(n22696), .B(n22695), .Z(n22700) );
  NAND U24346 ( .A(n22698), .B(n22697), .Z(n22699) );
  AND U24347 ( .A(n22700), .B(n22699), .Z(n22798) );
  XNOR U24348 ( .A(n22799), .B(n22798), .Z(n22727) );
  XOR U24349 ( .A(n22728), .B(n22727), .Z(n22730) );
  XOR U24350 ( .A(n22729), .B(n22730), .Z(n22808) );
  NANDN U24351 ( .A(n22702), .B(n22701), .Z(n22706) );
  NAND U24352 ( .A(n22704), .B(n22703), .Z(n22705) );
  AND U24353 ( .A(n22706), .B(n22705), .Z(n22806) );
  NAND U24354 ( .A(n22708), .B(n22707), .Z(n22712) );
  NAND U24355 ( .A(n22710), .B(n22709), .Z(n22711) );
  NAND U24356 ( .A(n22712), .B(n22711), .Z(n22805) );
  XNOR U24357 ( .A(n22808), .B(n22807), .Z(n22804) );
  NANDN U24358 ( .A(n22713), .B(n22714), .Z(n22719) );
  NOR U24359 ( .A(n22715), .B(n22714), .Z(n22717) );
  OR U24360 ( .A(n22717), .B(n22716), .Z(n22718) );
  AND U24361 ( .A(n22719), .B(n22718), .Z(n22802) );
  NAND U24362 ( .A(n22721), .B(n22720), .Z(n22725) );
  NANDN U24363 ( .A(n22723), .B(n22722), .Z(n22724) );
  AND U24364 ( .A(n22725), .B(n22724), .Z(n22803) );
  XOR U24365 ( .A(n22802), .B(n22803), .Z(n22726) );
  XNOR U24366 ( .A(n22804), .B(n22726), .Z(N495) );
  NAND U24367 ( .A(n22728), .B(n22727), .Z(n22732) );
  NAND U24368 ( .A(n22730), .B(n22729), .Z(n22731) );
  NAND U24369 ( .A(n22732), .B(n22731), .Z(n22903) );
  NAND U24370 ( .A(n22734), .B(n22733), .Z(n22738) );
  NAND U24371 ( .A(n22736), .B(n22735), .Z(n22737) );
  AND U24372 ( .A(n22738), .B(n22737), .Z(n22873) );
  NAND U24373 ( .A(n22740), .B(n22739), .Z(n22744) );
  NAND U24374 ( .A(n22742), .B(n22741), .Z(n22743) );
  AND U24375 ( .A(n22744), .B(n22743), .Z(n22879) );
  NAND U24376 ( .A(n22746), .B(n22745), .Z(n22750) );
  NANDN U24377 ( .A(n22748), .B(n22747), .Z(n22749) );
  AND U24378 ( .A(n22750), .B(n22749), .Z(n22877) );
  NAND U24379 ( .A(x[492]), .B(y[7911]), .Z(n23256) );
  NANDN U24380 ( .A(n23256), .B(n22751), .Z(n22755) );
  NAND U24381 ( .A(n22753), .B(n22752), .Z(n22754) );
  AND U24382 ( .A(n22755), .B(n22754), .Z(n22853) );
  AND U24383 ( .A(y[7908]), .B(x[491]), .Z(n22757) );
  NAND U24384 ( .A(y[7906]), .B(x[493]), .Z(n22756) );
  XNOR U24385 ( .A(n22757), .B(n22756), .Z(n22857) );
  AND U24386 ( .A(x[492]), .B(y[7907]), .Z(n22856) );
  XOR U24387 ( .A(n22857), .B(n22856), .Z(n22851) );
  AND U24388 ( .A(y[7904]), .B(x[495]), .Z(n22759) );
  NAND U24389 ( .A(y[7919]), .B(x[480]), .Z(n22758) );
  XNOR U24390 ( .A(n22759), .B(n22758), .Z(n22819) );
  ANDN U24391 ( .B(o[238]), .A(n22760), .Z(n22818) );
  XNOR U24392 ( .A(n22819), .B(n22818), .Z(n22850) );
  XOR U24393 ( .A(n22853), .B(n22852), .Z(n22885) );
  NAND U24394 ( .A(x[490]), .B(y[7916]), .Z(n23694) );
  NANDN U24395 ( .A(n23694), .B(n22761), .Z(n22764) );
  NAND U24396 ( .A(n23380), .B(n22762), .Z(n22763) );
  AND U24397 ( .A(n22764), .B(n22763), .Z(n22883) );
  AND U24398 ( .A(x[491]), .B(y[7912]), .Z(n23164) );
  NAND U24399 ( .A(n23164), .B(n22765), .Z(n22769) );
  NANDN U24400 ( .A(n22767), .B(n22766), .Z(n22768) );
  NAND U24401 ( .A(n22769), .B(n22768), .Z(n22882) );
  AND U24402 ( .A(x[494]), .B(y[7918]), .Z(n24552) );
  NAND U24403 ( .A(n24552), .B(n22817), .Z(n22773) );
  NAND U24404 ( .A(n22771), .B(n22770), .Z(n22772) );
  AND U24405 ( .A(n22773), .B(n22772), .Z(n22845) );
  AND U24406 ( .A(x[488]), .B(y[7915]), .Z(n22774) );
  NAND U24407 ( .A(n22775), .B(n22774), .Z(n22778) );
  NANDN U24408 ( .A(n22776), .B(n23058), .Z(n22777) );
  NAND U24409 ( .A(n22778), .B(n22777), .Z(n22844) );
  AND U24410 ( .A(y[7909]), .B(x[490]), .Z(n22780) );
  NAND U24411 ( .A(y[7915]), .B(x[484]), .Z(n22779) );
  XNOR U24412 ( .A(n22780), .B(n22779), .Z(n22825) );
  AND U24413 ( .A(x[487]), .B(y[7912]), .Z(n22824) );
  XOR U24414 ( .A(n22825), .B(n22824), .Z(n22832) );
  NAND U24415 ( .A(x[486]), .B(y[7913]), .Z(n22935) );
  XNOR U24416 ( .A(n22935), .B(n22830), .Z(n22831) );
  AND U24417 ( .A(y[7917]), .B(x[482]), .Z(n22782) );
  NAND U24418 ( .A(y[7910]), .B(x[489]), .Z(n22781) );
  XNOR U24419 ( .A(n22782), .B(n22781), .Z(n22835) );
  NAND U24420 ( .A(x[483]), .B(y[7916]), .Z(n22836) );
  AND U24421 ( .A(y[7918]), .B(x[481]), .Z(n22784) );
  NAND U24422 ( .A(y[7911]), .B(x[488]), .Z(n22783) );
  XNOR U24423 ( .A(n22784), .B(n22783), .Z(n22814) );
  AND U24424 ( .A(x[494]), .B(y[7905]), .Z(n22841) );
  XOR U24425 ( .A(o[239]), .B(n22841), .Z(n22813) );
  XOR U24426 ( .A(n22814), .B(n22813), .Z(n22864) );
  XOR U24427 ( .A(n22865), .B(n22864), .Z(n22867) );
  XOR U24428 ( .A(n22866), .B(n22867), .Z(n22846) );
  XOR U24429 ( .A(n22847), .B(n22846), .Z(n22889) );
  NAND U24430 ( .A(n23165), .B(n22785), .Z(n22789) );
  NAND U24431 ( .A(n22787), .B(n22786), .Z(n22788) );
  AND U24432 ( .A(n22789), .B(n22788), .Z(n22888) );
  NANDN U24433 ( .A(n22791), .B(n22790), .Z(n22795) );
  NAND U24434 ( .A(n22793), .B(n22792), .Z(n22794) );
  NAND U24435 ( .A(n22795), .B(n22794), .Z(n22891) );
  XOR U24436 ( .A(n22870), .B(n22871), .Z(n22872) );
  NAND U24437 ( .A(n22797), .B(n22796), .Z(n22801) );
  NAND U24438 ( .A(n22799), .B(n22798), .Z(n22800) );
  AND U24439 ( .A(n22801), .B(n22800), .Z(n22901) );
  XNOR U24440 ( .A(n22902), .B(n22901), .Z(n22904) );
  XOR U24441 ( .A(n22903), .B(n22904), .Z(n22897) );
  NANDN U24442 ( .A(n22806), .B(n22805), .Z(n22810) );
  NAND U24443 ( .A(n22808), .B(n22807), .Z(n22809) );
  NAND U24444 ( .A(n22810), .B(n22809), .Z(n22895) );
  IV U24445 ( .A(n22895), .Z(n22894) );
  XOR U24446 ( .A(n22896), .B(n22894), .Z(n22811) );
  XNOR U24447 ( .A(n22897), .B(n22811), .Z(N496) );
  AND U24448 ( .A(x[488]), .B(y[7918]), .Z(n23166) );
  NAND U24449 ( .A(n23166), .B(n22812), .Z(n22816) );
  NAND U24450 ( .A(n22814), .B(n22813), .Z(n22815) );
  AND U24451 ( .A(n22816), .B(n22815), .Z(n22965) );
  AND U24452 ( .A(x[495]), .B(y[7919]), .Z(n24984) );
  NAND U24453 ( .A(n24984), .B(n22817), .Z(n22821) );
  NAND U24454 ( .A(n22819), .B(n22818), .Z(n22820) );
  NAND U24455 ( .A(n22821), .B(n22820), .Z(n22964) );
  AND U24456 ( .A(x[490]), .B(y[7915]), .Z(n22823) );
  NAND U24457 ( .A(n22823), .B(n22822), .Z(n22827) );
  NAND U24458 ( .A(n22825), .B(n22824), .Z(n22826) );
  NAND U24459 ( .A(n22827), .B(n22826), .Z(n22922) );
  AND U24460 ( .A(x[480]), .B(y[7920]), .Z(n22944) );
  AND U24461 ( .A(x[496]), .B(y[7904]), .Z(n22945) );
  XOR U24462 ( .A(n22944), .B(n22945), .Z(n22947) );
  AND U24463 ( .A(x[495]), .B(y[7905]), .Z(n22932) );
  XOR U24464 ( .A(o[240]), .B(n22932), .Z(n22946) );
  XOR U24465 ( .A(n22947), .B(n22946), .Z(n22921) );
  NAND U24466 ( .A(y[7913]), .B(x[487]), .Z(n22828) );
  XNOR U24467 ( .A(n22829), .B(n22828), .Z(n22937) );
  AND U24468 ( .A(x[490]), .B(y[7910]), .Z(n22936) );
  XOR U24469 ( .A(n22937), .B(n22936), .Z(n22920) );
  XOR U24470 ( .A(n22921), .B(n22920), .Z(n22923) );
  XOR U24471 ( .A(n22922), .B(n22923), .Z(n22966) );
  XOR U24472 ( .A(n22967), .B(n22966), .Z(n22917) );
  NANDN U24473 ( .A(n22830), .B(n22935), .Z(n22834) );
  NANDN U24474 ( .A(n22832), .B(n22831), .Z(n22833) );
  AND U24475 ( .A(n22834), .B(n22833), .Z(n22915) );
  NAND U24476 ( .A(x[489]), .B(y[7917]), .Z(n23675) );
  NANDN U24477 ( .A(n23675), .B(n23254), .Z(n22838) );
  NANDN U24478 ( .A(n22836), .B(n22835), .Z(n22837) );
  AND U24479 ( .A(n22838), .B(n22837), .Z(n22955) );
  AND U24480 ( .A(y[7919]), .B(x[481]), .Z(n22840) );
  NAND U24481 ( .A(y[7912]), .B(x[488]), .Z(n22839) );
  XNOR U24482 ( .A(n22840), .B(n22839), .Z(n22941) );
  AND U24483 ( .A(o[239]), .B(n22841), .Z(n22940) );
  XOR U24484 ( .A(n22941), .B(n22940), .Z(n22953) );
  NAND U24485 ( .A(y[7906]), .B(x[494]), .Z(n22842) );
  XNOR U24486 ( .A(n22843), .B(n22842), .Z(n22976) );
  AND U24487 ( .A(x[484]), .B(y[7916]), .Z(n22977) );
  XOR U24488 ( .A(n22976), .B(n22977), .Z(n22952) );
  XOR U24489 ( .A(n22953), .B(n22952), .Z(n22954) );
  XOR U24490 ( .A(n22955), .B(n22954), .Z(n22914) );
  NANDN U24491 ( .A(n22845), .B(n22844), .Z(n22849) );
  NAND U24492 ( .A(n22847), .B(n22846), .Z(n22848) );
  NAND U24493 ( .A(n22849), .B(n22848), .Z(n22959) );
  NANDN U24494 ( .A(n22851), .B(n22850), .Z(n22855) );
  NAND U24495 ( .A(n22853), .B(n22852), .Z(n22854) );
  AND U24496 ( .A(n22855), .B(n22854), .Z(n22991) );
  AND U24497 ( .A(x[493]), .B(y[7908]), .Z(n22987) );
  NAND U24498 ( .A(n23502), .B(n22987), .Z(n22859) );
  NAND U24499 ( .A(n22857), .B(n22856), .Z(n22858) );
  AND U24500 ( .A(n22859), .B(n22858), .Z(n22973) );
  AND U24501 ( .A(y[7918]), .B(x[482]), .Z(n22861) );
  NAND U24502 ( .A(y[7911]), .B(x[489]), .Z(n22860) );
  XNOR U24503 ( .A(n22861), .B(n22860), .Z(n22980) );
  AND U24504 ( .A(x[483]), .B(y[7917]), .Z(n22981) );
  XOR U24505 ( .A(n22980), .B(n22981), .Z(n22971) );
  AND U24506 ( .A(x[492]), .B(y[7908]), .Z(n23663) );
  AND U24507 ( .A(y[7915]), .B(x[485]), .Z(n22863) );
  NAND U24508 ( .A(y[7907]), .B(x[493]), .Z(n22862) );
  XNOR U24509 ( .A(n22863), .B(n22862), .Z(n22927) );
  XOR U24510 ( .A(n23663), .B(n22927), .Z(n22970) );
  XOR U24511 ( .A(n22971), .B(n22970), .Z(n22972) );
  NAND U24512 ( .A(n22865), .B(n22864), .Z(n22869) );
  NAND U24513 ( .A(n22867), .B(n22866), .Z(n22868) );
  AND U24514 ( .A(n22869), .B(n22868), .Z(n22989) );
  XOR U24515 ( .A(n22988), .B(n22989), .Z(n22990) );
  XOR U24516 ( .A(n22961), .B(n22960), .Z(n22995) );
  NAND U24517 ( .A(n22871), .B(n22870), .Z(n22875) );
  NANDN U24518 ( .A(n22873), .B(n22872), .Z(n22874) );
  AND U24519 ( .A(n22875), .B(n22874), .Z(n22994) );
  NANDN U24520 ( .A(n22877), .B(n22876), .Z(n22881) );
  NANDN U24521 ( .A(n22879), .B(n22878), .Z(n22880) );
  AND U24522 ( .A(n22881), .B(n22880), .Z(n22911) );
  NANDN U24523 ( .A(n22883), .B(n22882), .Z(n22887) );
  NANDN U24524 ( .A(n22885), .B(n22884), .Z(n22886) );
  AND U24525 ( .A(n22887), .B(n22886), .Z(n22909) );
  NANDN U24526 ( .A(n22889), .B(n22888), .Z(n22893) );
  NANDN U24527 ( .A(n22891), .B(n22890), .Z(n22892) );
  AND U24528 ( .A(n22893), .B(n22892), .Z(n22908) );
  XNOR U24529 ( .A(n22997), .B(n22996), .Z(n23002) );
  OR U24530 ( .A(n22896), .B(n22894), .Z(n22900) );
  ANDN U24531 ( .B(n22896), .A(n22895), .Z(n22898) );
  OR U24532 ( .A(n22898), .B(n22897), .Z(n22899) );
  AND U24533 ( .A(n22900), .B(n22899), .Z(n23001) );
  NAND U24534 ( .A(n22902), .B(n22901), .Z(n22906) );
  NANDN U24535 ( .A(n22904), .B(n22903), .Z(n22905) );
  NAND U24536 ( .A(n22906), .B(n22905), .Z(n23000) );
  XNOR U24537 ( .A(n23001), .B(n23000), .Z(n22907) );
  XNOR U24538 ( .A(n23002), .B(n22907), .Z(N497) );
  NANDN U24539 ( .A(n22909), .B(n22908), .Z(n22913) );
  NANDN U24540 ( .A(n22911), .B(n22910), .Z(n22912) );
  AND U24541 ( .A(n22913), .B(n22912), .Z(n23104) );
  NANDN U24542 ( .A(n22915), .B(n22914), .Z(n22919) );
  NANDN U24543 ( .A(n22917), .B(n22916), .Z(n22918) );
  AND U24544 ( .A(n22919), .B(n22918), .Z(n23013) );
  NAND U24545 ( .A(n22921), .B(n22920), .Z(n22925) );
  NAND U24546 ( .A(n22923), .B(n22922), .Z(n22924) );
  AND U24547 ( .A(n22925), .B(n22924), .Z(n23095) );
  AND U24548 ( .A(x[493]), .B(y[7915]), .Z(n23922) );
  NAND U24549 ( .A(n23922), .B(n22926), .Z(n22929) );
  NAND U24550 ( .A(n22927), .B(n23663), .Z(n22928) );
  NAND U24551 ( .A(n22929), .B(n22928), .Z(n23043) );
  AND U24552 ( .A(y[7920]), .B(x[481]), .Z(n22931) );
  NAND U24553 ( .A(y[7912]), .B(x[489]), .Z(n22930) );
  XNOR U24554 ( .A(n22931), .B(n22930), .Z(n23064) );
  AND U24555 ( .A(o[240]), .B(n22932), .Z(n23063) );
  XOR U24556 ( .A(n23064), .B(n23063), .Z(n23041) );
  AND U24557 ( .A(y[7906]), .B(x[495]), .Z(n22934) );
  NAND U24558 ( .A(y[7909]), .B(x[492]), .Z(n22933) );
  XNOR U24559 ( .A(n22934), .B(n22933), .Z(n23016) );
  NAND U24560 ( .A(x[494]), .B(y[7907]), .Z(n23017) );
  XOR U24561 ( .A(n23041), .B(n23040), .Z(n23042) );
  XOR U24562 ( .A(n23043), .B(n23042), .Z(n23093) );
  AND U24563 ( .A(x[487]), .B(y[7914]), .Z(n23075) );
  NANDN U24564 ( .A(n22935), .B(n23075), .Z(n22939) );
  NAND U24565 ( .A(n22937), .B(n22936), .Z(n22938) );
  NAND U24566 ( .A(n22939), .B(n22938), .Z(n23053) );
  NAND U24567 ( .A(x[488]), .B(y[7919]), .Z(n23753) );
  AND U24568 ( .A(x[481]), .B(y[7912]), .Z(n23144) );
  NANDN U24569 ( .A(n23753), .B(n23144), .Z(n22943) );
  NAND U24570 ( .A(n22941), .B(n22940), .Z(n22942) );
  NAND U24571 ( .A(n22943), .B(n22942), .Z(n23052) );
  XOR U24572 ( .A(n23053), .B(n23052), .Z(n23055) );
  NAND U24573 ( .A(n22945), .B(n22944), .Z(n22949) );
  NAND U24574 ( .A(n22947), .B(n22946), .Z(n22948) );
  NAND U24575 ( .A(n22949), .B(n22948), .Z(n23049) );
  AND U24576 ( .A(x[480]), .B(y[7921]), .Z(n23030) );
  NAND U24577 ( .A(x[497]), .B(y[7904]), .Z(n23031) );
  AND U24578 ( .A(x[496]), .B(y[7905]), .Z(n23027) );
  XOR U24579 ( .A(o[241]), .B(n23027), .Z(n23032) );
  XOR U24580 ( .A(n23033), .B(n23032), .Z(n23047) );
  AND U24581 ( .A(y[7919]), .B(x[482]), .Z(n22951) );
  NAND U24582 ( .A(y[7911]), .B(x[490]), .Z(n22950) );
  XNOR U24583 ( .A(n22951), .B(n22950), .Z(n23068) );
  AND U24584 ( .A(x[483]), .B(y[7918]), .Z(n23069) );
  XOR U24585 ( .A(n23068), .B(n23069), .Z(n23046) );
  XOR U24586 ( .A(n23047), .B(n23046), .Z(n23048) );
  XOR U24587 ( .A(n23049), .B(n23048), .Z(n23054) );
  XOR U24588 ( .A(n23055), .B(n23054), .Z(n23092) );
  XOR U24589 ( .A(n23093), .B(n23092), .Z(n23094) );
  NAND U24590 ( .A(n22953), .B(n22952), .Z(n22957) );
  NANDN U24591 ( .A(n22955), .B(n22954), .Z(n22956) );
  AND U24592 ( .A(n22957), .B(n22956), .Z(n23011) );
  XOR U24593 ( .A(n23010), .B(n23011), .Z(n23012) );
  NANDN U24594 ( .A(n22959), .B(n22958), .Z(n22963) );
  NAND U24595 ( .A(n22961), .B(n22960), .Z(n22962) );
  AND U24596 ( .A(n22963), .B(n22962), .Z(n23007) );
  NANDN U24597 ( .A(n22965), .B(n22964), .Z(n22969) );
  NAND U24598 ( .A(n22967), .B(n22966), .Z(n22968) );
  AND U24599 ( .A(n22969), .B(n22968), .Z(n23089) );
  NAND U24600 ( .A(n22971), .B(n22970), .Z(n22975) );
  NANDN U24601 ( .A(n22973), .B(n22972), .Z(n22974) );
  AND U24602 ( .A(n22975), .B(n22974), .Z(n23087) );
  NAND U24603 ( .A(x[494]), .B(y[7909]), .Z(n23288) );
  NANDN U24604 ( .A(n23288), .B(n23502), .Z(n22979) );
  NAND U24605 ( .A(n22977), .B(n22976), .Z(n22978) );
  NAND U24606 ( .A(n22979), .B(n22978), .Z(n23081) );
  AND U24607 ( .A(x[489]), .B(y[7918]), .Z(n23903) );
  NANDN U24608 ( .A(n23067), .B(n23903), .Z(n22983) );
  NAND U24609 ( .A(n22981), .B(n22980), .Z(n22982) );
  NAND U24610 ( .A(n22983), .B(n22982), .Z(n23080) );
  XOR U24611 ( .A(n23081), .B(n23080), .Z(n23083) );
  AND U24612 ( .A(y[7916]), .B(x[485]), .Z(n23126) );
  NAND U24613 ( .A(y[7913]), .B(x[488]), .Z(n22984) );
  XNOR U24614 ( .A(n23126), .B(n22984), .Z(n23059) );
  XOR U24615 ( .A(n23059), .B(n22985), .Z(n23074) );
  XOR U24616 ( .A(n23075), .B(n23074), .Z(n23077) );
  NAND U24617 ( .A(y[7917]), .B(x[484]), .Z(n22986) );
  XNOR U24618 ( .A(n22987), .B(n22986), .Z(n23021) );
  AND U24619 ( .A(x[491]), .B(y[7910]), .Z(n23022) );
  XOR U24620 ( .A(n23021), .B(n23022), .Z(n23076) );
  XOR U24621 ( .A(n23077), .B(n23076), .Z(n23082) );
  XOR U24622 ( .A(n23083), .B(n23082), .Z(n23086) );
  NAND U24623 ( .A(n22989), .B(n22988), .Z(n22993) );
  NANDN U24624 ( .A(n22991), .B(n22990), .Z(n22992) );
  NAND U24625 ( .A(n22993), .B(n22992), .Z(n23004) );
  XOR U24626 ( .A(n23005), .B(n23004), .Z(n23006) );
  XOR U24627 ( .A(n23007), .B(n23006), .Z(n23101) );
  XOR U24628 ( .A(n23102), .B(n23101), .Z(n23103) );
  XOR U24629 ( .A(n23104), .B(n23103), .Z(n23100) );
  NANDN U24630 ( .A(n22995), .B(n22994), .Z(n22999) );
  NAND U24631 ( .A(n22997), .B(n22996), .Z(n22998) );
  NAND U24632 ( .A(n22999), .B(n22998), .Z(n23098) );
  XOR U24633 ( .A(n23098), .B(n23099), .Z(n23003) );
  XNOR U24634 ( .A(n23100), .B(n23003), .Z(N498) );
  NAND U24635 ( .A(n23005), .B(n23004), .Z(n23009) );
  NANDN U24636 ( .A(n23007), .B(n23006), .Z(n23008) );
  AND U24637 ( .A(n23009), .B(n23008), .Z(n23220) );
  NAND U24638 ( .A(n23011), .B(n23010), .Z(n23015) );
  NANDN U24639 ( .A(n23013), .B(n23012), .Z(n23014) );
  AND U24640 ( .A(n23015), .B(n23014), .Z(n23218) );
  AND U24641 ( .A(x[495]), .B(y[7909]), .Z(n23262) );
  AND U24642 ( .A(x[492]), .B(y[7906]), .Z(n23370) );
  NAND U24643 ( .A(n23262), .B(n23370), .Z(n23019) );
  NANDN U24644 ( .A(n23017), .B(n23016), .Z(n23018) );
  NAND U24645 ( .A(n23019), .B(n23018), .Z(n23193) );
  NAND U24646 ( .A(n24216), .B(n23020), .Z(n23024) );
  NAND U24647 ( .A(n23022), .B(n23021), .Z(n23023) );
  NAND U24648 ( .A(n23024), .B(n23023), .Z(n23183) );
  AND U24649 ( .A(y[7921]), .B(x[481]), .Z(n23026) );
  NAND U24650 ( .A(y[7912]), .B(x[490]), .Z(n23025) );
  XNOR U24651 ( .A(n23026), .B(n23025), .Z(n23146) );
  AND U24652 ( .A(o[241]), .B(n23027), .Z(n23145) );
  XOR U24653 ( .A(n23146), .B(n23145), .Z(n23181) );
  AND U24654 ( .A(y[7907]), .B(x[495]), .Z(n23029) );
  NAND U24655 ( .A(y[7913]), .B(x[489]), .Z(n23028) );
  XNOR U24656 ( .A(n23029), .B(n23028), .Z(n23136) );
  AND U24657 ( .A(x[494]), .B(y[7908]), .Z(n23137) );
  XOR U24658 ( .A(n23136), .B(n23137), .Z(n23180) );
  XOR U24659 ( .A(n23181), .B(n23180), .Z(n23182) );
  XOR U24660 ( .A(n23183), .B(n23182), .Z(n23192) );
  XOR U24661 ( .A(n23193), .B(n23192), .Z(n23195) );
  NANDN U24662 ( .A(n23031), .B(n23030), .Z(n23035) );
  NAND U24663 ( .A(n23033), .B(n23032), .Z(n23034) );
  AND U24664 ( .A(n23035), .B(n23034), .Z(n23205) );
  AND U24665 ( .A(y[7906]), .B(x[496]), .Z(n23037) );
  NAND U24666 ( .A(y[7911]), .B(x[491]), .Z(n23036) );
  XNOR U24667 ( .A(n23037), .B(n23036), .Z(n23132) );
  AND U24668 ( .A(x[482]), .B(y[7920]), .Z(n23133) );
  XOR U24669 ( .A(n23132), .B(n23133), .Z(n23204) );
  AND U24670 ( .A(y[7917]), .B(x[485]), .Z(n23270) );
  NAND U24671 ( .A(y[7916]), .B(x[486]), .Z(n23038) );
  XNOR U24672 ( .A(n23270), .B(n23038), .Z(n23129) );
  NAND U24673 ( .A(y[7918]), .B(x[484]), .Z(n23039) );
  XNOR U24674 ( .A(n23908), .B(n23039), .Z(n23167) );
  AND U24675 ( .A(x[487]), .B(y[7915]), .Z(n23168) );
  XOR U24676 ( .A(n23167), .B(n23168), .Z(n23128) );
  XOR U24677 ( .A(n23129), .B(n23128), .Z(n23206) );
  XOR U24678 ( .A(n23207), .B(n23206), .Z(n23194) );
  XOR U24679 ( .A(n23195), .B(n23194), .Z(n23115) );
  NAND U24680 ( .A(n23041), .B(n23040), .Z(n23045) );
  NAND U24681 ( .A(n23043), .B(n23042), .Z(n23044) );
  AND U24682 ( .A(n23045), .B(n23044), .Z(n23186) );
  NAND U24683 ( .A(n23047), .B(n23046), .Z(n23051) );
  NAND U24684 ( .A(n23049), .B(n23048), .Z(n23050) );
  AND U24685 ( .A(n23051), .B(n23050), .Z(n23187) );
  XOR U24686 ( .A(n23186), .B(n23187), .Z(n23188) );
  NAND U24687 ( .A(n23053), .B(n23052), .Z(n23057) );
  NAND U24688 ( .A(n23055), .B(n23054), .Z(n23056) );
  AND U24689 ( .A(n23057), .B(n23056), .Z(n23189) );
  XOR U24690 ( .A(n23188), .B(n23189), .Z(n23114) );
  AND U24691 ( .A(x[488]), .B(y[7916]), .Z(n23410) );
  NAND U24692 ( .A(n23410), .B(n23058), .Z(n23062) );
  NANDN U24693 ( .A(n23060), .B(n23059), .Z(n23061) );
  NAND U24694 ( .A(n23062), .B(n23061), .Z(n23199) );
  AND U24695 ( .A(x[489]), .B(y[7920]), .Z(n24056) );
  IV U24696 ( .A(n24056), .Z(n23932) );
  NANDN U24697 ( .A(n23932), .B(n23144), .Z(n23066) );
  NAND U24698 ( .A(n23064), .B(n23063), .Z(n23065) );
  NAND U24699 ( .A(n23066), .B(n23065), .Z(n23198) );
  XOR U24700 ( .A(n23199), .B(n23198), .Z(n23201) );
  AND U24701 ( .A(x[490]), .B(y[7919]), .Z(n23931) );
  NANDN U24702 ( .A(n23067), .B(n23931), .Z(n23071) );
  NAND U24703 ( .A(n23069), .B(n23068), .Z(n23070) );
  NAND U24704 ( .A(n23071), .B(n23070), .Z(n23177) );
  AND U24705 ( .A(x[480]), .B(y[7922]), .Z(n23149) );
  AND U24706 ( .A(x[498]), .B(y[7904]), .Z(n23150) );
  XOR U24707 ( .A(n23149), .B(n23150), .Z(n23152) );
  AND U24708 ( .A(x[497]), .B(y[7905]), .Z(n23171) );
  XOR U24709 ( .A(o[242]), .B(n23171), .Z(n23151) );
  XOR U24710 ( .A(n23152), .B(n23151), .Z(n23175) );
  AND U24711 ( .A(y[7909]), .B(x[493]), .Z(n23073) );
  NAND U24712 ( .A(y[7919]), .B(x[483]), .Z(n23072) );
  XNOR U24713 ( .A(n23073), .B(n23072), .Z(n23157) );
  AND U24714 ( .A(x[492]), .B(y[7910]), .Z(n23158) );
  XOR U24715 ( .A(n23157), .B(n23158), .Z(n23174) );
  XOR U24716 ( .A(n23175), .B(n23174), .Z(n23176) );
  XOR U24717 ( .A(n23177), .B(n23176), .Z(n23200) );
  XNOR U24718 ( .A(n23201), .B(n23200), .Z(n23121) );
  NAND U24719 ( .A(n23075), .B(n23074), .Z(n23079) );
  NAND U24720 ( .A(n23077), .B(n23076), .Z(n23078) );
  AND U24721 ( .A(n23079), .B(n23078), .Z(n23120) );
  XOR U24722 ( .A(n23121), .B(n23120), .Z(n23122) );
  NAND U24723 ( .A(n23081), .B(n23080), .Z(n23085) );
  NAND U24724 ( .A(n23083), .B(n23082), .Z(n23084) );
  AND U24725 ( .A(n23085), .B(n23084), .Z(n23123) );
  XOR U24726 ( .A(n23122), .B(n23123), .Z(n23116) );
  XOR U24727 ( .A(n23117), .B(n23116), .Z(n23111) );
  NANDN U24728 ( .A(n23087), .B(n23086), .Z(n23091) );
  NANDN U24729 ( .A(n23089), .B(n23088), .Z(n23090) );
  AND U24730 ( .A(n23091), .B(n23090), .Z(n23109) );
  NAND U24731 ( .A(n23093), .B(n23092), .Z(n23097) );
  NANDN U24732 ( .A(n23095), .B(n23094), .Z(n23096) );
  NAND U24733 ( .A(n23097), .B(n23096), .Z(n23108) );
  XOR U24734 ( .A(n23218), .B(n23217), .Z(n23219) );
  XNOR U24735 ( .A(n23220), .B(n23219), .Z(n23213) );
  NAND U24736 ( .A(n23102), .B(n23101), .Z(n23106) );
  NANDN U24737 ( .A(n23104), .B(n23103), .Z(n23105) );
  NAND U24738 ( .A(n23106), .B(n23105), .Z(n23211) );
  IV U24739 ( .A(n23211), .Z(n23210) );
  XOR U24740 ( .A(n23212), .B(n23210), .Z(n23107) );
  XNOR U24741 ( .A(n23213), .B(n23107), .Z(N499) );
  NANDN U24742 ( .A(n23109), .B(n23108), .Z(n23113) );
  NANDN U24743 ( .A(n23111), .B(n23110), .Z(n23112) );
  AND U24744 ( .A(n23113), .B(n23112), .Z(n23227) );
  NANDN U24745 ( .A(n23115), .B(n23114), .Z(n23119) );
  NAND U24746 ( .A(n23117), .B(n23116), .Z(n23118) );
  AND U24747 ( .A(n23119), .B(n23118), .Z(n23225) );
  NAND U24748 ( .A(n23121), .B(n23120), .Z(n23125) );
  NAND U24749 ( .A(n23123), .B(n23122), .Z(n23124) );
  NAND U24750 ( .A(n23125), .B(n23124), .Z(n23329) );
  AND U24751 ( .A(x[486]), .B(y[7917]), .Z(n23127) );
  NAND U24752 ( .A(n23127), .B(n23126), .Z(n23131) );
  NAND U24753 ( .A(n23129), .B(n23128), .Z(n23130) );
  NAND U24754 ( .A(n23131), .B(n23130), .Z(n23323) );
  AND U24755 ( .A(x[496]), .B(y[7911]), .Z(n23679) );
  NAND U24756 ( .A(n23679), .B(n23502), .Z(n23135) );
  NAND U24757 ( .A(n23133), .B(n23132), .Z(n23134) );
  NAND U24758 ( .A(n23135), .B(n23134), .Z(n23321) );
  AND U24759 ( .A(x[495]), .B(y[7913]), .Z(n23941) );
  NAND U24760 ( .A(n23941), .B(n23249), .Z(n23139) );
  NAND U24761 ( .A(n23137), .B(n23136), .Z(n23138) );
  NAND U24762 ( .A(n23139), .B(n23138), .Z(n23240) );
  AND U24763 ( .A(y[7922]), .B(x[481]), .Z(n23141) );
  NAND U24764 ( .A(y[7915]), .B(x[488]), .Z(n23140) );
  XNOR U24765 ( .A(n23141), .B(n23140), .Z(n23287) );
  AND U24766 ( .A(y[7910]), .B(x[493]), .Z(n23143) );
  NAND U24767 ( .A(y[7921]), .B(x[482]), .Z(n23142) );
  XNOR U24768 ( .A(n23143), .B(n23142), .Z(n23255) );
  XOR U24769 ( .A(n23238), .B(n23237), .Z(n23239) );
  XOR U24770 ( .A(n23240), .B(n23239), .Z(n23320) );
  XOR U24771 ( .A(n23321), .B(n23320), .Z(n23322) );
  XNOR U24772 ( .A(n23323), .B(n23322), .Z(n23327) );
  AND U24773 ( .A(x[490]), .B(y[7921]), .Z(n24307) );
  IV U24774 ( .A(n24307), .Z(n24416) );
  NANDN U24775 ( .A(n24416), .B(n23144), .Z(n23148) );
  NAND U24776 ( .A(n23146), .B(n23145), .Z(n23147) );
  NAND U24777 ( .A(n23148), .B(n23147), .Z(n23299) );
  NAND U24778 ( .A(n23150), .B(n23149), .Z(n23154) );
  NAND U24779 ( .A(n23152), .B(n23151), .Z(n23153) );
  NAND U24780 ( .A(n23154), .B(n23153), .Z(n23297) );
  AND U24781 ( .A(y[7907]), .B(x[496]), .Z(n23982) );
  NAND U24782 ( .A(y[7914]), .B(x[489]), .Z(n23155) );
  XNOR U24783 ( .A(n23982), .B(n23155), .Z(n23250) );
  AND U24784 ( .A(x[495]), .B(y[7908]), .Z(n23251) );
  XOR U24785 ( .A(n23250), .B(n23251), .Z(n23296) );
  XOR U24786 ( .A(n23297), .B(n23296), .Z(n23298) );
  XNOR U24787 ( .A(n23299), .B(n23298), .Z(n23316) );
  AND U24788 ( .A(x[493]), .B(y[7919]), .Z(n24579) );
  NANDN U24789 ( .A(n23156), .B(n24579), .Z(n23160) );
  NAND U24790 ( .A(n23158), .B(n23157), .Z(n23159) );
  NAND U24791 ( .A(n23160), .B(n23159), .Z(n23305) );
  AND U24792 ( .A(y[7913]), .B(x[490]), .Z(n23162) );
  NAND U24793 ( .A(y[7906]), .B(x[497]), .Z(n23161) );
  XNOR U24794 ( .A(n23162), .B(n23161), .Z(n23293) );
  AND U24795 ( .A(x[498]), .B(y[7905]), .Z(n23269) );
  XOR U24796 ( .A(o[243]), .B(n23269), .Z(n23292) );
  XOR U24797 ( .A(n23293), .B(n23292), .Z(n23303) );
  NAND U24798 ( .A(y[7920]), .B(x[483]), .Z(n23163) );
  XNOR U24799 ( .A(n23164), .B(n23163), .Z(n23263) );
  XOR U24800 ( .A(n23303), .B(n23302), .Z(n23304) );
  XNOR U24801 ( .A(n23305), .B(n23304), .Z(n23315) );
  NAND U24802 ( .A(n23166), .B(n23165), .Z(n23170) );
  NAND U24803 ( .A(n23168), .B(n23167), .Z(n23169) );
  AND U24804 ( .A(n23170), .B(n23169), .Z(n23246) );
  AND U24805 ( .A(x[480]), .B(y[7923]), .Z(n23274) );
  AND U24806 ( .A(x[499]), .B(y[7904]), .Z(n23275) );
  XOR U24807 ( .A(n23274), .B(n23275), .Z(n23277) );
  AND U24808 ( .A(o[242]), .B(n23171), .Z(n23276) );
  XOR U24809 ( .A(n23277), .B(n23276), .Z(n23244) );
  AND U24810 ( .A(x[484]), .B(y[7919]), .Z(n23424) );
  AND U24811 ( .A(y[7918]), .B(x[485]), .Z(n23173) );
  NAND U24812 ( .A(y[7917]), .B(x[486]), .Z(n23172) );
  XNOR U24813 ( .A(n23173), .B(n23172), .Z(n23271) );
  XOR U24814 ( .A(n23424), .B(n23271), .Z(n23243) );
  XOR U24815 ( .A(n23244), .B(n23243), .Z(n23245) );
  XOR U24816 ( .A(n23246), .B(n23245), .Z(n23314) );
  XOR U24817 ( .A(n23315), .B(n23314), .Z(n23317) );
  XNOR U24818 ( .A(n23316), .B(n23317), .Z(n23310) );
  NAND U24819 ( .A(n23175), .B(n23174), .Z(n23179) );
  NAND U24820 ( .A(n23177), .B(n23176), .Z(n23178) );
  NAND U24821 ( .A(n23179), .B(n23178), .Z(n23309) );
  NAND U24822 ( .A(n23181), .B(n23180), .Z(n23185) );
  NAND U24823 ( .A(n23183), .B(n23182), .Z(n23184) );
  NAND U24824 ( .A(n23185), .B(n23184), .Z(n23308) );
  XOR U24825 ( .A(n23309), .B(n23308), .Z(n23311) );
  XNOR U24826 ( .A(n23310), .B(n23311), .Z(n23326) );
  XOR U24827 ( .A(n23327), .B(n23326), .Z(n23328) );
  XNOR U24828 ( .A(n23329), .B(n23328), .Z(n23340) );
  NAND U24829 ( .A(n23187), .B(n23186), .Z(n23191) );
  NAND U24830 ( .A(n23189), .B(n23188), .Z(n23190) );
  AND U24831 ( .A(n23191), .B(n23190), .Z(n23339) );
  NAND U24832 ( .A(n23193), .B(n23192), .Z(n23197) );
  NAND U24833 ( .A(n23195), .B(n23194), .Z(n23196) );
  AND U24834 ( .A(n23197), .B(n23196), .Z(n23335) );
  NAND U24835 ( .A(n23199), .B(n23198), .Z(n23203) );
  NAND U24836 ( .A(n23201), .B(n23200), .Z(n23202) );
  AND U24837 ( .A(n23203), .B(n23202), .Z(n23333) );
  NANDN U24838 ( .A(n23205), .B(n23204), .Z(n23209) );
  NAND U24839 ( .A(n23207), .B(n23206), .Z(n23208) );
  NAND U24840 ( .A(n23209), .B(n23208), .Z(n23332) );
  XOR U24841 ( .A(n23339), .B(n23338), .Z(n23341) );
  XOR U24842 ( .A(n23340), .B(n23341), .Z(n23224) );
  XOR U24843 ( .A(n23225), .B(n23224), .Z(n23226) );
  XOR U24844 ( .A(n23227), .B(n23226), .Z(n23233) );
  OR U24845 ( .A(n23212), .B(n23210), .Z(n23216) );
  ANDN U24846 ( .B(n23212), .A(n23211), .Z(n23214) );
  OR U24847 ( .A(n23214), .B(n23213), .Z(n23215) );
  AND U24848 ( .A(n23216), .B(n23215), .Z(n23232) );
  NAND U24849 ( .A(n23218), .B(n23217), .Z(n23222) );
  NAND U24850 ( .A(n23220), .B(n23219), .Z(n23221) );
  NAND U24851 ( .A(n23222), .B(n23221), .Z(n23231) );
  IV U24852 ( .A(n23231), .Z(n23230) );
  XOR U24853 ( .A(n23232), .B(n23230), .Z(n23223) );
  XNOR U24854 ( .A(n23233), .B(n23223), .Z(N500) );
  NAND U24855 ( .A(n23225), .B(n23224), .Z(n23229) );
  NANDN U24856 ( .A(n23227), .B(n23226), .Z(n23228) );
  NAND U24857 ( .A(n23229), .B(n23228), .Z(n23352) );
  IV U24858 ( .A(n23352), .Z(n23351) );
  OR U24859 ( .A(n23232), .B(n23230), .Z(n23236) );
  ANDN U24860 ( .B(n23232), .A(n23231), .Z(n23234) );
  OR U24861 ( .A(n23234), .B(n23233), .Z(n23235) );
  AND U24862 ( .A(n23236), .B(n23235), .Z(n23353) );
  NAND U24863 ( .A(n23238), .B(n23237), .Z(n23242) );
  NAND U24864 ( .A(n23240), .B(n23239), .Z(n23241) );
  NAND U24865 ( .A(n23242), .B(n23241), .Z(n23359) );
  NAND U24866 ( .A(n23244), .B(n23243), .Z(n23248) );
  NANDN U24867 ( .A(n23246), .B(n23245), .Z(n23247) );
  NAND U24868 ( .A(n23248), .B(n23247), .Z(n23358) );
  XOR U24869 ( .A(n23359), .B(n23358), .Z(n23361) );
  AND U24870 ( .A(x[496]), .B(y[7914]), .Z(n24265) );
  NAND U24871 ( .A(n24265), .B(n23249), .Z(n23253) );
  NAND U24872 ( .A(n23251), .B(n23250), .Z(n23252) );
  NAND U24873 ( .A(n23253), .B(n23252), .Z(n23399) );
  AND U24874 ( .A(x[493]), .B(y[7921]), .Z(n24807) );
  NAND U24875 ( .A(n24807), .B(n23254), .Z(n23258) );
  NANDN U24876 ( .A(n23256), .B(n23255), .Z(n23257) );
  NAND U24877 ( .A(n23258), .B(n23257), .Z(n23444) );
  AND U24878 ( .A(y[7908]), .B(x[496]), .Z(n23260) );
  NAND U24879 ( .A(y[7914]), .B(x[490]), .Z(n23259) );
  XNOR U24880 ( .A(n23260), .B(n23259), .Z(n23405) );
  AND U24881 ( .A(x[482]), .B(y[7922]), .Z(n23406) );
  XOR U24882 ( .A(n23405), .B(n23406), .Z(n23442) );
  NAND U24883 ( .A(y[7915]), .B(x[489]), .Z(n23261) );
  XNOR U24884 ( .A(n23262), .B(n23261), .Z(n23381) );
  AND U24885 ( .A(x[494]), .B(y[7910]), .Z(n23382) );
  XOR U24886 ( .A(n23381), .B(n23382), .Z(n23441) );
  XOR U24887 ( .A(n23442), .B(n23441), .Z(n23443) );
  XOR U24888 ( .A(n23444), .B(n23443), .Z(n23398) );
  XOR U24889 ( .A(n23399), .B(n23398), .Z(n23401) );
  AND U24890 ( .A(x[491]), .B(y[7920]), .Z(n24419) );
  NAND U24891 ( .A(n23529), .B(n24419), .Z(n23266) );
  NANDN U24892 ( .A(n23264), .B(n23263), .Z(n23265) );
  NAND U24893 ( .A(n23266), .B(n23265), .Z(n23450) );
  AND U24894 ( .A(y[7913]), .B(x[491]), .Z(n23268) );
  NAND U24895 ( .A(y[7923]), .B(x[481]), .Z(n23267) );
  XNOR U24896 ( .A(n23268), .B(n23267), .Z(n23377) );
  AND U24897 ( .A(x[499]), .B(y[7905]), .Z(n23385) );
  XOR U24898 ( .A(o[244]), .B(n23385), .Z(n23376) );
  XOR U24899 ( .A(n23377), .B(n23376), .Z(n23448) );
  AND U24900 ( .A(x[480]), .B(y[7924]), .Z(n23429) );
  AND U24901 ( .A(x[500]), .B(y[7904]), .Z(n23430) );
  XOR U24902 ( .A(n23429), .B(n23430), .Z(n23432) );
  AND U24903 ( .A(o[243]), .B(n23269), .Z(n23431) );
  XOR U24904 ( .A(n23432), .B(n23431), .Z(n23447) );
  XOR U24905 ( .A(n23448), .B(n23447), .Z(n23449) );
  XOR U24906 ( .A(n23450), .B(n23449), .Z(n23400) );
  XOR U24907 ( .A(n23401), .B(n23400), .Z(n23360) );
  XNOR U24908 ( .A(n23361), .B(n23360), .Z(n23456) );
  NAND U24909 ( .A(x[486]), .B(y[7918]), .Z(n23365) );
  NANDN U24910 ( .A(n23365), .B(n23270), .Z(n23273) );
  NAND U24911 ( .A(n23271), .B(n23424), .Z(n23272) );
  NAND U24912 ( .A(n23273), .B(n23272), .Z(n23389) );
  NAND U24913 ( .A(n23275), .B(n23274), .Z(n23279) );
  NAND U24914 ( .A(n23277), .B(n23276), .Z(n23278) );
  NAND U24915 ( .A(n23279), .B(n23278), .Z(n23387) );
  AND U24916 ( .A(y[7906]), .B(x[498]), .Z(n23281) );
  NAND U24917 ( .A(y[7912]), .B(x[492]), .Z(n23280) );
  XNOR U24918 ( .A(n23281), .B(n23280), .Z(n23371) );
  AND U24919 ( .A(x[497]), .B(y[7907]), .Z(n23372) );
  XOR U24920 ( .A(n23371), .B(n23372), .Z(n23386) );
  XOR U24921 ( .A(n23387), .B(n23386), .Z(n23388) );
  XNOR U24922 ( .A(n23389), .B(n23388), .Z(n23393) );
  AND U24923 ( .A(y[7911]), .B(x[493]), .Z(n23283) );
  NAND U24924 ( .A(y[7921]), .B(x[483]), .Z(n23282) );
  XNOR U24925 ( .A(n23283), .B(n23282), .Z(n23411) );
  XNOR U24926 ( .A(n23411), .B(n23410), .Z(n23367) );
  AND U24927 ( .A(y[7919]), .B(x[485]), .Z(n23285) );
  NAND U24928 ( .A(y[7920]), .B(x[484]), .Z(n23284) );
  XNOR U24929 ( .A(n23285), .B(n23284), .Z(n23426) );
  AND U24930 ( .A(x[487]), .B(y[7917]), .Z(n23425) );
  XNOR U24931 ( .A(n23426), .B(n23425), .Z(n23364) );
  XOR U24932 ( .A(n23365), .B(n23364), .Z(n23366) );
  XNOR U24933 ( .A(n23367), .B(n23366), .Z(n23437) );
  AND U24934 ( .A(x[488]), .B(y[7922]), .Z(n24532) );
  AND U24935 ( .A(x[481]), .B(y[7915]), .Z(n23286) );
  NAND U24936 ( .A(n24532), .B(n23286), .Z(n23290) );
  NANDN U24937 ( .A(n23288), .B(n23287), .Z(n23289) );
  NAND U24938 ( .A(n23290), .B(n23289), .Z(n23436) );
  NAND U24939 ( .A(x[497]), .B(y[7913]), .Z(n24273) );
  NANDN U24940 ( .A(n24273), .B(n23291), .Z(n23295) );
  NAND U24941 ( .A(n23293), .B(n23292), .Z(n23294) );
  NAND U24942 ( .A(n23295), .B(n23294), .Z(n23435) );
  XOR U24943 ( .A(n23436), .B(n23435), .Z(n23438) );
  XNOR U24944 ( .A(n23437), .B(n23438), .Z(n23392) );
  XOR U24945 ( .A(n23393), .B(n23392), .Z(n23394) );
  NAND U24946 ( .A(n23297), .B(n23296), .Z(n23301) );
  NAND U24947 ( .A(n23299), .B(n23298), .Z(n23300) );
  AND U24948 ( .A(n23301), .B(n23300), .Z(n23395) );
  XOR U24949 ( .A(n23394), .B(n23395), .Z(n23453) );
  NAND U24950 ( .A(n23303), .B(n23302), .Z(n23307) );
  NAND U24951 ( .A(n23305), .B(n23304), .Z(n23306) );
  AND U24952 ( .A(n23307), .B(n23306), .Z(n23454) );
  XOR U24953 ( .A(n23453), .B(n23454), .Z(n23455) );
  XNOR U24954 ( .A(n23456), .B(n23455), .Z(n23460) );
  NAND U24955 ( .A(n23309), .B(n23308), .Z(n23313) );
  NAND U24956 ( .A(n23311), .B(n23310), .Z(n23312) );
  AND U24957 ( .A(n23313), .B(n23312), .Z(n23468) );
  NAND U24958 ( .A(n23315), .B(n23314), .Z(n23319) );
  NAND U24959 ( .A(n23317), .B(n23316), .Z(n23318) );
  AND U24960 ( .A(n23319), .B(n23318), .Z(n23466) );
  NAND U24961 ( .A(n23321), .B(n23320), .Z(n23325) );
  NAND U24962 ( .A(n23323), .B(n23322), .Z(n23324) );
  AND U24963 ( .A(n23325), .B(n23324), .Z(n23465) );
  XNOR U24964 ( .A(n23468), .B(n23467), .Z(n23459) );
  XOR U24965 ( .A(n23460), .B(n23459), .Z(n23462) );
  NAND U24966 ( .A(n23327), .B(n23326), .Z(n23331) );
  NAND U24967 ( .A(n23329), .B(n23328), .Z(n23330) );
  AND U24968 ( .A(n23331), .B(n23330), .Z(n23461) );
  XNOR U24969 ( .A(n23462), .B(n23461), .Z(n23348) );
  NANDN U24970 ( .A(n23333), .B(n23332), .Z(n23337) );
  NANDN U24971 ( .A(n23335), .B(n23334), .Z(n23336) );
  AND U24972 ( .A(n23337), .B(n23336), .Z(n23345) );
  NAND U24973 ( .A(n23339), .B(n23338), .Z(n23343) );
  NAND U24974 ( .A(n23341), .B(n23340), .Z(n23342) );
  AND U24975 ( .A(n23343), .B(n23342), .Z(n23346) );
  XOR U24976 ( .A(n23345), .B(n23346), .Z(n23347) );
  XOR U24977 ( .A(n23348), .B(n23347), .Z(n23354) );
  XNOR U24978 ( .A(n23353), .B(n23354), .Z(n23344) );
  XOR U24979 ( .A(n23351), .B(n23344), .Z(N501) );
  NAND U24980 ( .A(n23346), .B(n23345), .Z(n23350) );
  NAND U24981 ( .A(n23348), .B(n23347), .Z(n23349) );
  NAND U24982 ( .A(n23350), .B(n23349), .Z(n23595) );
  IV U24983 ( .A(n23595), .Z(n23593) );
  OR U24984 ( .A(n23353), .B(n23351), .Z(n23357) );
  ANDN U24985 ( .B(n23353), .A(n23352), .Z(n23355) );
  OR U24986 ( .A(n23355), .B(n23354), .Z(n23356) );
  AND U24987 ( .A(n23357), .B(n23356), .Z(n23594) );
  NAND U24988 ( .A(n23359), .B(n23358), .Z(n23363) );
  NAND U24989 ( .A(n23361), .B(n23360), .Z(n23362) );
  NAND U24990 ( .A(n23363), .B(n23362), .Z(n23481) );
  NAND U24991 ( .A(n23365), .B(n23364), .Z(n23369) );
  NAND U24992 ( .A(n23367), .B(n23366), .Z(n23368) );
  NAND U24993 ( .A(n23369), .B(n23368), .Z(n23570) );
  AND U24994 ( .A(x[498]), .B(y[7912]), .Z(n24272) );
  NAND U24995 ( .A(n24272), .B(n23370), .Z(n23374) );
  NAND U24996 ( .A(n23372), .B(n23371), .Z(n23373) );
  NAND U24997 ( .A(n23374), .B(n23373), .Z(n23552) );
  AND U24998 ( .A(x[491]), .B(y[7923]), .Z(n24864) );
  AND U24999 ( .A(x[481]), .B(y[7913]), .Z(n23375) );
  NAND U25000 ( .A(n24864), .B(n23375), .Z(n23379) );
  NAND U25001 ( .A(n23377), .B(n23376), .Z(n23378) );
  NAND U25002 ( .A(n23379), .B(n23378), .Z(n23551) );
  XOR U25003 ( .A(n23552), .B(n23551), .Z(n23554) );
  AND U25004 ( .A(x[495]), .B(y[7915]), .Z(n24260) );
  NAND U25005 ( .A(n24260), .B(n23380), .Z(n23384) );
  NAND U25006 ( .A(n23382), .B(n23381), .Z(n23383) );
  NAND U25007 ( .A(n23384), .B(n23383), .Z(n23516) );
  AND U25008 ( .A(x[480]), .B(y[7925]), .Z(n23535) );
  AND U25009 ( .A(x[501]), .B(y[7904]), .Z(n23536) );
  XOR U25010 ( .A(n23535), .B(n23536), .Z(n23538) );
  AND U25011 ( .A(o[244]), .B(n23385), .Z(n23537) );
  XOR U25012 ( .A(n23538), .B(n23537), .Z(n23514) );
  AND U25013 ( .A(x[485]), .B(y[7920]), .Z(n23522) );
  AND U25014 ( .A(x[496]), .B(y[7909]), .Z(n23521) );
  XOR U25015 ( .A(n23522), .B(n23521), .Z(n23520) );
  AND U25016 ( .A(x[495]), .B(y[7910]), .Z(n23519) );
  XOR U25017 ( .A(n23520), .B(n23519), .Z(n23513) );
  XOR U25018 ( .A(n23514), .B(n23513), .Z(n23515) );
  XOR U25019 ( .A(n23516), .B(n23515), .Z(n23553) );
  XNOR U25020 ( .A(n23554), .B(n23553), .Z(n23569) );
  XOR U25021 ( .A(n23570), .B(n23569), .Z(n23572) );
  NAND U25022 ( .A(n23387), .B(n23386), .Z(n23391) );
  NAND U25023 ( .A(n23389), .B(n23388), .Z(n23390) );
  AND U25024 ( .A(n23391), .B(n23390), .Z(n23571) );
  XNOR U25025 ( .A(n23572), .B(n23571), .Z(n23479) );
  NAND U25026 ( .A(n23393), .B(n23392), .Z(n23397) );
  NAND U25027 ( .A(n23395), .B(n23394), .Z(n23396) );
  AND U25028 ( .A(n23397), .B(n23396), .Z(n23478) );
  XOR U25029 ( .A(n23479), .B(n23478), .Z(n23480) );
  XNOR U25030 ( .A(n23481), .B(n23480), .Z(n23474) );
  NAND U25031 ( .A(n23399), .B(n23398), .Z(n23403) );
  NAND U25032 ( .A(n23401), .B(n23400), .Z(n23402) );
  NAND U25033 ( .A(n23403), .B(n23402), .Z(n23578) );
  NAND U25034 ( .A(n24265), .B(n23404), .Z(n23408) );
  NAND U25035 ( .A(n23406), .B(n23405), .Z(n23407) );
  NAND U25036 ( .A(n23408), .B(n23407), .Z(n23485) );
  NAND U25037 ( .A(n24807), .B(n23409), .Z(n23413) );
  NAND U25038 ( .A(n23411), .B(n23410), .Z(n23412) );
  NAND U25039 ( .A(n23413), .B(n23412), .Z(n23566) );
  AND U25040 ( .A(y[7906]), .B(x[499]), .Z(n23415) );
  NAND U25041 ( .A(y[7914]), .B(x[491]), .Z(n23414) );
  XNOR U25042 ( .A(n23415), .B(n23414), .Z(n23504) );
  AND U25043 ( .A(x[500]), .B(y[7905]), .Z(n23534) );
  XOR U25044 ( .A(o[245]), .B(n23534), .Z(n23503) );
  XOR U25045 ( .A(n23504), .B(n23503), .Z(n23564) );
  AND U25046 ( .A(y[7907]), .B(x[498]), .Z(n23417) );
  NAND U25047 ( .A(y[7915]), .B(x[490]), .Z(n23416) );
  XNOR U25048 ( .A(n23417), .B(n23416), .Z(n23542) );
  AND U25049 ( .A(x[481]), .B(y[7924]), .Z(n23543) );
  XOR U25050 ( .A(n23542), .B(n23543), .Z(n23563) );
  XOR U25051 ( .A(n23564), .B(n23563), .Z(n23565) );
  XOR U25052 ( .A(n23566), .B(n23565), .Z(n23484) );
  XOR U25053 ( .A(n23485), .B(n23484), .Z(n23487) );
  AND U25054 ( .A(x[487]), .B(y[7918]), .Z(n23751) );
  AND U25055 ( .A(y[7919]), .B(x[486]), .Z(n23419) );
  NAND U25056 ( .A(y[7911]), .B(x[494]), .Z(n23418) );
  XNOR U25057 ( .A(n23419), .B(n23418), .Z(n23546) );
  XNOR U25058 ( .A(n23751), .B(n23546), .Z(n23493) );
  NAND U25059 ( .A(x[489]), .B(y[7916]), .Z(n23491) );
  NAND U25060 ( .A(x[488]), .B(y[7917]), .Z(n23490) );
  XOR U25061 ( .A(n23491), .B(n23490), .Z(n23492) );
  XNOR U25062 ( .A(n23493), .B(n23492), .Z(n23509) );
  AND U25063 ( .A(y[7912]), .B(x[493]), .Z(n23421) );
  NAND U25064 ( .A(y[7922]), .B(x[483]), .Z(n23420) );
  XNOR U25065 ( .A(n23421), .B(n23420), .Z(n23530) );
  AND U25066 ( .A(x[484]), .B(y[7921]), .Z(n23531) );
  XOR U25067 ( .A(n23530), .B(n23531), .Z(n23508) );
  AND U25068 ( .A(y[7913]), .B(x[492]), .Z(n23423) );
  NAND U25069 ( .A(y[7908]), .B(x[497]), .Z(n23422) );
  XNOR U25070 ( .A(n23423), .B(n23422), .Z(n23496) );
  AND U25071 ( .A(x[482]), .B(y[7923]), .Z(n23497) );
  XOR U25072 ( .A(n23496), .B(n23497), .Z(n23507) );
  XOR U25073 ( .A(n23508), .B(n23507), .Z(n23510) );
  XOR U25074 ( .A(n23509), .B(n23510), .Z(n23560) );
  NAND U25075 ( .A(n23522), .B(n23424), .Z(n23428) );
  NAND U25076 ( .A(n23426), .B(n23425), .Z(n23427) );
  NAND U25077 ( .A(n23428), .B(n23427), .Z(n23558) );
  NAND U25078 ( .A(n23430), .B(n23429), .Z(n23434) );
  NAND U25079 ( .A(n23432), .B(n23431), .Z(n23433) );
  NAND U25080 ( .A(n23434), .B(n23433), .Z(n23557) );
  XOR U25081 ( .A(n23558), .B(n23557), .Z(n23559) );
  XOR U25082 ( .A(n23560), .B(n23559), .Z(n23486) );
  XOR U25083 ( .A(n23487), .B(n23486), .Z(n23576) );
  NAND U25084 ( .A(n23436), .B(n23435), .Z(n23440) );
  NAND U25085 ( .A(n23438), .B(n23437), .Z(n23439) );
  NAND U25086 ( .A(n23440), .B(n23439), .Z(n23583) );
  NAND U25087 ( .A(n23442), .B(n23441), .Z(n23446) );
  NAND U25088 ( .A(n23444), .B(n23443), .Z(n23445) );
  NAND U25089 ( .A(n23446), .B(n23445), .Z(n23582) );
  NAND U25090 ( .A(n23448), .B(n23447), .Z(n23452) );
  NAND U25091 ( .A(n23450), .B(n23449), .Z(n23451) );
  NAND U25092 ( .A(n23452), .B(n23451), .Z(n23581) );
  XOR U25093 ( .A(n23582), .B(n23581), .Z(n23584) );
  XOR U25094 ( .A(n23583), .B(n23584), .Z(n23575) );
  XOR U25095 ( .A(n23576), .B(n23575), .Z(n23577) );
  XNOR U25096 ( .A(n23578), .B(n23577), .Z(n23473) );
  NAND U25097 ( .A(n23454), .B(n23453), .Z(n23458) );
  NAND U25098 ( .A(n23456), .B(n23455), .Z(n23457) );
  NAND U25099 ( .A(n23458), .B(n23457), .Z(n23472) );
  XOR U25100 ( .A(n23473), .B(n23472), .Z(n23475) );
  XNOR U25101 ( .A(n23474), .B(n23475), .Z(n23589) );
  NAND U25102 ( .A(n23460), .B(n23459), .Z(n23464) );
  NAND U25103 ( .A(n23462), .B(n23461), .Z(n23463) );
  NAND U25104 ( .A(n23464), .B(n23463), .Z(n23588) );
  NANDN U25105 ( .A(n23466), .B(n23465), .Z(n23470) );
  NAND U25106 ( .A(n23468), .B(n23467), .Z(n23469) );
  AND U25107 ( .A(n23470), .B(n23469), .Z(n23587) );
  XOR U25108 ( .A(n23588), .B(n23587), .Z(n23590) );
  XOR U25109 ( .A(n23589), .B(n23590), .Z(n23596) );
  XNOR U25110 ( .A(n23594), .B(n23596), .Z(n23471) );
  XOR U25111 ( .A(n23593), .B(n23471), .Z(N502) );
  NAND U25112 ( .A(n23473), .B(n23472), .Z(n23477) );
  NAND U25113 ( .A(n23475), .B(n23474), .Z(n23476) );
  AND U25114 ( .A(n23477), .B(n23476), .Z(n23727) );
  NAND U25115 ( .A(n23479), .B(n23478), .Z(n23483) );
  NAND U25116 ( .A(n23481), .B(n23480), .Z(n23482) );
  NAND U25117 ( .A(n23483), .B(n23482), .Z(n23725) );
  NAND U25118 ( .A(n23485), .B(n23484), .Z(n23489) );
  NAND U25119 ( .A(n23487), .B(n23486), .Z(n23488) );
  AND U25120 ( .A(n23489), .B(n23488), .Z(n23718) );
  NAND U25121 ( .A(n23491), .B(n23490), .Z(n23495) );
  NAND U25122 ( .A(n23493), .B(n23492), .Z(n23494) );
  NAND U25123 ( .A(n23495), .B(n23494), .Z(n23712) );
  NANDN U25124 ( .A(n24273), .B(n23663), .Z(n23499) );
  NAND U25125 ( .A(n23497), .B(n23496), .Z(n23498) );
  NAND U25126 ( .A(n23499), .B(n23498), .Z(n23639) );
  AND U25127 ( .A(x[485]), .B(y[7921]), .Z(n23685) );
  AND U25128 ( .A(x[497]), .B(y[7909]), .Z(n23686) );
  XOR U25129 ( .A(n23685), .B(n23686), .Z(n23687) );
  AND U25130 ( .A(x[496]), .B(y[7910]), .Z(n23688) );
  XOR U25131 ( .A(n23687), .B(n23688), .Z(n23638) );
  AND U25132 ( .A(y[7908]), .B(x[498]), .Z(n23501) );
  NAND U25133 ( .A(y[7914]), .B(x[492]), .Z(n23500) );
  XNOR U25134 ( .A(n23501), .B(n23500), .Z(n23664) );
  AND U25135 ( .A(x[484]), .B(y[7922]), .Z(n23665) );
  XOR U25136 ( .A(n23664), .B(n23665), .Z(n23637) );
  XOR U25137 ( .A(n23638), .B(n23637), .Z(n23640) );
  XNOR U25138 ( .A(n23639), .B(n23640), .Z(n23709) );
  AND U25139 ( .A(x[499]), .B(y[7914]), .Z(n24701) );
  NAND U25140 ( .A(n24701), .B(n23502), .Z(n23506) );
  NAND U25141 ( .A(n23504), .B(n23503), .Z(n23505) );
  AND U25142 ( .A(n23506), .B(n23505), .Z(n23710) );
  XOR U25143 ( .A(n23709), .B(n23710), .Z(n23711) );
  XNOR U25144 ( .A(n23712), .B(n23711), .Z(n23715) );
  NAND U25145 ( .A(n23508), .B(n23507), .Z(n23512) );
  NAND U25146 ( .A(n23510), .B(n23509), .Z(n23511) );
  NAND U25147 ( .A(n23512), .B(n23511), .Z(n23698) );
  NAND U25148 ( .A(n23514), .B(n23513), .Z(n23518) );
  NAND U25149 ( .A(n23516), .B(n23515), .Z(n23517) );
  NAND U25150 ( .A(n23518), .B(n23517), .Z(n23697) );
  XOR U25151 ( .A(n23698), .B(n23697), .Z(n23700) );
  AND U25152 ( .A(n23520), .B(n23519), .Z(n23524) );
  NAND U25153 ( .A(n23522), .B(n23521), .Z(n23523) );
  NANDN U25154 ( .A(n23524), .B(n23523), .Z(n23660) );
  AND U25155 ( .A(y[7913]), .B(x[493]), .Z(n23526) );
  NAND U25156 ( .A(y[7906]), .B(x[500]), .Z(n23525) );
  XNOR U25157 ( .A(n23526), .B(n23525), .Z(n23681) );
  AND U25158 ( .A(x[482]), .B(y[7924]), .Z(n23682) );
  XOR U25159 ( .A(n23681), .B(n23682), .Z(n23658) );
  AND U25160 ( .A(y[7920]), .B(x[486]), .Z(n23528) );
  NAND U25161 ( .A(y[7911]), .B(x[495]), .Z(n23527) );
  XNOR U25162 ( .A(n23528), .B(n23527), .Z(n23693) );
  XOR U25163 ( .A(n23658), .B(n23657), .Z(n23659) );
  XOR U25164 ( .A(n23660), .B(n23659), .Z(n23704) );
  AND U25165 ( .A(x[493]), .B(y[7922]), .Z(n24900) );
  NAND U25166 ( .A(n23529), .B(n24900), .Z(n23533) );
  NAND U25167 ( .A(n23531), .B(n23530), .Z(n23532) );
  NAND U25168 ( .A(n23533), .B(n23532), .Z(n23628) );
  AND U25169 ( .A(x[481]), .B(y[7925]), .Z(n23651) );
  XOR U25170 ( .A(n23652), .B(n23651), .Z(n23650) );
  AND U25171 ( .A(o[245]), .B(n23534), .Z(n23649) );
  XOR U25172 ( .A(n23650), .B(n23649), .Z(n23626) );
  AND U25173 ( .A(x[494]), .B(y[7912]), .Z(n23643) );
  NAND U25174 ( .A(x[483]), .B(y[7923]), .Z(n23644) );
  NAND U25175 ( .A(x[499]), .B(y[7907]), .Z(n23646) );
  XOR U25176 ( .A(n23626), .B(n23625), .Z(n23627) );
  XOR U25177 ( .A(n23628), .B(n23627), .Z(n23703) );
  XOR U25178 ( .A(n23704), .B(n23703), .Z(n23706) );
  NAND U25179 ( .A(n23536), .B(n23535), .Z(n23540) );
  NAND U25180 ( .A(n23538), .B(n23537), .Z(n23539) );
  NAND U25181 ( .A(n23540), .B(n23539), .Z(n23620) );
  AND U25182 ( .A(x[498]), .B(y[7915]), .Z(n24704) );
  NAND U25183 ( .A(n24704), .B(n23541), .Z(n23545) );
  NAND U25184 ( .A(n23543), .B(n23542), .Z(n23544) );
  NAND U25185 ( .A(n23545), .B(n23544), .Z(n23619) );
  XOR U25186 ( .A(n23620), .B(n23619), .Z(n23622) );
  AND U25187 ( .A(x[494]), .B(y[7919]), .Z(n24714) );
  NAND U25188 ( .A(n24714), .B(n23692), .Z(n23548) );
  NAND U25189 ( .A(n23751), .B(n23546), .Z(n23547) );
  NAND U25190 ( .A(n23548), .B(n23547), .Z(n23634) );
  AND U25191 ( .A(x[480]), .B(y[7926]), .Z(n23668) );
  NAND U25192 ( .A(x[502]), .B(y[7904]), .Z(n23669) );
  NAND U25193 ( .A(x[501]), .B(y[7905]), .Z(n23691) );
  XOR U25194 ( .A(n23671), .B(n23670), .Z(n23632) );
  AND U25195 ( .A(y[7919]), .B(x[487]), .Z(n23550) );
  NAND U25196 ( .A(y[7918]), .B(x[488]), .Z(n23549) );
  XNOR U25197 ( .A(n23550), .B(n23549), .Z(n23674) );
  XOR U25198 ( .A(n23632), .B(n23631), .Z(n23633) );
  XOR U25199 ( .A(n23634), .B(n23633), .Z(n23621) );
  XOR U25200 ( .A(n23622), .B(n23621), .Z(n23705) );
  XOR U25201 ( .A(n23706), .B(n23705), .Z(n23699) );
  XOR U25202 ( .A(n23700), .B(n23699), .Z(n23716) );
  XOR U25203 ( .A(n23715), .B(n23716), .Z(n23717) );
  NAND U25204 ( .A(n23552), .B(n23551), .Z(n23556) );
  NAND U25205 ( .A(n23554), .B(n23553), .Z(n23555) );
  NAND U25206 ( .A(n23556), .B(n23555), .Z(n23616) );
  NAND U25207 ( .A(n23558), .B(n23557), .Z(n23562) );
  NAND U25208 ( .A(n23560), .B(n23559), .Z(n23561) );
  NAND U25209 ( .A(n23562), .B(n23561), .Z(n23614) );
  NAND U25210 ( .A(n23564), .B(n23563), .Z(n23568) );
  NAND U25211 ( .A(n23566), .B(n23565), .Z(n23567) );
  NAND U25212 ( .A(n23568), .B(n23567), .Z(n23613) );
  XOR U25213 ( .A(n23614), .B(n23613), .Z(n23615) );
  XNOR U25214 ( .A(n23616), .B(n23615), .Z(n23608) );
  NAND U25215 ( .A(n23570), .B(n23569), .Z(n23574) );
  NAND U25216 ( .A(n23572), .B(n23571), .Z(n23573) );
  NAND U25217 ( .A(n23574), .B(n23573), .Z(n23607) );
  XOR U25218 ( .A(n23608), .B(n23607), .Z(n23610) );
  XNOR U25219 ( .A(n23609), .B(n23610), .Z(n23603) );
  NAND U25220 ( .A(n23576), .B(n23575), .Z(n23580) );
  NAND U25221 ( .A(n23578), .B(n23577), .Z(n23579) );
  NAND U25222 ( .A(n23580), .B(n23579), .Z(n23602) );
  NAND U25223 ( .A(n23582), .B(n23581), .Z(n23586) );
  NAND U25224 ( .A(n23584), .B(n23583), .Z(n23585) );
  NAND U25225 ( .A(n23586), .B(n23585), .Z(n23601) );
  XOR U25226 ( .A(n23602), .B(n23601), .Z(n23604) );
  XOR U25227 ( .A(n23603), .B(n23604), .Z(n23724) );
  XOR U25228 ( .A(n23725), .B(n23724), .Z(n23726) );
  XNOR U25229 ( .A(n23727), .B(n23726), .Z(n23723) );
  NAND U25230 ( .A(n23588), .B(n23587), .Z(n23592) );
  NAND U25231 ( .A(n23590), .B(n23589), .Z(n23591) );
  NAND U25232 ( .A(n23592), .B(n23591), .Z(n23722) );
  NANDN U25233 ( .A(n23593), .B(n23594), .Z(n23599) );
  NOR U25234 ( .A(n23595), .B(n23594), .Z(n23597) );
  OR U25235 ( .A(n23597), .B(n23596), .Z(n23598) );
  AND U25236 ( .A(n23599), .B(n23598), .Z(n23721) );
  XOR U25237 ( .A(n23722), .B(n23721), .Z(n23600) );
  XNOR U25238 ( .A(n23723), .B(n23600), .Z(N503) );
  NAND U25239 ( .A(n23602), .B(n23601), .Z(n23606) );
  NAND U25240 ( .A(n23604), .B(n23603), .Z(n23605) );
  AND U25241 ( .A(n23606), .B(n23605), .Z(n23872) );
  NAND U25242 ( .A(n23608), .B(n23607), .Z(n23612) );
  NAND U25243 ( .A(n23610), .B(n23609), .Z(n23611) );
  NAND U25244 ( .A(n23612), .B(n23611), .Z(n23870) );
  NAND U25245 ( .A(n23614), .B(n23613), .Z(n23618) );
  NAND U25246 ( .A(n23616), .B(n23615), .Z(n23617) );
  NAND U25247 ( .A(n23618), .B(n23617), .Z(n23847) );
  NAND U25248 ( .A(n23620), .B(n23619), .Z(n23624) );
  NAND U25249 ( .A(n23622), .B(n23621), .Z(n23623) );
  NAND U25250 ( .A(n23624), .B(n23623), .Z(n23841) );
  NAND U25251 ( .A(n23626), .B(n23625), .Z(n23630) );
  NAND U25252 ( .A(n23628), .B(n23627), .Z(n23629) );
  NAND U25253 ( .A(n23630), .B(n23629), .Z(n23839) );
  NAND U25254 ( .A(n23632), .B(n23631), .Z(n23636) );
  NAND U25255 ( .A(n23634), .B(n23633), .Z(n23635) );
  NAND U25256 ( .A(n23636), .B(n23635), .Z(n23838) );
  XOR U25257 ( .A(n23839), .B(n23838), .Z(n23840) );
  XOR U25258 ( .A(n23841), .B(n23840), .Z(n23859) );
  NAND U25259 ( .A(n23638), .B(n23637), .Z(n23642) );
  NAND U25260 ( .A(n23640), .B(n23639), .Z(n23641) );
  NAND U25261 ( .A(n23642), .B(n23641), .Z(n23857) );
  NANDN U25262 ( .A(n23644), .B(n23643), .Z(n23648) );
  NANDN U25263 ( .A(n23646), .B(n23645), .Z(n23647) );
  NAND U25264 ( .A(n23648), .B(n23647), .Z(n23785) );
  AND U25265 ( .A(n23650), .B(n23649), .Z(n23654) );
  NAND U25266 ( .A(n23652), .B(n23651), .Z(n23653) );
  NANDN U25267 ( .A(n23654), .B(n23653), .Z(n23784) );
  XOR U25268 ( .A(n23785), .B(n23784), .Z(n23787) );
  AND U25269 ( .A(y[7920]), .B(x[487]), .Z(n23656) );
  NAND U25270 ( .A(y[7918]), .B(x[489]), .Z(n23655) );
  XNOR U25271 ( .A(n23656), .B(n23655), .Z(n23752) );
  NAND U25272 ( .A(x[490]), .B(y[7917]), .Z(n23791) );
  AND U25273 ( .A(x[486]), .B(y[7921]), .Z(n23743) );
  NAND U25274 ( .A(x[495]), .B(y[7912]), .Z(n23744) );
  NAND U25275 ( .A(x[491]), .B(y[7916]), .Z(n23746) );
  XOR U25276 ( .A(n23793), .B(n23792), .Z(n23786) );
  XOR U25277 ( .A(n23787), .B(n23786), .Z(n23856) );
  XOR U25278 ( .A(n23857), .B(n23856), .Z(n23858) );
  XOR U25279 ( .A(n23859), .B(n23858), .Z(n23845) );
  NAND U25280 ( .A(n23658), .B(n23657), .Z(n23662) );
  NAND U25281 ( .A(n23660), .B(n23659), .Z(n23661) );
  NAND U25282 ( .A(n23662), .B(n23661), .Z(n23779) );
  NAND U25283 ( .A(x[498]), .B(y[7914]), .Z(n24563) );
  NANDN U25284 ( .A(n24563), .B(n23663), .Z(n23667) );
  NAND U25285 ( .A(n23665), .B(n23664), .Z(n23666) );
  NAND U25286 ( .A(n23667), .B(n23666), .Z(n23827) );
  NANDN U25287 ( .A(n23669), .B(n23668), .Z(n23673) );
  NAND U25288 ( .A(n23671), .B(n23670), .Z(n23672) );
  NAND U25289 ( .A(n23673), .B(n23672), .Z(n23826) );
  XOR U25290 ( .A(n23827), .B(n23826), .Z(n23828) );
  NANDN U25291 ( .A(n23753), .B(n23751), .Z(n23677) );
  NANDN U25292 ( .A(n23675), .B(n23674), .Z(n23676) );
  NAND U25293 ( .A(n23677), .B(n23676), .Z(n23822) );
  AND U25294 ( .A(x[480]), .B(y[7927]), .Z(n23762) );
  NAND U25295 ( .A(x[503]), .B(y[7904]), .Z(n23763) );
  NAND U25296 ( .A(x[502]), .B(y[7905]), .Z(n23742) );
  XOR U25297 ( .A(n23765), .B(n23764), .Z(n23821) );
  NAND U25298 ( .A(y[7907]), .B(x[500]), .Z(n23678) );
  XNOR U25299 ( .A(n23679), .B(n23678), .Z(n23738) );
  NAND U25300 ( .A(x[499]), .B(y[7908]), .Z(n23739) );
  XOR U25301 ( .A(n23821), .B(n23820), .Z(n23823) );
  XOR U25302 ( .A(n23822), .B(n23823), .Z(n23829) );
  XOR U25303 ( .A(n23828), .B(n23829), .Z(n23778) );
  XOR U25304 ( .A(n23779), .B(n23778), .Z(n23781) );
  NAND U25305 ( .A(x[500]), .B(y[7913]), .Z(n24726) );
  AND U25306 ( .A(x[493]), .B(y[7906]), .Z(n23680) );
  NANDN U25307 ( .A(n24726), .B(n23680), .Z(n23684) );
  NAND U25308 ( .A(n23682), .B(n23681), .Z(n23683) );
  NAND U25309 ( .A(n23684), .B(n23683), .Z(n23773) );
  NAND U25310 ( .A(n23686), .B(n23685), .Z(n23690) );
  NAND U25311 ( .A(n23688), .B(n23687), .Z(n23689) );
  NAND U25312 ( .A(n23690), .B(n23689), .Z(n23834) );
  AND U25313 ( .A(x[493]), .B(y[7914]), .Z(n23809) );
  AND U25314 ( .A(x[482]), .B(y[7925]), .Z(n23808) );
  XOR U25315 ( .A(n23809), .B(n23808), .Z(n23811) );
  AND U25316 ( .A(x[501]), .B(y[7906]), .Z(n23810) );
  XOR U25317 ( .A(n23811), .B(n23810), .Z(n23833) );
  ANDN U25318 ( .B(o[246]), .A(n23691), .Z(n23759) );
  AND U25319 ( .A(x[492]), .B(y[7915]), .Z(n23757) );
  AND U25320 ( .A(x[481]), .B(y[7926]), .Z(n23756) );
  XOR U25321 ( .A(n23757), .B(n23756), .Z(n23758) );
  XOR U25322 ( .A(n23759), .B(n23758), .Z(n23832) );
  XOR U25323 ( .A(n23833), .B(n23832), .Z(n23835) );
  XOR U25324 ( .A(n23834), .B(n23835), .Z(n23772) );
  XOR U25325 ( .A(n23773), .B(n23772), .Z(n23775) );
  AND U25326 ( .A(x[495]), .B(y[7920]), .Z(n24894) );
  NAND U25327 ( .A(n24894), .B(n23692), .Z(n23696) );
  NANDN U25328 ( .A(n23694), .B(n23693), .Z(n23695) );
  NAND U25329 ( .A(n23696), .B(n23695), .Z(n23816) );
  AND U25330 ( .A(x[494]), .B(y[7913]), .Z(n23803) );
  AND U25331 ( .A(x[483]), .B(y[7924]), .Z(n23802) );
  XOR U25332 ( .A(n23803), .B(n23802), .Z(n23805) );
  AND U25333 ( .A(x[484]), .B(y[7923]), .Z(n23804) );
  XOR U25334 ( .A(n23805), .B(n23804), .Z(n23815) );
  AND U25335 ( .A(x[485]), .B(y[7922]), .Z(n23797) );
  AND U25336 ( .A(x[498]), .B(y[7909]), .Z(n23796) );
  XOR U25337 ( .A(n23797), .B(n23796), .Z(n23799) );
  AND U25338 ( .A(x[497]), .B(y[7910]), .Z(n23798) );
  XOR U25339 ( .A(n23799), .B(n23798), .Z(n23814) );
  XOR U25340 ( .A(n23815), .B(n23814), .Z(n23817) );
  XOR U25341 ( .A(n23816), .B(n23817), .Z(n23774) );
  XOR U25342 ( .A(n23775), .B(n23774), .Z(n23780) );
  XOR U25343 ( .A(n23781), .B(n23780), .Z(n23844) );
  XOR U25344 ( .A(n23845), .B(n23844), .Z(n23846) );
  XNOR U25345 ( .A(n23847), .B(n23846), .Z(n23733) );
  NAND U25346 ( .A(n23698), .B(n23697), .Z(n23702) );
  NAND U25347 ( .A(n23700), .B(n23699), .Z(n23701) );
  NAND U25348 ( .A(n23702), .B(n23701), .Z(n23853) );
  NAND U25349 ( .A(n23704), .B(n23703), .Z(n23708) );
  NAND U25350 ( .A(n23706), .B(n23705), .Z(n23707) );
  NAND U25351 ( .A(n23708), .B(n23707), .Z(n23851) );
  NAND U25352 ( .A(n23710), .B(n23709), .Z(n23714) );
  NAND U25353 ( .A(n23712), .B(n23711), .Z(n23713) );
  AND U25354 ( .A(n23714), .B(n23713), .Z(n23850) );
  XOR U25355 ( .A(n23851), .B(n23850), .Z(n23852) );
  XNOR U25356 ( .A(n23853), .B(n23852), .Z(n23731) );
  NAND U25357 ( .A(n23716), .B(n23715), .Z(n23720) );
  NANDN U25358 ( .A(n23718), .B(n23717), .Z(n23719) );
  AND U25359 ( .A(n23720), .B(n23719), .Z(n23732) );
  XOR U25360 ( .A(n23731), .B(n23732), .Z(n23734) );
  XOR U25361 ( .A(n23733), .B(n23734), .Z(n23869) );
  XOR U25362 ( .A(n23870), .B(n23869), .Z(n23871) );
  XNOR U25363 ( .A(n23872), .B(n23871), .Z(n23865) );
  NAND U25364 ( .A(n23725), .B(n23724), .Z(n23729) );
  NAND U25365 ( .A(n23727), .B(n23726), .Z(n23728) );
  AND U25366 ( .A(n23729), .B(n23728), .Z(n23864) );
  IV U25367 ( .A(n23864), .Z(n23862) );
  XOR U25368 ( .A(n23863), .B(n23862), .Z(n23730) );
  XNOR U25369 ( .A(n23865), .B(n23730), .Z(N504) );
  NAND U25370 ( .A(n23732), .B(n23731), .Z(n23736) );
  NAND U25371 ( .A(n23734), .B(n23733), .Z(n23735) );
  AND U25372 ( .A(n23736), .B(n23735), .Z(n23879) );
  AND U25373 ( .A(x[500]), .B(y[7911]), .Z(n23737) );
  NAND U25374 ( .A(n23737), .B(n23982), .Z(n23741) );
  NANDN U25375 ( .A(n23739), .B(n23738), .Z(n23740) );
  NAND U25376 ( .A(n23741), .B(n23740), .Z(n24007) );
  AND U25377 ( .A(x[502]), .B(y[7906]), .Z(n23913) );
  XOR U25378 ( .A(n23914), .B(n23913), .Z(n23916) );
  NAND U25379 ( .A(x[482]), .B(y[7926]), .Z(n23915) );
  ANDN U25380 ( .B(o[247]), .A(n23742), .Z(n23920) );
  AND U25381 ( .A(x[481]), .B(y[7927]), .Z(n23921) );
  XOR U25382 ( .A(n23922), .B(n23921), .Z(n23919) );
  XOR U25383 ( .A(n23920), .B(n23919), .Z(n24005) );
  XOR U25384 ( .A(n24006), .B(n24005), .Z(n24008) );
  XOR U25385 ( .A(n24007), .B(n24008), .Z(n23953) );
  NANDN U25386 ( .A(n23744), .B(n23743), .Z(n23748) );
  NANDN U25387 ( .A(n23746), .B(n23745), .Z(n23747) );
  NAND U25388 ( .A(n23748), .B(n23747), .Z(n24001) );
  AND U25389 ( .A(y[7912]), .B(x[496]), .Z(n23750) );
  NAND U25390 ( .A(y[7907]), .B(x[501]), .Z(n23749) );
  XNOR U25391 ( .A(n23750), .B(n23749), .Z(n23983) );
  NAND U25392 ( .A(x[485]), .B(y[7923]), .Z(n23984) );
  AND U25393 ( .A(x[486]), .B(y[7922]), .Z(n24227) );
  NAND U25394 ( .A(x[500]), .B(y[7908]), .Z(n24130) );
  AND U25395 ( .A(x[499]), .B(y[7909]), .Z(n23989) );
  XOR U25396 ( .A(n23990), .B(n23989), .Z(n23999) );
  XOR U25397 ( .A(n24000), .B(n23999), .Z(n24002) );
  XOR U25398 ( .A(n24001), .B(n24002), .Z(n23979) );
  NANDN U25399 ( .A(n23932), .B(n23751), .Z(n23755) );
  NANDN U25400 ( .A(n23753), .B(n23752), .Z(n23754) );
  NAND U25401 ( .A(n23755), .B(n23754), .Z(n23977) );
  NAND U25402 ( .A(n23757), .B(n23756), .Z(n23761) );
  NAND U25403 ( .A(n23759), .B(n23758), .Z(n23760) );
  NAND U25404 ( .A(n23761), .B(n23760), .Z(n23976) );
  XOR U25405 ( .A(n23977), .B(n23976), .Z(n23978) );
  XOR U25406 ( .A(n23979), .B(n23978), .Z(n23952) );
  XOR U25407 ( .A(n23953), .B(n23952), .Z(n23955) );
  NANDN U25408 ( .A(n23763), .B(n23762), .Z(n23767) );
  NAND U25409 ( .A(n23765), .B(n23764), .Z(n23766) );
  NAND U25410 ( .A(n23767), .B(n23766), .Z(n23934) );
  AND U25411 ( .A(x[483]), .B(y[7925]), .Z(n23940) );
  XOR U25412 ( .A(n23941), .B(n23940), .Z(n23943) );
  NAND U25413 ( .A(x[484]), .B(y[7924]), .Z(n23942) );
  XOR U25414 ( .A(n23934), .B(n23935), .Z(n23937) );
  AND U25415 ( .A(y[7919]), .B(x[489]), .Z(n23769) );
  NAND U25416 ( .A(y[7918]), .B(x[490]), .Z(n23768) );
  XNOR U25417 ( .A(n23769), .B(n23768), .Z(n23905) );
  AND U25418 ( .A(y[7914]), .B(x[494]), .Z(n23771) );
  NAND U25419 ( .A(y[7920]), .B(x[488]), .Z(n23770) );
  XNOR U25420 ( .A(n23771), .B(n23770), .Z(n23909) );
  NAND U25421 ( .A(x[491]), .B(y[7917]), .Z(n23910) );
  XOR U25422 ( .A(n23905), .B(n23904), .Z(n23936) );
  XOR U25423 ( .A(n23937), .B(n23936), .Z(n23954) );
  XOR U25424 ( .A(n23955), .B(n23954), .Z(n23898) );
  NAND U25425 ( .A(n23773), .B(n23772), .Z(n23777) );
  NAND U25426 ( .A(n23775), .B(n23774), .Z(n23776) );
  AND U25427 ( .A(n23777), .B(n23776), .Z(n23897) );
  NAND U25428 ( .A(n23779), .B(n23778), .Z(n23783) );
  NAND U25429 ( .A(n23781), .B(n23780), .Z(n23782) );
  NAND U25430 ( .A(n23783), .B(n23782), .Z(n23900) );
  NAND U25431 ( .A(n23785), .B(n23784), .Z(n23789) );
  NAND U25432 ( .A(n23787), .B(n23786), .Z(n23788) );
  AND U25433 ( .A(n23789), .B(n23788), .Z(n23961) );
  NANDN U25434 ( .A(n23791), .B(n23790), .Z(n23795) );
  NAND U25435 ( .A(n23793), .B(n23792), .Z(n23794) );
  AND U25436 ( .A(n23795), .B(n23794), .Z(n23959) );
  NAND U25437 ( .A(n23797), .B(n23796), .Z(n23801) );
  NAND U25438 ( .A(n23799), .B(n23798), .Z(n23800) );
  NAND U25439 ( .A(n23801), .B(n23800), .Z(n23995) );
  AND U25440 ( .A(x[480]), .B(y[7928]), .Z(n23946) );
  NAND U25441 ( .A(x[504]), .B(y[7904]), .Z(n23947) );
  NAND U25442 ( .A(x[503]), .B(y[7905]), .Z(n23933) );
  XOR U25443 ( .A(n23949), .B(n23948), .Z(n23994) );
  AND U25444 ( .A(x[487]), .B(y[7921]), .Z(n23925) );
  NAND U25445 ( .A(x[498]), .B(y[7910]), .Z(n23926) );
  AND U25446 ( .A(x[497]), .B(y[7911]), .Z(n23927) );
  XOR U25447 ( .A(n23928), .B(n23927), .Z(n23993) );
  XOR U25448 ( .A(n23994), .B(n23993), .Z(n23996) );
  XOR U25449 ( .A(n23995), .B(n23996), .Z(n23972) );
  NAND U25450 ( .A(n23803), .B(n23802), .Z(n23807) );
  NAND U25451 ( .A(n23805), .B(n23804), .Z(n23806) );
  NAND U25452 ( .A(n23807), .B(n23806), .Z(n23971) );
  NAND U25453 ( .A(n23809), .B(n23808), .Z(n23813) );
  NAND U25454 ( .A(n23811), .B(n23810), .Z(n23812) );
  NAND U25455 ( .A(n23813), .B(n23812), .Z(n23970) );
  XNOR U25456 ( .A(n23971), .B(n23970), .Z(n23973) );
  NAND U25457 ( .A(n23815), .B(n23814), .Z(n23819) );
  NAND U25458 ( .A(n23817), .B(n23816), .Z(n23818) );
  AND U25459 ( .A(n23819), .B(n23818), .Z(n24012) );
  NAND U25460 ( .A(n23821), .B(n23820), .Z(n23825) );
  NAND U25461 ( .A(n23823), .B(n23822), .Z(n23824) );
  AND U25462 ( .A(n23825), .B(n23824), .Z(n24011) );
  XOR U25463 ( .A(n24012), .B(n24011), .Z(n24014) );
  NAND U25464 ( .A(n23827), .B(n23826), .Z(n23831) );
  NAND U25465 ( .A(n23829), .B(n23828), .Z(n23830) );
  AND U25466 ( .A(n23831), .B(n23830), .Z(n24013) );
  XOR U25467 ( .A(n24014), .B(n24013), .Z(n23964) );
  NAND U25468 ( .A(n23833), .B(n23832), .Z(n23837) );
  NAND U25469 ( .A(n23835), .B(n23834), .Z(n23836) );
  NAND U25470 ( .A(n23837), .B(n23836), .Z(n23965) );
  XOR U25471 ( .A(n23966), .B(n23967), .Z(n23891) );
  NAND U25472 ( .A(n23839), .B(n23838), .Z(n23843) );
  NAND U25473 ( .A(n23841), .B(n23840), .Z(n23842) );
  AND U25474 ( .A(n23843), .B(n23842), .Z(n23892) );
  XOR U25475 ( .A(n23891), .B(n23892), .Z(n23893) );
  XOR U25476 ( .A(n23894), .B(n23893), .Z(n23877) );
  NAND U25477 ( .A(n23845), .B(n23844), .Z(n23849) );
  NAND U25478 ( .A(n23847), .B(n23846), .Z(n23848) );
  NAND U25479 ( .A(n23849), .B(n23848), .Z(n23888) );
  NAND U25480 ( .A(n23851), .B(n23850), .Z(n23855) );
  NAND U25481 ( .A(n23853), .B(n23852), .Z(n23854) );
  NAND U25482 ( .A(n23855), .B(n23854), .Z(n23886) );
  NAND U25483 ( .A(n23857), .B(n23856), .Z(n23861) );
  NAND U25484 ( .A(n23859), .B(n23858), .Z(n23860) );
  NAND U25485 ( .A(n23861), .B(n23860), .Z(n23885) );
  XOR U25486 ( .A(n23886), .B(n23885), .Z(n23887) );
  XOR U25487 ( .A(n23888), .B(n23887), .Z(n23876) );
  XNOR U25488 ( .A(n23879), .B(n23878), .Z(n23884) );
  NANDN U25489 ( .A(n23862), .B(n23863), .Z(n23868) );
  NOR U25490 ( .A(n23864), .B(n23863), .Z(n23866) );
  OR U25491 ( .A(n23866), .B(n23865), .Z(n23867) );
  AND U25492 ( .A(n23868), .B(n23867), .Z(n23882) );
  NAND U25493 ( .A(n23870), .B(n23869), .Z(n23874) );
  NAND U25494 ( .A(n23872), .B(n23871), .Z(n23873) );
  AND U25495 ( .A(n23874), .B(n23873), .Z(n23883) );
  XOR U25496 ( .A(n23882), .B(n23883), .Z(n23875) );
  XNOR U25497 ( .A(n23884), .B(n23875), .Z(N505) );
  NANDN U25498 ( .A(n23877), .B(n23876), .Z(n23881) );
  NAND U25499 ( .A(n23879), .B(n23878), .Z(n23880) );
  NAND U25500 ( .A(n23881), .B(n23880), .Z(n24025) );
  IV U25501 ( .A(n24025), .Z(n24024) );
  NAND U25502 ( .A(n23886), .B(n23885), .Z(n23890) );
  NAND U25503 ( .A(n23888), .B(n23887), .Z(n23889) );
  AND U25504 ( .A(n23890), .B(n23889), .Z(n24021) );
  NAND U25505 ( .A(n23892), .B(n23891), .Z(n23896) );
  NAND U25506 ( .A(n23894), .B(n23893), .Z(n23895) );
  NAND U25507 ( .A(n23896), .B(n23895), .Z(n24019) );
  NANDN U25508 ( .A(n23898), .B(n23897), .Z(n23902) );
  NANDN U25509 ( .A(n23900), .B(n23899), .Z(n23901) );
  NAND U25510 ( .A(n23902), .B(n23901), .Z(n24031) );
  IV U25511 ( .A(n23931), .Z(n24055) );
  NANDN U25512 ( .A(n24055), .B(n23903), .Z(n23907) );
  NAND U25513 ( .A(n23905), .B(n23904), .Z(n23906) );
  NAND U25514 ( .A(n23907), .B(n23906), .Z(n24079) );
  AND U25515 ( .A(x[494]), .B(y[7920]), .Z(n25000) );
  NAND U25516 ( .A(n25000), .B(n23908), .Z(n23912) );
  NANDN U25517 ( .A(n23910), .B(n23909), .Z(n23911) );
  AND U25518 ( .A(n23912), .B(n23911), .Z(n24108) );
  AND U25519 ( .A(x[491]), .B(y[7918]), .Z(n24127) );
  AND U25520 ( .A(x[492]), .B(y[7917]), .Z(n24125) );
  NAND U25521 ( .A(x[487]), .B(y[7922]), .Z(n24124) );
  NAND U25522 ( .A(x[504]), .B(y[7905]), .Z(n24123) );
  XNOR U25523 ( .A(o[249]), .B(n24123), .Z(n24093) );
  NAND U25524 ( .A(x[481]), .B(y[7928]), .Z(n24094) );
  NAND U25525 ( .A(x[493]), .B(y[7916]), .Z(n24096) );
  XOR U25526 ( .A(n24105), .B(n24106), .Z(n24107) );
  XOR U25527 ( .A(n24079), .B(n24080), .Z(n24082) );
  NAND U25528 ( .A(n23914), .B(n23913), .Z(n23918) );
  ANDN U25529 ( .B(n23916), .A(n23915), .Z(n23917) );
  ANDN U25530 ( .B(n23918), .A(n23917), .Z(n24068) );
  AND U25531 ( .A(n23920), .B(n23919), .Z(n23924) );
  NAND U25532 ( .A(n23922), .B(n23921), .Z(n23923) );
  NANDN U25533 ( .A(n23924), .B(n23923), .Z(n24067) );
  NANDN U25534 ( .A(n23926), .B(n23925), .Z(n23930) );
  NAND U25535 ( .A(n23928), .B(n23927), .Z(n23929) );
  AND U25536 ( .A(n23930), .B(n23929), .Z(n24064) );
  AND U25537 ( .A(x[488]), .B(y[7921]), .Z(n24058) );
  XNOR U25538 ( .A(n23932), .B(n23931), .Z(n24057) );
  ANDN U25539 ( .B(o[248]), .A(n23933), .Z(n24052) );
  AND U25540 ( .A(x[505]), .B(y[7904]), .Z(n24050) );
  NAND U25541 ( .A(x[480]), .B(y[7929]), .Z(n24049) );
  XOR U25542 ( .A(n24052), .B(n24051), .Z(n24061) );
  XOR U25543 ( .A(n24062), .B(n24061), .Z(n24063) );
  XOR U25544 ( .A(n24070), .B(n24069), .Z(n24081) );
  XOR U25545 ( .A(n24082), .B(n24081), .Z(n24162) );
  NAND U25546 ( .A(n23935), .B(n23934), .Z(n23939) );
  NAND U25547 ( .A(n23937), .B(n23936), .Z(n23938) );
  AND U25548 ( .A(n23939), .B(n23938), .Z(n24159) );
  NAND U25549 ( .A(n23941), .B(n23940), .Z(n23945) );
  ANDN U25550 ( .B(n23943), .A(n23942), .Z(n23944) );
  ANDN U25551 ( .B(n23945), .A(n23944), .Z(n24144) );
  NANDN U25552 ( .A(n23947), .B(n23946), .Z(n23951) );
  NAND U25553 ( .A(n23949), .B(n23948), .Z(n23950) );
  AND U25554 ( .A(n23951), .B(n23950), .Z(n24142) );
  AND U25555 ( .A(x[494]), .B(y[7915]), .Z(n24099) );
  NAND U25556 ( .A(x[482]), .B(y[7927]), .Z(n24100) );
  NAND U25557 ( .A(x[483]), .B(y[7926]), .Z(n24102) );
  NAND U25558 ( .A(n23953), .B(n23952), .Z(n23957) );
  NAND U25559 ( .A(n23955), .B(n23954), .Z(n23956) );
  AND U25560 ( .A(n23957), .B(n23956), .Z(n24165) );
  XOR U25561 ( .A(n24166), .B(n24165), .Z(n24168) );
  NANDN U25562 ( .A(n23959), .B(n23958), .Z(n23963) );
  NANDN U25563 ( .A(n23961), .B(n23960), .Z(n23962) );
  AND U25564 ( .A(n23963), .B(n23962), .Z(n24167) );
  XOR U25565 ( .A(n24168), .B(n24167), .Z(n24032) );
  XOR U25566 ( .A(n24031), .B(n24032), .Z(n24033) );
  NANDN U25567 ( .A(n23965), .B(n23964), .Z(n23969) );
  NAND U25568 ( .A(n23967), .B(n23966), .Z(n23968) );
  NAND U25569 ( .A(n23969), .B(n23968), .Z(n24039) );
  NAND U25570 ( .A(n23971), .B(n23970), .Z(n23975) );
  NANDN U25571 ( .A(n23973), .B(n23972), .Z(n23974) );
  NAND U25572 ( .A(n23975), .B(n23974), .Z(n24044) );
  NAND U25573 ( .A(n23977), .B(n23976), .Z(n23981) );
  NAND U25574 ( .A(n23979), .B(n23978), .Z(n23980) );
  NAND U25575 ( .A(n23981), .B(n23980), .Z(n24043) );
  XOR U25576 ( .A(n24044), .B(n24043), .Z(n24045) );
  NAND U25577 ( .A(x[501]), .B(y[7912]), .Z(n24870) );
  NANDN U25578 ( .A(n24870), .B(n23982), .Z(n23986) );
  NANDN U25579 ( .A(n23984), .B(n23983), .Z(n23985) );
  AND U25580 ( .A(n23986), .B(n23985), .Z(n24150) );
  AND U25581 ( .A(x[502]), .B(y[7907]), .Z(n24120) );
  AND U25582 ( .A(x[485]), .B(y[7924]), .Z(n24118) );
  NAND U25583 ( .A(x[497]), .B(y[7912]), .Z(n24117) );
  AND U25584 ( .A(y[7909]), .B(x[500]), .Z(n23988) );
  NAND U25585 ( .A(y[7908]), .B(x[501]), .Z(n23987) );
  XNOR U25586 ( .A(n23988), .B(n23987), .Z(n24131) );
  NAND U25587 ( .A(x[499]), .B(y[7910]), .Z(n24132) );
  XOR U25588 ( .A(n24147), .B(n24148), .Z(n24149) );
  NANDN U25589 ( .A(n24130), .B(n24227), .Z(n23992) );
  NAND U25590 ( .A(n23990), .B(n23989), .Z(n23991) );
  AND U25591 ( .A(n23992), .B(n23991), .Z(n24156) );
  AND U25592 ( .A(x[495]), .B(y[7914]), .Z(n24138) );
  AND U25593 ( .A(x[498]), .B(y[7911]), .Z(n24136) );
  NAND U25594 ( .A(x[486]), .B(y[7923]), .Z(n24135) );
  AND U25595 ( .A(x[503]), .B(y[7906]), .Z(n24114) );
  AND U25596 ( .A(x[484]), .B(y[7925]), .Z(n24112) );
  NAND U25597 ( .A(x[496]), .B(y[7913]), .Z(n24111) );
  XOR U25598 ( .A(n24114), .B(n24113), .Z(n24153) );
  XOR U25599 ( .A(n24154), .B(n24153), .Z(n24155) );
  XOR U25600 ( .A(n24156), .B(n24155), .Z(n24073) );
  NAND U25601 ( .A(n23994), .B(n23993), .Z(n23998) );
  NAND U25602 ( .A(n23996), .B(n23995), .Z(n23997) );
  AND U25603 ( .A(n23998), .B(n23997), .Z(n24075) );
  XNOR U25604 ( .A(n24076), .B(n24075), .Z(n24087) );
  NAND U25605 ( .A(n24000), .B(n23999), .Z(n24004) );
  NAND U25606 ( .A(n24002), .B(n24001), .Z(n24003) );
  NAND U25607 ( .A(n24004), .B(n24003), .Z(n24086) );
  NAND U25608 ( .A(n24006), .B(n24005), .Z(n24010) );
  NAND U25609 ( .A(n24008), .B(n24007), .Z(n24009) );
  NAND U25610 ( .A(n24010), .B(n24009), .Z(n24085) );
  XNOR U25611 ( .A(n24086), .B(n24085), .Z(n24088) );
  XNOR U25612 ( .A(n24045), .B(n24046), .Z(n24038) );
  NAND U25613 ( .A(n24012), .B(n24011), .Z(n24016) );
  NAND U25614 ( .A(n24014), .B(n24013), .Z(n24015) );
  NAND U25615 ( .A(n24016), .B(n24015), .Z(n24037) );
  XOR U25616 ( .A(n24039), .B(n24040), .Z(n24034) );
  XNOR U25617 ( .A(n24033), .B(n24034), .Z(n24018) );
  XOR U25618 ( .A(n24019), .B(n24018), .Z(n24020) );
  XOR U25619 ( .A(n24021), .B(n24020), .Z(n24027) );
  XNOR U25620 ( .A(n24026), .B(n24027), .Z(n24017) );
  XOR U25621 ( .A(n24024), .B(n24017), .Z(N506) );
  NAND U25622 ( .A(n24019), .B(n24018), .Z(n24023) );
  NAND U25623 ( .A(n24021), .B(n24020), .Z(n24022) );
  NAND U25624 ( .A(n24023), .B(n24022), .Z(n24180) );
  IV U25625 ( .A(n24180), .Z(n24178) );
  OR U25626 ( .A(n24026), .B(n24024), .Z(n24030) );
  ANDN U25627 ( .B(n24026), .A(n24025), .Z(n24028) );
  OR U25628 ( .A(n24028), .B(n24027), .Z(n24029) );
  AND U25629 ( .A(n24030), .B(n24029), .Z(n24179) );
  NAND U25630 ( .A(n24032), .B(n24031), .Z(n24036) );
  NANDN U25631 ( .A(n24034), .B(n24033), .Z(n24035) );
  AND U25632 ( .A(n24036), .B(n24035), .Z(n24173) );
  NANDN U25633 ( .A(n24038), .B(n24037), .Z(n24042) );
  NANDN U25634 ( .A(n24040), .B(n24039), .Z(n24041) );
  AND U25635 ( .A(n24042), .B(n24041), .Z(n24172) );
  XOR U25636 ( .A(n24173), .B(n24172), .Z(n24175) );
  NAND U25637 ( .A(n24044), .B(n24043), .Z(n24048) );
  NANDN U25638 ( .A(n24046), .B(n24045), .Z(n24047) );
  NAND U25639 ( .A(n24048), .B(n24047), .Z(n24329) );
  AND U25640 ( .A(x[482]), .B(y[7928]), .Z(n24259) );
  XOR U25641 ( .A(n24260), .B(n24259), .Z(n24262) );
  NAND U25642 ( .A(x[504]), .B(y[7906]), .Z(n24261) );
  XNOR U25643 ( .A(n24262), .B(n24261), .Z(n24295) );
  NANDN U25644 ( .A(n24050), .B(n24049), .Z(n24054) );
  NANDN U25645 ( .A(n24052), .B(n24051), .Z(n24053) );
  NAND U25646 ( .A(n24054), .B(n24053), .Z(n24296) );
  NANDN U25647 ( .A(n24056), .B(n24055), .Z(n24060) );
  NANDN U25648 ( .A(n24058), .B(n24057), .Z(n24059) );
  AND U25649 ( .A(n24060), .B(n24059), .Z(n24297) );
  XOR U25650 ( .A(n24298), .B(n24297), .Z(n24204) );
  NAND U25651 ( .A(n24062), .B(n24061), .Z(n24066) );
  NANDN U25652 ( .A(n24064), .B(n24063), .Z(n24065) );
  AND U25653 ( .A(n24066), .B(n24065), .Z(n24203) );
  NANDN U25654 ( .A(n24068), .B(n24067), .Z(n24072) );
  NAND U25655 ( .A(n24070), .B(n24069), .Z(n24071) );
  NAND U25656 ( .A(n24072), .B(n24071), .Z(n24206) );
  NANDN U25657 ( .A(n24074), .B(n24073), .Z(n24078) );
  NAND U25658 ( .A(n24076), .B(n24075), .Z(n24077) );
  NAND U25659 ( .A(n24078), .B(n24077), .Z(n24191) );
  NAND U25660 ( .A(n24080), .B(n24079), .Z(n24084) );
  NAND U25661 ( .A(n24082), .B(n24081), .Z(n24083) );
  AND U25662 ( .A(n24084), .B(n24083), .Z(n24192) );
  XNOR U25663 ( .A(n24191), .B(n24192), .Z(n24194) );
  NAND U25664 ( .A(n24086), .B(n24085), .Z(n24090) );
  NANDN U25665 ( .A(n24088), .B(n24087), .Z(n24089) );
  NAND U25666 ( .A(n24090), .B(n24089), .Z(n24243) );
  AND U25667 ( .A(y[7924]), .B(x[486]), .Z(n24092) );
  NAND U25668 ( .A(y[7922]), .B(x[488]), .Z(n24091) );
  XNOR U25669 ( .A(n24092), .B(n24091), .Z(n24228) );
  NAND U25670 ( .A(x[489]), .B(y[7921]), .Z(n24229) );
  XNOR U25671 ( .A(n24228), .B(n24229), .Z(n24210) );
  AND U25672 ( .A(x[487]), .B(y[7923]), .Z(n24209) );
  XOR U25673 ( .A(n24210), .B(n24209), .Z(n24212) );
  AND U25674 ( .A(x[492]), .B(y[7918]), .Z(n24428) );
  AND U25675 ( .A(x[485]), .B(y[7925]), .Z(n24310) );
  XOR U25676 ( .A(n24428), .B(n24310), .Z(n24312) );
  AND U25677 ( .A(x[490]), .B(y[7920]), .Z(n24311) );
  XOR U25678 ( .A(n24312), .B(n24311), .Z(n24211) );
  XOR U25679 ( .A(n24212), .B(n24211), .Z(n24286) );
  NANDN U25680 ( .A(n24094), .B(n24093), .Z(n24098) );
  NANDN U25681 ( .A(n24096), .B(n24095), .Z(n24097) );
  AND U25682 ( .A(n24098), .B(n24097), .Z(n24284) );
  NANDN U25683 ( .A(n24100), .B(n24099), .Z(n24104) );
  NANDN U25684 ( .A(n24102), .B(n24101), .Z(n24103) );
  NAND U25685 ( .A(n24104), .B(n24103), .Z(n24283) );
  XOR U25686 ( .A(n24286), .B(n24285), .Z(n24322) );
  NAND U25687 ( .A(n24106), .B(n24105), .Z(n24110) );
  NANDN U25688 ( .A(n24108), .B(n24107), .Z(n24109) );
  AND U25689 ( .A(n24110), .B(n24109), .Z(n24321) );
  NANDN U25690 ( .A(n24112), .B(n24111), .Z(n24116) );
  NANDN U25691 ( .A(n24114), .B(n24113), .Z(n24115) );
  AND U25692 ( .A(n24116), .B(n24115), .Z(n24247) );
  NANDN U25693 ( .A(n24118), .B(n24117), .Z(n24122) );
  NANDN U25694 ( .A(n24120), .B(n24119), .Z(n24121) );
  NAND U25695 ( .A(n24122), .B(n24121), .Z(n24248) );
  ANDN U25696 ( .B(o[249]), .A(n24123), .Z(n24221) );
  NAND U25697 ( .A(x[494]), .B(y[7916]), .Z(n24222) );
  XNOR U25698 ( .A(n24221), .B(n24222), .Z(n24223) );
  NAND U25699 ( .A(x[481]), .B(y[7929]), .Z(n24224) );
  XNOR U25700 ( .A(n24223), .B(n24224), .Z(n24301) );
  NAND U25701 ( .A(x[505]), .B(y[7905]), .Z(n24232) );
  XNOR U25702 ( .A(o[250]), .B(n24232), .Z(n24315) );
  NAND U25703 ( .A(x[506]), .B(y[7904]), .Z(n24316) );
  XNOR U25704 ( .A(n24315), .B(n24316), .Z(n24317) );
  NAND U25705 ( .A(x[480]), .B(y[7930]), .Z(n24318) );
  XOR U25706 ( .A(n24317), .B(n24318), .Z(n24302) );
  NANDN U25707 ( .A(n24125), .B(n24124), .Z(n24129) );
  NANDN U25708 ( .A(n24127), .B(n24126), .Z(n24128) );
  NAND U25709 ( .A(n24129), .B(n24128), .Z(n24304) );
  XOR U25710 ( .A(n24250), .B(n24249), .Z(n24292) );
  AND U25711 ( .A(x[501]), .B(y[7909]), .Z(n24215) );
  NANDN U25712 ( .A(n24130), .B(n24215), .Z(n24134) );
  NANDN U25713 ( .A(n24132), .B(n24131), .Z(n24133) );
  AND U25714 ( .A(n24134), .B(n24133), .Z(n24280) );
  XOR U25715 ( .A(n24216), .B(n24215), .Z(n24218) );
  NAND U25716 ( .A(x[500]), .B(y[7910]), .Z(n24217) );
  XNOR U25717 ( .A(n24218), .B(n24217), .Z(n24277) );
  NAND U25718 ( .A(x[503]), .B(y[7907]), .Z(n24266) );
  XNOR U25719 ( .A(n24265), .B(n24266), .Z(n24267) );
  NAND U25720 ( .A(x[502]), .B(y[7908]), .Z(n24268) );
  XOR U25721 ( .A(n24267), .B(n24268), .Z(n24278) );
  AND U25722 ( .A(x[484]), .B(y[7926]), .Z(n24271) );
  XOR U25723 ( .A(n24272), .B(n24271), .Z(n24274) );
  XNOR U25724 ( .A(n24274), .B(n24273), .Z(n24253) );
  AND U25725 ( .A(x[491]), .B(y[7919]), .Z(n24233) );
  NAND U25726 ( .A(x[499]), .B(y[7911]), .Z(n24234) );
  XNOR U25727 ( .A(n24233), .B(n24234), .Z(n24235) );
  NAND U25728 ( .A(x[483]), .B(y[7927]), .Z(n24236) );
  XOR U25729 ( .A(n24235), .B(n24236), .Z(n24254) );
  NANDN U25730 ( .A(n24136), .B(n24135), .Z(n24140) );
  NANDN U25731 ( .A(n24138), .B(n24137), .Z(n24139) );
  AND U25732 ( .A(n24140), .B(n24139), .Z(n24255) );
  XNOR U25733 ( .A(n24256), .B(n24255), .Z(n24289) );
  XOR U25734 ( .A(n24290), .B(n24289), .Z(n24291) );
  XOR U25735 ( .A(n24324), .B(n24323), .Z(n24242) );
  NANDN U25736 ( .A(n24142), .B(n24141), .Z(n24146) );
  NANDN U25737 ( .A(n24144), .B(n24143), .Z(n24145) );
  AND U25738 ( .A(n24146), .B(n24145), .Z(n24200) );
  NAND U25739 ( .A(n24148), .B(n24147), .Z(n24152) );
  NANDN U25740 ( .A(n24150), .B(n24149), .Z(n24151) );
  AND U25741 ( .A(n24152), .B(n24151), .Z(n24198) );
  NAND U25742 ( .A(n24154), .B(n24153), .Z(n24158) );
  NANDN U25743 ( .A(n24156), .B(n24155), .Z(n24157) );
  NAND U25744 ( .A(n24158), .B(n24157), .Z(n24197) );
  XOR U25745 ( .A(n24243), .B(n24244), .Z(n24327) );
  XOR U25746 ( .A(n24329), .B(n24330), .Z(n24188) );
  NANDN U25747 ( .A(n24160), .B(n24159), .Z(n24164) );
  NANDN U25748 ( .A(n24162), .B(n24161), .Z(n24163) );
  AND U25749 ( .A(n24164), .B(n24163), .Z(n24186) );
  NAND U25750 ( .A(n24166), .B(n24165), .Z(n24170) );
  NAND U25751 ( .A(n24168), .B(n24167), .Z(n24169) );
  AND U25752 ( .A(n24170), .B(n24169), .Z(n24185) );
  XOR U25753 ( .A(n24186), .B(n24185), .Z(n24187) );
  XOR U25754 ( .A(n24188), .B(n24187), .Z(n24174) );
  XOR U25755 ( .A(n24175), .B(n24174), .Z(n24181) );
  XNOR U25756 ( .A(n24179), .B(n24181), .Z(n24171) );
  XOR U25757 ( .A(n24178), .B(n24171), .Z(N507) );
  NAND U25758 ( .A(n24173), .B(n24172), .Z(n24177) );
  NAND U25759 ( .A(n24175), .B(n24174), .Z(n24176) );
  AND U25760 ( .A(n24177), .B(n24176), .Z(n24340) );
  NANDN U25761 ( .A(n24178), .B(n24179), .Z(n24184) );
  NOR U25762 ( .A(n24180), .B(n24179), .Z(n24182) );
  OR U25763 ( .A(n24182), .B(n24181), .Z(n24183) );
  AND U25764 ( .A(n24184), .B(n24183), .Z(n24341) );
  NAND U25765 ( .A(n24186), .B(n24185), .Z(n24190) );
  NAND U25766 ( .A(n24188), .B(n24187), .Z(n24189) );
  NAND U25767 ( .A(n24190), .B(n24189), .Z(n24336) );
  NAND U25768 ( .A(n24192), .B(n24191), .Z(n24196) );
  NANDN U25769 ( .A(n24194), .B(n24193), .Z(n24195) );
  NAND U25770 ( .A(n24196), .B(n24195), .Z(n24350) );
  NANDN U25771 ( .A(n24198), .B(n24197), .Z(n24202) );
  NANDN U25772 ( .A(n24200), .B(n24199), .Z(n24201) );
  AND U25773 ( .A(n24202), .B(n24201), .Z(n24358) );
  NANDN U25774 ( .A(n24204), .B(n24203), .Z(n24208) );
  NANDN U25775 ( .A(n24206), .B(n24205), .Z(n24207) );
  AND U25776 ( .A(n24208), .B(n24207), .Z(n24356) );
  NAND U25777 ( .A(n24210), .B(n24209), .Z(n24214) );
  NAND U25778 ( .A(n24212), .B(n24211), .Z(n24213) );
  AND U25779 ( .A(n24214), .B(n24213), .Z(n24479) );
  NAND U25780 ( .A(n24216), .B(n24215), .Z(n24220) );
  ANDN U25781 ( .B(n24218), .A(n24217), .Z(n24219) );
  ANDN U25782 ( .B(n24220), .A(n24219), .Z(n24442) );
  NANDN U25783 ( .A(n24222), .B(n24221), .Z(n24226) );
  NANDN U25784 ( .A(n24224), .B(n24223), .Z(n24225) );
  NAND U25785 ( .A(n24226), .B(n24225), .Z(n24441) );
  XNOR U25786 ( .A(n24442), .B(n24441), .Z(n24443) );
  AND U25787 ( .A(x[488]), .B(y[7924]), .Z(n24391) );
  NAND U25788 ( .A(n24391), .B(n24227), .Z(n24231) );
  NANDN U25789 ( .A(n24229), .B(n24228), .Z(n24230) );
  AND U25790 ( .A(n24231), .B(n24230), .Z(n24407) );
  AND U25791 ( .A(x[494]), .B(y[7917]), .Z(n24437) );
  NAND U25792 ( .A(x[481]), .B(y[7930]), .Z(n24438) );
  XNOR U25793 ( .A(n24437), .B(n24438), .Z(n24440) );
  ANDN U25794 ( .B(o[250]), .A(n24232), .Z(n24439) );
  XOR U25795 ( .A(n24440), .B(n24439), .Z(n24404) );
  AND U25796 ( .A(x[497]), .B(y[7914]), .Z(n24373) );
  NAND U25797 ( .A(x[484]), .B(y[7927]), .Z(n24374) );
  XNOR U25798 ( .A(n24373), .B(n24374), .Z(n24375) );
  NAND U25799 ( .A(x[485]), .B(y[7926]), .Z(n24376) );
  XOR U25800 ( .A(n24375), .B(n24376), .Z(n24405) );
  XNOR U25801 ( .A(n24404), .B(n24405), .Z(n24406) );
  XOR U25802 ( .A(n24407), .B(n24406), .Z(n24444) );
  XNOR U25803 ( .A(n24443), .B(n24444), .Z(n24476) );
  NANDN U25804 ( .A(n24234), .B(n24233), .Z(n24238) );
  NANDN U25805 ( .A(n24236), .B(n24235), .Z(n24237) );
  AND U25806 ( .A(n24238), .B(n24237), .Z(n24450) );
  AND U25807 ( .A(y[7907]), .B(x[504]), .Z(n24240) );
  NAND U25808 ( .A(y[7911]), .B(x[500]), .Z(n24239) );
  XNOR U25809 ( .A(n24240), .B(n24239), .Z(n24362) );
  NAND U25810 ( .A(x[487]), .B(y[7924]), .Z(n24363) );
  XNOR U25811 ( .A(n24362), .B(n24363), .Z(n24447) );
  AND U25812 ( .A(x[488]), .B(y[7923]), .Z(n24422) );
  NAND U25813 ( .A(x[503]), .B(y[7908]), .Z(n24423) );
  XNOR U25814 ( .A(n24422), .B(n24423), .Z(n24424) );
  NAND U25815 ( .A(x[502]), .B(y[7909]), .Z(n24425) );
  XOR U25816 ( .A(n24424), .B(n24425), .Z(n24448) );
  XNOR U25817 ( .A(n24447), .B(n24448), .Z(n24449) );
  XOR U25818 ( .A(n24450), .B(n24449), .Z(n24477) );
  XOR U25819 ( .A(n24356), .B(n24355), .Z(n24357) );
  XOR U25820 ( .A(n24358), .B(n24357), .Z(n24349) );
  XOR U25821 ( .A(n24350), .B(n24349), .Z(n24352) );
  NANDN U25822 ( .A(n24242), .B(n24241), .Z(n24246) );
  NAND U25823 ( .A(n24244), .B(n24243), .Z(n24245) );
  AND U25824 ( .A(n24246), .B(n24245), .Z(n24346) );
  NANDN U25825 ( .A(n24248), .B(n24247), .Z(n24252) );
  NAND U25826 ( .A(n24250), .B(n24249), .Z(n24251) );
  AND U25827 ( .A(n24252), .B(n24251), .Z(n24467) );
  NANDN U25828 ( .A(n24254), .B(n24253), .Z(n24258) );
  NAND U25829 ( .A(n24256), .B(n24255), .Z(n24257) );
  AND U25830 ( .A(n24258), .B(n24257), .Z(n24465) );
  NAND U25831 ( .A(n24260), .B(n24259), .Z(n24264) );
  ANDN U25832 ( .B(n24262), .A(n24261), .Z(n24263) );
  ANDN U25833 ( .B(n24264), .A(n24263), .Z(n24399) );
  NANDN U25834 ( .A(n24266), .B(n24265), .Z(n24270) );
  NANDN U25835 ( .A(n24268), .B(n24267), .Z(n24269) );
  NAND U25836 ( .A(n24270), .B(n24269), .Z(n24398) );
  XNOR U25837 ( .A(n24399), .B(n24398), .Z(n24400) );
  NAND U25838 ( .A(n24272), .B(n24271), .Z(n24276) );
  ANDN U25839 ( .B(n24274), .A(n24273), .Z(n24275) );
  ANDN U25840 ( .B(n24276), .A(n24275), .Z(n24413) );
  AND U25841 ( .A(x[480]), .B(y[7931]), .Z(n24379) );
  NAND U25842 ( .A(x[507]), .B(y[7904]), .Z(n24380) );
  XNOR U25843 ( .A(n24379), .B(n24380), .Z(n24382) );
  AND U25844 ( .A(x[506]), .B(y[7905]), .Z(n24389) );
  XOR U25845 ( .A(o[251]), .B(n24389), .Z(n24381) );
  XOR U25846 ( .A(n24382), .B(n24381), .Z(n24410) );
  AND U25847 ( .A(x[489]), .B(y[7922]), .Z(n24383) );
  NAND U25848 ( .A(x[501]), .B(y[7910]), .Z(n24384) );
  XNOR U25849 ( .A(n24383), .B(n24384), .Z(n24385) );
  NAND U25850 ( .A(x[498]), .B(y[7913]), .Z(n24386) );
  XOR U25851 ( .A(n24385), .B(n24386), .Z(n24411) );
  XNOR U25852 ( .A(n24410), .B(n24411), .Z(n24412) );
  XOR U25853 ( .A(n24413), .B(n24412), .Z(n24401) );
  XNOR U25854 ( .A(n24400), .B(n24401), .Z(n24464) );
  NANDN U25855 ( .A(n24278), .B(n24277), .Z(n24282) );
  NANDN U25856 ( .A(n24280), .B(n24279), .Z(n24281) );
  AND U25857 ( .A(n24282), .B(n24281), .Z(n24482) );
  NANDN U25858 ( .A(n24284), .B(n24283), .Z(n24288) );
  NAND U25859 ( .A(n24286), .B(n24285), .Z(n24287) );
  NAND U25860 ( .A(n24288), .B(n24287), .Z(n24483) );
  XOR U25861 ( .A(n24484), .B(n24485), .Z(n24343) );
  NAND U25862 ( .A(n24290), .B(n24289), .Z(n24294) );
  NANDN U25863 ( .A(n24292), .B(n24291), .Z(n24293) );
  AND U25864 ( .A(n24294), .B(n24293), .Z(n24471) );
  NANDN U25865 ( .A(n24296), .B(n24295), .Z(n24300) );
  NAND U25866 ( .A(n24298), .B(n24297), .Z(n24299) );
  AND U25867 ( .A(n24300), .B(n24299), .Z(n24461) );
  NANDN U25868 ( .A(n24302), .B(n24301), .Z(n24306) );
  NANDN U25869 ( .A(n24304), .B(n24303), .Z(n24305) );
  AND U25870 ( .A(n24306), .B(n24305), .Z(n24459) );
  AND U25871 ( .A(x[499]), .B(y[7912]), .Z(n24366) );
  NAND U25872 ( .A(x[505]), .B(y[7906]), .Z(n24367) );
  XNOR U25873 ( .A(n24366), .B(n24367), .Z(n24368) );
  NAND U25874 ( .A(x[486]), .B(y[7925]), .Z(n24369) );
  XNOR U25875 ( .A(n24368), .B(n24369), .Z(n24453) );
  AND U25876 ( .A(x[495]), .B(y[7916]), .Z(n24431) );
  NAND U25877 ( .A(x[482]), .B(y[7929]), .Z(n24432) );
  XNOR U25878 ( .A(n24431), .B(n24432), .Z(n24433) );
  NAND U25879 ( .A(x[483]), .B(y[7928]), .Z(n24434) );
  XOR U25880 ( .A(n24433), .B(n24434), .Z(n24454) );
  XNOR U25881 ( .A(n24453), .B(n24454), .Z(n24456) );
  AND U25882 ( .A(x[496]), .B(y[7915]), .Z(n24417) );
  XOR U25883 ( .A(n24417), .B(n24307), .Z(n24418) );
  XOR U25884 ( .A(n24419), .B(n24418), .Z(n24429) );
  AND U25885 ( .A(y[7918]), .B(x[493]), .Z(n24309) );
  NAND U25886 ( .A(y[7919]), .B(x[492]), .Z(n24308) );
  XNOR U25887 ( .A(n24309), .B(n24308), .Z(n24430) );
  XOR U25888 ( .A(n24429), .B(n24430), .Z(n24455) );
  XOR U25889 ( .A(n24456), .B(n24455), .Z(n24394) );
  NAND U25890 ( .A(n24428), .B(n24310), .Z(n24314) );
  AND U25891 ( .A(n24312), .B(n24311), .Z(n24313) );
  ANDN U25892 ( .B(n24314), .A(n24313), .Z(n24393) );
  NANDN U25893 ( .A(n24316), .B(n24315), .Z(n24320) );
  NANDN U25894 ( .A(n24318), .B(n24317), .Z(n24319) );
  NAND U25895 ( .A(n24320), .B(n24319), .Z(n24392) );
  XOR U25896 ( .A(n24393), .B(n24392), .Z(n24395) );
  XNOR U25897 ( .A(n24394), .B(n24395), .Z(n24458) );
  XOR U25898 ( .A(n24471), .B(n24470), .Z(n24472) );
  NANDN U25899 ( .A(n24322), .B(n24321), .Z(n24326) );
  NAND U25900 ( .A(n24324), .B(n24323), .Z(n24325) );
  NAND U25901 ( .A(n24326), .B(n24325), .Z(n24473) );
  XOR U25902 ( .A(n24346), .B(n24345), .Z(n24351) );
  XOR U25903 ( .A(n24352), .B(n24351), .Z(n24335) );
  NANDN U25904 ( .A(n24328), .B(n24327), .Z(n24332) );
  NAND U25905 ( .A(n24330), .B(n24329), .Z(n24331) );
  NAND U25906 ( .A(n24332), .B(n24331), .Z(n24334) );
  XOR U25907 ( .A(n24336), .B(n24337), .Z(n24342) );
  XNOR U25908 ( .A(n24341), .B(n24342), .Z(n24333) );
  XOR U25909 ( .A(n24340), .B(n24333), .Z(N508) );
  NANDN U25910 ( .A(n24335), .B(n24334), .Z(n24339) );
  NAND U25911 ( .A(n24337), .B(n24336), .Z(n24338) );
  AND U25912 ( .A(n24339), .B(n24338), .Z(n24634) );
  NANDN U25913 ( .A(n24344), .B(n24343), .Z(n24348) );
  NAND U25914 ( .A(n24346), .B(n24345), .Z(n24347) );
  AND U25915 ( .A(n24348), .B(n24347), .Z(n24638) );
  NAND U25916 ( .A(n24350), .B(n24349), .Z(n24354) );
  NAND U25917 ( .A(n24352), .B(n24351), .Z(n24353) );
  AND U25918 ( .A(n24354), .B(n24353), .Z(n24637) );
  XOR U25919 ( .A(n24638), .B(n24637), .Z(n24640) );
  NAND U25920 ( .A(n24356), .B(n24355), .Z(n24360) );
  NANDN U25921 ( .A(n24358), .B(n24357), .Z(n24359) );
  AND U25922 ( .A(n24360), .B(n24359), .Z(n24490) );
  AND U25923 ( .A(x[504]), .B(y[7911]), .Z(n24882) );
  AND U25924 ( .A(x[500]), .B(y[7907]), .Z(n24361) );
  NAND U25925 ( .A(n24882), .B(n24361), .Z(n24365) );
  NANDN U25926 ( .A(n24363), .B(n24362), .Z(n24364) );
  AND U25927 ( .A(n24365), .B(n24364), .Z(n24633) );
  AND U25928 ( .A(x[505]), .B(y[7907]), .Z(n24551) );
  XOR U25929 ( .A(n24552), .B(n24551), .Z(n24550) );
  NAND U25930 ( .A(x[481]), .B(y[7931]), .Z(n24549) );
  AND U25931 ( .A(x[496]), .B(y[7916]), .Z(n24543) );
  NAND U25932 ( .A(x[504]), .B(y[7908]), .Z(n24544) );
  NAND U25933 ( .A(x[482]), .B(y[7930]), .Z(n24546) );
  XOR U25934 ( .A(n24631), .B(n24630), .Z(n24632) );
  XOR U25935 ( .A(n24633), .B(n24632), .Z(n24609) );
  NANDN U25936 ( .A(n24367), .B(n24366), .Z(n24371) );
  NANDN U25937 ( .A(n24369), .B(n24368), .Z(n24370) );
  AND U25938 ( .A(n24371), .B(n24370), .Z(n24629) );
  NAND U25939 ( .A(x[483]), .B(y[7929]), .Z(n24580) );
  NAND U25940 ( .A(x[503]), .B(y[7909]), .Z(n24582) );
  IV U25941 ( .A(n24582), .Z(n24372) );
  XOR U25942 ( .A(n24581), .B(n24372), .Z(n24627) );
  AND U25943 ( .A(x[485]), .B(y[7927]), .Z(n24566) );
  NAND U25944 ( .A(x[501]), .B(y[7911]), .Z(n24567) );
  NAND U25945 ( .A(x[500]), .B(y[7912]), .Z(n24569) );
  XOR U25946 ( .A(n24627), .B(n24626), .Z(n24628) );
  XOR U25947 ( .A(n24629), .B(n24628), .Z(n24606) );
  NANDN U25948 ( .A(n24374), .B(n24373), .Z(n24378) );
  NANDN U25949 ( .A(n24376), .B(n24375), .Z(n24377) );
  AND U25950 ( .A(n24378), .B(n24377), .Z(n24621) );
  XNOR U25951 ( .A(n24621), .B(n24620), .Z(n24623) );
  NANDN U25952 ( .A(n24384), .B(n24383), .Z(n24388) );
  NANDN U25953 ( .A(n24386), .B(n24385), .Z(n24387) );
  NAND U25954 ( .A(n24388), .B(n24387), .Z(n24516) );
  AND U25955 ( .A(n24389), .B(o[251]), .Z(n24529) );
  AND U25956 ( .A(x[480]), .B(y[7932]), .Z(n24527) );
  AND U25957 ( .A(x[508]), .B(y[7904]), .Z(n24526) );
  XOR U25958 ( .A(n24527), .B(n24526), .Z(n24528) );
  XOR U25959 ( .A(n24529), .B(n24528), .Z(n24515) );
  NAND U25960 ( .A(y[7922]), .B(x[490]), .Z(n24390) );
  XNOR U25961 ( .A(n24391), .B(n24390), .Z(n24534) );
  AND U25962 ( .A(x[489]), .B(y[7923]), .Z(n24533) );
  XOR U25963 ( .A(n24534), .B(n24533), .Z(n24514) );
  XOR U25964 ( .A(n24515), .B(n24514), .Z(n24517) );
  XOR U25965 ( .A(n24516), .B(n24517), .Z(n24622) );
  XNOR U25966 ( .A(n24623), .B(n24622), .Z(n24607) );
  XOR U25967 ( .A(n24606), .B(n24607), .Z(n24608) );
  XNOR U25968 ( .A(n24609), .B(n24608), .Z(n24508) );
  NANDN U25969 ( .A(n24393), .B(n24392), .Z(n24397) );
  NANDN U25970 ( .A(n24395), .B(n24394), .Z(n24396) );
  AND U25971 ( .A(n24397), .B(n24396), .Z(n24511) );
  NANDN U25972 ( .A(n24399), .B(n24398), .Z(n24403) );
  NANDN U25973 ( .A(n24401), .B(n24400), .Z(n24402) );
  AND U25974 ( .A(n24403), .B(n24402), .Z(n24613) );
  NANDN U25975 ( .A(n24405), .B(n24404), .Z(n24409) );
  NANDN U25976 ( .A(n24407), .B(n24406), .Z(n24408) );
  AND U25977 ( .A(n24409), .B(n24408), .Z(n24611) );
  NANDN U25978 ( .A(n24411), .B(n24410), .Z(n24415) );
  NANDN U25979 ( .A(n24413), .B(n24412), .Z(n24414) );
  NAND U25980 ( .A(n24415), .B(n24414), .Z(n24610) );
  XNOR U25981 ( .A(n24611), .B(n24610), .Z(n24612) );
  XNOR U25982 ( .A(n24613), .B(n24612), .Z(n24510) );
  XNOR U25983 ( .A(n24511), .B(n24510), .Z(n24513) );
  NANDN U25984 ( .A(n24417), .B(n24416), .Z(n24421) );
  NANDN U25985 ( .A(n24419), .B(n24418), .Z(n24420) );
  AND U25986 ( .A(n24421), .B(n24420), .Z(n24576) );
  AND U25987 ( .A(x[487]), .B(y[7925]), .Z(n24556) );
  AND U25988 ( .A(x[492]), .B(y[7920]), .Z(n24555) );
  XOR U25989 ( .A(n24556), .B(n24555), .Z(n24558) );
  AND U25990 ( .A(x[491]), .B(y[7921]), .Z(n24557) );
  XOR U25991 ( .A(n24558), .B(n24557), .Z(n24574) );
  AND U25992 ( .A(x[507]), .B(y[7905]), .Z(n24572) );
  XOR U25993 ( .A(o[252]), .B(n24572), .Z(n24586) );
  AND U25994 ( .A(x[506]), .B(y[7906]), .Z(n24585) );
  XOR U25995 ( .A(n24586), .B(n24585), .Z(n24588) );
  AND U25996 ( .A(x[495]), .B(y[7917]), .Z(n24587) );
  XNOR U25997 ( .A(n24588), .B(n24587), .Z(n24573) );
  NANDN U25998 ( .A(n24423), .B(n24422), .Z(n24427) );
  NANDN U25999 ( .A(n24425), .B(n24424), .Z(n24426) );
  AND U26000 ( .A(n24427), .B(n24426), .Z(n24597) );
  AND U26001 ( .A(x[497]), .B(y[7915]), .Z(n24521) );
  AND U26002 ( .A(x[502]), .B(y[7910]), .Z(n24520) );
  XOR U26003 ( .A(n24521), .B(n24520), .Z(n24523) );
  AND U26004 ( .A(x[484]), .B(y[7928]), .Z(n24522) );
  XOR U26005 ( .A(n24523), .B(n24522), .Z(n24595) );
  AND U26006 ( .A(x[486]), .B(y[7926]), .Z(n24743) );
  NAND U26007 ( .A(x[499]), .B(y[7913]), .Z(n24561) );
  XOR U26008 ( .A(n24595), .B(n24594), .Z(n24596) );
  XOR U26009 ( .A(n24617), .B(n24616), .Z(n24619) );
  NANDN U26010 ( .A(n24432), .B(n24431), .Z(n24436) );
  NANDN U26011 ( .A(n24434), .B(n24433), .Z(n24435) );
  AND U26012 ( .A(n24436), .B(n24435), .Z(n24538) );
  XOR U26013 ( .A(n24619), .B(n24618), .Z(n24512) );
  XOR U26014 ( .A(n24513), .B(n24512), .Z(n24509) );
  NANDN U26015 ( .A(n24442), .B(n24441), .Z(n24446) );
  NANDN U26016 ( .A(n24444), .B(n24443), .Z(n24445) );
  AND U26017 ( .A(n24446), .B(n24445), .Z(n24603) );
  NANDN U26018 ( .A(n24448), .B(n24447), .Z(n24452) );
  NANDN U26019 ( .A(n24450), .B(n24449), .Z(n24451) );
  AND U26020 ( .A(n24452), .B(n24451), .Z(n24601) );
  XNOR U26021 ( .A(n24601), .B(n24600), .Z(n24602) );
  XOR U26022 ( .A(n24603), .B(n24602), .Z(n24507) );
  XOR U26023 ( .A(n24509), .B(n24507), .Z(n24457) );
  XNOR U26024 ( .A(n24508), .B(n24457), .Z(n24504) );
  NANDN U26025 ( .A(n24459), .B(n24458), .Z(n24463) );
  NANDN U26026 ( .A(n24461), .B(n24460), .Z(n24462) );
  AND U26027 ( .A(n24463), .B(n24462), .Z(n24502) );
  NANDN U26028 ( .A(n24465), .B(n24464), .Z(n24469) );
  NANDN U26029 ( .A(n24467), .B(n24466), .Z(n24468) );
  NAND U26030 ( .A(n24469), .B(n24468), .Z(n24501) );
  XOR U26031 ( .A(n24504), .B(n24503), .Z(n24489) );
  NAND U26032 ( .A(n24471), .B(n24470), .Z(n24475) );
  NANDN U26033 ( .A(n24473), .B(n24472), .Z(n24474) );
  AND U26034 ( .A(n24475), .B(n24474), .Z(n24498) );
  NANDN U26035 ( .A(n24477), .B(n24476), .Z(n24481) );
  NANDN U26036 ( .A(n24479), .B(n24478), .Z(n24480) );
  AND U26037 ( .A(n24481), .B(n24480), .Z(n24496) );
  NANDN U26038 ( .A(n24483), .B(n24482), .Z(n24487) );
  NAND U26039 ( .A(n24485), .B(n24484), .Z(n24486) );
  AND U26040 ( .A(n24487), .B(n24486), .Z(n24495) );
  XOR U26041 ( .A(n24492), .B(n24491), .Z(n24639) );
  XOR U26042 ( .A(n24640), .B(n24639), .Z(n24636) );
  XNOR U26043 ( .A(n24635), .B(n24636), .Z(n24488) );
  XOR U26044 ( .A(n24634), .B(n24488), .Z(N509) );
  NANDN U26045 ( .A(n24490), .B(n24489), .Z(n24494) );
  NAND U26046 ( .A(n24492), .B(n24491), .Z(n24493) );
  AND U26047 ( .A(n24494), .B(n24493), .Z(n24650) );
  NANDN U26048 ( .A(n24496), .B(n24495), .Z(n24500) );
  NANDN U26049 ( .A(n24498), .B(n24497), .Z(n24499) );
  AND U26050 ( .A(n24500), .B(n24499), .Z(n24648) );
  NANDN U26051 ( .A(n24502), .B(n24501), .Z(n24506) );
  NAND U26052 ( .A(n24504), .B(n24503), .Z(n24505) );
  AND U26053 ( .A(n24506), .B(n24505), .Z(n24654) );
  NAND U26054 ( .A(n24515), .B(n24514), .Z(n24519) );
  NAND U26055 ( .A(n24517), .B(n24516), .Z(n24518) );
  AND U26056 ( .A(n24519), .B(n24518), .Z(n24774) );
  NAND U26057 ( .A(n24521), .B(n24520), .Z(n24525) );
  NAND U26058 ( .A(n24523), .B(n24522), .Z(n24524) );
  NAND U26059 ( .A(n24525), .B(n24524), .Z(n24811) );
  NAND U26060 ( .A(n24527), .B(n24526), .Z(n24531) );
  NAND U26061 ( .A(n24529), .B(n24528), .Z(n24530) );
  NAND U26062 ( .A(n24531), .B(n24530), .Z(n24810) );
  XOR U26063 ( .A(n24811), .B(n24810), .Z(n24812) );
  AND U26064 ( .A(y[7924]), .B(x[490]), .Z(n24808) );
  NAND U26065 ( .A(n24808), .B(n24532), .Z(n24536) );
  NAND U26066 ( .A(n24534), .B(n24533), .Z(n24535) );
  NAND U26067 ( .A(n24536), .B(n24535), .Z(n24782) );
  AND U26068 ( .A(x[502]), .B(y[7911]), .Z(n24721) );
  AND U26069 ( .A(x[492]), .B(y[7921]), .Z(n24865) );
  AND U26070 ( .A(x[481]), .B(y[7932]), .Z(n24719) );
  XOR U26071 ( .A(n24865), .B(n24719), .Z(n24720) );
  XOR U26072 ( .A(n24721), .B(n24720), .Z(n24781) );
  AND U26073 ( .A(x[495]), .B(y[7918]), .Z(n24724) );
  XOR U26074 ( .A(n24781), .B(n24780), .Z(n24783) );
  XNOR U26075 ( .A(n24782), .B(n24783), .Z(n24813) );
  NANDN U26076 ( .A(n24538), .B(n24537), .Z(n24542) );
  NANDN U26077 ( .A(n24540), .B(n24539), .Z(n24541) );
  AND U26078 ( .A(n24542), .B(n24541), .Z(n24776) );
  XOR U26079 ( .A(n24777), .B(n24776), .Z(n24771) );
  NANDN U26080 ( .A(n24544), .B(n24543), .Z(n24548) );
  NANDN U26081 ( .A(n24546), .B(n24545), .Z(n24547) );
  NAND U26082 ( .A(n24548), .B(n24547), .Z(n24787) );
  ANDN U26083 ( .B(n24550), .A(n24549), .Z(n24554) );
  NAND U26084 ( .A(n24552), .B(n24551), .Z(n24553) );
  NANDN U26085 ( .A(n24554), .B(n24553), .Z(n24786) );
  XOR U26086 ( .A(n24787), .B(n24786), .Z(n24788) );
  NAND U26087 ( .A(n24556), .B(n24555), .Z(n24560) );
  NAND U26088 ( .A(n24558), .B(n24557), .Z(n24559) );
  NAND U26089 ( .A(n24560), .B(n24559), .Z(n24685) );
  AND U26090 ( .A(x[491]), .B(y[7922]), .Z(n24740) );
  AND U26091 ( .A(x[483]), .B(y[7930]), .Z(n24738) );
  AND U26092 ( .A(x[497]), .B(y[7916]), .Z(n24737) );
  XOR U26093 ( .A(n24738), .B(n24737), .Z(n24739) );
  XOR U26094 ( .A(n24740), .B(n24739), .Z(n24684) );
  AND U26095 ( .A(x[503]), .B(y[7910]), .Z(n24734) );
  AND U26096 ( .A(x[493]), .B(y[7920]), .Z(n24732) );
  AND U26097 ( .A(x[504]), .B(y[7909]), .Z(n24934) );
  XOR U26098 ( .A(n24732), .B(n24934), .Z(n24733) );
  XOR U26099 ( .A(n24734), .B(n24733), .Z(n24683) );
  XOR U26100 ( .A(n24684), .B(n24683), .Z(n24686) );
  XNOR U26101 ( .A(n24685), .B(n24686), .Z(n24789) );
  NANDN U26102 ( .A(n24561), .B(n24743), .Z(n24565) );
  NANDN U26103 ( .A(n24563), .B(n24562), .Z(n24564) );
  NAND U26104 ( .A(n24565), .B(n24564), .Z(n24795) );
  AND U26105 ( .A(x[508]), .B(y[7905]), .Z(n24731) );
  XOR U26106 ( .A(o[253]), .B(n24731), .Z(n24803) );
  AND U26107 ( .A(x[480]), .B(y[7933]), .Z(n24801) );
  AND U26108 ( .A(x[509]), .B(y[7904]), .Z(n24800) );
  XOR U26109 ( .A(n24801), .B(n24800), .Z(n24802) );
  XOR U26110 ( .A(n24803), .B(n24802), .Z(n24793) );
  AND U26111 ( .A(x[505]), .B(y[7908]), .Z(n24716) );
  AND U26112 ( .A(x[506]), .B(y[7907]), .Z(n24713) );
  XOR U26113 ( .A(n24714), .B(n24713), .Z(n24715) );
  XOR U26114 ( .A(n24716), .B(n24715), .Z(n24792) );
  XOR U26115 ( .A(n24793), .B(n24792), .Z(n24794) );
  XNOR U26116 ( .A(n24795), .B(n24794), .Z(n24763) );
  NANDN U26117 ( .A(n24567), .B(n24566), .Z(n24571) );
  NANDN U26118 ( .A(n24569), .B(n24568), .Z(n24570) );
  NAND U26119 ( .A(n24571), .B(n24570), .Z(n24752) );
  AND U26120 ( .A(n24572), .B(o[252]), .Z(n24692) );
  AND U26121 ( .A(x[496]), .B(y[7917]), .Z(n24690) );
  AND U26122 ( .A(x[507]), .B(y[7906]), .Z(n24689) );
  XOR U26123 ( .A(n24690), .B(n24689), .Z(n24691) );
  XOR U26124 ( .A(n24692), .B(n24691), .Z(n24751) );
  AND U26125 ( .A(x[482]), .B(y[7931]), .Z(n24702) );
  XOR U26126 ( .A(n24702), .B(n24701), .Z(n24703) );
  XOR U26127 ( .A(n24704), .B(n24703), .Z(n24750) );
  XOR U26128 ( .A(n24751), .B(n24750), .Z(n24753) );
  XNOR U26129 ( .A(n24752), .B(n24753), .Z(n24762) );
  XOR U26130 ( .A(n24763), .B(n24762), .Z(n24764) );
  NANDN U26131 ( .A(n24574), .B(n24573), .Z(n24578) );
  NANDN U26132 ( .A(n24576), .B(n24575), .Z(n24577) );
  AND U26133 ( .A(n24578), .B(n24577), .Z(n24678) );
  NANDN U26134 ( .A(n24580), .B(n24579), .Z(n24584) );
  NANDN U26135 ( .A(n24582), .B(n24581), .Z(n24583) );
  NAND U26136 ( .A(n24584), .B(n24583), .Z(n24708) );
  NAND U26137 ( .A(n24586), .B(n24585), .Z(n24590) );
  NAND U26138 ( .A(n24588), .B(n24587), .Z(n24589) );
  NAND U26139 ( .A(n24590), .B(n24589), .Z(n24707) );
  XOR U26140 ( .A(n24708), .B(n24707), .Z(n24710) );
  AND U26141 ( .A(x[488]), .B(y[7925]), .Z(n24745) );
  AND U26142 ( .A(y[7927]), .B(x[486]), .Z(n24592) );
  NAND U26143 ( .A(y[7926]), .B(x[487]), .Z(n24591) );
  XNOR U26144 ( .A(n24592), .B(n24591), .Z(n24744) );
  XOR U26145 ( .A(n24745), .B(n24744), .Z(n24798) );
  NAND U26146 ( .A(x[489]), .B(y[7924]), .Z(n24877) );
  AND U26147 ( .A(x[485]), .B(y[7928]), .Z(n24698) );
  AND U26148 ( .A(x[484]), .B(y[7929]), .Z(n24696) );
  AND U26149 ( .A(x[490]), .B(y[7923]), .Z(n24695) );
  XOR U26150 ( .A(n24696), .B(n24695), .Z(n24697) );
  XNOR U26151 ( .A(n24698), .B(n24697), .Z(n24799) );
  XOR U26152 ( .A(n24877), .B(n24799), .Z(n24593) );
  XOR U26153 ( .A(n24798), .B(n24593), .Z(n24709) );
  XNOR U26154 ( .A(n24710), .B(n24709), .Z(n24677) );
  XOR U26155 ( .A(n24680), .B(n24679), .Z(n24769) );
  NAND U26156 ( .A(n24595), .B(n24594), .Z(n24599) );
  NANDN U26157 ( .A(n24597), .B(n24596), .Z(n24598) );
  NAND U26158 ( .A(n24599), .B(n24598), .Z(n24768) );
  XNOR U26159 ( .A(n24672), .B(n24671), .Z(n24673) );
  NANDN U26160 ( .A(n24601), .B(n24600), .Z(n24605) );
  NANDN U26161 ( .A(n24603), .B(n24602), .Z(n24604) );
  AND U26162 ( .A(n24605), .B(n24604), .Z(n24666) );
  XNOR U26163 ( .A(n24666), .B(n24665), .Z(n24667) );
  NANDN U26164 ( .A(n24611), .B(n24610), .Z(n24615) );
  NANDN U26165 ( .A(n24613), .B(n24612), .Z(n24614) );
  AND U26166 ( .A(n24615), .B(n24614), .Z(n24662) );
  NANDN U26167 ( .A(n24621), .B(n24620), .Z(n24625) );
  NAND U26168 ( .A(n24623), .B(n24622), .Z(n24624) );
  AND U26169 ( .A(n24625), .B(n24624), .Z(n24759) );
  XNOR U26170 ( .A(n24660), .B(n24659), .Z(n24661) );
  XOR U26171 ( .A(n24662), .B(n24661), .Z(n24668) );
  XOR U26172 ( .A(n24667), .B(n24668), .Z(n24674) );
  XOR U26173 ( .A(n24673), .B(n24674), .Z(n24656) );
  XOR U26174 ( .A(n24650), .B(n24649), .Z(n24646) );
  NAND U26175 ( .A(n24638), .B(n24637), .Z(n24642) );
  NAND U26176 ( .A(n24640), .B(n24639), .Z(n24641) );
  NAND U26177 ( .A(n24642), .B(n24641), .Z(n24644) );
  XOR U26178 ( .A(n24645), .B(n24644), .Z(n24643) );
  XNOR U26179 ( .A(n24646), .B(n24643), .Z(N510) );
  NANDN U26180 ( .A(n24648), .B(n24647), .Z(n24652) );
  NANDN U26181 ( .A(n24650), .B(n24649), .Z(n24651) );
  AND U26182 ( .A(n24652), .B(n24651), .Z(n25071) );
  NANDN U26183 ( .A(n24654), .B(n24653), .Z(n24658) );
  NANDN U26184 ( .A(n24656), .B(n24655), .Z(n24657) );
  AND U26185 ( .A(n24658), .B(n24657), .Z(n25088) );
  NANDN U26186 ( .A(n24660), .B(n24659), .Z(n24664) );
  NANDN U26187 ( .A(n24662), .B(n24661), .Z(n24663) );
  AND U26188 ( .A(n24664), .B(n24663), .Z(n24817) );
  NANDN U26189 ( .A(n24666), .B(n24665), .Z(n24670) );
  NANDN U26190 ( .A(n24668), .B(n24667), .Z(n24669) );
  AND U26191 ( .A(n24670), .B(n24669), .Z(n24819) );
  NANDN U26192 ( .A(n24672), .B(n24671), .Z(n24676) );
  NANDN U26193 ( .A(n24674), .B(n24673), .Z(n24675) );
  AND U26194 ( .A(n24676), .B(n24675), .Z(n24818) );
  XOR U26195 ( .A(n24819), .B(n24818), .Z(n24816) );
  XOR U26196 ( .A(n24817), .B(n24816), .Z(n25090) );
  NANDN U26197 ( .A(n24678), .B(n24677), .Z(n24682) );
  NAND U26198 ( .A(n24680), .B(n24679), .Z(n24681) );
  AND U26199 ( .A(n24682), .B(n24681), .Z(n25057) );
  NAND U26200 ( .A(n24684), .B(n24683), .Z(n24688) );
  NAND U26201 ( .A(n24686), .B(n24685), .Z(n24687) );
  AND U26202 ( .A(n24688), .B(n24687), .Z(n24825) );
  NAND U26203 ( .A(n24690), .B(n24689), .Z(n24694) );
  NAND U26204 ( .A(n24692), .B(n24691), .Z(n24693) );
  NAND U26205 ( .A(n24694), .B(n24693), .Z(n24835) );
  NAND U26206 ( .A(n24696), .B(n24695), .Z(n24700) );
  NAND U26207 ( .A(n24698), .B(n24697), .Z(n24699) );
  NAND U26208 ( .A(n24700), .B(n24699), .Z(n24838) );
  AND U26209 ( .A(x[486]), .B(y[7928]), .Z(n24944) );
  AND U26210 ( .A(x[485]), .B(y[7929]), .Z(n24946) );
  AND U26211 ( .A(x[499]), .B(y[7915]), .Z(n24945) );
  XOR U26212 ( .A(n24946), .B(n24945), .Z(n24943) );
  XNOR U26213 ( .A(n24944), .B(n24943), .Z(n24978) );
  AND U26214 ( .A(x[484]), .B(y[7930]), .Z(n24938) );
  AND U26215 ( .A(x[483]), .B(y[7931]), .Z(n24940) );
  AND U26216 ( .A(x[498]), .B(y[7916]), .Z(n24939) );
  XOR U26217 ( .A(n24940), .B(n24939), .Z(n24937) );
  XOR U26218 ( .A(n24938), .B(n24937), .Z(n24975) );
  NAND U26219 ( .A(n24702), .B(n24701), .Z(n24706) );
  NAND U26220 ( .A(n24704), .B(n24703), .Z(n24705) );
  AND U26221 ( .A(n24706), .B(n24705), .Z(n24976) );
  XOR U26222 ( .A(n24978), .B(n24977), .Z(n24837) );
  XOR U26223 ( .A(n24838), .B(n24837), .Z(n24836) );
  XOR U26224 ( .A(n24835), .B(n24836), .Z(n24826) );
  NAND U26225 ( .A(n24708), .B(n24707), .Z(n24712) );
  NAND U26226 ( .A(n24710), .B(n24709), .Z(n24711) );
  AND U26227 ( .A(n24712), .B(n24711), .Z(n24822) );
  XOR U26228 ( .A(n24823), .B(n24822), .Z(n25060) );
  AND U26229 ( .A(n24714), .B(n24713), .Z(n24718) );
  NAND U26230 ( .A(n24716), .B(n24715), .Z(n24717) );
  NANDN U26231 ( .A(n24718), .B(n24717), .Z(n24855) );
  AND U26232 ( .A(n24865), .B(n24719), .Z(n24723) );
  NAND U26233 ( .A(n24721), .B(n24720), .Z(n24722) );
  NANDN U26234 ( .A(n24723), .B(n24722), .Z(n24858) );
  NANDN U26235 ( .A(n24870), .B(n24724), .Z(n24728) );
  NANDN U26236 ( .A(n24726), .B(n24725), .Z(n24727) );
  AND U26237 ( .A(n24728), .B(n24727), .Z(n24842) );
  AND U26238 ( .A(x[503]), .B(y[7911]), .Z(n24932) );
  AND U26239 ( .A(y[7910]), .B(x[504]), .Z(n24730) );
  AND U26240 ( .A(y[7909]), .B(x[505]), .Z(n24729) );
  XOR U26241 ( .A(n24730), .B(n24729), .Z(n24931) );
  XOR U26242 ( .A(n24932), .B(n24931), .Z(n24844) );
  AND U26243 ( .A(n24731), .B(o[253]), .Z(n25004) );
  AND U26244 ( .A(x[508]), .B(y[7906]), .Z(n25006) );
  AND U26245 ( .A(x[496]), .B(y[7918]), .Z(n25005) );
  XOR U26246 ( .A(n25006), .B(n25005), .Z(n25003) );
  XNOR U26247 ( .A(n25004), .B(n25003), .Z(n24843) );
  XNOR U26248 ( .A(n24842), .B(n24841), .Z(n24857) );
  XOR U26249 ( .A(n24858), .B(n24857), .Z(n24856) );
  XOR U26250 ( .A(n24855), .B(n24856), .Z(n25040) );
  NAND U26251 ( .A(n24732), .B(n24934), .Z(n24736) );
  NAND U26252 ( .A(n24734), .B(n24733), .Z(n24735) );
  NAND U26253 ( .A(n24736), .B(n24735), .Z(n24832) );
  NAND U26254 ( .A(n24738), .B(n24737), .Z(n24742) );
  NAND U26255 ( .A(n24740), .B(n24739), .Z(n24741) );
  AND U26256 ( .A(n24742), .B(n24741), .Z(n24970) );
  AND U26257 ( .A(x[480]), .B(y[7934]), .Z(n24860) );
  AND U26258 ( .A(x[509]), .B(y[7905]), .Z(n24880) );
  XOR U26259 ( .A(o[254]), .B(n24880), .Z(n24862) );
  AND U26260 ( .A(x[510]), .B(y[7904]), .Z(n24861) );
  XOR U26261 ( .A(n24862), .B(n24861), .Z(n24859) );
  XOR U26262 ( .A(n24860), .B(n24859), .Z(n24972) );
  AND U26263 ( .A(x[500]), .B(y[7914]), .Z(n24999) );
  XOR U26264 ( .A(n25000), .B(n24999), .Z(n24998) );
  AND U26265 ( .A(x[488]), .B(y[7926]), .Z(n24997) );
  XNOR U26266 ( .A(n24998), .B(n24997), .Z(n24971) );
  XNOR U26267 ( .A(n24970), .B(n24969), .Z(n24831) );
  XOR U26268 ( .A(n24832), .B(n24831), .Z(n24829) );
  AND U26269 ( .A(x[487]), .B(y[7927]), .Z(n24869) );
  NAND U26270 ( .A(n24743), .B(n24869), .Z(n24747) );
  NAND U26271 ( .A(n24745), .B(n24744), .Z(n24746) );
  AND U26272 ( .A(n24747), .B(n24746), .Z(n24851) );
  AND U26273 ( .A(x[501]), .B(y[7913]), .Z(n24749) );
  AND U26274 ( .A(y[7912]), .B(x[502]), .Z(n24748) );
  XOR U26275 ( .A(n24749), .B(n24748), .Z(n24868) );
  XOR U26276 ( .A(n24869), .B(n24868), .Z(n24854) );
  AND U26277 ( .A(x[497]), .B(y[7917]), .Z(n24990) );
  AND U26278 ( .A(x[482]), .B(y[7932]), .Z(n24992) );
  AND U26279 ( .A(x[506]), .B(y[7908]), .Z(n24991) );
  XOR U26280 ( .A(n24992), .B(n24991), .Z(n24989) );
  XNOR U26281 ( .A(n24990), .B(n24989), .Z(n24853) );
  XNOR U26282 ( .A(n24851), .B(n24852), .Z(n24830) );
  XNOR U26283 ( .A(n24829), .B(n24830), .Z(n25042) );
  NAND U26284 ( .A(n24751), .B(n24750), .Z(n24755) );
  NAND U26285 ( .A(n24753), .B(n24752), .Z(n24754) );
  NAND U26286 ( .A(n24755), .B(n24754), .Z(n25041) );
  XOR U26287 ( .A(n25042), .B(n25041), .Z(n25039) );
  XOR U26288 ( .A(n25040), .B(n25039), .Z(n25059) );
  XNOR U26289 ( .A(n25057), .B(n25058), .Z(n25052) );
  NANDN U26290 ( .A(n24757), .B(n24756), .Z(n24761) );
  NANDN U26291 ( .A(n24759), .B(n24758), .Z(n24760) );
  AND U26292 ( .A(n24761), .B(n24760), .Z(n25054) );
  NAND U26293 ( .A(n24763), .B(n24762), .Z(n24767) );
  NANDN U26294 ( .A(n24765), .B(n24764), .Z(n24766) );
  NAND U26295 ( .A(n24767), .B(n24766), .Z(n25053) );
  XOR U26296 ( .A(n25054), .B(n25053), .Z(n25051) );
  XOR U26297 ( .A(n25052), .B(n25051), .Z(n25075) );
  NANDN U26298 ( .A(n24769), .B(n24768), .Z(n24773) );
  NANDN U26299 ( .A(n24771), .B(n24770), .Z(n24772) );
  NAND U26300 ( .A(n24773), .B(n24772), .Z(n25077) );
  NANDN U26301 ( .A(n24775), .B(n24774), .Z(n24779) );
  NAND U26302 ( .A(n24777), .B(n24776), .Z(n24778) );
  AND U26303 ( .A(n24779), .B(n24778), .Z(n25033) );
  NAND U26304 ( .A(n24781), .B(n24780), .Z(n24785) );
  NAND U26305 ( .A(n24783), .B(n24782), .Z(n24784) );
  AND U26306 ( .A(n24785), .B(n24784), .Z(n25024) );
  NAND U26307 ( .A(n24787), .B(n24786), .Z(n24791) );
  NANDN U26308 ( .A(n24789), .B(n24788), .Z(n24790) );
  AND U26309 ( .A(n24791), .B(n24790), .Z(n25023) );
  XOR U26310 ( .A(n25024), .B(n25023), .Z(n25022) );
  NAND U26311 ( .A(n24793), .B(n24792), .Z(n24797) );
  NAND U26312 ( .A(n24795), .B(n24794), .Z(n24796) );
  AND U26313 ( .A(n24797), .B(n24796), .Z(n25021) );
  XOR U26314 ( .A(n25022), .B(n25021), .Z(n25036) );
  NAND U26315 ( .A(n24801), .B(n24800), .Z(n24805) );
  NAND U26316 ( .A(n24803), .B(n24802), .Z(n24804) );
  NAND U26317 ( .A(n24805), .B(n24804), .Z(n24847) );
  AND U26318 ( .A(y[7922]), .B(x[492]), .Z(n24806) );
  XOR U26319 ( .A(n24807), .B(n24806), .Z(n24863) );
  XOR U26320 ( .A(n24864), .B(n24863), .Z(n24876) );
  AND U26321 ( .A(x[489]), .B(y[7925]), .Z(n24809) );
  XOR U26322 ( .A(n24809), .B(n24808), .Z(n24875) );
  XOR U26323 ( .A(n24876), .B(n24875), .Z(n24850) );
  AND U26324 ( .A(x[507]), .B(y[7907]), .Z(n24986) );
  AND U26325 ( .A(x[481]), .B(y[7933]), .Z(n24985) );
  XOR U26326 ( .A(n24986), .B(n24985), .Z(n24983) );
  XOR U26327 ( .A(n24984), .B(n24983), .Z(n24849) );
  XOR U26328 ( .A(n24850), .B(n24849), .Z(n24848) );
  XOR U26329 ( .A(n24847), .B(n24848), .Z(n25018) );
  NAND U26330 ( .A(n24811), .B(n24810), .Z(n24815) );
  NANDN U26331 ( .A(n24813), .B(n24812), .Z(n24814) );
  AND U26332 ( .A(n24815), .B(n24814), .Z(n25016) );
  XNOR U26333 ( .A(n25015), .B(n25016), .Z(n25035) );
  XNOR U26334 ( .A(n25033), .B(n25034), .Z(n25078) );
  XOR U26335 ( .A(n25077), .B(n25078), .Z(n25076) );
  XOR U26336 ( .A(n25075), .B(n25076), .Z(n25089) );
  XOR U26337 ( .A(n25088), .B(n25087), .Z(n25069) );
  XNOR U26338 ( .A(n25070), .B(n25069), .Z(N511) );
  NAND U26339 ( .A(n24817), .B(n24816), .Z(n24821) );
  NAND U26340 ( .A(n24819), .B(n24818), .Z(n24820) );
  AND U26341 ( .A(n24821), .B(n24820), .Z(n25086) );
  IV U26342 ( .A(n24822), .Z(n24824) );
  NANDN U26343 ( .A(n24824), .B(n24823), .Z(n24828) );
  NANDN U26344 ( .A(n24826), .B(n24825), .Z(n24827) );
  AND U26345 ( .A(n24828), .B(n24827), .Z(n25068) );
  NANDN U26346 ( .A(n24830), .B(n24829), .Z(n24834) );
  NAND U26347 ( .A(n24832), .B(n24831), .Z(n24833) );
  AND U26348 ( .A(n24834), .B(n24833), .Z(n25050) );
  NAND U26349 ( .A(n24836), .B(n24835), .Z(n24840) );
  NAND U26350 ( .A(n24838), .B(n24837), .Z(n24839) );
  AND U26351 ( .A(n24840), .B(n24839), .Z(n25032) );
  NAND U26352 ( .A(n24842), .B(n24841), .Z(n24846) );
  NANDN U26353 ( .A(n24844), .B(n24843), .Z(n24845) );
  AND U26354 ( .A(n24846), .B(n24845), .Z(n25014) );
  NAND U26355 ( .A(n24864), .B(n24863), .Z(n24867) );
  NAND U26356 ( .A(n24865), .B(n24900), .Z(n24866) );
  AND U26357 ( .A(n24867), .B(n24866), .Z(n24874) );
  NAND U26358 ( .A(n24869), .B(n24868), .Z(n24872) );
  AND U26359 ( .A(x[502]), .B(y[7913]), .Z(n24881) );
  NANDN U26360 ( .A(n24870), .B(n24881), .Z(n24871) );
  NAND U26361 ( .A(n24872), .B(n24871), .Z(n24873) );
  NAND U26362 ( .A(n24876), .B(n24875), .Z(n24879) );
  AND U26363 ( .A(x[490]), .B(y[7925]), .Z(n24899) );
  NANDN U26364 ( .A(n24877), .B(n24899), .Z(n24878) );
  AND U26365 ( .A(n24879), .B(n24878), .Z(n24930) );
  AND U26366 ( .A(y[7904]), .B(x[511]), .Z(n24888) );
  AND U26367 ( .A(n24880), .B(o[254]), .Z(n24886) );
  XOR U26368 ( .A(n24881), .B(o[255]), .Z(n24884) );
  AND U26369 ( .A(x[505]), .B(y[7910]), .Z(n24933) );
  XNOR U26370 ( .A(n24882), .B(n24933), .Z(n24883) );
  XNOR U26371 ( .A(n24884), .B(n24883), .Z(n24885) );
  XNOR U26372 ( .A(n24886), .B(n24885), .Z(n24887) );
  XNOR U26373 ( .A(n24888), .B(n24887), .Z(n24928) );
  AND U26374 ( .A(y[7905]), .B(x[510]), .Z(n24890) );
  NAND U26375 ( .A(y[7926]), .B(x[489]), .Z(n24889) );
  XNOR U26376 ( .A(n24890), .B(n24889), .Z(n24898) );
  AND U26377 ( .A(y[7906]), .B(x[509]), .Z(n24896) );
  AND U26378 ( .A(y[7934]), .B(x[481]), .Z(n24892) );
  NAND U26379 ( .A(y[7907]), .B(x[508]), .Z(n24891) );
  XNOR U26380 ( .A(n24892), .B(n24891), .Z(n24893) );
  XNOR U26381 ( .A(n24894), .B(n24893), .Z(n24895) );
  XNOR U26382 ( .A(n24896), .B(n24895), .Z(n24897) );
  XOR U26383 ( .A(n24898), .B(n24897), .Z(n24902) );
  XNOR U26384 ( .A(n24900), .B(n24899), .Z(n24901) );
  XNOR U26385 ( .A(n24902), .B(n24901), .Z(n24918) );
  AND U26386 ( .A(y[7924]), .B(x[491]), .Z(n24904) );
  NAND U26387 ( .A(y[7923]), .B(x[492]), .Z(n24903) );
  XNOR U26388 ( .A(n24904), .B(n24903), .Z(n24908) );
  AND U26389 ( .A(y[7927]), .B(x[488]), .Z(n24906) );
  NAND U26390 ( .A(y[7909]), .B(x[506]), .Z(n24905) );
  XNOR U26391 ( .A(n24906), .B(n24905), .Z(n24907) );
  XOR U26392 ( .A(n24908), .B(n24907), .Z(n24916) );
  AND U26393 ( .A(y[7919]), .B(x[496]), .Z(n24910) );
  NAND U26394 ( .A(y[7935]), .B(x[480]), .Z(n24909) );
  XNOR U26395 ( .A(n24910), .B(n24909), .Z(n24914) );
  AND U26396 ( .A(y[7921]), .B(x[494]), .Z(n24912) );
  NAND U26397 ( .A(y[7915]), .B(x[500]), .Z(n24911) );
  XNOR U26398 ( .A(n24912), .B(n24911), .Z(n24913) );
  XNOR U26399 ( .A(n24914), .B(n24913), .Z(n24915) );
  XNOR U26400 ( .A(n24916), .B(n24915), .Z(n24917) );
  XOR U26401 ( .A(n24918), .B(n24917), .Z(n24926) );
  AND U26402 ( .A(y[7930]), .B(x[485]), .Z(n24920) );
  NAND U26403 ( .A(y[7931]), .B(x[484]), .Z(n24919) );
  XNOR U26404 ( .A(n24920), .B(n24919), .Z(n24924) );
  AND U26405 ( .A(y[7929]), .B(x[486]), .Z(n24922) );
  NAND U26406 ( .A(y[7928]), .B(x[487]), .Z(n24921) );
  XNOR U26407 ( .A(n24922), .B(n24921), .Z(n24923) );
  XNOR U26408 ( .A(n24924), .B(n24923), .Z(n24925) );
  XNOR U26409 ( .A(n24926), .B(n24925), .Z(n24927) );
  XNOR U26410 ( .A(n24928), .B(n24927), .Z(n24929) );
  NAND U26411 ( .A(n24932), .B(n24931), .Z(n24936) );
  NAND U26412 ( .A(n24934), .B(n24933), .Z(n24935) );
  AND U26413 ( .A(n24936), .B(n24935), .Z(n24968) );
  NAND U26414 ( .A(n24938), .B(n24937), .Z(n24942) );
  NAND U26415 ( .A(n24940), .B(n24939), .Z(n24941) );
  AND U26416 ( .A(n24942), .B(n24941), .Z(n24950) );
  NAND U26417 ( .A(n24944), .B(n24943), .Z(n24948) );
  NAND U26418 ( .A(n24946), .B(n24945), .Z(n24947) );
  NAND U26419 ( .A(n24948), .B(n24947), .Z(n24949) );
  XNOR U26420 ( .A(n24950), .B(n24949), .Z(n24966) );
  AND U26421 ( .A(y[7932]), .B(x[483]), .Z(n24952) );
  NAND U26422 ( .A(y[7917]), .B(x[498]), .Z(n24951) );
  XNOR U26423 ( .A(n24952), .B(n24951), .Z(n24956) );
  AND U26424 ( .A(y[7916]), .B(x[499]), .Z(n24954) );
  NAND U26425 ( .A(y[7914]), .B(x[501]), .Z(n24953) );
  XNOR U26426 ( .A(n24954), .B(n24953), .Z(n24955) );
  XOR U26427 ( .A(n24956), .B(n24955), .Z(n24964) );
  AND U26428 ( .A(y[7933]), .B(x[482]), .Z(n24958) );
  NAND U26429 ( .A(y[7918]), .B(x[497]), .Z(n24957) );
  XNOR U26430 ( .A(n24958), .B(n24957), .Z(n24962) );
  AND U26431 ( .A(y[7908]), .B(x[507]), .Z(n24960) );
  NAND U26432 ( .A(y[7912]), .B(x[503]), .Z(n24959) );
  XNOR U26433 ( .A(n24960), .B(n24959), .Z(n24961) );
  XNOR U26434 ( .A(n24962), .B(n24961), .Z(n24963) );
  XNOR U26435 ( .A(n24964), .B(n24963), .Z(n24965) );
  XNOR U26436 ( .A(n24966), .B(n24965), .Z(n24967) );
  NAND U26437 ( .A(n24970), .B(n24969), .Z(n24974) );
  NANDN U26438 ( .A(n24972), .B(n24971), .Z(n24973) );
  AND U26439 ( .A(n24974), .B(n24973), .Z(n24982) );
  ANDN U26440 ( .B(n24976), .A(n24975), .Z(n24980) );
  ANDN U26441 ( .B(n24978), .A(n24977), .Z(n24979) );
  OR U26442 ( .A(n24980), .B(n24979), .Z(n24981) );
  NAND U26443 ( .A(n24984), .B(n24983), .Z(n24988) );
  NAND U26444 ( .A(n24986), .B(n24985), .Z(n24987) );
  AND U26445 ( .A(n24988), .B(n24987), .Z(n24996) );
  NAND U26446 ( .A(n24990), .B(n24989), .Z(n24994) );
  NAND U26447 ( .A(n24992), .B(n24991), .Z(n24993) );
  NAND U26448 ( .A(n24994), .B(n24993), .Z(n24995) );
  NAND U26449 ( .A(n24998), .B(n24997), .Z(n25002) );
  NAND U26450 ( .A(n25000), .B(n24999), .Z(n25001) );
  AND U26451 ( .A(n25002), .B(n25001), .Z(n25010) );
  NAND U26452 ( .A(n25004), .B(n25003), .Z(n25008) );
  NAND U26453 ( .A(n25006), .B(n25005), .Z(n25007) );
  NAND U26454 ( .A(n25008), .B(n25007), .Z(n25009) );
  XNOR U26455 ( .A(n25012), .B(n25011), .Z(n25013) );
  XNOR U26456 ( .A(n25014), .B(n25013), .Z(n25030) );
  NAND U26457 ( .A(n25016), .B(n25015), .Z(n25020) );
  NANDN U26458 ( .A(n25018), .B(n25017), .Z(n25019) );
  AND U26459 ( .A(n25020), .B(n25019), .Z(n25028) );
  NAND U26460 ( .A(n25024), .B(n25023), .Z(n25025) );
  NAND U26461 ( .A(n25026), .B(n25025), .Z(n25027) );
  XNOR U26462 ( .A(n25028), .B(n25027), .Z(n25029) );
  XNOR U26463 ( .A(n25030), .B(n25029), .Z(n25031) );
  XNOR U26464 ( .A(n25032), .B(n25031), .Z(n25048) );
  NANDN U26465 ( .A(n25034), .B(n25033), .Z(n25038) );
  NANDN U26466 ( .A(n25036), .B(n25035), .Z(n25037) );
  AND U26467 ( .A(n25038), .B(n25037), .Z(n25046) );
  NAND U26468 ( .A(n25040), .B(n25039), .Z(n25044) );
  NAND U26469 ( .A(n25042), .B(n25041), .Z(n25043) );
  NAND U26470 ( .A(n25044), .B(n25043), .Z(n25045) );
  XNOR U26471 ( .A(n25046), .B(n25045), .Z(n25047) );
  XNOR U26472 ( .A(n25048), .B(n25047), .Z(n25049) );
  XNOR U26473 ( .A(n25050), .B(n25049), .Z(n25066) );
  NANDN U26474 ( .A(n25052), .B(n25051), .Z(n25056) );
  NAND U26475 ( .A(n25054), .B(n25053), .Z(n25055) );
  AND U26476 ( .A(n25056), .B(n25055), .Z(n25064) );
  NANDN U26477 ( .A(n25058), .B(n25057), .Z(n25062) );
  NANDN U26478 ( .A(n25060), .B(n25059), .Z(n25061) );
  NAND U26479 ( .A(n25062), .B(n25061), .Z(n25063) );
  XNOR U26480 ( .A(n25064), .B(n25063), .Z(n25065) );
  XNOR U26481 ( .A(n25066), .B(n25065), .Z(n25067) );
  XNOR U26482 ( .A(n25068), .B(n25067), .Z(n25084) );
  NAND U26483 ( .A(n25070), .B(n25069), .Z(n25074) );
  NANDN U26484 ( .A(n25072), .B(n25071), .Z(n25073) );
  AND U26485 ( .A(n25074), .B(n25073), .Z(n25082) );
  NAND U26486 ( .A(n25076), .B(n25075), .Z(n25080) );
  NAND U26487 ( .A(n25078), .B(n25077), .Z(n25079) );
  NAND U26488 ( .A(n25080), .B(n25079), .Z(n25081) );
  XNOR U26489 ( .A(n25082), .B(n25081), .Z(n25083) );
  XNOR U26490 ( .A(n25084), .B(n25083), .Z(n25085) );
  XNOR U26491 ( .A(n25086), .B(n25085), .Z(n25094) );
  NANDN U26492 ( .A(n25088), .B(n25087), .Z(n25092) );
  NANDN U26493 ( .A(n25090), .B(n25089), .Z(n25091) );
  NAND U26494 ( .A(n25092), .B(n25091), .Z(n25093) );
  XNOR U26495 ( .A(n25094), .B(n25093), .Z(N512) );
  AND U26496 ( .A(x[480]), .B(y[7936]), .Z(n25741) );
  XOR U26497 ( .A(n25741), .B(o[256]), .Z(N545) );
  AND U26498 ( .A(x[481]), .B(y[7936]), .Z(n25103) );
  AND U26499 ( .A(x[480]), .B(y[7937]), .Z(n25102) );
  XNOR U26500 ( .A(n25102), .B(o[257]), .Z(n25095) );
  XNOR U26501 ( .A(n25103), .B(n25095), .Z(n25097) );
  NAND U26502 ( .A(n25741), .B(o[256]), .Z(n25096) );
  XNOR U26503 ( .A(n25097), .B(n25096), .Z(N546) );
  NANDN U26504 ( .A(n25103), .B(n25095), .Z(n25099) );
  NAND U26505 ( .A(n25097), .B(n25096), .Z(n25098) );
  AND U26506 ( .A(n25099), .B(n25098), .Z(n25109) );
  AND U26507 ( .A(x[480]), .B(y[7938]), .Z(n25116) );
  XNOR U26508 ( .A(n25116), .B(o[258]), .Z(n25108) );
  XNOR U26509 ( .A(n25109), .B(n25108), .Z(n25111) );
  AND U26510 ( .A(y[7936]), .B(x[482]), .Z(n25101) );
  NAND U26511 ( .A(y[7937]), .B(x[481]), .Z(n25100) );
  XNOR U26512 ( .A(n25101), .B(n25100), .Z(n25105) );
  AND U26513 ( .A(n25102), .B(o[257]), .Z(n25104) );
  XNOR U26514 ( .A(n25105), .B(n25104), .Z(n25110) );
  XNOR U26515 ( .A(n25111), .B(n25110), .Z(N547) );
  AND U26516 ( .A(x[482]), .B(y[7937]), .Z(n25123) );
  NAND U26517 ( .A(n25123), .B(n25103), .Z(n25107) );
  NAND U26518 ( .A(n25105), .B(n25104), .Z(n25106) );
  AND U26519 ( .A(n25107), .B(n25106), .Z(n25126) );
  NANDN U26520 ( .A(n25109), .B(n25108), .Z(n25113) );
  NAND U26521 ( .A(n25111), .B(n25110), .Z(n25112) );
  AND U26522 ( .A(n25113), .B(n25112), .Z(n25125) );
  XNOR U26523 ( .A(n25126), .B(n25125), .Z(n25128) );
  AND U26524 ( .A(x[481]), .B(y[7938]), .Z(n25241) );
  XOR U26525 ( .A(n25123), .B(o[259]), .Z(n25131) );
  XOR U26526 ( .A(n25241), .B(n25131), .Z(n25133) );
  AND U26527 ( .A(y[7936]), .B(x[483]), .Z(n25115) );
  NAND U26528 ( .A(y[7939]), .B(x[480]), .Z(n25114) );
  XNOR U26529 ( .A(n25115), .B(n25114), .Z(n25118) );
  AND U26530 ( .A(n25116), .B(o[258]), .Z(n25117) );
  XOR U26531 ( .A(n25118), .B(n25117), .Z(n25132) );
  XOR U26532 ( .A(n25133), .B(n25132), .Z(n25127) );
  XOR U26533 ( .A(n25128), .B(n25127), .Z(N548) );
  AND U26534 ( .A(x[483]), .B(y[7939]), .Z(n25176) );
  NAND U26535 ( .A(n25741), .B(n25176), .Z(n25120) );
  NAND U26536 ( .A(n25118), .B(n25117), .Z(n25119) );
  NAND U26537 ( .A(n25120), .B(n25119), .Z(n25154) );
  AND U26538 ( .A(y[7940]), .B(x[480]), .Z(n25122) );
  NAND U26539 ( .A(y[7936]), .B(x[484]), .Z(n25121) );
  XNOR U26540 ( .A(n25122), .B(n25121), .Z(n25147) );
  AND U26541 ( .A(n25123), .B(o[259]), .Z(n25148) );
  XOR U26542 ( .A(n25147), .B(n25148), .Z(n25152) );
  AND U26543 ( .A(y[7938]), .B(x[482]), .Z(n25297) );
  NAND U26544 ( .A(y[7939]), .B(x[481]), .Z(n25124) );
  XNOR U26545 ( .A(n25297), .B(n25124), .Z(n25144) );
  AND U26546 ( .A(x[483]), .B(y[7937]), .Z(n25139) );
  XOR U26547 ( .A(o[260]), .B(n25139), .Z(n25143) );
  XOR U26548 ( .A(n25144), .B(n25143), .Z(n25151) );
  XOR U26549 ( .A(n25152), .B(n25151), .Z(n25153) );
  XOR U26550 ( .A(n25154), .B(n25153), .Z(n25158) );
  NANDN U26551 ( .A(n25126), .B(n25125), .Z(n25130) );
  NAND U26552 ( .A(n25128), .B(n25127), .Z(n25129) );
  NAND U26553 ( .A(n25130), .B(n25129), .Z(n25159) );
  NAND U26554 ( .A(n25241), .B(n25131), .Z(n25135) );
  NAND U26555 ( .A(n25133), .B(n25132), .Z(n25134) );
  NAND U26556 ( .A(n25135), .B(n25134), .Z(n25160) );
  IV U26557 ( .A(n25160), .Z(n25157) );
  XOR U26558 ( .A(n25159), .B(n25157), .Z(n25136) );
  XNOR U26559 ( .A(n25158), .B(n25136), .Z(N549) );
  AND U26560 ( .A(y[7938]), .B(x[483]), .Z(n25138) );
  NAND U26561 ( .A(y[7940]), .B(x[481]), .Z(n25137) );
  XNOR U26562 ( .A(n25138), .B(n25137), .Z(n25163) );
  AND U26563 ( .A(x[484]), .B(y[7937]), .Z(n25174) );
  XOR U26564 ( .A(n25174), .B(o[261]), .Z(n25162) );
  XNOR U26565 ( .A(n25163), .B(n25162), .Z(n25166) );
  AND U26566 ( .A(x[482]), .B(y[7939]), .Z(n25250) );
  AND U26567 ( .A(o[260]), .B(n25139), .Z(n25168) );
  AND U26568 ( .A(y[7936]), .B(x[485]), .Z(n25141) );
  NAND U26569 ( .A(y[7941]), .B(x[480]), .Z(n25140) );
  XNOR U26570 ( .A(n25141), .B(n25140), .Z(n25169) );
  XOR U26571 ( .A(n25168), .B(n25169), .Z(n25167) );
  XNOR U26572 ( .A(n25250), .B(n25167), .Z(n25142) );
  XOR U26573 ( .A(n25166), .B(n25142), .Z(n25184) );
  NAND U26574 ( .A(n25250), .B(n25241), .Z(n25146) );
  NAND U26575 ( .A(n25144), .B(n25143), .Z(n25145) );
  NAND U26576 ( .A(n25146), .B(n25145), .Z(n25182) );
  AND U26577 ( .A(x[484]), .B(y[7940]), .Z(n25943) );
  NAND U26578 ( .A(n25943), .B(n25741), .Z(n25150) );
  NAND U26579 ( .A(n25148), .B(n25147), .Z(n25149) );
  NAND U26580 ( .A(n25150), .B(n25149), .Z(n25181) );
  XOR U26581 ( .A(n25182), .B(n25181), .Z(n25183) );
  XNOR U26582 ( .A(n25184), .B(n25183), .Z(n25180) );
  NAND U26583 ( .A(n25152), .B(n25151), .Z(n25156) );
  NAND U26584 ( .A(n25154), .B(n25153), .Z(n25155) );
  NAND U26585 ( .A(n25156), .B(n25155), .Z(n25179) );
  XOR U26586 ( .A(n25179), .B(n25178), .Z(n25161) );
  XNOR U26587 ( .A(n25180), .B(n25161), .Z(N550) );
  AND U26588 ( .A(x[483]), .B(y[7940]), .Z(n25251) );
  NAND U26589 ( .A(n25251), .B(n25241), .Z(n25165) );
  NAND U26590 ( .A(n25163), .B(n25162), .Z(n25164) );
  NAND U26591 ( .A(n25165), .B(n25164), .Z(n25219) );
  XOR U26592 ( .A(n25219), .B(n25220), .Z(n25222) );
  AND U26593 ( .A(x[485]), .B(y[7941]), .Z(n25421) );
  NAND U26594 ( .A(n25741), .B(n25421), .Z(n25171) );
  NAND U26595 ( .A(n25169), .B(n25168), .Z(n25170) );
  NAND U26596 ( .A(n25171), .B(n25170), .Z(n25189) );
  AND U26597 ( .A(y[7936]), .B(x[486]), .Z(n25173) );
  NAND U26598 ( .A(y[7942]), .B(x[480]), .Z(n25172) );
  XNOR U26599 ( .A(n25173), .B(n25172), .Z(n25195) );
  AND U26600 ( .A(n25174), .B(o[261]), .Z(n25196) );
  XOR U26601 ( .A(n25195), .B(n25196), .Z(n25188) );
  XOR U26602 ( .A(n25189), .B(n25188), .Z(n25191) );
  NAND U26603 ( .A(y[7940]), .B(x[482]), .Z(n25175) );
  XNOR U26604 ( .A(n25176), .B(n25175), .Z(n25200) );
  AND U26605 ( .A(y[7941]), .B(x[481]), .Z(n25442) );
  NAND U26606 ( .A(y[7938]), .B(x[484]), .Z(n25177) );
  XNOR U26607 ( .A(n25442), .B(n25177), .Z(n25204) );
  AND U26608 ( .A(x[485]), .B(y[7937]), .Z(n25211) );
  XOR U26609 ( .A(o[262]), .B(n25211), .Z(n25203) );
  XOR U26610 ( .A(n25204), .B(n25203), .Z(n25199) );
  XOR U26611 ( .A(n25200), .B(n25199), .Z(n25190) );
  XOR U26612 ( .A(n25191), .B(n25190), .Z(n25221) );
  XOR U26613 ( .A(n25222), .B(n25221), .Z(n25215) );
  NAND U26614 ( .A(n25182), .B(n25181), .Z(n25186) );
  NAND U26615 ( .A(n25184), .B(n25183), .Z(n25185) );
  AND U26616 ( .A(n25186), .B(n25185), .Z(n25214) );
  IV U26617 ( .A(n25214), .Z(n25212) );
  XOR U26618 ( .A(n25213), .B(n25212), .Z(n25187) );
  XNOR U26619 ( .A(n25215), .B(n25187), .Z(N551) );
  NAND U26620 ( .A(n25189), .B(n25188), .Z(n25193) );
  NAND U26621 ( .A(n25191), .B(n25190), .Z(n25192) );
  AND U26622 ( .A(n25193), .B(n25192), .Z(n25229) );
  AND U26623 ( .A(y[7938]), .B(x[485]), .Z(n25320) );
  NAND U26624 ( .A(y[7942]), .B(x[481]), .Z(n25194) );
  XNOR U26625 ( .A(n25320), .B(n25194), .Z(n25243) );
  AND U26626 ( .A(x[486]), .B(y[7937]), .Z(n25247) );
  XOR U26627 ( .A(o[263]), .B(n25247), .Z(n25242) );
  XNOR U26628 ( .A(n25243), .B(n25242), .Z(n25262) );
  AND U26629 ( .A(x[486]), .B(y[7942]), .Z(n25462) );
  NAND U26630 ( .A(n25741), .B(n25462), .Z(n25198) );
  NAND U26631 ( .A(n25196), .B(n25195), .Z(n25197) );
  AND U26632 ( .A(n25198), .B(n25197), .Z(n25261) );
  XOR U26633 ( .A(n25262), .B(n25261), .Z(n25263) );
  NAND U26634 ( .A(n25250), .B(n25251), .Z(n25202) );
  NAND U26635 ( .A(n25200), .B(n25199), .Z(n25201) );
  AND U26636 ( .A(n25202), .B(n25201), .Z(n25264) );
  XOR U26637 ( .A(n25263), .B(n25264), .Z(n25227) );
  AND U26638 ( .A(x[484]), .B(y[7941]), .Z(n25746) );
  NAND U26639 ( .A(n25746), .B(n25241), .Z(n25206) );
  NAND U26640 ( .A(n25204), .B(n25203), .Z(n25205) );
  AND U26641 ( .A(n25206), .B(n25205), .Z(n25238) );
  AND U26642 ( .A(y[7941]), .B(x[482]), .Z(n25208) );
  NAND U26643 ( .A(y[7939]), .B(x[484]), .Z(n25207) );
  XNOR U26644 ( .A(n25208), .B(n25207), .Z(n25252) );
  XNOR U26645 ( .A(n25252), .B(n25251), .Z(n25236) );
  AND U26646 ( .A(y[7936]), .B(x[487]), .Z(n25210) );
  NAND U26647 ( .A(y[7943]), .B(x[480]), .Z(n25209) );
  XNOR U26648 ( .A(n25210), .B(n25209), .Z(n25256) );
  AND U26649 ( .A(o[262]), .B(n25211), .Z(n25255) );
  XNOR U26650 ( .A(n25256), .B(n25255), .Z(n25235) );
  XOR U26651 ( .A(n25236), .B(n25235), .Z(n25237) );
  XOR U26652 ( .A(n25238), .B(n25237), .Z(n25226) );
  XOR U26653 ( .A(n25227), .B(n25226), .Z(n25228) );
  XNOR U26654 ( .A(n25229), .B(n25228), .Z(n25234) );
  NANDN U26655 ( .A(n25212), .B(n25213), .Z(n25218) );
  NOR U26656 ( .A(n25214), .B(n25213), .Z(n25216) );
  OR U26657 ( .A(n25216), .B(n25215), .Z(n25217) );
  AND U26658 ( .A(n25218), .B(n25217), .Z(n25233) );
  NAND U26659 ( .A(n25220), .B(n25219), .Z(n25224) );
  NAND U26660 ( .A(n25222), .B(n25221), .Z(n25223) );
  AND U26661 ( .A(n25224), .B(n25223), .Z(n25232) );
  XOR U26662 ( .A(n25233), .B(n25232), .Z(n25225) );
  XNOR U26663 ( .A(n25234), .B(n25225), .Z(N552) );
  NAND U26664 ( .A(n25227), .B(n25226), .Z(n25231) );
  NAND U26665 ( .A(n25229), .B(n25228), .Z(n25230) );
  AND U26666 ( .A(n25231), .B(n25230), .Z(n25275) );
  NAND U26667 ( .A(n25236), .B(n25235), .Z(n25240) );
  NAND U26668 ( .A(n25238), .B(n25237), .Z(n25239) );
  AND U26669 ( .A(n25240), .B(n25239), .Z(n25310) );
  AND U26670 ( .A(x[485]), .B(y[7942]), .Z(n25413) );
  NAND U26671 ( .A(n25413), .B(n25241), .Z(n25245) );
  NAND U26672 ( .A(n25243), .B(n25242), .Z(n25244) );
  NAND U26673 ( .A(n25245), .B(n25244), .Z(n25308) );
  AND U26674 ( .A(y[7939]), .B(x[485]), .Z(n25846) );
  NAND U26675 ( .A(y[7943]), .B(x[481]), .Z(n25246) );
  XNOR U26676 ( .A(n25846), .B(n25246), .Z(n25289) );
  AND U26677 ( .A(o[263]), .B(n25247), .Z(n25288) );
  XOR U26678 ( .A(n25289), .B(n25288), .Z(n25294) );
  NAND U26679 ( .A(x[483]), .B(y[7941]), .Z(n26070) );
  AND U26680 ( .A(y[7938]), .B(x[486]), .Z(n25249) );
  NAND U26681 ( .A(y[7942]), .B(x[482]), .Z(n25248) );
  XNOR U26682 ( .A(n25249), .B(n25248), .Z(n25298) );
  XNOR U26683 ( .A(n25943), .B(n25298), .Z(n25292) );
  XOR U26684 ( .A(n26070), .B(n25292), .Z(n25293) );
  XOR U26685 ( .A(n25294), .B(n25293), .Z(n25307) );
  XOR U26686 ( .A(n25308), .B(n25307), .Z(n25309) );
  XNOR U26687 ( .A(n25310), .B(n25309), .Z(n25271) );
  NAND U26688 ( .A(n25250), .B(n25746), .Z(n25254) );
  NAND U26689 ( .A(n25252), .B(n25251), .Z(n25253) );
  NAND U26690 ( .A(n25254), .B(n25253), .Z(n25304) );
  AND U26691 ( .A(x[487]), .B(y[7943]), .Z(n25624) );
  NAND U26692 ( .A(n25741), .B(n25624), .Z(n25258) );
  NAND U26693 ( .A(n25256), .B(n25255), .Z(n25257) );
  NAND U26694 ( .A(n25258), .B(n25257), .Z(n25302) );
  AND U26695 ( .A(y[7936]), .B(x[488]), .Z(n25260) );
  NAND U26696 ( .A(y[7944]), .B(x[480]), .Z(n25259) );
  XNOR U26697 ( .A(n25260), .B(n25259), .Z(n25279) );
  AND U26698 ( .A(x[487]), .B(y[7937]), .Z(n25284) );
  XOR U26699 ( .A(o[264]), .B(n25284), .Z(n25278) );
  XOR U26700 ( .A(n25279), .B(n25278), .Z(n25301) );
  XOR U26701 ( .A(n25302), .B(n25301), .Z(n25303) );
  XNOR U26702 ( .A(n25304), .B(n25303), .Z(n25269) );
  NAND U26703 ( .A(n25262), .B(n25261), .Z(n25266) );
  NAND U26704 ( .A(n25264), .B(n25263), .Z(n25265) );
  NAND U26705 ( .A(n25266), .B(n25265), .Z(n25268) );
  XOR U26706 ( .A(n25269), .B(n25268), .Z(n25270) );
  XOR U26707 ( .A(n25271), .B(n25270), .Z(n25276) );
  XNOR U26708 ( .A(n25274), .B(n25276), .Z(n25267) );
  XOR U26709 ( .A(n25275), .B(n25267), .Z(N553) );
  NAND U26710 ( .A(n25269), .B(n25268), .Z(n25273) );
  NAND U26711 ( .A(n25271), .B(n25270), .Z(n25272) );
  NAND U26712 ( .A(n25273), .B(n25272), .Z(n25364) );
  IV U26713 ( .A(n25364), .Z(n25362) );
  AND U26714 ( .A(x[488]), .B(y[7944]), .Z(n25277) );
  NAND U26715 ( .A(n25277), .B(n25741), .Z(n25281) );
  NAND U26716 ( .A(n25279), .B(n25278), .Z(n25280) );
  AND U26717 ( .A(n25281), .B(n25280), .Z(n25349) );
  AND U26718 ( .A(y[7940]), .B(x[485]), .Z(n25283) );
  NAND U26719 ( .A(y[7938]), .B(x[487]), .Z(n25282) );
  XNOR U26720 ( .A(n25283), .B(n25282), .Z(n25322) );
  AND U26721 ( .A(o[264]), .B(n25284), .Z(n25321) );
  XOR U26722 ( .A(n25322), .B(n25321), .Z(n25347) );
  AND U26723 ( .A(y[7936]), .B(x[489]), .Z(n25286) );
  NAND U26724 ( .A(y[7945]), .B(x[480]), .Z(n25285) );
  XNOR U26725 ( .A(n25286), .B(n25285), .Z(n25329) );
  AND U26726 ( .A(x[488]), .B(y[7937]), .Z(n25338) );
  XOR U26727 ( .A(o[265]), .B(n25338), .Z(n25328) );
  XNOR U26728 ( .A(n25329), .B(n25328), .Z(n25346) );
  XNOR U26729 ( .A(n25349), .B(n25348), .Z(n25343) );
  AND U26730 ( .A(y[7939]), .B(x[486]), .Z(n25689) );
  NAND U26731 ( .A(y[7944]), .B(x[481]), .Z(n25287) );
  XNOR U26732 ( .A(n25689), .B(n25287), .Z(n25333) );
  XNOR U26733 ( .A(n25746), .B(n25333), .Z(n25352) );
  NAND U26734 ( .A(x[482]), .B(y[7943]), .Z(n25988) );
  AND U26735 ( .A(x[483]), .B(y[7942]), .Z(n25699) );
  XOR U26736 ( .A(n25988), .B(n25699), .Z(n25353) );
  XOR U26737 ( .A(n25352), .B(n25353), .Z(n25341) );
  NAND U26738 ( .A(x[485]), .B(y[7943]), .Z(n25538) );
  AND U26739 ( .A(x[481]), .B(y[7939]), .Z(n25332) );
  NANDN U26740 ( .A(n25538), .B(n25332), .Z(n25291) );
  NAND U26741 ( .A(n25289), .B(n25288), .Z(n25290) );
  NAND U26742 ( .A(n25291), .B(n25290), .Z(n25340) );
  XOR U26743 ( .A(n25341), .B(n25340), .Z(n25342) );
  XNOR U26744 ( .A(n25343), .B(n25342), .Z(n25316) );
  NAND U26745 ( .A(n26070), .B(n25292), .Z(n25296) );
  NANDN U26746 ( .A(n25294), .B(n25293), .Z(n25295) );
  NAND U26747 ( .A(n25296), .B(n25295), .Z(n25315) );
  NAND U26748 ( .A(n25462), .B(n25297), .Z(n25300) );
  NAND U26749 ( .A(n25943), .B(n25298), .Z(n25299) );
  AND U26750 ( .A(n25300), .B(n25299), .Z(n25314) );
  XOR U26751 ( .A(n25315), .B(n25314), .Z(n25317) );
  XNOR U26752 ( .A(n25316), .B(n25317), .Z(n25358) );
  NAND U26753 ( .A(n25302), .B(n25301), .Z(n25306) );
  NAND U26754 ( .A(n25304), .B(n25303), .Z(n25305) );
  NAND U26755 ( .A(n25306), .B(n25305), .Z(n25357) );
  NAND U26756 ( .A(n25308), .B(n25307), .Z(n25312) );
  NAND U26757 ( .A(n25310), .B(n25309), .Z(n25311) );
  NAND U26758 ( .A(n25312), .B(n25311), .Z(n25356) );
  XOR U26759 ( .A(n25357), .B(n25356), .Z(n25359) );
  XOR U26760 ( .A(n25358), .B(n25359), .Z(n25365) );
  XNOR U26761 ( .A(n25363), .B(n25365), .Z(n25313) );
  XOR U26762 ( .A(n25362), .B(n25313), .Z(N554) );
  NAND U26763 ( .A(n25315), .B(n25314), .Z(n25319) );
  NAND U26764 ( .A(n25317), .B(n25316), .Z(n25318) );
  NAND U26765 ( .A(n25319), .B(n25318), .Z(n25373) );
  AND U26766 ( .A(x[487]), .B(y[7940]), .Z(n25415) );
  NAND U26767 ( .A(n25415), .B(n25320), .Z(n25324) );
  NAND U26768 ( .A(n25322), .B(n25321), .Z(n25323) );
  AND U26769 ( .A(n25324), .B(n25323), .Z(n25428) );
  AND U26770 ( .A(y[7939]), .B(x[487]), .Z(n25326) );
  NAND U26771 ( .A(y[7942]), .B(x[484]), .Z(n25325) );
  XNOR U26772 ( .A(n25326), .B(n25325), .Z(n25399) );
  AND U26773 ( .A(x[486]), .B(y[7940]), .Z(n25398) );
  XNOR U26774 ( .A(n25399), .B(n25398), .Z(n25426) );
  AND U26775 ( .A(x[488]), .B(y[7938]), .Z(n25598) );
  AND U26776 ( .A(x[489]), .B(y[7937]), .Z(n25409) );
  XOR U26777 ( .A(o[266]), .B(n25409), .Z(n25420) );
  XOR U26778 ( .A(n25598), .B(n25420), .Z(n25422) );
  XNOR U26779 ( .A(n25422), .B(n25421), .Z(n25425) );
  XOR U26780 ( .A(n25426), .B(n25425), .Z(n25427) );
  XNOR U26781 ( .A(n25428), .B(n25427), .Z(n25387) );
  AND U26782 ( .A(x[489]), .B(y[7945]), .Z(n25327) );
  NAND U26783 ( .A(n25327), .B(n25741), .Z(n25331) );
  NAND U26784 ( .A(n25329), .B(n25328), .Z(n25330) );
  NAND U26785 ( .A(n25331), .B(n25330), .Z(n25385) );
  AND U26786 ( .A(x[486]), .B(y[7944]), .Z(n25634) );
  NAND U26787 ( .A(n25634), .B(n25332), .Z(n25335) );
  NAND U26788 ( .A(n25333), .B(n25746), .Z(n25334) );
  NAND U26789 ( .A(n25335), .B(n25334), .Z(n25394) );
  AND U26790 ( .A(y[7936]), .B(x[490]), .Z(n25337) );
  NAND U26791 ( .A(y[7946]), .B(x[480]), .Z(n25336) );
  XNOR U26792 ( .A(n25337), .B(n25336), .Z(n25404) );
  AND U26793 ( .A(o[265]), .B(n25338), .Z(n25403) );
  XOR U26794 ( .A(n25404), .B(n25403), .Z(n25392) );
  AND U26795 ( .A(y[7943]), .B(x[483]), .Z(n26293) );
  NAND U26796 ( .A(y[7945]), .B(x[481]), .Z(n25339) );
  XNOR U26797 ( .A(n26293), .B(n25339), .Z(n25416) );
  AND U26798 ( .A(x[482]), .B(y[7944]), .Z(n25417) );
  XOR U26799 ( .A(n25416), .B(n25417), .Z(n25391) );
  XOR U26800 ( .A(n25392), .B(n25391), .Z(n25393) );
  XNOR U26801 ( .A(n25394), .B(n25393), .Z(n25386) );
  XOR U26802 ( .A(n25385), .B(n25386), .Z(n25388) );
  XOR U26803 ( .A(n25387), .B(n25388), .Z(n25371) );
  NAND U26804 ( .A(n25341), .B(n25340), .Z(n25345) );
  NAND U26805 ( .A(n25343), .B(n25342), .Z(n25344) );
  NAND U26806 ( .A(n25345), .B(n25344), .Z(n25381) );
  NANDN U26807 ( .A(n25347), .B(n25346), .Z(n25351) );
  NAND U26808 ( .A(n25349), .B(n25348), .Z(n25350) );
  AND U26809 ( .A(n25351), .B(n25350), .Z(n25380) );
  NANDN U26810 ( .A(n25353), .B(n25352), .Z(n25355) );
  ANDN U26811 ( .B(n25988), .A(n25699), .Z(n25354) );
  ANDN U26812 ( .B(n25355), .A(n25354), .Z(n25379) );
  XOR U26813 ( .A(n25380), .B(n25379), .Z(n25382) );
  XNOR U26814 ( .A(n25381), .B(n25382), .Z(n25370) );
  XOR U26815 ( .A(n25371), .B(n25370), .Z(n25372) );
  XOR U26816 ( .A(n25373), .B(n25372), .Z(n25378) );
  NAND U26817 ( .A(n25357), .B(n25356), .Z(n25361) );
  NAND U26818 ( .A(n25359), .B(n25358), .Z(n25360) );
  NAND U26819 ( .A(n25361), .B(n25360), .Z(n25377) );
  NANDN U26820 ( .A(n25362), .B(n25363), .Z(n25368) );
  NOR U26821 ( .A(n25364), .B(n25363), .Z(n25366) );
  OR U26822 ( .A(n25366), .B(n25365), .Z(n25367) );
  AND U26823 ( .A(n25368), .B(n25367), .Z(n25376) );
  XOR U26824 ( .A(n25377), .B(n25376), .Z(n25369) );
  XNOR U26825 ( .A(n25378), .B(n25369), .Z(N555) );
  NAND U26826 ( .A(n25371), .B(n25370), .Z(n25375) );
  NAND U26827 ( .A(n25373), .B(n25372), .Z(n25374) );
  NAND U26828 ( .A(n25375), .B(n25374), .Z(n25489) );
  IV U26829 ( .A(n25489), .Z(n25487) );
  NAND U26830 ( .A(n25380), .B(n25379), .Z(n25384) );
  NAND U26831 ( .A(n25382), .B(n25381), .Z(n25383) );
  NAND U26832 ( .A(n25384), .B(n25383), .Z(n25496) );
  NANDN U26833 ( .A(n25386), .B(n25385), .Z(n25390) );
  NANDN U26834 ( .A(n25388), .B(n25387), .Z(n25389) );
  NAND U26835 ( .A(n25390), .B(n25389), .Z(n25495) );
  NAND U26836 ( .A(n25392), .B(n25391), .Z(n25396) );
  NAND U26837 ( .A(n25394), .B(n25393), .Z(n25395) );
  NAND U26838 ( .A(n25396), .B(n25395), .Z(n25483) );
  AND U26839 ( .A(x[487]), .B(y[7942]), .Z(n25533) );
  AND U26840 ( .A(x[484]), .B(y[7939]), .Z(n25397) );
  NAND U26841 ( .A(n25533), .B(n25397), .Z(n25401) );
  NAND U26842 ( .A(n25399), .B(n25398), .Z(n25400) );
  NAND U26843 ( .A(n25401), .B(n25400), .Z(n25481) );
  AND U26844 ( .A(x[490]), .B(y[7946]), .Z(n25402) );
  NAND U26845 ( .A(n25402), .B(n25741), .Z(n25406) );
  NAND U26846 ( .A(n25404), .B(n25403), .Z(n25405) );
  NAND U26847 ( .A(n25406), .B(n25405), .Z(n25477) );
  AND U26848 ( .A(y[7936]), .B(x[491]), .Z(n25408) );
  NAND U26849 ( .A(y[7947]), .B(x[480]), .Z(n25407) );
  XNOR U26850 ( .A(n25408), .B(n25407), .Z(n25453) );
  AND U26851 ( .A(o[266]), .B(n25409), .Z(n25452) );
  XOR U26852 ( .A(n25453), .B(n25452), .Z(n25476) );
  AND U26853 ( .A(y[7941]), .B(x[486]), .Z(n25411) );
  NAND U26854 ( .A(y[7946]), .B(x[481]), .Z(n25410) );
  XNOR U26855 ( .A(n25411), .B(n25410), .Z(n25444) );
  AND U26856 ( .A(x[490]), .B(y[7937]), .Z(n25463) );
  XOR U26857 ( .A(o[267]), .B(n25463), .Z(n25443) );
  XOR U26858 ( .A(n25444), .B(n25443), .Z(n25475) );
  XOR U26859 ( .A(n25476), .B(n25475), .Z(n25478) );
  XOR U26860 ( .A(n25477), .B(n25478), .Z(n25482) );
  XNOR U26861 ( .A(n25481), .B(n25482), .Z(n25484) );
  XOR U26862 ( .A(n25483), .B(n25484), .Z(n25466) );
  NAND U26863 ( .A(x[483]), .B(y[7944]), .Z(n26450) );
  NAND U26864 ( .A(y[7945]), .B(x[482]), .Z(n25412) );
  XNOR U26865 ( .A(n25413), .B(n25412), .Z(n25439) );
  AND U26866 ( .A(x[484]), .B(y[7943]), .Z(n25438) );
  XNOR U26867 ( .A(n25439), .B(n25438), .Z(n25470) );
  XOR U26868 ( .A(n26450), .B(n25470), .Z(n25472) );
  NAND U26869 ( .A(y[7938]), .B(x[489]), .Z(n25414) );
  XNOR U26870 ( .A(n25415), .B(n25414), .Z(n25458) );
  AND U26871 ( .A(x[488]), .B(y[7939]), .Z(n25457) );
  XNOR U26872 ( .A(n25458), .B(n25457), .Z(n25471) );
  XNOR U26873 ( .A(n25472), .B(n25471), .Z(n25435) );
  NAND U26874 ( .A(x[483]), .B(y[7945]), .Z(n25529) );
  AND U26875 ( .A(x[481]), .B(y[7943]), .Z(n25736) );
  NANDN U26876 ( .A(n25529), .B(n25736), .Z(n25419) );
  NAND U26877 ( .A(n25417), .B(n25416), .Z(n25418) );
  NAND U26878 ( .A(n25419), .B(n25418), .Z(n25433) );
  NAND U26879 ( .A(n25598), .B(n25420), .Z(n25424) );
  NAND U26880 ( .A(n25422), .B(n25421), .Z(n25423) );
  NAND U26881 ( .A(n25424), .B(n25423), .Z(n25432) );
  XOR U26882 ( .A(n25433), .B(n25432), .Z(n25434) );
  XNOR U26883 ( .A(n25435), .B(n25434), .Z(n25465) );
  NAND U26884 ( .A(n25426), .B(n25425), .Z(n25430) );
  NAND U26885 ( .A(n25428), .B(n25427), .Z(n25429) );
  NAND U26886 ( .A(n25430), .B(n25429), .Z(n25464) );
  XOR U26887 ( .A(n25465), .B(n25464), .Z(n25467) );
  XNOR U26888 ( .A(n25466), .B(n25467), .Z(n25494) );
  XOR U26889 ( .A(n25495), .B(n25494), .Z(n25497) );
  XOR U26890 ( .A(n25496), .B(n25497), .Z(n25490) );
  XNOR U26891 ( .A(n25488), .B(n25490), .Z(n25431) );
  XOR U26892 ( .A(n25487), .B(n25431), .Z(N556) );
  NAND U26893 ( .A(n25433), .B(n25432), .Z(n25437) );
  NAND U26894 ( .A(n25435), .B(n25434), .Z(n25436) );
  NAND U26895 ( .A(n25437), .B(n25436), .Z(n25569) );
  AND U26896 ( .A(x[482]), .B(y[7942]), .Z(n26147) );
  AND U26897 ( .A(x[485]), .B(y[7945]), .Z(n25981) );
  NAND U26898 ( .A(n26147), .B(n25981), .Z(n25441) );
  NAND U26899 ( .A(n25439), .B(n25438), .Z(n25440) );
  NAND U26900 ( .A(n25441), .B(n25440), .Z(n25517) );
  AND U26901 ( .A(x[486]), .B(y[7946]), .Z(n25753) );
  NAND U26902 ( .A(n25753), .B(n25442), .Z(n25446) );
  NAND U26903 ( .A(n25444), .B(n25443), .Z(n25445) );
  NAND U26904 ( .A(n25446), .B(n25445), .Z(n25516) );
  XOR U26905 ( .A(n25517), .B(n25516), .Z(n25519) );
  AND U26906 ( .A(x[489]), .B(y[7939]), .Z(n26142) );
  AND U26907 ( .A(y[7938]), .B(x[490]), .Z(n26197) );
  NAND U26908 ( .A(y[7944]), .B(x[484]), .Z(n25447) );
  XOR U26909 ( .A(n26197), .B(n25447), .Z(n25560) );
  NAND U26910 ( .A(x[487]), .B(y[7941]), .Z(n25537) );
  XOR U26911 ( .A(n25538), .B(n25537), .Z(n25540) );
  AND U26912 ( .A(y[7936]), .B(x[492]), .Z(n25449) );
  NAND U26913 ( .A(y[7948]), .B(x[480]), .Z(n25448) );
  XNOR U26914 ( .A(n25449), .B(n25448), .Z(n25554) );
  AND U26915 ( .A(x[491]), .B(y[7937]), .Z(n25534) );
  XOR U26916 ( .A(o[268]), .B(n25534), .Z(n25553) );
  XOR U26917 ( .A(n25554), .B(n25553), .Z(n25523) );
  AND U26918 ( .A(y[7946]), .B(x[482]), .Z(n25451) );
  NAND U26919 ( .A(y[7940]), .B(x[488]), .Z(n25450) );
  XNOR U26920 ( .A(n25451), .B(n25450), .Z(n25528) );
  XOR U26921 ( .A(n25523), .B(n25522), .Z(n25525) );
  XOR U26922 ( .A(n25524), .B(n25525), .Z(n25518) );
  XOR U26923 ( .A(n25519), .B(n25518), .Z(n25568) );
  AND U26924 ( .A(x[491]), .B(y[7947]), .Z(n26537) );
  NAND U26925 ( .A(n26537), .B(n25741), .Z(n25455) );
  NAND U26926 ( .A(n25453), .B(n25452), .Z(n25454) );
  NAND U26927 ( .A(n25455), .B(n25454), .Z(n25546) );
  AND U26928 ( .A(x[487]), .B(y[7938]), .Z(n25675) );
  AND U26929 ( .A(x[489]), .B(y[7940]), .Z(n25456) );
  NAND U26930 ( .A(n25675), .B(n25456), .Z(n25460) );
  NAND U26931 ( .A(n25458), .B(n25457), .Z(n25459) );
  NAND U26932 ( .A(n25460), .B(n25459), .Z(n25544) );
  NAND U26933 ( .A(y[7947]), .B(x[481]), .Z(n25461) );
  XNOR U26934 ( .A(n25462), .B(n25461), .Z(n25550) );
  AND U26935 ( .A(o[267]), .B(n25463), .Z(n25549) );
  XOR U26936 ( .A(n25550), .B(n25549), .Z(n25543) );
  XOR U26937 ( .A(n25544), .B(n25543), .Z(n25545) );
  XOR U26938 ( .A(n25546), .B(n25545), .Z(n25567) );
  XOR U26939 ( .A(n25568), .B(n25567), .Z(n25570) );
  XNOR U26940 ( .A(n25569), .B(n25570), .Z(n25502) );
  NAND U26941 ( .A(n25465), .B(n25464), .Z(n25469) );
  NAND U26942 ( .A(n25467), .B(n25466), .Z(n25468) );
  NAND U26943 ( .A(n25469), .B(n25468), .Z(n25501) );
  XOR U26944 ( .A(n25502), .B(n25501), .Z(n25504) );
  IV U26945 ( .A(n26450), .Z(n26156) );
  NANDN U26946 ( .A(n26156), .B(n25470), .Z(n25474) );
  NAND U26947 ( .A(n25472), .B(n25471), .Z(n25473) );
  NAND U26948 ( .A(n25474), .B(n25473), .Z(n25510) );
  NAND U26949 ( .A(n25476), .B(n25475), .Z(n25480) );
  NAND U26950 ( .A(n25478), .B(n25477), .Z(n25479) );
  AND U26951 ( .A(n25480), .B(n25479), .Z(n25511) );
  XOR U26952 ( .A(n25510), .B(n25511), .Z(n25513) );
  NAND U26953 ( .A(n25482), .B(n25481), .Z(n25486) );
  NANDN U26954 ( .A(n25484), .B(n25483), .Z(n25485) );
  AND U26955 ( .A(n25486), .B(n25485), .Z(n25512) );
  XOR U26956 ( .A(n25513), .B(n25512), .Z(n25503) );
  XNOR U26957 ( .A(n25504), .B(n25503), .Z(n25509) );
  NANDN U26958 ( .A(n25487), .B(n25488), .Z(n25493) );
  NOR U26959 ( .A(n25489), .B(n25488), .Z(n25491) );
  OR U26960 ( .A(n25491), .B(n25490), .Z(n25492) );
  AND U26961 ( .A(n25493), .B(n25492), .Z(n25508) );
  NAND U26962 ( .A(n25495), .B(n25494), .Z(n25499) );
  NAND U26963 ( .A(n25497), .B(n25496), .Z(n25498) );
  AND U26964 ( .A(n25499), .B(n25498), .Z(n25507) );
  XOR U26965 ( .A(n25508), .B(n25507), .Z(n25500) );
  XNOR U26966 ( .A(n25509), .B(n25500), .Z(N557) );
  NAND U26967 ( .A(n25502), .B(n25501), .Z(n25506) );
  NAND U26968 ( .A(n25504), .B(n25503), .Z(n25505) );
  AND U26969 ( .A(n25506), .B(n25505), .Z(n25648) );
  NAND U26970 ( .A(n25511), .B(n25510), .Z(n25515) );
  NAND U26971 ( .A(n25513), .B(n25512), .Z(n25514) );
  NAND U26972 ( .A(n25515), .B(n25514), .Z(n25643) );
  NAND U26973 ( .A(n25517), .B(n25516), .Z(n25521) );
  NAND U26974 ( .A(n25519), .B(n25518), .Z(n25520) );
  AND U26975 ( .A(n25521), .B(n25520), .Z(n25575) );
  NAND U26976 ( .A(n25523), .B(n25522), .Z(n25527) );
  NAND U26977 ( .A(n25525), .B(n25524), .Z(n25526) );
  NAND U26978 ( .A(n25527), .B(n25526), .Z(n25582) );
  AND U26979 ( .A(y[7946]), .B(x[488]), .Z(n26794) );
  AND U26980 ( .A(x[482]), .B(y[7940]), .Z(n25685) );
  NAND U26981 ( .A(n26794), .B(n25685), .Z(n25531) );
  NANDN U26982 ( .A(n25529), .B(n25528), .Z(n25530) );
  NAND U26983 ( .A(n25531), .B(n25530), .Z(n25613) );
  NAND U26984 ( .A(y[7948]), .B(x[481]), .Z(n25532) );
  XNOR U26985 ( .A(n25533), .B(n25532), .Z(n25604) );
  AND U26986 ( .A(o[268]), .B(n25534), .Z(n25603) );
  XOR U26987 ( .A(n25604), .B(n25603), .Z(n25611) );
  AND U26988 ( .A(x[486]), .B(y[7943]), .Z(n26577) );
  AND U26989 ( .A(y[7947]), .B(x[482]), .Z(n25536) );
  NAND U26990 ( .A(y[7940]), .B(x[489]), .Z(n25535) );
  XNOR U26991 ( .A(n25536), .B(n25535), .Z(n25617) );
  XOR U26992 ( .A(n26577), .B(n25617), .Z(n25610) );
  XOR U26993 ( .A(n25611), .B(n25610), .Z(n25612) );
  XOR U26994 ( .A(n25613), .B(n25612), .Z(n25581) );
  NAND U26995 ( .A(n25538), .B(n25537), .Z(n25542) );
  ANDN U26996 ( .B(n25540), .A(n25539), .Z(n25541) );
  ANDN U26997 ( .B(n25542), .A(n25541), .Z(n25580) );
  XOR U26998 ( .A(n25581), .B(n25580), .Z(n25583) );
  XOR U26999 ( .A(n25582), .B(n25583), .Z(n25574) );
  NAND U27000 ( .A(n25544), .B(n25543), .Z(n25548) );
  NAND U27001 ( .A(n25546), .B(n25545), .Z(n25547) );
  AND U27002 ( .A(n25548), .B(n25547), .Z(n25589) );
  NAND U27003 ( .A(x[486]), .B(y[7947]), .Z(n25983) );
  AND U27004 ( .A(x[481]), .B(y[7942]), .Z(n25602) );
  NANDN U27005 ( .A(n25983), .B(n25602), .Z(n25552) );
  NAND U27006 ( .A(n25550), .B(n25549), .Z(n25551) );
  NAND U27007 ( .A(n25552), .B(n25551), .Z(n25595) );
  AND U27008 ( .A(x[492]), .B(y[7948]), .Z(n26800) );
  NAND U27009 ( .A(n26800), .B(n25741), .Z(n25556) );
  NAND U27010 ( .A(n25554), .B(n25553), .Z(n25555) );
  NAND U27011 ( .A(n25556), .B(n25555), .Z(n25593) );
  AND U27012 ( .A(x[490]), .B(y[7939]), .Z(n26462) );
  AND U27013 ( .A(y[7938]), .B(x[491]), .Z(n26423) );
  NAND U27014 ( .A(y[7941]), .B(x[488]), .Z(n25557) );
  XNOR U27015 ( .A(n26423), .B(n25557), .Z(n25599) );
  XOR U27016 ( .A(n26462), .B(n25599), .Z(n25592) );
  XOR U27017 ( .A(n25593), .B(n25592), .Z(n25594) );
  XOR U27018 ( .A(n25595), .B(n25594), .Z(n25587) );
  AND U27019 ( .A(x[490]), .B(y[7944]), .Z(n25559) );
  AND U27020 ( .A(x[484]), .B(y[7938]), .Z(n25558) );
  NAND U27021 ( .A(n25559), .B(n25558), .Z(n25562) );
  NANDN U27022 ( .A(n25560), .B(n26142), .Z(n25561) );
  AND U27023 ( .A(n25562), .B(n25561), .Z(n25638) );
  AND U27024 ( .A(y[7936]), .B(x[493]), .Z(n25564) );
  NAND U27025 ( .A(y[7949]), .B(x[480]), .Z(n25563) );
  XNOR U27026 ( .A(n25564), .B(n25563), .Z(n25630) );
  AND U27027 ( .A(x[492]), .B(y[7937]), .Z(n25622) );
  XOR U27028 ( .A(o[269]), .B(n25622), .Z(n25629) );
  XOR U27029 ( .A(n25630), .B(n25629), .Z(n25636) );
  AND U27030 ( .A(y[7944]), .B(x[485]), .Z(n25566) );
  NAND U27031 ( .A(y[7946]), .B(x[483]), .Z(n25565) );
  XNOR U27032 ( .A(n25566), .B(n25565), .Z(n25625) );
  AND U27033 ( .A(x[484]), .B(y[7945]), .Z(n25626) );
  XOR U27034 ( .A(n25625), .B(n25626), .Z(n25635) );
  XOR U27035 ( .A(n25636), .B(n25635), .Z(n25637) );
  XOR U27036 ( .A(n25587), .B(n25586), .Z(n25588) );
  XNOR U27037 ( .A(n25577), .B(n25576), .Z(n25642) );
  NAND U27038 ( .A(n25568), .B(n25567), .Z(n25572) );
  NAND U27039 ( .A(n25570), .B(n25569), .Z(n25571) );
  AND U27040 ( .A(n25572), .B(n25571), .Z(n25641) );
  XOR U27041 ( .A(n25642), .B(n25641), .Z(n25644) );
  XOR U27042 ( .A(n25643), .B(n25644), .Z(n25649) );
  XNOR U27043 ( .A(n25647), .B(n25649), .Z(n25573) );
  XOR U27044 ( .A(n25648), .B(n25573), .Z(N558) );
  NANDN U27045 ( .A(n25575), .B(n25574), .Z(n25579) );
  NAND U27046 ( .A(n25577), .B(n25576), .Z(n25578) );
  AND U27047 ( .A(n25579), .B(n25578), .Z(n25727) );
  NAND U27048 ( .A(n25581), .B(n25580), .Z(n25585) );
  NAND U27049 ( .A(n25583), .B(n25582), .Z(n25584) );
  NAND U27050 ( .A(n25585), .B(n25584), .Z(n25726) );
  NAND U27051 ( .A(n25587), .B(n25586), .Z(n25591) );
  NANDN U27052 ( .A(n25589), .B(n25588), .Z(n25590) );
  AND U27053 ( .A(n25591), .B(n25590), .Z(n25654) );
  NAND U27054 ( .A(n25593), .B(n25592), .Z(n25597) );
  NAND U27055 ( .A(n25595), .B(n25594), .Z(n25596) );
  AND U27056 ( .A(n25597), .B(n25596), .Z(n25660) );
  AND U27057 ( .A(x[491]), .B(y[7941]), .Z(n25767) );
  NAND U27058 ( .A(n25767), .B(n25598), .Z(n25601) );
  NAND U27059 ( .A(n25599), .B(n26462), .Z(n25600) );
  NAND U27060 ( .A(n25601), .B(n25600), .Z(n25715) );
  NAND U27061 ( .A(x[487]), .B(y[7948]), .Z(n26158) );
  NANDN U27062 ( .A(n26158), .B(n25602), .Z(n25606) );
  NAND U27063 ( .A(n25604), .B(n25603), .Z(n25605) );
  NAND U27064 ( .A(n25606), .B(n25605), .Z(n25714) );
  XOR U27065 ( .A(n25715), .B(n25714), .Z(n25717) );
  AND U27066 ( .A(x[484]), .B(y[7946]), .Z(n26079) );
  AND U27067 ( .A(y[7947]), .B(x[483]), .Z(n25608) );
  NAND U27068 ( .A(y[7942]), .B(x[488]), .Z(n25607) );
  XNOR U27069 ( .A(n25608), .B(n25607), .Z(n25700) );
  XOR U27070 ( .A(n25981), .B(n25700), .Z(n25709) );
  XOR U27071 ( .A(n26079), .B(n25709), .Z(n25711) );
  AND U27072 ( .A(x[489]), .B(y[7941]), .Z(n26264) );
  AND U27073 ( .A(y[7948]), .B(x[482]), .Z(n25609) );
  AND U27074 ( .A(y[7940]), .B(x[490]), .Z(n26288) );
  XOR U27075 ( .A(n25609), .B(n26288), .Z(n25686) );
  XOR U27076 ( .A(n26264), .B(n25686), .Z(n25710) );
  XOR U27077 ( .A(n25711), .B(n25710), .Z(n25716) );
  XNOR U27078 ( .A(n25717), .B(n25716), .Z(n25658) );
  NAND U27079 ( .A(n25611), .B(n25610), .Z(n25615) );
  NAND U27080 ( .A(n25613), .B(n25612), .Z(n25614) );
  AND U27081 ( .A(n25615), .B(n25614), .Z(n25657) );
  XOR U27082 ( .A(n25658), .B(n25657), .Z(n25659) );
  XOR U27083 ( .A(n25660), .B(n25659), .Z(n25652) );
  AND U27084 ( .A(x[489]), .B(y[7947]), .Z(n25616) );
  NAND U27085 ( .A(n25616), .B(n25685), .Z(n25619) );
  NAND U27086 ( .A(n25617), .B(n26577), .Z(n25618) );
  NAND U27087 ( .A(n25619), .B(n25618), .Z(n25672) );
  AND U27088 ( .A(y[7936]), .B(x[494]), .Z(n25621) );
  NAND U27089 ( .A(y[7950]), .B(x[480]), .Z(n25620) );
  XNOR U27090 ( .A(n25621), .B(n25620), .Z(n25695) );
  AND U27091 ( .A(o[269]), .B(n25622), .Z(n25694) );
  XOR U27092 ( .A(n25695), .B(n25694), .Z(n25670) );
  NAND U27093 ( .A(y[7938]), .B(x[492]), .Z(n25623) );
  XNOR U27094 ( .A(n25624), .B(n25623), .Z(n25677) );
  AND U27095 ( .A(x[493]), .B(y[7937]), .Z(n25684) );
  XOR U27096 ( .A(o[270]), .B(n25684), .Z(n25676) );
  XOR U27097 ( .A(n25677), .B(n25676), .Z(n25669) );
  XOR U27098 ( .A(n25670), .B(n25669), .Z(n25671) );
  XNOR U27099 ( .A(n25672), .B(n25671), .Z(n25721) );
  AND U27100 ( .A(x[485]), .B(y[7946]), .Z(n25754) );
  NANDN U27101 ( .A(n26450), .B(n25754), .Z(n25628) );
  NAND U27102 ( .A(n25626), .B(n25625), .Z(n25627) );
  AND U27103 ( .A(n25628), .B(n25627), .Z(n25666) );
  AND U27104 ( .A(x[493]), .B(y[7949]), .Z(n27200) );
  NAND U27105 ( .A(n27200), .B(n25741), .Z(n25632) );
  NAND U27106 ( .A(n25630), .B(n25629), .Z(n25631) );
  NAND U27107 ( .A(n25632), .B(n25631), .Z(n25664) );
  NAND U27108 ( .A(y[7939]), .B(x[491]), .Z(n25633) );
  XNOR U27109 ( .A(n25634), .B(n25633), .Z(n25691) );
  AND U27110 ( .A(x[481]), .B(y[7949]), .Z(n25690) );
  XOR U27111 ( .A(n25691), .B(n25690), .Z(n25663) );
  XOR U27112 ( .A(n25664), .B(n25663), .Z(n25665) );
  XOR U27113 ( .A(n25666), .B(n25665), .Z(n25720) );
  XOR U27114 ( .A(n25721), .B(n25720), .Z(n25723) );
  NAND U27115 ( .A(n25636), .B(n25635), .Z(n25640) );
  NANDN U27116 ( .A(n25638), .B(n25637), .Z(n25639) );
  AND U27117 ( .A(n25640), .B(n25639), .Z(n25722) );
  XNOR U27118 ( .A(n25723), .B(n25722), .Z(n25651) );
  XNOR U27119 ( .A(n25729), .B(n25728), .Z(n25734) );
  NAND U27120 ( .A(n25642), .B(n25641), .Z(n25646) );
  NAND U27121 ( .A(n25644), .B(n25643), .Z(n25645) );
  AND U27122 ( .A(n25646), .B(n25645), .Z(n25732) );
  XNOR U27123 ( .A(n25732), .B(n25733), .Z(n25650) );
  XNOR U27124 ( .A(n25734), .B(n25650), .Z(N559) );
  NANDN U27125 ( .A(n25652), .B(n25651), .Z(n25656) );
  NANDN U27126 ( .A(n25654), .B(n25653), .Z(n25655) );
  AND U27127 ( .A(n25656), .B(n25655), .Z(n25824) );
  NAND U27128 ( .A(n25658), .B(n25657), .Z(n25662) );
  NAND U27129 ( .A(n25660), .B(n25659), .Z(n25661) );
  NAND U27130 ( .A(n25662), .B(n25661), .Z(n25797) );
  NAND U27131 ( .A(n25664), .B(n25663), .Z(n25668) );
  NANDN U27132 ( .A(n25666), .B(n25665), .Z(n25667) );
  NAND U27133 ( .A(n25668), .B(n25667), .Z(n25802) );
  NAND U27134 ( .A(n25670), .B(n25669), .Z(n25674) );
  NAND U27135 ( .A(n25672), .B(n25671), .Z(n25673) );
  NAND U27136 ( .A(n25674), .B(n25673), .Z(n25800) );
  NAND U27137 ( .A(x[492]), .B(y[7943]), .Z(n26149) );
  NANDN U27138 ( .A(n26149), .B(n25675), .Z(n25679) );
  NAND U27139 ( .A(n25677), .B(n25676), .Z(n25678) );
  AND U27140 ( .A(n25679), .B(n25678), .Z(n25777) );
  AND U27141 ( .A(y[7940]), .B(x[491]), .Z(n25681) );
  NAND U27142 ( .A(y[7938]), .B(x[493]), .Z(n25680) );
  XNOR U27143 ( .A(n25681), .B(n25680), .Z(n25781) );
  AND U27144 ( .A(x[492]), .B(y[7939]), .Z(n25780) );
  XNOR U27145 ( .A(n25781), .B(n25780), .Z(n25775) );
  AND U27146 ( .A(y[7936]), .B(x[495]), .Z(n25683) );
  NAND U27147 ( .A(y[7951]), .B(x[480]), .Z(n25682) );
  XNOR U27148 ( .A(n25683), .B(n25682), .Z(n25743) );
  AND U27149 ( .A(o[270]), .B(n25684), .Z(n25742) );
  XNOR U27150 ( .A(n25743), .B(n25742), .Z(n25774) );
  XOR U27151 ( .A(n25775), .B(n25774), .Z(n25776) );
  XNOR U27152 ( .A(n25777), .B(n25776), .Z(n25808) );
  NAND U27153 ( .A(x[490]), .B(y[7948]), .Z(n26579) );
  NANDN U27154 ( .A(n26579), .B(n25685), .Z(n25688) );
  NAND U27155 ( .A(n26264), .B(n25686), .Z(n25687) );
  NAND U27156 ( .A(n25688), .B(n25687), .Z(n25807) );
  AND U27157 ( .A(x[491]), .B(y[7944]), .Z(n26078) );
  NAND U27158 ( .A(n26078), .B(n25689), .Z(n25693) );
  NAND U27159 ( .A(n25691), .B(n25690), .Z(n25692) );
  NAND U27160 ( .A(n25693), .B(n25692), .Z(n25806) );
  XNOR U27161 ( .A(n25807), .B(n25806), .Z(n25809) );
  XOR U27162 ( .A(n25800), .B(n25801), .Z(n25803) );
  XOR U27163 ( .A(n25802), .B(n25803), .Z(n25794) );
  AND U27164 ( .A(x[494]), .B(y[7950]), .Z(n27457) );
  NAND U27165 ( .A(n27457), .B(n25741), .Z(n25697) );
  NAND U27166 ( .A(n25695), .B(n25694), .Z(n25696) );
  NAND U27167 ( .A(n25697), .B(n25696), .Z(n25769) );
  AND U27168 ( .A(x[488]), .B(y[7947]), .Z(n25698) );
  NAND U27169 ( .A(n25699), .B(n25698), .Z(n25702) );
  NAND U27170 ( .A(n25700), .B(n25981), .Z(n25701) );
  NAND U27171 ( .A(n25702), .B(n25701), .Z(n25768) );
  XOR U27172 ( .A(n25769), .B(n25768), .Z(n25771) );
  AND U27173 ( .A(y[7941]), .B(x[490]), .Z(n25704) );
  NAND U27174 ( .A(y[7947]), .B(x[484]), .Z(n25703) );
  XNOR U27175 ( .A(n25704), .B(n25703), .Z(n25749) );
  AND U27176 ( .A(x[487]), .B(y[7944]), .Z(n25748) );
  XNOR U27177 ( .A(n25749), .B(n25748), .Z(n25756) );
  NAND U27178 ( .A(x[486]), .B(y[7945]), .Z(n25855) );
  XNOR U27179 ( .A(n25855), .B(n25754), .Z(n25755) );
  XNOR U27180 ( .A(n25756), .B(n25755), .Z(n25790) );
  AND U27181 ( .A(y[7949]), .B(x[482]), .Z(n25706) );
  NAND U27182 ( .A(y[7942]), .B(x[489]), .Z(n25705) );
  XNOR U27183 ( .A(n25706), .B(n25705), .Z(n25759) );
  AND U27184 ( .A(x[483]), .B(y[7948]), .Z(n25760) );
  XOR U27185 ( .A(n25759), .B(n25760), .Z(n25789) );
  AND U27186 ( .A(y[7950]), .B(x[481]), .Z(n25708) );
  NAND U27187 ( .A(y[7943]), .B(x[488]), .Z(n25707) );
  XNOR U27188 ( .A(n25708), .B(n25707), .Z(n25738) );
  AND U27189 ( .A(x[494]), .B(y[7937]), .Z(n25765) );
  XOR U27190 ( .A(o[271]), .B(n25765), .Z(n25737) );
  XOR U27191 ( .A(n25738), .B(n25737), .Z(n25788) );
  XOR U27192 ( .A(n25789), .B(n25788), .Z(n25791) );
  XOR U27193 ( .A(n25790), .B(n25791), .Z(n25770) );
  XOR U27194 ( .A(n25771), .B(n25770), .Z(n25813) );
  NAND U27195 ( .A(n26079), .B(n25709), .Z(n25713) );
  NAND U27196 ( .A(n25711), .B(n25710), .Z(n25712) );
  AND U27197 ( .A(n25713), .B(n25712), .Z(n25812) );
  NAND U27198 ( .A(n25715), .B(n25714), .Z(n25719) );
  NAND U27199 ( .A(n25717), .B(n25716), .Z(n25718) );
  AND U27200 ( .A(n25719), .B(n25718), .Z(n25814) );
  XOR U27201 ( .A(n25815), .B(n25814), .Z(n25795) );
  XOR U27202 ( .A(n25794), .B(n25795), .Z(n25796) );
  XNOR U27203 ( .A(n25797), .B(n25796), .Z(n25821) );
  NAND U27204 ( .A(n25721), .B(n25720), .Z(n25725) );
  NAND U27205 ( .A(n25723), .B(n25722), .Z(n25724) );
  AND U27206 ( .A(n25725), .B(n25724), .Z(n25822) );
  XOR U27207 ( .A(n25821), .B(n25822), .Z(n25823) );
  XOR U27208 ( .A(n25824), .B(n25823), .Z(n25820) );
  NANDN U27209 ( .A(n25727), .B(n25726), .Z(n25731) );
  NAND U27210 ( .A(n25729), .B(n25728), .Z(n25730) );
  NAND U27211 ( .A(n25731), .B(n25730), .Z(n25818) );
  XOR U27212 ( .A(n25818), .B(n25819), .Z(n25735) );
  XNOR U27213 ( .A(n25820), .B(n25735), .Z(N560) );
  AND U27214 ( .A(x[488]), .B(y[7950]), .Z(n26080) );
  NAND U27215 ( .A(n26080), .B(n25736), .Z(n25740) );
  NAND U27216 ( .A(n25738), .B(n25737), .Z(n25739) );
  NAND U27217 ( .A(n25740), .B(n25739), .Z(n25885) );
  AND U27218 ( .A(x[495]), .B(y[7951]), .Z(n27804) );
  NAND U27219 ( .A(n27804), .B(n25741), .Z(n25745) );
  NAND U27220 ( .A(n25743), .B(n25742), .Z(n25744) );
  NAND U27221 ( .A(n25745), .B(n25744), .Z(n25884) );
  XOR U27222 ( .A(n25885), .B(n25884), .Z(n25887) );
  AND U27223 ( .A(x[490]), .B(y[7947]), .Z(n25747) );
  NAND U27224 ( .A(n25747), .B(n25746), .Z(n25751) );
  NAND U27225 ( .A(n25749), .B(n25748), .Z(n25750) );
  NAND U27226 ( .A(n25751), .B(n25750), .Z(n25842) );
  AND U27227 ( .A(x[480]), .B(y[7952]), .Z(n25864) );
  AND U27228 ( .A(x[496]), .B(y[7936]), .Z(n25865) );
  XOR U27229 ( .A(n25864), .B(n25865), .Z(n25866) );
  NAND U27230 ( .A(x[495]), .B(y[7937]), .Z(n25852) );
  XNOR U27231 ( .A(o[272]), .B(n25852), .Z(n25867) );
  XOR U27232 ( .A(n25866), .B(n25867), .Z(n25841) );
  NAND U27233 ( .A(y[7945]), .B(x[487]), .Z(n25752) );
  XNOR U27234 ( .A(n25753), .B(n25752), .Z(n25857) );
  AND U27235 ( .A(x[490]), .B(y[7942]), .Z(n25856) );
  XOR U27236 ( .A(n25857), .B(n25856), .Z(n25840) );
  XOR U27237 ( .A(n25841), .B(n25840), .Z(n25843) );
  XOR U27238 ( .A(n25842), .B(n25843), .Z(n25886) );
  XOR U27239 ( .A(n25887), .B(n25886), .Z(n25837) );
  NANDN U27240 ( .A(n25754), .B(n25855), .Z(n25758) );
  NAND U27241 ( .A(n25756), .B(n25755), .Z(n25757) );
  AND U27242 ( .A(n25758), .B(n25757), .Z(n25835) );
  NAND U27243 ( .A(x[489]), .B(y[7949]), .Z(n26560) );
  NANDN U27244 ( .A(n26560), .B(n26147), .Z(n25762) );
  NAND U27245 ( .A(n25760), .B(n25759), .Z(n25761) );
  AND U27246 ( .A(n25762), .B(n25761), .Z(n25875) );
  AND U27247 ( .A(y[7951]), .B(x[481]), .Z(n25764) );
  NAND U27248 ( .A(y[7944]), .B(x[488]), .Z(n25763) );
  XNOR U27249 ( .A(n25764), .B(n25763), .Z(n25861) );
  AND U27250 ( .A(o[271]), .B(n25765), .Z(n25860) );
  XOR U27251 ( .A(n25861), .B(n25860), .Z(n25872) );
  NAND U27252 ( .A(y[7938]), .B(x[494]), .Z(n25766) );
  XNOR U27253 ( .A(n25767), .B(n25766), .Z(n25896) );
  NAND U27254 ( .A(x[484]), .B(y[7948]), .Z(n25897) );
  XOR U27255 ( .A(n25896), .B(n25897), .Z(n25873) );
  XOR U27256 ( .A(n25875), .B(n25874), .Z(n25834) );
  NAND U27257 ( .A(n25769), .B(n25768), .Z(n25773) );
  NAND U27258 ( .A(n25771), .B(n25770), .Z(n25772) );
  NAND U27259 ( .A(n25773), .B(n25772), .Z(n25879) );
  NAND U27260 ( .A(n25775), .B(n25774), .Z(n25779) );
  NAND U27261 ( .A(n25777), .B(n25776), .Z(n25778) );
  AND U27262 ( .A(n25779), .B(n25778), .Z(n25910) );
  AND U27263 ( .A(x[493]), .B(y[7940]), .Z(n25906) );
  NAND U27264 ( .A(n25906), .B(n26423), .Z(n25783) );
  NAND U27265 ( .A(n25781), .B(n25780), .Z(n25782) );
  NAND U27266 ( .A(n25783), .B(n25782), .Z(n25893) );
  AND U27267 ( .A(y[7950]), .B(x[482]), .Z(n25785) );
  NAND U27268 ( .A(y[7943]), .B(x[489]), .Z(n25784) );
  XNOR U27269 ( .A(n25785), .B(n25784), .Z(n25900) );
  NAND U27270 ( .A(x[483]), .B(y[7949]), .Z(n25901) );
  XNOR U27271 ( .A(n25900), .B(n25901), .Z(n25891) );
  AND U27272 ( .A(x[492]), .B(y[7940]), .Z(n26548) );
  AND U27273 ( .A(y[7947]), .B(x[485]), .Z(n25787) );
  NAND U27274 ( .A(y[7939]), .B(x[493]), .Z(n25786) );
  XNOR U27275 ( .A(n25787), .B(n25786), .Z(n25847) );
  XOR U27276 ( .A(n26548), .B(n25847), .Z(n25890) );
  XOR U27277 ( .A(n25891), .B(n25890), .Z(n25892) );
  XNOR U27278 ( .A(n25893), .B(n25892), .Z(n25907) );
  NAND U27279 ( .A(n25789), .B(n25788), .Z(n25793) );
  NAND U27280 ( .A(n25791), .B(n25790), .Z(n25792) );
  AND U27281 ( .A(n25793), .B(n25792), .Z(n25908) );
  XOR U27282 ( .A(n25907), .B(n25908), .Z(n25909) );
  XNOR U27283 ( .A(n25881), .B(n25880), .Z(n25921) );
  NAND U27284 ( .A(n25795), .B(n25794), .Z(n25799) );
  NAND U27285 ( .A(n25797), .B(n25796), .Z(n25798) );
  AND U27286 ( .A(n25799), .B(n25798), .Z(n25920) );
  XOR U27287 ( .A(n25921), .B(n25920), .Z(n25923) );
  NANDN U27288 ( .A(n25801), .B(n25800), .Z(n25805) );
  NANDN U27289 ( .A(n25803), .B(n25802), .Z(n25804) );
  NAND U27290 ( .A(n25805), .B(n25804), .Z(n25830) );
  NAND U27291 ( .A(n25807), .B(n25806), .Z(n25811) );
  NANDN U27292 ( .A(n25809), .B(n25808), .Z(n25810) );
  NAND U27293 ( .A(n25811), .B(n25810), .Z(n25828) );
  NANDN U27294 ( .A(n25813), .B(n25812), .Z(n25817) );
  NAND U27295 ( .A(n25815), .B(n25814), .Z(n25816) );
  AND U27296 ( .A(n25817), .B(n25816), .Z(n25829) );
  XOR U27297 ( .A(n25828), .B(n25829), .Z(n25831) );
  XOR U27298 ( .A(n25830), .B(n25831), .Z(n25922) );
  XNOR U27299 ( .A(n25923), .B(n25922), .Z(n25916) );
  NAND U27300 ( .A(n25822), .B(n25821), .Z(n25826) );
  NANDN U27301 ( .A(n25824), .B(n25823), .Z(n25825) );
  NAND U27302 ( .A(n25826), .B(n25825), .Z(n25914) );
  IV U27303 ( .A(n25914), .Z(n25913) );
  XOR U27304 ( .A(n25915), .B(n25913), .Z(n25827) );
  XNOR U27305 ( .A(n25916), .B(n25827), .Z(N561) );
  NAND U27306 ( .A(n25829), .B(n25828), .Z(n25833) );
  NAND U27307 ( .A(n25831), .B(n25830), .Z(n25832) );
  NAND U27308 ( .A(n25833), .B(n25832), .Z(n26024) );
  NANDN U27309 ( .A(n25835), .B(n25834), .Z(n25839) );
  NANDN U27310 ( .A(n25837), .B(n25836), .Z(n25838) );
  AND U27311 ( .A(n25839), .B(n25838), .Z(n25936) );
  NAND U27312 ( .A(n25841), .B(n25840), .Z(n25845) );
  NAND U27313 ( .A(n25843), .B(n25842), .Z(n25844) );
  NAND U27314 ( .A(n25845), .B(n25844), .Z(n26012) );
  AND U27315 ( .A(x[493]), .B(y[7947]), .Z(n26808) );
  NAND U27316 ( .A(n26808), .B(n25846), .Z(n25849) );
  NAND U27317 ( .A(n25847), .B(n26548), .Z(n25848) );
  NAND U27318 ( .A(n25849), .B(n25848), .Z(n25966) );
  AND U27319 ( .A(y[7952]), .B(x[481]), .Z(n25851) );
  NAND U27320 ( .A(y[7944]), .B(x[489]), .Z(n25850) );
  XNOR U27321 ( .A(n25851), .B(n25850), .Z(n25987) );
  ANDN U27322 ( .B(o[272]), .A(n25852), .Z(n25986) );
  XOR U27323 ( .A(n25987), .B(n25986), .Z(n25964) );
  AND U27324 ( .A(y[7938]), .B(x[495]), .Z(n25854) );
  NAND U27325 ( .A(y[7941]), .B(x[492]), .Z(n25853) );
  XNOR U27326 ( .A(n25854), .B(n25853), .Z(n25939) );
  AND U27327 ( .A(x[494]), .B(y[7939]), .Z(n25940) );
  XOR U27328 ( .A(n25939), .B(n25940), .Z(n25963) );
  XOR U27329 ( .A(n25964), .B(n25963), .Z(n25965) );
  XOR U27330 ( .A(n25966), .B(n25965), .Z(n26010) );
  AND U27331 ( .A(x[487]), .B(y[7946]), .Z(n25994) );
  NANDN U27332 ( .A(n25855), .B(n25994), .Z(n25859) );
  NAND U27333 ( .A(n25857), .B(n25856), .Z(n25858) );
  NAND U27334 ( .A(n25859), .B(n25858), .Z(n25976) );
  NAND U27335 ( .A(x[488]), .B(y[7951]), .Z(n26708) );
  AND U27336 ( .A(x[481]), .B(y[7944]), .Z(n26060) );
  NANDN U27337 ( .A(n26708), .B(n26060), .Z(n25863) );
  NAND U27338 ( .A(n25861), .B(n25860), .Z(n25862) );
  NAND U27339 ( .A(n25863), .B(n25862), .Z(n25975) );
  XOR U27340 ( .A(n25976), .B(n25975), .Z(n25978) );
  NAND U27341 ( .A(n25865), .B(n25864), .Z(n25869) );
  NAND U27342 ( .A(n25867), .B(n25866), .Z(n25868) );
  NAND U27343 ( .A(n25869), .B(n25868), .Z(n25972) );
  AND U27344 ( .A(x[480]), .B(y[7953]), .Z(n25953) );
  AND U27345 ( .A(x[497]), .B(y[7936]), .Z(n25954) );
  XOR U27346 ( .A(n25953), .B(n25954), .Z(n25955) );
  NAND U27347 ( .A(x[496]), .B(y[7937]), .Z(n25950) );
  XNOR U27348 ( .A(o[273]), .B(n25950), .Z(n25956) );
  XOR U27349 ( .A(n25955), .B(n25956), .Z(n25969) );
  AND U27350 ( .A(y[7951]), .B(x[482]), .Z(n25871) );
  NAND U27351 ( .A(y[7943]), .B(x[490]), .Z(n25870) );
  XNOR U27352 ( .A(n25871), .B(n25870), .Z(n25989) );
  NAND U27353 ( .A(x[483]), .B(y[7950]), .Z(n25990) );
  XNOR U27354 ( .A(n25989), .B(n25990), .Z(n25970) );
  XOR U27355 ( .A(n25969), .B(n25970), .Z(n25971) );
  XOR U27356 ( .A(n25972), .B(n25971), .Z(n25977) );
  XOR U27357 ( .A(n25978), .B(n25977), .Z(n26009) );
  XOR U27358 ( .A(n26010), .B(n26009), .Z(n26011) );
  XNOR U27359 ( .A(n26012), .B(n26011), .Z(n25933) );
  NANDN U27360 ( .A(n25873), .B(n25872), .Z(n25877) );
  NANDN U27361 ( .A(n25875), .B(n25874), .Z(n25876) );
  AND U27362 ( .A(n25877), .B(n25876), .Z(n25934) );
  XOR U27363 ( .A(n25933), .B(n25934), .Z(n25935) );
  NANDN U27364 ( .A(n25879), .B(n25878), .Z(n25883) );
  NAND U27365 ( .A(n25881), .B(n25880), .Z(n25882) );
  AND U27366 ( .A(n25883), .B(n25882), .Z(n25930) );
  NAND U27367 ( .A(n25885), .B(n25884), .Z(n25889) );
  NAND U27368 ( .A(n25887), .B(n25886), .Z(n25888) );
  NAND U27369 ( .A(n25889), .B(n25888), .Z(n26006) );
  NAND U27370 ( .A(n25891), .B(n25890), .Z(n25895) );
  NAND U27371 ( .A(n25893), .B(n25892), .Z(n25894) );
  NAND U27372 ( .A(n25895), .B(n25894), .Z(n26004) );
  NAND U27373 ( .A(x[494]), .B(y[7941]), .Z(n26194) );
  NANDN U27374 ( .A(n26194), .B(n26423), .Z(n25899) );
  NANDN U27375 ( .A(n25897), .B(n25896), .Z(n25898) );
  AND U27376 ( .A(n25899), .B(n25898), .Z(n25998) );
  AND U27377 ( .A(x[489]), .B(y[7950]), .Z(n26789) );
  NANDN U27378 ( .A(n25988), .B(n26789), .Z(n25903) );
  NANDN U27379 ( .A(n25901), .B(n25900), .Z(n25902) );
  NAND U27380 ( .A(n25903), .B(n25902), .Z(n25997) );
  XNOR U27381 ( .A(n25998), .B(n25997), .Z(n25999) );
  AND U27382 ( .A(y[7948]), .B(x[485]), .Z(n26047) );
  NAND U27383 ( .A(y[7945]), .B(x[488]), .Z(n25904) );
  XNOR U27384 ( .A(n26047), .B(n25904), .Z(n25982) );
  XOR U27385 ( .A(n25994), .B(n25993), .Z(n25995) );
  NAND U27386 ( .A(y[7949]), .B(x[484]), .Z(n25905) );
  XNOR U27387 ( .A(n25906), .B(n25905), .Z(n25944) );
  NAND U27388 ( .A(x[491]), .B(y[7942]), .Z(n25945) );
  XOR U27389 ( .A(n25944), .B(n25945), .Z(n25996) );
  XOR U27390 ( .A(n25995), .B(n25996), .Z(n26000) );
  XNOR U27391 ( .A(n25999), .B(n26000), .Z(n26003) );
  XOR U27392 ( .A(n26004), .B(n26003), .Z(n26005) );
  XNOR U27393 ( .A(n26006), .B(n26005), .Z(n25928) );
  NAND U27394 ( .A(n25908), .B(n25907), .Z(n25912) );
  NANDN U27395 ( .A(n25910), .B(n25909), .Z(n25911) );
  NAND U27396 ( .A(n25912), .B(n25911), .Z(n25927) );
  XOR U27397 ( .A(n25928), .B(n25927), .Z(n25929) );
  XOR U27398 ( .A(n25930), .B(n25929), .Z(n26022) );
  XOR U27399 ( .A(n26024), .B(n26025), .Z(n26018) );
  OR U27400 ( .A(n25915), .B(n25913), .Z(n25919) );
  ANDN U27401 ( .B(n25915), .A(n25914), .Z(n25917) );
  OR U27402 ( .A(n25917), .B(n25916), .Z(n25918) );
  AND U27403 ( .A(n25919), .B(n25918), .Z(n26016) );
  NAND U27404 ( .A(n25921), .B(n25920), .Z(n25925) );
  NAND U27405 ( .A(n25923), .B(n25922), .Z(n25924) );
  AND U27406 ( .A(n25925), .B(n25924), .Z(n26017) );
  IV U27407 ( .A(n26017), .Z(n26015) );
  XOR U27408 ( .A(n26016), .B(n26015), .Z(n25926) );
  XNOR U27409 ( .A(n26018), .B(n25926), .Z(N562) );
  NAND U27410 ( .A(n25928), .B(n25927), .Z(n25932) );
  NANDN U27411 ( .A(n25930), .B(n25929), .Z(n25931) );
  AND U27412 ( .A(n25932), .B(n25931), .Z(n26123) );
  NAND U27413 ( .A(n25934), .B(n25933), .Z(n25938) );
  NANDN U27414 ( .A(n25936), .B(n25935), .Z(n25937) );
  AND U27415 ( .A(n25938), .B(n25937), .Z(n26121) );
  AND U27416 ( .A(x[495]), .B(y[7941]), .Z(n26155) );
  AND U27417 ( .A(x[492]), .B(y[7938]), .Z(n26254) );
  NAND U27418 ( .A(n26155), .B(n26254), .Z(n25942) );
  NAND U27419 ( .A(n25940), .B(n25939), .Z(n25941) );
  AND U27420 ( .A(n25942), .B(n25941), .Z(n26103) );
  NAND U27421 ( .A(n27200), .B(n25943), .Z(n25947) );
  NANDN U27422 ( .A(n25945), .B(n25944), .Z(n25946) );
  NAND U27423 ( .A(n25947), .B(n25946), .Z(n26094) );
  AND U27424 ( .A(y[7953]), .B(x[481]), .Z(n25949) );
  NAND U27425 ( .A(y[7944]), .B(x[490]), .Z(n25948) );
  XNOR U27426 ( .A(n25949), .B(n25948), .Z(n26062) );
  ANDN U27427 ( .B(o[273]), .A(n25950), .Z(n26061) );
  XOR U27428 ( .A(n26062), .B(n26061), .Z(n26093) );
  AND U27429 ( .A(y[7939]), .B(x[495]), .Z(n25952) );
  NAND U27430 ( .A(y[7945]), .B(x[489]), .Z(n25951) );
  XNOR U27431 ( .A(n25952), .B(n25951), .Z(n26053) );
  AND U27432 ( .A(x[494]), .B(y[7940]), .Z(n26052) );
  XOR U27433 ( .A(n26053), .B(n26052), .Z(n26092) );
  XOR U27434 ( .A(n26093), .B(n26092), .Z(n26095) );
  XOR U27435 ( .A(n26094), .B(n26095), .Z(n26102) );
  NAND U27436 ( .A(n25954), .B(n25953), .Z(n25958) );
  NAND U27437 ( .A(n25956), .B(n25955), .Z(n25957) );
  AND U27438 ( .A(n25958), .B(n25957), .Z(n26115) );
  AND U27439 ( .A(y[7938]), .B(x[496]), .Z(n25960) );
  NAND U27440 ( .A(y[7943]), .B(x[491]), .Z(n25959) );
  XNOR U27441 ( .A(n25960), .B(n25959), .Z(n26051) );
  AND U27442 ( .A(x[482]), .B(y[7952]), .Z(n26050) );
  XOR U27443 ( .A(n26051), .B(n26050), .Z(n26114) );
  AND U27444 ( .A(y[7949]), .B(x[485]), .Z(n26176) );
  NAND U27445 ( .A(y[7948]), .B(x[486]), .Z(n25961) );
  XNOR U27446 ( .A(n26176), .B(n25961), .Z(n26049) );
  NAND U27447 ( .A(y[7950]), .B(x[484]), .Z(n25962) );
  XNOR U27448 ( .A(n26794), .B(n25962), .Z(n26082) );
  AND U27449 ( .A(x[487]), .B(y[7947]), .Z(n26081) );
  XOR U27450 ( .A(n26082), .B(n26081), .Z(n26048) );
  XOR U27451 ( .A(n26049), .B(n26048), .Z(n26116) );
  XOR U27452 ( .A(n26117), .B(n26116), .Z(n26104) );
  XNOR U27453 ( .A(n26105), .B(n26104), .Z(n26036) );
  NAND U27454 ( .A(n25964), .B(n25963), .Z(n25968) );
  NAND U27455 ( .A(n25966), .B(n25965), .Z(n25967) );
  AND U27456 ( .A(n25968), .B(n25967), .Z(n26096) );
  NAND U27457 ( .A(n25970), .B(n25969), .Z(n25974) );
  NAND U27458 ( .A(n25972), .B(n25971), .Z(n25973) );
  NAND U27459 ( .A(n25974), .B(n25973), .Z(n26097) );
  NAND U27460 ( .A(n25976), .B(n25975), .Z(n25980) );
  NAND U27461 ( .A(n25978), .B(n25977), .Z(n25979) );
  NAND U27462 ( .A(n25980), .B(n25979), .Z(n26099) );
  XOR U27463 ( .A(n26036), .B(n26035), .Z(n26038) );
  AND U27464 ( .A(x[488]), .B(y[7948]), .Z(n26294) );
  NAND U27465 ( .A(n26294), .B(n25981), .Z(n25985) );
  NANDN U27466 ( .A(n25983), .B(n25982), .Z(n25984) );
  AND U27467 ( .A(n25985), .B(n25984), .Z(n26109) );
  NAND U27468 ( .A(x[489]), .B(y[7952]), .Z(n26937) );
  NAND U27469 ( .A(x[490]), .B(y[7951]), .Z(n26936) );
  AND U27470 ( .A(x[480]), .B(y[7954]), .Z(n26063) );
  NAND U27471 ( .A(x[498]), .B(y[7936]), .Z(n26064) );
  XNOR U27472 ( .A(n26063), .B(n26064), .Z(n26065) );
  NAND U27473 ( .A(x[497]), .B(y[7937]), .Z(n26085) );
  XOR U27474 ( .A(o[274]), .B(n26085), .Z(n26066) );
  XNOR U27475 ( .A(n26065), .B(n26066), .Z(n26089) );
  AND U27476 ( .A(y[7941]), .B(x[493]), .Z(n25992) );
  NAND U27477 ( .A(y[7951]), .B(x[483]), .Z(n25991) );
  XNOR U27478 ( .A(n25992), .B(n25991), .Z(n26072) );
  AND U27479 ( .A(x[492]), .B(y[7942]), .Z(n26071) );
  XOR U27480 ( .A(n26072), .B(n26071), .Z(n26088) );
  XOR U27481 ( .A(n26089), .B(n26088), .Z(n26091) );
  XOR U27482 ( .A(n26090), .B(n26091), .Z(n26110) );
  XOR U27483 ( .A(n26111), .B(n26110), .Z(n26042) );
  XNOR U27484 ( .A(n26042), .B(n26041), .Z(n26043) );
  NANDN U27485 ( .A(n25998), .B(n25997), .Z(n26002) );
  NANDN U27486 ( .A(n26000), .B(n25999), .Z(n26001) );
  NAND U27487 ( .A(n26002), .B(n26001), .Z(n26044) );
  XNOR U27488 ( .A(n26043), .B(n26044), .Z(n26037) );
  XNOR U27489 ( .A(n26038), .B(n26037), .Z(n26032) );
  NAND U27490 ( .A(n26004), .B(n26003), .Z(n26008) );
  NAND U27491 ( .A(n26006), .B(n26005), .Z(n26007) );
  NAND U27492 ( .A(n26008), .B(n26007), .Z(n26030) );
  NAND U27493 ( .A(n26010), .B(n26009), .Z(n26014) );
  NAND U27494 ( .A(n26012), .B(n26011), .Z(n26013) );
  NAND U27495 ( .A(n26014), .B(n26013), .Z(n26029) );
  XOR U27496 ( .A(n26030), .B(n26029), .Z(n26031) );
  XOR U27497 ( .A(n26032), .B(n26031), .Z(n26120) );
  XOR U27498 ( .A(n26121), .B(n26120), .Z(n26122) );
  XNOR U27499 ( .A(n26123), .B(n26122), .Z(n26128) );
  NANDN U27500 ( .A(n26015), .B(n26016), .Z(n26021) );
  NOR U27501 ( .A(n26017), .B(n26016), .Z(n26019) );
  OR U27502 ( .A(n26019), .B(n26018), .Z(n26020) );
  AND U27503 ( .A(n26021), .B(n26020), .Z(n26127) );
  NANDN U27504 ( .A(n26023), .B(n26022), .Z(n26027) );
  NAND U27505 ( .A(n26025), .B(n26024), .Z(n26026) );
  NAND U27506 ( .A(n26027), .B(n26026), .Z(n26126) );
  XOR U27507 ( .A(n26127), .B(n26126), .Z(n26028) );
  XNOR U27508 ( .A(n26128), .B(n26028), .Z(N563) );
  NAND U27509 ( .A(n26030), .B(n26029), .Z(n26034) );
  NAND U27510 ( .A(n26032), .B(n26031), .Z(n26033) );
  AND U27511 ( .A(n26034), .B(n26033), .Z(n26238) );
  NAND U27512 ( .A(n26036), .B(n26035), .Z(n26040) );
  NAND U27513 ( .A(n26038), .B(n26037), .Z(n26039) );
  AND U27514 ( .A(n26040), .B(n26039), .Z(n26236) );
  NANDN U27515 ( .A(n26042), .B(n26041), .Z(n26046) );
  NANDN U27516 ( .A(n26044), .B(n26043), .Z(n26045) );
  NAND U27517 ( .A(n26046), .B(n26045), .Z(n26219) );
  AND U27518 ( .A(x[496]), .B(y[7943]), .Z(n26564) );
  AND U27519 ( .A(x[495]), .B(y[7945]), .Z(n26821) );
  NAND U27520 ( .A(n26821), .B(n26142), .Z(n26055) );
  NAND U27521 ( .A(n26053), .B(n26052), .Z(n26054) );
  NAND U27522 ( .A(n26055), .B(n26054), .Z(n26133) );
  AND U27523 ( .A(y[7954]), .B(x[481]), .Z(n26057) );
  NAND U27524 ( .A(y[7947]), .B(x[488]), .Z(n26056) );
  XNOR U27525 ( .A(n26057), .B(n26056), .Z(n26193) );
  AND U27526 ( .A(y[7942]), .B(x[493]), .Z(n26059) );
  NAND U27527 ( .A(y[7953]), .B(x[482]), .Z(n26058) );
  XNOR U27528 ( .A(n26059), .B(n26058), .Z(n26148) );
  XOR U27529 ( .A(n26131), .B(n26130), .Z(n26132) );
  XOR U27530 ( .A(n26133), .B(n26132), .Z(n26213) );
  XOR U27531 ( .A(n26212), .B(n26213), .Z(n26215) );
  XOR U27532 ( .A(n26214), .B(n26215), .Z(n26217) );
  AND U27533 ( .A(x[490]), .B(y[7953]), .Z(n27280) );
  IV U27534 ( .A(n27280), .Z(n27153) );
  NANDN U27535 ( .A(n26064), .B(n26063), .Z(n26068) );
  NANDN U27536 ( .A(n26066), .B(n26065), .Z(n26067) );
  NAND U27537 ( .A(n26068), .B(n26067), .Z(n26171) );
  AND U27538 ( .A(y[7939]), .B(x[496]), .Z(n26872) );
  NAND U27539 ( .A(y[7946]), .B(x[489]), .Z(n26069) );
  XNOR U27540 ( .A(n26872), .B(n26069), .Z(n26143) );
  AND U27541 ( .A(x[495]), .B(y[7940]), .Z(n26144) );
  XOR U27542 ( .A(n26143), .B(n26144), .Z(n26170) );
  XOR U27543 ( .A(n26171), .B(n26170), .Z(n26172) );
  XOR U27544 ( .A(n26173), .B(n26172), .Z(n26209) );
  AND U27545 ( .A(x[493]), .B(y[7951]), .Z(n27485) );
  NANDN U27546 ( .A(n26070), .B(n27485), .Z(n26074) );
  NAND U27547 ( .A(n26072), .B(n26071), .Z(n26073) );
  NAND U27548 ( .A(n26074), .B(n26073), .Z(n26167) );
  AND U27549 ( .A(y[7945]), .B(x[490]), .Z(n26076) );
  NAND U27550 ( .A(y[7938]), .B(x[497]), .Z(n26075) );
  XNOR U27551 ( .A(n26076), .B(n26075), .Z(n26199) );
  AND U27552 ( .A(x[498]), .B(y[7937]), .Z(n26163) );
  XOR U27553 ( .A(o[275]), .B(n26163), .Z(n26198) );
  XOR U27554 ( .A(n26199), .B(n26198), .Z(n26165) );
  NAND U27555 ( .A(y[7952]), .B(x[483]), .Z(n26077) );
  XNOR U27556 ( .A(n26078), .B(n26077), .Z(n26157) );
  XOR U27557 ( .A(n26165), .B(n26164), .Z(n26166) );
  XOR U27558 ( .A(n26167), .B(n26166), .Z(n26207) );
  NAND U27559 ( .A(n26080), .B(n26079), .Z(n26084) );
  NAND U27560 ( .A(n26082), .B(n26081), .Z(n26083) );
  AND U27561 ( .A(n26084), .B(n26083), .Z(n26139) );
  AND U27562 ( .A(x[480]), .B(y[7955]), .Z(n26180) );
  AND U27563 ( .A(x[499]), .B(y[7936]), .Z(n26181) );
  XOR U27564 ( .A(n26180), .B(n26181), .Z(n26183) );
  ANDN U27565 ( .B(o[274]), .A(n26085), .Z(n26182) );
  XOR U27566 ( .A(n26183), .B(n26182), .Z(n26137) );
  AND U27567 ( .A(x[484]), .B(y[7951]), .Z(n26308) );
  AND U27568 ( .A(y[7950]), .B(x[485]), .Z(n26087) );
  NAND U27569 ( .A(y[7949]), .B(x[486]), .Z(n26086) );
  XNOR U27570 ( .A(n26087), .B(n26086), .Z(n26177) );
  XOR U27571 ( .A(n26308), .B(n26177), .Z(n26136) );
  XOR U27572 ( .A(n26137), .B(n26136), .Z(n26138) );
  XOR U27573 ( .A(n26139), .B(n26138), .Z(n26206) );
  XNOR U27574 ( .A(n26207), .B(n26206), .Z(n26208) );
  XOR U27575 ( .A(n26209), .B(n26208), .Z(n26204) );
  XOR U27576 ( .A(n26202), .B(n26203), .Z(n26205) );
  XOR U27577 ( .A(n26204), .B(n26205), .Z(n26216) );
  XOR U27578 ( .A(n26217), .B(n26216), .Z(n26218) );
  XNOR U27579 ( .A(n26219), .B(n26218), .Z(n26228) );
  NANDN U27580 ( .A(n26097), .B(n26096), .Z(n26101) );
  NANDN U27581 ( .A(n26099), .B(n26098), .Z(n26100) );
  AND U27582 ( .A(n26101), .B(n26100), .Z(n26227) );
  NANDN U27583 ( .A(n26103), .B(n26102), .Z(n26107) );
  NAND U27584 ( .A(n26105), .B(n26104), .Z(n26106) );
  AND U27585 ( .A(n26107), .B(n26106), .Z(n26223) );
  NANDN U27586 ( .A(n26109), .B(n26108), .Z(n26113) );
  NAND U27587 ( .A(n26111), .B(n26110), .Z(n26112) );
  AND U27588 ( .A(n26113), .B(n26112), .Z(n26221) );
  NANDN U27589 ( .A(n26115), .B(n26114), .Z(n26119) );
  NAND U27590 ( .A(n26117), .B(n26116), .Z(n26118) );
  NAND U27591 ( .A(n26119), .B(n26118), .Z(n26220) );
  XOR U27592 ( .A(n26227), .B(n26226), .Z(n26229) );
  XOR U27593 ( .A(n26228), .B(n26229), .Z(n26235) );
  XOR U27594 ( .A(n26236), .B(n26235), .Z(n26237) );
  XOR U27595 ( .A(n26238), .B(n26237), .Z(n26234) );
  NAND U27596 ( .A(n26121), .B(n26120), .Z(n26125) );
  NAND U27597 ( .A(n26123), .B(n26122), .Z(n26124) );
  NAND U27598 ( .A(n26125), .B(n26124), .Z(n26232) );
  XOR U27599 ( .A(n26232), .B(n26233), .Z(n26129) );
  XNOR U27600 ( .A(n26234), .B(n26129), .Z(N564) );
  NAND U27601 ( .A(n26131), .B(n26130), .Z(n26135) );
  NAND U27602 ( .A(n26133), .B(n26132), .Z(n26134) );
  NAND U27603 ( .A(n26135), .B(n26134), .Z(n26243) );
  NAND U27604 ( .A(n26137), .B(n26136), .Z(n26141) );
  NANDN U27605 ( .A(n26139), .B(n26138), .Z(n26140) );
  NAND U27606 ( .A(n26141), .B(n26140), .Z(n26242) );
  XOR U27607 ( .A(n26243), .B(n26242), .Z(n26245) );
  AND U27608 ( .A(x[496]), .B(y[7946]), .Z(n27112) );
  NAND U27609 ( .A(n27112), .B(n26142), .Z(n26146) );
  NAND U27610 ( .A(n26144), .B(n26143), .Z(n26145) );
  NAND U27611 ( .A(n26146), .B(n26145), .Z(n26283) );
  AND U27612 ( .A(x[493]), .B(y[7953]), .Z(n27725) );
  NAND U27613 ( .A(n27725), .B(n26147), .Z(n26151) );
  NANDN U27614 ( .A(n26149), .B(n26148), .Z(n26150) );
  NAND U27615 ( .A(n26151), .B(n26150), .Z(n26328) );
  AND U27616 ( .A(y[7940]), .B(x[496]), .Z(n26153) );
  NAND U27617 ( .A(y[7946]), .B(x[490]), .Z(n26152) );
  XNOR U27618 ( .A(n26153), .B(n26152), .Z(n26289) );
  AND U27619 ( .A(x[482]), .B(y[7954]), .Z(n26290) );
  XOR U27620 ( .A(n26289), .B(n26290), .Z(n26326) );
  NAND U27621 ( .A(y[7947]), .B(x[489]), .Z(n26154) );
  XNOR U27622 ( .A(n26155), .B(n26154), .Z(n26265) );
  AND U27623 ( .A(x[494]), .B(y[7942]), .Z(n26266) );
  XOR U27624 ( .A(n26265), .B(n26266), .Z(n26325) );
  XOR U27625 ( .A(n26326), .B(n26325), .Z(n26327) );
  XOR U27626 ( .A(n26328), .B(n26327), .Z(n26282) );
  XOR U27627 ( .A(n26283), .B(n26282), .Z(n26285) );
  NAND U27628 ( .A(x[491]), .B(y[7952]), .Z(n27281) );
  NANDN U27629 ( .A(n27281), .B(n26156), .Z(n26160) );
  NANDN U27630 ( .A(n26158), .B(n26157), .Z(n26159) );
  NAND U27631 ( .A(n26160), .B(n26159), .Z(n26334) );
  AND U27632 ( .A(y[7945]), .B(x[491]), .Z(n26162) );
  NAND U27633 ( .A(y[7955]), .B(x[481]), .Z(n26161) );
  XNOR U27634 ( .A(n26162), .B(n26161), .Z(n26261) );
  AND U27635 ( .A(x[499]), .B(y[7937]), .Z(n26269) );
  XOR U27636 ( .A(o[276]), .B(n26269), .Z(n26260) );
  XOR U27637 ( .A(n26261), .B(n26260), .Z(n26332) );
  AND U27638 ( .A(x[480]), .B(y[7956]), .Z(n26313) );
  AND U27639 ( .A(x[500]), .B(y[7936]), .Z(n26314) );
  XOR U27640 ( .A(n26313), .B(n26314), .Z(n26316) );
  AND U27641 ( .A(o[275]), .B(n26163), .Z(n26315) );
  XOR U27642 ( .A(n26316), .B(n26315), .Z(n26331) );
  XOR U27643 ( .A(n26332), .B(n26331), .Z(n26333) );
  XOR U27644 ( .A(n26334), .B(n26333), .Z(n26284) );
  XOR U27645 ( .A(n26285), .B(n26284), .Z(n26244) );
  XNOR U27646 ( .A(n26245), .B(n26244), .Z(n26340) );
  NAND U27647 ( .A(n26165), .B(n26164), .Z(n26169) );
  NAND U27648 ( .A(n26167), .B(n26166), .Z(n26168) );
  AND U27649 ( .A(n26169), .B(n26168), .Z(n26338) );
  NAND U27650 ( .A(n26171), .B(n26170), .Z(n26175) );
  NAND U27651 ( .A(n26173), .B(n26172), .Z(n26174) );
  AND U27652 ( .A(n26175), .B(n26174), .Z(n26279) );
  NAND U27653 ( .A(x[486]), .B(y[7950]), .Z(n26249) );
  NANDN U27654 ( .A(n26249), .B(n26176), .Z(n26179) );
  NAND U27655 ( .A(n26177), .B(n26308), .Z(n26178) );
  NAND U27656 ( .A(n26179), .B(n26178), .Z(n26273) );
  NAND U27657 ( .A(n26181), .B(n26180), .Z(n26185) );
  NAND U27658 ( .A(n26183), .B(n26182), .Z(n26184) );
  NAND U27659 ( .A(n26185), .B(n26184), .Z(n26271) );
  AND U27660 ( .A(y[7938]), .B(x[498]), .Z(n26187) );
  NAND U27661 ( .A(y[7944]), .B(x[492]), .Z(n26186) );
  XNOR U27662 ( .A(n26187), .B(n26186), .Z(n26255) );
  AND U27663 ( .A(x[497]), .B(y[7939]), .Z(n26256) );
  XOR U27664 ( .A(n26255), .B(n26256), .Z(n26270) );
  XOR U27665 ( .A(n26271), .B(n26270), .Z(n26272) );
  XNOR U27666 ( .A(n26273), .B(n26272), .Z(n26277) );
  AND U27667 ( .A(y[7943]), .B(x[493]), .Z(n26189) );
  NAND U27668 ( .A(y[7953]), .B(x[483]), .Z(n26188) );
  XNOR U27669 ( .A(n26189), .B(n26188), .Z(n26295) );
  XNOR U27670 ( .A(n26295), .B(n26294), .Z(n26251) );
  AND U27671 ( .A(y[7951]), .B(x[485]), .Z(n26191) );
  NAND U27672 ( .A(y[7952]), .B(x[484]), .Z(n26190) );
  XNOR U27673 ( .A(n26191), .B(n26190), .Z(n26310) );
  AND U27674 ( .A(x[487]), .B(y[7949]), .Z(n26309) );
  XNOR U27675 ( .A(n26310), .B(n26309), .Z(n26248) );
  XOR U27676 ( .A(n26249), .B(n26248), .Z(n26250) );
  XNOR U27677 ( .A(n26251), .B(n26250), .Z(n26321) );
  AND U27678 ( .A(x[488]), .B(y[7954]), .Z(n27437) );
  AND U27679 ( .A(x[481]), .B(y[7947]), .Z(n26192) );
  NAND U27680 ( .A(n27437), .B(n26192), .Z(n26196) );
  NANDN U27681 ( .A(n26194), .B(n26193), .Z(n26195) );
  NAND U27682 ( .A(n26196), .B(n26195), .Z(n26320) );
  NAND U27683 ( .A(x[497]), .B(y[7945]), .Z(n27120) );
  NANDN U27684 ( .A(n27120), .B(n26197), .Z(n26201) );
  NAND U27685 ( .A(n26199), .B(n26198), .Z(n26200) );
  NAND U27686 ( .A(n26201), .B(n26200), .Z(n26319) );
  XOR U27687 ( .A(n26320), .B(n26319), .Z(n26322) );
  XNOR U27688 ( .A(n26321), .B(n26322), .Z(n26276) );
  XOR U27689 ( .A(n26277), .B(n26276), .Z(n26278) );
  XOR U27690 ( .A(n26279), .B(n26278), .Z(n26337) );
  XOR U27691 ( .A(n26338), .B(n26337), .Z(n26339) );
  XOR U27692 ( .A(n26340), .B(n26339), .Z(n26344) );
  NANDN U27693 ( .A(n26207), .B(n26206), .Z(n26211) );
  NANDN U27694 ( .A(n26209), .B(n26208), .Z(n26210) );
  AND U27695 ( .A(n26211), .B(n26210), .Z(n26350) );
  XNOR U27696 ( .A(n26350), .B(n26349), .Z(n26351) );
  XNOR U27697 ( .A(n26352), .B(n26351), .Z(n26343) );
  XNOR U27698 ( .A(n26344), .B(n26343), .Z(n26346) );
  XOR U27699 ( .A(n26346), .B(n26345), .Z(n26358) );
  NANDN U27700 ( .A(n26221), .B(n26220), .Z(n26225) );
  NANDN U27701 ( .A(n26223), .B(n26222), .Z(n26224) );
  AND U27702 ( .A(n26225), .B(n26224), .Z(n26355) );
  NAND U27703 ( .A(n26227), .B(n26226), .Z(n26231) );
  NAND U27704 ( .A(n26229), .B(n26228), .Z(n26230) );
  NAND U27705 ( .A(n26231), .B(n26230), .Z(n26356) );
  XOR U27706 ( .A(n26358), .B(n26357), .Z(n26364) );
  NAND U27707 ( .A(n26236), .B(n26235), .Z(n26240) );
  NANDN U27708 ( .A(n26238), .B(n26237), .Z(n26239) );
  AND U27709 ( .A(n26240), .B(n26239), .Z(n26363) );
  IV U27710 ( .A(n26363), .Z(n26361) );
  XOR U27711 ( .A(n26362), .B(n26361), .Z(n26241) );
  XNOR U27712 ( .A(n26364), .B(n26241), .Z(N565) );
  NAND U27713 ( .A(n26243), .B(n26242), .Z(n26247) );
  NAND U27714 ( .A(n26245), .B(n26244), .Z(n26246) );
  NAND U27715 ( .A(n26247), .B(n26246), .Z(n26378) );
  NAND U27716 ( .A(n26249), .B(n26248), .Z(n26253) );
  NAND U27717 ( .A(n26251), .B(n26250), .Z(n26252) );
  NAND U27718 ( .A(n26253), .B(n26252), .Z(n26400) );
  AND U27719 ( .A(x[498]), .B(y[7944]), .Z(n27118) );
  NAND U27720 ( .A(n27118), .B(n26254), .Z(n26258) );
  NAND U27721 ( .A(n26256), .B(n26255), .Z(n26257) );
  NAND U27722 ( .A(n26258), .B(n26257), .Z(n26382) );
  AND U27723 ( .A(x[491]), .B(y[7955]), .Z(n27866) );
  AND U27724 ( .A(x[481]), .B(y[7945]), .Z(n26259) );
  NAND U27725 ( .A(n27866), .B(n26259), .Z(n26263) );
  NAND U27726 ( .A(n26261), .B(n26260), .Z(n26262) );
  NAND U27727 ( .A(n26263), .B(n26262), .Z(n26381) );
  XOR U27728 ( .A(n26382), .B(n26381), .Z(n26384) );
  AND U27729 ( .A(x[495]), .B(y[7947]), .Z(n27106) );
  NAND U27730 ( .A(n27106), .B(n26264), .Z(n26268) );
  NAND U27731 ( .A(n26266), .B(n26265), .Z(n26267) );
  NAND U27732 ( .A(n26268), .B(n26267), .Z(n26437) );
  AND U27733 ( .A(o[276]), .B(n26269), .Z(n26459) );
  AND U27734 ( .A(x[480]), .B(y[7957]), .Z(n26456) );
  AND U27735 ( .A(x[501]), .B(y[7936]), .Z(n26457) );
  XOR U27736 ( .A(n26456), .B(n26457), .Z(n26458) );
  XOR U27737 ( .A(n26459), .B(n26458), .Z(n26435) );
  AND U27738 ( .A(x[485]), .B(y[7952]), .Z(n26443) );
  AND U27739 ( .A(x[496]), .B(y[7941]), .Z(n26442) );
  XOR U27740 ( .A(n26443), .B(n26442), .Z(n26441) );
  AND U27741 ( .A(x[495]), .B(y[7942]), .Z(n26440) );
  XOR U27742 ( .A(n26441), .B(n26440), .Z(n26434) );
  XOR U27743 ( .A(n26435), .B(n26434), .Z(n26436) );
  XOR U27744 ( .A(n26437), .B(n26436), .Z(n26383) );
  XNOR U27745 ( .A(n26384), .B(n26383), .Z(n26399) );
  XOR U27746 ( .A(n26400), .B(n26399), .Z(n26402) );
  NAND U27747 ( .A(n26271), .B(n26270), .Z(n26275) );
  NAND U27748 ( .A(n26273), .B(n26272), .Z(n26274) );
  AND U27749 ( .A(n26275), .B(n26274), .Z(n26401) );
  XNOR U27750 ( .A(n26402), .B(n26401), .Z(n26376) );
  NAND U27751 ( .A(n26277), .B(n26276), .Z(n26281) );
  NAND U27752 ( .A(n26279), .B(n26278), .Z(n26280) );
  AND U27753 ( .A(n26281), .B(n26280), .Z(n26375) );
  XOR U27754 ( .A(n26376), .B(n26375), .Z(n26377) );
  XNOR U27755 ( .A(n26378), .B(n26377), .Z(n26371) );
  NAND U27756 ( .A(n26283), .B(n26282), .Z(n26287) );
  NAND U27757 ( .A(n26285), .B(n26284), .Z(n26286) );
  NAND U27758 ( .A(n26287), .B(n26286), .Z(n26475) );
  NAND U27759 ( .A(n27112), .B(n26288), .Z(n26292) );
  NAND U27760 ( .A(n26290), .B(n26289), .Z(n26291) );
  NAND U27761 ( .A(n26292), .B(n26291), .Z(n26406) );
  NAND U27762 ( .A(n27725), .B(n26293), .Z(n26297) );
  NAND U27763 ( .A(n26295), .B(n26294), .Z(n26296) );
  NAND U27764 ( .A(n26297), .B(n26296), .Z(n26396) );
  AND U27765 ( .A(y[7938]), .B(x[499]), .Z(n26299) );
  NAND U27766 ( .A(y[7946]), .B(x[491]), .Z(n26298) );
  XNOR U27767 ( .A(n26299), .B(n26298), .Z(n26425) );
  AND U27768 ( .A(x[500]), .B(y[7937]), .Z(n26455) );
  XOR U27769 ( .A(o[277]), .B(n26455), .Z(n26424) );
  XOR U27770 ( .A(n26425), .B(n26424), .Z(n26394) );
  AND U27771 ( .A(y[7939]), .B(x[498]), .Z(n26301) );
  NAND U27772 ( .A(y[7947]), .B(x[490]), .Z(n26300) );
  XNOR U27773 ( .A(n26301), .B(n26300), .Z(n26463) );
  AND U27774 ( .A(x[481]), .B(y[7956]), .Z(n26464) );
  XOR U27775 ( .A(n26463), .B(n26464), .Z(n26393) );
  XOR U27776 ( .A(n26394), .B(n26393), .Z(n26395) );
  XOR U27777 ( .A(n26396), .B(n26395), .Z(n26405) );
  XOR U27778 ( .A(n26406), .B(n26405), .Z(n26408) );
  AND U27779 ( .A(x[487]), .B(y[7950]), .Z(n26706) );
  AND U27780 ( .A(y[7951]), .B(x[486]), .Z(n26303) );
  NAND U27781 ( .A(y[7943]), .B(x[494]), .Z(n26302) );
  XNOR U27782 ( .A(n26303), .B(n26302), .Z(n26467) );
  XNOR U27783 ( .A(n26706), .B(n26467), .Z(n26414) );
  NAND U27784 ( .A(x[489]), .B(y[7948]), .Z(n26412) );
  NAND U27785 ( .A(x[488]), .B(y[7949]), .Z(n26411) );
  XOR U27786 ( .A(n26412), .B(n26411), .Z(n26413) );
  XNOR U27787 ( .A(n26414), .B(n26413), .Z(n26430) );
  AND U27788 ( .A(y[7945]), .B(x[492]), .Z(n26305) );
  NAND U27789 ( .A(y[7940]), .B(x[497]), .Z(n26304) );
  XNOR U27790 ( .A(n26305), .B(n26304), .Z(n26417) );
  AND U27791 ( .A(x[482]), .B(y[7955]), .Z(n26418) );
  XOR U27792 ( .A(n26417), .B(n26418), .Z(n26429) );
  AND U27793 ( .A(y[7944]), .B(x[493]), .Z(n26307) );
  NAND U27794 ( .A(y[7954]), .B(x[483]), .Z(n26306) );
  XNOR U27795 ( .A(n26307), .B(n26306), .Z(n26451) );
  AND U27796 ( .A(x[484]), .B(y[7953]), .Z(n26452) );
  XOR U27797 ( .A(n26451), .B(n26452), .Z(n26428) );
  XOR U27798 ( .A(n26429), .B(n26428), .Z(n26431) );
  XOR U27799 ( .A(n26430), .B(n26431), .Z(n26390) );
  NAND U27800 ( .A(n26443), .B(n26308), .Z(n26312) );
  NAND U27801 ( .A(n26310), .B(n26309), .Z(n26311) );
  NAND U27802 ( .A(n26312), .B(n26311), .Z(n26388) );
  NAND U27803 ( .A(n26314), .B(n26313), .Z(n26318) );
  NAND U27804 ( .A(n26316), .B(n26315), .Z(n26317) );
  NAND U27805 ( .A(n26318), .B(n26317), .Z(n26387) );
  XOR U27806 ( .A(n26388), .B(n26387), .Z(n26389) );
  XOR U27807 ( .A(n26390), .B(n26389), .Z(n26407) );
  XOR U27808 ( .A(n26408), .B(n26407), .Z(n26473) );
  NAND U27809 ( .A(n26320), .B(n26319), .Z(n26324) );
  NAND U27810 ( .A(n26322), .B(n26321), .Z(n26323) );
  NAND U27811 ( .A(n26324), .B(n26323), .Z(n26480) );
  NAND U27812 ( .A(n26326), .B(n26325), .Z(n26330) );
  NAND U27813 ( .A(n26328), .B(n26327), .Z(n26329) );
  NAND U27814 ( .A(n26330), .B(n26329), .Z(n26479) );
  NAND U27815 ( .A(n26332), .B(n26331), .Z(n26336) );
  NAND U27816 ( .A(n26334), .B(n26333), .Z(n26335) );
  NAND U27817 ( .A(n26336), .B(n26335), .Z(n26478) );
  XOR U27818 ( .A(n26479), .B(n26478), .Z(n26481) );
  XOR U27819 ( .A(n26480), .B(n26481), .Z(n26472) );
  XOR U27820 ( .A(n26473), .B(n26472), .Z(n26474) );
  XNOR U27821 ( .A(n26475), .B(n26474), .Z(n26370) );
  NAND U27822 ( .A(n26338), .B(n26337), .Z(n26342) );
  NAND U27823 ( .A(n26340), .B(n26339), .Z(n26341) );
  NAND U27824 ( .A(n26342), .B(n26341), .Z(n26369) );
  XOR U27825 ( .A(n26370), .B(n26369), .Z(n26372) );
  XOR U27826 ( .A(n26371), .B(n26372), .Z(n26487) );
  NANDN U27827 ( .A(n26344), .B(n26343), .Z(n26348) );
  NAND U27828 ( .A(n26346), .B(n26345), .Z(n26347) );
  NAND U27829 ( .A(n26348), .B(n26347), .Z(n26484) );
  NANDN U27830 ( .A(n26350), .B(n26349), .Z(n26354) );
  NAND U27831 ( .A(n26352), .B(n26351), .Z(n26353) );
  AND U27832 ( .A(n26354), .B(n26353), .Z(n26485) );
  XOR U27833 ( .A(n26484), .B(n26485), .Z(n26486) );
  XNOR U27834 ( .A(n26487), .B(n26486), .Z(n26490) );
  NANDN U27835 ( .A(n26356), .B(n26355), .Z(n26360) );
  NANDN U27836 ( .A(n26358), .B(n26357), .Z(n26359) );
  NAND U27837 ( .A(n26360), .B(n26359), .Z(n26488) );
  NANDN U27838 ( .A(n26361), .B(n26362), .Z(n26367) );
  NOR U27839 ( .A(n26363), .B(n26362), .Z(n26365) );
  OR U27840 ( .A(n26365), .B(n26364), .Z(n26366) );
  AND U27841 ( .A(n26367), .B(n26366), .Z(n26489) );
  XOR U27842 ( .A(n26488), .B(n26489), .Z(n26368) );
  XNOR U27843 ( .A(n26490), .B(n26368), .Z(N566) );
  NAND U27844 ( .A(n26370), .B(n26369), .Z(n26374) );
  NAND U27845 ( .A(n26372), .B(n26371), .Z(n26373) );
  AND U27846 ( .A(n26374), .B(n26373), .Z(n26622) );
  NAND U27847 ( .A(n26376), .B(n26375), .Z(n26380) );
  NAND U27848 ( .A(n26378), .B(n26377), .Z(n26379) );
  NAND U27849 ( .A(n26380), .B(n26379), .Z(n26620) );
  NAND U27850 ( .A(n26382), .B(n26381), .Z(n26386) );
  NAND U27851 ( .A(n26384), .B(n26383), .Z(n26385) );
  NAND U27852 ( .A(n26386), .B(n26385), .Z(n26501) );
  NAND U27853 ( .A(n26388), .B(n26387), .Z(n26392) );
  NAND U27854 ( .A(n26390), .B(n26389), .Z(n26391) );
  NAND U27855 ( .A(n26392), .B(n26391), .Z(n26499) );
  NAND U27856 ( .A(n26394), .B(n26393), .Z(n26398) );
  NAND U27857 ( .A(n26396), .B(n26395), .Z(n26397) );
  NAND U27858 ( .A(n26398), .B(n26397), .Z(n26498) );
  XOR U27859 ( .A(n26499), .B(n26498), .Z(n26500) );
  XOR U27860 ( .A(n26501), .B(n26500), .Z(n26606) );
  NAND U27861 ( .A(n26400), .B(n26399), .Z(n26404) );
  NAND U27862 ( .A(n26402), .B(n26401), .Z(n26403) );
  AND U27863 ( .A(n26404), .B(n26403), .Z(n26607) );
  XOR U27864 ( .A(n26606), .B(n26607), .Z(n26609) );
  NAND U27865 ( .A(n26406), .B(n26405), .Z(n26410) );
  NAND U27866 ( .A(n26408), .B(n26407), .Z(n26409) );
  NAND U27867 ( .A(n26410), .B(n26409), .Z(n26603) );
  NAND U27868 ( .A(n26412), .B(n26411), .Z(n26416) );
  NAND U27869 ( .A(n26414), .B(n26413), .Z(n26415) );
  NAND U27870 ( .A(n26416), .B(n26415), .Z(n26597) );
  NANDN U27871 ( .A(n27120), .B(n26548), .Z(n26420) );
  NAND U27872 ( .A(n26418), .B(n26417), .Z(n26419) );
  NAND U27873 ( .A(n26420), .B(n26419), .Z(n26524) );
  AND U27874 ( .A(x[485]), .B(y[7953]), .Z(n26570) );
  AND U27875 ( .A(x[497]), .B(y[7941]), .Z(n26571) );
  XOR U27876 ( .A(n26570), .B(n26571), .Z(n26572) );
  AND U27877 ( .A(x[496]), .B(y[7942]), .Z(n26573) );
  XOR U27878 ( .A(n26572), .B(n26573), .Z(n26523) );
  AND U27879 ( .A(y[7940]), .B(x[498]), .Z(n26422) );
  NAND U27880 ( .A(y[7946]), .B(x[492]), .Z(n26421) );
  XNOR U27881 ( .A(n26422), .B(n26421), .Z(n26549) );
  AND U27882 ( .A(x[484]), .B(y[7954]), .Z(n26550) );
  XOR U27883 ( .A(n26549), .B(n26550), .Z(n26522) );
  XOR U27884 ( .A(n26523), .B(n26522), .Z(n26525) );
  XNOR U27885 ( .A(n26524), .B(n26525), .Z(n26594) );
  NAND U27886 ( .A(x[499]), .B(y[7946]), .Z(n27624) );
  NANDN U27887 ( .A(n27624), .B(n26423), .Z(n26427) );
  NAND U27888 ( .A(n26425), .B(n26424), .Z(n26426) );
  AND U27889 ( .A(n26427), .B(n26426), .Z(n26595) );
  XOR U27890 ( .A(n26594), .B(n26595), .Z(n26596) );
  XNOR U27891 ( .A(n26597), .B(n26596), .Z(n26600) );
  NAND U27892 ( .A(n26429), .B(n26428), .Z(n26433) );
  NAND U27893 ( .A(n26431), .B(n26430), .Z(n26432) );
  NAND U27894 ( .A(n26433), .B(n26432), .Z(n26583) );
  NAND U27895 ( .A(n26435), .B(n26434), .Z(n26439) );
  NAND U27896 ( .A(n26437), .B(n26436), .Z(n26438) );
  NAND U27897 ( .A(n26439), .B(n26438), .Z(n26582) );
  XOR U27898 ( .A(n26583), .B(n26582), .Z(n26585) );
  AND U27899 ( .A(n26441), .B(n26440), .Z(n26445) );
  NAND U27900 ( .A(n26443), .B(n26442), .Z(n26444) );
  NANDN U27901 ( .A(n26445), .B(n26444), .Z(n26545) );
  AND U27902 ( .A(y[7945]), .B(x[493]), .Z(n26447) );
  NAND U27903 ( .A(y[7938]), .B(x[500]), .Z(n26446) );
  XNOR U27904 ( .A(n26447), .B(n26446), .Z(n26566) );
  AND U27905 ( .A(x[482]), .B(y[7956]), .Z(n26567) );
  XOR U27906 ( .A(n26566), .B(n26567), .Z(n26543) );
  AND U27907 ( .A(y[7952]), .B(x[486]), .Z(n26449) );
  NAND U27908 ( .A(y[7943]), .B(x[495]), .Z(n26448) );
  XNOR U27909 ( .A(n26449), .B(n26448), .Z(n26578) );
  XOR U27910 ( .A(n26543), .B(n26542), .Z(n26544) );
  XOR U27911 ( .A(n26545), .B(n26544), .Z(n26589) );
  AND U27912 ( .A(x[493]), .B(y[7954]), .Z(n27901) );
  NANDN U27913 ( .A(n26450), .B(n27901), .Z(n26454) );
  NAND U27914 ( .A(n26452), .B(n26451), .Z(n26453) );
  NAND U27915 ( .A(n26454), .B(n26453), .Z(n26513) );
  AND U27916 ( .A(x[481]), .B(y[7957]), .Z(n26536) );
  XOR U27917 ( .A(n26537), .B(n26536), .Z(n26535) );
  AND U27918 ( .A(o[277]), .B(n26455), .Z(n26534) );
  XOR U27919 ( .A(n26535), .B(n26534), .Z(n26511) );
  AND U27920 ( .A(x[494]), .B(y[7944]), .Z(n26528) );
  AND U27921 ( .A(x[483]), .B(y[7955]), .Z(n26529) );
  XOR U27922 ( .A(n26528), .B(n26529), .Z(n26530) );
  AND U27923 ( .A(x[499]), .B(y[7939]), .Z(n26531) );
  XOR U27924 ( .A(n26530), .B(n26531), .Z(n26510) );
  XOR U27925 ( .A(n26511), .B(n26510), .Z(n26512) );
  XOR U27926 ( .A(n26513), .B(n26512), .Z(n26588) );
  XOR U27927 ( .A(n26589), .B(n26588), .Z(n26591) );
  NAND U27928 ( .A(n26457), .B(n26456), .Z(n26461) );
  NAND U27929 ( .A(n26459), .B(n26458), .Z(n26460) );
  NAND U27930 ( .A(n26461), .B(n26460), .Z(n26505) );
  AND U27931 ( .A(x[498]), .B(y[7947]), .Z(n27626) );
  NAND U27932 ( .A(n27626), .B(n26462), .Z(n26466) );
  NAND U27933 ( .A(n26464), .B(n26463), .Z(n26465) );
  NAND U27934 ( .A(n26466), .B(n26465), .Z(n26504) );
  XOR U27935 ( .A(n26505), .B(n26504), .Z(n26507) );
  AND U27936 ( .A(x[494]), .B(y[7951]), .Z(n27636) );
  NAND U27937 ( .A(n27636), .B(n26577), .Z(n26469) );
  NAND U27938 ( .A(n26706), .B(n26467), .Z(n26468) );
  NAND U27939 ( .A(n26469), .B(n26468), .Z(n26519) );
  AND U27940 ( .A(x[480]), .B(y[7958]), .Z(n26553) );
  NAND U27941 ( .A(x[502]), .B(y[7936]), .Z(n26554) );
  AND U27942 ( .A(x[501]), .B(y[7937]), .Z(n26576) );
  XOR U27943 ( .A(o[278]), .B(n26576), .Z(n26555) );
  XOR U27944 ( .A(n26556), .B(n26555), .Z(n26517) );
  AND U27945 ( .A(y[7951]), .B(x[487]), .Z(n26471) );
  NAND U27946 ( .A(y[7950]), .B(x[488]), .Z(n26470) );
  XNOR U27947 ( .A(n26471), .B(n26470), .Z(n26559) );
  XOR U27948 ( .A(n26517), .B(n26516), .Z(n26518) );
  XOR U27949 ( .A(n26519), .B(n26518), .Z(n26506) );
  XOR U27950 ( .A(n26507), .B(n26506), .Z(n26590) );
  XOR U27951 ( .A(n26591), .B(n26590), .Z(n26584) );
  XOR U27952 ( .A(n26585), .B(n26584), .Z(n26601) );
  XOR U27953 ( .A(n26600), .B(n26601), .Z(n26602) );
  XOR U27954 ( .A(n26603), .B(n26602), .Z(n26608) );
  XOR U27955 ( .A(n26609), .B(n26608), .Z(n26495) );
  NAND U27956 ( .A(n26473), .B(n26472), .Z(n26477) );
  NAND U27957 ( .A(n26475), .B(n26474), .Z(n26476) );
  NAND U27958 ( .A(n26477), .B(n26476), .Z(n26493) );
  NAND U27959 ( .A(n26479), .B(n26478), .Z(n26483) );
  NAND U27960 ( .A(n26481), .B(n26480), .Z(n26482) );
  NAND U27961 ( .A(n26483), .B(n26482), .Z(n26492) );
  XOR U27962 ( .A(n26493), .B(n26492), .Z(n26494) );
  XOR U27963 ( .A(n26495), .B(n26494), .Z(n26619) );
  XOR U27964 ( .A(n26620), .B(n26619), .Z(n26621) );
  XNOR U27965 ( .A(n26622), .B(n26621), .Z(n26613) );
  IV U27966 ( .A(n26615), .Z(n26612) );
  XOR U27967 ( .A(n26612), .B(n26616), .Z(n26491) );
  XNOR U27968 ( .A(n26613), .B(n26491), .Z(N567) );
  NAND U27969 ( .A(n26493), .B(n26492), .Z(n26497) );
  NAND U27970 ( .A(n26495), .B(n26494), .Z(n26496) );
  AND U27971 ( .A(n26497), .B(n26496), .Z(n26767) );
  NAND U27972 ( .A(n26499), .B(n26498), .Z(n26503) );
  NAND U27973 ( .A(n26501), .B(n26500), .Z(n26502) );
  NAND U27974 ( .A(n26503), .B(n26502), .Z(n26742) );
  NAND U27975 ( .A(n26505), .B(n26504), .Z(n26509) );
  NAND U27976 ( .A(n26507), .B(n26506), .Z(n26508) );
  NAND U27977 ( .A(n26509), .B(n26508), .Z(n26689) );
  NAND U27978 ( .A(n26511), .B(n26510), .Z(n26515) );
  NAND U27979 ( .A(n26513), .B(n26512), .Z(n26514) );
  NAND U27980 ( .A(n26515), .B(n26514), .Z(n26687) );
  NAND U27981 ( .A(n26517), .B(n26516), .Z(n26521) );
  NAND U27982 ( .A(n26519), .B(n26518), .Z(n26520) );
  NAND U27983 ( .A(n26521), .B(n26520), .Z(n26686) );
  XOR U27984 ( .A(n26687), .B(n26686), .Z(n26688) );
  XOR U27985 ( .A(n26689), .B(n26688), .Z(n26754) );
  NAND U27986 ( .A(n26523), .B(n26522), .Z(n26527) );
  NAND U27987 ( .A(n26525), .B(n26524), .Z(n26526) );
  NAND U27988 ( .A(n26527), .B(n26526), .Z(n26752) );
  NAND U27989 ( .A(n26529), .B(n26528), .Z(n26533) );
  NAND U27990 ( .A(n26531), .B(n26530), .Z(n26532) );
  NAND U27991 ( .A(n26533), .B(n26532), .Z(n26633) );
  AND U27992 ( .A(n26535), .B(n26534), .Z(n26539) );
  NAND U27993 ( .A(n26537), .B(n26536), .Z(n26538) );
  NANDN U27994 ( .A(n26539), .B(n26538), .Z(n26632) );
  XOR U27995 ( .A(n26633), .B(n26632), .Z(n26635) );
  AND U27996 ( .A(y[7952]), .B(x[487]), .Z(n26541) );
  NAND U27997 ( .A(y[7950]), .B(x[489]), .Z(n26540) );
  XNOR U27998 ( .A(n26541), .B(n26540), .Z(n26707) );
  AND U27999 ( .A(x[490]), .B(y[7949]), .Z(n26639) );
  XOR U28000 ( .A(n26638), .B(n26639), .Z(n26641) );
  AND U28001 ( .A(x[486]), .B(y[7953]), .Z(n26698) );
  AND U28002 ( .A(x[495]), .B(y[7944]), .Z(n26699) );
  XOR U28003 ( .A(n26698), .B(n26699), .Z(n26700) );
  AND U28004 ( .A(x[491]), .B(y[7948]), .Z(n26701) );
  XOR U28005 ( .A(n26700), .B(n26701), .Z(n26640) );
  XOR U28006 ( .A(n26641), .B(n26640), .Z(n26634) );
  XOR U28007 ( .A(n26635), .B(n26634), .Z(n26751) );
  XOR U28008 ( .A(n26752), .B(n26751), .Z(n26753) );
  XOR U28009 ( .A(n26754), .B(n26753), .Z(n26740) );
  NAND U28010 ( .A(n26543), .B(n26542), .Z(n26547) );
  NAND U28011 ( .A(n26545), .B(n26544), .Z(n26546) );
  NAND U28012 ( .A(n26547), .B(n26546), .Z(n26734) );
  AND U28013 ( .A(x[498]), .B(y[7946]), .Z(n27467) );
  NAND U28014 ( .A(n27467), .B(n26548), .Z(n26552) );
  NAND U28015 ( .A(n26550), .B(n26549), .Z(n26551) );
  NAND U28016 ( .A(n26552), .B(n26551), .Z(n26675) );
  NANDN U28017 ( .A(n26554), .B(n26553), .Z(n26558) );
  NAND U28018 ( .A(n26556), .B(n26555), .Z(n26557) );
  NAND U28019 ( .A(n26558), .B(n26557), .Z(n26674) );
  XOR U28020 ( .A(n26675), .B(n26674), .Z(n26676) );
  NANDN U28021 ( .A(n26708), .B(n26706), .Z(n26562) );
  NANDN U28022 ( .A(n26560), .B(n26559), .Z(n26561) );
  NAND U28023 ( .A(n26562), .B(n26561), .Z(n26670) );
  AND U28024 ( .A(x[480]), .B(y[7959]), .Z(n26717) );
  AND U28025 ( .A(x[503]), .B(y[7936]), .Z(n26718) );
  XOR U28026 ( .A(n26717), .B(n26718), .Z(n26720) );
  AND U28027 ( .A(x[502]), .B(y[7937]), .Z(n26697) );
  XOR U28028 ( .A(o[279]), .B(n26697), .Z(n26719) );
  XOR U28029 ( .A(n26720), .B(n26719), .Z(n26669) );
  NAND U28030 ( .A(y[7939]), .B(x[500]), .Z(n26563) );
  XNOR U28031 ( .A(n26564), .B(n26563), .Z(n26693) );
  AND U28032 ( .A(x[499]), .B(y[7940]), .Z(n26694) );
  XOR U28033 ( .A(n26693), .B(n26694), .Z(n26668) );
  XOR U28034 ( .A(n26669), .B(n26668), .Z(n26671) );
  XOR U28035 ( .A(n26670), .B(n26671), .Z(n26677) );
  XOR U28036 ( .A(n26676), .B(n26677), .Z(n26733) );
  XOR U28037 ( .A(n26734), .B(n26733), .Z(n26736) );
  NAND U28038 ( .A(x[500]), .B(y[7945]), .Z(n27648) );
  AND U28039 ( .A(x[493]), .B(y[7938]), .Z(n26565) );
  NANDN U28040 ( .A(n27648), .B(n26565), .Z(n26569) );
  NAND U28041 ( .A(n26567), .B(n26566), .Z(n26568) );
  NAND U28042 ( .A(n26569), .B(n26568), .Z(n26728) );
  NAND U28043 ( .A(n26571), .B(n26570), .Z(n26575) );
  NAND U28044 ( .A(n26573), .B(n26572), .Z(n26574) );
  NAND U28045 ( .A(n26575), .B(n26574), .Z(n26682) );
  AND U28046 ( .A(x[493]), .B(y[7946]), .Z(n26656) );
  AND U28047 ( .A(x[482]), .B(y[7957]), .Z(n26657) );
  XOR U28048 ( .A(n26656), .B(n26657), .Z(n26658) );
  AND U28049 ( .A(x[501]), .B(y[7938]), .Z(n26659) );
  XOR U28050 ( .A(n26658), .B(n26659), .Z(n26681) );
  AND U28051 ( .A(x[492]), .B(y[7947]), .Z(n26711) );
  AND U28052 ( .A(x[481]), .B(y[7958]), .Z(n26712) );
  XOR U28053 ( .A(n26711), .B(n26712), .Z(n26714) );
  AND U28054 ( .A(o[278]), .B(n26576), .Z(n26713) );
  XOR U28055 ( .A(n26714), .B(n26713), .Z(n26680) );
  XOR U28056 ( .A(n26681), .B(n26680), .Z(n26683) );
  XOR U28057 ( .A(n26682), .B(n26683), .Z(n26727) );
  XOR U28058 ( .A(n26728), .B(n26727), .Z(n26730) );
  AND U28059 ( .A(x[495]), .B(y[7952]), .Z(n27889) );
  NAND U28060 ( .A(n27889), .B(n26577), .Z(n26581) );
  NANDN U28061 ( .A(n26579), .B(n26578), .Z(n26580) );
  NAND U28062 ( .A(n26581), .B(n26580), .Z(n26664) );
  AND U28063 ( .A(x[494]), .B(y[7945]), .Z(n26650) );
  AND U28064 ( .A(x[483]), .B(y[7956]), .Z(n26651) );
  XOR U28065 ( .A(n26650), .B(n26651), .Z(n26652) );
  AND U28066 ( .A(x[484]), .B(y[7955]), .Z(n26653) );
  XOR U28067 ( .A(n26652), .B(n26653), .Z(n26663) );
  AND U28068 ( .A(x[485]), .B(y[7954]), .Z(n26644) );
  AND U28069 ( .A(x[498]), .B(y[7941]), .Z(n26645) );
  XOR U28070 ( .A(n26644), .B(n26645), .Z(n26647) );
  AND U28071 ( .A(x[497]), .B(y[7942]), .Z(n26646) );
  XOR U28072 ( .A(n26647), .B(n26646), .Z(n26662) );
  XOR U28073 ( .A(n26663), .B(n26662), .Z(n26665) );
  XOR U28074 ( .A(n26664), .B(n26665), .Z(n26729) );
  XOR U28075 ( .A(n26730), .B(n26729), .Z(n26735) );
  XOR U28076 ( .A(n26736), .B(n26735), .Z(n26739) );
  XOR U28077 ( .A(n26740), .B(n26739), .Z(n26741) );
  XNOR U28078 ( .A(n26742), .B(n26741), .Z(n26628) );
  NAND U28079 ( .A(n26583), .B(n26582), .Z(n26587) );
  NAND U28080 ( .A(n26585), .B(n26584), .Z(n26586) );
  NAND U28081 ( .A(n26587), .B(n26586), .Z(n26748) );
  NAND U28082 ( .A(n26589), .B(n26588), .Z(n26593) );
  NAND U28083 ( .A(n26591), .B(n26590), .Z(n26592) );
  NAND U28084 ( .A(n26593), .B(n26592), .Z(n26746) );
  NAND U28085 ( .A(n26595), .B(n26594), .Z(n26599) );
  NAND U28086 ( .A(n26597), .B(n26596), .Z(n26598) );
  AND U28087 ( .A(n26599), .B(n26598), .Z(n26745) );
  XOR U28088 ( .A(n26746), .B(n26745), .Z(n26747) );
  XNOR U28089 ( .A(n26748), .B(n26747), .Z(n26626) );
  NAND U28090 ( .A(n26601), .B(n26600), .Z(n26605) );
  NAND U28091 ( .A(n26603), .B(n26602), .Z(n26604) );
  AND U28092 ( .A(n26605), .B(n26604), .Z(n26627) );
  XOR U28093 ( .A(n26626), .B(n26627), .Z(n26629) );
  XOR U28094 ( .A(n26628), .B(n26629), .Z(n26764) );
  NAND U28095 ( .A(n26607), .B(n26606), .Z(n26611) );
  NAND U28096 ( .A(n26609), .B(n26608), .Z(n26610) );
  AND U28097 ( .A(n26611), .B(n26610), .Z(n26765) );
  XOR U28098 ( .A(n26764), .B(n26765), .Z(n26766) );
  XNOR U28099 ( .A(n26767), .B(n26766), .Z(n26760) );
  NOR U28100 ( .A(n26612), .B(n26616), .Z(n26614) );
  OR U28101 ( .A(n26614), .B(n26613), .Z(n26618) );
  ANDN U28102 ( .B(n26616), .A(n26615), .Z(n26617) );
  ANDN U28103 ( .B(n26618), .A(n26617), .Z(n26758) );
  NAND U28104 ( .A(n26620), .B(n26619), .Z(n26624) );
  NAND U28105 ( .A(n26622), .B(n26621), .Z(n26623) );
  AND U28106 ( .A(n26624), .B(n26623), .Z(n26759) );
  IV U28107 ( .A(n26759), .Z(n26757) );
  XOR U28108 ( .A(n26758), .B(n26757), .Z(n26625) );
  XNOR U28109 ( .A(n26760), .B(n26625), .Z(N568) );
  NAND U28110 ( .A(n26627), .B(n26626), .Z(n26631) );
  NAND U28111 ( .A(n26629), .B(n26628), .Z(n26630) );
  AND U28112 ( .A(n26631), .B(n26630), .Z(n26908) );
  NAND U28113 ( .A(n26633), .B(n26632), .Z(n26637) );
  NAND U28114 ( .A(n26635), .B(n26634), .Z(n26636) );
  NAND U28115 ( .A(n26637), .B(n26636), .Z(n26845) );
  NAND U28116 ( .A(n26639), .B(n26638), .Z(n26643) );
  NAND U28117 ( .A(n26641), .B(n26640), .Z(n26642) );
  NAND U28118 ( .A(n26643), .B(n26642), .Z(n26843) );
  NAND U28119 ( .A(n26645), .B(n26644), .Z(n26649) );
  NAND U28120 ( .A(n26647), .B(n26646), .Z(n26648) );
  NAND U28121 ( .A(n26649), .B(n26648), .Z(n26869) );
  AND U28122 ( .A(x[480]), .B(y[7960]), .Z(n26824) );
  AND U28123 ( .A(x[504]), .B(y[7936]), .Z(n26825) );
  XOR U28124 ( .A(n26824), .B(n26825), .Z(n26827) );
  AND U28125 ( .A(x[503]), .B(y[7937]), .Z(n26817) );
  XOR U28126 ( .A(o[280]), .B(n26817), .Z(n26826) );
  XOR U28127 ( .A(n26827), .B(n26826), .Z(n26867) );
  AND U28128 ( .A(x[487]), .B(y[7953]), .Z(n26811) );
  NAND U28129 ( .A(x[498]), .B(y[7942]), .Z(n26812) );
  NAND U28130 ( .A(x[497]), .B(y[7943]), .Z(n26814) );
  XOR U28131 ( .A(n26867), .B(n26866), .Z(n26868) );
  XOR U28132 ( .A(n26869), .B(n26868), .Z(n26857) );
  NAND U28133 ( .A(n26651), .B(n26650), .Z(n26655) );
  NAND U28134 ( .A(n26653), .B(n26652), .Z(n26654) );
  NAND U28135 ( .A(n26655), .B(n26654), .Z(n26855) );
  NAND U28136 ( .A(n26657), .B(n26656), .Z(n26661) );
  NAND U28137 ( .A(n26659), .B(n26658), .Z(n26660) );
  NAND U28138 ( .A(n26661), .B(n26660), .Z(n26854) );
  XOR U28139 ( .A(n26855), .B(n26854), .Z(n26856) );
  XOR U28140 ( .A(n26857), .B(n26856), .Z(n26842) );
  XOR U28141 ( .A(n26843), .B(n26842), .Z(n26844) );
  XNOR U28142 ( .A(n26845), .B(n26844), .Z(n26850) );
  NAND U28143 ( .A(n26663), .B(n26662), .Z(n26667) );
  NAND U28144 ( .A(n26665), .B(n26664), .Z(n26666) );
  AND U28145 ( .A(n26667), .B(n26666), .Z(n26897) );
  NAND U28146 ( .A(n26669), .B(n26668), .Z(n26673) );
  NAND U28147 ( .A(n26671), .B(n26670), .Z(n26672) );
  AND U28148 ( .A(n26673), .B(n26672), .Z(n26896) );
  XOR U28149 ( .A(n26897), .B(n26896), .Z(n26899) );
  NAND U28150 ( .A(n26675), .B(n26674), .Z(n26679) );
  NAND U28151 ( .A(n26677), .B(n26676), .Z(n26678) );
  AND U28152 ( .A(n26679), .B(n26678), .Z(n26898) );
  XOR U28153 ( .A(n26899), .B(n26898), .Z(n26848) );
  NAND U28154 ( .A(n26681), .B(n26680), .Z(n26685) );
  NAND U28155 ( .A(n26683), .B(n26682), .Z(n26684) );
  NAND U28156 ( .A(n26685), .B(n26684), .Z(n26849) );
  XOR U28157 ( .A(n26850), .B(n26851), .Z(n26777) );
  NAND U28158 ( .A(n26687), .B(n26686), .Z(n26691) );
  NAND U28159 ( .A(n26689), .B(n26688), .Z(n26690) );
  AND U28160 ( .A(n26691), .B(n26690), .Z(n26778) );
  XOR U28161 ( .A(n26777), .B(n26778), .Z(n26780) );
  AND U28162 ( .A(x[500]), .B(y[7943]), .Z(n26692) );
  NAND U28163 ( .A(n26692), .B(n26872), .Z(n26696) );
  NAND U28164 ( .A(n26694), .B(n26693), .Z(n26695) );
  NAND U28165 ( .A(n26696), .B(n26695), .Z(n26893) );
  AND U28166 ( .A(x[502]), .B(y[7938]), .Z(n26799) );
  XOR U28167 ( .A(n26800), .B(n26799), .Z(n26802) );
  NAND U28168 ( .A(x[482]), .B(y[7958]), .Z(n26801) );
  AND U28169 ( .A(x[481]), .B(y[7959]), .Z(n26807) );
  XOR U28170 ( .A(n26808), .B(n26807), .Z(n26806) );
  AND U28171 ( .A(o[279]), .B(n26697), .Z(n26805) );
  XOR U28172 ( .A(n26806), .B(n26805), .Z(n26890) );
  XOR U28173 ( .A(n26891), .B(n26890), .Z(n26892) );
  XOR U28174 ( .A(n26893), .B(n26892), .Z(n26837) );
  NAND U28175 ( .A(n26699), .B(n26698), .Z(n26703) );
  NAND U28176 ( .A(n26701), .B(n26700), .Z(n26702) );
  NAND U28177 ( .A(n26703), .B(n26702), .Z(n26887) );
  AND U28178 ( .A(y[7944]), .B(x[496]), .Z(n26705) );
  NAND U28179 ( .A(y[7939]), .B(x[501]), .Z(n26704) );
  XNOR U28180 ( .A(n26705), .B(n26704), .Z(n26873) );
  AND U28181 ( .A(x[485]), .B(y[7955]), .Z(n26874) );
  XOR U28182 ( .A(n26873), .B(n26874), .Z(n26885) );
  AND U28183 ( .A(x[486]), .B(y[7954]), .Z(n27211) );
  NAND U28184 ( .A(x[500]), .B(y[7940]), .Z(n26879) );
  IV U28185 ( .A(n26879), .Z(n27011) );
  XOR U28186 ( .A(n27211), .B(n27011), .Z(n26880) );
  AND U28187 ( .A(x[499]), .B(y[7941]), .Z(n26881) );
  XOR U28188 ( .A(n26880), .B(n26881), .Z(n26884) );
  XOR U28189 ( .A(n26885), .B(n26884), .Z(n26886) );
  XOR U28190 ( .A(n26887), .B(n26886), .Z(n26863) );
  NANDN U28191 ( .A(n26937), .B(n26706), .Z(n26710) );
  NANDN U28192 ( .A(n26708), .B(n26707), .Z(n26709) );
  NAND U28193 ( .A(n26710), .B(n26709), .Z(n26861) );
  NAND U28194 ( .A(n26712), .B(n26711), .Z(n26716) );
  NAND U28195 ( .A(n26714), .B(n26713), .Z(n26715) );
  NAND U28196 ( .A(n26716), .B(n26715), .Z(n26860) );
  XOR U28197 ( .A(n26861), .B(n26860), .Z(n26862) );
  XOR U28198 ( .A(n26863), .B(n26862), .Z(n26836) );
  XOR U28199 ( .A(n26837), .B(n26836), .Z(n26839) );
  NAND U28200 ( .A(n26718), .B(n26717), .Z(n26722) );
  NAND U28201 ( .A(n26720), .B(n26719), .Z(n26721) );
  AND U28202 ( .A(n26722), .B(n26721), .Z(n26831) );
  AND U28203 ( .A(x[483]), .B(y[7957]), .Z(n26820) );
  XOR U28204 ( .A(n26821), .B(n26820), .Z(n26819) );
  AND U28205 ( .A(x[484]), .B(y[7956]), .Z(n26818) );
  XOR U28206 ( .A(n26819), .B(n26818), .Z(n26830) );
  AND U28207 ( .A(y[7951]), .B(x[489]), .Z(n26724) );
  NAND U28208 ( .A(y[7950]), .B(x[490]), .Z(n26723) );
  XNOR U28209 ( .A(n26724), .B(n26723), .Z(n26791) );
  AND U28210 ( .A(y[7946]), .B(x[494]), .Z(n26726) );
  NAND U28211 ( .A(y[7952]), .B(x[488]), .Z(n26725) );
  XNOR U28212 ( .A(n26726), .B(n26725), .Z(n26795) );
  AND U28213 ( .A(x[491]), .B(y[7949]), .Z(n26796) );
  XOR U28214 ( .A(n26795), .B(n26796), .Z(n26790) );
  XOR U28215 ( .A(n26791), .B(n26790), .Z(n26832) );
  XOR U28216 ( .A(n26833), .B(n26832), .Z(n26838) );
  XOR U28217 ( .A(n26839), .B(n26838), .Z(n26784) );
  NAND U28218 ( .A(n26728), .B(n26727), .Z(n26732) );
  NAND U28219 ( .A(n26730), .B(n26729), .Z(n26731) );
  AND U28220 ( .A(n26732), .B(n26731), .Z(n26783) );
  NAND U28221 ( .A(n26734), .B(n26733), .Z(n26738) );
  NAND U28222 ( .A(n26736), .B(n26735), .Z(n26737) );
  NAND U28223 ( .A(n26738), .B(n26737), .Z(n26786) );
  XNOR U28224 ( .A(n26780), .B(n26779), .Z(n26906) );
  NAND U28225 ( .A(n26740), .B(n26739), .Z(n26744) );
  NAND U28226 ( .A(n26742), .B(n26741), .Z(n26743) );
  NAND U28227 ( .A(n26744), .B(n26743), .Z(n26774) );
  NAND U28228 ( .A(n26746), .B(n26745), .Z(n26750) );
  NAND U28229 ( .A(n26748), .B(n26747), .Z(n26749) );
  NAND U28230 ( .A(n26750), .B(n26749), .Z(n26772) );
  NAND U28231 ( .A(n26752), .B(n26751), .Z(n26756) );
  NAND U28232 ( .A(n26754), .B(n26753), .Z(n26755) );
  NAND U28233 ( .A(n26756), .B(n26755), .Z(n26771) );
  XOR U28234 ( .A(n26772), .B(n26771), .Z(n26773) );
  XOR U28235 ( .A(n26774), .B(n26773), .Z(n26905) );
  XOR U28236 ( .A(n26906), .B(n26905), .Z(n26907) );
  XNOR U28237 ( .A(n26908), .B(n26907), .Z(n26904) );
  NANDN U28238 ( .A(n26757), .B(n26758), .Z(n26763) );
  NOR U28239 ( .A(n26759), .B(n26758), .Z(n26761) );
  OR U28240 ( .A(n26761), .B(n26760), .Z(n26762) );
  AND U28241 ( .A(n26763), .B(n26762), .Z(n26902) );
  NAND U28242 ( .A(n26765), .B(n26764), .Z(n26769) );
  NAND U28243 ( .A(n26767), .B(n26766), .Z(n26768) );
  AND U28244 ( .A(n26769), .B(n26768), .Z(n26903) );
  XOR U28245 ( .A(n26902), .B(n26903), .Z(n26770) );
  XNOR U28246 ( .A(n26904), .B(n26770), .Z(N569) );
  NAND U28247 ( .A(n26772), .B(n26771), .Z(n26776) );
  NAND U28248 ( .A(n26774), .B(n26773), .Z(n26775) );
  AND U28249 ( .A(n26776), .B(n26775), .Z(n27062) );
  NAND U28250 ( .A(n26778), .B(n26777), .Z(n26782) );
  NAND U28251 ( .A(n26780), .B(n26779), .Z(n26781) );
  NAND U28252 ( .A(n26782), .B(n26781), .Z(n27060) );
  NANDN U28253 ( .A(n26784), .B(n26783), .Z(n26788) );
  NANDN U28254 ( .A(n26786), .B(n26785), .Z(n26787) );
  AND U28255 ( .A(n26788), .B(n26787), .Z(n26913) );
  NANDN U28256 ( .A(n26936), .B(n26789), .Z(n26793) );
  NAND U28257 ( .A(n26791), .B(n26790), .Z(n26792) );
  NAND U28258 ( .A(n26793), .B(n26792), .Z(n26961) );
  AND U28259 ( .A(x[494]), .B(y[7952]), .Z(n27835) );
  NAND U28260 ( .A(n27835), .B(n26794), .Z(n26798) );
  NAND U28261 ( .A(n26796), .B(n26795), .Z(n26797) );
  NAND U28262 ( .A(n26798), .B(n26797), .Z(n26988) );
  NAND U28263 ( .A(x[491]), .B(y[7950]), .Z(n27007) );
  NAND U28264 ( .A(x[492]), .B(y[7949]), .Z(n27006) );
  NAND U28265 ( .A(x[487]), .B(y[7954]), .Z(n27005) );
  XOR U28266 ( .A(n27006), .B(n27005), .Z(n27008) );
  XNOR U28267 ( .A(n27007), .B(n27008), .Z(n26987) );
  AND U28268 ( .A(x[504]), .B(y[7937]), .Z(n27004) );
  XOR U28269 ( .A(o[281]), .B(n27004), .Z(n26975) );
  AND U28270 ( .A(x[481]), .B(y[7960]), .Z(n26974) );
  XOR U28271 ( .A(n26975), .B(n26974), .Z(n26977) );
  AND U28272 ( .A(x[493]), .B(y[7948]), .Z(n26976) );
  XOR U28273 ( .A(n26977), .B(n26976), .Z(n26986) );
  XOR U28274 ( .A(n26987), .B(n26986), .Z(n26989) );
  XOR U28275 ( .A(n26988), .B(n26989), .Z(n26960) );
  XOR U28276 ( .A(n26961), .B(n26960), .Z(n26963) );
  NAND U28277 ( .A(n26800), .B(n26799), .Z(n26804) );
  ANDN U28278 ( .B(n26802), .A(n26801), .Z(n26803) );
  ANDN U28279 ( .B(n26804), .A(n26803), .Z(n26949) );
  AND U28280 ( .A(n26806), .B(n26805), .Z(n26810) );
  NAND U28281 ( .A(n26808), .B(n26807), .Z(n26809) );
  NANDN U28282 ( .A(n26810), .B(n26809), .Z(n26948) );
  NANDN U28283 ( .A(n26812), .B(n26811), .Z(n26816) );
  NANDN U28284 ( .A(n26814), .B(n26813), .Z(n26815) );
  AND U28285 ( .A(n26816), .B(n26815), .Z(n26945) );
  NAND U28286 ( .A(x[488]), .B(y[7953]), .Z(n26938) );
  XOR U28287 ( .A(n26937), .B(n26936), .Z(n26939) );
  XNOR U28288 ( .A(n26938), .B(n26939), .Z(n26943) );
  NAND U28289 ( .A(n26817), .B(o[280]), .Z(n26932) );
  NAND U28290 ( .A(x[505]), .B(y[7936]), .Z(n26931) );
  NAND U28291 ( .A(x[480]), .B(y[7961]), .Z(n26930) );
  XNOR U28292 ( .A(n26931), .B(n26930), .Z(n26933) );
  XOR U28293 ( .A(n26932), .B(n26933), .Z(n26942) );
  XOR U28294 ( .A(n26943), .B(n26942), .Z(n26944) );
  XOR U28295 ( .A(n26951), .B(n26950), .Z(n26962) );
  XOR U28296 ( .A(n26963), .B(n26962), .Z(n27043) );
  AND U28297 ( .A(n26819), .B(n26818), .Z(n26823) );
  NAND U28298 ( .A(n26821), .B(n26820), .Z(n26822) );
  NANDN U28299 ( .A(n26823), .B(n26822), .Z(n27025) );
  NAND U28300 ( .A(n26825), .B(n26824), .Z(n26829) );
  NAND U28301 ( .A(n26827), .B(n26826), .Z(n26828) );
  NAND U28302 ( .A(n26829), .B(n26828), .Z(n27023) );
  AND U28303 ( .A(x[494]), .B(y[7947]), .Z(n26981) );
  AND U28304 ( .A(x[482]), .B(y[7959]), .Z(n26980) );
  XOR U28305 ( .A(n26981), .B(n26980), .Z(n26983) );
  AND U28306 ( .A(x[483]), .B(y[7958]), .Z(n26982) );
  XOR U28307 ( .A(n26983), .B(n26982), .Z(n27022) );
  XOR U28308 ( .A(n27023), .B(n27022), .Z(n27024) );
  XNOR U28309 ( .A(n27025), .B(n27024), .Z(n27040) );
  NANDN U28310 ( .A(n26831), .B(n26830), .Z(n26835) );
  NAND U28311 ( .A(n26833), .B(n26832), .Z(n26834) );
  AND U28312 ( .A(n26835), .B(n26834), .Z(n27041) );
  XOR U28313 ( .A(n27040), .B(n27041), .Z(n27042) );
  NAND U28314 ( .A(n26837), .B(n26836), .Z(n26841) );
  NAND U28315 ( .A(n26839), .B(n26838), .Z(n26840) );
  AND U28316 ( .A(n26841), .B(n26840), .Z(n27047) );
  XOR U28317 ( .A(n27046), .B(n27047), .Z(n27048) );
  NAND U28318 ( .A(n26843), .B(n26842), .Z(n26847) );
  NAND U28319 ( .A(n26845), .B(n26844), .Z(n26846) );
  AND U28320 ( .A(n26847), .B(n26846), .Z(n27049) );
  XOR U28321 ( .A(n27048), .B(n27049), .Z(n26912) );
  NANDN U28322 ( .A(n26849), .B(n26848), .Z(n26853) );
  NAND U28323 ( .A(n26851), .B(n26850), .Z(n26852) );
  NAND U28324 ( .A(n26853), .B(n26852), .Z(n26920) );
  NAND U28325 ( .A(n26855), .B(n26854), .Z(n26859) );
  NAND U28326 ( .A(n26857), .B(n26856), .Z(n26858) );
  NAND U28327 ( .A(n26859), .B(n26858), .Z(n26925) );
  NAND U28328 ( .A(n26861), .B(n26860), .Z(n26865) );
  NAND U28329 ( .A(n26863), .B(n26862), .Z(n26864) );
  NAND U28330 ( .A(n26865), .B(n26864), .Z(n26924) );
  XOR U28331 ( .A(n26925), .B(n26924), .Z(n26927) );
  NAND U28332 ( .A(n26867), .B(n26866), .Z(n26871) );
  NAND U28333 ( .A(n26869), .B(n26868), .Z(n26870) );
  AND U28334 ( .A(n26871), .B(n26870), .Z(n26957) );
  NAND U28335 ( .A(x[501]), .B(y[7944]), .Z(n27790) );
  NANDN U28336 ( .A(n27790), .B(n26872), .Z(n26876) );
  NAND U28337 ( .A(n26874), .B(n26873), .Z(n26875) );
  NAND U28338 ( .A(n26876), .B(n26875), .Z(n27031) );
  NAND U28339 ( .A(x[502]), .B(y[7939]), .Z(n27000) );
  NAND U28340 ( .A(x[485]), .B(y[7956]), .Z(n26999) );
  NAND U28341 ( .A(x[497]), .B(y[7944]), .Z(n26998) );
  XOR U28342 ( .A(n26999), .B(n26998), .Z(n27001) );
  XNOR U28343 ( .A(n27000), .B(n27001), .Z(n27028) );
  AND U28344 ( .A(y[7941]), .B(x[500]), .Z(n26878) );
  NAND U28345 ( .A(y[7940]), .B(x[501]), .Z(n26877) );
  XNOR U28346 ( .A(n26878), .B(n26877), .Z(n27013) );
  AND U28347 ( .A(x[499]), .B(y[7942]), .Z(n27012) );
  XOR U28348 ( .A(n27013), .B(n27012), .Z(n27029) );
  XOR U28349 ( .A(n27028), .B(n27029), .Z(n27030) );
  XNOR U28350 ( .A(n27031), .B(n27030), .Z(n26955) );
  NANDN U28351 ( .A(n26879), .B(n27211), .Z(n26883) );
  NAND U28352 ( .A(n26881), .B(n26880), .Z(n26882) );
  AND U28353 ( .A(n26883), .B(n26882), .Z(n27037) );
  NAND U28354 ( .A(x[495]), .B(y[7946]), .Z(n27018) );
  NAND U28355 ( .A(x[498]), .B(y[7943]), .Z(n27017) );
  NAND U28356 ( .A(x[486]), .B(y[7955]), .Z(n27016) );
  XOR U28357 ( .A(n27017), .B(n27016), .Z(n27019) );
  XNOR U28358 ( .A(n27018), .B(n27019), .Z(n27035) );
  NAND U28359 ( .A(x[503]), .B(y[7938]), .Z(n26994) );
  NAND U28360 ( .A(x[484]), .B(y[7957]), .Z(n26993) );
  NAND U28361 ( .A(x[496]), .B(y[7945]), .Z(n26992) );
  XNOR U28362 ( .A(n26993), .B(n26992), .Z(n26995) );
  XOR U28363 ( .A(n26994), .B(n26995), .Z(n27034) );
  XOR U28364 ( .A(n27035), .B(n27034), .Z(n27036) );
  XOR U28365 ( .A(n27037), .B(n27036), .Z(n26954) );
  XOR U28366 ( .A(n26955), .B(n26954), .Z(n26956) );
  XNOR U28367 ( .A(n26957), .B(n26956), .Z(n26969) );
  NAND U28368 ( .A(n26885), .B(n26884), .Z(n26889) );
  NAND U28369 ( .A(n26887), .B(n26886), .Z(n26888) );
  NAND U28370 ( .A(n26889), .B(n26888), .Z(n26967) );
  NAND U28371 ( .A(n26891), .B(n26890), .Z(n26895) );
  NAND U28372 ( .A(n26893), .B(n26892), .Z(n26894) );
  NAND U28373 ( .A(n26895), .B(n26894), .Z(n26966) );
  XOR U28374 ( .A(n26967), .B(n26966), .Z(n26968) );
  XOR U28375 ( .A(n26969), .B(n26968), .Z(n26926) );
  XOR U28376 ( .A(n26927), .B(n26926), .Z(n26919) );
  NAND U28377 ( .A(n26897), .B(n26896), .Z(n26901) );
  NAND U28378 ( .A(n26899), .B(n26898), .Z(n26900) );
  NAND U28379 ( .A(n26901), .B(n26900), .Z(n26918) );
  XOR U28380 ( .A(n26920), .B(n26921), .Z(n26914) );
  XOR U28381 ( .A(n26915), .B(n26914), .Z(n27059) );
  XOR U28382 ( .A(n27060), .B(n27059), .Z(n27061) );
  XNOR U28383 ( .A(n27062), .B(n27061), .Z(n27055) );
  NAND U28384 ( .A(n26906), .B(n26905), .Z(n26910) );
  NAND U28385 ( .A(n26908), .B(n26907), .Z(n26909) );
  AND U28386 ( .A(n26910), .B(n26909), .Z(n27054) );
  IV U28387 ( .A(n27054), .Z(n27052) );
  XOR U28388 ( .A(n27053), .B(n27052), .Z(n26911) );
  XNOR U28389 ( .A(n27055), .B(n26911), .Z(N570) );
  NANDN U28390 ( .A(n26913), .B(n26912), .Z(n26917) );
  NAND U28391 ( .A(n26915), .B(n26914), .Z(n26916) );
  AND U28392 ( .A(n26917), .B(n26916), .Z(n27066) );
  NANDN U28393 ( .A(n26919), .B(n26918), .Z(n26923) );
  NAND U28394 ( .A(n26921), .B(n26920), .Z(n26922) );
  NAND U28395 ( .A(n26923), .B(n26922), .Z(n27067) );
  NAND U28396 ( .A(n26925), .B(n26924), .Z(n26929) );
  NAND U28397 ( .A(n26927), .B(n26926), .Z(n26928) );
  NAND U28398 ( .A(n26929), .B(n26928), .Z(n27084) );
  AND U28399 ( .A(x[482]), .B(y[7960]), .Z(n27105) );
  XOR U28400 ( .A(n27106), .B(n27105), .Z(n27108) );
  AND U28401 ( .A(x[504]), .B(y[7938]), .Z(n27107) );
  XOR U28402 ( .A(n27108), .B(n27107), .Z(n27142) );
  NAND U28403 ( .A(n26931), .B(n26930), .Z(n26935) );
  NANDN U28404 ( .A(n26933), .B(n26932), .Z(n26934) );
  AND U28405 ( .A(n26935), .B(n26934), .Z(n27141) );
  XOR U28406 ( .A(n27142), .B(n27141), .Z(n27144) );
  NAND U28407 ( .A(n26937), .B(n26936), .Z(n26941) );
  NAND U28408 ( .A(n26939), .B(n26938), .Z(n26940) );
  AND U28409 ( .A(n26941), .B(n26940), .Z(n27143) );
  XOR U28410 ( .A(n27144), .B(n27143), .Z(n27180) );
  NAND U28411 ( .A(n26943), .B(n26942), .Z(n26947) );
  NANDN U28412 ( .A(n26945), .B(n26944), .Z(n26946) );
  AND U28413 ( .A(n26947), .B(n26946), .Z(n27179) );
  NANDN U28414 ( .A(n26949), .B(n26948), .Z(n26953) );
  NAND U28415 ( .A(n26951), .B(n26950), .Z(n26952) );
  NAND U28416 ( .A(n26953), .B(n26952), .Z(n27182) );
  NAND U28417 ( .A(n26955), .B(n26954), .Z(n26959) );
  NAND U28418 ( .A(n26957), .B(n26956), .Z(n26958) );
  NAND U28419 ( .A(n26959), .B(n26958), .Z(n27174) );
  NAND U28420 ( .A(n26961), .B(n26960), .Z(n26965) );
  NAND U28421 ( .A(n26963), .B(n26962), .Z(n26964) );
  AND U28422 ( .A(n26965), .B(n26964), .Z(n27173) );
  XOR U28423 ( .A(n27174), .B(n27173), .Z(n27175) );
  XNOR U28424 ( .A(n27176), .B(n27175), .Z(n27082) );
  NAND U28425 ( .A(n26967), .B(n26966), .Z(n26971) );
  NAND U28426 ( .A(n26969), .B(n26968), .Z(n26970) );
  NAND U28427 ( .A(n26971), .B(n26970), .Z(n27090) );
  AND U28428 ( .A(x[492]), .B(y[7950]), .Z(n27291) );
  AND U28429 ( .A(x[485]), .B(y[7957]), .Z(n27156) );
  XOR U28430 ( .A(n27291), .B(n27156), .Z(n27158) );
  AND U28431 ( .A(x[490]), .B(y[7952]), .Z(n27157) );
  XOR U28432 ( .A(n27158), .B(n27157), .Z(n27188) );
  AND U28433 ( .A(x[487]), .B(y[7955]), .Z(n27186) );
  AND U28434 ( .A(y[7956]), .B(x[486]), .Z(n26973) );
  NAND U28435 ( .A(y[7954]), .B(x[488]), .Z(n26972) );
  XNOR U28436 ( .A(n26973), .B(n26972), .Z(n27213) );
  AND U28437 ( .A(x[489]), .B(y[7953]), .Z(n27212) );
  XOR U28438 ( .A(n27213), .B(n27212), .Z(n27185) );
  XOR U28439 ( .A(n27186), .B(n27185), .Z(n27187) );
  XOR U28440 ( .A(n27188), .B(n27187), .Z(n27131) );
  NAND U28441 ( .A(n26975), .B(n26974), .Z(n26979) );
  NAND U28442 ( .A(n26977), .B(n26976), .Z(n26978) );
  NAND U28443 ( .A(n26979), .B(n26978), .Z(n27130) );
  NAND U28444 ( .A(n26981), .B(n26980), .Z(n26985) );
  NAND U28445 ( .A(n26983), .B(n26982), .Z(n26984) );
  NAND U28446 ( .A(n26985), .B(n26984), .Z(n27129) );
  XOR U28447 ( .A(n27130), .B(n27129), .Z(n27132) );
  XNOR U28448 ( .A(n27131), .B(n27132), .Z(n27168) );
  NAND U28449 ( .A(n26987), .B(n26986), .Z(n26991) );
  NAND U28450 ( .A(n26989), .B(n26988), .Z(n26990) );
  AND U28451 ( .A(n26991), .B(n26990), .Z(n27167) );
  XOR U28452 ( .A(n27168), .B(n27167), .Z(n27170) );
  NAND U28453 ( .A(n26993), .B(n26992), .Z(n26997) );
  NANDN U28454 ( .A(n26995), .B(n26994), .Z(n26996) );
  AND U28455 ( .A(n26997), .B(n26996), .Z(n27094) );
  NAND U28456 ( .A(n26999), .B(n26998), .Z(n27003) );
  NAND U28457 ( .A(n27001), .B(n27000), .Z(n27002) );
  AND U28458 ( .A(n27003), .B(n27002), .Z(n27093) );
  XOR U28459 ( .A(n27094), .B(n27093), .Z(n27096) );
  AND U28460 ( .A(o[281]), .B(n27004), .Z(n27205) );
  NAND U28461 ( .A(x[494]), .B(y[7948]), .Z(n27206) );
  NAND U28462 ( .A(x[481]), .B(y[7961]), .Z(n27208) );
  NAND U28463 ( .A(x[505]), .B(y[7937]), .Z(n27216) );
  AND U28464 ( .A(x[506]), .B(y[7936]), .Z(n27161) );
  XOR U28465 ( .A(n27162), .B(n27161), .Z(n27164) );
  AND U28466 ( .A(x[480]), .B(y[7962]), .Z(n27163) );
  XOR U28467 ( .A(n27164), .B(n27163), .Z(n27147) );
  XOR U28468 ( .A(n27148), .B(n27147), .Z(n27150) );
  NAND U28469 ( .A(n27006), .B(n27005), .Z(n27010) );
  NAND U28470 ( .A(n27008), .B(n27007), .Z(n27009) );
  AND U28471 ( .A(n27010), .B(n27009), .Z(n27149) );
  XOR U28472 ( .A(n27150), .B(n27149), .Z(n27095) );
  XNOR U28473 ( .A(n27096), .B(n27095), .Z(n27138) );
  NAND U28474 ( .A(x[501]), .B(y[7941]), .Z(n27199) );
  NANDN U28475 ( .A(n27199), .B(n27011), .Z(n27015) );
  NAND U28476 ( .A(n27013), .B(n27012), .Z(n27014) );
  NAND U28477 ( .A(n27015), .B(n27014), .Z(n27125) );
  XNOR U28478 ( .A(n27200), .B(n27199), .Z(n27201) );
  NAND U28479 ( .A(x[500]), .B(y[7942]), .Z(n27202) );
  AND U28480 ( .A(x[503]), .B(y[7939]), .Z(n27111) );
  XOR U28481 ( .A(n27112), .B(n27111), .Z(n27114) );
  AND U28482 ( .A(x[502]), .B(y[7940]), .Z(n27113) );
  XOR U28483 ( .A(n27114), .B(n27113), .Z(n27123) );
  XOR U28484 ( .A(n27124), .B(n27123), .Z(n27126) );
  XNOR U28485 ( .A(n27125), .B(n27126), .Z(n27136) );
  AND U28486 ( .A(x[484]), .B(y[7958]), .Z(n27117) );
  XOR U28487 ( .A(n27118), .B(n27117), .Z(n27119) );
  XNOR U28488 ( .A(n27119), .B(n27120), .Z(n27100) );
  AND U28489 ( .A(x[483]), .B(y[7959]), .Z(n27191) );
  NAND U28490 ( .A(x[499]), .B(y[7943]), .Z(n27192) );
  AND U28491 ( .A(x[491]), .B(y[7951]), .Z(n27193) );
  XOR U28492 ( .A(n27194), .B(n27193), .Z(n27099) );
  XOR U28493 ( .A(n27100), .B(n27099), .Z(n27102) );
  NAND U28494 ( .A(n27017), .B(n27016), .Z(n27021) );
  NAND U28495 ( .A(n27019), .B(n27018), .Z(n27020) );
  AND U28496 ( .A(n27021), .B(n27020), .Z(n27101) );
  XNOR U28497 ( .A(n27102), .B(n27101), .Z(n27135) );
  XOR U28498 ( .A(n27136), .B(n27135), .Z(n27137) );
  XOR U28499 ( .A(n27138), .B(n27137), .Z(n27169) );
  XNOR U28500 ( .A(n27170), .B(n27169), .Z(n27088) );
  NAND U28501 ( .A(n27023), .B(n27022), .Z(n27027) );
  NAND U28502 ( .A(n27025), .B(n27024), .Z(n27026) );
  AND U28503 ( .A(n27027), .B(n27026), .Z(n27220) );
  NAND U28504 ( .A(n27029), .B(n27028), .Z(n27033) );
  NAND U28505 ( .A(n27031), .B(n27030), .Z(n27032) );
  AND U28506 ( .A(n27033), .B(n27032), .Z(n27218) );
  NAND U28507 ( .A(n27035), .B(n27034), .Z(n27039) );
  NANDN U28508 ( .A(n27037), .B(n27036), .Z(n27038) );
  NAND U28509 ( .A(n27039), .B(n27038), .Z(n27217) );
  XOR U28510 ( .A(n27088), .B(n27087), .Z(n27089) );
  XOR U28511 ( .A(n27090), .B(n27089), .Z(n27081) );
  XOR U28512 ( .A(n27082), .B(n27081), .Z(n27083) );
  XOR U28513 ( .A(n27084), .B(n27083), .Z(n27078) );
  NAND U28514 ( .A(n27041), .B(n27040), .Z(n27045) );
  NANDN U28515 ( .A(n27043), .B(n27042), .Z(n27044) );
  AND U28516 ( .A(n27045), .B(n27044), .Z(n27075) );
  NAND U28517 ( .A(n27047), .B(n27046), .Z(n27051) );
  NAND U28518 ( .A(n27049), .B(n27048), .Z(n27050) );
  AND U28519 ( .A(n27051), .B(n27050), .Z(n27076) );
  XOR U28520 ( .A(n27075), .B(n27076), .Z(n27077) );
  XOR U28521 ( .A(n27078), .B(n27077), .Z(n27068) );
  XNOR U28522 ( .A(n27069), .B(n27068), .Z(n27074) );
  NANDN U28523 ( .A(n27052), .B(n27053), .Z(n27058) );
  NOR U28524 ( .A(n27054), .B(n27053), .Z(n27056) );
  OR U28525 ( .A(n27056), .B(n27055), .Z(n27057) );
  AND U28526 ( .A(n27058), .B(n27057), .Z(n27072) );
  NAND U28527 ( .A(n27060), .B(n27059), .Z(n27064) );
  NAND U28528 ( .A(n27062), .B(n27061), .Z(n27063) );
  AND U28529 ( .A(n27064), .B(n27063), .Z(n27073) );
  XOR U28530 ( .A(n27072), .B(n27073), .Z(n27065) );
  XNOR U28531 ( .A(n27074), .B(n27065), .Z(N571) );
  NANDN U28532 ( .A(n27067), .B(n27066), .Z(n27071) );
  NAND U28533 ( .A(n27069), .B(n27068), .Z(n27070) );
  NAND U28534 ( .A(n27071), .B(n27070), .Z(n27231) );
  IV U28535 ( .A(n27231), .Z(n27230) );
  NAND U28536 ( .A(n27076), .B(n27075), .Z(n27080) );
  NAND U28537 ( .A(n27078), .B(n27077), .Z(n27079) );
  AND U28538 ( .A(n27080), .B(n27079), .Z(n27227) );
  NAND U28539 ( .A(n27082), .B(n27081), .Z(n27086) );
  NAND U28540 ( .A(n27084), .B(n27083), .Z(n27085) );
  AND U28541 ( .A(n27086), .B(n27085), .Z(n27225) );
  NAND U28542 ( .A(n27088), .B(n27087), .Z(n27092) );
  NAND U28543 ( .A(n27090), .B(n27089), .Z(n27091) );
  NAND U28544 ( .A(n27092), .B(n27091), .Z(n27239) );
  NAND U28545 ( .A(n27094), .B(n27093), .Z(n27098) );
  NAND U28546 ( .A(n27096), .B(n27095), .Z(n27097) );
  NAND U28547 ( .A(n27098), .B(n27097), .Z(n27366) );
  NAND U28548 ( .A(n27100), .B(n27099), .Z(n27104) );
  NAND U28549 ( .A(n27102), .B(n27101), .Z(n27103) );
  NAND U28550 ( .A(n27104), .B(n27103), .Z(n27364) );
  AND U28551 ( .A(n27106), .B(n27105), .Z(n27110) );
  NAND U28552 ( .A(n27108), .B(n27107), .Z(n27109) );
  NANDN U28553 ( .A(n27110), .B(n27109), .Z(n27262) );
  NAND U28554 ( .A(n27112), .B(n27111), .Z(n27116) );
  NAND U28555 ( .A(n27114), .B(n27113), .Z(n27115) );
  NAND U28556 ( .A(n27116), .B(n27115), .Z(n27261) );
  XOR U28557 ( .A(n27262), .B(n27261), .Z(n27263) );
  AND U28558 ( .A(n27118), .B(n27117), .Z(n27122) );
  NANDN U28559 ( .A(n27120), .B(n27119), .Z(n27121) );
  NANDN U28560 ( .A(n27122), .B(n27121), .Z(n27275) );
  AND U28561 ( .A(x[480]), .B(y[7963]), .Z(n27344) );
  AND U28562 ( .A(x[507]), .B(y[7936]), .Z(n27343) );
  XOR U28563 ( .A(n27344), .B(n27343), .Z(n27346) );
  AND U28564 ( .A(x[506]), .B(y[7937]), .Z(n27355) );
  XOR U28565 ( .A(n27355), .B(o[283]), .Z(n27345) );
  XOR U28566 ( .A(n27346), .B(n27345), .Z(n27274) );
  AND U28567 ( .A(x[489]), .B(y[7954]), .Z(n27350) );
  AND U28568 ( .A(x[501]), .B(y[7942]), .Z(n27349) );
  XOR U28569 ( .A(n27350), .B(n27349), .Z(n27352) );
  AND U28570 ( .A(x[498]), .B(y[7945]), .Z(n27351) );
  XOR U28571 ( .A(n27352), .B(n27351), .Z(n27273) );
  XOR U28572 ( .A(n27274), .B(n27273), .Z(n27276) );
  XNOR U28573 ( .A(n27275), .B(n27276), .Z(n27264) );
  XOR U28574 ( .A(n27364), .B(n27365), .Z(n27367) );
  XOR U28575 ( .A(n27366), .B(n27367), .Z(n27385) );
  NAND U28576 ( .A(n27124), .B(n27123), .Z(n27128) );
  NAND U28577 ( .A(n27126), .B(n27125), .Z(n27127) );
  AND U28578 ( .A(n27128), .B(n27127), .Z(n27383) );
  NAND U28579 ( .A(n27130), .B(n27129), .Z(n27134) );
  NAND U28580 ( .A(n27132), .B(n27131), .Z(n27133) );
  AND U28581 ( .A(n27134), .B(n27133), .Z(n27382) );
  XOR U28582 ( .A(n27383), .B(n27382), .Z(n27384) );
  NAND U28583 ( .A(n27136), .B(n27135), .Z(n27140) );
  NAND U28584 ( .A(n27138), .B(n27137), .Z(n27139) );
  AND U28585 ( .A(n27140), .B(n27139), .Z(n27370) );
  NAND U28586 ( .A(n27142), .B(n27141), .Z(n27146) );
  NAND U28587 ( .A(n27144), .B(n27143), .Z(n27145) );
  NAND U28588 ( .A(n27146), .B(n27145), .Z(n27360) );
  NAND U28589 ( .A(n27148), .B(n27147), .Z(n27152) );
  NAND U28590 ( .A(n27150), .B(n27149), .Z(n27151) );
  NAND U28591 ( .A(n27152), .B(n27151), .Z(n27358) );
  AND U28592 ( .A(x[499]), .B(y[7944]), .Z(n27332) );
  AND U28593 ( .A(x[505]), .B(y[7938]), .Z(n27331) );
  XOR U28594 ( .A(n27332), .B(n27331), .Z(n27334) );
  AND U28595 ( .A(x[486]), .B(y[7957]), .Z(n27333) );
  XOR U28596 ( .A(n27334), .B(n27333), .Z(n27321) );
  AND U28597 ( .A(x[495]), .B(y[7948]), .Z(n27297) );
  AND U28598 ( .A(x[482]), .B(y[7961]), .Z(n27296) );
  XOR U28599 ( .A(n27297), .B(n27296), .Z(n27299) );
  AND U28600 ( .A(x[483]), .B(y[7960]), .Z(n27298) );
  XOR U28601 ( .A(n27299), .B(n27298), .Z(n27320) );
  XOR U28602 ( .A(n27321), .B(n27320), .Z(n27322) );
  NAND U28603 ( .A(x[496]), .B(y[7947]), .Z(n27279) );
  XOR U28604 ( .A(n27279), .B(n27153), .Z(n27282) );
  XOR U28605 ( .A(n27281), .B(n27282), .Z(n27293) );
  AND U28606 ( .A(y[7950]), .B(x[493]), .Z(n27155) );
  AND U28607 ( .A(y[7951]), .B(x[492]), .Z(n27154) );
  XOR U28608 ( .A(n27155), .B(n27154), .Z(n27292) );
  XNOR U28609 ( .A(n27322), .B(n27323), .Z(n27258) );
  AND U28610 ( .A(n27291), .B(n27156), .Z(n27160) );
  NAND U28611 ( .A(n27158), .B(n27157), .Z(n27159) );
  NANDN U28612 ( .A(n27160), .B(n27159), .Z(n27256) );
  NAND U28613 ( .A(n27162), .B(n27161), .Z(n27166) );
  NAND U28614 ( .A(n27164), .B(n27163), .Z(n27165) );
  NAND U28615 ( .A(n27166), .B(n27165), .Z(n27255) );
  XOR U28616 ( .A(n27256), .B(n27255), .Z(n27257) );
  XOR U28617 ( .A(n27258), .B(n27257), .Z(n27359) );
  XNOR U28618 ( .A(n27358), .B(n27359), .Z(n27361) );
  XNOR U28619 ( .A(n27370), .B(n27371), .Z(n27373) );
  NAND U28620 ( .A(n27168), .B(n27167), .Z(n27172) );
  NAND U28621 ( .A(n27170), .B(n27169), .Z(n27171) );
  AND U28622 ( .A(n27172), .B(n27171), .Z(n27372) );
  XOR U28623 ( .A(n27373), .B(n27372), .Z(n27237) );
  XNOR U28624 ( .A(n27238), .B(n27237), .Z(n27240) );
  XOR U28625 ( .A(n27239), .B(n27240), .Z(n27245) );
  NAND U28626 ( .A(n27174), .B(n27173), .Z(n27178) );
  NAND U28627 ( .A(n27176), .B(n27175), .Z(n27177) );
  NAND U28628 ( .A(n27178), .B(n27177), .Z(n27244) );
  NANDN U28629 ( .A(n27180), .B(n27179), .Z(n27184) );
  NANDN U28630 ( .A(n27182), .B(n27181), .Z(n27183) );
  NAND U28631 ( .A(n27184), .B(n27183), .Z(n27249) );
  NAND U28632 ( .A(n27186), .B(n27185), .Z(n27190) );
  NAND U28633 ( .A(n27188), .B(n27187), .Z(n27189) );
  AND U28634 ( .A(n27190), .B(n27189), .Z(n27378) );
  NANDN U28635 ( .A(n27192), .B(n27191), .Z(n27196) );
  NAND U28636 ( .A(n27194), .B(n27193), .Z(n27195) );
  NAND U28637 ( .A(n27196), .B(n27195), .Z(n27316) );
  AND U28638 ( .A(y[7939]), .B(x[504]), .Z(n27198) );
  NAND U28639 ( .A(y[7943]), .B(x[500]), .Z(n27197) );
  XNOR U28640 ( .A(n27198), .B(n27197), .Z(n27328) );
  AND U28641 ( .A(x[487]), .B(y[7956]), .Z(n27327) );
  XOR U28642 ( .A(n27328), .B(n27327), .Z(n27315) );
  AND U28643 ( .A(x[488]), .B(y[7955]), .Z(n27286) );
  AND U28644 ( .A(x[503]), .B(y[7940]), .Z(n27285) );
  XOR U28645 ( .A(n27286), .B(n27285), .Z(n27288) );
  AND U28646 ( .A(x[502]), .B(y[7941]), .Z(n27287) );
  XOR U28647 ( .A(n27288), .B(n27287), .Z(n27314) );
  XOR U28648 ( .A(n27315), .B(n27314), .Z(n27317) );
  XOR U28649 ( .A(n27316), .B(n27317), .Z(n27377) );
  ANDN U28650 ( .B(n27200), .A(n27199), .Z(n27204) );
  NANDN U28651 ( .A(n27202), .B(n27201), .Z(n27203) );
  NANDN U28652 ( .A(n27204), .B(n27203), .Z(n27309) );
  NANDN U28653 ( .A(n27206), .B(n27205), .Z(n27210) );
  NANDN U28654 ( .A(n27208), .B(n27207), .Z(n27209) );
  NAND U28655 ( .A(n27210), .B(n27209), .Z(n27308) );
  XOR U28656 ( .A(n27309), .B(n27308), .Z(n27310) );
  AND U28657 ( .A(y[7956]), .B(x[488]), .Z(n27357) );
  NAND U28658 ( .A(n27357), .B(n27211), .Z(n27215) );
  NAND U28659 ( .A(n27213), .B(n27212), .Z(n27214) );
  NAND U28660 ( .A(n27215), .B(n27214), .Z(n27269) );
  AND U28661 ( .A(x[494]), .B(y[7949]), .Z(n27303) );
  AND U28662 ( .A(x[481]), .B(y[7962]), .Z(n27302) );
  XOR U28663 ( .A(n27303), .B(n27302), .Z(n27305) );
  ANDN U28664 ( .B(o[282]), .A(n27216), .Z(n27304) );
  XOR U28665 ( .A(n27305), .B(n27304), .Z(n27268) );
  AND U28666 ( .A(x[497]), .B(y[7946]), .Z(n27338) );
  AND U28667 ( .A(x[484]), .B(y[7959]), .Z(n27337) );
  XOR U28668 ( .A(n27338), .B(n27337), .Z(n27340) );
  AND U28669 ( .A(x[485]), .B(y[7958]), .Z(n27339) );
  XOR U28670 ( .A(n27340), .B(n27339), .Z(n27267) );
  XOR U28671 ( .A(n27268), .B(n27267), .Z(n27270) );
  XOR U28672 ( .A(n27269), .B(n27270), .Z(n27311) );
  XNOR U28673 ( .A(n27310), .B(n27311), .Z(n27376) );
  XNOR U28674 ( .A(n27378), .B(n27379), .Z(n27250) );
  XOR U28675 ( .A(n27249), .B(n27250), .Z(n27252) );
  NANDN U28676 ( .A(n27218), .B(n27217), .Z(n27222) );
  NANDN U28677 ( .A(n27220), .B(n27219), .Z(n27221) );
  AND U28678 ( .A(n27222), .B(n27221), .Z(n27251) );
  XOR U28679 ( .A(n27252), .B(n27251), .Z(n27243) );
  XOR U28680 ( .A(n27244), .B(n27243), .Z(n27246) );
  XOR U28681 ( .A(n27245), .B(n27246), .Z(n27224) );
  XOR U28682 ( .A(n27225), .B(n27224), .Z(n27226) );
  XOR U28683 ( .A(n27227), .B(n27226), .Z(n27233) );
  XNOR U28684 ( .A(n27232), .B(n27233), .Z(n27223) );
  XOR U28685 ( .A(n27230), .B(n27223), .Z(N572) );
  NAND U28686 ( .A(n27225), .B(n27224), .Z(n27229) );
  NAND U28687 ( .A(n27227), .B(n27226), .Z(n27228) );
  NAND U28688 ( .A(n27229), .B(n27228), .Z(n27554) );
  IV U28689 ( .A(n27554), .Z(n27552) );
  OR U28690 ( .A(n27232), .B(n27230), .Z(n27236) );
  ANDN U28691 ( .B(n27232), .A(n27231), .Z(n27234) );
  OR U28692 ( .A(n27234), .B(n27233), .Z(n27235) );
  AND U28693 ( .A(n27236), .B(n27235), .Z(n27553) );
  NAND U28694 ( .A(n27238), .B(n27237), .Z(n27242) );
  NANDN U28695 ( .A(n27240), .B(n27239), .Z(n27241) );
  NAND U28696 ( .A(n27242), .B(n27241), .Z(n27547) );
  NAND U28697 ( .A(n27244), .B(n27243), .Z(n27248) );
  NAND U28698 ( .A(n27246), .B(n27245), .Z(n27247) );
  AND U28699 ( .A(n27248), .B(n27247), .Z(n27546) );
  XOR U28700 ( .A(n27547), .B(n27546), .Z(n27549) );
  NAND U28701 ( .A(n27250), .B(n27249), .Z(n27254) );
  NAND U28702 ( .A(n27252), .B(n27251), .Z(n27253) );
  AND U28703 ( .A(n27254), .B(n27253), .Z(n27389) );
  NAND U28704 ( .A(n27256), .B(n27255), .Z(n27260) );
  NAND U28705 ( .A(n27258), .B(n27257), .Z(n27259) );
  NAND U28706 ( .A(n27260), .B(n27259), .Z(n27413) );
  NAND U28707 ( .A(n27262), .B(n27261), .Z(n27266) );
  NANDN U28708 ( .A(n27264), .B(n27263), .Z(n27265) );
  NAND U28709 ( .A(n27266), .B(n27265), .Z(n27518) );
  NAND U28710 ( .A(n27268), .B(n27267), .Z(n27272) );
  NAND U28711 ( .A(n27270), .B(n27269), .Z(n27271) );
  NAND U28712 ( .A(n27272), .B(n27271), .Z(n27517) );
  NAND U28713 ( .A(n27274), .B(n27273), .Z(n27278) );
  NAND U28714 ( .A(n27276), .B(n27275), .Z(n27277) );
  NAND U28715 ( .A(n27278), .B(n27277), .Z(n27516) );
  XOR U28716 ( .A(n27517), .B(n27516), .Z(n27519) );
  XOR U28717 ( .A(n27518), .B(n27519), .Z(n27414) );
  XOR U28718 ( .A(n27413), .B(n27414), .Z(n27416) );
  NANDN U28719 ( .A(n27280), .B(n27279), .Z(n27284) );
  NAND U28720 ( .A(n27282), .B(n27281), .Z(n27283) );
  NAND U28721 ( .A(n27284), .B(n27283), .Z(n27480) );
  AND U28722 ( .A(x[487]), .B(y[7957]), .Z(n27461) );
  AND U28723 ( .A(x[492]), .B(y[7952]), .Z(n27460) );
  XOR U28724 ( .A(n27461), .B(n27460), .Z(n27463) );
  AND U28725 ( .A(x[491]), .B(y[7953]), .Z(n27462) );
  XOR U28726 ( .A(n27463), .B(n27462), .Z(n27479) );
  AND U28727 ( .A(x[507]), .B(y[7937]), .Z(n27477) );
  XOR U28728 ( .A(o[284]), .B(n27477), .Z(n27491) );
  AND U28729 ( .A(x[506]), .B(y[7938]), .Z(n27490) );
  XOR U28730 ( .A(n27491), .B(n27490), .Z(n27493) );
  AND U28731 ( .A(x[495]), .B(y[7949]), .Z(n27492) );
  XNOR U28732 ( .A(n27493), .B(n27492), .Z(n27478) );
  XOR U28733 ( .A(n27480), .B(n27481), .Z(n27523) );
  NAND U28734 ( .A(n27286), .B(n27285), .Z(n27290) );
  NAND U28735 ( .A(n27288), .B(n27287), .Z(n27289) );
  NAND U28736 ( .A(n27290), .B(n27289), .Z(n27500) );
  AND U28737 ( .A(x[497]), .B(y[7947]), .Z(n27426) );
  AND U28738 ( .A(x[502]), .B(y[7942]), .Z(n27425) );
  XOR U28739 ( .A(n27426), .B(n27425), .Z(n27428) );
  AND U28740 ( .A(x[484]), .B(y[7960]), .Z(n27427) );
  XOR U28741 ( .A(n27428), .B(n27427), .Z(n27499) );
  AND U28742 ( .A(x[486]), .B(y[7958]), .Z(n27665) );
  AND U28743 ( .A(x[499]), .B(y[7945]), .Z(n27466) );
  XOR U28744 ( .A(n27665), .B(n27466), .Z(n27468) );
  XOR U28745 ( .A(n27468), .B(n27467), .Z(n27498) );
  XOR U28746 ( .A(n27499), .B(n27498), .Z(n27501) );
  XOR U28747 ( .A(n27500), .B(n27501), .Z(n27522) );
  NAND U28748 ( .A(n27485), .B(n27291), .Z(n27295) );
  NANDN U28749 ( .A(n27293), .B(n27292), .Z(n27294) );
  NAND U28750 ( .A(n27295), .B(n27294), .Z(n27444) );
  NAND U28751 ( .A(n27297), .B(n27296), .Z(n27301) );
  NAND U28752 ( .A(n27299), .B(n27298), .Z(n27300) );
  NAND U28753 ( .A(n27301), .B(n27300), .Z(n27443) );
  NAND U28754 ( .A(n27303), .B(n27302), .Z(n27307) );
  NAND U28755 ( .A(n27305), .B(n27304), .Z(n27306) );
  NAND U28756 ( .A(n27307), .B(n27306), .Z(n27442) );
  XOR U28757 ( .A(n27443), .B(n27442), .Z(n27445) );
  XOR U28758 ( .A(n27444), .B(n27445), .Z(n27524) );
  XOR U28759 ( .A(n27525), .B(n27524), .Z(n27415) );
  XNOR U28760 ( .A(n27416), .B(n27415), .Z(n27410) );
  NAND U28761 ( .A(n27309), .B(n27308), .Z(n27313) );
  NAND U28762 ( .A(n27311), .B(n27310), .Z(n27312) );
  NAND U28763 ( .A(n27313), .B(n27312), .Z(n27506) );
  NAND U28764 ( .A(n27315), .B(n27314), .Z(n27319) );
  NAND U28765 ( .A(n27317), .B(n27316), .Z(n27318) );
  NAND U28766 ( .A(n27319), .B(n27318), .Z(n27505) );
  NAND U28767 ( .A(n27321), .B(n27320), .Z(n27325) );
  NANDN U28768 ( .A(n27323), .B(n27322), .Z(n27324) );
  NAND U28769 ( .A(n27325), .B(n27324), .Z(n27504) );
  XOR U28770 ( .A(n27505), .B(n27504), .Z(n27507) );
  XOR U28771 ( .A(n27506), .B(n27507), .Z(n27408) );
  AND U28772 ( .A(x[504]), .B(y[7943]), .Z(n27879) );
  AND U28773 ( .A(x[500]), .B(y[7939]), .Z(n27326) );
  NAND U28774 ( .A(n27879), .B(n27326), .Z(n27330) );
  NAND U28775 ( .A(n27328), .B(n27327), .Z(n27329) );
  NAND U28776 ( .A(n27330), .B(n27329), .Z(n27542) );
  AND U28777 ( .A(x[505]), .B(y[7939]), .Z(n27456) );
  XOR U28778 ( .A(n27457), .B(n27456), .Z(n27455) );
  AND U28779 ( .A(x[481]), .B(y[7963]), .Z(n27454) );
  XOR U28780 ( .A(n27455), .B(n27454), .Z(n27541) );
  AND U28781 ( .A(x[496]), .B(y[7948]), .Z(n27449) );
  AND U28782 ( .A(x[504]), .B(y[7940]), .Z(n27448) );
  XOR U28783 ( .A(n27449), .B(n27448), .Z(n27451) );
  AND U28784 ( .A(x[482]), .B(y[7962]), .Z(n27450) );
  XOR U28785 ( .A(n27451), .B(n27450), .Z(n27540) );
  XOR U28786 ( .A(n27541), .B(n27540), .Z(n27543) );
  XOR U28787 ( .A(n27542), .B(n27543), .Z(n27513) );
  NAND U28788 ( .A(n27332), .B(n27331), .Z(n27336) );
  NAND U28789 ( .A(n27334), .B(n27333), .Z(n27335) );
  NAND U28790 ( .A(n27336), .B(n27335), .Z(n27536) );
  AND U28791 ( .A(x[483]), .B(y[7961]), .Z(n27484) );
  XOR U28792 ( .A(n27485), .B(n27484), .Z(n27487) );
  AND U28793 ( .A(x[503]), .B(y[7941]), .Z(n27486) );
  XOR U28794 ( .A(n27487), .B(n27486), .Z(n27535) );
  AND U28795 ( .A(x[485]), .B(y[7959]), .Z(n27472) );
  AND U28796 ( .A(x[501]), .B(y[7943]), .Z(n27471) );
  XOR U28797 ( .A(n27472), .B(n27471), .Z(n27474) );
  AND U28798 ( .A(x[500]), .B(y[7944]), .Z(n27473) );
  XOR U28799 ( .A(n27474), .B(n27473), .Z(n27534) );
  XOR U28800 ( .A(n27535), .B(n27534), .Z(n27537) );
  XOR U28801 ( .A(n27536), .B(n27537), .Z(n27511) );
  NAND U28802 ( .A(n27338), .B(n27337), .Z(n27342) );
  NAND U28803 ( .A(n27340), .B(n27339), .Z(n27341) );
  NAND U28804 ( .A(n27342), .B(n27341), .Z(n27529) );
  NAND U28805 ( .A(n27344), .B(n27343), .Z(n27348) );
  NAND U28806 ( .A(n27346), .B(n27345), .Z(n27347) );
  NAND U28807 ( .A(n27348), .B(n27347), .Z(n27528) );
  XOR U28808 ( .A(n27529), .B(n27528), .Z(n27531) );
  NAND U28809 ( .A(n27350), .B(n27349), .Z(n27354) );
  NAND U28810 ( .A(n27352), .B(n27351), .Z(n27353) );
  NAND U28811 ( .A(n27354), .B(n27353), .Z(n27421) );
  AND U28812 ( .A(n27355), .B(o[283]), .Z(n27434) );
  AND U28813 ( .A(x[480]), .B(y[7964]), .Z(n27432) );
  AND U28814 ( .A(x[508]), .B(y[7936]), .Z(n27431) );
  XOR U28815 ( .A(n27432), .B(n27431), .Z(n27433) );
  XOR U28816 ( .A(n27434), .B(n27433), .Z(n27420) );
  NAND U28817 ( .A(y[7954]), .B(x[490]), .Z(n27356) );
  XNOR U28818 ( .A(n27357), .B(n27356), .Z(n27439) );
  AND U28819 ( .A(x[489]), .B(y[7955]), .Z(n27438) );
  XOR U28820 ( .A(n27439), .B(n27438), .Z(n27419) );
  XOR U28821 ( .A(n27420), .B(n27419), .Z(n27422) );
  XOR U28822 ( .A(n27421), .B(n27422), .Z(n27530) );
  XNOR U28823 ( .A(n27531), .B(n27530), .Z(n27510) );
  XNOR U28824 ( .A(n27410), .B(n27409), .Z(n27403) );
  NAND U28825 ( .A(n27359), .B(n27358), .Z(n27363) );
  NANDN U28826 ( .A(n27361), .B(n27360), .Z(n27362) );
  NAND U28827 ( .A(n27363), .B(n27362), .Z(n27402) );
  NAND U28828 ( .A(n27365), .B(n27364), .Z(n27369) );
  NAND U28829 ( .A(n27367), .B(n27366), .Z(n27368) );
  NAND U28830 ( .A(n27369), .B(n27368), .Z(n27401) );
  XNOR U28831 ( .A(n27402), .B(n27401), .Z(n27404) );
  XNOR U28832 ( .A(n27389), .B(n27390), .Z(n27391) );
  NANDN U28833 ( .A(n27371), .B(n27370), .Z(n27375) );
  NAND U28834 ( .A(n27373), .B(n27372), .Z(n27374) );
  NAND U28835 ( .A(n27375), .B(n27374), .Z(n27397) );
  NANDN U28836 ( .A(n27377), .B(n27376), .Z(n27381) );
  NANDN U28837 ( .A(n27379), .B(n27378), .Z(n27380) );
  AND U28838 ( .A(n27381), .B(n27380), .Z(n27396) );
  NAND U28839 ( .A(n27383), .B(n27382), .Z(n27387) );
  NANDN U28840 ( .A(n27385), .B(n27384), .Z(n27386) );
  AND U28841 ( .A(n27387), .B(n27386), .Z(n27395) );
  XOR U28842 ( .A(n27396), .B(n27395), .Z(n27398) );
  XNOR U28843 ( .A(n27397), .B(n27398), .Z(n27392) );
  XOR U28844 ( .A(n27549), .B(n27548), .Z(n27555) );
  XNOR U28845 ( .A(n27553), .B(n27555), .Z(n27388) );
  XOR U28846 ( .A(n27552), .B(n27388), .Z(N573) );
  NANDN U28847 ( .A(n27390), .B(n27389), .Z(n27394) );
  NANDN U28848 ( .A(n27392), .B(n27391), .Z(n27393) );
  NAND U28849 ( .A(n27394), .B(n27393), .Z(n27565) );
  NAND U28850 ( .A(n27396), .B(n27395), .Z(n27400) );
  NAND U28851 ( .A(n27398), .B(n27397), .Z(n27399) );
  NAND U28852 ( .A(n27400), .B(n27399), .Z(n27563) );
  NAND U28853 ( .A(n27402), .B(n27401), .Z(n27406) );
  NANDN U28854 ( .A(n27404), .B(n27403), .Z(n27405) );
  NAND U28855 ( .A(n27406), .B(n27405), .Z(n27569) );
  NANDN U28856 ( .A(n27408), .B(n27407), .Z(n27412) );
  NAND U28857 ( .A(n27410), .B(n27409), .Z(n27411) );
  AND U28858 ( .A(n27412), .B(n27411), .Z(n27570) );
  XOR U28859 ( .A(n27569), .B(n27570), .Z(n27572) );
  NAND U28860 ( .A(n27414), .B(n27413), .Z(n27418) );
  NAND U28861 ( .A(n27416), .B(n27415), .Z(n27417) );
  NAND U28862 ( .A(n27418), .B(n27417), .Z(n27587) );
  NAND U28863 ( .A(n27420), .B(n27419), .Z(n27424) );
  NAND U28864 ( .A(n27422), .B(n27421), .Z(n27423) );
  AND U28865 ( .A(n27424), .B(n27423), .Z(n27691) );
  NAND U28866 ( .A(n27426), .B(n27425), .Z(n27430) );
  NAND U28867 ( .A(n27428), .B(n27427), .Z(n27429) );
  NAND U28868 ( .A(n27430), .B(n27429), .Z(n27729) );
  NAND U28869 ( .A(n27432), .B(n27431), .Z(n27436) );
  NAND U28870 ( .A(n27434), .B(n27433), .Z(n27435) );
  NAND U28871 ( .A(n27436), .B(n27435), .Z(n27728) );
  XOR U28872 ( .A(n27729), .B(n27728), .Z(n27730) );
  AND U28873 ( .A(y[7956]), .B(x[490]), .Z(n27726) );
  NAND U28874 ( .A(n27726), .B(n27437), .Z(n27441) );
  NAND U28875 ( .A(n27439), .B(n27438), .Z(n27440) );
  NAND U28876 ( .A(n27441), .B(n27440), .Z(n27699) );
  AND U28877 ( .A(x[502]), .B(y[7943]), .Z(n27643) );
  AND U28878 ( .A(x[492]), .B(y[7953]), .Z(n27864) );
  AND U28879 ( .A(x[481]), .B(y[7964]), .Z(n27641) );
  XOR U28880 ( .A(n27864), .B(n27641), .Z(n27642) );
  XOR U28881 ( .A(n27643), .B(n27642), .Z(n27698) );
  AND U28882 ( .A(x[495]), .B(y[7950]), .Z(n27646) );
  XOR U28883 ( .A(n27698), .B(n27697), .Z(n27700) );
  XNOR U28884 ( .A(n27699), .B(n27700), .Z(n27731) );
  NAND U28885 ( .A(n27443), .B(n27442), .Z(n27447) );
  NAND U28886 ( .A(n27445), .B(n27444), .Z(n27446) );
  AND U28887 ( .A(n27447), .B(n27446), .Z(n27693) );
  XOR U28888 ( .A(n27694), .B(n27693), .Z(n27688) );
  NAND U28889 ( .A(n27449), .B(n27448), .Z(n27453) );
  NAND U28890 ( .A(n27451), .B(n27450), .Z(n27452) );
  NAND U28891 ( .A(n27453), .B(n27452), .Z(n27704) );
  AND U28892 ( .A(n27455), .B(n27454), .Z(n27459) );
  NAND U28893 ( .A(n27457), .B(n27456), .Z(n27458) );
  NANDN U28894 ( .A(n27459), .B(n27458), .Z(n27703) );
  XOR U28895 ( .A(n27704), .B(n27703), .Z(n27705) );
  NAND U28896 ( .A(n27461), .B(n27460), .Z(n27465) );
  NAND U28897 ( .A(n27463), .B(n27462), .Z(n27464) );
  NAND U28898 ( .A(n27465), .B(n27464), .Z(n27607) );
  AND U28899 ( .A(x[491]), .B(y[7954]), .Z(n27662) );
  AND U28900 ( .A(x[483]), .B(y[7962]), .Z(n27660) );
  AND U28901 ( .A(x[497]), .B(y[7948]), .Z(n27659) );
  XOR U28902 ( .A(n27660), .B(n27659), .Z(n27661) );
  XOR U28903 ( .A(n27662), .B(n27661), .Z(n27606) );
  AND U28904 ( .A(x[503]), .B(y[7942]), .Z(n27656) );
  AND U28905 ( .A(x[493]), .B(y[7952]), .Z(n27654) );
  AND U28906 ( .A(x[504]), .B(y[7941]), .Z(n27811) );
  XOR U28907 ( .A(n27654), .B(n27811), .Z(n27655) );
  XOR U28908 ( .A(n27656), .B(n27655), .Z(n27605) );
  XOR U28909 ( .A(n27606), .B(n27605), .Z(n27608) );
  XNOR U28910 ( .A(n27607), .B(n27608), .Z(n27706) );
  NAND U28911 ( .A(n27665), .B(n27466), .Z(n27470) );
  NAND U28912 ( .A(n27468), .B(n27467), .Z(n27469) );
  NAND U28913 ( .A(n27470), .B(n27469), .Z(n27712) );
  AND U28914 ( .A(x[505]), .B(y[7940]), .Z(n27638) );
  AND U28915 ( .A(x[506]), .B(y[7939]), .Z(n27635) );
  XOR U28916 ( .A(n27636), .B(n27635), .Z(n27637) );
  XOR U28917 ( .A(n27638), .B(n27637), .Z(n27710) );
  AND U28918 ( .A(x[508]), .B(y[7937]), .Z(n27653) );
  XOR U28919 ( .A(o[285]), .B(n27653), .Z(n27721) );
  AND U28920 ( .A(x[480]), .B(y[7965]), .Z(n27719) );
  AND U28921 ( .A(x[509]), .B(y[7936]), .Z(n27718) );
  XOR U28922 ( .A(n27719), .B(n27718), .Z(n27720) );
  XNOR U28923 ( .A(n27721), .B(n27720), .Z(n27709) );
  XOR U28924 ( .A(n27712), .B(n27711), .Z(n27593) );
  NAND U28925 ( .A(n27472), .B(n27471), .Z(n27476) );
  NAND U28926 ( .A(n27474), .B(n27473), .Z(n27475) );
  NAND U28927 ( .A(n27476), .B(n27475), .Z(n27674) );
  AND U28928 ( .A(n27477), .B(o[284]), .Z(n27614) );
  AND U28929 ( .A(x[496]), .B(y[7949]), .Z(n27612) );
  AND U28930 ( .A(x[507]), .B(y[7938]), .Z(n27611) );
  XOR U28931 ( .A(n27612), .B(n27611), .Z(n27613) );
  XOR U28932 ( .A(n27614), .B(n27613), .Z(n27673) );
  AND U28933 ( .A(x[482]), .B(y[7963]), .Z(n27623) );
  XOR U28934 ( .A(n27626), .B(n27625), .Z(n27672) );
  XOR U28935 ( .A(n27673), .B(n27672), .Z(n27675) );
  XOR U28936 ( .A(n27674), .B(n27675), .Z(n27594) );
  NANDN U28937 ( .A(n27479), .B(n27478), .Z(n27483) );
  NAND U28938 ( .A(n27481), .B(n27480), .Z(n27482) );
  NAND U28939 ( .A(n27483), .B(n27482), .Z(n27599) );
  NAND U28940 ( .A(n27485), .B(n27484), .Z(n27489) );
  NAND U28941 ( .A(n27487), .B(n27486), .Z(n27488) );
  NAND U28942 ( .A(n27489), .B(n27488), .Z(n27630) );
  NAND U28943 ( .A(n27491), .B(n27490), .Z(n27495) );
  NAND U28944 ( .A(n27493), .B(n27492), .Z(n27494) );
  NAND U28945 ( .A(n27495), .B(n27494), .Z(n27629) );
  XOR U28946 ( .A(n27630), .B(n27629), .Z(n27631) );
  AND U28947 ( .A(x[488]), .B(y[7957]), .Z(n27667) );
  AND U28948 ( .A(y[7959]), .B(x[486]), .Z(n27497) );
  NAND U28949 ( .A(y[7958]), .B(x[487]), .Z(n27496) );
  XNOR U28950 ( .A(n27497), .B(n27496), .Z(n27666) );
  XNOR U28951 ( .A(n27667), .B(n27666), .Z(n27716) );
  AND U28952 ( .A(x[485]), .B(y[7960]), .Z(n27620) );
  AND U28953 ( .A(x[484]), .B(y[7961]), .Z(n27618) );
  AND U28954 ( .A(x[490]), .B(y[7955]), .Z(n27617) );
  XOR U28955 ( .A(n27618), .B(n27617), .Z(n27619) );
  XOR U28956 ( .A(n27620), .B(n27619), .Z(n27717) );
  NAND U28957 ( .A(x[489]), .B(y[7956]), .Z(n27873) );
  IV U28958 ( .A(n27873), .Z(n27715) );
  XNOR U28959 ( .A(n27601), .B(n27602), .Z(n27686) );
  NAND U28960 ( .A(n27499), .B(n27498), .Z(n27503) );
  NAND U28961 ( .A(n27501), .B(n27500), .Z(n27502) );
  NAND U28962 ( .A(n27503), .B(n27502), .Z(n27685) );
  XOR U28963 ( .A(n27587), .B(n27588), .Z(n27590) );
  NAND U28964 ( .A(n27505), .B(n27504), .Z(n27509) );
  NAND U28965 ( .A(n27507), .B(n27506), .Z(n27508) );
  NAND U28966 ( .A(n27509), .B(n27508), .Z(n27581) );
  NANDN U28967 ( .A(n27511), .B(n27510), .Z(n27515) );
  NANDN U28968 ( .A(n27513), .B(n27512), .Z(n27514) );
  AND U28969 ( .A(n27515), .B(n27514), .Z(n27582) );
  XOR U28970 ( .A(n27581), .B(n27582), .Z(n27584) );
  NAND U28971 ( .A(n27517), .B(n27516), .Z(n27521) );
  NAND U28972 ( .A(n27519), .B(n27518), .Z(n27520) );
  NAND U28973 ( .A(n27521), .B(n27520), .Z(n27577) );
  NANDN U28974 ( .A(n27523), .B(n27522), .Z(n27527) );
  NAND U28975 ( .A(n27525), .B(n27524), .Z(n27526) );
  NAND U28976 ( .A(n27527), .B(n27526), .Z(n27575) );
  NAND U28977 ( .A(n27529), .B(n27528), .Z(n27533) );
  NAND U28978 ( .A(n27531), .B(n27530), .Z(n27532) );
  NAND U28979 ( .A(n27533), .B(n27532), .Z(n27680) );
  NAND U28980 ( .A(n27535), .B(n27534), .Z(n27539) );
  NAND U28981 ( .A(n27537), .B(n27536), .Z(n27538) );
  NAND U28982 ( .A(n27539), .B(n27538), .Z(n27679) );
  NAND U28983 ( .A(n27541), .B(n27540), .Z(n27545) );
  NAND U28984 ( .A(n27543), .B(n27542), .Z(n27544) );
  NAND U28985 ( .A(n27545), .B(n27544), .Z(n27678) );
  XOR U28986 ( .A(n27679), .B(n27678), .Z(n27681) );
  XOR U28987 ( .A(n27680), .B(n27681), .Z(n27576) );
  XOR U28988 ( .A(n27575), .B(n27576), .Z(n27578) );
  XOR U28989 ( .A(n27577), .B(n27578), .Z(n27583) );
  XOR U28990 ( .A(n27584), .B(n27583), .Z(n27589) );
  XOR U28991 ( .A(n27590), .B(n27589), .Z(n27571) );
  XOR U28992 ( .A(n27572), .B(n27571), .Z(n27564) );
  XNOR U28993 ( .A(n27563), .B(n27564), .Z(n27566) );
  XOR U28994 ( .A(n27565), .B(n27566), .Z(n27562) );
  NAND U28995 ( .A(n27547), .B(n27546), .Z(n27551) );
  NAND U28996 ( .A(n27549), .B(n27548), .Z(n27550) );
  NAND U28997 ( .A(n27551), .B(n27550), .Z(n27561) );
  NANDN U28998 ( .A(n27552), .B(n27553), .Z(n27558) );
  NOR U28999 ( .A(n27554), .B(n27553), .Z(n27556) );
  OR U29000 ( .A(n27556), .B(n27555), .Z(n27557) );
  AND U29001 ( .A(n27558), .B(n27557), .Z(n27560) );
  XOR U29002 ( .A(n27561), .B(n27560), .Z(n27559) );
  XNOR U29003 ( .A(n27562), .B(n27559), .Z(N574) );
  NAND U29004 ( .A(n27564), .B(n27563), .Z(n27568) );
  NANDN U29005 ( .A(n27566), .B(n27565), .Z(n27567) );
  NAND U29006 ( .A(n27568), .B(n27567), .Z(n27737) );
  NAND U29007 ( .A(n27570), .B(n27569), .Z(n27574) );
  NAND U29008 ( .A(n27572), .B(n27571), .Z(n27573) );
  NAND U29009 ( .A(n27574), .B(n27573), .Z(n28023) );
  NAND U29010 ( .A(n27576), .B(n27575), .Z(n27580) );
  NAND U29011 ( .A(n27578), .B(n27577), .Z(n27579) );
  AND U29012 ( .A(n27580), .B(n27579), .Z(n28029) );
  NAND U29013 ( .A(n27582), .B(n27581), .Z(n27586) );
  NAND U29014 ( .A(n27584), .B(n27583), .Z(n27585) );
  AND U29015 ( .A(n27586), .B(n27585), .Z(n28027) );
  NAND U29016 ( .A(n27588), .B(n27587), .Z(n27592) );
  NAND U29017 ( .A(n27590), .B(n27589), .Z(n27591) );
  AND U29018 ( .A(n27592), .B(n27591), .Z(n28026) );
  XOR U29019 ( .A(n28027), .B(n28026), .Z(n28028) );
  XOR U29020 ( .A(n28029), .B(n28028), .Z(n28020) );
  NANDN U29021 ( .A(n27594), .B(n27593), .Z(n27598) );
  NANDN U29022 ( .A(n27596), .B(n27595), .Z(n27597) );
  AND U29023 ( .A(n27598), .B(n27597), .Z(n28009) );
  NANDN U29024 ( .A(n27600), .B(n27599), .Z(n27604) );
  NANDN U29025 ( .A(n27602), .B(n27601), .Z(n27603) );
  AND U29026 ( .A(n27604), .B(n27603), .Z(n28000) );
  NAND U29027 ( .A(n27606), .B(n27605), .Z(n27610) );
  NAND U29028 ( .A(n27608), .B(n27607), .Z(n27609) );
  AND U29029 ( .A(n27610), .B(n27609), .Z(n27984) );
  NAND U29030 ( .A(n27612), .B(n27611), .Z(n27616) );
  NAND U29031 ( .A(n27614), .B(n27613), .Z(n27615) );
  NAND U29032 ( .A(n27616), .B(n27615), .Z(n27942) );
  NAND U29033 ( .A(n27618), .B(n27617), .Z(n27622) );
  NAND U29034 ( .A(n27620), .B(n27619), .Z(n27621) );
  NAND U29035 ( .A(n27622), .B(n27621), .Z(n27945) );
  AND U29036 ( .A(x[486]), .B(y[7960]), .Z(n27798) );
  AND U29037 ( .A(x[485]), .B(y[7961]), .Z(n27800) );
  AND U29038 ( .A(x[499]), .B(y[7947]), .Z(n27799) );
  XOR U29039 ( .A(n27800), .B(n27799), .Z(n27797) );
  XNOR U29040 ( .A(n27798), .B(n27797), .Z(n27752) );
  AND U29041 ( .A(x[484]), .B(y[7962]), .Z(n27859) );
  AND U29042 ( .A(x[483]), .B(y[7963]), .Z(n27861) );
  AND U29043 ( .A(x[498]), .B(y[7948]), .Z(n27860) );
  XOR U29044 ( .A(n27861), .B(n27860), .Z(n27858) );
  XOR U29045 ( .A(n27859), .B(n27858), .Z(n27755) );
  NANDN U29046 ( .A(n27624), .B(n27623), .Z(n27628) );
  NAND U29047 ( .A(n27626), .B(n27625), .Z(n27627) );
  AND U29048 ( .A(n27628), .B(n27627), .Z(n27754) );
  XOR U29049 ( .A(n27752), .B(n27753), .Z(n27944) );
  XOR U29050 ( .A(n27945), .B(n27944), .Z(n27943) );
  XOR U29051 ( .A(n27942), .B(n27943), .Z(n27985) );
  NAND U29052 ( .A(n27630), .B(n27629), .Z(n27634) );
  NANDN U29053 ( .A(n27632), .B(n27631), .Z(n27633) );
  AND U29054 ( .A(n27634), .B(n27633), .Z(n27982) );
  XOR U29055 ( .A(n27983), .B(n27982), .Z(n28003) );
  AND U29056 ( .A(n27636), .B(n27635), .Z(n27640) );
  NAND U29057 ( .A(n27638), .B(n27637), .Z(n27639) );
  NANDN U29058 ( .A(n27640), .B(n27639), .Z(n27936) );
  AND U29059 ( .A(n27864), .B(n27641), .Z(n27645) );
  NAND U29060 ( .A(n27643), .B(n27642), .Z(n27644) );
  NANDN U29061 ( .A(n27645), .B(n27644), .Z(n27939) );
  NANDN U29062 ( .A(n27790), .B(n27646), .Z(n27650) );
  NANDN U29063 ( .A(n27648), .B(n27647), .Z(n27649) );
  AND U29064 ( .A(n27650), .B(n27649), .Z(n27773) );
  AND U29065 ( .A(x[503]), .B(y[7943]), .Z(n27810) );
  AND U29066 ( .A(y[7942]), .B(x[504]), .Z(n27652) );
  AND U29067 ( .A(y[7941]), .B(x[505]), .Z(n27651) );
  XOR U29068 ( .A(n27652), .B(n27651), .Z(n27809) );
  XOR U29069 ( .A(n27810), .B(n27809), .Z(n27775) );
  AND U29070 ( .A(n27653), .B(o[285]), .Z(n27843) );
  AND U29071 ( .A(x[508]), .B(y[7938]), .Z(n27841) );
  AND U29072 ( .A(x[496]), .B(y[7950]), .Z(n27840) );
  XOR U29073 ( .A(n27841), .B(n27840), .Z(n27842) );
  XNOR U29074 ( .A(n27843), .B(n27842), .Z(n27774) );
  XNOR U29075 ( .A(n27773), .B(n27772), .Z(n27938) );
  XOR U29076 ( .A(n27939), .B(n27938), .Z(n27937) );
  XOR U29077 ( .A(n27936), .B(n27937), .Z(n27741) );
  NAND U29078 ( .A(n27654), .B(n27811), .Z(n27658) );
  NAND U29079 ( .A(n27656), .B(n27655), .Z(n27657) );
  NAND U29080 ( .A(n27658), .B(n27657), .Z(n27967) );
  NAND U29081 ( .A(n27660), .B(n27659), .Z(n27664) );
  NAND U29082 ( .A(n27662), .B(n27661), .Z(n27663) );
  AND U29083 ( .A(n27664), .B(n27663), .Z(n27765) );
  AND U29084 ( .A(x[480]), .B(y[7966]), .Z(n27855) );
  AND U29085 ( .A(x[509]), .B(y[7937]), .Z(n27876) );
  XOR U29086 ( .A(o[286]), .B(n27876), .Z(n27853) );
  AND U29087 ( .A(x[510]), .B(y[7936]), .Z(n27852) );
  XOR U29088 ( .A(n27853), .B(n27852), .Z(n27854) );
  XOR U29089 ( .A(n27855), .B(n27854), .Z(n27767) );
  AND U29090 ( .A(x[500]), .B(y[7946]), .Z(n27834) );
  XOR U29091 ( .A(n27835), .B(n27834), .Z(n27837) );
  AND U29092 ( .A(x[488]), .B(y[7958]), .Z(n27836) );
  XNOR U29093 ( .A(n27837), .B(n27836), .Z(n27766) );
  XNOR U29094 ( .A(n27765), .B(n27764), .Z(n27966) );
  XOR U29095 ( .A(n27967), .B(n27966), .Z(n27964) );
  AND U29096 ( .A(x[487]), .B(y[7959]), .Z(n27792) );
  NAND U29097 ( .A(n27665), .B(n27792), .Z(n27669) );
  NAND U29098 ( .A(n27667), .B(n27666), .Z(n27668) );
  AND U29099 ( .A(n27669), .B(n27668), .Z(n27758) );
  AND U29100 ( .A(x[501]), .B(y[7945]), .Z(n27671) );
  AND U29101 ( .A(y[7944]), .B(x[502]), .Z(n27670) );
  XOR U29102 ( .A(n27671), .B(n27670), .Z(n27791) );
  XOR U29103 ( .A(n27792), .B(n27791), .Z(n27761) );
  AND U29104 ( .A(x[497]), .B(y[7949]), .Z(n27787) );
  AND U29105 ( .A(x[482]), .B(y[7964]), .Z(n27785) );
  AND U29106 ( .A(x[506]), .B(y[7940]), .Z(n27784) );
  XOR U29107 ( .A(n27785), .B(n27784), .Z(n27786) );
  XNOR U29108 ( .A(n27787), .B(n27786), .Z(n27760) );
  XNOR U29109 ( .A(n27758), .B(n27759), .Z(n27965) );
  NAND U29110 ( .A(n27673), .B(n27672), .Z(n27677) );
  NAND U29111 ( .A(n27675), .B(n27674), .Z(n27676) );
  NAND U29112 ( .A(n27677), .B(n27676), .Z(n27742) );
  XOR U29113 ( .A(n27743), .B(n27742), .Z(n27740) );
  XOR U29114 ( .A(n27741), .B(n27740), .Z(n28002) );
  XNOR U29115 ( .A(n28000), .B(n28001), .Z(n28011) );
  NAND U29116 ( .A(n27679), .B(n27678), .Z(n27683) );
  NAND U29117 ( .A(n27681), .B(n27680), .Z(n27682) );
  NAND U29118 ( .A(n27683), .B(n27682), .Z(n28008) );
  XOR U29119 ( .A(n28011), .B(n28008), .Z(n27684) );
  XOR U29120 ( .A(n28009), .B(n27684), .Z(n27995) );
  NANDN U29121 ( .A(n27686), .B(n27685), .Z(n27690) );
  NANDN U29122 ( .A(n27688), .B(n27687), .Z(n27689) );
  NAND U29123 ( .A(n27690), .B(n27689), .Z(n27996) );
  NANDN U29124 ( .A(n27692), .B(n27691), .Z(n27696) );
  NAND U29125 ( .A(n27694), .B(n27693), .Z(n27695) );
  AND U29126 ( .A(n27696), .B(n27695), .Z(n27976) );
  NAND U29127 ( .A(n27698), .B(n27697), .Z(n27702) );
  NAND U29128 ( .A(n27700), .B(n27699), .Z(n27701) );
  AND U29129 ( .A(n27702), .B(n27701), .Z(n27961) );
  NAND U29130 ( .A(n27704), .B(n27703), .Z(n27708) );
  NANDN U29131 ( .A(n27706), .B(n27705), .Z(n27707) );
  AND U29132 ( .A(n27708), .B(n27707), .Z(n27960) );
  XOR U29133 ( .A(n27961), .B(n27960), .Z(n27959) );
  NANDN U29134 ( .A(n27710), .B(n27709), .Z(n27714) );
  OR U29135 ( .A(n27712), .B(n27711), .Z(n27713) );
  NAND U29136 ( .A(n27714), .B(n27713), .Z(n27958) );
  XOR U29137 ( .A(n27959), .B(n27958), .Z(n27979) );
  NAND U29138 ( .A(n27719), .B(n27718), .Z(n27723) );
  NAND U29139 ( .A(n27721), .B(n27720), .Z(n27722) );
  NAND U29140 ( .A(n27723), .B(n27722), .Z(n27778) );
  AND U29141 ( .A(y[7954]), .B(x[492]), .Z(n27724) );
  XOR U29142 ( .A(n27725), .B(n27724), .Z(n27865) );
  XOR U29143 ( .A(n27866), .B(n27865), .Z(n27872) );
  AND U29144 ( .A(x[489]), .B(y[7957]), .Z(n27727) );
  XOR U29145 ( .A(n27727), .B(n27726), .Z(n27871) );
  XOR U29146 ( .A(n27872), .B(n27871), .Z(n27781) );
  AND U29147 ( .A(x[507]), .B(y[7939]), .Z(n27806) );
  AND U29148 ( .A(x[481]), .B(y[7965]), .Z(n27805) );
  XOR U29149 ( .A(n27806), .B(n27805), .Z(n27803) );
  XOR U29150 ( .A(n27804), .B(n27803), .Z(n27780) );
  XOR U29151 ( .A(n27781), .B(n27780), .Z(n27779) );
  XOR U29152 ( .A(n27778), .B(n27779), .Z(n27749) );
  NAND U29153 ( .A(n27729), .B(n27728), .Z(n27733) );
  NANDN U29154 ( .A(n27731), .B(n27730), .Z(n27732) );
  AND U29155 ( .A(n27733), .B(n27732), .Z(n27746) );
  XNOR U29156 ( .A(n27747), .B(n27746), .Z(n27978) );
  XNOR U29157 ( .A(n27976), .B(n27977), .Z(n27997) );
  XOR U29158 ( .A(n27996), .B(n27997), .Z(n27994) );
  XOR U29159 ( .A(n27995), .B(n27994), .Z(n28021) );
  XOR U29160 ( .A(n28023), .B(n28022), .Z(n27734) );
  XNOR U29161 ( .A(n27735), .B(n27734), .Z(N575) );
  NAND U29162 ( .A(n27735), .B(n27734), .Z(n27739) );
  NANDN U29163 ( .A(n27737), .B(n27736), .Z(n27738) );
  AND U29164 ( .A(n27739), .B(n27738), .Z(n28019) );
  NAND U29165 ( .A(n27741), .B(n27740), .Z(n27745) );
  NAND U29166 ( .A(n27743), .B(n27742), .Z(n27744) );
  AND U29167 ( .A(n27745), .B(n27744), .Z(n27993) );
  NAND U29168 ( .A(n27747), .B(n27746), .Z(n27751) );
  NANDN U29169 ( .A(n27749), .B(n27748), .Z(n27750) );
  AND U29170 ( .A(n27751), .B(n27750), .Z(n27975) );
  NANDN U29171 ( .A(n27753), .B(n27752), .Z(n27757) );
  NANDN U29172 ( .A(n27755), .B(n27754), .Z(n27756) );
  AND U29173 ( .A(n27757), .B(n27756), .Z(n27957) );
  NANDN U29174 ( .A(n27759), .B(n27758), .Z(n27763) );
  NANDN U29175 ( .A(n27761), .B(n27760), .Z(n27762) );
  AND U29176 ( .A(n27763), .B(n27762), .Z(n27771) );
  NAND U29177 ( .A(n27765), .B(n27764), .Z(n27769) );
  NANDN U29178 ( .A(n27767), .B(n27766), .Z(n27768) );
  NAND U29179 ( .A(n27769), .B(n27768), .Z(n27770) );
  XNOR U29180 ( .A(n27771), .B(n27770), .Z(n27955) );
  NAND U29181 ( .A(n27773), .B(n27772), .Z(n27777) );
  NANDN U29182 ( .A(n27775), .B(n27774), .Z(n27776) );
  AND U29183 ( .A(n27777), .B(n27776), .Z(n27953) );
  NAND U29184 ( .A(n27779), .B(n27778), .Z(n27783) );
  NAND U29185 ( .A(n27781), .B(n27780), .Z(n27782) );
  AND U29186 ( .A(n27783), .B(n27782), .Z(n27935) );
  AND U29187 ( .A(n27785), .B(n27784), .Z(n27789) );
  AND U29188 ( .A(n27787), .B(n27786), .Z(n27788) );
  NOR U29189 ( .A(n27789), .B(n27788), .Z(n27796) );
  AND U29190 ( .A(x[502]), .B(y[7945]), .Z(n27877) );
  NANDN U29191 ( .A(n27790), .B(n27877), .Z(n27794) );
  NAND U29192 ( .A(n27792), .B(n27791), .Z(n27793) );
  AND U29193 ( .A(n27794), .B(n27793), .Z(n27795) );
  XNOR U29194 ( .A(n27796), .B(n27795), .Z(n27851) );
  NAND U29195 ( .A(n27798), .B(n27797), .Z(n27802) );
  NAND U29196 ( .A(n27800), .B(n27799), .Z(n27801) );
  AND U29197 ( .A(n27802), .B(n27801), .Z(n27833) );
  NAND U29198 ( .A(n27804), .B(n27803), .Z(n27808) );
  NAND U29199 ( .A(n27806), .B(n27805), .Z(n27807) );
  AND U29200 ( .A(n27808), .B(n27807), .Z(n27815) );
  NAND U29201 ( .A(n27810), .B(n27809), .Z(n27813) );
  AND U29202 ( .A(x[505]), .B(y[7942]), .Z(n27878) );
  NAND U29203 ( .A(n27811), .B(n27878), .Z(n27812) );
  NAND U29204 ( .A(n27813), .B(n27812), .Z(n27814) );
  XNOR U29205 ( .A(n27815), .B(n27814), .Z(n27831) );
  AND U29206 ( .A(y[7955]), .B(x[492]), .Z(n27817) );
  NAND U29207 ( .A(y[7941]), .B(x[506]), .Z(n27816) );
  XNOR U29208 ( .A(n27817), .B(n27816), .Z(n27821) );
  AND U29209 ( .A(y[7956]), .B(x[491]), .Z(n27819) );
  NAND U29210 ( .A(y[7967]), .B(x[480]), .Z(n27818) );
  XNOR U29211 ( .A(n27819), .B(n27818), .Z(n27820) );
  XOR U29212 ( .A(n27821), .B(n27820), .Z(n27829) );
  AND U29213 ( .A(y[7953]), .B(x[494]), .Z(n27823) );
  NAND U29214 ( .A(y[7958]), .B(x[489]), .Z(n27822) );
  XNOR U29215 ( .A(n27823), .B(n27822), .Z(n27827) );
  AND U29216 ( .A(y[7936]), .B(x[511]), .Z(n27825) );
  NAND U29217 ( .A(y[7963]), .B(x[484]), .Z(n27824) );
  XNOR U29218 ( .A(n27825), .B(n27824), .Z(n27826) );
  XNOR U29219 ( .A(n27827), .B(n27826), .Z(n27828) );
  XNOR U29220 ( .A(n27829), .B(n27828), .Z(n27830) );
  XNOR U29221 ( .A(n27831), .B(n27830), .Z(n27832) );
  XNOR U29222 ( .A(n27833), .B(n27832), .Z(n27849) );
  AND U29223 ( .A(n27835), .B(n27834), .Z(n27839) );
  AND U29224 ( .A(n27837), .B(n27836), .Z(n27838) );
  NOR U29225 ( .A(n27839), .B(n27838), .Z(n27847) );
  NAND U29226 ( .A(n27841), .B(n27840), .Z(n27845) );
  NAND U29227 ( .A(n27843), .B(n27842), .Z(n27844) );
  AND U29228 ( .A(n27845), .B(n27844), .Z(n27846) );
  XNOR U29229 ( .A(n27847), .B(n27846), .Z(n27848) );
  XNOR U29230 ( .A(n27849), .B(n27848), .Z(n27850) );
  XNOR U29231 ( .A(n27851), .B(n27850), .Z(n27933) );
  AND U29232 ( .A(n27853), .B(n27852), .Z(n27857) );
  AND U29233 ( .A(n27855), .B(n27854), .Z(n27856) );
  NOR U29234 ( .A(n27857), .B(n27856), .Z(n27931) );
  NAND U29235 ( .A(n27859), .B(n27858), .Z(n27863) );
  NAND U29236 ( .A(n27861), .B(n27860), .Z(n27862) );
  AND U29237 ( .A(n27863), .B(n27862), .Z(n27870) );
  NAND U29238 ( .A(n27864), .B(n27901), .Z(n27868) );
  NAND U29239 ( .A(n27866), .B(n27865), .Z(n27867) );
  AND U29240 ( .A(n27868), .B(n27867), .Z(n27869) );
  XNOR U29241 ( .A(n27870), .B(n27869), .Z(n27929) );
  NAND U29242 ( .A(n27872), .B(n27871), .Z(n27875) );
  AND U29243 ( .A(x[490]), .B(y[7957]), .Z(n27900) );
  NANDN U29244 ( .A(n27873), .B(n27900), .Z(n27874) );
  AND U29245 ( .A(n27875), .B(n27874), .Z(n27927) );
  AND U29246 ( .A(y[7962]), .B(x[485]), .Z(n27885) );
  AND U29247 ( .A(n27876), .B(o[286]), .Z(n27883) );
  XOR U29248 ( .A(n27877), .B(o[287]), .Z(n27881) );
  XNOR U29249 ( .A(n27879), .B(n27878), .Z(n27880) );
  XNOR U29250 ( .A(n27881), .B(n27880), .Z(n27882) );
  XNOR U29251 ( .A(n27883), .B(n27882), .Z(n27884) );
  XNOR U29252 ( .A(n27885), .B(n27884), .Z(n27925) );
  AND U29253 ( .A(y[7950]), .B(x[497]), .Z(n27891) );
  AND U29254 ( .A(y[7966]), .B(x[481]), .Z(n27887) );
  NAND U29255 ( .A(y[7939]), .B(x[508]), .Z(n27886) );
  XNOR U29256 ( .A(n27887), .B(n27886), .Z(n27888) );
  XNOR U29257 ( .A(n27889), .B(n27888), .Z(n27890) );
  XNOR U29258 ( .A(n27891), .B(n27890), .Z(n27915) );
  AND U29259 ( .A(y[7946]), .B(x[501]), .Z(n27893) );
  NAND U29260 ( .A(y[7959]), .B(x[488]), .Z(n27892) );
  XNOR U29261 ( .A(n27893), .B(n27892), .Z(n27905) );
  AND U29262 ( .A(y[7948]), .B(x[499]), .Z(n27895) );
  NAND U29263 ( .A(y[7944]), .B(x[503]), .Z(n27894) );
  XNOR U29264 ( .A(n27895), .B(n27894), .Z(n27899) );
  AND U29265 ( .A(y[7940]), .B(x[507]), .Z(n27897) );
  NAND U29266 ( .A(y[7965]), .B(x[482]), .Z(n27896) );
  XNOR U29267 ( .A(n27897), .B(n27896), .Z(n27898) );
  XOR U29268 ( .A(n27899), .B(n27898), .Z(n27903) );
  XNOR U29269 ( .A(n27901), .B(n27900), .Z(n27902) );
  XNOR U29270 ( .A(n27903), .B(n27902), .Z(n27904) );
  XOR U29271 ( .A(n27905), .B(n27904), .Z(n27913) );
  AND U29272 ( .A(y[7961]), .B(x[486]), .Z(n27907) );
  NAND U29273 ( .A(y[7960]), .B(x[487]), .Z(n27906) );
  XNOR U29274 ( .A(n27907), .B(n27906), .Z(n27911) );
  AND U29275 ( .A(y[7964]), .B(x[483]), .Z(n27909) );
  NAND U29276 ( .A(y[7949]), .B(x[498]), .Z(n27908) );
  XNOR U29277 ( .A(n27909), .B(n27908), .Z(n27910) );
  XNOR U29278 ( .A(n27911), .B(n27910), .Z(n27912) );
  XNOR U29279 ( .A(n27913), .B(n27912), .Z(n27914) );
  XOR U29280 ( .A(n27915), .B(n27914), .Z(n27923) );
  AND U29281 ( .A(y[7951]), .B(x[496]), .Z(n27917) );
  NAND U29282 ( .A(y[7947]), .B(x[500]), .Z(n27916) );
  XNOR U29283 ( .A(n27917), .B(n27916), .Z(n27921) );
  AND U29284 ( .A(y[7937]), .B(x[510]), .Z(n27919) );
  NAND U29285 ( .A(y[7938]), .B(x[509]), .Z(n27918) );
  XNOR U29286 ( .A(n27919), .B(n27918), .Z(n27920) );
  XNOR U29287 ( .A(n27921), .B(n27920), .Z(n27922) );
  XNOR U29288 ( .A(n27923), .B(n27922), .Z(n27924) );
  XNOR U29289 ( .A(n27925), .B(n27924), .Z(n27926) );
  XNOR U29290 ( .A(n27927), .B(n27926), .Z(n27928) );
  XOR U29291 ( .A(n27929), .B(n27928), .Z(n27930) );
  XNOR U29292 ( .A(n27931), .B(n27930), .Z(n27932) );
  XNOR U29293 ( .A(n27933), .B(n27932), .Z(n27934) );
  XNOR U29294 ( .A(n27935), .B(n27934), .Z(n27951) );
  NAND U29295 ( .A(n27937), .B(n27936), .Z(n27941) );
  NAND U29296 ( .A(n27939), .B(n27938), .Z(n27940) );
  AND U29297 ( .A(n27941), .B(n27940), .Z(n27949) );
  NAND U29298 ( .A(n27943), .B(n27942), .Z(n27947) );
  NAND U29299 ( .A(n27945), .B(n27944), .Z(n27946) );
  NAND U29300 ( .A(n27947), .B(n27946), .Z(n27948) );
  XNOR U29301 ( .A(n27949), .B(n27948), .Z(n27950) );
  XNOR U29302 ( .A(n27951), .B(n27950), .Z(n27952) );
  XNOR U29303 ( .A(n27953), .B(n27952), .Z(n27954) );
  XNOR U29304 ( .A(n27955), .B(n27954), .Z(n27956) );
  XNOR U29305 ( .A(n27957), .B(n27956), .Z(n27973) );
  NAND U29306 ( .A(n27959), .B(n27958), .Z(n27963) );
  NAND U29307 ( .A(n27961), .B(n27960), .Z(n27962) );
  AND U29308 ( .A(n27963), .B(n27962), .Z(n27971) );
  NANDN U29309 ( .A(n27965), .B(n27964), .Z(n27969) );
  NAND U29310 ( .A(n27967), .B(n27966), .Z(n27968) );
  NAND U29311 ( .A(n27969), .B(n27968), .Z(n27970) );
  XNOR U29312 ( .A(n27971), .B(n27970), .Z(n27972) );
  XNOR U29313 ( .A(n27973), .B(n27972), .Z(n27974) );
  XNOR U29314 ( .A(n27975), .B(n27974), .Z(n27991) );
  NANDN U29315 ( .A(n27977), .B(n27976), .Z(n27981) );
  NANDN U29316 ( .A(n27979), .B(n27978), .Z(n27980) );
  AND U29317 ( .A(n27981), .B(n27980), .Z(n27989) );
  NAND U29318 ( .A(n27983), .B(n27982), .Z(n27987) );
  NANDN U29319 ( .A(n27985), .B(n27984), .Z(n27986) );
  NAND U29320 ( .A(n27987), .B(n27986), .Z(n27988) );
  XNOR U29321 ( .A(n27989), .B(n27988), .Z(n27990) );
  XNOR U29322 ( .A(n27991), .B(n27990), .Z(n27992) );
  XNOR U29323 ( .A(n27993), .B(n27992), .Z(n28017) );
  NAND U29324 ( .A(n27995), .B(n27994), .Z(n27999) );
  NAND U29325 ( .A(n27997), .B(n27996), .Z(n27998) );
  AND U29326 ( .A(n27999), .B(n27998), .Z(n28007) );
  NANDN U29327 ( .A(n28001), .B(n28000), .Z(n28005) );
  NANDN U29328 ( .A(n28003), .B(n28002), .Z(n28004) );
  NAND U29329 ( .A(n28005), .B(n28004), .Z(n28006) );
  XNOR U29330 ( .A(n28007), .B(n28006), .Z(n28015) );
  OR U29331 ( .A(n28008), .B(n28009), .Z(n28013) );
  AND U29332 ( .A(n28009), .B(n28008), .Z(n28010) );
  OR U29333 ( .A(n28011), .B(n28010), .Z(n28012) );
  NAND U29334 ( .A(n28013), .B(n28012), .Z(n28014) );
  XNOR U29335 ( .A(n28015), .B(n28014), .Z(n28016) );
  XNOR U29336 ( .A(n28017), .B(n28016), .Z(n28018) );
  XNOR U29337 ( .A(n28019), .B(n28018), .Z(n28035) );
  ANDN U29338 ( .B(n28021), .A(n28020), .Z(n28025) );
  ANDN U29339 ( .B(n28023), .A(n28022), .Z(n28024) );
  NOR U29340 ( .A(n28025), .B(n28024), .Z(n28033) );
  NAND U29341 ( .A(n28027), .B(n28026), .Z(n28031) );
  NAND U29342 ( .A(n28029), .B(n28028), .Z(n28030) );
  AND U29343 ( .A(n28031), .B(n28030), .Z(n28032) );
  XNOR U29344 ( .A(n28033), .B(n28032), .Z(n28034) );
  XNOR U29345 ( .A(n28035), .B(n28034), .Z(N576) );
  AND U29346 ( .A(x[480]), .B(y[7968]), .Z(n28679) );
  XOR U29347 ( .A(n28679), .B(o[288]), .Z(N609) );
  AND U29348 ( .A(x[481]), .B(y[7968]), .Z(n28044) );
  AND U29349 ( .A(x[480]), .B(y[7969]), .Z(n28043) );
  XNOR U29350 ( .A(n28043), .B(o[289]), .Z(n28036) );
  XNOR U29351 ( .A(n28044), .B(n28036), .Z(n28038) );
  NAND U29352 ( .A(n28679), .B(o[288]), .Z(n28037) );
  XNOR U29353 ( .A(n28038), .B(n28037), .Z(N610) );
  NANDN U29354 ( .A(n28044), .B(n28036), .Z(n28040) );
  NAND U29355 ( .A(n28038), .B(n28037), .Z(n28039) );
  AND U29356 ( .A(n28040), .B(n28039), .Z(n28050) );
  AND U29357 ( .A(x[480]), .B(y[7970]), .Z(n28058) );
  XNOR U29358 ( .A(n28058), .B(o[290]), .Z(n28049) );
  XNOR U29359 ( .A(n28050), .B(n28049), .Z(n28052) );
  AND U29360 ( .A(y[7968]), .B(x[482]), .Z(n28042) );
  NAND U29361 ( .A(y[7969]), .B(x[481]), .Z(n28041) );
  XNOR U29362 ( .A(n28042), .B(n28041), .Z(n28046) );
  AND U29363 ( .A(n28043), .B(o[289]), .Z(n28045) );
  XNOR U29364 ( .A(n28046), .B(n28045), .Z(n28051) );
  XNOR U29365 ( .A(n28052), .B(n28051), .Z(N611) );
  AND U29366 ( .A(x[482]), .B(y[7969]), .Z(n28055) );
  IV U29367 ( .A(n28055), .Z(n28063) );
  NANDN U29368 ( .A(n28063), .B(n28044), .Z(n28048) );
  NAND U29369 ( .A(n28046), .B(n28045), .Z(n28047) );
  AND U29370 ( .A(n28048), .B(n28047), .Z(n28071) );
  NANDN U29371 ( .A(n28050), .B(n28049), .Z(n28054) );
  NAND U29372 ( .A(n28052), .B(n28051), .Z(n28053) );
  AND U29373 ( .A(n28054), .B(n28053), .Z(n28070) );
  XNOR U29374 ( .A(n28071), .B(n28070), .Z(n28073) );
  AND U29375 ( .A(x[481]), .B(y[7970]), .Z(n28161) );
  XOR U29376 ( .A(o[291]), .B(n28055), .Z(n28067) );
  XOR U29377 ( .A(n28161), .B(n28067), .Z(n28069) );
  AND U29378 ( .A(y[7968]), .B(x[483]), .Z(n28057) );
  NAND U29379 ( .A(y[7971]), .B(x[480]), .Z(n28056) );
  XNOR U29380 ( .A(n28057), .B(n28056), .Z(n28060) );
  AND U29381 ( .A(n28058), .B(o[290]), .Z(n28059) );
  XOR U29382 ( .A(n28060), .B(n28059), .Z(n28068) );
  XOR U29383 ( .A(n28069), .B(n28068), .Z(n28072) );
  XOR U29384 ( .A(n28073), .B(n28072), .Z(N612) );
  AND U29385 ( .A(x[483]), .B(y[7971]), .Z(n28118) );
  NAND U29386 ( .A(n28679), .B(n28118), .Z(n28062) );
  NAND U29387 ( .A(n28060), .B(n28059), .Z(n28061) );
  NAND U29388 ( .A(n28062), .B(n28061), .Z(n28092) );
  ANDN U29389 ( .B(o[291]), .A(n28063), .Z(n28086) );
  AND U29390 ( .A(x[480]), .B(y[7972]), .Z(n28065) );
  AND U29391 ( .A(y[7968]), .B(x[484]), .Z(n28064) );
  XOR U29392 ( .A(n28065), .B(n28064), .Z(n28085) );
  XOR U29393 ( .A(n28086), .B(n28085), .Z(n28091) );
  AND U29394 ( .A(x[482]), .B(y[7970]), .Z(n28196) );
  NAND U29395 ( .A(y[7971]), .B(x[481]), .Z(n28066) );
  XNOR U29396 ( .A(n28196), .B(n28066), .Z(n28084) );
  AND U29397 ( .A(x[483]), .B(y[7969]), .Z(n28079) );
  XOR U29398 ( .A(n28079), .B(o[292]), .Z(n28083) );
  XOR U29399 ( .A(n28084), .B(n28083), .Z(n28090) );
  XOR U29400 ( .A(n28091), .B(n28090), .Z(n28093) );
  XNOR U29401 ( .A(n28092), .B(n28093), .Z(n28089) );
  NANDN U29402 ( .A(n28071), .B(n28070), .Z(n28075) );
  NAND U29403 ( .A(n28073), .B(n28072), .Z(n28074) );
  NAND U29404 ( .A(n28075), .B(n28074), .Z(n28088) );
  XOR U29405 ( .A(n28087), .B(n28088), .Z(n28076) );
  XNOR U29406 ( .A(n28089), .B(n28076), .Z(N613) );
  AND U29407 ( .A(y[7968]), .B(x[485]), .Z(n28078) );
  NAND U29408 ( .A(y[7973]), .B(x[480]), .Z(n28077) );
  XNOR U29409 ( .A(n28078), .B(n28077), .Z(n28110) );
  AND U29410 ( .A(n28079), .B(o[292]), .Z(n28111) );
  XOR U29411 ( .A(n28110), .B(n28111), .Z(n28109) );
  NAND U29412 ( .A(x[482]), .B(y[7971]), .Z(n28169) );
  AND U29413 ( .A(y[7970]), .B(x[483]), .Z(n28081) );
  NAND U29414 ( .A(y[7972]), .B(x[481]), .Z(n28080) );
  XNOR U29415 ( .A(n28081), .B(n28080), .Z(n28105) );
  AND U29416 ( .A(x[484]), .B(y[7969]), .Z(n28116) );
  XOR U29417 ( .A(n28116), .B(o[293]), .Z(n28104) );
  XOR U29418 ( .A(n28105), .B(n28104), .Z(n28108) );
  XOR U29419 ( .A(n28169), .B(n28108), .Z(n28082) );
  XNOR U29420 ( .A(n28109), .B(n28082), .Z(n28100) );
  AND U29421 ( .A(x[484]), .B(y[7972]), .Z(n28883) );
  XOR U29422 ( .A(n28097), .B(n28098), .Z(n28099) );
  XNOR U29423 ( .A(n28100), .B(n28099), .Z(n28103) );
  NAND U29424 ( .A(n28091), .B(n28090), .Z(n28095) );
  NAND U29425 ( .A(n28093), .B(n28092), .Z(n28094) );
  NAND U29426 ( .A(n28095), .B(n28094), .Z(n28101) );
  XNOR U29427 ( .A(n28102), .B(n28101), .Z(n28096) );
  XNOR U29428 ( .A(n28103), .B(n28096), .Z(N614) );
  AND U29429 ( .A(x[483]), .B(y[7972]), .Z(n28170) );
  NAND U29430 ( .A(n28170), .B(n28161), .Z(n28107) );
  NAND U29431 ( .A(n28105), .B(n28104), .Z(n28106) );
  NAND U29432 ( .A(n28107), .B(n28106), .Z(n28146) );
  XOR U29433 ( .A(n28146), .B(n28145), .Z(n28148) );
  AND U29434 ( .A(x[485]), .B(y[7973]), .Z(n28339) );
  NAND U29435 ( .A(n28679), .B(n28339), .Z(n28113) );
  NAND U29436 ( .A(n28111), .B(n28110), .Z(n28112) );
  NAND U29437 ( .A(n28113), .B(n28112), .Z(n28122) );
  AND U29438 ( .A(y[7968]), .B(x[486]), .Z(n28115) );
  NAND U29439 ( .A(y[7974]), .B(x[480]), .Z(n28114) );
  XNOR U29440 ( .A(n28115), .B(n28114), .Z(n28128) );
  AND U29441 ( .A(n28116), .B(o[293]), .Z(n28129) );
  XOR U29442 ( .A(n28128), .B(n28129), .Z(n28121) );
  XOR U29443 ( .A(n28122), .B(n28121), .Z(n28124) );
  NAND U29444 ( .A(y[7972]), .B(x[482]), .Z(n28117) );
  XNOR U29445 ( .A(n28118), .B(n28117), .Z(n28133) );
  AND U29446 ( .A(y[7973]), .B(x[481]), .Z(n28372) );
  NAND U29447 ( .A(y[7970]), .B(x[484]), .Z(n28119) );
  XNOR U29448 ( .A(n28372), .B(n28119), .Z(n28137) );
  AND U29449 ( .A(x[485]), .B(y[7969]), .Z(n28144) );
  XOR U29450 ( .A(o[294]), .B(n28144), .Z(n28136) );
  XOR U29451 ( .A(n28137), .B(n28136), .Z(n28132) );
  XOR U29452 ( .A(n28133), .B(n28132), .Z(n28123) );
  XOR U29453 ( .A(n28124), .B(n28123), .Z(n28147) );
  XOR U29454 ( .A(n28148), .B(n28147), .Z(n28153) );
  XOR U29455 ( .A(n28151), .B(n28153), .Z(n28120) );
  XOR U29456 ( .A(n28152), .B(n28120), .Z(N615) );
  NAND U29457 ( .A(n28122), .B(n28121), .Z(n28126) );
  NAND U29458 ( .A(n28124), .B(n28123), .Z(n28125) );
  AND U29459 ( .A(n28126), .B(n28125), .Z(n28192) );
  AND U29460 ( .A(y[7970]), .B(x[485]), .Z(n28261) );
  NAND U29461 ( .A(y[7974]), .B(x[481]), .Z(n28127) );
  XNOR U29462 ( .A(n28261), .B(n28127), .Z(n28163) );
  AND U29463 ( .A(x[486]), .B(y[7969]), .Z(n28166) );
  XOR U29464 ( .A(o[295]), .B(n28166), .Z(n28162) );
  XNOR U29465 ( .A(n28163), .B(n28162), .Z(n28181) );
  AND U29466 ( .A(x[486]), .B(y[7974]), .Z(n28392) );
  NAND U29467 ( .A(n28679), .B(n28392), .Z(n28131) );
  NAND U29468 ( .A(n28129), .B(n28128), .Z(n28130) );
  AND U29469 ( .A(n28131), .B(n28130), .Z(n28180) );
  XOR U29470 ( .A(n28181), .B(n28180), .Z(n28182) );
  NANDN U29471 ( .A(n28169), .B(n28170), .Z(n28135) );
  NAND U29472 ( .A(n28133), .B(n28132), .Z(n28134) );
  AND U29473 ( .A(n28135), .B(n28134), .Z(n28183) );
  XOR U29474 ( .A(n28182), .B(n28183), .Z(n28190) );
  AND U29475 ( .A(x[484]), .B(y[7973]), .Z(n28684) );
  NAND U29476 ( .A(n28684), .B(n28161), .Z(n28139) );
  NAND U29477 ( .A(n28137), .B(n28136), .Z(n28138) );
  AND U29478 ( .A(n28139), .B(n28138), .Z(n28158) );
  AND U29479 ( .A(y[7973]), .B(x[482]), .Z(n28141) );
  NAND U29480 ( .A(y[7971]), .B(x[484]), .Z(n28140) );
  XNOR U29481 ( .A(n28141), .B(n28140), .Z(n28171) );
  XNOR U29482 ( .A(n28171), .B(n28170), .Z(n28156) );
  AND U29483 ( .A(y[7968]), .B(x[487]), .Z(n28143) );
  NAND U29484 ( .A(y[7975]), .B(x[480]), .Z(n28142) );
  XNOR U29485 ( .A(n28143), .B(n28142), .Z(n28175) );
  AND U29486 ( .A(o[294]), .B(n28144), .Z(n28174) );
  XNOR U29487 ( .A(n28175), .B(n28174), .Z(n28155) );
  XOR U29488 ( .A(n28156), .B(n28155), .Z(n28157) );
  XOR U29489 ( .A(n28158), .B(n28157), .Z(n28189) );
  XOR U29490 ( .A(n28190), .B(n28189), .Z(n28191) );
  XOR U29491 ( .A(n28192), .B(n28191), .Z(n28188) );
  NAND U29492 ( .A(n28146), .B(n28145), .Z(n28150) );
  NAND U29493 ( .A(n28148), .B(n28147), .Z(n28149) );
  NAND U29494 ( .A(n28150), .B(n28149), .Z(n28187) );
  XOR U29495 ( .A(n28187), .B(n28186), .Z(n28154) );
  XNOR U29496 ( .A(n28188), .B(n28154), .Z(N616) );
  NAND U29497 ( .A(n28156), .B(n28155), .Z(n28160) );
  NAND U29498 ( .A(n28158), .B(n28157), .Z(n28159) );
  AND U29499 ( .A(n28160), .B(n28159), .Z(n28229) );
  AND U29500 ( .A(x[485]), .B(y[7974]), .Z(n28330) );
  NAND U29501 ( .A(n28330), .B(n28161), .Z(n28165) );
  NAND U29502 ( .A(n28163), .B(n28162), .Z(n28164) );
  AND U29503 ( .A(n28165), .B(n28164), .Z(n28227) );
  AND U29504 ( .A(o[295]), .B(n28166), .Z(n28216) );
  AND U29505 ( .A(y[7971]), .B(x[485]), .Z(n28788) );
  NAND U29506 ( .A(y[7975]), .B(x[481]), .Z(n28167) );
  XNOR U29507 ( .A(n28788), .B(n28167), .Z(n28217) );
  XNOR U29508 ( .A(n28216), .B(n28217), .Z(n28201) );
  NAND U29509 ( .A(x[483]), .B(y[7973]), .Z(n29019) );
  AND U29510 ( .A(x[486]), .B(y[7970]), .Z(n28168) );
  AND U29511 ( .A(y[7974]), .B(x[482]), .Z(n29113) );
  XOR U29512 ( .A(n28168), .B(n29113), .Z(n28197) );
  XOR U29513 ( .A(n28883), .B(n28197), .Z(n28200) );
  XOR U29514 ( .A(n28201), .B(n28202), .Z(n28226) );
  XOR U29515 ( .A(n28229), .B(n28228), .Z(n28242) );
  NANDN U29516 ( .A(n28169), .B(n28684), .Z(n28173) );
  NAND U29517 ( .A(n28171), .B(n28170), .Z(n28172) );
  AND U29518 ( .A(n28173), .B(n28172), .Z(n28223) );
  AND U29519 ( .A(x[487]), .B(y[7975]), .Z(n28568) );
  NAND U29520 ( .A(n28679), .B(n28568), .Z(n28177) );
  NAND U29521 ( .A(n28175), .B(n28174), .Z(n28176) );
  AND U29522 ( .A(n28177), .B(n28176), .Z(n28221) );
  AND U29523 ( .A(y[7968]), .B(x[488]), .Z(n28179) );
  NAND U29524 ( .A(y[7976]), .B(x[480]), .Z(n28178) );
  XNOR U29525 ( .A(n28179), .B(n28178), .Z(n28207) );
  AND U29526 ( .A(x[487]), .B(y[7969]), .Z(n28210) );
  XOR U29527 ( .A(o[296]), .B(n28210), .Z(n28206) );
  XOR U29528 ( .A(n28207), .B(n28206), .Z(n28220) );
  NAND U29529 ( .A(n28181), .B(n28180), .Z(n28185) );
  NAND U29530 ( .A(n28183), .B(n28182), .Z(n28184) );
  NAND U29531 ( .A(n28185), .B(n28184), .Z(n28239) );
  XOR U29532 ( .A(n28240), .B(n28239), .Z(n28241) );
  XOR U29533 ( .A(n28242), .B(n28241), .Z(n28235) );
  NAND U29534 ( .A(n28190), .B(n28189), .Z(n28194) );
  NAND U29535 ( .A(n28192), .B(n28191), .Z(n28193) );
  NAND U29536 ( .A(n28194), .B(n28193), .Z(n28234) );
  IV U29537 ( .A(n28234), .Z(n28232) );
  XOR U29538 ( .A(n28233), .B(n28232), .Z(n28195) );
  XNOR U29539 ( .A(n28235), .B(n28195), .Z(N617) );
  NAND U29540 ( .A(n28392), .B(n28196), .Z(n28199) );
  NAND U29541 ( .A(n28883), .B(n28197), .Z(n28198) );
  NAND U29542 ( .A(n28199), .B(n28198), .Z(n28255) );
  NANDN U29543 ( .A(n28200), .B(n29019), .Z(n28204) );
  NANDN U29544 ( .A(n28202), .B(n28201), .Z(n28203) );
  AND U29545 ( .A(n28204), .B(n28203), .Z(n28256) );
  XOR U29546 ( .A(n28255), .B(n28256), .Z(n28257) );
  AND U29547 ( .A(x[488]), .B(y[7976]), .Z(n28205) );
  NAND U29548 ( .A(n28205), .B(n28679), .Z(n28209) );
  NAND U29549 ( .A(n28207), .B(n28206), .Z(n28208) );
  AND U29550 ( .A(n28209), .B(n28208), .Z(n28290) );
  AND U29551 ( .A(o[296]), .B(n28210), .Z(n28263) );
  AND U29552 ( .A(y[7972]), .B(x[485]), .Z(n28212) );
  NAND U29553 ( .A(y[7970]), .B(x[487]), .Z(n28211) );
  XNOR U29554 ( .A(n28212), .B(n28211), .Z(n28262) );
  XNOR U29555 ( .A(n28263), .B(n28262), .Z(n28288) );
  AND U29556 ( .A(y[7968]), .B(x[489]), .Z(n28214) );
  NAND U29557 ( .A(y[7977]), .B(x[480]), .Z(n28213) );
  XNOR U29558 ( .A(n28214), .B(n28213), .Z(n28270) );
  AND U29559 ( .A(x[488]), .B(y[7969]), .Z(n28277) );
  XOR U29560 ( .A(o[297]), .B(n28277), .Z(n28269) );
  XNOR U29561 ( .A(n28270), .B(n28269), .Z(n28287) );
  XOR U29562 ( .A(n28288), .B(n28287), .Z(n28289) );
  XNOR U29563 ( .A(n28290), .B(n28289), .Z(n28284) );
  AND U29564 ( .A(y[7971]), .B(x[486]), .Z(n28623) );
  NAND U29565 ( .A(y[7976]), .B(x[481]), .Z(n28215) );
  XNOR U29566 ( .A(n28623), .B(n28215), .Z(n28274) );
  XNOR U29567 ( .A(n28684), .B(n28274), .Z(n28294) );
  AND U29568 ( .A(x[482]), .B(y[7975]), .Z(n28926) );
  NAND U29569 ( .A(x[483]), .B(y[7974]), .Z(n28633) );
  XNOR U29570 ( .A(n28926), .B(n28633), .Z(n28293) );
  XNOR U29571 ( .A(n28294), .B(n28293), .Z(n28282) );
  NAND U29572 ( .A(x[485]), .B(y[7975]), .Z(n28472) );
  AND U29573 ( .A(x[481]), .B(y[7971]), .Z(n28273) );
  NANDN U29574 ( .A(n28472), .B(n28273), .Z(n28219) );
  NAND U29575 ( .A(n28217), .B(n28216), .Z(n28218) );
  NAND U29576 ( .A(n28219), .B(n28218), .Z(n28281) );
  XOR U29577 ( .A(n28282), .B(n28281), .Z(n28283) );
  XNOR U29578 ( .A(n28284), .B(n28283), .Z(n28258) );
  XNOR U29579 ( .A(n28257), .B(n28258), .Z(n28249) );
  NANDN U29580 ( .A(n28221), .B(n28220), .Z(n28225) );
  NANDN U29581 ( .A(n28223), .B(n28222), .Z(n28224) );
  AND U29582 ( .A(n28225), .B(n28224), .Z(n28247) );
  NANDN U29583 ( .A(n28227), .B(n28226), .Z(n28231) );
  NAND U29584 ( .A(n28229), .B(n28228), .Z(n28230) );
  NAND U29585 ( .A(n28231), .B(n28230), .Z(n28246) );
  XNOR U29586 ( .A(n28249), .B(n28248), .Z(n28254) );
  NANDN U29587 ( .A(n28232), .B(n28233), .Z(n28238) );
  NOR U29588 ( .A(n28234), .B(n28233), .Z(n28236) );
  OR U29589 ( .A(n28236), .B(n28235), .Z(n28237) );
  AND U29590 ( .A(n28238), .B(n28237), .Z(n28252) );
  NAND U29591 ( .A(n28240), .B(n28239), .Z(n28244) );
  NANDN U29592 ( .A(n28242), .B(n28241), .Z(n28243) );
  AND U29593 ( .A(n28244), .B(n28243), .Z(n28253) );
  XOR U29594 ( .A(n28252), .B(n28253), .Z(n28245) );
  XNOR U29595 ( .A(n28254), .B(n28245), .Z(N618) );
  NANDN U29596 ( .A(n28247), .B(n28246), .Z(n28251) );
  NAND U29597 ( .A(n28249), .B(n28248), .Z(n28250) );
  NAND U29598 ( .A(n28251), .B(n28250), .Z(n28349) );
  IV U29599 ( .A(n28349), .Z(n28348) );
  NAND U29600 ( .A(n28256), .B(n28255), .Z(n28260) );
  NANDN U29601 ( .A(n28258), .B(n28257), .Z(n28259) );
  AND U29602 ( .A(n28260), .B(n28259), .Z(n28357) );
  AND U29603 ( .A(x[487]), .B(y[7972]), .Z(n28332) );
  NAND U29604 ( .A(n28332), .B(n28261), .Z(n28265) );
  NAND U29605 ( .A(n28263), .B(n28262), .Z(n28264) );
  AND U29606 ( .A(n28265), .B(n28264), .Z(n28345) );
  AND U29607 ( .A(y[7971]), .B(x[487]), .Z(n28267) );
  NAND U29608 ( .A(y[7974]), .B(x[484]), .Z(n28266) );
  XNOR U29609 ( .A(n28267), .B(n28266), .Z(n28316) );
  AND U29610 ( .A(x[486]), .B(y[7972]), .Z(n28315) );
  XNOR U29611 ( .A(n28316), .B(n28315), .Z(n28343) );
  AND U29612 ( .A(x[488]), .B(y[7970]), .Z(n28532) );
  NAND U29613 ( .A(x[489]), .B(y[7969]), .Z(n28326) );
  XOR U29614 ( .A(n28532), .B(n28337), .Z(n28338) );
  XNOR U29615 ( .A(n28339), .B(n28338), .Z(n28342) );
  XOR U29616 ( .A(n28343), .B(n28342), .Z(n28344) );
  XNOR U29617 ( .A(n28345), .B(n28344), .Z(n28305) );
  AND U29618 ( .A(x[489]), .B(y[7977]), .Z(n28268) );
  NAND U29619 ( .A(n28268), .B(n28679), .Z(n28272) );
  NAND U29620 ( .A(n28270), .B(n28269), .Z(n28271) );
  NAND U29621 ( .A(n28272), .B(n28271), .Z(n28303) );
  AND U29622 ( .A(x[486]), .B(y[7976]), .Z(n28559) );
  NAND U29623 ( .A(n28559), .B(n28273), .Z(n28276) );
  NAND U29624 ( .A(n28684), .B(n28274), .Z(n28275) );
  NAND U29625 ( .A(n28276), .B(n28275), .Z(n28311) );
  AND U29626 ( .A(o[297]), .B(n28277), .Z(n28321) );
  AND U29627 ( .A(y[7968]), .B(x[490]), .Z(n28279) );
  AND U29628 ( .A(y[7978]), .B(x[480]), .Z(n28278) );
  XOR U29629 ( .A(n28279), .B(n28278), .Z(n28320) );
  XOR U29630 ( .A(n28321), .B(n28320), .Z(n28309) );
  AND U29631 ( .A(y[7975]), .B(x[483]), .Z(n29249) );
  NAND U29632 ( .A(y[7977]), .B(x[481]), .Z(n28280) );
  XNOR U29633 ( .A(n29249), .B(n28280), .Z(n28333) );
  AND U29634 ( .A(x[482]), .B(y[7976]), .Z(n28334) );
  XOR U29635 ( .A(n28333), .B(n28334), .Z(n28308) );
  XOR U29636 ( .A(n28309), .B(n28308), .Z(n28310) );
  XOR U29637 ( .A(n28311), .B(n28310), .Z(n28302) );
  XOR U29638 ( .A(n28303), .B(n28302), .Z(n28304) );
  XOR U29639 ( .A(n28305), .B(n28304), .Z(n28356) );
  NAND U29640 ( .A(n28282), .B(n28281), .Z(n28286) );
  NAND U29641 ( .A(n28284), .B(n28283), .Z(n28285) );
  NAND U29642 ( .A(n28286), .B(n28285), .Z(n28299) );
  NAND U29643 ( .A(n28288), .B(n28287), .Z(n28292) );
  NAND U29644 ( .A(n28290), .B(n28289), .Z(n28291) );
  AND U29645 ( .A(n28292), .B(n28291), .Z(n28296) );
  XOR U29646 ( .A(n28296), .B(n28297), .Z(n28298) );
  XNOR U29647 ( .A(n28299), .B(n28298), .Z(n28355) );
  XNOR U29648 ( .A(n28357), .B(n28358), .Z(n28351) );
  XNOR U29649 ( .A(n28350), .B(n28351), .Z(n28295) );
  XOR U29650 ( .A(n28348), .B(n28295), .Z(N619) );
  NAND U29651 ( .A(n28297), .B(n28296), .Z(n28301) );
  NAND U29652 ( .A(n28299), .B(n28298), .Z(n28300) );
  AND U29653 ( .A(n28301), .B(n28300), .Z(n28427) );
  NAND U29654 ( .A(n28303), .B(n28302), .Z(n28307) );
  NAND U29655 ( .A(n28305), .B(n28304), .Z(n28306) );
  NAND U29656 ( .A(n28307), .B(n28306), .Z(n28425) );
  NAND U29657 ( .A(n28309), .B(n28308), .Z(n28313) );
  NAND U29658 ( .A(n28311), .B(n28310), .Z(n28312) );
  NAND U29659 ( .A(n28313), .B(n28312), .Z(n28413) );
  AND U29660 ( .A(x[487]), .B(y[7974]), .Z(n28467) );
  AND U29661 ( .A(x[484]), .B(y[7971]), .Z(n28314) );
  NAND U29662 ( .A(n28467), .B(n28314), .Z(n28318) );
  NAND U29663 ( .A(n28316), .B(n28315), .Z(n28317) );
  NAND U29664 ( .A(n28318), .B(n28317), .Z(n28411) );
  AND U29665 ( .A(x[490]), .B(y[7978]), .Z(n28319) );
  NAND U29666 ( .A(n28319), .B(n28679), .Z(n28323) );
  NAND U29667 ( .A(n28321), .B(n28320), .Z(n28322) );
  NAND U29668 ( .A(n28323), .B(n28322), .Z(n28407) );
  AND U29669 ( .A(y[7968]), .B(x[491]), .Z(n28325) );
  NAND U29670 ( .A(y[7979]), .B(x[480]), .Z(n28324) );
  XNOR U29671 ( .A(n28325), .B(n28324), .Z(n28383) );
  ANDN U29672 ( .B(o[298]), .A(n28326), .Z(n28382) );
  XOR U29673 ( .A(n28383), .B(n28382), .Z(n28406) );
  AND U29674 ( .A(y[7973]), .B(x[486]), .Z(n28328) );
  NAND U29675 ( .A(y[7978]), .B(x[481]), .Z(n28327) );
  XNOR U29676 ( .A(n28328), .B(n28327), .Z(n28374) );
  AND U29677 ( .A(x[490]), .B(y[7969]), .Z(n28393) );
  XOR U29678 ( .A(o[299]), .B(n28393), .Z(n28373) );
  XOR U29679 ( .A(n28374), .B(n28373), .Z(n28405) );
  XOR U29680 ( .A(n28406), .B(n28405), .Z(n28408) );
  XNOR U29681 ( .A(n28407), .B(n28408), .Z(n28412) );
  XOR U29682 ( .A(n28413), .B(n28414), .Z(n28396) );
  AND U29683 ( .A(x[483]), .B(y[7976]), .Z(n29378) );
  NAND U29684 ( .A(y[7977]), .B(x[482]), .Z(n28329) );
  XNOR U29685 ( .A(n28330), .B(n28329), .Z(n28369) );
  AND U29686 ( .A(x[484]), .B(y[7975]), .Z(n28368) );
  XNOR U29687 ( .A(n28369), .B(n28368), .Z(n28400) );
  XNOR U29688 ( .A(n29378), .B(n28400), .Z(n28402) );
  NAND U29689 ( .A(y[7970]), .B(x[489]), .Z(n28331) );
  XNOR U29690 ( .A(n28332), .B(n28331), .Z(n28388) );
  AND U29691 ( .A(x[488]), .B(y[7971]), .Z(n28387) );
  XNOR U29692 ( .A(n28388), .B(n28387), .Z(n28401) );
  XNOR U29693 ( .A(n28402), .B(n28401), .Z(n28365) );
  AND U29694 ( .A(x[483]), .B(y[7977]), .Z(n28463) );
  AND U29695 ( .A(x[481]), .B(y[7975]), .Z(n28674) );
  NAND U29696 ( .A(n28463), .B(n28674), .Z(n28336) );
  NAND U29697 ( .A(n28334), .B(n28333), .Z(n28335) );
  NAND U29698 ( .A(n28336), .B(n28335), .Z(n28363) );
  NAND U29699 ( .A(n28532), .B(n28337), .Z(n28341) );
  NAND U29700 ( .A(n28339), .B(n28338), .Z(n28340) );
  NAND U29701 ( .A(n28341), .B(n28340), .Z(n28362) );
  XOR U29702 ( .A(n28363), .B(n28362), .Z(n28364) );
  XNOR U29703 ( .A(n28365), .B(n28364), .Z(n28395) );
  NAND U29704 ( .A(n28343), .B(n28342), .Z(n28347) );
  NAND U29705 ( .A(n28345), .B(n28344), .Z(n28346) );
  NAND U29706 ( .A(n28347), .B(n28346), .Z(n28394) );
  XOR U29707 ( .A(n28395), .B(n28394), .Z(n28397) );
  XNOR U29708 ( .A(n28396), .B(n28397), .Z(n28424) );
  XOR U29709 ( .A(n28425), .B(n28424), .Z(n28426) );
  XOR U29710 ( .A(n28427), .B(n28426), .Z(n28420) );
  OR U29711 ( .A(n28350), .B(n28348), .Z(n28354) );
  ANDN U29712 ( .B(n28350), .A(n28349), .Z(n28352) );
  OR U29713 ( .A(n28352), .B(n28351), .Z(n28353) );
  AND U29714 ( .A(n28354), .B(n28353), .Z(n28419) );
  NANDN U29715 ( .A(n28356), .B(n28355), .Z(n28360) );
  NANDN U29716 ( .A(n28358), .B(n28357), .Z(n28359) );
  AND U29717 ( .A(n28360), .B(n28359), .Z(n28418) );
  IV U29718 ( .A(n28418), .Z(n28417) );
  XOR U29719 ( .A(n28419), .B(n28417), .Z(n28361) );
  XNOR U29720 ( .A(n28420), .B(n28361), .Z(N620) );
  NAND U29721 ( .A(n28363), .B(n28362), .Z(n28367) );
  NAND U29722 ( .A(n28365), .B(n28364), .Z(n28366) );
  NAND U29723 ( .A(n28367), .B(n28366), .Z(n28503) );
  AND U29724 ( .A(x[485]), .B(y[7977]), .Z(n28919) );
  NAND U29725 ( .A(n29113), .B(n28919), .Z(n28371) );
  NAND U29726 ( .A(n28369), .B(n28368), .Z(n28370) );
  AND U29727 ( .A(n28371), .B(n28370), .Z(n28451) );
  AND U29728 ( .A(x[486]), .B(y[7978]), .Z(n28691) );
  NAND U29729 ( .A(n28691), .B(n28372), .Z(n28376) );
  NAND U29730 ( .A(n28374), .B(n28373), .Z(n28375) );
  NAND U29731 ( .A(n28376), .B(n28375), .Z(n28450) );
  AND U29732 ( .A(x[489]), .B(y[7971]), .Z(n29108) );
  AND U29733 ( .A(y[7970]), .B(x[490]), .Z(n29150) );
  NAND U29734 ( .A(y[7976]), .B(x[484]), .Z(n28377) );
  XOR U29735 ( .A(n29150), .B(n28377), .Z(n28494) );
  NAND U29736 ( .A(x[487]), .B(y[7973]), .Z(n28471) );
  XOR U29737 ( .A(n28472), .B(n28471), .Z(n28474) );
  AND U29738 ( .A(y[7968]), .B(x[492]), .Z(n28379) );
  NAND U29739 ( .A(y[7980]), .B(x[480]), .Z(n28378) );
  XNOR U29740 ( .A(n28379), .B(n28378), .Z(n28488) );
  AND U29741 ( .A(x[491]), .B(y[7969]), .Z(n28468) );
  XOR U29742 ( .A(o[300]), .B(n28468), .Z(n28487) );
  XOR U29743 ( .A(n28488), .B(n28487), .Z(n28457) );
  AND U29744 ( .A(y[7978]), .B(x[482]), .Z(n28381) );
  NAND U29745 ( .A(y[7972]), .B(x[488]), .Z(n28380) );
  XNOR U29746 ( .A(n28381), .B(n28380), .Z(n28462) );
  XOR U29747 ( .A(n28462), .B(n28463), .Z(n28456) );
  XOR U29748 ( .A(n28457), .B(n28456), .Z(n28459) );
  XOR U29749 ( .A(n28458), .B(n28459), .Z(n28452) );
  XOR U29750 ( .A(n28453), .B(n28452), .Z(n28502) );
  AND U29751 ( .A(x[491]), .B(y[7979]), .Z(n29501) );
  NAND U29752 ( .A(n29501), .B(n28679), .Z(n28385) );
  NAND U29753 ( .A(n28383), .B(n28382), .Z(n28384) );
  AND U29754 ( .A(n28385), .B(n28384), .Z(n28480) );
  AND U29755 ( .A(x[487]), .B(y[7970]), .Z(n28609) );
  AND U29756 ( .A(x[489]), .B(y[7972]), .Z(n28386) );
  NAND U29757 ( .A(n28609), .B(n28386), .Z(n28390) );
  NAND U29758 ( .A(n28388), .B(n28387), .Z(n28389) );
  AND U29759 ( .A(n28390), .B(n28389), .Z(n28478) );
  NAND U29760 ( .A(y[7979]), .B(x[481]), .Z(n28391) );
  XNOR U29761 ( .A(n28392), .B(n28391), .Z(n28484) );
  AND U29762 ( .A(o[299]), .B(n28393), .Z(n28483) );
  XOR U29763 ( .A(n28484), .B(n28483), .Z(n28477) );
  XOR U29764 ( .A(n28502), .B(n28501), .Z(n28504) );
  XNOR U29765 ( .A(n28503), .B(n28504), .Z(n28432) );
  NAND U29766 ( .A(n28395), .B(n28394), .Z(n28399) );
  NAND U29767 ( .A(n28397), .B(n28396), .Z(n28398) );
  NAND U29768 ( .A(n28399), .B(n28398), .Z(n28431) );
  XOR U29769 ( .A(n28432), .B(n28431), .Z(n28434) );
  NANDN U29770 ( .A(n29378), .B(n28400), .Z(n28404) );
  NAND U29771 ( .A(n28402), .B(n28401), .Z(n28403) );
  NAND U29772 ( .A(n28404), .B(n28403), .Z(n28444) );
  NAND U29773 ( .A(n28406), .B(n28405), .Z(n28410) );
  NAND U29774 ( .A(n28408), .B(n28407), .Z(n28409) );
  AND U29775 ( .A(n28410), .B(n28409), .Z(n28445) );
  XOR U29776 ( .A(n28444), .B(n28445), .Z(n28447) );
  NANDN U29777 ( .A(n28412), .B(n28411), .Z(n28416) );
  NANDN U29778 ( .A(n28414), .B(n28413), .Z(n28415) );
  AND U29779 ( .A(n28416), .B(n28415), .Z(n28446) );
  XOR U29780 ( .A(n28447), .B(n28446), .Z(n28433) );
  XNOR U29781 ( .A(n28434), .B(n28433), .Z(n28441) );
  OR U29782 ( .A(n28419), .B(n28417), .Z(n28423) );
  ANDN U29783 ( .B(n28419), .A(n28418), .Z(n28421) );
  OR U29784 ( .A(n28421), .B(n28420), .Z(n28422) );
  AND U29785 ( .A(n28423), .B(n28422), .Z(n28438) );
  NAND U29786 ( .A(n28425), .B(n28424), .Z(n28429) );
  NANDN U29787 ( .A(n28427), .B(n28426), .Z(n28428) );
  AND U29788 ( .A(n28429), .B(n28428), .Z(n28439) );
  IV U29789 ( .A(n28439), .Z(n28437) );
  XOR U29790 ( .A(n28438), .B(n28437), .Z(n28430) );
  XNOR U29791 ( .A(n28441), .B(n28430), .Z(N621) );
  NAND U29792 ( .A(n28432), .B(n28431), .Z(n28436) );
  NAND U29793 ( .A(n28434), .B(n28433), .Z(n28435) );
  AND U29794 ( .A(n28436), .B(n28435), .Z(n28576) );
  NANDN U29795 ( .A(n28437), .B(n28438), .Z(n28443) );
  NOR U29796 ( .A(n28439), .B(n28438), .Z(n28440) );
  OR U29797 ( .A(n28441), .B(n28440), .Z(n28442) );
  AND U29798 ( .A(n28443), .B(n28442), .Z(n28575) );
  NAND U29799 ( .A(n28445), .B(n28444), .Z(n28449) );
  NAND U29800 ( .A(n28447), .B(n28446), .Z(n28448) );
  NAND U29801 ( .A(n28449), .B(n28448), .Z(n28580) );
  NANDN U29802 ( .A(n28451), .B(n28450), .Z(n28455) );
  NAND U29803 ( .A(n28453), .B(n28452), .Z(n28454) );
  AND U29804 ( .A(n28455), .B(n28454), .Z(n28509) );
  NAND U29805 ( .A(n28457), .B(n28456), .Z(n28461) );
  NAND U29806 ( .A(n28459), .B(n28458), .Z(n28460) );
  NAND U29807 ( .A(n28461), .B(n28460), .Z(n28516) );
  AND U29808 ( .A(y[7978]), .B(x[488]), .Z(n29789) );
  AND U29809 ( .A(x[482]), .B(y[7972]), .Z(n28619) );
  NAND U29810 ( .A(n29789), .B(n28619), .Z(n28465) );
  NAND U29811 ( .A(n28463), .B(n28462), .Z(n28464) );
  NAND U29812 ( .A(n28465), .B(n28464), .Z(n28547) );
  NAND U29813 ( .A(y[7980]), .B(x[481]), .Z(n28466) );
  XNOR U29814 ( .A(n28467), .B(n28466), .Z(n28538) );
  AND U29815 ( .A(o[300]), .B(n28468), .Z(n28537) );
  XOR U29816 ( .A(n28538), .B(n28537), .Z(n28545) );
  AND U29817 ( .A(x[486]), .B(y[7975]), .Z(n29541) );
  AND U29818 ( .A(y[7979]), .B(x[482]), .Z(n28470) );
  NAND U29819 ( .A(y[7972]), .B(x[489]), .Z(n28469) );
  XNOR U29820 ( .A(n28470), .B(n28469), .Z(n28561) );
  XOR U29821 ( .A(n29541), .B(n28561), .Z(n28544) );
  XOR U29822 ( .A(n28545), .B(n28544), .Z(n28546) );
  XOR U29823 ( .A(n28547), .B(n28546), .Z(n28515) );
  NAND U29824 ( .A(n28472), .B(n28471), .Z(n28476) );
  ANDN U29825 ( .B(n28474), .A(n28473), .Z(n28475) );
  ANDN U29826 ( .B(n28476), .A(n28475), .Z(n28514) );
  XOR U29827 ( .A(n28515), .B(n28514), .Z(n28517) );
  XOR U29828 ( .A(n28516), .B(n28517), .Z(n28508) );
  NANDN U29829 ( .A(n28478), .B(n28477), .Z(n28482) );
  NANDN U29830 ( .A(n28480), .B(n28479), .Z(n28481) );
  AND U29831 ( .A(n28482), .B(n28481), .Z(n28523) );
  AND U29832 ( .A(x[486]), .B(y[7979]), .Z(n28920) );
  AND U29833 ( .A(x[481]), .B(y[7974]), .Z(n28536) );
  NAND U29834 ( .A(n28920), .B(n28536), .Z(n28486) );
  NAND U29835 ( .A(n28484), .B(n28483), .Z(n28485) );
  NAND U29836 ( .A(n28486), .B(n28485), .Z(n28529) );
  AND U29837 ( .A(x[492]), .B(y[7980]), .Z(n29795) );
  NAND U29838 ( .A(n29795), .B(n28679), .Z(n28490) );
  NAND U29839 ( .A(n28488), .B(n28487), .Z(n28489) );
  NAND U29840 ( .A(n28490), .B(n28489), .Z(n28527) );
  AND U29841 ( .A(x[490]), .B(y[7971]), .Z(n29390) );
  AND U29842 ( .A(y[7970]), .B(x[491]), .Z(n29351) );
  NAND U29843 ( .A(y[7973]), .B(x[488]), .Z(n28491) );
  XNOR U29844 ( .A(n29351), .B(n28491), .Z(n28533) );
  XOR U29845 ( .A(n29390), .B(n28533), .Z(n28526) );
  XOR U29846 ( .A(n28527), .B(n28526), .Z(n28528) );
  XOR U29847 ( .A(n28529), .B(n28528), .Z(n28521) );
  AND U29848 ( .A(x[490]), .B(y[7976]), .Z(n28493) );
  AND U29849 ( .A(x[484]), .B(y[7970]), .Z(n28492) );
  NAND U29850 ( .A(n28493), .B(n28492), .Z(n28496) );
  NANDN U29851 ( .A(n28494), .B(n29108), .Z(n28495) );
  AND U29852 ( .A(n28496), .B(n28495), .Z(n28572) );
  AND U29853 ( .A(y[7968]), .B(x[493]), .Z(n28498) );
  NAND U29854 ( .A(y[7981]), .B(x[480]), .Z(n28497) );
  XNOR U29855 ( .A(n28498), .B(n28497), .Z(n28555) );
  AND U29856 ( .A(x[492]), .B(y[7969]), .Z(n28566) );
  XOR U29857 ( .A(o[301]), .B(n28566), .Z(n28554) );
  XOR U29858 ( .A(n28555), .B(n28554), .Z(n28570) );
  AND U29859 ( .A(y[7976]), .B(x[485]), .Z(n28500) );
  NAND U29860 ( .A(y[7978]), .B(x[483]), .Z(n28499) );
  XNOR U29861 ( .A(n28500), .B(n28499), .Z(n28550) );
  AND U29862 ( .A(x[484]), .B(y[7977]), .Z(n28551) );
  XOR U29863 ( .A(n28550), .B(n28551), .Z(n28569) );
  XOR U29864 ( .A(n28570), .B(n28569), .Z(n28571) );
  XOR U29865 ( .A(n28521), .B(n28520), .Z(n28522) );
  XOR U29866 ( .A(n28511), .B(n28510), .Z(n28579) );
  NAND U29867 ( .A(n28502), .B(n28501), .Z(n28506) );
  NAND U29868 ( .A(n28504), .B(n28503), .Z(n28505) );
  AND U29869 ( .A(n28506), .B(n28505), .Z(n28578) );
  XOR U29870 ( .A(n28580), .B(n28581), .Z(n28577) );
  XNOR U29871 ( .A(n28575), .B(n28577), .Z(n28507) );
  XOR U29872 ( .A(n28576), .B(n28507), .Z(N622) );
  NANDN U29873 ( .A(n28509), .B(n28508), .Z(n28513) );
  NAND U29874 ( .A(n28511), .B(n28510), .Z(n28512) );
  AND U29875 ( .A(n28513), .B(n28512), .Z(n28668) );
  NAND U29876 ( .A(n28515), .B(n28514), .Z(n28519) );
  NAND U29877 ( .A(n28517), .B(n28516), .Z(n28518) );
  NAND U29878 ( .A(n28519), .B(n28518), .Z(n28667) );
  NAND U29879 ( .A(n28521), .B(n28520), .Z(n28525) );
  NANDN U29880 ( .A(n28523), .B(n28522), .Z(n28524) );
  AND U29881 ( .A(n28525), .B(n28524), .Z(n28588) );
  NAND U29882 ( .A(n28527), .B(n28526), .Z(n28531) );
  NAND U29883 ( .A(n28529), .B(n28528), .Z(n28530) );
  AND U29884 ( .A(n28531), .B(n28530), .Z(n28594) );
  AND U29885 ( .A(x[491]), .B(y[7973]), .Z(n28705) );
  NAND U29886 ( .A(n28705), .B(n28532), .Z(n28535) );
  NAND U29887 ( .A(n28533), .B(n29390), .Z(n28534) );
  NAND U29888 ( .A(n28535), .B(n28534), .Z(n28649) );
  NAND U29889 ( .A(x[487]), .B(y[7980]), .Z(n29123) );
  NANDN U29890 ( .A(n29123), .B(n28536), .Z(n28540) );
  NAND U29891 ( .A(n28538), .B(n28537), .Z(n28539) );
  NAND U29892 ( .A(n28540), .B(n28539), .Z(n28648) );
  XOR U29893 ( .A(n28649), .B(n28648), .Z(n28651) );
  AND U29894 ( .A(x[484]), .B(y[7978]), .Z(n29028) );
  AND U29895 ( .A(y[7979]), .B(x[483]), .Z(n28542) );
  NAND U29896 ( .A(y[7974]), .B(x[488]), .Z(n28541) );
  XNOR U29897 ( .A(n28542), .B(n28541), .Z(n28634) );
  XOR U29898 ( .A(n28919), .B(n28634), .Z(n28643) );
  XOR U29899 ( .A(n29028), .B(n28643), .Z(n28645) );
  AND U29900 ( .A(x[489]), .B(y[7973]), .Z(n29214) );
  AND U29901 ( .A(y[7980]), .B(x[482]), .Z(n28543) );
  AND U29902 ( .A(y[7972]), .B(x[490]), .Z(n29244) );
  XOR U29903 ( .A(n28543), .B(n29244), .Z(n28620) );
  XOR U29904 ( .A(n29214), .B(n28620), .Z(n28644) );
  XOR U29905 ( .A(n28645), .B(n28644), .Z(n28650) );
  XNOR U29906 ( .A(n28651), .B(n28650), .Z(n28592) );
  NAND U29907 ( .A(n28545), .B(n28544), .Z(n28549) );
  NAND U29908 ( .A(n28547), .B(n28546), .Z(n28548) );
  AND U29909 ( .A(n28549), .B(n28548), .Z(n28591) );
  XOR U29910 ( .A(n28592), .B(n28591), .Z(n28593) );
  XOR U29911 ( .A(n28594), .B(n28593), .Z(n28586) );
  NAND U29912 ( .A(x[485]), .B(y[7978]), .Z(n28692) );
  NANDN U29913 ( .A(n28692), .B(n29378), .Z(n28553) );
  NAND U29914 ( .A(n28551), .B(n28550), .Z(n28552) );
  NAND U29915 ( .A(n28553), .B(n28552), .Z(n28600) );
  AND U29916 ( .A(x[493]), .B(y[7981]), .Z(n30129) );
  NAND U29917 ( .A(n30129), .B(n28679), .Z(n28557) );
  NAND U29918 ( .A(n28555), .B(n28554), .Z(n28556) );
  NAND U29919 ( .A(n28557), .B(n28556), .Z(n28598) );
  NAND U29920 ( .A(y[7971]), .B(x[491]), .Z(n28558) );
  XNOR U29921 ( .A(n28559), .B(n28558), .Z(n28624) );
  AND U29922 ( .A(x[481]), .B(y[7981]), .Z(n28625) );
  XOR U29923 ( .A(n28624), .B(n28625), .Z(n28597) );
  XOR U29924 ( .A(n28598), .B(n28597), .Z(n28599) );
  XNOR U29925 ( .A(n28600), .B(n28599), .Z(n28655) );
  AND U29926 ( .A(x[489]), .B(y[7979]), .Z(n28560) );
  NAND U29927 ( .A(n28560), .B(n28619), .Z(n28563) );
  NAND U29928 ( .A(n28561), .B(n29541), .Z(n28562) );
  AND U29929 ( .A(n28563), .B(n28562), .Z(n28606) );
  AND U29930 ( .A(y[7968]), .B(x[494]), .Z(n28565) );
  NAND U29931 ( .A(y[7982]), .B(x[480]), .Z(n28564) );
  XNOR U29932 ( .A(n28565), .B(n28564), .Z(n28629) );
  AND U29933 ( .A(o[301]), .B(n28566), .Z(n28628) );
  XOR U29934 ( .A(n28629), .B(n28628), .Z(n28604) );
  NAND U29935 ( .A(y[7970]), .B(x[492]), .Z(n28567) );
  XNOR U29936 ( .A(n28568), .B(n28567), .Z(n28610) );
  NAND U29937 ( .A(x[493]), .B(y[7969]), .Z(n28618) );
  XNOR U29938 ( .A(o[302]), .B(n28618), .Z(n28611) );
  XOR U29939 ( .A(n28610), .B(n28611), .Z(n28603) );
  XOR U29940 ( .A(n28604), .B(n28603), .Z(n28605) );
  XOR U29941 ( .A(n28606), .B(n28605), .Z(n28654) );
  XOR U29942 ( .A(n28655), .B(n28654), .Z(n28657) );
  NAND U29943 ( .A(n28570), .B(n28569), .Z(n28574) );
  NANDN U29944 ( .A(n28572), .B(n28571), .Z(n28573) );
  AND U29945 ( .A(n28574), .B(n28573), .Z(n28656) );
  XNOR U29946 ( .A(n28657), .B(n28656), .Z(n28585) );
  XNOR U29947 ( .A(n28670), .B(n28669), .Z(n28663) );
  NANDN U29948 ( .A(n28579), .B(n28578), .Z(n28583) );
  NAND U29949 ( .A(n28581), .B(n28580), .Z(n28582) );
  AND U29950 ( .A(n28583), .B(n28582), .Z(n28661) );
  IV U29951 ( .A(n28661), .Z(n28660) );
  XOR U29952 ( .A(n28662), .B(n28660), .Z(n28584) );
  XNOR U29953 ( .A(n28663), .B(n28584), .Z(N623) );
  NANDN U29954 ( .A(n28586), .B(n28585), .Z(n28590) );
  NANDN U29955 ( .A(n28588), .B(n28587), .Z(n28589) );
  AND U29956 ( .A(n28590), .B(n28589), .Z(n28766) );
  NAND U29957 ( .A(n28592), .B(n28591), .Z(n28596) );
  NAND U29958 ( .A(n28594), .B(n28593), .Z(n28595) );
  NAND U29959 ( .A(n28596), .B(n28595), .Z(n28735) );
  NAND U29960 ( .A(n28598), .B(n28597), .Z(n28602) );
  NAND U29961 ( .A(n28600), .B(n28599), .Z(n28601) );
  NAND U29962 ( .A(n28602), .B(n28601), .Z(n28741) );
  NAND U29963 ( .A(n28604), .B(n28603), .Z(n28608) );
  NANDN U29964 ( .A(n28606), .B(n28605), .Z(n28607) );
  NAND U29965 ( .A(n28608), .B(n28607), .Z(n28739) );
  NAND U29966 ( .A(x[492]), .B(y[7975]), .Z(n29115) );
  NANDN U29967 ( .A(n29115), .B(n28609), .Z(n28613) );
  NAND U29968 ( .A(n28611), .B(n28610), .Z(n28612) );
  AND U29969 ( .A(n28613), .B(n28612), .Z(n28715) );
  AND U29970 ( .A(y[7972]), .B(x[491]), .Z(n28615) );
  NAND U29971 ( .A(y[7970]), .B(x[493]), .Z(n28614) );
  XNOR U29972 ( .A(n28615), .B(n28614), .Z(n28719) );
  AND U29973 ( .A(x[492]), .B(y[7971]), .Z(n28718) );
  XNOR U29974 ( .A(n28719), .B(n28718), .Z(n28713) );
  AND U29975 ( .A(y[7968]), .B(x[495]), .Z(n28617) );
  NAND U29976 ( .A(y[7983]), .B(x[480]), .Z(n28616) );
  XNOR U29977 ( .A(n28617), .B(n28616), .Z(n28681) );
  ANDN U29978 ( .B(o[302]), .A(n28618), .Z(n28680) );
  XNOR U29979 ( .A(n28681), .B(n28680), .Z(n28712) );
  XOR U29980 ( .A(n28713), .B(n28712), .Z(n28714) );
  XNOR U29981 ( .A(n28715), .B(n28714), .Z(n28747) );
  NAND U29982 ( .A(x[490]), .B(y[7980]), .Z(n29543) );
  NANDN U29983 ( .A(n29543), .B(n28619), .Z(n28622) );
  NAND U29984 ( .A(n29214), .B(n28620), .Z(n28621) );
  NAND U29985 ( .A(n28622), .B(n28621), .Z(n28745) );
  AND U29986 ( .A(x[491]), .B(y[7976]), .Z(n29027) );
  NAND U29987 ( .A(n29027), .B(n28623), .Z(n28627) );
  NAND U29988 ( .A(n28625), .B(n28624), .Z(n28626) );
  NAND U29989 ( .A(n28627), .B(n28626), .Z(n28744) );
  XOR U29990 ( .A(n28745), .B(n28744), .Z(n28746) );
  XOR U29991 ( .A(n28747), .B(n28746), .Z(n28738) );
  XOR U29992 ( .A(n28739), .B(n28738), .Z(n28740) );
  XNOR U29993 ( .A(n28741), .B(n28740), .Z(n28732) );
  AND U29994 ( .A(x[494]), .B(y[7982]), .Z(n30403) );
  NAND U29995 ( .A(n30403), .B(n28679), .Z(n28631) );
  NAND U29996 ( .A(n28629), .B(n28628), .Z(n28630) );
  NAND U29997 ( .A(n28631), .B(n28630), .Z(n28707) );
  AND U29998 ( .A(x[488]), .B(y[7979]), .Z(n28632) );
  NANDN U29999 ( .A(n28633), .B(n28632), .Z(n28636) );
  NAND U30000 ( .A(n28634), .B(n28919), .Z(n28635) );
  NAND U30001 ( .A(n28636), .B(n28635), .Z(n28706) );
  XOR U30002 ( .A(n28707), .B(n28706), .Z(n28709) );
  AND U30003 ( .A(y[7973]), .B(x[490]), .Z(n28638) );
  NAND U30004 ( .A(y[7979]), .B(x[484]), .Z(n28637) );
  XNOR U30005 ( .A(n28638), .B(n28637), .Z(n28687) );
  AND U30006 ( .A(x[487]), .B(y[7976]), .Z(n28686) );
  XNOR U30007 ( .A(n28687), .B(n28686), .Z(n28694) );
  AND U30008 ( .A(x[486]), .B(y[7977]), .Z(n28797) );
  XNOR U30009 ( .A(n28797), .B(n28692), .Z(n28693) );
  XOR U30010 ( .A(n28694), .B(n28693), .Z(n28729) );
  AND U30011 ( .A(y[7981]), .B(x[482]), .Z(n28640) );
  NAND U30012 ( .A(y[7974]), .B(x[489]), .Z(n28639) );
  XNOR U30013 ( .A(n28640), .B(n28639), .Z(n28697) );
  AND U30014 ( .A(x[483]), .B(y[7980]), .Z(n28698) );
  XOR U30015 ( .A(n28697), .B(n28698), .Z(n28727) );
  AND U30016 ( .A(y[7982]), .B(x[481]), .Z(n28642) );
  NAND U30017 ( .A(y[7975]), .B(x[488]), .Z(n28641) );
  XNOR U30018 ( .A(n28642), .B(n28641), .Z(n28676) );
  NAND U30019 ( .A(x[494]), .B(y[7969]), .Z(n28703) );
  XNOR U30020 ( .A(o[303]), .B(n28703), .Z(n28675) );
  XOR U30021 ( .A(n28676), .B(n28675), .Z(n28726) );
  XOR U30022 ( .A(n28727), .B(n28726), .Z(n28728) );
  XNOR U30023 ( .A(n28709), .B(n28708), .Z(n28751) );
  NAND U30024 ( .A(n29028), .B(n28643), .Z(n28647) );
  NAND U30025 ( .A(n28645), .B(n28644), .Z(n28646) );
  AND U30026 ( .A(n28647), .B(n28646), .Z(n28750) );
  XOR U30027 ( .A(n28751), .B(n28750), .Z(n28752) );
  NAND U30028 ( .A(n28649), .B(n28648), .Z(n28653) );
  NAND U30029 ( .A(n28651), .B(n28650), .Z(n28652) );
  AND U30030 ( .A(n28653), .B(n28652), .Z(n28753) );
  XOR U30031 ( .A(n28752), .B(n28753), .Z(n28733) );
  XOR U30032 ( .A(n28732), .B(n28733), .Z(n28734) );
  XNOR U30033 ( .A(n28735), .B(n28734), .Z(n28763) );
  NAND U30034 ( .A(n28655), .B(n28654), .Z(n28659) );
  NAND U30035 ( .A(n28657), .B(n28656), .Z(n28658) );
  AND U30036 ( .A(n28659), .B(n28658), .Z(n28764) );
  XOR U30037 ( .A(n28763), .B(n28764), .Z(n28765) );
  XOR U30038 ( .A(n28766), .B(n28765), .Z(n28759) );
  OR U30039 ( .A(n28662), .B(n28660), .Z(n28666) );
  ANDN U30040 ( .B(n28662), .A(n28661), .Z(n28664) );
  OR U30041 ( .A(n28664), .B(n28663), .Z(n28665) );
  AND U30042 ( .A(n28666), .B(n28665), .Z(n28758) );
  NANDN U30043 ( .A(n28668), .B(n28667), .Z(n28672) );
  NAND U30044 ( .A(n28670), .B(n28669), .Z(n28671) );
  NAND U30045 ( .A(n28672), .B(n28671), .Z(n28757) );
  IV U30046 ( .A(n28757), .Z(n28756) );
  XOR U30047 ( .A(n28758), .B(n28756), .Z(n28673) );
  XNOR U30048 ( .A(n28759), .B(n28673), .Z(N624) );
  AND U30049 ( .A(x[488]), .B(y[7982]), .Z(n29029) );
  NAND U30050 ( .A(n29029), .B(n28674), .Z(n28678) );
  NAND U30051 ( .A(n28676), .B(n28675), .Z(n28677) );
  AND U30052 ( .A(n28678), .B(n28677), .Z(n28825) );
  AND U30053 ( .A(x[495]), .B(y[7983]), .Z(n30864) );
  NAND U30054 ( .A(n30864), .B(n28679), .Z(n28683) );
  NAND U30055 ( .A(n28681), .B(n28680), .Z(n28682) );
  NAND U30056 ( .A(n28683), .B(n28682), .Z(n28824) );
  XNOR U30057 ( .A(n28825), .B(n28824), .Z(n28827) );
  AND U30058 ( .A(x[490]), .B(y[7979]), .Z(n28685) );
  NAND U30059 ( .A(n28685), .B(n28684), .Z(n28689) );
  NAND U30060 ( .A(n28687), .B(n28686), .Z(n28688) );
  NAND U30061 ( .A(n28689), .B(n28688), .Z(n28784) );
  AND U30062 ( .A(x[480]), .B(y[7984]), .Z(n28804) );
  NAND U30063 ( .A(x[496]), .B(y[7968]), .Z(n28805) );
  XNOR U30064 ( .A(n28804), .B(n28805), .Z(n28806) );
  NAND U30065 ( .A(x[495]), .B(y[7969]), .Z(n28794) );
  XOR U30066 ( .A(o[304]), .B(n28794), .Z(n28807) );
  XNOR U30067 ( .A(n28806), .B(n28807), .Z(n28783) );
  NAND U30068 ( .A(y[7977]), .B(x[487]), .Z(n28690) );
  XNOR U30069 ( .A(n28691), .B(n28690), .Z(n28799) );
  AND U30070 ( .A(x[490]), .B(y[7974]), .Z(n28798) );
  XOR U30071 ( .A(n28799), .B(n28798), .Z(n28782) );
  XOR U30072 ( .A(n28783), .B(n28782), .Z(n28785) );
  XOR U30073 ( .A(n28784), .B(n28785), .Z(n28826) );
  XNOR U30074 ( .A(n28827), .B(n28826), .Z(n28779) );
  NANDN U30075 ( .A(n28797), .B(n28692), .Z(n28696) );
  NAND U30076 ( .A(n28694), .B(n28693), .Z(n28695) );
  NAND U30077 ( .A(n28696), .B(n28695), .Z(n28777) );
  NAND U30078 ( .A(x[489]), .B(y[7981]), .Z(n29513) );
  NANDN U30079 ( .A(n29513), .B(n29113), .Z(n28700) );
  NAND U30080 ( .A(n28698), .B(n28697), .Z(n28699) );
  NAND U30081 ( .A(n28700), .B(n28699), .Z(n28814) );
  AND U30082 ( .A(y[7983]), .B(x[481]), .Z(n28702) );
  NAND U30083 ( .A(y[7976]), .B(x[488]), .Z(n28701) );
  XNOR U30084 ( .A(n28702), .B(n28701), .Z(n28803) );
  ANDN U30085 ( .B(o[303]), .A(n28703), .Z(n28802) );
  XOR U30086 ( .A(n28803), .B(n28802), .Z(n28813) );
  NAND U30087 ( .A(y[7970]), .B(x[494]), .Z(n28704) );
  XNOR U30088 ( .A(n28705), .B(n28704), .Z(n28836) );
  NAND U30089 ( .A(x[484]), .B(y[7980]), .Z(n28837) );
  XNOR U30090 ( .A(n28836), .B(n28837), .Z(n28812) );
  XOR U30091 ( .A(n28813), .B(n28812), .Z(n28815) );
  XNOR U30092 ( .A(n28814), .B(n28815), .Z(n28776) );
  XOR U30093 ( .A(n28777), .B(n28776), .Z(n28778) );
  XOR U30094 ( .A(n28779), .B(n28778), .Z(n28818) );
  NAND U30095 ( .A(n28707), .B(n28706), .Z(n28711) );
  NAND U30096 ( .A(n28709), .B(n28708), .Z(n28710) );
  AND U30097 ( .A(n28711), .B(n28710), .Z(n28819) );
  XOR U30098 ( .A(n28818), .B(n28819), .Z(n28821) );
  NAND U30099 ( .A(n28713), .B(n28712), .Z(n28717) );
  NAND U30100 ( .A(n28715), .B(n28714), .Z(n28716) );
  NAND U30101 ( .A(n28717), .B(n28716), .Z(n28849) );
  AND U30102 ( .A(x[493]), .B(y[7972]), .Z(n28846) );
  NAND U30103 ( .A(n29351), .B(n28846), .Z(n28721) );
  NAND U30104 ( .A(n28719), .B(n28718), .Z(n28720) );
  AND U30105 ( .A(n28721), .B(n28720), .Z(n28833) );
  AND U30106 ( .A(y[7982]), .B(x[482]), .Z(n28723) );
  NAND U30107 ( .A(y[7975]), .B(x[489]), .Z(n28722) );
  XNOR U30108 ( .A(n28723), .B(n28722), .Z(n28840) );
  NAND U30109 ( .A(x[483]), .B(y[7981]), .Z(n28841) );
  XNOR U30110 ( .A(n28840), .B(n28841), .Z(n28830) );
  AND U30111 ( .A(x[492]), .B(y[7972]), .Z(n29518) );
  AND U30112 ( .A(y[7979]), .B(x[485]), .Z(n28725) );
  NAND U30113 ( .A(y[7971]), .B(x[493]), .Z(n28724) );
  XOR U30114 ( .A(n28725), .B(n28724), .Z(n28789) );
  XOR U30115 ( .A(n29518), .B(n28789), .Z(n28831) );
  XNOR U30116 ( .A(n28830), .B(n28831), .Z(n28832) );
  XOR U30117 ( .A(n28833), .B(n28832), .Z(n28847) );
  NAND U30118 ( .A(n28727), .B(n28726), .Z(n28731) );
  NANDN U30119 ( .A(n28729), .B(n28728), .Z(n28730) );
  AND U30120 ( .A(n28731), .B(n28730), .Z(n28848) );
  XOR U30121 ( .A(n28847), .B(n28848), .Z(n28850) );
  XOR U30122 ( .A(n28849), .B(n28850), .Z(n28820) );
  XNOR U30123 ( .A(n28821), .B(n28820), .Z(n28861) );
  NAND U30124 ( .A(n28733), .B(n28732), .Z(n28737) );
  NAND U30125 ( .A(n28735), .B(n28734), .Z(n28736) );
  AND U30126 ( .A(n28737), .B(n28736), .Z(n28860) );
  XOR U30127 ( .A(n28861), .B(n28860), .Z(n28863) );
  NAND U30128 ( .A(n28739), .B(n28738), .Z(n28743) );
  NAND U30129 ( .A(n28741), .B(n28740), .Z(n28742) );
  NAND U30130 ( .A(n28743), .B(n28742), .Z(n28773) );
  NAND U30131 ( .A(n28745), .B(n28744), .Z(n28749) );
  NAND U30132 ( .A(n28747), .B(n28746), .Z(n28748) );
  NAND U30133 ( .A(n28749), .B(n28748), .Z(n28771) );
  NAND U30134 ( .A(n28751), .B(n28750), .Z(n28755) );
  NAND U30135 ( .A(n28753), .B(n28752), .Z(n28754) );
  AND U30136 ( .A(n28755), .B(n28754), .Z(n28770) );
  XOR U30137 ( .A(n28771), .B(n28770), .Z(n28772) );
  XOR U30138 ( .A(n28773), .B(n28772), .Z(n28862) );
  XNOR U30139 ( .A(n28863), .B(n28862), .Z(n28856) );
  OR U30140 ( .A(n28758), .B(n28756), .Z(n28762) );
  ANDN U30141 ( .B(n28758), .A(n28757), .Z(n28760) );
  OR U30142 ( .A(n28760), .B(n28759), .Z(n28761) );
  AND U30143 ( .A(n28762), .B(n28761), .Z(n28855) );
  NAND U30144 ( .A(n28764), .B(n28763), .Z(n28768) );
  NANDN U30145 ( .A(n28766), .B(n28765), .Z(n28767) );
  NAND U30146 ( .A(n28768), .B(n28767), .Z(n28854) );
  IV U30147 ( .A(n28854), .Z(n28853) );
  XOR U30148 ( .A(n28855), .B(n28853), .Z(n28769) );
  XNOR U30149 ( .A(n28856), .B(n28769), .Z(N625) );
  NAND U30150 ( .A(n28771), .B(n28770), .Z(n28775) );
  NAND U30151 ( .A(n28773), .B(n28772), .Z(n28774) );
  NAND U30152 ( .A(n28775), .B(n28774), .Z(n28960) );
  NAND U30153 ( .A(n28777), .B(n28776), .Z(n28781) );
  NAND U30154 ( .A(n28779), .B(n28778), .Z(n28780) );
  NAND U30155 ( .A(n28781), .B(n28780), .Z(n28875) );
  NAND U30156 ( .A(n28783), .B(n28782), .Z(n28787) );
  NAND U30157 ( .A(n28785), .B(n28784), .Z(n28786) );
  AND U30158 ( .A(n28787), .B(n28786), .Z(n28954) );
  AND U30159 ( .A(x[493]), .B(y[7979]), .Z(n29803) );
  NAND U30160 ( .A(n29803), .B(n28788), .Z(n28791) );
  NANDN U30161 ( .A(n28789), .B(n29518), .Z(n28790) );
  AND U30162 ( .A(n28791), .B(n28790), .Z(n28906) );
  AND U30163 ( .A(y[7984]), .B(x[481]), .Z(n28793) );
  NAND U30164 ( .A(y[7976]), .B(x[489]), .Z(n28792) );
  XNOR U30165 ( .A(n28793), .B(n28792), .Z(n28925) );
  ANDN U30166 ( .B(o[304]), .A(n28794), .Z(n28924) );
  XOR U30167 ( .A(n28925), .B(n28924), .Z(n28904) );
  AND U30168 ( .A(y[7970]), .B(x[495]), .Z(n28796) );
  NAND U30169 ( .A(y[7973]), .B(x[492]), .Z(n28795) );
  XNOR U30170 ( .A(n28796), .B(n28795), .Z(n28880) );
  AND U30171 ( .A(x[494]), .B(y[7971]), .Z(n28879) );
  XOR U30172 ( .A(n28880), .B(n28879), .Z(n28903) );
  XOR U30173 ( .A(n28904), .B(n28903), .Z(n28905) );
  XNOR U30174 ( .A(n28906), .B(n28905), .Z(n28951) );
  NAND U30175 ( .A(x[487]), .B(y[7978]), .Z(n28934) );
  NANDN U30176 ( .A(n28934), .B(n28797), .Z(n28801) );
  NAND U30177 ( .A(n28799), .B(n28798), .Z(n28800) );
  AND U30178 ( .A(n28801), .B(n28800), .Z(n28914) );
  AND U30179 ( .A(x[488]), .B(y[7983]), .Z(n29601) );
  AND U30180 ( .A(x[481]), .B(y[7976]), .Z(n29007) );
  XNOR U30181 ( .A(n28914), .B(n28913), .Z(n28915) );
  NANDN U30182 ( .A(n28805), .B(n28804), .Z(n28809) );
  NANDN U30183 ( .A(n28807), .B(n28806), .Z(n28808) );
  AND U30184 ( .A(n28809), .B(n28808), .Z(n28910) );
  AND U30185 ( .A(x[480]), .B(y[7985]), .Z(n28894) );
  AND U30186 ( .A(x[497]), .B(y[7968]), .Z(n28893) );
  XOR U30187 ( .A(n28894), .B(n28893), .Z(n28896) );
  AND U30188 ( .A(x[496]), .B(y[7969]), .Z(n28890) );
  XOR U30189 ( .A(n28890), .B(o[305]), .Z(n28895) );
  XOR U30190 ( .A(n28896), .B(n28895), .Z(n28907) );
  AND U30191 ( .A(y[7983]), .B(x[482]), .Z(n28811) );
  NAND U30192 ( .A(y[7975]), .B(x[490]), .Z(n28810) );
  XNOR U30193 ( .A(n28811), .B(n28810), .Z(n28927) );
  NAND U30194 ( .A(x[483]), .B(y[7982]), .Z(n28928) );
  XOR U30195 ( .A(n28927), .B(n28928), .Z(n28908) );
  XNOR U30196 ( .A(n28907), .B(n28908), .Z(n28909) );
  XOR U30197 ( .A(n28910), .B(n28909), .Z(n28916) );
  XOR U30198 ( .A(n28915), .B(n28916), .Z(n28952) );
  XNOR U30199 ( .A(n28951), .B(n28952), .Z(n28953) );
  XOR U30200 ( .A(n28954), .B(n28953), .Z(n28873) );
  NAND U30201 ( .A(n28813), .B(n28812), .Z(n28817) );
  NAND U30202 ( .A(n28815), .B(n28814), .Z(n28816) );
  AND U30203 ( .A(n28817), .B(n28816), .Z(n28874) );
  XNOR U30204 ( .A(n28873), .B(n28874), .Z(n28876) );
  NAND U30205 ( .A(n28819), .B(n28818), .Z(n28823) );
  NAND U30206 ( .A(n28821), .B(n28820), .Z(n28822) );
  NAND U30207 ( .A(n28823), .B(n28822), .Z(n28869) );
  NANDN U30208 ( .A(n28825), .B(n28824), .Z(n28829) );
  NAND U30209 ( .A(n28827), .B(n28826), .Z(n28828) );
  AND U30210 ( .A(n28829), .B(n28828), .Z(n28948) );
  NANDN U30211 ( .A(n28831), .B(n28830), .Z(n28835) );
  NANDN U30212 ( .A(n28833), .B(n28832), .Z(n28834) );
  AND U30213 ( .A(n28835), .B(n28834), .Z(n28946) );
  NAND U30214 ( .A(x[494]), .B(y[7973]), .Z(n29147) );
  NANDN U30215 ( .A(n29147), .B(n29351), .Z(n28839) );
  NANDN U30216 ( .A(n28837), .B(n28836), .Z(n28838) );
  AND U30217 ( .A(n28839), .B(n28838), .Z(n28940) );
  AND U30218 ( .A(x[489]), .B(y[7982]), .Z(n29784) );
  NAND U30219 ( .A(n28926), .B(n29784), .Z(n28843) );
  NANDN U30220 ( .A(n28841), .B(n28840), .Z(n28842) );
  NAND U30221 ( .A(n28843), .B(n28842), .Z(n28939) );
  XNOR U30222 ( .A(n28940), .B(n28939), .Z(n28941) );
  AND U30223 ( .A(x[485]), .B(y[7980]), .Z(n28989) );
  NAND U30224 ( .A(y[7977]), .B(x[488]), .Z(n28844) );
  XNOR U30225 ( .A(n28989), .B(n28844), .Z(n28921) );
  XOR U30226 ( .A(n28921), .B(n28920), .Z(n28933) );
  NAND U30227 ( .A(y[7981]), .B(x[484]), .Z(n28845) );
  XNOR U30228 ( .A(n28846), .B(n28845), .Z(n28884) );
  NAND U30229 ( .A(x[491]), .B(y[7974]), .Z(n28885) );
  XOR U30230 ( .A(n28884), .B(n28885), .Z(n28936) );
  XOR U30231 ( .A(n28935), .B(n28936), .Z(n28942) );
  XNOR U30232 ( .A(n28941), .B(n28942), .Z(n28945) );
  XNOR U30233 ( .A(n28946), .B(n28945), .Z(n28947) );
  XOR U30234 ( .A(n28948), .B(n28947), .Z(n28868) );
  NAND U30235 ( .A(n28848), .B(n28847), .Z(n28852) );
  NAND U30236 ( .A(n28850), .B(n28849), .Z(n28851) );
  NAND U30237 ( .A(n28852), .B(n28851), .Z(n28867) );
  XNOR U30238 ( .A(n28868), .B(n28867), .Z(n28870) );
  XOR U30239 ( .A(n28869), .B(n28870), .Z(n28957) );
  XOR U30240 ( .A(n28958), .B(n28957), .Z(n28959) );
  XOR U30241 ( .A(n28960), .B(n28959), .Z(n28966) );
  OR U30242 ( .A(n28855), .B(n28853), .Z(n28859) );
  ANDN U30243 ( .B(n28855), .A(n28854), .Z(n28857) );
  OR U30244 ( .A(n28857), .B(n28856), .Z(n28858) );
  AND U30245 ( .A(n28859), .B(n28858), .Z(n28964) );
  NAND U30246 ( .A(n28861), .B(n28860), .Z(n28865) );
  NAND U30247 ( .A(n28863), .B(n28862), .Z(n28864) );
  AND U30248 ( .A(n28865), .B(n28864), .Z(n28965) );
  IV U30249 ( .A(n28965), .Z(n28963) );
  XOR U30250 ( .A(n28964), .B(n28963), .Z(n28866) );
  XNOR U30251 ( .A(n28966), .B(n28866), .Z(N626) );
  NAND U30252 ( .A(n28868), .B(n28867), .Z(n28872) );
  NANDN U30253 ( .A(n28870), .B(n28869), .Z(n28871) );
  AND U30254 ( .A(n28872), .B(n28871), .Z(n29076) );
  NAND U30255 ( .A(n28874), .B(n28873), .Z(n28878) );
  NANDN U30256 ( .A(n28876), .B(n28875), .Z(n28877) );
  AND U30257 ( .A(n28878), .B(n28877), .Z(n29074) );
  AND U30258 ( .A(x[495]), .B(y[7973]), .Z(n29121) );
  AND U30259 ( .A(x[492]), .B(y[7970]), .Z(n29204) );
  NAND U30260 ( .A(n29121), .B(n29204), .Z(n28882) );
  NAND U30261 ( .A(n28880), .B(n28879), .Z(n28881) );
  NAND U30262 ( .A(n28882), .B(n28881), .Z(n29055) );
  NAND U30263 ( .A(n30129), .B(n28883), .Z(n28887) );
  NANDN U30264 ( .A(n28885), .B(n28884), .Z(n28886) );
  AND U30265 ( .A(n28887), .B(n28886), .Z(n29046) );
  AND U30266 ( .A(y[7985]), .B(x[481]), .Z(n28889) );
  NAND U30267 ( .A(y[7976]), .B(x[490]), .Z(n28888) );
  XNOR U30268 ( .A(n28889), .B(n28888), .Z(n29008) );
  NAND U30269 ( .A(n28890), .B(o[305]), .Z(n29009) );
  XNOR U30270 ( .A(n29008), .B(n29009), .Z(n29043) );
  AND U30271 ( .A(y[7971]), .B(x[495]), .Z(n28892) );
  NAND U30272 ( .A(y[7977]), .B(x[489]), .Z(n28891) );
  XNOR U30273 ( .A(n28892), .B(n28891), .Z(n28999) );
  NAND U30274 ( .A(x[494]), .B(y[7972]), .Z(n29000) );
  XOR U30275 ( .A(n28999), .B(n29000), .Z(n29044) );
  XNOR U30276 ( .A(n29043), .B(n29044), .Z(n29045) );
  XNOR U30277 ( .A(n29046), .B(n29045), .Z(n29056) );
  XOR U30278 ( .A(n29055), .B(n29056), .Z(n29058) );
  NAND U30279 ( .A(n28894), .B(n28893), .Z(n28898) );
  NAND U30280 ( .A(n28896), .B(n28895), .Z(n28897) );
  NAND U30281 ( .A(n28898), .B(n28897), .Z(n29067) );
  AND U30282 ( .A(y[7970]), .B(x[496]), .Z(n28900) );
  NAND U30283 ( .A(y[7975]), .B(x[491]), .Z(n28899) );
  XNOR U30284 ( .A(n28900), .B(n28899), .Z(n28995) );
  NAND U30285 ( .A(x[482]), .B(y[7984]), .Z(n28996) );
  XNOR U30286 ( .A(n28995), .B(n28996), .Z(n29068) );
  XOR U30287 ( .A(n29067), .B(n29068), .Z(n29070) );
  AND U30288 ( .A(y[7981]), .B(x[485]), .Z(n29129) );
  NAND U30289 ( .A(y[7980]), .B(x[486]), .Z(n28901) );
  XNOR U30290 ( .A(n29129), .B(n28901), .Z(n28992) );
  NAND U30291 ( .A(y[7982]), .B(x[484]), .Z(n28902) );
  XNOR U30292 ( .A(n29789), .B(n28902), .Z(n29030) );
  AND U30293 ( .A(x[487]), .B(y[7979]), .Z(n29031) );
  XOR U30294 ( .A(n29030), .B(n29031), .Z(n28991) );
  XOR U30295 ( .A(n28992), .B(n28991), .Z(n29069) );
  XOR U30296 ( .A(n29070), .B(n29069), .Z(n29057) );
  XOR U30297 ( .A(n29058), .B(n29057), .Z(n28978) );
  NANDN U30298 ( .A(n28908), .B(n28907), .Z(n28912) );
  NANDN U30299 ( .A(n28910), .B(n28909), .Z(n28911) );
  AND U30300 ( .A(n28912), .B(n28911), .Z(n29049) );
  XOR U30301 ( .A(n29050), .B(n29049), .Z(n29052) );
  NANDN U30302 ( .A(n28914), .B(n28913), .Z(n28918) );
  NANDN U30303 ( .A(n28916), .B(n28915), .Z(n28917) );
  AND U30304 ( .A(n28918), .B(n28917), .Z(n29051) );
  XOR U30305 ( .A(n29052), .B(n29051), .Z(n28977) );
  XNOR U30306 ( .A(n28978), .B(n28977), .Z(n28980) );
  AND U30307 ( .A(x[488]), .B(y[7980]), .Z(n29250) );
  NAND U30308 ( .A(n29250), .B(n28919), .Z(n28923) );
  NAND U30309 ( .A(n28921), .B(n28920), .Z(n28922) );
  NAND U30310 ( .A(n28923), .B(n28922), .Z(n29062) );
  AND U30311 ( .A(x[489]), .B(y[7984]), .Z(n29912) );
  XOR U30312 ( .A(n29062), .B(n29061), .Z(n29064) );
  AND U30313 ( .A(x[490]), .B(y[7983]), .Z(n29812) );
  IV U30314 ( .A(n29812), .Z(n29911) );
  NANDN U30315 ( .A(n29911), .B(n28926), .Z(n28930) );
  NANDN U30316 ( .A(n28928), .B(n28927), .Z(n28929) );
  AND U30317 ( .A(n28930), .B(n28929), .Z(n29040) );
  AND U30318 ( .A(x[480]), .B(y[7986]), .Z(n29012) );
  NAND U30319 ( .A(x[498]), .B(y[7968]), .Z(n29013) );
  XNOR U30320 ( .A(n29012), .B(n29013), .Z(n29014) );
  NAND U30321 ( .A(x[497]), .B(y[7969]), .Z(n29034) );
  XOR U30322 ( .A(o[306]), .B(n29034), .Z(n29015) );
  XNOR U30323 ( .A(n29014), .B(n29015), .Z(n29037) );
  AND U30324 ( .A(y[7973]), .B(x[493]), .Z(n28932) );
  NAND U30325 ( .A(y[7983]), .B(x[483]), .Z(n28931) );
  XNOR U30326 ( .A(n28932), .B(n28931), .Z(n29020) );
  NAND U30327 ( .A(x[492]), .B(y[7974]), .Z(n29021) );
  XOR U30328 ( .A(n29020), .B(n29021), .Z(n29038) );
  XNOR U30329 ( .A(n29037), .B(n29038), .Z(n29039) );
  XNOR U30330 ( .A(n29040), .B(n29039), .Z(n29063) );
  XOR U30331 ( .A(n29064), .B(n29063), .Z(n28984) );
  NANDN U30332 ( .A(n28934), .B(n28933), .Z(n28938) );
  NANDN U30333 ( .A(n28936), .B(n28935), .Z(n28937) );
  AND U30334 ( .A(n28938), .B(n28937), .Z(n28983) );
  XNOR U30335 ( .A(n28984), .B(n28983), .Z(n28985) );
  NANDN U30336 ( .A(n28940), .B(n28939), .Z(n28944) );
  NANDN U30337 ( .A(n28942), .B(n28941), .Z(n28943) );
  NAND U30338 ( .A(n28944), .B(n28943), .Z(n28986) );
  XNOR U30339 ( .A(n28985), .B(n28986), .Z(n28979) );
  XOR U30340 ( .A(n28980), .B(n28979), .Z(n28973) );
  NANDN U30341 ( .A(n28946), .B(n28945), .Z(n28950) );
  NANDN U30342 ( .A(n28948), .B(n28947), .Z(n28949) );
  AND U30343 ( .A(n28950), .B(n28949), .Z(n28972) );
  NANDN U30344 ( .A(n28952), .B(n28951), .Z(n28956) );
  NANDN U30345 ( .A(n28954), .B(n28953), .Z(n28955) );
  NAND U30346 ( .A(n28956), .B(n28955), .Z(n28971) );
  XOR U30347 ( .A(n28972), .B(n28971), .Z(n28974) );
  XOR U30348 ( .A(n28973), .B(n28974), .Z(n29073) );
  XOR U30349 ( .A(n29074), .B(n29073), .Z(n29075) );
  XNOR U30350 ( .A(n29076), .B(n29075), .Z(n29081) );
  NAND U30351 ( .A(n28958), .B(n28957), .Z(n28962) );
  NAND U30352 ( .A(n28960), .B(n28959), .Z(n28961) );
  NAND U30353 ( .A(n28962), .B(n28961), .Z(n29080) );
  NANDN U30354 ( .A(n28963), .B(n28964), .Z(n28969) );
  NOR U30355 ( .A(n28965), .B(n28964), .Z(n28967) );
  OR U30356 ( .A(n28967), .B(n28966), .Z(n28968) );
  AND U30357 ( .A(n28969), .B(n28968), .Z(n29079) );
  XOR U30358 ( .A(n29080), .B(n29079), .Z(n28970) );
  XNOR U30359 ( .A(n29081), .B(n28970), .Z(N627) );
  NANDN U30360 ( .A(n28972), .B(n28971), .Z(n28976) );
  OR U30361 ( .A(n28974), .B(n28973), .Z(n28975) );
  AND U30362 ( .A(n28976), .B(n28975), .Z(n29089) );
  NANDN U30363 ( .A(n28978), .B(n28977), .Z(n28982) );
  NAND U30364 ( .A(n28980), .B(n28979), .Z(n28981) );
  AND U30365 ( .A(n28982), .B(n28981), .Z(n29087) );
  NANDN U30366 ( .A(n28984), .B(n28983), .Z(n28988) );
  NANDN U30367 ( .A(n28986), .B(n28985), .Z(n28987) );
  AND U30368 ( .A(n28988), .B(n28987), .Z(n29093) );
  AND U30369 ( .A(x[486]), .B(y[7981]), .Z(n28990) );
  NAND U30370 ( .A(n28990), .B(n28989), .Z(n28994) );
  NAND U30371 ( .A(n28992), .B(n28991), .Z(n28993) );
  AND U30372 ( .A(n28994), .B(n28993), .Z(n29181) );
  AND U30373 ( .A(x[496]), .B(y[7975]), .Z(n29517) );
  NAND U30374 ( .A(n29517), .B(n29351), .Z(n28998) );
  NANDN U30375 ( .A(n28996), .B(n28995), .Z(n28997) );
  AND U30376 ( .A(n28998), .B(n28997), .Z(n29180) );
  AND U30377 ( .A(x[495]), .B(y[7977]), .Z(n29817) );
  NAND U30378 ( .A(n29817), .B(n29108), .Z(n29002) );
  NANDN U30379 ( .A(n29000), .B(n28999), .Z(n29001) );
  NAND U30380 ( .A(n29002), .B(n29001), .Z(n29099) );
  AND U30381 ( .A(y[7986]), .B(x[481]), .Z(n29004) );
  NAND U30382 ( .A(y[7979]), .B(x[488]), .Z(n29003) );
  XNOR U30383 ( .A(n29004), .B(n29003), .Z(n29146) );
  AND U30384 ( .A(y[7974]), .B(x[493]), .Z(n29006) );
  NAND U30385 ( .A(y[7985]), .B(x[482]), .Z(n29005) );
  XNOR U30386 ( .A(n29006), .B(n29005), .Z(n29114) );
  XOR U30387 ( .A(n29097), .B(n29096), .Z(n29098) );
  XOR U30388 ( .A(n29099), .B(n29098), .Z(n29179) );
  XOR U30389 ( .A(n29180), .B(n29179), .Z(n29182) );
  XOR U30390 ( .A(n29181), .B(n29182), .Z(n29091) );
  AND U30391 ( .A(x[490]), .B(y[7985]), .Z(n30230) );
  NAND U30392 ( .A(n30230), .B(n29007), .Z(n29011) );
  NANDN U30393 ( .A(n29009), .B(n29008), .Z(n29010) );
  NAND U30394 ( .A(n29011), .B(n29010), .Z(n29158) );
  NANDN U30395 ( .A(n29013), .B(n29012), .Z(n29017) );
  NANDN U30396 ( .A(n29015), .B(n29014), .Z(n29016) );
  NAND U30397 ( .A(n29017), .B(n29016), .Z(n29156) );
  AND U30398 ( .A(y[7971]), .B(x[496]), .Z(n29755) );
  NAND U30399 ( .A(y[7978]), .B(x[489]), .Z(n29018) );
  XNOR U30400 ( .A(n29755), .B(n29018), .Z(n29109) );
  NAND U30401 ( .A(x[495]), .B(y[7972]), .Z(n29110) );
  XOR U30402 ( .A(n29156), .B(n29155), .Z(n29157) );
  XNOR U30403 ( .A(n29158), .B(n29157), .Z(n29175) );
  AND U30404 ( .A(x[493]), .B(y[7983]), .Z(n30430) );
  NANDN U30405 ( .A(n29019), .B(n30430), .Z(n29023) );
  NANDN U30406 ( .A(n29021), .B(n29020), .Z(n29022) );
  NAND U30407 ( .A(n29023), .B(n29022), .Z(n29164) );
  AND U30408 ( .A(y[7977]), .B(x[490]), .Z(n29025) );
  NAND U30409 ( .A(y[7970]), .B(x[497]), .Z(n29024) );
  XNOR U30410 ( .A(n29025), .B(n29024), .Z(n29152) );
  AND U30411 ( .A(x[498]), .B(y[7969]), .Z(n29128) );
  XOR U30412 ( .A(o[307]), .B(n29128), .Z(n29151) );
  XOR U30413 ( .A(n29152), .B(n29151), .Z(n29162) );
  NAND U30414 ( .A(y[7984]), .B(x[483]), .Z(n29026) );
  XNOR U30415 ( .A(n29027), .B(n29026), .Z(n29122) );
  XOR U30416 ( .A(n29162), .B(n29161), .Z(n29163) );
  XNOR U30417 ( .A(n29164), .B(n29163), .Z(n29174) );
  NAND U30418 ( .A(n29029), .B(n29028), .Z(n29033) );
  NAND U30419 ( .A(n29031), .B(n29030), .Z(n29032) );
  AND U30420 ( .A(n29033), .B(n29032), .Z(n29105) );
  AND U30421 ( .A(x[480]), .B(y[7987]), .Z(n29133) );
  AND U30422 ( .A(x[499]), .B(y[7968]), .Z(n29134) );
  XOR U30423 ( .A(n29133), .B(n29134), .Z(n29136) );
  ANDN U30424 ( .B(o[306]), .A(n29034), .Z(n29135) );
  XOR U30425 ( .A(n29136), .B(n29135), .Z(n29103) );
  AND U30426 ( .A(x[484]), .B(y[7983]), .Z(n29264) );
  AND U30427 ( .A(y[7982]), .B(x[485]), .Z(n29036) );
  NAND U30428 ( .A(y[7981]), .B(x[486]), .Z(n29035) );
  XNOR U30429 ( .A(n29036), .B(n29035), .Z(n29130) );
  XOR U30430 ( .A(n29264), .B(n29130), .Z(n29102) );
  XOR U30431 ( .A(n29103), .B(n29102), .Z(n29104) );
  XOR U30432 ( .A(n29105), .B(n29104), .Z(n29173) );
  XNOR U30433 ( .A(n29174), .B(n29173), .Z(n29176) );
  XOR U30434 ( .A(n29175), .B(n29176), .Z(n29169) );
  NANDN U30435 ( .A(n29038), .B(n29037), .Z(n29042) );
  NANDN U30436 ( .A(n29040), .B(n29039), .Z(n29041) );
  AND U30437 ( .A(n29042), .B(n29041), .Z(n29168) );
  NANDN U30438 ( .A(n29044), .B(n29043), .Z(n29048) );
  NANDN U30439 ( .A(n29046), .B(n29045), .Z(n29047) );
  NAND U30440 ( .A(n29048), .B(n29047), .Z(n29167) );
  XOR U30441 ( .A(n29168), .B(n29167), .Z(n29170) );
  XOR U30442 ( .A(n29169), .B(n29170), .Z(n29090) );
  XNOR U30443 ( .A(n29091), .B(n29090), .Z(n29092) );
  XOR U30444 ( .A(n29093), .B(n29092), .Z(n29193) );
  NAND U30445 ( .A(n29050), .B(n29049), .Z(n29054) );
  NAND U30446 ( .A(n29052), .B(n29051), .Z(n29053) );
  AND U30447 ( .A(n29054), .B(n29053), .Z(n29191) );
  NAND U30448 ( .A(n29056), .B(n29055), .Z(n29060) );
  NAND U30449 ( .A(n29058), .B(n29057), .Z(n29059) );
  NAND U30450 ( .A(n29060), .B(n29059), .Z(n29187) );
  NAND U30451 ( .A(n29062), .B(n29061), .Z(n29066) );
  NAND U30452 ( .A(n29064), .B(n29063), .Z(n29065) );
  NAND U30453 ( .A(n29066), .B(n29065), .Z(n29186) );
  NAND U30454 ( .A(n29068), .B(n29067), .Z(n29072) );
  NAND U30455 ( .A(n29070), .B(n29069), .Z(n29071) );
  NAND U30456 ( .A(n29072), .B(n29071), .Z(n29185) );
  XNOR U30457 ( .A(n29186), .B(n29185), .Z(n29188) );
  XNOR U30458 ( .A(n29191), .B(n29192), .Z(n29194) );
  XOR U30459 ( .A(n29193), .B(n29194), .Z(n29086) );
  XOR U30460 ( .A(n29087), .B(n29086), .Z(n29088) );
  XNOR U30461 ( .A(n29089), .B(n29088), .Z(n29085) );
  NAND U30462 ( .A(n29074), .B(n29073), .Z(n29078) );
  NAND U30463 ( .A(n29076), .B(n29075), .Z(n29077) );
  AND U30464 ( .A(n29078), .B(n29077), .Z(n29084) );
  XNOR U30465 ( .A(n29084), .B(n29083), .Z(n29082) );
  XNOR U30466 ( .A(n29085), .B(n29082), .Z(N628) );
  NANDN U30467 ( .A(n29091), .B(n29090), .Z(n29095) );
  NANDN U30468 ( .A(n29093), .B(n29092), .Z(n29094) );
  AND U30469 ( .A(n29095), .B(n29094), .Z(n29301) );
  NAND U30470 ( .A(n29097), .B(n29096), .Z(n29101) );
  NAND U30471 ( .A(n29099), .B(n29098), .Z(n29100) );
  NAND U30472 ( .A(n29101), .B(n29100), .Z(n29199) );
  NAND U30473 ( .A(n29103), .B(n29102), .Z(n29107) );
  NANDN U30474 ( .A(n29105), .B(n29104), .Z(n29106) );
  NAND U30475 ( .A(n29107), .B(n29106), .Z(n29198) );
  XOR U30476 ( .A(n29199), .B(n29198), .Z(n29201) );
  AND U30477 ( .A(x[496]), .B(y[7978]), .Z(n30046) );
  NAND U30478 ( .A(n30046), .B(n29108), .Z(n29112) );
  NANDN U30479 ( .A(n29110), .B(n29109), .Z(n29111) );
  AND U30480 ( .A(n29112), .B(n29111), .Z(n29239) );
  AND U30481 ( .A(x[493]), .B(y[7985]), .Z(n30673) );
  NAND U30482 ( .A(n30673), .B(n29113), .Z(n29117) );
  NANDN U30483 ( .A(n29115), .B(n29114), .Z(n29116) );
  AND U30484 ( .A(n29117), .B(n29116), .Z(n29284) );
  AND U30485 ( .A(y[7972]), .B(x[496]), .Z(n29119) );
  NAND U30486 ( .A(y[7978]), .B(x[490]), .Z(n29118) );
  XNOR U30487 ( .A(n29119), .B(n29118), .Z(n29245) );
  AND U30488 ( .A(x[482]), .B(y[7986]), .Z(n29246) );
  XOR U30489 ( .A(n29245), .B(n29246), .Z(n29282) );
  NAND U30490 ( .A(y[7979]), .B(x[489]), .Z(n29120) );
  XNOR U30491 ( .A(n29121), .B(n29120), .Z(n29215) );
  AND U30492 ( .A(x[494]), .B(y[7974]), .Z(n29216) );
  XOR U30493 ( .A(n29215), .B(n29216), .Z(n29281) );
  XOR U30494 ( .A(n29282), .B(n29281), .Z(n29283) );
  AND U30495 ( .A(x[491]), .B(y[7984]), .Z(n30232) );
  IV U30496 ( .A(n30232), .Z(n30094) );
  NANDN U30497 ( .A(n30094), .B(n29378), .Z(n29125) );
  NANDN U30498 ( .A(n29123), .B(n29122), .Z(n29124) );
  AND U30499 ( .A(n29125), .B(n29124), .Z(n29290) );
  AND U30500 ( .A(y[7977]), .B(x[491]), .Z(n29127) );
  NAND U30501 ( .A(y[7987]), .B(x[481]), .Z(n29126) );
  XNOR U30502 ( .A(n29127), .B(n29126), .Z(n29211) );
  AND U30503 ( .A(x[499]), .B(y[7969]), .Z(n29219) );
  XOR U30504 ( .A(o[308]), .B(n29219), .Z(n29210) );
  XOR U30505 ( .A(n29211), .B(n29210), .Z(n29288) );
  AND U30506 ( .A(x[480]), .B(y[7988]), .Z(n29269) );
  AND U30507 ( .A(x[500]), .B(y[7968]), .Z(n29270) );
  XOR U30508 ( .A(n29269), .B(n29270), .Z(n29272) );
  AND U30509 ( .A(o[307]), .B(n29128), .Z(n29271) );
  XOR U30510 ( .A(n29272), .B(n29271), .Z(n29287) );
  XOR U30511 ( .A(n29288), .B(n29287), .Z(n29289) );
  XOR U30512 ( .A(n29241), .B(n29240), .Z(n29200) );
  XNOR U30513 ( .A(n29201), .B(n29200), .Z(n29296) );
  NAND U30514 ( .A(x[486]), .B(y[7982]), .Z(n29221) );
  NANDN U30515 ( .A(n29221), .B(n29129), .Z(n29132) );
  NAND U30516 ( .A(n29130), .B(n29264), .Z(n29131) );
  NAND U30517 ( .A(n29132), .B(n29131), .Z(n29229) );
  NAND U30518 ( .A(n29134), .B(n29133), .Z(n29138) );
  NAND U30519 ( .A(n29136), .B(n29135), .Z(n29137) );
  NAND U30520 ( .A(n29138), .B(n29137), .Z(n29227) );
  AND U30521 ( .A(y[7970]), .B(x[498]), .Z(n29140) );
  NAND U30522 ( .A(y[7976]), .B(x[492]), .Z(n29139) );
  XNOR U30523 ( .A(n29140), .B(n29139), .Z(n29205) );
  AND U30524 ( .A(x[497]), .B(y[7971]), .Z(n29206) );
  XOR U30525 ( .A(n29205), .B(n29206), .Z(n29226) );
  XOR U30526 ( .A(n29227), .B(n29226), .Z(n29228) );
  XNOR U30527 ( .A(n29229), .B(n29228), .Z(n29233) );
  AND U30528 ( .A(y[7975]), .B(x[493]), .Z(n29142) );
  NAND U30529 ( .A(y[7985]), .B(x[483]), .Z(n29141) );
  XNOR U30530 ( .A(n29142), .B(n29141), .Z(n29251) );
  XNOR U30531 ( .A(n29251), .B(n29250), .Z(n29223) );
  AND U30532 ( .A(y[7983]), .B(x[485]), .Z(n29144) );
  NAND U30533 ( .A(y[7984]), .B(x[484]), .Z(n29143) );
  XNOR U30534 ( .A(n29144), .B(n29143), .Z(n29266) );
  AND U30535 ( .A(x[487]), .B(y[7981]), .Z(n29265) );
  XNOR U30536 ( .A(n29266), .B(n29265), .Z(n29220) );
  XOR U30537 ( .A(n29221), .B(n29220), .Z(n29222) );
  XNOR U30538 ( .A(n29223), .B(n29222), .Z(n29277) );
  AND U30539 ( .A(x[488]), .B(y[7986]), .Z(n30383) );
  AND U30540 ( .A(x[481]), .B(y[7979]), .Z(n29145) );
  NAND U30541 ( .A(n30383), .B(n29145), .Z(n29149) );
  NANDN U30542 ( .A(n29147), .B(n29146), .Z(n29148) );
  AND U30543 ( .A(n29149), .B(n29148), .Z(n29276) );
  NAND U30544 ( .A(x[497]), .B(y[7977]), .Z(n30054) );
  NANDN U30545 ( .A(n30054), .B(n29150), .Z(n29154) );
  NAND U30546 ( .A(n29152), .B(n29151), .Z(n29153) );
  NAND U30547 ( .A(n29154), .B(n29153), .Z(n29275) );
  XNOR U30548 ( .A(n29277), .B(n29278), .Z(n29232) );
  XOR U30549 ( .A(n29233), .B(n29232), .Z(n29234) );
  NAND U30550 ( .A(n29156), .B(n29155), .Z(n29160) );
  NAND U30551 ( .A(n29158), .B(n29157), .Z(n29159) );
  AND U30552 ( .A(n29160), .B(n29159), .Z(n29235) );
  XOR U30553 ( .A(n29234), .B(n29235), .Z(n29293) );
  NAND U30554 ( .A(n29162), .B(n29161), .Z(n29166) );
  NAND U30555 ( .A(n29164), .B(n29163), .Z(n29165) );
  AND U30556 ( .A(n29166), .B(n29165), .Z(n29294) );
  XOR U30557 ( .A(n29293), .B(n29294), .Z(n29295) );
  XNOR U30558 ( .A(n29296), .B(n29295), .Z(n29300) );
  NANDN U30559 ( .A(n29168), .B(n29167), .Z(n29172) );
  NANDN U30560 ( .A(n29170), .B(n29169), .Z(n29171) );
  AND U30561 ( .A(n29172), .B(n29171), .Z(n29308) );
  NAND U30562 ( .A(n29174), .B(n29173), .Z(n29178) );
  NANDN U30563 ( .A(n29176), .B(n29175), .Z(n29177) );
  AND U30564 ( .A(n29178), .B(n29177), .Z(n29306) );
  NANDN U30565 ( .A(n29180), .B(n29179), .Z(n29184) );
  OR U30566 ( .A(n29182), .B(n29181), .Z(n29183) );
  AND U30567 ( .A(n29184), .B(n29183), .Z(n29305) );
  XNOR U30568 ( .A(n29306), .B(n29305), .Z(n29307) );
  XNOR U30569 ( .A(n29308), .B(n29307), .Z(n29299) );
  XNOR U30570 ( .A(n29300), .B(n29299), .Z(n29302) );
  XNOR U30571 ( .A(n29301), .B(n29302), .Z(n29317) );
  NAND U30572 ( .A(n29186), .B(n29185), .Z(n29190) );
  NANDN U30573 ( .A(n29188), .B(n29187), .Z(n29189) );
  AND U30574 ( .A(n29190), .B(n29189), .Z(n29315) );
  NANDN U30575 ( .A(n29192), .B(n29191), .Z(n29196) );
  NAND U30576 ( .A(n29194), .B(n29193), .Z(n29195) );
  AND U30577 ( .A(n29196), .B(n29195), .Z(n29314) );
  XOR U30578 ( .A(n29315), .B(n29314), .Z(n29316) );
  XOR U30579 ( .A(n29311), .B(n29313), .Z(n29197) );
  XNOR U30580 ( .A(n29312), .B(n29197), .Z(N629) );
  NAND U30581 ( .A(n29199), .B(n29198), .Z(n29203) );
  NAND U30582 ( .A(n29201), .B(n29200), .Z(n29202) );
  NAND U30583 ( .A(n29203), .B(n29202), .Z(n29330) );
  AND U30584 ( .A(x[498]), .B(y[7976]), .Z(n30053) );
  NAND U30585 ( .A(n30053), .B(n29204), .Z(n29208) );
  NAND U30586 ( .A(n29206), .B(n29205), .Z(n29207) );
  NAND U30587 ( .A(n29208), .B(n29207), .Z(n29407) );
  AND U30588 ( .A(x[491]), .B(y[7987]), .Z(n30738) );
  AND U30589 ( .A(x[481]), .B(y[7977]), .Z(n29209) );
  NAND U30590 ( .A(n30738), .B(n29209), .Z(n29213) );
  NAND U30591 ( .A(n29211), .B(n29210), .Z(n29212) );
  NAND U30592 ( .A(n29213), .B(n29212), .Z(n29406) );
  XOR U30593 ( .A(n29407), .B(n29406), .Z(n29409) );
  AND U30594 ( .A(x[495]), .B(y[7979]), .Z(n30041) );
  NAND U30595 ( .A(n30041), .B(n29214), .Z(n29218) );
  NAND U30596 ( .A(n29216), .B(n29215), .Z(n29217) );
  NAND U30597 ( .A(n29218), .B(n29217), .Z(n29365) );
  AND U30598 ( .A(x[480]), .B(y[7989]), .Z(n29384) );
  AND U30599 ( .A(x[501]), .B(y[7968]), .Z(n29385) );
  XOR U30600 ( .A(n29384), .B(n29385), .Z(n29387) );
  AND U30601 ( .A(o[308]), .B(n29219), .Z(n29386) );
  XOR U30602 ( .A(n29387), .B(n29386), .Z(n29363) );
  AND U30603 ( .A(x[485]), .B(y[7984]), .Z(n29371) );
  AND U30604 ( .A(x[496]), .B(y[7973]), .Z(n29370) );
  XOR U30605 ( .A(n29371), .B(n29370), .Z(n29369) );
  AND U30606 ( .A(x[495]), .B(y[7974]), .Z(n29368) );
  XOR U30607 ( .A(n29369), .B(n29368), .Z(n29362) );
  XOR U30608 ( .A(n29363), .B(n29362), .Z(n29364) );
  XOR U30609 ( .A(n29365), .B(n29364), .Z(n29408) );
  XOR U30610 ( .A(n29409), .B(n29408), .Z(n29401) );
  NAND U30611 ( .A(n29221), .B(n29220), .Z(n29225) );
  NAND U30612 ( .A(n29223), .B(n29222), .Z(n29224) );
  NAND U30613 ( .A(n29225), .B(n29224), .Z(n29400) );
  NAND U30614 ( .A(n29227), .B(n29226), .Z(n29231) );
  NAND U30615 ( .A(n29229), .B(n29228), .Z(n29230) );
  AND U30616 ( .A(n29231), .B(n29230), .Z(n29402) );
  XNOR U30617 ( .A(n29403), .B(n29402), .Z(n29328) );
  NAND U30618 ( .A(n29233), .B(n29232), .Z(n29237) );
  NAND U30619 ( .A(n29235), .B(n29234), .Z(n29236) );
  AND U30620 ( .A(n29237), .B(n29236), .Z(n29327) );
  XOR U30621 ( .A(n29328), .B(n29327), .Z(n29329) );
  XNOR U30622 ( .A(n29330), .B(n29329), .Z(n29323) );
  NANDN U30623 ( .A(n29239), .B(n29238), .Z(n29243) );
  NAND U30624 ( .A(n29241), .B(n29240), .Z(n29242) );
  NAND U30625 ( .A(n29243), .B(n29242), .Z(n29427) );
  NAND U30626 ( .A(n30046), .B(n29244), .Z(n29248) );
  NAND U30627 ( .A(n29246), .B(n29245), .Z(n29247) );
  NAND U30628 ( .A(n29248), .B(n29247), .Z(n29334) );
  NAND U30629 ( .A(n30673), .B(n29249), .Z(n29253) );
  NAND U30630 ( .A(n29251), .B(n29250), .Z(n29252) );
  NAND U30631 ( .A(n29253), .B(n29252), .Z(n29421) );
  AND U30632 ( .A(y[7970]), .B(x[499]), .Z(n29255) );
  NAND U30633 ( .A(y[7978]), .B(x[491]), .Z(n29254) );
  XNOR U30634 ( .A(n29255), .B(n29254), .Z(n29353) );
  AND U30635 ( .A(x[500]), .B(y[7969]), .Z(n29383) );
  XOR U30636 ( .A(o[309]), .B(n29383), .Z(n29352) );
  XOR U30637 ( .A(n29353), .B(n29352), .Z(n29419) );
  AND U30638 ( .A(y[7971]), .B(x[498]), .Z(n29257) );
  NAND U30639 ( .A(y[7979]), .B(x[490]), .Z(n29256) );
  XNOR U30640 ( .A(n29257), .B(n29256), .Z(n29391) );
  AND U30641 ( .A(x[481]), .B(y[7988]), .Z(n29392) );
  XOR U30642 ( .A(n29391), .B(n29392), .Z(n29418) );
  XOR U30643 ( .A(n29419), .B(n29418), .Z(n29420) );
  XOR U30644 ( .A(n29421), .B(n29420), .Z(n29333) );
  XOR U30645 ( .A(n29334), .B(n29333), .Z(n29336) );
  AND U30646 ( .A(x[487]), .B(y[7982]), .Z(n29600) );
  AND U30647 ( .A(y[7983]), .B(x[486]), .Z(n29259) );
  NAND U30648 ( .A(y[7975]), .B(x[494]), .Z(n29258) );
  XNOR U30649 ( .A(n29259), .B(n29258), .Z(n29395) );
  XNOR U30650 ( .A(n29600), .B(n29395), .Z(n29342) );
  NAND U30651 ( .A(x[489]), .B(y[7980]), .Z(n29340) );
  NAND U30652 ( .A(x[488]), .B(y[7981]), .Z(n29339) );
  XOR U30653 ( .A(n29340), .B(n29339), .Z(n29341) );
  XNOR U30654 ( .A(n29342), .B(n29341), .Z(n29358) );
  AND U30655 ( .A(y[7977]), .B(x[492]), .Z(n29261) );
  NAND U30656 ( .A(y[7972]), .B(x[497]), .Z(n29260) );
  XNOR U30657 ( .A(n29261), .B(n29260), .Z(n29345) );
  AND U30658 ( .A(x[482]), .B(y[7987]), .Z(n29346) );
  XOR U30659 ( .A(n29345), .B(n29346), .Z(n29357) );
  AND U30660 ( .A(y[7976]), .B(x[493]), .Z(n29263) );
  NAND U30661 ( .A(y[7986]), .B(x[483]), .Z(n29262) );
  XNOR U30662 ( .A(n29263), .B(n29262), .Z(n29379) );
  AND U30663 ( .A(x[484]), .B(y[7985]), .Z(n29380) );
  XOR U30664 ( .A(n29379), .B(n29380), .Z(n29356) );
  XOR U30665 ( .A(n29357), .B(n29356), .Z(n29359) );
  XOR U30666 ( .A(n29358), .B(n29359), .Z(n29415) );
  NAND U30667 ( .A(n29371), .B(n29264), .Z(n29268) );
  NAND U30668 ( .A(n29266), .B(n29265), .Z(n29267) );
  NAND U30669 ( .A(n29268), .B(n29267), .Z(n29413) );
  NAND U30670 ( .A(n29270), .B(n29269), .Z(n29274) );
  NAND U30671 ( .A(n29272), .B(n29271), .Z(n29273) );
  NAND U30672 ( .A(n29274), .B(n29273), .Z(n29412) );
  XOR U30673 ( .A(n29413), .B(n29412), .Z(n29414) );
  XOR U30674 ( .A(n29415), .B(n29414), .Z(n29335) );
  XOR U30675 ( .A(n29336), .B(n29335), .Z(n29425) );
  NANDN U30676 ( .A(n29276), .B(n29275), .Z(n29280) );
  NAND U30677 ( .A(n29278), .B(n29277), .Z(n29279) );
  NAND U30678 ( .A(n29280), .B(n29279), .Z(n29432) );
  NAND U30679 ( .A(n29282), .B(n29281), .Z(n29286) );
  NANDN U30680 ( .A(n29284), .B(n29283), .Z(n29285) );
  NAND U30681 ( .A(n29286), .B(n29285), .Z(n29431) );
  NAND U30682 ( .A(n29288), .B(n29287), .Z(n29292) );
  NANDN U30683 ( .A(n29290), .B(n29289), .Z(n29291) );
  NAND U30684 ( .A(n29292), .B(n29291), .Z(n29430) );
  XOR U30685 ( .A(n29431), .B(n29430), .Z(n29433) );
  XOR U30686 ( .A(n29432), .B(n29433), .Z(n29424) );
  XOR U30687 ( .A(n29425), .B(n29424), .Z(n29426) );
  XNOR U30688 ( .A(n29427), .B(n29426), .Z(n29322) );
  NAND U30689 ( .A(n29294), .B(n29293), .Z(n29298) );
  NAND U30690 ( .A(n29296), .B(n29295), .Z(n29297) );
  NAND U30691 ( .A(n29298), .B(n29297), .Z(n29321) );
  XOR U30692 ( .A(n29322), .B(n29321), .Z(n29324) );
  XNOR U30693 ( .A(n29323), .B(n29324), .Z(n29445) );
  NAND U30694 ( .A(n29300), .B(n29299), .Z(n29304) );
  NANDN U30695 ( .A(n29302), .B(n29301), .Z(n29303) );
  AND U30696 ( .A(n29304), .B(n29303), .Z(n29444) );
  NANDN U30697 ( .A(n29306), .B(n29305), .Z(n29310) );
  NAND U30698 ( .A(n29308), .B(n29307), .Z(n29309) );
  AND U30699 ( .A(n29310), .B(n29309), .Z(n29443) );
  XOR U30700 ( .A(n29444), .B(n29443), .Z(n29446) );
  XOR U30701 ( .A(n29445), .B(n29446), .Z(n29439) );
  NAND U30702 ( .A(n29315), .B(n29314), .Z(n29319) );
  NANDN U30703 ( .A(n29317), .B(n29316), .Z(n29318) );
  AND U30704 ( .A(n29319), .B(n29318), .Z(n29437) );
  IV U30705 ( .A(n29437), .Z(n29436) );
  XOR U30706 ( .A(n29438), .B(n29436), .Z(n29320) );
  XNOR U30707 ( .A(n29439), .B(n29320), .Z(N630) );
  NAND U30708 ( .A(n29322), .B(n29321), .Z(n29326) );
  NAND U30709 ( .A(n29324), .B(n29323), .Z(n29325) );
  AND U30710 ( .A(n29326), .B(n29325), .Z(n29576) );
  NAND U30711 ( .A(n29328), .B(n29327), .Z(n29332) );
  NAND U30712 ( .A(n29330), .B(n29329), .Z(n29331) );
  NAND U30713 ( .A(n29332), .B(n29331), .Z(n29574) );
  NAND U30714 ( .A(n29334), .B(n29333), .Z(n29338) );
  NAND U30715 ( .A(n29336), .B(n29335), .Z(n29337) );
  NAND U30716 ( .A(n29338), .B(n29337), .Z(n29567) );
  NAND U30717 ( .A(n29340), .B(n29339), .Z(n29344) );
  NAND U30718 ( .A(n29342), .B(n29341), .Z(n29343) );
  NAND U30719 ( .A(n29344), .B(n29343), .Z(n29561) );
  NANDN U30720 ( .A(n30054), .B(n29518), .Z(n29348) );
  NAND U30721 ( .A(n29346), .B(n29345), .Z(n29347) );
  NAND U30722 ( .A(n29348), .B(n29347), .Z(n29488) );
  AND U30723 ( .A(x[485]), .B(y[7985]), .Z(n29534) );
  AND U30724 ( .A(x[497]), .B(y[7973]), .Z(n29535) );
  XOR U30725 ( .A(n29534), .B(n29535), .Z(n29536) );
  AND U30726 ( .A(x[496]), .B(y[7974]), .Z(n29537) );
  XOR U30727 ( .A(n29536), .B(n29537), .Z(n29487) );
  AND U30728 ( .A(y[7972]), .B(x[498]), .Z(n29350) );
  NAND U30729 ( .A(y[7978]), .B(x[492]), .Z(n29349) );
  XNOR U30730 ( .A(n29350), .B(n29349), .Z(n29519) );
  AND U30731 ( .A(x[484]), .B(y[7986]), .Z(n29520) );
  XOR U30732 ( .A(n29519), .B(n29520), .Z(n29486) );
  XOR U30733 ( .A(n29487), .B(n29486), .Z(n29489) );
  XNOR U30734 ( .A(n29488), .B(n29489), .Z(n29558) );
  AND U30735 ( .A(x[499]), .B(y[7978]), .Z(n30563) );
  NAND U30736 ( .A(n30563), .B(n29351), .Z(n29355) );
  NAND U30737 ( .A(n29353), .B(n29352), .Z(n29354) );
  AND U30738 ( .A(n29355), .B(n29354), .Z(n29559) );
  XOR U30739 ( .A(n29558), .B(n29559), .Z(n29560) );
  XNOR U30740 ( .A(n29561), .B(n29560), .Z(n29564) );
  NAND U30741 ( .A(n29357), .B(n29356), .Z(n29361) );
  NAND U30742 ( .A(n29359), .B(n29358), .Z(n29360) );
  NAND U30743 ( .A(n29361), .B(n29360), .Z(n29547) );
  NAND U30744 ( .A(n29363), .B(n29362), .Z(n29367) );
  NAND U30745 ( .A(n29365), .B(n29364), .Z(n29366) );
  NAND U30746 ( .A(n29367), .B(n29366), .Z(n29546) );
  XOR U30747 ( .A(n29547), .B(n29546), .Z(n29549) );
  AND U30748 ( .A(n29369), .B(n29368), .Z(n29373) );
  NAND U30749 ( .A(n29371), .B(n29370), .Z(n29372) );
  NANDN U30750 ( .A(n29373), .B(n29372), .Z(n29509) );
  AND U30751 ( .A(y[7977]), .B(x[493]), .Z(n29375) );
  NAND U30752 ( .A(y[7970]), .B(x[500]), .Z(n29374) );
  XNOR U30753 ( .A(n29375), .B(n29374), .Z(n29530) );
  AND U30754 ( .A(x[482]), .B(y[7988]), .Z(n29531) );
  XOR U30755 ( .A(n29530), .B(n29531), .Z(n29507) );
  AND U30756 ( .A(y[7984]), .B(x[486]), .Z(n29377) );
  NAND U30757 ( .A(y[7975]), .B(x[495]), .Z(n29376) );
  XNOR U30758 ( .A(n29377), .B(n29376), .Z(n29542) );
  XOR U30759 ( .A(n29507), .B(n29506), .Z(n29508) );
  XOR U30760 ( .A(n29509), .B(n29508), .Z(n29553) );
  AND U30761 ( .A(x[493]), .B(y[7986]), .Z(n30813) );
  NAND U30762 ( .A(n29378), .B(n30813), .Z(n29382) );
  NAND U30763 ( .A(n29380), .B(n29379), .Z(n29381) );
  NAND U30764 ( .A(n29382), .B(n29381), .Z(n29477) );
  AND U30765 ( .A(x[481]), .B(y[7989]), .Z(n29500) );
  XOR U30766 ( .A(n29501), .B(n29500), .Z(n29499) );
  AND U30767 ( .A(o[309]), .B(n29383), .Z(n29498) );
  XOR U30768 ( .A(n29499), .B(n29498), .Z(n29475) );
  AND U30769 ( .A(x[494]), .B(y[7976]), .Z(n29492) );
  AND U30770 ( .A(x[483]), .B(y[7987]), .Z(n29493) );
  XOR U30771 ( .A(n29492), .B(n29493), .Z(n29494) );
  AND U30772 ( .A(x[499]), .B(y[7971]), .Z(n29495) );
  XOR U30773 ( .A(n29494), .B(n29495), .Z(n29474) );
  XOR U30774 ( .A(n29475), .B(n29474), .Z(n29476) );
  XOR U30775 ( .A(n29477), .B(n29476), .Z(n29552) );
  XOR U30776 ( .A(n29553), .B(n29552), .Z(n29555) );
  NAND U30777 ( .A(n29385), .B(n29384), .Z(n29389) );
  NAND U30778 ( .A(n29387), .B(n29386), .Z(n29388) );
  NAND U30779 ( .A(n29389), .B(n29388), .Z(n29469) );
  AND U30780 ( .A(x[498]), .B(y[7979]), .Z(n30566) );
  NAND U30781 ( .A(n30566), .B(n29390), .Z(n29394) );
  NAND U30782 ( .A(n29392), .B(n29391), .Z(n29393) );
  NAND U30783 ( .A(n29394), .B(n29393), .Z(n29468) );
  XOR U30784 ( .A(n29469), .B(n29468), .Z(n29471) );
  AND U30785 ( .A(x[494]), .B(y[7983]), .Z(n30582) );
  NAND U30786 ( .A(n30582), .B(n29541), .Z(n29397) );
  NAND U30787 ( .A(n29600), .B(n29395), .Z(n29396) );
  NAND U30788 ( .A(n29397), .B(n29396), .Z(n29483) );
  AND U30789 ( .A(x[480]), .B(y[7990]), .Z(n29523) );
  AND U30790 ( .A(x[502]), .B(y[7968]), .Z(n29524) );
  XOR U30791 ( .A(n29523), .B(n29524), .Z(n29526) );
  AND U30792 ( .A(x[501]), .B(y[7969]), .Z(n29540) );
  XOR U30793 ( .A(o[310]), .B(n29540), .Z(n29525) );
  XOR U30794 ( .A(n29526), .B(n29525), .Z(n29481) );
  AND U30795 ( .A(y[7983]), .B(x[487]), .Z(n29399) );
  NAND U30796 ( .A(y[7982]), .B(x[488]), .Z(n29398) );
  XNOR U30797 ( .A(n29399), .B(n29398), .Z(n29512) );
  XOR U30798 ( .A(n29481), .B(n29480), .Z(n29482) );
  XOR U30799 ( .A(n29483), .B(n29482), .Z(n29470) );
  XOR U30800 ( .A(n29471), .B(n29470), .Z(n29554) );
  XOR U30801 ( .A(n29555), .B(n29554), .Z(n29548) );
  XOR U30802 ( .A(n29549), .B(n29548), .Z(n29565) );
  XOR U30803 ( .A(n29564), .B(n29565), .Z(n29566) );
  XNOR U30804 ( .A(n29567), .B(n29566), .Z(n29458) );
  NANDN U30805 ( .A(n29401), .B(n29400), .Z(n29405) );
  NAND U30806 ( .A(n29403), .B(n29402), .Z(n29404) );
  AND U30807 ( .A(n29405), .B(n29404), .Z(n29457) );
  NAND U30808 ( .A(n29407), .B(n29406), .Z(n29411) );
  NAND U30809 ( .A(n29409), .B(n29408), .Z(n29410) );
  AND U30810 ( .A(n29411), .B(n29410), .Z(n29465) );
  NAND U30811 ( .A(n29413), .B(n29412), .Z(n29417) );
  NAND U30812 ( .A(n29415), .B(n29414), .Z(n29416) );
  NAND U30813 ( .A(n29417), .B(n29416), .Z(n29463) );
  NAND U30814 ( .A(n29419), .B(n29418), .Z(n29423) );
  NAND U30815 ( .A(n29421), .B(n29420), .Z(n29422) );
  NAND U30816 ( .A(n29423), .B(n29422), .Z(n29462) );
  XOR U30817 ( .A(n29463), .B(n29462), .Z(n29464) );
  XOR U30818 ( .A(n29465), .B(n29464), .Z(n29456) );
  XNOR U30819 ( .A(n29458), .B(n29459), .Z(n29452) );
  NAND U30820 ( .A(n29425), .B(n29424), .Z(n29429) );
  NAND U30821 ( .A(n29427), .B(n29426), .Z(n29428) );
  AND U30822 ( .A(n29429), .B(n29428), .Z(n29451) );
  NAND U30823 ( .A(n29431), .B(n29430), .Z(n29435) );
  NAND U30824 ( .A(n29433), .B(n29432), .Z(n29434) );
  NAND U30825 ( .A(n29435), .B(n29434), .Z(n29450) );
  XOR U30826 ( .A(n29452), .B(n29453), .Z(n29573) );
  XOR U30827 ( .A(n29574), .B(n29573), .Z(n29575) );
  XNOR U30828 ( .A(n29576), .B(n29575), .Z(n29570) );
  OR U30829 ( .A(n29438), .B(n29436), .Z(n29442) );
  ANDN U30830 ( .B(n29438), .A(n29437), .Z(n29440) );
  OR U30831 ( .A(n29440), .B(n29439), .Z(n29441) );
  AND U30832 ( .A(n29442), .B(n29441), .Z(n29571) );
  NANDN U30833 ( .A(n29444), .B(n29443), .Z(n29448) );
  NANDN U30834 ( .A(n29446), .B(n29445), .Z(n29447) );
  AND U30835 ( .A(n29448), .B(n29447), .Z(n29572) );
  XOR U30836 ( .A(n29571), .B(n29572), .Z(n29449) );
  XNOR U30837 ( .A(n29570), .B(n29449), .Z(N631) );
  NANDN U30838 ( .A(n29451), .B(n29450), .Z(n29455) );
  NAND U30839 ( .A(n29453), .B(n29452), .Z(n29454) );
  AND U30840 ( .A(n29455), .B(n29454), .Z(n29714) );
  NANDN U30841 ( .A(n29457), .B(n29456), .Z(n29461) );
  NAND U30842 ( .A(n29459), .B(n29458), .Z(n29460) );
  AND U30843 ( .A(n29461), .B(n29460), .Z(n29712) );
  NAND U30844 ( .A(n29463), .B(n29462), .Z(n29467) );
  NANDN U30845 ( .A(n29465), .B(n29464), .Z(n29466) );
  NAND U30846 ( .A(n29467), .B(n29466), .Z(n29696) );
  NAND U30847 ( .A(n29469), .B(n29468), .Z(n29473) );
  NAND U30848 ( .A(n29471), .B(n29470), .Z(n29472) );
  NAND U30849 ( .A(n29473), .B(n29472), .Z(n29690) );
  NAND U30850 ( .A(n29475), .B(n29474), .Z(n29479) );
  NAND U30851 ( .A(n29477), .B(n29476), .Z(n29478) );
  NAND U30852 ( .A(n29479), .B(n29478), .Z(n29688) );
  NAND U30853 ( .A(n29481), .B(n29480), .Z(n29485) );
  NAND U30854 ( .A(n29483), .B(n29482), .Z(n29484) );
  NAND U30855 ( .A(n29485), .B(n29484), .Z(n29687) );
  XOR U30856 ( .A(n29688), .B(n29687), .Z(n29689) );
  XOR U30857 ( .A(n29690), .B(n29689), .Z(n29708) );
  NAND U30858 ( .A(n29487), .B(n29486), .Z(n29491) );
  NAND U30859 ( .A(n29489), .B(n29488), .Z(n29490) );
  NAND U30860 ( .A(n29491), .B(n29490), .Z(n29706) );
  NAND U30861 ( .A(n29493), .B(n29492), .Z(n29497) );
  NAND U30862 ( .A(n29495), .B(n29494), .Z(n29496) );
  NAND U30863 ( .A(n29497), .B(n29496), .Z(n29634) );
  AND U30864 ( .A(n29499), .B(n29498), .Z(n29503) );
  NAND U30865 ( .A(n29501), .B(n29500), .Z(n29502) );
  NANDN U30866 ( .A(n29503), .B(n29502), .Z(n29633) );
  XOR U30867 ( .A(n29634), .B(n29633), .Z(n29636) );
  AND U30868 ( .A(y[7984]), .B(x[487]), .Z(n29505) );
  NAND U30869 ( .A(y[7982]), .B(x[489]), .Z(n29504) );
  XNOR U30870 ( .A(n29505), .B(n29504), .Z(n29602) );
  XOR U30871 ( .A(n29601), .B(n29602), .Z(n29639) );
  AND U30872 ( .A(x[490]), .B(y[7981]), .Z(n29640) );
  XOR U30873 ( .A(n29639), .B(n29640), .Z(n29642) );
  AND U30874 ( .A(x[486]), .B(y[7985]), .Z(n29592) );
  AND U30875 ( .A(x[495]), .B(y[7976]), .Z(n29593) );
  XOR U30876 ( .A(n29592), .B(n29593), .Z(n29594) );
  AND U30877 ( .A(x[491]), .B(y[7980]), .Z(n29595) );
  XOR U30878 ( .A(n29594), .B(n29595), .Z(n29641) );
  XOR U30879 ( .A(n29642), .B(n29641), .Z(n29635) );
  XOR U30880 ( .A(n29636), .B(n29635), .Z(n29705) );
  XOR U30881 ( .A(n29706), .B(n29705), .Z(n29707) );
  XOR U30882 ( .A(n29708), .B(n29707), .Z(n29694) );
  NAND U30883 ( .A(n29507), .B(n29506), .Z(n29511) );
  NAND U30884 ( .A(n29509), .B(n29508), .Z(n29510) );
  NAND U30885 ( .A(n29511), .B(n29510), .Z(n29628) );
  NAND U30886 ( .A(n29600), .B(n29601), .Z(n29515) );
  NANDN U30887 ( .A(n29513), .B(n29512), .Z(n29514) );
  AND U30888 ( .A(n29515), .B(n29514), .Z(n29678) );
  AND U30889 ( .A(x[480]), .B(y[7991]), .Z(n29611) );
  AND U30890 ( .A(x[503]), .B(y[7968]), .Z(n29612) );
  XOR U30891 ( .A(n29611), .B(n29612), .Z(n29614) );
  AND U30892 ( .A(x[502]), .B(y[7969]), .Z(n29591) );
  XOR U30893 ( .A(o[311]), .B(n29591), .Z(n29613) );
  XOR U30894 ( .A(n29614), .B(n29613), .Z(n29676) );
  NAND U30895 ( .A(y[7971]), .B(x[500]), .Z(n29516) );
  XNOR U30896 ( .A(n29517), .B(n29516), .Z(n29587) );
  AND U30897 ( .A(x[499]), .B(y[7972]), .Z(n29588) );
  XOR U30898 ( .A(n29587), .B(n29588), .Z(n29675) );
  XOR U30899 ( .A(n29676), .B(n29675), .Z(n29677) );
  NAND U30900 ( .A(x[498]), .B(y[7978]), .Z(n30414) );
  NANDN U30901 ( .A(n30414), .B(n29518), .Z(n29522) );
  NAND U30902 ( .A(n29520), .B(n29519), .Z(n29521) );
  AND U30903 ( .A(n29522), .B(n29521), .Z(n29664) );
  NAND U30904 ( .A(n29524), .B(n29523), .Z(n29528) );
  NAND U30905 ( .A(n29526), .B(n29525), .Z(n29527) );
  NAND U30906 ( .A(n29528), .B(n29527), .Z(n29663) );
  XOR U30907 ( .A(n29666), .B(n29665), .Z(n29627) );
  XOR U30908 ( .A(n29628), .B(n29627), .Z(n29630) );
  NAND U30909 ( .A(x[500]), .B(y[7977]), .Z(n30594) );
  AND U30910 ( .A(x[493]), .B(y[7970]), .Z(n29529) );
  NANDN U30911 ( .A(n30594), .B(n29529), .Z(n29533) );
  NAND U30912 ( .A(n29531), .B(n29530), .Z(n29532) );
  NAND U30913 ( .A(n29533), .B(n29532), .Z(n29622) );
  NAND U30914 ( .A(n29535), .B(n29534), .Z(n29539) );
  NAND U30915 ( .A(n29537), .B(n29536), .Z(n29538) );
  AND U30916 ( .A(n29539), .B(n29538), .Z(n29684) );
  AND U30917 ( .A(x[493]), .B(y[7978]), .Z(n29657) );
  AND U30918 ( .A(x[482]), .B(y[7989]), .Z(n29658) );
  XOR U30919 ( .A(n29657), .B(n29658), .Z(n29659) );
  AND U30920 ( .A(x[501]), .B(y[7970]), .Z(n29660) );
  XOR U30921 ( .A(n29659), .B(n29660), .Z(n29682) );
  AND U30922 ( .A(x[492]), .B(y[7979]), .Z(n29605) );
  AND U30923 ( .A(x[481]), .B(y[7990]), .Z(n29606) );
  XOR U30924 ( .A(n29605), .B(n29606), .Z(n29608) );
  AND U30925 ( .A(o[310]), .B(n29540), .Z(n29607) );
  XOR U30926 ( .A(n29608), .B(n29607), .Z(n29681) );
  XOR U30927 ( .A(n29682), .B(n29681), .Z(n29683) );
  XOR U30928 ( .A(n29622), .B(n29621), .Z(n29624) );
  AND U30929 ( .A(x[495]), .B(y[7984]), .Z(n30807) );
  NAND U30930 ( .A(n30807), .B(n29541), .Z(n29545) );
  NANDN U30931 ( .A(n29543), .B(n29542), .Z(n29544) );
  AND U30932 ( .A(n29545), .B(n29544), .Z(n29672) );
  AND U30933 ( .A(x[494]), .B(y[7977]), .Z(n29651) );
  AND U30934 ( .A(x[483]), .B(y[7988]), .Z(n29652) );
  XOR U30935 ( .A(n29651), .B(n29652), .Z(n29653) );
  AND U30936 ( .A(x[484]), .B(y[7987]), .Z(n29654) );
  XOR U30937 ( .A(n29653), .B(n29654), .Z(n29670) );
  AND U30938 ( .A(x[485]), .B(y[7986]), .Z(n29645) );
  AND U30939 ( .A(x[498]), .B(y[7973]), .Z(n29646) );
  XOR U30940 ( .A(n29645), .B(n29646), .Z(n29647) );
  AND U30941 ( .A(x[497]), .B(y[7974]), .Z(n29648) );
  XOR U30942 ( .A(n29647), .B(n29648), .Z(n29669) );
  XOR U30943 ( .A(n29670), .B(n29669), .Z(n29671) );
  XOR U30944 ( .A(n29624), .B(n29623), .Z(n29629) );
  XOR U30945 ( .A(n29630), .B(n29629), .Z(n29693) );
  XOR U30946 ( .A(n29694), .B(n29693), .Z(n29695) );
  XNOR U30947 ( .A(n29696), .B(n29695), .Z(n29582) );
  NAND U30948 ( .A(n29547), .B(n29546), .Z(n29551) );
  NAND U30949 ( .A(n29549), .B(n29548), .Z(n29550) );
  NAND U30950 ( .A(n29551), .B(n29550), .Z(n29702) );
  NAND U30951 ( .A(n29553), .B(n29552), .Z(n29557) );
  NAND U30952 ( .A(n29555), .B(n29554), .Z(n29556) );
  NAND U30953 ( .A(n29557), .B(n29556), .Z(n29700) );
  NAND U30954 ( .A(n29559), .B(n29558), .Z(n29563) );
  NAND U30955 ( .A(n29561), .B(n29560), .Z(n29562) );
  AND U30956 ( .A(n29563), .B(n29562), .Z(n29699) );
  XOR U30957 ( .A(n29700), .B(n29699), .Z(n29701) );
  XNOR U30958 ( .A(n29702), .B(n29701), .Z(n29580) );
  NAND U30959 ( .A(n29565), .B(n29564), .Z(n29569) );
  NAND U30960 ( .A(n29567), .B(n29566), .Z(n29568) );
  AND U30961 ( .A(n29569), .B(n29568), .Z(n29581) );
  XOR U30962 ( .A(n29580), .B(n29581), .Z(n29583) );
  XOR U30963 ( .A(n29582), .B(n29583), .Z(n29711) );
  XNOR U30964 ( .A(n29714), .B(n29713), .Z(n29720) );
  NAND U30965 ( .A(n29574), .B(n29573), .Z(n29578) );
  NAND U30966 ( .A(n29576), .B(n29575), .Z(n29577) );
  AND U30967 ( .A(n29578), .B(n29577), .Z(n29719) );
  IV U30968 ( .A(n29719), .Z(n29717) );
  XOR U30969 ( .A(n29718), .B(n29717), .Z(n29579) );
  XNOR U30970 ( .A(n29720), .B(n29579), .Z(N632) );
  NAND U30971 ( .A(n29581), .B(n29580), .Z(n29585) );
  NAND U30972 ( .A(n29583), .B(n29582), .Z(n29584) );
  AND U30973 ( .A(n29585), .B(n29584), .Z(n29859) );
  AND U30974 ( .A(x[500]), .B(y[7975]), .Z(n29586) );
  NAND U30975 ( .A(n29586), .B(n29755), .Z(n29590) );
  NAND U30976 ( .A(n29588), .B(n29587), .Z(n29589) );
  NAND U30977 ( .A(n29590), .B(n29589), .Z(n29775) );
  AND U30978 ( .A(x[502]), .B(y[7970]), .Z(n29794) );
  XOR U30979 ( .A(n29795), .B(n29794), .Z(n29797) );
  AND U30980 ( .A(x[482]), .B(y[7990]), .Z(n29796) );
  XOR U30981 ( .A(n29797), .B(n29796), .Z(n29773) );
  AND U30982 ( .A(x[481]), .B(y[7991]), .Z(n29802) );
  XOR U30983 ( .A(n29803), .B(n29802), .Z(n29801) );
  AND U30984 ( .A(o[311]), .B(n29591), .Z(n29800) );
  XOR U30985 ( .A(n29801), .B(n29800), .Z(n29772) );
  XOR U30986 ( .A(n29773), .B(n29772), .Z(n29774) );
  XOR U30987 ( .A(n29775), .B(n29774), .Z(n29833) );
  NAND U30988 ( .A(n29593), .B(n29592), .Z(n29597) );
  NAND U30989 ( .A(n29595), .B(n29594), .Z(n29596) );
  NAND U30990 ( .A(n29597), .B(n29596), .Z(n29769) );
  AND U30991 ( .A(y[7976]), .B(x[496]), .Z(n29599) );
  NAND U30992 ( .A(y[7971]), .B(x[501]), .Z(n29598) );
  XNOR U30993 ( .A(n29599), .B(n29598), .Z(n29756) );
  AND U30994 ( .A(x[485]), .B(y[7987]), .Z(n29757) );
  XOR U30995 ( .A(n29756), .B(n29757), .Z(n29767) );
  AND U30996 ( .A(x[486]), .B(y[7986]), .Z(n30140) );
  NAND U30997 ( .A(x[500]), .B(y[7972]), .Z(n29986) );
  AND U30998 ( .A(x[499]), .B(y[7973]), .Z(n29763) );
  XOR U30999 ( .A(n29762), .B(n29763), .Z(n29766) );
  XOR U31000 ( .A(n29767), .B(n29766), .Z(n29768) );
  XOR U31001 ( .A(n29769), .B(n29768), .Z(n29746) );
  NAND U31002 ( .A(n29912), .B(n29600), .Z(n29604) );
  NAND U31003 ( .A(n29602), .B(n29601), .Z(n29603) );
  NAND U31004 ( .A(n29604), .B(n29603), .Z(n29744) );
  NAND U31005 ( .A(n29606), .B(n29605), .Z(n29610) );
  NAND U31006 ( .A(n29608), .B(n29607), .Z(n29609) );
  NAND U31007 ( .A(n29610), .B(n29609), .Z(n29743) );
  XOR U31008 ( .A(n29744), .B(n29743), .Z(n29745) );
  XOR U31009 ( .A(n29746), .B(n29745), .Z(n29832) );
  XOR U31010 ( .A(n29833), .B(n29832), .Z(n29835) );
  NAND U31011 ( .A(n29612), .B(n29611), .Z(n29616) );
  NAND U31012 ( .A(n29614), .B(n29613), .Z(n29615) );
  AND U31013 ( .A(n29616), .B(n29615), .Z(n29827) );
  AND U31014 ( .A(x[483]), .B(y[7989]), .Z(n29816) );
  XOR U31015 ( .A(n29817), .B(n29816), .Z(n29815) );
  AND U31016 ( .A(x[484]), .B(y[7988]), .Z(n29814) );
  XOR U31017 ( .A(n29815), .B(n29814), .Z(n29826) );
  AND U31018 ( .A(y[7983]), .B(x[489]), .Z(n29618) );
  NAND U31019 ( .A(y[7982]), .B(x[490]), .Z(n29617) );
  XNOR U31020 ( .A(n29618), .B(n29617), .Z(n29786) );
  AND U31021 ( .A(y[7978]), .B(x[494]), .Z(n29620) );
  NAND U31022 ( .A(y[7984]), .B(x[488]), .Z(n29619) );
  XNOR U31023 ( .A(n29620), .B(n29619), .Z(n29790) );
  NAND U31024 ( .A(x[491]), .B(y[7981]), .Z(n29791) );
  XOR U31025 ( .A(n29786), .B(n29785), .Z(n29828) );
  XOR U31026 ( .A(n29829), .B(n29828), .Z(n29834) );
  XNOR U31027 ( .A(n29835), .B(n29834), .Z(n29845) );
  NAND U31028 ( .A(n29622), .B(n29621), .Z(n29626) );
  NAND U31029 ( .A(n29624), .B(n29623), .Z(n29625) );
  AND U31030 ( .A(n29626), .B(n29625), .Z(n29844) );
  XOR U31031 ( .A(n29845), .B(n29844), .Z(n29846) );
  NAND U31032 ( .A(n29628), .B(n29627), .Z(n29632) );
  NAND U31033 ( .A(n29630), .B(n29629), .Z(n29631) );
  AND U31034 ( .A(n29632), .B(n29631), .Z(n29847) );
  XOR U31035 ( .A(n29846), .B(n29847), .Z(n29853) );
  NAND U31036 ( .A(n29634), .B(n29633), .Z(n29638) );
  NAND U31037 ( .A(n29636), .B(n29635), .Z(n29637) );
  NAND U31038 ( .A(n29638), .B(n29637), .Z(n29841) );
  NAND U31039 ( .A(n29640), .B(n29639), .Z(n29644) );
  NAND U31040 ( .A(n29642), .B(n29641), .Z(n29643) );
  NAND U31041 ( .A(n29644), .B(n29643), .Z(n29839) );
  NAND U31042 ( .A(n29646), .B(n29645), .Z(n29650) );
  NAND U31043 ( .A(n29648), .B(n29647), .Z(n29649) );
  NAND U31044 ( .A(n29650), .B(n29649), .Z(n29752) );
  AND U31045 ( .A(x[480]), .B(y[7992]), .Z(n29820) );
  NAND U31046 ( .A(x[504]), .B(y[7968]), .Z(n29821) );
  NAND U31047 ( .A(x[503]), .B(y[7969]), .Z(n29813) );
  XOR U31048 ( .A(o[312]), .B(n29813), .Z(n29823) );
  AND U31049 ( .A(x[487]), .B(y[7985]), .Z(n29806) );
  NAND U31050 ( .A(x[498]), .B(y[7974]), .Z(n29807) );
  NAND U31051 ( .A(x[497]), .B(y[7975]), .Z(n29809) );
  XOR U31052 ( .A(n29750), .B(n29749), .Z(n29751) );
  XOR U31053 ( .A(n29752), .B(n29751), .Z(n29740) );
  NAND U31054 ( .A(n29652), .B(n29651), .Z(n29656) );
  NAND U31055 ( .A(n29654), .B(n29653), .Z(n29655) );
  NAND U31056 ( .A(n29656), .B(n29655), .Z(n29738) );
  NAND U31057 ( .A(n29658), .B(n29657), .Z(n29662) );
  NAND U31058 ( .A(n29660), .B(n29659), .Z(n29661) );
  NAND U31059 ( .A(n29662), .B(n29661), .Z(n29737) );
  XOR U31060 ( .A(n29738), .B(n29737), .Z(n29739) );
  XOR U31061 ( .A(n29740), .B(n29739), .Z(n29838) );
  XOR U31062 ( .A(n29839), .B(n29838), .Z(n29840) );
  XNOR U31063 ( .A(n29841), .B(n29840), .Z(n29780) );
  NANDN U31064 ( .A(n29664), .B(n29663), .Z(n29668) );
  NAND U31065 ( .A(n29666), .B(n29665), .Z(n29667) );
  AND U31066 ( .A(n29668), .B(n29667), .Z(n29734) );
  NAND U31067 ( .A(n29670), .B(n29669), .Z(n29674) );
  NANDN U31068 ( .A(n29672), .B(n29671), .Z(n29673) );
  AND U31069 ( .A(n29674), .B(n29673), .Z(n29731) );
  NAND U31070 ( .A(n29676), .B(n29675), .Z(n29680) );
  NANDN U31071 ( .A(n29678), .B(n29677), .Z(n29679) );
  AND U31072 ( .A(n29680), .B(n29679), .Z(n29732) );
  XOR U31073 ( .A(n29731), .B(n29732), .Z(n29733) );
  XOR U31074 ( .A(n29734), .B(n29733), .Z(n29778) );
  NAND U31075 ( .A(n29682), .B(n29681), .Z(n29686) );
  NANDN U31076 ( .A(n29684), .B(n29683), .Z(n29685) );
  AND U31077 ( .A(n29686), .B(n29685), .Z(n29779) );
  XOR U31078 ( .A(n29778), .B(n29779), .Z(n29781) );
  XOR U31079 ( .A(n29780), .B(n29781), .Z(n29850) );
  NAND U31080 ( .A(n29688), .B(n29687), .Z(n29692) );
  NAND U31081 ( .A(n29690), .B(n29689), .Z(n29691) );
  AND U31082 ( .A(n29692), .B(n29691), .Z(n29851) );
  XOR U31083 ( .A(n29850), .B(n29851), .Z(n29852) );
  XNOR U31084 ( .A(n29853), .B(n29852), .Z(n29857) );
  NAND U31085 ( .A(n29694), .B(n29693), .Z(n29698) );
  NAND U31086 ( .A(n29696), .B(n29695), .Z(n29697) );
  NAND U31087 ( .A(n29698), .B(n29697), .Z(n29728) );
  NAND U31088 ( .A(n29700), .B(n29699), .Z(n29704) );
  NAND U31089 ( .A(n29702), .B(n29701), .Z(n29703) );
  NAND U31090 ( .A(n29704), .B(n29703), .Z(n29726) );
  NAND U31091 ( .A(n29706), .B(n29705), .Z(n29710) );
  NAND U31092 ( .A(n29708), .B(n29707), .Z(n29709) );
  NAND U31093 ( .A(n29710), .B(n29709), .Z(n29725) );
  XOR U31094 ( .A(n29726), .B(n29725), .Z(n29727) );
  XOR U31095 ( .A(n29728), .B(n29727), .Z(n29856) );
  XOR U31096 ( .A(n29857), .B(n29856), .Z(n29858) );
  XOR U31097 ( .A(n29859), .B(n29858), .Z(n29864) );
  NANDN U31098 ( .A(n29712), .B(n29711), .Z(n29716) );
  NAND U31099 ( .A(n29714), .B(n29713), .Z(n29715) );
  NAND U31100 ( .A(n29716), .B(n29715), .Z(n29862) );
  NANDN U31101 ( .A(n29717), .B(n29718), .Z(n29723) );
  NOR U31102 ( .A(n29719), .B(n29718), .Z(n29721) );
  OR U31103 ( .A(n29721), .B(n29720), .Z(n29722) );
  AND U31104 ( .A(n29723), .B(n29722), .Z(n29863) );
  XOR U31105 ( .A(n29862), .B(n29863), .Z(n29724) );
  XNOR U31106 ( .A(n29864), .B(n29724), .Z(N633) );
  NAND U31107 ( .A(n29726), .B(n29725), .Z(n29730) );
  NAND U31108 ( .A(n29728), .B(n29727), .Z(n29729) );
  AND U31109 ( .A(n29730), .B(n29729), .Z(n29869) );
  NAND U31110 ( .A(n29732), .B(n29731), .Z(n29736) );
  NAND U31111 ( .A(n29734), .B(n29733), .Z(n29735) );
  AND U31112 ( .A(n29736), .B(n29735), .Z(n29882) );
  NAND U31113 ( .A(n29738), .B(n29737), .Z(n29742) );
  NAND U31114 ( .A(n29740), .B(n29739), .Z(n29741) );
  NAND U31115 ( .A(n29742), .B(n29741), .Z(n29900) );
  NAND U31116 ( .A(n29744), .B(n29743), .Z(n29748) );
  NAND U31117 ( .A(n29746), .B(n29745), .Z(n29747) );
  NAND U31118 ( .A(n29748), .B(n29747), .Z(n29899) );
  XOR U31119 ( .A(n29900), .B(n29899), .Z(n29902) );
  NAND U31120 ( .A(n29750), .B(n29749), .Z(n29754) );
  NAND U31121 ( .A(n29752), .B(n29751), .Z(n29753) );
  AND U31122 ( .A(n29754), .B(n29753), .Z(n29932) );
  NAND U31123 ( .A(x[501]), .B(y[7976]), .Z(n30777) );
  NANDN U31124 ( .A(n30777), .B(n29755), .Z(n29759) );
  NAND U31125 ( .A(n29757), .B(n29756), .Z(n29758) );
  AND U31126 ( .A(n29759), .B(n29758), .Z(n30006) );
  AND U31127 ( .A(x[502]), .B(y[7971]), .Z(n29975) );
  AND U31128 ( .A(x[485]), .B(y[7988]), .Z(n29974) );
  NAND U31129 ( .A(x[497]), .B(y[7976]), .Z(n29973) );
  XOR U31130 ( .A(n29974), .B(n29973), .Z(n29976) );
  XOR U31131 ( .A(n29975), .B(n29976), .Z(n30004) );
  AND U31132 ( .A(y[7973]), .B(x[500]), .Z(n29761) );
  NAND U31133 ( .A(y[7972]), .B(x[501]), .Z(n29760) );
  XNOR U31134 ( .A(n29761), .B(n29760), .Z(n29988) );
  AND U31135 ( .A(x[499]), .B(y[7974]), .Z(n29987) );
  XOR U31136 ( .A(n29988), .B(n29987), .Z(n30003) );
  NANDN U31137 ( .A(n29986), .B(n30140), .Z(n29765) );
  NAND U31138 ( .A(n29763), .B(n29762), .Z(n29764) );
  AND U31139 ( .A(n29765), .B(n29764), .Z(n30012) );
  AND U31140 ( .A(x[495]), .B(y[7978]), .Z(n29993) );
  AND U31141 ( .A(x[498]), .B(y[7975]), .Z(n29992) );
  NAND U31142 ( .A(x[486]), .B(y[7987]), .Z(n29991) );
  XOR U31143 ( .A(n29992), .B(n29991), .Z(n29994) );
  XOR U31144 ( .A(n29993), .B(n29994), .Z(n30010) );
  AND U31145 ( .A(x[503]), .B(y[7970]), .Z(n29969) );
  AND U31146 ( .A(x[484]), .B(y[7989]), .Z(n29968) );
  NAND U31147 ( .A(x[496]), .B(y[7977]), .Z(n29967) );
  XOR U31148 ( .A(n29968), .B(n29967), .Z(n29970) );
  XNOR U31149 ( .A(n29969), .B(n29970), .Z(n30009) );
  XOR U31150 ( .A(n30012), .B(n30011), .Z(n29929) );
  XOR U31151 ( .A(n29930), .B(n29929), .Z(n29931) );
  XNOR U31152 ( .A(n29932), .B(n29931), .Z(n29944) );
  NAND U31153 ( .A(n29767), .B(n29766), .Z(n29771) );
  NAND U31154 ( .A(n29769), .B(n29768), .Z(n29770) );
  NAND U31155 ( .A(n29771), .B(n29770), .Z(n29942) );
  NAND U31156 ( .A(n29773), .B(n29772), .Z(n29777) );
  NAND U31157 ( .A(n29775), .B(n29774), .Z(n29776) );
  NAND U31158 ( .A(n29777), .B(n29776), .Z(n29941) );
  XOR U31159 ( .A(n29942), .B(n29941), .Z(n29943) );
  XOR U31160 ( .A(n29944), .B(n29943), .Z(n29901) );
  XNOR U31161 ( .A(n29902), .B(n29901), .Z(n29881) );
  NAND U31162 ( .A(n29779), .B(n29778), .Z(n29783) );
  NAND U31163 ( .A(n29781), .B(n29780), .Z(n29782) );
  NAND U31164 ( .A(n29783), .B(n29782), .Z(n29883) );
  XNOR U31165 ( .A(n29884), .B(n29883), .Z(n29878) );
  NANDN U31166 ( .A(n29911), .B(n29784), .Z(n29788) );
  NAND U31167 ( .A(n29786), .B(n29785), .Z(n29787) );
  NAND U31168 ( .A(n29788), .B(n29787), .Z(n29936) );
  AND U31169 ( .A(x[494]), .B(y[7984]), .Z(n30734) );
  NAND U31170 ( .A(n30734), .B(n29789), .Z(n29793) );
  NANDN U31171 ( .A(n29791), .B(n29790), .Z(n29792) );
  NAND U31172 ( .A(n29793), .B(n29792), .Z(n29963) );
  AND U31173 ( .A(x[491]), .B(y[7982]), .Z(n29983) );
  AND U31174 ( .A(x[492]), .B(y[7981]), .Z(n29981) );
  NAND U31175 ( .A(x[487]), .B(y[7986]), .Z(n29980) );
  XNOR U31176 ( .A(n29981), .B(n29980), .Z(n29982) );
  XOR U31177 ( .A(n29983), .B(n29982), .Z(n29961) );
  NAND U31178 ( .A(x[504]), .B(y[7969]), .Z(n29979) );
  XNOR U31179 ( .A(o[313]), .B(n29979), .Z(n29950) );
  AND U31180 ( .A(x[481]), .B(y[7992]), .Z(n29949) );
  XOR U31181 ( .A(n29950), .B(n29949), .Z(n29952) );
  AND U31182 ( .A(x[493]), .B(y[7980]), .Z(n29951) );
  XOR U31183 ( .A(n29952), .B(n29951), .Z(n29962) );
  XOR U31184 ( .A(n29961), .B(n29962), .Z(n29964) );
  XOR U31185 ( .A(n29963), .B(n29964), .Z(n29935) );
  XOR U31186 ( .A(n29936), .B(n29935), .Z(n29938) );
  NAND U31187 ( .A(n29795), .B(n29794), .Z(n29799) );
  AND U31188 ( .A(n29797), .B(n29796), .Z(n29798) );
  ANDN U31189 ( .B(n29799), .A(n29798), .Z(n29924) );
  AND U31190 ( .A(n29801), .B(n29800), .Z(n29805) );
  NAND U31191 ( .A(n29803), .B(n29802), .Z(n29804) );
  NANDN U31192 ( .A(n29805), .B(n29804), .Z(n29923) );
  NANDN U31193 ( .A(n29807), .B(n29806), .Z(n29811) );
  NANDN U31194 ( .A(n29809), .B(n29808), .Z(n29810) );
  AND U31195 ( .A(n29811), .B(n29810), .Z(n29920) );
  AND U31196 ( .A(x[488]), .B(y[7985]), .Z(n29914) );
  XOR U31197 ( .A(n29912), .B(n29812), .Z(n29913) );
  XOR U31198 ( .A(n29914), .B(n29913), .Z(n29918) );
  ANDN U31199 ( .B(o[312]), .A(n29813), .Z(n29907) );
  AND U31200 ( .A(x[505]), .B(y[7968]), .Z(n29906) );
  NAND U31201 ( .A(x[480]), .B(y[7993]), .Z(n29905) );
  XOR U31202 ( .A(n29906), .B(n29905), .Z(n29908) );
  XNOR U31203 ( .A(n29907), .B(n29908), .Z(n29917) );
  XOR U31204 ( .A(n29918), .B(n29917), .Z(n29919) );
  XOR U31205 ( .A(n29926), .B(n29925), .Z(n29937) );
  XOR U31206 ( .A(n29938), .B(n29937), .Z(n29890) );
  AND U31207 ( .A(n29815), .B(n29814), .Z(n29819) );
  NAND U31208 ( .A(n29817), .B(n29816), .Z(n29818) );
  NANDN U31209 ( .A(n29819), .B(n29818), .Z(n30000) );
  NANDN U31210 ( .A(n29821), .B(n29820), .Z(n29825) );
  NANDN U31211 ( .A(n29823), .B(n29822), .Z(n29824) );
  NAND U31212 ( .A(n29825), .B(n29824), .Z(n29998) );
  AND U31213 ( .A(x[494]), .B(y[7979]), .Z(n29956) );
  AND U31214 ( .A(x[482]), .B(y[7991]), .Z(n29955) );
  XOR U31215 ( .A(n29956), .B(n29955), .Z(n29958) );
  AND U31216 ( .A(x[483]), .B(y[7990]), .Z(n29957) );
  XOR U31217 ( .A(n29958), .B(n29957), .Z(n29997) );
  XOR U31218 ( .A(n29998), .B(n29997), .Z(n29999) );
  XNOR U31219 ( .A(n30000), .B(n29999), .Z(n29887) );
  NANDN U31220 ( .A(n29827), .B(n29826), .Z(n29831) );
  NAND U31221 ( .A(n29829), .B(n29828), .Z(n29830) );
  AND U31222 ( .A(n29831), .B(n29830), .Z(n29888) );
  XOR U31223 ( .A(n29887), .B(n29888), .Z(n29889) );
  NAND U31224 ( .A(n29833), .B(n29832), .Z(n29837) );
  NAND U31225 ( .A(n29835), .B(n29834), .Z(n29836) );
  AND U31226 ( .A(n29837), .B(n29836), .Z(n29894) );
  XOR U31227 ( .A(n29893), .B(n29894), .Z(n29896) );
  NAND U31228 ( .A(n29839), .B(n29838), .Z(n29843) );
  NAND U31229 ( .A(n29841), .B(n29840), .Z(n29842) );
  AND U31230 ( .A(n29843), .B(n29842), .Z(n29895) );
  XNOR U31231 ( .A(n29896), .B(n29895), .Z(n29876) );
  NAND U31232 ( .A(n29845), .B(n29844), .Z(n29849) );
  NAND U31233 ( .A(n29847), .B(n29846), .Z(n29848) );
  AND U31234 ( .A(n29849), .B(n29848), .Z(n29875) );
  XOR U31235 ( .A(n29876), .B(n29875), .Z(n29877) );
  XNOR U31236 ( .A(n29878), .B(n29877), .Z(n29867) );
  NAND U31237 ( .A(n29851), .B(n29850), .Z(n29855) );
  NAND U31238 ( .A(n29853), .B(n29852), .Z(n29854) );
  NAND U31239 ( .A(n29855), .B(n29854), .Z(n29866) );
  XOR U31240 ( .A(n29867), .B(n29866), .Z(n29868) );
  XOR U31241 ( .A(n29869), .B(n29868), .Z(n29874) );
  NAND U31242 ( .A(n29857), .B(n29856), .Z(n29861) );
  NAND U31243 ( .A(n29859), .B(n29858), .Z(n29860) );
  NAND U31244 ( .A(n29861), .B(n29860), .Z(n29873) );
  XOR U31245 ( .A(n29873), .B(n29872), .Z(n29865) );
  XNOR U31246 ( .A(n29874), .B(n29865), .Z(N634) );
  NAND U31247 ( .A(n29867), .B(n29866), .Z(n29871) );
  NAND U31248 ( .A(n29869), .B(n29868), .Z(n29870) );
  NAND U31249 ( .A(n29871), .B(n29870), .Z(n30172) );
  IV U31250 ( .A(n30172), .Z(n30170) );
  NAND U31251 ( .A(n29876), .B(n29875), .Z(n29880) );
  NAND U31252 ( .A(n29878), .B(n29877), .Z(n29879) );
  NAND U31253 ( .A(n29880), .B(n29879), .Z(n30165) );
  NANDN U31254 ( .A(n29882), .B(n29881), .Z(n29886) );
  NAND U31255 ( .A(n29884), .B(n29883), .Z(n29885) );
  AND U31256 ( .A(n29886), .B(n29885), .Z(n30164) );
  XOR U31257 ( .A(n30165), .B(n30164), .Z(n30167) );
  NAND U31258 ( .A(n29888), .B(n29887), .Z(n29892) );
  NANDN U31259 ( .A(n29890), .B(n29889), .Z(n29891) );
  AND U31260 ( .A(n29892), .B(n29891), .Z(n30016) );
  NAND U31261 ( .A(n29894), .B(n29893), .Z(n29898) );
  NAND U31262 ( .A(n29896), .B(n29895), .Z(n29897) );
  AND U31263 ( .A(n29898), .B(n29897), .Z(n30017) );
  XOR U31264 ( .A(n30016), .B(n30017), .Z(n30019) );
  NAND U31265 ( .A(n29900), .B(n29899), .Z(n29904) );
  NAND U31266 ( .A(n29902), .B(n29901), .Z(n29903) );
  NAND U31267 ( .A(n29904), .B(n29903), .Z(n30161) );
  AND U31268 ( .A(x[482]), .B(y[7992]), .Z(n30040) );
  XOR U31269 ( .A(n30041), .B(n30040), .Z(n30043) );
  NAND U31270 ( .A(x[504]), .B(y[7970]), .Z(n30042) );
  XNOR U31271 ( .A(n30043), .B(n30042), .Z(n30082) );
  NANDN U31272 ( .A(n29906), .B(n29905), .Z(n29910) );
  OR U31273 ( .A(n29908), .B(n29907), .Z(n29909) );
  NAND U31274 ( .A(n29910), .B(n29909), .Z(n30083) );
  XNOR U31275 ( .A(n30082), .B(n30083), .Z(n30085) );
  NANDN U31276 ( .A(n29912), .B(n29911), .Z(n29916) );
  NANDN U31277 ( .A(n29914), .B(n29913), .Z(n29915) );
  AND U31278 ( .A(n29916), .B(n29915), .Z(n30084) );
  XOR U31279 ( .A(n30085), .B(n30084), .Z(n30147) );
  NAND U31280 ( .A(n29918), .B(n29917), .Z(n29922) );
  NANDN U31281 ( .A(n29920), .B(n29919), .Z(n29921) );
  AND U31282 ( .A(n29922), .B(n29921), .Z(n30146) );
  NANDN U31283 ( .A(n29924), .B(n29923), .Z(n29928) );
  NAND U31284 ( .A(n29926), .B(n29925), .Z(n29927) );
  NAND U31285 ( .A(n29928), .B(n29927), .Z(n30149) );
  NAND U31286 ( .A(n29930), .B(n29929), .Z(n29934) );
  NAND U31287 ( .A(n29932), .B(n29931), .Z(n29933) );
  NAND U31288 ( .A(n29934), .B(n29933), .Z(n30153) );
  NAND U31289 ( .A(n29936), .B(n29935), .Z(n29940) );
  NAND U31290 ( .A(n29938), .B(n29937), .Z(n29939) );
  AND U31291 ( .A(n29940), .B(n29939), .Z(n30152) );
  XOR U31292 ( .A(n30153), .B(n30152), .Z(n30154) );
  XNOR U31293 ( .A(n30155), .B(n30154), .Z(n30159) );
  NAND U31294 ( .A(n29942), .B(n29941), .Z(n29946) );
  NAND U31295 ( .A(n29944), .B(n29943), .Z(n29945) );
  NAND U31296 ( .A(n29946), .B(n29945), .Z(n30025) );
  AND U31297 ( .A(y[7988]), .B(x[486]), .Z(n29948) );
  NAND U31298 ( .A(y[7986]), .B(x[488]), .Z(n29947) );
  XNOR U31299 ( .A(n29948), .B(n29947), .Z(n30141) );
  NAND U31300 ( .A(x[489]), .B(y[7985]), .Z(n30142) );
  XNOR U31301 ( .A(n30141), .B(n30142), .Z(n30114) );
  AND U31302 ( .A(x[487]), .B(y[7987]), .Z(n30115) );
  XOR U31303 ( .A(n30114), .B(n30115), .Z(n30116) );
  AND U31304 ( .A(x[492]), .B(y[7982]), .Z(n30241) );
  AND U31305 ( .A(x[485]), .B(y[7989]), .Z(n30097) );
  XOR U31306 ( .A(n30241), .B(n30097), .Z(n30099) );
  NAND U31307 ( .A(x[490]), .B(y[7984]), .Z(n30098) );
  XNOR U31308 ( .A(n30099), .B(n30098), .Z(n30117) );
  XOR U31309 ( .A(n30116), .B(n30117), .Z(n30066) );
  NAND U31310 ( .A(n29950), .B(n29949), .Z(n29954) );
  NAND U31311 ( .A(n29952), .B(n29951), .Z(n29953) );
  NAND U31312 ( .A(n29954), .B(n29953), .Z(n30065) );
  NAND U31313 ( .A(n29956), .B(n29955), .Z(n29960) );
  NAND U31314 ( .A(n29958), .B(n29957), .Z(n29959) );
  NAND U31315 ( .A(n29960), .B(n29959), .Z(n30064) );
  XNOR U31316 ( .A(n30065), .B(n30064), .Z(n30067) );
  NAND U31317 ( .A(n29962), .B(n29961), .Z(n29966) );
  NAND U31318 ( .A(n29964), .B(n29963), .Z(n29965) );
  AND U31319 ( .A(n29966), .B(n29965), .Z(n30070) );
  NANDN U31320 ( .A(n29968), .B(n29967), .Z(n29972) );
  OR U31321 ( .A(n29970), .B(n29969), .Z(n29971) );
  AND U31322 ( .A(n29972), .B(n29971), .Z(n30028) );
  NANDN U31323 ( .A(n29974), .B(n29973), .Z(n29978) );
  OR U31324 ( .A(n29976), .B(n29975), .Z(n29977) );
  NAND U31325 ( .A(n29978), .B(n29977), .Z(n30029) );
  XNOR U31326 ( .A(n30028), .B(n30029), .Z(n30030) );
  ANDN U31327 ( .B(o[313]), .A(n29979), .Z(n30134) );
  NAND U31328 ( .A(x[494]), .B(y[7980]), .Z(n30135) );
  XNOR U31329 ( .A(n30134), .B(n30135), .Z(n30136) );
  NAND U31330 ( .A(x[481]), .B(y[7993]), .Z(n30137) );
  XNOR U31331 ( .A(n30136), .B(n30137), .Z(n30088) );
  NAND U31332 ( .A(x[505]), .B(y[7969]), .Z(n30145) );
  XNOR U31333 ( .A(o[314]), .B(n30145), .Z(n30102) );
  NAND U31334 ( .A(x[506]), .B(y[7968]), .Z(n30103) );
  XNOR U31335 ( .A(n30102), .B(n30103), .Z(n30104) );
  NAND U31336 ( .A(x[480]), .B(y[7994]), .Z(n30105) );
  XOR U31337 ( .A(n30104), .B(n30105), .Z(n30089) );
  XNOR U31338 ( .A(n30088), .B(n30089), .Z(n30090) );
  NANDN U31339 ( .A(n29981), .B(n29980), .Z(n29985) );
  NANDN U31340 ( .A(n29983), .B(n29982), .Z(n29984) );
  NAND U31341 ( .A(n29985), .B(n29984), .Z(n30091) );
  XOR U31342 ( .A(n30090), .B(n30091), .Z(n30031) );
  XOR U31343 ( .A(n30030), .B(n30031), .Z(n30078) );
  AND U31344 ( .A(x[501]), .B(y[7973]), .Z(n30128) );
  NANDN U31345 ( .A(n29986), .B(n30128), .Z(n29990) );
  NAND U31346 ( .A(n29988), .B(n29987), .Z(n29989) );
  NAND U31347 ( .A(n29990), .B(n29989), .Z(n30060) );
  XOR U31348 ( .A(n30129), .B(n30128), .Z(n30131) );
  NAND U31349 ( .A(x[500]), .B(y[7974]), .Z(n30130) );
  XNOR U31350 ( .A(n30131), .B(n30130), .Z(n30059) );
  NAND U31351 ( .A(x[503]), .B(y[7971]), .Z(n30047) );
  XNOR U31352 ( .A(n30046), .B(n30047), .Z(n30049) );
  AND U31353 ( .A(x[502]), .B(y[7972]), .Z(n30048) );
  XOR U31354 ( .A(n30049), .B(n30048), .Z(n30058) );
  XOR U31355 ( .A(n30059), .B(n30058), .Z(n30061) );
  XOR U31356 ( .A(n30060), .B(n30061), .Z(n30077) );
  AND U31357 ( .A(x[484]), .B(y[7990]), .Z(n30052) );
  XOR U31358 ( .A(n30053), .B(n30052), .Z(n30055) );
  AND U31359 ( .A(x[491]), .B(y[7983]), .Z(n30120) );
  NAND U31360 ( .A(x[483]), .B(y[7991]), .Z(n30121) );
  XNOR U31361 ( .A(n30120), .B(n30121), .Z(n30122) );
  NAND U31362 ( .A(x[499]), .B(y[7975]), .Z(n30123) );
  XOR U31363 ( .A(n30122), .B(n30123), .Z(n30035) );
  XNOR U31364 ( .A(n30034), .B(n30035), .Z(n30037) );
  NANDN U31365 ( .A(n29992), .B(n29991), .Z(n29996) );
  OR U31366 ( .A(n29994), .B(n29993), .Z(n29995) );
  AND U31367 ( .A(n29996), .B(n29995), .Z(n30036) );
  XNOR U31368 ( .A(n30037), .B(n30036), .Z(n30076) );
  XOR U31369 ( .A(n30078), .B(n30079), .Z(n30072) );
  XNOR U31370 ( .A(n30073), .B(n30072), .Z(n30023) );
  NAND U31371 ( .A(n29998), .B(n29997), .Z(n30002) );
  NAND U31372 ( .A(n30000), .B(n29999), .Z(n30001) );
  NAND U31373 ( .A(n30002), .B(n30001), .Z(n30111) );
  NANDN U31374 ( .A(n30004), .B(n30003), .Z(n30008) );
  NANDN U31375 ( .A(n30006), .B(n30005), .Z(n30007) );
  NAND U31376 ( .A(n30008), .B(n30007), .Z(n30109) );
  NANDN U31377 ( .A(n30010), .B(n30009), .Z(n30014) );
  NANDN U31378 ( .A(n30012), .B(n30011), .Z(n30013) );
  NAND U31379 ( .A(n30014), .B(n30013), .Z(n30108) );
  XOR U31380 ( .A(n30109), .B(n30108), .Z(n30110) );
  XOR U31381 ( .A(n30111), .B(n30110), .Z(n30022) );
  XOR U31382 ( .A(n30023), .B(n30022), .Z(n30024) );
  XOR U31383 ( .A(n30025), .B(n30024), .Z(n30158) );
  XOR U31384 ( .A(n30159), .B(n30158), .Z(n30160) );
  XOR U31385 ( .A(n30161), .B(n30160), .Z(n30018) );
  XOR U31386 ( .A(n30019), .B(n30018), .Z(n30166) );
  XOR U31387 ( .A(n30167), .B(n30166), .Z(n30173) );
  XNOR U31388 ( .A(n30171), .B(n30173), .Z(n30015) );
  XOR U31389 ( .A(n30170), .B(n30015), .Z(N635) );
  NAND U31390 ( .A(n30017), .B(n30016), .Z(n30021) );
  NAND U31391 ( .A(n30019), .B(n30018), .Z(n30020) );
  AND U31392 ( .A(n30021), .B(n30020), .Z(n30181) );
  NAND U31393 ( .A(n30023), .B(n30022), .Z(n30027) );
  NAND U31394 ( .A(n30025), .B(n30024), .Z(n30026) );
  NAND U31395 ( .A(n30027), .B(n30026), .Z(n30195) );
  NANDN U31396 ( .A(n30029), .B(n30028), .Z(n30033) );
  NANDN U31397 ( .A(n30031), .B(n30030), .Z(n30032) );
  AND U31398 ( .A(n30033), .B(n30032), .Z(n30313) );
  NANDN U31399 ( .A(n30035), .B(n30034), .Z(n30039) );
  NAND U31400 ( .A(n30037), .B(n30036), .Z(n30038) );
  AND U31401 ( .A(n30039), .B(n30038), .Z(n30311) );
  NAND U31402 ( .A(n30041), .B(n30040), .Z(n30045) );
  ANDN U31403 ( .B(n30043), .A(n30042), .Z(n30044) );
  ANDN U31404 ( .B(n30045), .A(n30044), .Z(n30212) );
  NANDN U31405 ( .A(n30047), .B(n30046), .Z(n30051) );
  NAND U31406 ( .A(n30049), .B(n30048), .Z(n30050) );
  NAND U31407 ( .A(n30051), .B(n30050), .Z(n30211) );
  XNOR U31408 ( .A(n30212), .B(n30211), .Z(n30213) );
  NAND U31409 ( .A(n30053), .B(n30052), .Z(n30057) );
  ANDN U31410 ( .B(n30055), .A(n30054), .Z(n30056) );
  ANDN U31411 ( .B(n30057), .A(n30056), .Z(n30226) );
  AND U31412 ( .A(x[480]), .B(y[7995]), .Z(n30289) );
  NAND U31413 ( .A(x[507]), .B(y[7968]), .Z(n30290) );
  XNOR U31414 ( .A(n30289), .B(n30290), .Z(n30291) );
  AND U31415 ( .A(x[506]), .B(y[7969]), .Z(n30301) );
  XNOR U31416 ( .A(o[315]), .B(n30301), .Z(n30292) );
  XNOR U31417 ( .A(n30291), .B(n30292), .Z(n30223) );
  AND U31418 ( .A(x[489]), .B(y[7986]), .Z(n30295) );
  NAND U31419 ( .A(x[501]), .B(y[7974]), .Z(n30296) );
  XNOR U31420 ( .A(n30295), .B(n30296), .Z(n30297) );
  NAND U31421 ( .A(x[498]), .B(y[7977]), .Z(n30298) );
  XOR U31422 ( .A(n30297), .B(n30298), .Z(n30224) );
  XNOR U31423 ( .A(n30223), .B(n30224), .Z(n30225) );
  XOR U31424 ( .A(n30226), .B(n30225), .Z(n30214) );
  XNOR U31425 ( .A(n30213), .B(n30214), .Z(n30310) );
  XNOR U31426 ( .A(n30311), .B(n30310), .Z(n30312) );
  XOR U31427 ( .A(n30313), .B(n30312), .Z(n30330) );
  NAND U31428 ( .A(n30059), .B(n30058), .Z(n30063) );
  NAND U31429 ( .A(n30061), .B(n30060), .Z(n30062) );
  AND U31430 ( .A(n30063), .B(n30062), .Z(n30329) );
  NAND U31431 ( .A(n30065), .B(n30064), .Z(n30069) );
  NANDN U31432 ( .A(n30067), .B(n30066), .Z(n30068) );
  AND U31433 ( .A(n30069), .B(n30068), .Z(n30328) );
  XOR U31434 ( .A(n30329), .B(n30328), .Z(n30331) );
  XOR U31435 ( .A(n30330), .B(n30331), .Z(n30194) );
  NANDN U31436 ( .A(n30071), .B(n30070), .Z(n30075) );
  NAND U31437 ( .A(n30073), .B(n30072), .Z(n30074) );
  AND U31438 ( .A(n30075), .B(n30074), .Z(n30319) );
  NANDN U31439 ( .A(n30077), .B(n30076), .Z(n30081) );
  NAND U31440 ( .A(n30079), .B(n30078), .Z(n30080) );
  AND U31441 ( .A(n30081), .B(n30080), .Z(n30317) );
  NANDN U31442 ( .A(n30083), .B(n30082), .Z(n30087) );
  NAND U31443 ( .A(n30085), .B(n30084), .Z(n30086) );
  AND U31444 ( .A(n30087), .B(n30086), .Z(n30307) );
  NANDN U31445 ( .A(n30089), .B(n30088), .Z(n30093) );
  NANDN U31446 ( .A(n30091), .B(n30090), .Z(n30092) );
  AND U31447 ( .A(n30093), .B(n30092), .Z(n30305) );
  AND U31448 ( .A(x[499]), .B(y[7976]), .Z(n30277) );
  NAND U31449 ( .A(x[505]), .B(y[7970]), .Z(n30278) );
  XNOR U31450 ( .A(n30277), .B(n30278), .Z(n30279) );
  NAND U31451 ( .A(x[486]), .B(y[7989]), .Z(n30280) );
  XNOR U31452 ( .A(n30279), .B(n30280), .Z(n30266) );
  AND U31453 ( .A(x[495]), .B(y[7980]), .Z(n30246) );
  NAND U31454 ( .A(x[482]), .B(y[7993]), .Z(n30247) );
  NAND U31455 ( .A(x[483]), .B(y[7992]), .Z(n30249) );
  XNOR U31456 ( .A(n30266), .B(n30267), .Z(n30268) );
  NAND U31457 ( .A(x[496]), .B(y[7979]), .Z(n30229) );
  XNOR U31458 ( .A(n30229), .B(n30230), .Z(n30231) );
  XNOR U31459 ( .A(n30094), .B(n30231), .Z(n30242) );
  AND U31460 ( .A(y[7982]), .B(x[493]), .Z(n30096) );
  NAND U31461 ( .A(y[7983]), .B(x[492]), .Z(n30095) );
  XNOR U31462 ( .A(n30096), .B(n30095), .Z(n30243) );
  XNOR U31463 ( .A(n30242), .B(n30243), .Z(n30269) );
  XNOR U31464 ( .A(n30268), .B(n30269), .Z(n30207) );
  NAND U31465 ( .A(n30241), .B(n30097), .Z(n30101) );
  ANDN U31466 ( .B(n30099), .A(n30098), .Z(n30100) );
  ANDN U31467 ( .B(n30101), .A(n30100), .Z(n30206) );
  NANDN U31468 ( .A(n30103), .B(n30102), .Z(n30107) );
  NANDN U31469 ( .A(n30105), .B(n30104), .Z(n30106) );
  NAND U31470 ( .A(n30107), .B(n30106), .Z(n30205) );
  XOR U31471 ( .A(n30206), .B(n30205), .Z(n30208) );
  XNOR U31472 ( .A(n30207), .B(n30208), .Z(n30304) );
  XNOR U31473 ( .A(n30305), .B(n30304), .Z(n30306) );
  XNOR U31474 ( .A(n30307), .B(n30306), .Z(n30316) );
  XOR U31475 ( .A(n30317), .B(n30316), .Z(n30318) );
  XOR U31476 ( .A(n30319), .B(n30318), .Z(n30193) );
  XOR U31477 ( .A(n30195), .B(n30196), .Z(n30190) );
  NAND U31478 ( .A(n30109), .B(n30108), .Z(n30113) );
  NAND U31479 ( .A(n30111), .B(n30110), .Z(n30112) );
  NAND U31480 ( .A(n30113), .B(n30112), .Z(n30201) );
  NAND U31481 ( .A(n30115), .B(n30114), .Z(n30119) );
  NAND U31482 ( .A(n30117), .B(n30116), .Z(n30118) );
  AND U31483 ( .A(n30119), .B(n30118), .Z(n30324) );
  NANDN U31484 ( .A(n30121), .B(n30120), .Z(n30125) );
  NANDN U31485 ( .A(n30123), .B(n30122), .Z(n30124) );
  AND U31486 ( .A(n30125), .B(n30124), .Z(n30265) );
  AND U31487 ( .A(y[7971]), .B(x[504]), .Z(n30127) );
  NAND U31488 ( .A(y[7975]), .B(x[500]), .Z(n30126) );
  XNOR U31489 ( .A(n30127), .B(n30126), .Z(n30273) );
  NAND U31490 ( .A(x[487]), .B(y[7988]), .Z(n30274) );
  XNOR U31491 ( .A(n30273), .B(n30274), .Z(n30263) );
  AND U31492 ( .A(x[488]), .B(y[7987]), .Z(n30235) );
  AND U31493 ( .A(x[503]), .B(y[7972]), .Z(n30236) );
  XOR U31494 ( .A(n30235), .B(n30236), .Z(n30237) );
  AND U31495 ( .A(x[502]), .B(y[7973]), .Z(n30238) );
  XOR U31496 ( .A(n30237), .B(n30238), .Z(n30262) );
  XOR U31497 ( .A(n30263), .B(n30262), .Z(n30264) );
  XOR U31498 ( .A(n30265), .B(n30264), .Z(n30322) );
  NAND U31499 ( .A(n30129), .B(n30128), .Z(n30133) );
  ANDN U31500 ( .B(n30131), .A(n30130), .Z(n30132) );
  ANDN U31501 ( .B(n30133), .A(n30132), .Z(n30259) );
  NANDN U31502 ( .A(n30135), .B(n30134), .Z(n30139) );
  NANDN U31503 ( .A(n30137), .B(n30136), .Z(n30138) );
  NAND U31504 ( .A(n30139), .B(n30138), .Z(n30258) );
  XNOR U31505 ( .A(n30259), .B(n30258), .Z(n30261) );
  AND U31506 ( .A(y[7988]), .B(x[488]), .Z(n30303) );
  NAND U31507 ( .A(n30140), .B(n30303), .Z(n30144) );
  NANDN U31508 ( .A(n30142), .B(n30141), .Z(n30143) );
  NAND U31509 ( .A(n30144), .B(n30143), .Z(n30219) );
  AND U31510 ( .A(x[494]), .B(y[7981]), .Z(n30252) );
  NAND U31511 ( .A(x[481]), .B(y[7994]), .Z(n30253) );
  ANDN U31512 ( .B(o[314]), .A(n30145), .Z(n30254) );
  XOR U31513 ( .A(n30255), .B(n30254), .Z(n30218) );
  AND U31514 ( .A(x[497]), .B(y[7978]), .Z(n30283) );
  NAND U31515 ( .A(x[484]), .B(y[7991]), .Z(n30284) );
  XNOR U31516 ( .A(n30283), .B(n30284), .Z(n30286) );
  AND U31517 ( .A(x[485]), .B(y[7990]), .Z(n30285) );
  XOR U31518 ( .A(n30286), .B(n30285), .Z(n30217) );
  XOR U31519 ( .A(n30218), .B(n30217), .Z(n30220) );
  XOR U31520 ( .A(n30219), .B(n30220), .Z(n30260) );
  XOR U31521 ( .A(n30261), .B(n30260), .Z(n30323) );
  XNOR U31522 ( .A(n30324), .B(n30325), .Z(n30200) );
  NANDN U31523 ( .A(n30147), .B(n30146), .Z(n30151) );
  NANDN U31524 ( .A(n30149), .B(n30148), .Z(n30150) );
  AND U31525 ( .A(n30151), .B(n30150), .Z(n30199) );
  XOR U31526 ( .A(n30201), .B(n30202), .Z(n30187) );
  NAND U31527 ( .A(n30153), .B(n30152), .Z(n30157) );
  NAND U31528 ( .A(n30155), .B(n30154), .Z(n30156) );
  AND U31529 ( .A(n30157), .B(n30156), .Z(n30188) );
  XOR U31530 ( .A(n30187), .B(n30188), .Z(n30189) );
  XNOR U31531 ( .A(n30190), .B(n30189), .Z(n30179) );
  NAND U31532 ( .A(n30159), .B(n30158), .Z(n30163) );
  NAND U31533 ( .A(n30161), .B(n30160), .Z(n30162) );
  AND U31534 ( .A(n30163), .B(n30162), .Z(n30178) );
  XOR U31535 ( .A(n30179), .B(n30178), .Z(n30180) );
  XOR U31536 ( .A(n30181), .B(n30180), .Z(n30186) );
  NAND U31537 ( .A(n30165), .B(n30164), .Z(n30169) );
  NAND U31538 ( .A(n30167), .B(n30166), .Z(n30168) );
  NAND U31539 ( .A(n30169), .B(n30168), .Z(n30185) );
  NANDN U31540 ( .A(n30170), .B(n30171), .Z(n30176) );
  NOR U31541 ( .A(n30172), .B(n30171), .Z(n30174) );
  OR U31542 ( .A(n30174), .B(n30173), .Z(n30175) );
  AND U31543 ( .A(n30176), .B(n30175), .Z(n30184) );
  XOR U31544 ( .A(n30185), .B(n30184), .Z(n30177) );
  XNOR U31545 ( .A(n30186), .B(n30177), .Z(N636) );
  NAND U31546 ( .A(n30179), .B(n30178), .Z(n30183) );
  NAND U31547 ( .A(n30181), .B(n30180), .Z(n30182) );
  NAND U31548 ( .A(n30183), .B(n30182), .Z(n30500) );
  IV U31549 ( .A(n30500), .Z(n30498) );
  NAND U31550 ( .A(n30188), .B(n30187), .Z(n30192) );
  NAND U31551 ( .A(n30190), .B(n30189), .Z(n30191) );
  NAND U31552 ( .A(n30192), .B(n30191), .Z(n30493) );
  NANDN U31553 ( .A(n30194), .B(n30193), .Z(n30198) );
  NAND U31554 ( .A(n30196), .B(n30195), .Z(n30197) );
  NAND U31555 ( .A(n30198), .B(n30197), .Z(n30492) );
  XOR U31556 ( .A(n30493), .B(n30492), .Z(n30495) );
  NANDN U31557 ( .A(n30200), .B(n30199), .Z(n30204) );
  NAND U31558 ( .A(n30202), .B(n30201), .Z(n30203) );
  NAND U31559 ( .A(n30204), .B(n30203), .Z(n30335) );
  NANDN U31560 ( .A(n30206), .B(n30205), .Z(n30210) );
  NANDN U31561 ( .A(n30208), .B(n30207), .Z(n30209) );
  AND U31562 ( .A(n30210), .B(n30209), .Z(n30360) );
  NANDN U31563 ( .A(n30212), .B(n30211), .Z(n30216) );
  NANDN U31564 ( .A(n30214), .B(n30213), .Z(n30215) );
  AND U31565 ( .A(n30216), .B(n30215), .Z(n30465) );
  NAND U31566 ( .A(n30218), .B(n30217), .Z(n30222) );
  NAND U31567 ( .A(n30220), .B(n30219), .Z(n30221) );
  AND U31568 ( .A(n30222), .B(n30221), .Z(n30463) );
  NANDN U31569 ( .A(n30224), .B(n30223), .Z(n30228) );
  NANDN U31570 ( .A(n30226), .B(n30225), .Z(n30227) );
  NAND U31571 ( .A(n30228), .B(n30227), .Z(n30462) );
  XNOR U31572 ( .A(n30463), .B(n30462), .Z(n30464) );
  XNOR U31573 ( .A(n30465), .B(n30464), .Z(n30359) );
  XNOR U31574 ( .A(n30360), .B(n30359), .Z(n30362) );
  NANDN U31575 ( .A(n30230), .B(n30229), .Z(n30234) );
  NANDN U31576 ( .A(n30232), .B(n30231), .Z(n30233) );
  AND U31577 ( .A(n30234), .B(n30233), .Z(n30427) );
  AND U31578 ( .A(x[487]), .B(y[7989]), .Z(n30407) );
  AND U31579 ( .A(x[492]), .B(y[7984]), .Z(n30406) );
  XOR U31580 ( .A(n30407), .B(n30406), .Z(n30409) );
  AND U31581 ( .A(x[491]), .B(y[7985]), .Z(n30408) );
  XOR U31582 ( .A(n30409), .B(n30408), .Z(n30425) );
  AND U31583 ( .A(x[507]), .B(y[7969]), .Z(n30423) );
  XOR U31584 ( .A(o[316]), .B(n30423), .Z(n30437) );
  AND U31585 ( .A(x[506]), .B(y[7970]), .Z(n30436) );
  XOR U31586 ( .A(n30437), .B(n30436), .Z(n30439) );
  AND U31587 ( .A(x[495]), .B(y[7981]), .Z(n30438) );
  XNOR U31588 ( .A(n30439), .B(n30438), .Z(n30424) );
  NAND U31589 ( .A(n30236), .B(n30235), .Z(n30240) );
  NAND U31590 ( .A(n30238), .B(n30237), .Z(n30239) );
  AND U31591 ( .A(n30240), .B(n30239), .Z(n30447) );
  AND U31592 ( .A(x[497]), .B(y[7979]), .Z(n30372) );
  AND U31593 ( .A(x[502]), .B(y[7974]), .Z(n30371) );
  XOR U31594 ( .A(n30372), .B(n30371), .Z(n30374) );
  AND U31595 ( .A(x[484]), .B(y[7992]), .Z(n30373) );
  XOR U31596 ( .A(n30374), .B(n30373), .Z(n30445) );
  AND U31597 ( .A(x[486]), .B(y[7990]), .Z(n30611) );
  NAND U31598 ( .A(x[499]), .B(y[7977]), .Z(n30412) );
  XOR U31599 ( .A(n30445), .B(n30444), .Z(n30446) );
  XOR U31600 ( .A(n30469), .B(n30468), .Z(n30470) );
  NAND U31601 ( .A(n30430), .B(n30241), .Z(n30245) );
  NAND U31602 ( .A(n30243), .B(n30242), .Z(n30244) );
  AND U31603 ( .A(n30245), .B(n30244), .Z(n30368) );
  NANDN U31604 ( .A(n30247), .B(n30246), .Z(n30251) );
  NANDN U31605 ( .A(n30249), .B(n30248), .Z(n30250) );
  AND U31606 ( .A(n30251), .B(n30250), .Z(n30366) );
  NANDN U31607 ( .A(n30253), .B(n30252), .Z(n30257) );
  NAND U31608 ( .A(n30255), .B(n30254), .Z(n30256) );
  NAND U31609 ( .A(n30257), .B(n30256), .Z(n30365) );
  XNOR U31610 ( .A(n30470), .B(n30471), .Z(n30361) );
  XOR U31611 ( .A(n30362), .B(n30361), .Z(n30355) );
  NANDN U31612 ( .A(n30267), .B(n30266), .Z(n30271) );
  NANDN U31613 ( .A(n30269), .B(n30268), .Z(n30270) );
  NAND U31614 ( .A(n30271), .B(n30270), .Z(n30450) );
  XOR U31615 ( .A(n30451), .B(n30450), .Z(n30453) );
  XOR U31616 ( .A(n30452), .B(n30453), .Z(n30354) );
  AND U31617 ( .A(x[504]), .B(y[7975]), .Z(n30795) );
  AND U31618 ( .A(x[500]), .B(y[7971]), .Z(n30272) );
  NAND U31619 ( .A(n30795), .B(n30272), .Z(n30276) );
  NANDN U31620 ( .A(n30274), .B(n30273), .Z(n30275) );
  AND U31621 ( .A(n30276), .B(n30275), .Z(n30489) );
  AND U31622 ( .A(x[505]), .B(y[7971]), .Z(n30402) );
  XOR U31623 ( .A(n30403), .B(n30402), .Z(n30401) );
  NAND U31624 ( .A(x[481]), .B(y[7995]), .Z(n30400) );
  AND U31625 ( .A(x[496]), .B(y[7980]), .Z(n30394) );
  NAND U31626 ( .A(x[504]), .B(y[7972]), .Z(n30395) );
  NAND U31627 ( .A(x[482]), .B(y[7994]), .Z(n30397) );
  XOR U31628 ( .A(n30487), .B(n30486), .Z(n30488) );
  NANDN U31629 ( .A(n30278), .B(n30277), .Z(n30282) );
  NANDN U31630 ( .A(n30280), .B(n30279), .Z(n30281) );
  AND U31631 ( .A(n30282), .B(n30281), .Z(n30483) );
  NAND U31632 ( .A(x[483]), .B(y[7993]), .Z(n30431) );
  NAND U31633 ( .A(x[503]), .B(y[7973]), .Z(n30433) );
  AND U31634 ( .A(x[485]), .B(y[7991]), .Z(n30417) );
  NAND U31635 ( .A(x[501]), .B(y[7975]), .Z(n30418) );
  NAND U31636 ( .A(x[500]), .B(y[7976]), .Z(n30420) );
  XOR U31637 ( .A(n30481), .B(n30480), .Z(n30482) );
  NANDN U31638 ( .A(n30284), .B(n30283), .Z(n30288) );
  NAND U31639 ( .A(n30286), .B(n30285), .Z(n30287) );
  AND U31640 ( .A(n30288), .B(n30287), .Z(n30475) );
  NANDN U31641 ( .A(n30290), .B(n30289), .Z(n30294) );
  NANDN U31642 ( .A(n30292), .B(n30291), .Z(n30293) );
  NAND U31643 ( .A(n30294), .B(n30293), .Z(n30474) );
  NANDN U31644 ( .A(n30296), .B(n30295), .Z(n30300) );
  NANDN U31645 ( .A(n30298), .B(n30297), .Z(n30299) );
  NAND U31646 ( .A(n30300), .B(n30299), .Z(n30390) );
  AND U31647 ( .A(n30301), .B(o[315]), .Z(n30380) );
  AND U31648 ( .A(x[480]), .B(y[7996]), .Z(n30378) );
  AND U31649 ( .A(x[508]), .B(y[7968]), .Z(n30377) );
  XOR U31650 ( .A(n30378), .B(n30377), .Z(n30379) );
  XOR U31651 ( .A(n30380), .B(n30379), .Z(n30389) );
  NAND U31652 ( .A(y[7986]), .B(x[490]), .Z(n30302) );
  XNOR U31653 ( .A(n30303), .B(n30302), .Z(n30385) );
  AND U31654 ( .A(x[489]), .B(y[7987]), .Z(n30384) );
  XOR U31655 ( .A(n30385), .B(n30384), .Z(n30388) );
  XOR U31656 ( .A(n30389), .B(n30388), .Z(n30391) );
  XOR U31657 ( .A(n30390), .B(n30391), .Z(n30476) );
  XNOR U31658 ( .A(n30477), .B(n30476), .Z(n30456) );
  XOR U31659 ( .A(n30457), .B(n30456), .Z(n30458) );
  XOR U31660 ( .A(n30459), .B(n30458), .Z(n30353) );
  XOR U31661 ( .A(n30354), .B(n30353), .Z(n30356) );
  XOR U31662 ( .A(n30355), .B(n30356), .Z(n30350) );
  NANDN U31663 ( .A(n30305), .B(n30304), .Z(n30309) );
  NANDN U31664 ( .A(n30307), .B(n30306), .Z(n30308) );
  AND U31665 ( .A(n30309), .B(n30308), .Z(n30348) );
  NANDN U31666 ( .A(n30311), .B(n30310), .Z(n30315) );
  NANDN U31667 ( .A(n30313), .B(n30312), .Z(n30314) );
  NAND U31668 ( .A(n30315), .B(n30314), .Z(n30347) );
  XNOR U31669 ( .A(n30348), .B(n30347), .Z(n30349) );
  XNOR U31670 ( .A(n30350), .B(n30349), .Z(n30336) );
  XOR U31671 ( .A(n30335), .B(n30336), .Z(n30337) );
  NAND U31672 ( .A(n30317), .B(n30316), .Z(n30321) );
  NAND U31673 ( .A(n30319), .B(n30318), .Z(n30320) );
  NAND U31674 ( .A(n30321), .B(n30320), .Z(n30343) );
  NANDN U31675 ( .A(n30323), .B(n30322), .Z(n30327) );
  NANDN U31676 ( .A(n30325), .B(n30324), .Z(n30326) );
  AND U31677 ( .A(n30327), .B(n30326), .Z(n30342) );
  NAND U31678 ( .A(n30329), .B(n30328), .Z(n30333) );
  NAND U31679 ( .A(n30331), .B(n30330), .Z(n30332) );
  AND U31680 ( .A(n30333), .B(n30332), .Z(n30341) );
  XOR U31681 ( .A(n30342), .B(n30341), .Z(n30344) );
  XNOR U31682 ( .A(n30343), .B(n30344), .Z(n30338) );
  XOR U31683 ( .A(n30495), .B(n30494), .Z(n30501) );
  XNOR U31684 ( .A(n30499), .B(n30501), .Z(n30334) );
  XOR U31685 ( .A(n30498), .B(n30334), .Z(N637) );
  NAND U31686 ( .A(n30336), .B(n30335), .Z(n30340) );
  NANDN U31687 ( .A(n30338), .B(n30337), .Z(n30339) );
  NAND U31688 ( .A(n30340), .B(n30339), .Z(n30511) );
  NAND U31689 ( .A(n30342), .B(n30341), .Z(n30346) );
  NAND U31690 ( .A(n30344), .B(n30343), .Z(n30345) );
  NAND U31691 ( .A(n30346), .B(n30345), .Z(n30509) );
  NANDN U31692 ( .A(n30348), .B(n30347), .Z(n30352) );
  NANDN U31693 ( .A(n30350), .B(n30349), .Z(n30351) );
  AND U31694 ( .A(n30352), .B(n30351), .Z(n30516) );
  NANDN U31695 ( .A(n30354), .B(n30353), .Z(n30358) );
  OR U31696 ( .A(n30356), .B(n30355), .Z(n30357) );
  AND U31697 ( .A(n30358), .B(n30357), .Z(n30515) );
  XNOR U31698 ( .A(n30516), .B(n30515), .Z(n30518) );
  NANDN U31699 ( .A(n30360), .B(n30359), .Z(n30364) );
  NAND U31700 ( .A(n30362), .B(n30361), .Z(n30363) );
  AND U31701 ( .A(n30364), .B(n30363), .Z(n30528) );
  NANDN U31702 ( .A(n30366), .B(n30365), .Z(n30370) );
  NANDN U31703 ( .A(n30368), .B(n30367), .Z(n30369) );
  AND U31704 ( .A(n30370), .B(n30369), .Z(n30640) );
  NAND U31705 ( .A(n30372), .B(n30371), .Z(n30376) );
  NAND U31706 ( .A(n30374), .B(n30373), .Z(n30375) );
  NAND U31707 ( .A(n30376), .B(n30375), .Z(n30677) );
  NAND U31708 ( .A(n30378), .B(n30377), .Z(n30382) );
  NAND U31709 ( .A(n30380), .B(n30379), .Z(n30381) );
  NAND U31710 ( .A(n30382), .B(n30381), .Z(n30676) );
  XOR U31711 ( .A(n30677), .B(n30676), .Z(n30678) );
  AND U31712 ( .A(y[7988]), .B(x[490]), .Z(n30674) );
  NAND U31713 ( .A(n30383), .B(n30674), .Z(n30387) );
  NAND U31714 ( .A(n30385), .B(n30384), .Z(n30386) );
  NAND U31715 ( .A(n30387), .B(n30386), .Z(n30645) );
  AND U31716 ( .A(x[502]), .B(y[7975]), .Z(n30589) );
  AND U31717 ( .A(x[492]), .B(y[7985]), .Z(n30740) );
  AND U31718 ( .A(x[481]), .B(y[7996]), .Z(n30587) );
  XOR U31719 ( .A(n30740), .B(n30587), .Z(n30588) );
  XOR U31720 ( .A(n30589), .B(n30588), .Z(n30644) );
  AND U31721 ( .A(x[495]), .B(y[7982]), .Z(n30592) );
  XOR U31722 ( .A(n30644), .B(n30643), .Z(n30646) );
  XNOR U31723 ( .A(n30645), .B(n30646), .Z(n30679) );
  NAND U31724 ( .A(n30389), .B(n30388), .Z(n30393) );
  NAND U31725 ( .A(n30391), .B(n30390), .Z(n30392) );
  AND U31726 ( .A(n30393), .B(n30392), .Z(n30637) );
  XOR U31727 ( .A(n30640), .B(n30639), .Z(n30634) );
  NANDN U31728 ( .A(n30395), .B(n30394), .Z(n30399) );
  NANDN U31729 ( .A(n30397), .B(n30396), .Z(n30398) );
  NAND U31730 ( .A(n30399), .B(n30398), .Z(n30650) );
  ANDN U31731 ( .B(n30401), .A(n30400), .Z(n30405) );
  NAND U31732 ( .A(n30403), .B(n30402), .Z(n30404) );
  NANDN U31733 ( .A(n30405), .B(n30404), .Z(n30649) );
  XOR U31734 ( .A(n30650), .B(n30649), .Z(n30651) );
  NAND U31735 ( .A(n30407), .B(n30406), .Z(n30411) );
  NAND U31736 ( .A(n30409), .B(n30408), .Z(n30410) );
  NAND U31737 ( .A(n30411), .B(n30410), .Z(n30553) );
  AND U31738 ( .A(x[491]), .B(y[7986]), .Z(n30608) );
  AND U31739 ( .A(x[483]), .B(y[7994]), .Z(n30606) );
  AND U31740 ( .A(x[497]), .B(y[7980]), .Z(n30605) );
  XOR U31741 ( .A(n30606), .B(n30605), .Z(n30607) );
  XOR U31742 ( .A(n30608), .B(n30607), .Z(n30552) );
  AND U31743 ( .A(x[503]), .B(y[7974]), .Z(n30602) );
  AND U31744 ( .A(x[493]), .B(y[7984]), .Z(n30600) );
  AND U31745 ( .A(x[504]), .B(y[7973]), .Z(n30853) );
  XOR U31746 ( .A(n30600), .B(n30853), .Z(n30601) );
  XOR U31747 ( .A(n30602), .B(n30601), .Z(n30551) );
  XOR U31748 ( .A(n30552), .B(n30551), .Z(n30554) );
  XNOR U31749 ( .A(n30553), .B(n30554), .Z(n30652) );
  NANDN U31750 ( .A(n30412), .B(n30611), .Z(n30416) );
  NANDN U31751 ( .A(n30414), .B(n30413), .Z(n30415) );
  AND U31752 ( .A(n30416), .B(n30415), .Z(n30657) );
  AND U31753 ( .A(x[505]), .B(y[7972]), .Z(n30584) );
  AND U31754 ( .A(x[506]), .B(y[7971]), .Z(n30581) );
  XOR U31755 ( .A(n30582), .B(n30581), .Z(n30583) );
  XOR U31756 ( .A(n30584), .B(n30583), .Z(n30656) );
  AND U31757 ( .A(x[508]), .B(y[7969]), .Z(n30599) );
  XOR U31758 ( .A(o[317]), .B(n30599), .Z(n30669) );
  AND U31759 ( .A(x[480]), .B(y[7997]), .Z(n30667) );
  AND U31760 ( .A(x[509]), .B(y[7968]), .Z(n30666) );
  XOR U31761 ( .A(n30667), .B(n30666), .Z(n30668) );
  XNOR U31762 ( .A(n30669), .B(n30668), .Z(n30655) );
  XNOR U31763 ( .A(n30657), .B(n30658), .Z(n30539) );
  NANDN U31764 ( .A(n30418), .B(n30417), .Z(n30422) );
  NANDN U31765 ( .A(n30420), .B(n30419), .Z(n30421) );
  NAND U31766 ( .A(n30422), .B(n30421), .Z(n30620) );
  AND U31767 ( .A(o[316]), .B(n30423), .Z(n30572) );
  AND U31768 ( .A(x[496]), .B(y[7981]), .Z(n30570) );
  AND U31769 ( .A(x[507]), .B(y[7970]), .Z(n30569) );
  XOR U31770 ( .A(n30570), .B(n30569), .Z(n30571) );
  XOR U31771 ( .A(n30572), .B(n30571), .Z(n30619) );
  AND U31772 ( .A(x[482]), .B(y[7995]), .Z(n30564) );
  XOR U31773 ( .A(n30564), .B(n30563), .Z(n30565) );
  XOR U31774 ( .A(n30566), .B(n30565), .Z(n30618) );
  XOR U31775 ( .A(n30619), .B(n30618), .Z(n30621) );
  XOR U31776 ( .A(n30620), .B(n30621), .Z(n30540) );
  NANDN U31777 ( .A(n30425), .B(n30424), .Z(n30429) );
  NANDN U31778 ( .A(n30427), .B(n30426), .Z(n30428) );
  AND U31779 ( .A(n30429), .B(n30428), .Z(n30546) );
  NANDN U31780 ( .A(n30431), .B(n30430), .Z(n30435) );
  NANDN U31781 ( .A(n30433), .B(n30432), .Z(n30434) );
  NAND U31782 ( .A(n30435), .B(n30434), .Z(n30576) );
  NAND U31783 ( .A(n30437), .B(n30436), .Z(n30441) );
  NAND U31784 ( .A(n30439), .B(n30438), .Z(n30440) );
  NAND U31785 ( .A(n30441), .B(n30440), .Z(n30575) );
  XOR U31786 ( .A(n30576), .B(n30575), .Z(n30578) );
  AND U31787 ( .A(x[489]), .B(y[7988]), .Z(n30790) );
  AND U31788 ( .A(x[488]), .B(y[7989]), .Z(n30613) );
  AND U31789 ( .A(y[7991]), .B(x[486]), .Z(n30443) );
  NAND U31790 ( .A(y[7990]), .B(x[487]), .Z(n30442) );
  XNOR U31791 ( .A(n30443), .B(n30442), .Z(n30612) );
  XOR U31792 ( .A(n30613), .B(n30612), .Z(n30661) );
  XOR U31793 ( .A(n30790), .B(n30661), .Z(n30663) );
  AND U31794 ( .A(x[485]), .B(y[7992]), .Z(n30560) );
  AND U31795 ( .A(x[484]), .B(y[7993]), .Z(n30558) );
  AND U31796 ( .A(x[490]), .B(y[7987]), .Z(n30557) );
  XOR U31797 ( .A(n30558), .B(n30557), .Z(n30559) );
  XOR U31798 ( .A(n30560), .B(n30559), .Z(n30662) );
  XOR U31799 ( .A(n30663), .B(n30662), .Z(n30577) );
  XNOR U31800 ( .A(n30578), .B(n30577), .Z(n30545) );
  XOR U31801 ( .A(n30548), .B(n30547), .Z(n30632) );
  NAND U31802 ( .A(n30445), .B(n30444), .Z(n30449) );
  NANDN U31803 ( .A(n30447), .B(n30446), .Z(n30448) );
  NAND U31804 ( .A(n30449), .B(n30448), .Z(n30631) );
  XNOR U31805 ( .A(n30528), .B(n30527), .Z(n30529) );
  NANDN U31806 ( .A(n30451), .B(n30450), .Z(n30455) );
  OR U31807 ( .A(n30453), .B(n30452), .Z(n30454) );
  AND U31808 ( .A(n30455), .B(n30454), .Z(n30522) );
  NAND U31809 ( .A(n30457), .B(n30456), .Z(n30461) );
  NAND U31810 ( .A(n30459), .B(n30458), .Z(n30460) );
  AND U31811 ( .A(n30461), .B(n30460), .Z(n30521) );
  XNOR U31812 ( .A(n30522), .B(n30521), .Z(n30523) );
  NANDN U31813 ( .A(n30463), .B(n30462), .Z(n30467) );
  NANDN U31814 ( .A(n30465), .B(n30464), .Z(n30466) );
  NAND U31815 ( .A(n30467), .B(n30466), .Z(n30535) );
  NAND U31816 ( .A(n30469), .B(n30468), .Z(n30473) );
  NANDN U31817 ( .A(n30471), .B(n30470), .Z(n30472) );
  NAND U31818 ( .A(n30473), .B(n30472), .Z(n30533) );
  NANDN U31819 ( .A(n30475), .B(n30474), .Z(n30479) );
  NAND U31820 ( .A(n30477), .B(n30476), .Z(n30478) );
  AND U31821 ( .A(n30479), .B(n30478), .Z(n30627) );
  NAND U31822 ( .A(n30481), .B(n30480), .Z(n30485) );
  NANDN U31823 ( .A(n30483), .B(n30482), .Z(n30484) );
  AND U31824 ( .A(n30485), .B(n30484), .Z(n30625) );
  NAND U31825 ( .A(n30487), .B(n30486), .Z(n30491) );
  NANDN U31826 ( .A(n30489), .B(n30488), .Z(n30490) );
  NAND U31827 ( .A(n30491), .B(n30490), .Z(n30624) );
  XOR U31828 ( .A(n30533), .B(n30534), .Z(n30536) );
  XNOR U31829 ( .A(n30535), .B(n30536), .Z(n30524) );
  XOR U31830 ( .A(n30523), .B(n30524), .Z(n30530) );
  XNOR U31831 ( .A(n30529), .B(n30530), .Z(n30517) );
  XOR U31832 ( .A(n30518), .B(n30517), .Z(n30510) );
  XNOR U31833 ( .A(n30509), .B(n30510), .Z(n30512) );
  XOR U31834 ( .A(n30511), .B(n30512), .Z(n30508) );
  NAND U31835 ( .A(n30493), .B(n30492), .Z(n30497) );
  NAND U31836 ( .A(n30495), .B(n30494), .Z(n30496) );
  NAND U31837 ( .A(n30497), .B(n30496), .Z(n30507) );
  NANDN U31838 ( .A(n30498), .B(n30499), .Z(n30504) );
  NOR U31839 ( .A(n30500), .B(n30499), .Z(n30502) );
  OR U31840 ( .A(n30502), .B(n30501), .Z(n30503) );
  AND U31841 ( .A(n30504), .B(n30503), .Z(n30506) );
  XOR U31842 ( .A(n30507), .B(n30506), .Z(n30505) );
  XNOR U31843 ( .A(n30508), .B(n30505), .Z(N638) );
  NAND U31844 ( .A(n30510), .B(n30509), .Z(n30514) );
  NANDN U31845 ( .A(n30512), .B(n30511), .Z(n30513) );
  NAND U31846 ( .A(n30514), .B(n30513), .Z(n30969) );
  NANDN U31847 ( .A(n30516), .B(n30515), .Z(n30520) );
  NAND U31848 ( .A(n30518), .B(n30517), .Z(n30519) );
  AND U31849 ( .A(n30520), .B(n30519), .Z(n30683) );
  NANDN U31850 ( .A(n30522), .B(n30521), .Z(n30526) );
  NANDN U31851 ( .A(n30524), .B(n30523), .Z(n30525) );
  AND U31852 ( .A(n30526), .B(n30525), .Z(n30975) );
  NANDN U31853 ( .A(n30528), .B(n30527), .Z(n30532) );
  NANDN U31854 ( .A(n30530), .B(n30529), .Z(n30531) );
  AND U31855 ( .A(n30532), .B(n30531), .Z(n30974) );
  XOR U31856 ( .A(n30975), .B(n30974), .Z(n30973) );
  NAND U31857 ( .A(n30534), .B(n30533), .Z(n30538) );
  NAND U31858 ( .A(n30536), .B(n30535), .Z(n30537) );
  AND U31859 ( .A(n30538), .B(n30537), .Z(n30972) );
  XOR U31860 ( .A(n30973), .B(n30972), .Z(n30685) );
  NANDN U31861 ( .A(n30540), .B(n30539), .Z(n30544) );
  NANDN U31862 ( .A(n30542), .B(n30541), .Z(n30543) );
  AND U31863 ( .A(n30544), .B(n30543), .Z(n30959) );
  NANDN U31864 ( .A(n30546), .B(n30545), .Z(n30550) );
  NAND U31865 ( .A(n30548), .B(n30547), .Z(n30549) );
  AND U31866 ( .A(n30550), .B(n30549), .Z(n30946) );
  NAND U31867 ( .A(n30552), .B(n30551), .Z(n30556) );
  NAND U31868 ( .A(n30554), .B(n30553), .Z(n30555) );
  AND U31869 ( .A(n30556), .B(n30555), .Z(n30690) );
  NAND U31870 ( .A(n30558), .B(n30557), .Z(n30562) );
  NAND U31871 ( .A(n30560), .B(n30559), .Z(n30561) );
  NAND U31872 ( .A(n30562), .B(n30561), .Z(n30703) );
  AND U31873 ( .A(x[486]), .B(y[7992]), .Z(n30857) );
  AND U31874 ( .A(x[485]), .B(y[7993]), .Z(n30859) );
  AND U31875 ( .A(x[499]), .B(y[7979]), .Z(n30858) );
  XOR U31876 ( .A(n30859), .B(n30858), .Z(n30856) );
  XNOR U31877 ( .A(n30857), .B(n30856), .Z(n30706) );
  AND U31878 ( .A(x[484]), .B(y[7994]), .Z(n30781) );
  AND U31879 ( .A(x[483]), .B(y[7995]), .Z(n30783) );
  AND U31880 ( .A(x[498]), .B(y[7980]), .Z(n30782) );
  XOR U31881 ( .A(n30783), .B(n30782), .Z(n30780) );
  XOR U31882 ( .A(n30781), .B(n30780), .Z(n30709) );
  NAND U31883 ( .A(n30564), .B(n30563), .Z(n30568) );
  NAND U31884 ( .A(n30566), .B(n30565), .Z(n30567) );
  AND U31885 ( .A(n30568), .B(n30567), .Z(n30708) );
  XOR U31886 ( .A(n30706), .B(n30707), .Z(n30702) );
  XOR U31887 ( .A(n30703), .B(n30702), .Z(n30701) );
  NAND U31888 ( .A(n30570), .B(n30569), .Z(n30574) );
  NAND U31889 ( .A(n30572), .B(n30571), .Z(n30573) );
  NAND U31890 ( .A(n30574), .B(n30573), .Z(n30700) );
  XOR U31891 ( .A(n30701), .B(n30700), .Z(n30691) );
  NAND U31892 ( .A(n30576), .B(n30575), .Z(n30580) );
  NAND U31893 ( .A(n30578), .B(n30577), .Z(n30579) );
  AND U31894 ( .A(n30580), .B(n30579), .Z(n30688) );
  XOR U31895 ( .A(n30689), .B(n30688), .Z(n30949) );
  AND U31896 ( .A(n30582), .B(n30581), .Z(n30586) );
  NAND U31897 ( .A(n30584), .B(n30583), .Z(n30585) );
  NANDN U31898 ( .A(n30586), .B(n30585), .Z(n30726) );
  AND U31899 ( .A(n30740), .B(n30587), .Z(n30591) );
  NAND U31900 ( .A(n30589), .B(n30588), .Z(n30590) );
  NANDN U31901 ( .A(n30591), .B(n30590), .Z(n30729) );
  NANDN U31902 ( .A(n30777), .B(n30592), .Z(n30596) );
  NANDN U31903 ( .A(n30594), .B(n30593), .Z(n30595) );
  AND U31904 ( .A(n30596), .B(n30595), .Z(n30889) );
  AND U31905 ( .A(x[503]), .B(y[7975]), .Z(n30851) );
  AND U31906 ( .A(y[7974]), .B(x[504]), .Z(n30598) );
  AND U31907 ( .A(y[7973]), .B(x[505]), .Z(n30597) );
  XOR U31908 ( .A(n30598), .B(n30597), .Z(n30850) );
  XOR U31909 ( .A(n30851), .B(n30850), .Z(n30891) );
  AND U31910 ( .A(n30599), .B(o[317]), .Z(n30871) );
  AND U31911 ( .A(x[508]), .B(y[7970]), .Z(n30873) );
  AND U31912 ( .A(x[496]), .B(y[7982]), .Z(n30872) );
  XOR U31913 ( .A(n30873), .B(n30872), .Z(n30870) );
  XNOR U31914 ( .A(n30871), .B(n30870), .Z(n30890) );
  XNOR U31915 ( .A(n30889), .B(n30888), .Z(n30728) );
  XOR U31916 ( .A(n30729), .B(n30728), .Z(n30727) );
  XOR U31917 ( .A(n30726), .B(n30727), .Z(n30929) );
  NAND U31918 ( .A(n30600), .B(n30853), .Z(n30604) );
  NAND U31919 ( .A(n30602), .B(n30601), .Z(n30603) );
  NAND U31920 ( .A(n30604), .B(n30603), .Z(n30697) );
  NAND U31921 ( .A(n30606), .B(n30605), .Z(n30610) );
  NAND U31922 ( .A(n30608), .B(n30607), .Z(n30609) );
  AND U31923 ( .A(n30610), .B(n30609), .Z(n30883) );
  AND U31924 ( .A(x[480]), .B(y[7998]), .Z(n30770) );
  AND U31925 ( .A(x[509]), .B(y[7969]), .Z(n30793) );
  XOR U31926 ( .A(o[318]), .B(n30793), .Z(n30772) );
  AND U31927 ( .A(x[510]), .B(y[7968]), .Z(n30771) );
  XOR U31928 ( .A(n30772), .B(n30771), .Z(n30769) );
  XOR U31929 ( .A(n30770), .B(n30769), .Z(n30885) );
  AND U31930 ( .A(x[500]), .B(y[7978]), .Z(n30735) );
  XOR U31931 ( .A(n30735), .B(n30734), .Z(n30733) );
  AND U31932 ( .A(x[488]), .B(y[7990]), .Z(n30732) );
  XNOR U31933 ( .A(n30733), .B(n30732), .Z(n30884) );
  XNOR U31934 ( .A(n30883), .B(n30882), .Z(n30696) );
  XOR U31935 ( .A(n30697), .B(n30696), .Z(n30694) );
  AND U31936 ( .A(x[487]), .B(y[7991]), .Z(n30776) );
  NAND U31937 ( .A(n30611), .B(n30776), .Z(n30615) );
  NAND U31938 ( .A(n30613), .B(n30612), .Z(n30614) );
  AND U31939 ( .A(n30615), .B(n30614), .Z(n30718) );
  AND U31940 ( .A(y[7977]), .B(x[501]), .Z(n30617) );
  AND U31941 ( .A(y[7976]), .B(x[502]), .Z(n30616) );
  XOR U31942 ( .A(n30617), .B(n30616), .Z(n30775) );
  XOR U31943 ( .A(n30776), .B(n30775), .Z(n30721) );
  AND U31944 ( .A(x[497]), .B(y[7981]), .Z(n30744) );
  AND U31945 ( .A(x[482]), .B(y[7996]), .Z(n30746) );
  AND U31946 ( .A(x[506]), .B(y[7972]), .Z(n30745) );
  XOR U31947 ( .A(n30746), .B(n30745), .Z(n30743) );
  XNOR U31948 ( .A(n30744), .B(n30743), .Z(n30720) );
  XNOR U31949 ( .A(n30718), .B(n30719), .Z(n30695) );
  NAND U31950 ( .A(n30619), .B(n30618), .Z(n30623) );
  NAND U31951 ( .A(n30621), .B(n30620), .Z(n30622) );
  NAND U31952 ( .A(n30623), .B(n30622), .Z(n30930) );
  XOR U31953 ( .A(n30931), .B(n30930), .Z(n30928) );
  XOR U31954 ( .A(n30929), .B(n30928), .Z(n30948) );
  XNOR U31955 ( .A(n30946), .B(n30947), .Z(n30961) );
  NANDN U31956 ( .A(n30625), .B(n30624), .Z(n30629) );
  NANDN U31957 ( .A(n30627), .B(n30626), .Z(n30628) );
  NAND U31958 ( .A(n30629), .B(n30628), .Z(n30958) );
  XOR U31959 ( .A(n30961), .B(n30958), .Z(n30630) );
  XOR U31960 ( .A(n30959), .B(n30630), .Z(n30940) );
  NANDN U31961 ( .A(n30632), .B(n30631), .Z(n30636) );
  NANDN U31962 ( .A(n30634), .B(n30633), .Z(n30635) );
  NAND U31963 ( .A(n30636), .B(n30635), .Z(n30942) );
  NANDN U31964 ( .A(n30638), .B(n30637), .Z(n30642) );
  NAND U31965 ( .A(n30640), .B(n30639), .Z(n30641) );
  AND U31966 ( .A(n30642), .B(n30641), .Z(n30923) );
  NAND U31967 ( .A(n30644), .B(n30643), .Z(n30648) );
  NAND U31968 ( .A(n30646), .B(n30645), .Z(n30647) );
  AND U31969 ( .A(n30648), .B(n30647), .Z(n30913) );
  NAND U31970 ( .A(n30650), .B(n30649), .Z(n30654) );
  NANDN U31971 ( .A(n30652), .B(n30651), .Z(n30653) );
  AND U31972 ( .A(n30654), .B(n30653), .Z(n30912) );
  XOR U31973 ( .A(n30913), .B(n30912), .Z(n30911) );
  NANDN U31974 ( .A(n30656), .B(n30655), .Z(n30660) );
  NANDN U31975 ( .A(n30658), .B(n30657), .Z(n30659) );
  NAND U31976 ( .A(n30660), .B(n30659), .Z(n30910) );
  XOR U31977 ( .A(n30911), .B(n30910), .Z(n30925) );
  NAND U31978 ( .A(n30790), .B(n30661), .Z(n30665) );
  NAND U31979 ( .A(n30663), .B(n30662), .Z(n30664) );
  AND U31980 ( .A(n30665), .B(n30664), .Z(n30906) );
  NAND U31981 ( .A(n30667), .B(n30666), .Z(n30671) );
  NAND U31982 ( .A(n30669), .B(n30668), .Z(n30670) );
  NAND U31983 ( .A(n30671), .B(n30670), .Z(n30712) );
  NAND U31984 ( .A(y[7986]), .B(x[492]), .Z(n30672) );
  XNOR U31985 ( .A(n30673), .B(n30672), .Z(n30739) );
  XOR U31986 ( .A(n30739), .B(n30738), .Z(n30789) );
  AND U31987 ( .A(y[7989]), .B(x[489]), .Z(n30675) );
  XOR U31988 ( .A(n30675), .B(n30674), .Z(n30788) );
  XOR U31989 ( .A(n30789), .B(n30788), .Z(n30715) );
  AND U31990 ( .A(x[507]), .B(y[7971]), .Z(n30867) );
  AND U31991 ( .A(x[481]), .B(y[7997]), .Z(n30866) );
  XOR U31992 ( .A(n30867), .B(n30866), .Z(n30865) );
  XOR U31993 ( .A(n30865), .B(n30864), .Z(n30714) );
  XOR U31994 ( .A(n30715), .B(n30714), .Z(n30713) );
  XOR U31995 ( .A(n30712), .B(n30713), .Z(n30907) );
  NAND U31996 ( .A(n30677), .B(n30676), .Z(n30681) );
  NANDN U31997 ( .A(n30679), .B(n30678), .Z(n30680) );
  AND U31998 ( .A(n30681), .B(n30680), .Z(n30904) );
  XNOR U31999 ( .A(n30905), .B(n30904), .Z(n30924) );
  XOR U32000 ( .A(n30923), .B(n30922), .Z(n30943) );
  XNOR U32001 ( .A(n30942), .B(n30943), .Z(n30941) );
  XOR U32002 ( .A(n30683), .B(n30682), .Z(n30966) );
  XNOR U32003 ( .A(n30967), .B(n30966), .Z(N639) );
  NANDN U32004 ( .A(n30683), .B(n30682), .Z(n30687) );
  NANDN U32005 ( .A(n30685), .B(n30684), .Z(n30686) );
  AND U32006 ( .A(n30687), .B(n30686), .Z(n30983) );
  NAND U32007 ( .A(n30689), .B(n30688), .Z(n30693) );
  NANDN U32008 ( .A(n30691), .B(n30690), .Z(n30692) );
  AND U32009 ( .A(n30693), .B(n30692), .Z(n30957) );
  NANDN U32010 ( .A(n30695), .B(n30694), .Z(n30699) );
  NAND U32011 ( .A(n30697), .B(n30696), .Z(n30698) );
  AND U32012 ( .A(n30699), .B(n30698), .Z(n30939) );
  NAND U32013 ( .A(n30701), .B(n30700), .Z(n30705) );
  NAND U32014 ( .A(n30703), .B(n30702), .Z(n30704) );
  AND U32015 ( .A(n30705), .B(n30704), .Z(n30921) );
  NANDN U32016 ( .A(n30707), .B(n30706), .Z(n30711) );
  NANDN U32017 ( .A(n30709), .B(n30708), .Z(n30710) );
  AND U32018 ( .A(n30711), .B(n30710), .Z(n30903) );
  NAND U32019 ( .A(n30713), .B(n30712), .Z(n30717) );
  NAND U32020 ( .A(n30715), .B(n30714), .Z(n30716) );
  AND U32021 ( .A(n30717), .B(n30716), .Z(n30725) );
  NANDN U32022 ( .A(n30719), .B(n30718), .Z(n30723) );
  NANDN U32023 ( .A(n30721), .B(n30720), .Z(n30722) );
  NAND U32024 ( .A(n30723), .B(n30722), .Z(n30724) );
  XNOR U32025 ( .A(n30725), .B(n30724), .Z(n30901) );
  NAND U32026 ( .A(n30727), .B(n30726), .Z(n30731) );
  NAND U32027 ( .A(n30729), .B(n30728), .Z(n30730) );
  AND U32028 ( .A(n30731), .B(n30730), .Z(n30899) );
  NAND U32029 ( .A(n30733), .B(n30732), .Z(n30737) );
  NAND U32030 ( .A(n30735), .B(n30734), .Z(n30736) );
  AND U32031 ( .A(n30737), .B(n30736), .Z(n30768) );
  NAND U32032 ( .A(n30739), .B(n30738), .Z(n30742) );
  NAND U32033 ( .A(n30740), .B(n30813), .Z(n30741) );
  AND U32034 ( .A(n30742), .B(n30741), .Z(n30750) );
  NAND U32035 ( .A(n30744), .B(n30743), .Z(n30748) );
  NAND U32036 ( .A(n30746), .B(n30745), .Z(n30747) );
  NAND U32037 ( .A(n30748), .B(n30747), .Z(n30749) );
  XNOR U32038 ( .A(n30750), .B(n30749), .Z(n30766) );
  AND U32039 ( .A(y[7968]), .B(x[511]), .Z(n30752) );
  NAND U32040 ( .A(y[7995]), .B(x[484]), .Z(n30751) );
  XNOR U32041 ( .A(n30752), .B(n30751), .Z(n30756) );
  AND U32042 ( .A(y[7985]), .B(x[494]), .Z(n30754) );
  NAND U32043 ( .A(y[7990]), .B(x[489]), .Z(n30753) );
  XNOR U32044 ( .A(n30754), .B(n30753), .Z(n30755) );
  XOR U32045 ( .A(n30756), .B(n30755), .Z(n30764) );
  AND U32046 ( .A(y[7994]), .B(x[485]), .Z(n30758) );
  NAND U32047 ( .A(y[7992]), .B(x[487]), .Z(n30757) );
  XNOR U32048 ( .A(n30758), .B(n30757), .Z(n30762) );
  AND U32049 ( .A(y[7993]), .B(x[486]), .Z(n30760) );
  NAND U32050 ( .A(y[7981]), .B(x[498]), .Z(n30759) );
  XNOR U32051 ( .A(n30760), .B(n30759), .Z(n30761) );
  XNOR U32052 ( .A(n30762), .B(n30761), .Z(n30763) );
  XNOR U32053 ( .A(n30764), .B(n30763), .Z(n30765) );
  XNOR U32054 ( .A(n30766), .B(n30765), .Z(n30767) );
  XNOR U32055 ( .A(n30768), .B(n30767), .Z(n30849) );
  NAND U32056 ( .A(n30770), .B(n30769), .Z(n30774) );
  NAND U32057 ( .A(n30772), .B(n30771), .Z(n30773) );
  AND U32058 ( .A(n30774), .B(n30773), .Z(n30847) );
  NAND U32059 ( .A(n30776), .B(n30775), .Z(n30779) );
  AND U32060 ( .A(x[502]), .B(y[7977]), .Z(n30794) );
  NANDN U32061 ( .A(n30777), .B(n30794), .Z(n30778) );
  AND U32062 ( .A(n30779), .B(n30778), .Z(n30787) );
  NAND U32063 ( .A(n30781), .B(n30780), .Z(n30785) );
  NAND U32064 ( .A(n30783), .B(n30782), .Z(n30784) );
  NAND U32065 ( .A(n30785), .B(n30784), .Z(n30786) );
  XNOR U32066 ( .A(n30787), .B(n30786), .Z(n30845) );
  NAND U32067 ( .A(n30789), .B(n30788), .Z(n30792) );
  AND U32068 ( .A(x[490]), .B(y[7989]), .Z(n30812) );
  NAND U32069 ( .A(n30790), .B(n30812), .Z(n30791) );
  AND U32070 ( .A(n30792), .B(n30791), .Z(n30843) );
  AND U32071 ( .A(y[7997]), .B(x[482]), .Z(n30801) );
  AND U32072 ( .A(n30793), .B(o[318]), .Z(n30799) );
  XOR U32073 ( .A(n30794), .B(o[319]), .Z(n30797) );
  AND U32074 ( .A(x[505]), .B(y[7974]), .Z(n30852) );
  XNOR U32075 ( .A(n30795), .B(n30852), .Z(n30796) );
  XNOR U32076 ( .A(n30797), .B(n30796), .Z(n30798) );
  XNOR U32077 ( .A(n30799), .B(n30798), .Z(n30800) );
  XNOR U32078 ( .A(n30801), .B(n30800), .Z(n30841) );
  AND U32079 ( .A(y[7978]), .B(x[501]), .Z(n30803) );
  NAND U32080 ( .A(y[7991]), .B(x[488]), .Z(n30802) );
  XNOR U32081 ( .A(n30803), .B(n30802), .Z(n30811) );
  AND U32082 ( .A(y[7980]), .B(x[499]), .Z(n30809) );
  AND U32083 ( .A(y[7988]), .B(x[491]), .Z(n30805) );
  NAND U32084 ( .A(y[7987]), .B(x[492]), .Z(n30804) );
  XNOR U32085 ( .A(n30805), .B(n30804), .Z(n30806) );
  XNOR U32086 ( .A(n30807), .B(n30806), .Z(n30808) );
  XNOR U32087 ( .A(n30809), .B(n30808), .Z(n30810) );
  XOR U32088 ( .A(n30811), .B(n30810), .Z(n30815) );
  XNOR U32089 ( .A(n30813), .B(n30812), .Z(n30814) );
  XNOR U32090 ( .A(n30815), .B(n30814), .Z(n30831) );
  AND U32091 ( .A(y[7969]), .B(x[510]), .Z(n30817) );
  NAND U32092 ( .A(y[7970]), .B(x[509]), .Z(n30816) );
  XNOR U32093 ( .A(n30817), .B(n30816), .Z(n30821) );
  AND U32094 ( .A(y[7983]), .B(x[496]), .Z(n30819) );
  NAND U32095 ( .A(y[7979]), .B(x[500]), .Z(n30818) );
  XNOR U32096 ( .A(n30819), .B(n30818), .Z(n30820) );
  XOR U32097 ( .A(n30821), .B(n30820), .Z(n30829) );
  AND U32098 ( .A(y[7973]), .B(x[506]), .Z(n30823) );
  NAND U32099 ( .A(y[7971]), .B(x[508]), .Z(n30822) );
  XNOR U32100 ( .A(n30823), .B(n30822), .Z(n30827) );
  AND U32101 ( .A(y[7998]), .B(x[481]), .Z(n30825) );
  NAND U32102 ( .A(y[7999]), .B(x[480]), .Z(n30824) );
  XNOR U32103 ( .A(n30825), .B(n30824), .Z(n30826) );
  XNOR U32104 ( .A(n30827), .B(n30826), .Z(n30828) );
  XNOR U32105 ( .A(n30829), .B(n30828), .Z(n30830) );
  XOR U32106 ( .A(n30831), .B(n30830), .Z(n30839) );
  AND U32107 ( .A(y[7972]), .B(x[507]), .Z(n30833) );
  NAND U32108 ( .A(y[7982]), .B(x[497]), .Z(n30832) );
  XNOR U32109 ( .A(n30833), .B(n30832), .Z(n30837) );
  AND U32110 ( .A(y[7976]), .B(x[503]), .Z(n30835) );
  NAND U32111 ( .A(y[7996]), .B(x[483]), .Z(n30834) );
  XNOR U32112 ( .A(n30835), .B(n30834), .Z(n30836) );
  XNOR U32113 ( .A(n30837), .B(n30836), .Z(n30838) );
  XNOR U32114 ( .A(n30839), .B(n30838), .Z(n30840) );
  XNOR U32115 ( .A(n30841), .B(n30840), .Z(n30842) );
  XNOR U32116 ( .A(n30843), .B(n30842), .Z(n30844) );
  XNOR U32117 ( .A(n30845), .B(n30844), .Z(n30846) );
  XNOR U32118 ( .A(n30847), .B(n30846), .Z(n30848) );
  XOR U32119 ( .A(n30849), .B(n30848), .Z(n30881) );
  NAND U32120 ( .A(n30851), .B(n30850), .Z(n30855) );
  NAND U32121 ( .A(n30853), .B(n30852), .Z(n30854) );
  AND U32122 ( .A(n30855), .B(n30854), .Z(n30863) );
  NAND U32123 ( .A(n30857), .B(n30856), .Z(n30861) );
  NAND U32124 ( .A(n30859), .B(n30858), .Z(n30860) );
  NAND U32125 ( .A(n30861), .B(n30860), .Z(n30862) );
  XNOR U32126 ( .A(n30863), .B(n30862), .Z(n30879) );
  NAND U32127 ( .A(n30865), .B(n30864), .Z(n30869) );
  NAND U32128 ( .A(n30867), .B(n30866), .Z(n30868) );
  AND U32129 ( .A(n30869), .B(n30868), .Z(n30877) );
  NAND U32130 ( .A(n30871), .B(n30870), .Z(n30875) );
  NAND U32131 ( .A(n30873), .B(n30872), .Z(n30874) );
  NAND U32132 ( .A(n30875), .B(n30874), .Z(n30876) );
  XNOR U32133 ( .A(n30877), .B(n30876), .Z(n30878) );
  XNOR U32134 ( .A(n30879), .B(n30878), .Z(n30880) );
  XNOR U32135 ( .A(n30881), .B(n30880), .Z(n30897) );
  NAND U32136 ( .A(n30883), .B(n30882), .Z(n30887) );
  NANDN U32137 ( .A(n30885), .B(n30884), .Z(n30886) );
  AND U32138 ( .A(n30887), .B(n30886), .Z(n30895) );
  NAND U32139 ( .A(n30889), .B(n30888), .Z(n30893) );
  NANDN U32140 ( .A(n30891), .B(n30890), .Z(n30892) );
  NAND U32141 ( .A(n30893), .B(n30892), .Z(n30894) );
  XNOR U32142 ( .A(n30895), .B(n30894), .Z(n30896) );
  XNOR U32143 ( .A(n30897), .B(n30896), .Z(n30898) );
  XNOR U32144 ( .A(n30899), .B(n30898), .Z(n30900) );
  XNOR U32145 ( .A(n30901), .B(n30900), .Z(n30902) );
  XNOR U32146 ( .A(n30903), .B(n30902), .Z(n30919) );
  NAND U32147 ( .A(n30905), .B(n30904), .Z(n30909) );
  NANDN U32148 ( .A(n30907), .B(n30906), .Z(n30908) );
  AND U32149 ( .A(n30909), .B(n30908), .Z(n30917) );
  NAND U32150 ( .A(n30911), .B(n30910), .Z(n30915) );
  NAND U32151 ( .A(n30913), .B(n30912), .Z(n30914) );
  NAND U32152 ( .A(n30915), .B(n30914), .Z(n30916) );
  XNOR U32153 ( .A(n30917), .B(n30916), .Z(n30918) );
  XNOR U32154 ( .A(n30919), .B(n30918), .Z(n30920) );
  XNOR U32155 ( .A(n30921), .B(n30920), .Z(n30937) );
  NAND U32156 ( .A(n30923), .B(n30922), .Z(n30927) );
  NANDN U32157 ( .A(n30925), .B(n30924), .Z(n30926) );
  AND U32158 ( .A(n30927), .B(n30926), .Z(n30935) );
  NAND U32159 ( .A(n30929), .B(n30928), .Z(n30933) );
  NAND U32160 ( .A(n30931), .B(n30930), .Z(n30932) );
  NAND U32161 ( .A(n30933), .B(n30932), .Z(n30934) );
  XNOR U32162 ( .A(n30935), .B(n30934), .Z(n30936) );
  XNOR U32163 ( .A(n30937), .B(n30936), .Z(n30938) );
  XNOR U32164 ( .A(n30939), .B(n30938), .Z(n30955) );
  NANDN U32165 ( .A(n30941), .B(n30940), .Z(n30945) );
  NAND U32166 ( .A(n30943), .B(n30942), .Z(n30944) );
  AND U32167 ( .A(n30945), .B(n30944), .Z(n30953) );
  NANDN U32168 ( .A(n30947), .B(n30946), .Z(n30951) );
  NANDN U32169 ( .A(n30949), .B(n30948), .Z(n30950) );
  NAND U32170 ( .A(n30951), .B(n30950), .Z(n30952) );
  XNOR U32171 ( .A(n30953), .B(n30952), .Z(n30954) );
  XNOR U32172 ( .A(n30955), .B(n30954), .Z(n30956) );
  XNOR U32173 ( .A(n30957), .B(n30956), .Z(n30965) );
  OR U32174 ( .A(n30958), .B(n30959), .Z(n30963) );
  AND U32175 ( .A(n30959), .B(n30958), .Z(n30960) );
  OR U32176 ( .A(n30961), .B(n30960), .Z(n30962) );
  NAND U32177 ( .A(n30963), .B(n30962), .Z(n30964) );
  XNOR U32178 ( .A(n30965), .B(n30964), .Z(n30981) );
  NAND U32179 ( .A(n30967), .B(n30966), .Z(n30971) );
  NANDN U32180 ( .A(n30969), .B(n30968), .Z(n30970) );
  AND U32181 ( .A(n30971), .B(n30970), .Z(n30979) );
  NAND U32182 ( .A(n30973), .B(n30972), .Z(n30977) );
  NAND U32183 ( .A(n30975), .B(n30974), .Z(n30976) );
  NAND U32184 ( .A(n30977), .B(n30976), .Z(n30978) );
  XNOR U32185 ( .A(n30979), .B(n30978), .Z(n30980) );
  XNOR U32186 ( .A(n30981), .B(n30980), .Z(n30982) );
  XNOR U32187 ( .A(n30983), .B(n30982), .Z(N640) );
  AND U32188 ( .A(x[480]), .B(y[8000]), .Z(n31603) );
  XOR U32189 ( .A(n31603), .B(o[320]), .Z(N673) );
  NAND U32190 ( .A(x[481]), .B(y[8000]), .Z(n30993) );
  AND U32191 ( .A(x[480]), .B(y[8001]), .Z(n30989) );
  XNOR U32192 ( .A(n30989), .B(o[321]), .Z(n30984) );
  XOR U32193 ( .A(n30993), .B(n30984), .Z(n30986) );
  NAND U32194 ( .A(n31603), .B(o[320]), .Z(n30985) );
  XNOR U32195 ( .A(n30986), .B(n30985), .Z(N674) );
  AND U32196 ( .A(x[480]), .B(y[8002]), .Z(n30992) );
  XNOR U32197 ( .A(n30992), .B(o[322]), .Z(n30998) );
  XNOR U32198 ( .A(n30999), .B(n30998), .Z(n31001) );
  AND U32199 ( .A(y[8000]), .B(x[482]), .Z(n30988) );
  NAND U32200 ( .A(y[8001]), .B(x[481]), .Z(n30987) );
  XNOR U32201 ( .A(n30988), .B(n30987), .Z(n30995) );
  AND U32202 ( .A(n30989), .B(o[321]), .Z(n30994) );
  XNOR U32203 ( .A(n30995), .B(n30994), .Z(n31000) );
  XNOR U32204 ( .A(n31001), .B(n31000), .Z(N675) );
  AND U32205 ( .A(x[481]), .B(y[8002]), .Z(n31120) );
  AND U32206 ( .A(x[482]), .B(y[8001]), .Z(n31009) );
  XOR U32207 ( .A(o[323]), .B(n31009), .Z(n31016) );
  XOR U32208 ( .A(n31120), .B(n31016), .Z(n31018) );
  AND U32209 ( .A(y[8000]), .B(x[483]), .Z(n30991) );
  NAND U32210 ( .A(y[8003]), .B(x[480]), .Z(n30990) );
  XNOR U32211 ( .A(n30991), .B(n30990), .Z(n31005) );
  AND U32212 ( .A(n30992), .B(o[322]), .Z(n31006) );
  XOR U32213 ( .A(n31005), .B(n31006), .Z(n31017) );
  XNOR U32214 ( .A(n31018), .B(n31017), .Z(n31015) );
  NANDN U32215 ( .A(n30993), .B(n31009), .Z(n30997) );
  NAND U32216 ( .A(n30995), .B(n30994), .Z(n30996) );
  NAND U32217 ( .A(n30997), .B(n30996), .Z(n31013) );
  NANDN U32218 ( .A(n30999), .B(n30998), .Z(n31003) );
  NAND U32219 ( .A(n31001), .B(n31000), .Z(n31002) );
  AND U32220 ( .A(n31003), .B(n31002), .Z(n31014) );
  XOR U32221 ( .A(n31013), .B(n31014), .Z(n31004) );
  XNOR U32222 ( .A(n31015), .B(n31004), .Z(N676) );
  AND U32223 ( .A(x[483]), .B(y[8003]), .Z(n31077) );
  NAND U32224 ( .A(n31603), .B(n31077), .Z(n31008) );
  NAND U32225 ( .A(n31006), .B(n31005), .Z(n31007) );
  AND U32226 ( .A(n31008), .B(n31007), .Z(n31045) );
  AND U32227 ( .A(o[323]), .B(n31009), .Z(n31032) );
  AND U32228 ( .A(x[480]), .B(y[8004]), .Z(n31011) );
  AND U32229 ( .A(y[8000]), .B(x[484]), .Z(n31010) );
  XOR U32230 ( .A(n31011), .B(n31010), .Z(n31031) );
  XOR U32231 ( .A(n31032), .B(n31031), .Z(n31043) );
  AND U32232 ( .A(y[8002]), .B(x[482]), .Z(n31157) );
  NAND U32233 ( .A(y[8003]), .B(x[481]), .Z(n31012) );
  XNOR U32234 ( .A(n31157), .B(n31012), .Z(n31028) );
  AND U32235 ( .A(x[483]), .B(y[8001]), .Z(n31026) );
  XOR U32236 ( .A(n31026), .B(o[324]), .Z(n31027) );
  XOR U32237 ( .A(n31028), .B(n31027), .Z(n31042) );
  XOR U32238 ( .A(n31043), .B(n31042), .Z(n31044) );
  XOR U32239 ( .A(n31045), .B(n31044), .Z(n31038) );
  NAND U32240 ( .A(n31120), .B(n31016), .Z(n31020) );
  NAND U32241 ( .A(n31018), .B(n31017), .Z(n31019) );
  NAND U32242 ( .A(n31020), .B(n31019), .Z(n31036) );
  IV U32243 ( .A(n31036), .Z(n31035) );
  XOR U32244 ( .A(n31037), .B(n31035), .Z(n31021) );
  XNOR U32245 ( .A(n31038), .B(n31021), .Z(N677) );
  AND U32246 ( .A(x[482]), .B(y[8003]), .Z(n31129) );
  AND U32247 ( .A(y[8002]), .B(x[483]), .Z(n31023) );
  NAND U32248 ( .A(y[8004]), .B(x[481]), .Z(n31022) );
  XNOR U32249 ( .A(n31023), .B(n31022), .Z(n31063) );
  NAND U32250 ( .A(x[484]), .B(y[8001]), .Z(n31075) );
  XOR U32251 ( .A(n31063), .B(n31062), .Z(n31066) );
  XOR U32252 ( .A(n31129), .B(n31066), .Z(n31068) );
  AND U32253 ( .A(y[8000]), .B(x[485]), .Z(n31025) );
  NAND U32254 ( .A(y[8005]), .B(x[480]), .Z(n31024) );
  XNOR U32255 ( .A(n31025), .B(n31024), .Z(n31070) );
  AND U32256 ( .A(n31026), .B(o[324]), .Z(n31069) );
  XOR U32257 ( .A(n31070), .B(n31069), .Z(n31067) );
  XOR U32258 ( .A(n31068), .B(n31067), .Z(n31058) );
  NAND U32259 ( .A(n31129), .B(n31120), .Z(n31030) );
  NAND U32260 ( .A(n31028), .B(n31027), .Z(n31029) );
  NAND U32261 ( .A(n31030), .B(n31029), .Z(n31057) );
  AND U32262 ( .A(x[484]), .B(y[8004]), .Z(n31811) );
  NAND U32263 ( .A(n31811), .B(n31603), .Z(n31034) );
  NAND U32264 ( .A(n31032), .B(n31031), .Z(n31033) );
  NAND U32265 ( .A(n31034), .B(n31033), .Z(n31056) );
  XNOR U32266 ( .A(n31057), .B(n31056), .Z(n31059) );
  OR U32267 ( .A(n31037), .B(n31035), .Z(n31041) );
  ANDN U32268 ( .B(n31037), .A(n31036), .Z(n31039) );
  OR U32269 ( .A(n31039), .B(n31038), .Z(n31040) );
  AND U32270 ( .A(n31041), .B(n31040), .Z(n31050) );
  NAND U32271 ( .A(n31043), .B(n31042), .Z(n31047) );
  NANDN U32272 ( .A(n31045), .B(n31044), .Z(n31046) );
  AND U32273 ( .A(n31047), .B(n31046), .Z(n31051) );
  IV U32274 ( .A(n31051), .Z(n31049) );
  XOR U32275 ( .A(n31050), .B(n31049), .Z(n31048) );
  XNOR U32276 ( .A(n31052), .B(n31048), .Z(N678) );
  NANDN U32277 ( .A(n31049), .B(n31050), .Z(n31055) );
  NOR U32278 ( .A(n31051), .B(n31050), .Z(n31053) );
  OR U32279 ( .A(n31053), .B(n31052), .Z(n31054) );
  AND U32280 ( .A(n31055), .B(n31054), .Z(n31104) );
  NAND U32281 ( .A(n31057), .B(n31056), .Z(n31061) );
  NANDN U32282 ( .A(n31059), .B(n31058), .Z(n31060) );
  AND U32283 ( .A(n31061), .B(n31060), .Z(n31103) );
  XNOR U32284 ( .A(n31104), .B(n31103), .Z(n31106) );
  AND U32285 ( .A(x[483]), .B(y[8004]), .Z(n31130) );
  NAND U32286 ( .A(n31130), .B(n31120), .Z(n31065) );
  NAND U32287 ( .A(n31063), .B(n31062), .Z(n31064) );
  NAND U32288 ( .A(n31065), .B(n31064), .Z(n31109) );
  XOR U32289 ( .A(n31109), .B(n31110), .Z(n31112) );
  AND U32290 ( .A(x[485]), .B(y[8005]), .Z(n31304) );
  NAND U32291 ( .A(n31603), .B(n31304), .Z(n31072) );
  NAND U32292 ( .A(n31070), .B(n31069), .Z(n31071) );
  AND U32293 ( .A(n31072), .B(n31071), .Z(n31080) );
  AND U32294 ( .A(y[8000]), .B(x[486]), .Z(n31074) );
  NAND U32295 ( .A(y[8006]), .B(x[480]), .Z(n31073) );
  XNOR U32296 ( .A(n31074), .B(n31073), .Z(n31087) );
  ANDN U32297 ( .B(o[325]), .A(n31075), .Z(n31086) );
  XOR U32298 ( .A(n31087), .B(n31086), .Z(n31079) );
  NAND U32299 ( .A(y[8004]), .B(x[482]), .Z(n31076) );
  XNOR U32300 ( .A(n31077), .B(n31076), .Z(n31091) );
  AND U32301 ( .A(x[481]), .B(y[8005]), .Z(n31325) );
  NAND U32302 ( .A(y[8002]), .B(x[484]), .Z(n31078) );
  XNOR U32303 ( .A(n31325), .B(n31078), .Z(n31095) );
  NAND U32304 ( .A(x[485]), .B(y[8001]), .Z(n31102) );
  XOR U32305 ( .A(n31095), .B(n31094), .Z(n31090) );
  XOR U32306 ( .A(n31091), .B(n31090), .Z(n31081) );
  XOR U32307 ( .A(n31082), .B(n31081), .Z(n31111) );
  XNOR U32308 ( .A(n31112), .B(n31111), .Z(n31105) );
  XNOR U32309 ( .A(n31106), .B(n31105), .Z(N679) );
  NANDN U32310 ( .A(n31080), .B(n31079), .Z(n31084) );
  NAND U32311 ( .A(n31082), .B(n31081), .Z(n31083) );
  AND U32312 ( .A(n31084), .B(n31083), .Z(n31149) );
  AND U32313 ( .A(y[8002]), .B(x[485]), .Z(n31207) );
  NAND U32314 ( .A(y[8006]), .B(x[481]), .Z(n31085) );
  XNOR U32315 ( .A(n31207), .B(n31085), .Z(n31122) );
  AND U32316 ( .A(x[486]), .B(y[8001]), .Z(n31126) );
  XOR U32317 ( .A(o[327]), .B(n31126), .Z(n31121) );
  XOR U32318 ( .A(n31122), .B(n31121), .Z(n31141) );
  AND U32319 ( .A(x[486]), .B(y[8006]), .Z(n31346) );
  NAND U32320 ( .A(n31603), .B(n31346), .Z(n31089) );
  NAND U32321 ( .A(n31087), .B(n31086), .Z(n31088) );
  AND U32322 ( .A(n31089), .B(n31088), .Z(n31140) );
  NAND U32323 ( .A(n31129), .B(n31130), .Z(n31093) );
  NAND U32324 ( .A(n31091), .B(n31090), .Z(n31092) );
  AND U32325 ( .A(n31093), .B(n31092), .Z(n31142) );
  XOR U32326 ( .A(n31143), .B(n31142), .Z(n31147) );
  AND U32327 ( .A(x[484]), .B(y[8005]), .Z(n31608) );
  NAND U32328 ( .A(n31608), .B(n31120), .Z(n31097) );
  NAND U32329 ( .A(n31095), .B(n31094), .Z(n31096) );
  AND U32330 ( .A(n31097), .B(n31096), .Z(n31117) );
  AND U32331 ( .A(y[8005]), .B(x[482]), .Z(n31099) );
  NAND U32332 ( .A(y[8003]), .B(x[484]), .Z(n31098) );
  XNOR U32333 ( .A(n31099), .B(n31098), .Z(n31131) );
  XOR U32334 ( .A(n31131), .B(n31130), .Z(n31115) );
  AND U32335 ( .A(y[8000]), .B(x[487]), .Z(n31101) );
  NAND U32336 ( .A(y[8007]), .B(x[480]), .Z(n31100) );
  XNOR U32337 ( .A(n31101), .B(n31100), .Z(n31135) );
  ANDN U32338 ( .B(o[326]), .A(n31102), .Z(n31134) );
  XNOR U32339 ( .A(n31135), .B(n31134), .Z(n31114) );
  XOR U32340 ( .A(n31117), .B(n31116), .Z(n31146) );
  XOR U32341 ( .A(n31147), .B(n31146), .Z(n31148) );
  XNOR U32342 ( .A(n31149), .B(n31148), .Z(n31155) );
  NANDN U32343 ( .A(n31104), .B(n31103), .Z(n31108) );
  NAND U32344 ( .A(n31106), .B(n31105), .Z(n31107) );
  NAND U32345 ( .A(n31108), .B(n31107), .Z(n31153) );
  IV U32346 ( .A(n31154), .Z(n31152) );
  XOR U32347 ( .A(n31153), .B(n31152), .Z(n31113) );
  XNOR U32348 ( .A(n31155), .B(n31113), .Z(N680) );
  NANDN U32349 ( .A(n31115), .B(n31114), .Z(n31119) );
  NAND U32350 ( .A(n31117), .B(n31116), .Z(n31118) );
  AND U32351 ( .A(n31119), .B(n31118), .Z(n31188) );
  AND U32352 ( .A(x[485]), .B(y[8006]), .Z(n31296) );
  NAND U32353 ( .A(n31296), .B(n31120), .Z(n31124) );
  NAND U32354 ( .A(n31122), .B(n31121), .Z(n31123) );
  AND U32355 ( .A(n31124), .B(n31123), .Z(n31186) );
  AND U32356 ( .A(y[8003]), .B(x[485]), .Z(n31717) );
  NAND U32357 ( .A(y[8007]), .B(x[481]), .Z(n31125) );
  XNOR U32358 ( .A(n31717), .B(n31125), .Z(n31176) );
  AND U32359 ( .A(o[327]), .B(n31126), .Z(n31175) );
  XOR U32360 ( .A(n31176), .B(n31175), .Z(n31163) );
  NAND U32361 ( .A(x[483]), .B(y[8005]), .Z(n31947) );
  AND U32362 ( .A(y[8002]), .B(x[486]), .Z(n31128) );
  NAND U32363 ( .A(y[8006]), .B(x[482]), .Z(n31127) );
  XNOR U32364 ( .A(n31128), .B(n31127), .Z(n31158) );
  XNOR U32365 ( .A(n31811), .B(n31158), .Z(n31161) );
  XOR U32366 ( .A(n31947), .B(n31161), .Z(n31162) );
  XOR U32367 ( .A(n31163), .B(n31162), .Z(n31185) );
  XNOR U32368 ( .A(n31188), .B(n31187), .Z(n31196) );
  NAND U32369 ( .A(n31608), .B(n31129), .Z(n31133) );
  NAND U32370 ( .A(n31131), .B(n31130), .Z(n31132) );
  AND U32371 ( .A(n31133), .B(n31132), .Z(n31182) );
  AND U32372 ( .A(x[487]), .B(y[8007]), .Z(n31495) );
  NAND U32373 ( .A(n31603), .B(n31495), .Z(n31137) );
  NAND U32374 ( .A(n31135), .B(n31134), .Z(n31136) );
  AND U32375 ( .A(n31137), .B(n31136), .Z(n31180) );
  AND U32376 ( .A(y[8000]), .B(x[488]), .Z(n31139) );
  NAND U32377 ( .A(y[8008]), .B(x[480]), .Z(n31138) );
  XNOR U32378 ( .A(n31139), .B(n31138), .Z(n31166) );
  AND U32379 ( .A(x[487]), .B(y[8001]), .Z(n31171) );
  XOR U32380 ( .A(o[328]), .B(n31171), .Z(n31165) );
  XOR U32381 ( .A(n31166), .B(n31165), .Z(n31179) );
  NANDN U32382 ( .A(n31141), .B(n31140), .Z(n31145) );
  NAND U32383 ( .A(n31143), .B(n31142), .Z(n31144) );
  NAND U32384 ( .A(n31145), .B(n31144), .Z(n31194) );
  XOR U32385 ( .A(n31196), .B(n31197), .Z(n31193) );
  NAND U32386 ( .A(n31147), .B(n31146), .Z(n31151) );
  NAND U32387 ( .A(n31149), .B(n31148), .Z(n31150) );
  NAND U32388 ( .A(n31151), .B(n31150), .Z(n31191) );
  XOR U32389 ( .A(n31191), .B(n31192), .Z(n31156) );
  XNOR U32390 ( .A(n31193), .B(n31156), .Z(N681) );
  NAND U32391 ( .A(n31346), .B(n31157), .Z(n31160) );
  NAND U32392 ( .A(n31811), .B(n31158), .Z(n31159) );
  NAND U32393 ( .A(n31160), .B(n31159), .Z(n31202) );
  XOR U32394 ( .A(n31202), .B(n31201), .Z(n31204) );
  AND U32395 ( .A(x[488]), .B(y[8008]), .Z(n31164) );
  NAND U32396 ( .A(n31164), .B(n31603), .Z(n31168) );
  NAND U32397 ( .A(n31166), .B(n31165), .Z(n31167) );
  AND U32398 ( .A(n31168), .B(n31167), .Z(n31236) );
  AND U32399 ( .A(y[8004]), .B(x[485]), .Z(n31170) );
  NAND U32400 ( .A(y[8002]), .B(x[487]), .Z(n31169) );
  XNOR U32401 ( .A(n31170), .B(n31169), .Z(n31209) );
  AND U32402 ( .A(o[328]), .B(n31171), .Z(n31208) );
  XNOR U32403 ( .A(n31209), .B(n31208), .Z(n31234) );
  AND U32404 ( .A(y[8000]), .B(x[489]), .Z(n31173) );
  NAND U32405 ( .A(y[8009]), .B(x[480]), .Z(n31172) );
  XNOR U32406 ( .A(n31173), .B(n31172), .Z(n31216) );
  NAND U32407 ( .A(x[488]), .B(y[8001]), .Z(n31223) );
  XNOR U32408 ( .A(n31216), .B(n31215), .Z(n31233) );
  XOR U32409 ( .A(n31234), .B(n31233), .Z(n31235) );
  XNOR U32410 ( .A(n31236), .B(n31235), .Z(n31230) );
  AND U32411 ( .A(y[8003]), .B(x[486]), .Z(n31556) );
  NAND U32412 ( .A(y[8008]), .B(x[481]), .Z(n31174) );
  XNOR U32413 ( .A(n31556), .B(n31174), .Z(n31220) );
  XNOR U32414 ( .A(n31608), .B(n31220), .Z(n31240) );
  NAND U32415 ( .A(x[482]), .B(y[8007]), .Z(n31858) );
  AND U32416 ( .A(x[483]), .B(y[8006]), .Z(n31563) );
  XNOR U32417 ( .A(n31858), .B(n31563), .Z(n31239) );
  XNOR U32418 ( .A(n31240), .B(n31239), .Z(n31228) );
  NAND U32419 ( .A(x[485]), .B(y[8007]), .Z(n31412) );
  AND U32420 ( .A(x[481]), .B(y[8003]), .Z(n31219) );
  NANDN U32421 ( .A(n31412), .B(n31219), .Z(n31178) );
  NAND U32422 ( .A(n31176), .B(n31175), .Z(n31177) );
  NAND U32423 ( .A(n31178), .B(n31177), .Z(n31227) );
  XOR U32424 ( .A(n31228), .B(n31227), .Z(n31229) );
  XOR U32425 ( .A(n31230), .B(n31229), .Z(n31203) );
  XOR U32426 ( .A(n31204), .B(n31203), .Z(n31246) );
  NANDN U32427 ( .A(n31180), .B(n31179), .Z(n31184) );
  NANDN U32428 ( .A(n31182), .B(n31181), .Z(n31183) );
  AND U32429 ( .A(n31184), .B(n31183), .Z(n31244) );
  NANDN U32430 ( .A(n31186), .B(n31185), .Z(n31190) );
  NAND U32431 ( .A(n31188), .B(n31187), .Z(n31189) );
  NAND U32432 ( .A(n31190), .B(n31189), .Z(n31243) );
  XNOR U32433 ( .A(n31246), .B(n31245), .Z(n31251) );
  NANDN U32434 ( .A(n31195), .B(n31194), .Z(n31199) );
  NANDN U32435 ( .A(n31197), .B(n31196), .Z(n31198) );
  AND U32436 ( .A(n31199), .B(n31198), .Z(n31249) );
  XOR U32437 ( .A(n31250), .B(n31249), .Z(n31200) );
  XNOR U32438 ( .A(n31251), .B(n31200), .Z(N682) );
  NAND U32439 ( .A(n31202), .B(n31201), .Z(n31206) );
  NAND U32440 ( .A(n31204), .B(n31203), .Z(n31205) );
  AND U32441 ( .A(n31206), .B(n31205), .Z(n31256) );
  AND U32442 ( .A(x[487]), .B(y[8004]), .Z(n31298) );
  NAND U32443 ( .A(n31298), .B(n31207), .Z(n31211) );
  NAND U32444 ( .A(n31209), .B(n31208), .Z(n31210) );
  AND U32445 ( .A(n31211), .B(n31210), .Z(n31311) );
  AND U32446 ( .A(y[8003]), .B(x[487]), .Z(n31213) );
  NAND U32447 ( .A(y[8006]), .B(x[484]), .Z(n31212) );
  XNOR U32448 ( .A(n31213), .B(n31212), .Z(n31282) );
  AND U32449 ( .A(x[486]), .B(y[8004]), .Z(n31281) );
  XOR U32450 ( .A(n31282), .B(n31281), .Z(n31309) );
  AND U32451 ( .A(x[488]), .B(y[8002]), .Z(n31475) );
  AND U32452 ( .A(x[489]), .B(y[8001]), .Z(n31292) );
  XOR U32453 ( .A(n31292), .B(o[330]), .Z(n31303) );
  XOR U32454 ( .A(n31475), .B(n31303), .Z(n31305) );
  XNOR U32455 ( .A(n31305), .B(n31304), .Z(n31308) );
  XNOR U32456 ( .A(n31311), .B(n31310), .Z(n31271) );
  AND U32457 ( .A(x[489]), .B(y[8009]), .Z(n31214) );
  NAND U32458 ( .A(n31214), .B(n31603), .Z(n31218) );
  NAND U32459 ( .A(n31216), .B(n31215), .Z(n31217) );
  NAND U32460 ( .A(n31218), .B(n31217), .Z(n31269) );
  AND U32461 ( .A(x[486]), .B(y[8008]), .Z(n31501) );
  NAND U32462 ( .A(n31501), .B(n31219), .Z(n31222) );
  NAND U32463 ( .A(n31608), .B(n31220), .Z(n31221) );
  NAND U32464 ( .A(n31222), .B(n31221), .Z(n31276) );
  ANDN U32465 ( .B(o[329]), .A(n31223), .Z(n31287) );
  AND U32466 ( .A(y[8000]), .B(x[490]), .Z(n31225) );
  AND U32467 ( .A(y[8010]), .B(x[480]), .Z(n31224) );
  XOR U32468 ( .A(n31225), .B(n31224), .Z(n31286) );
  XOR U32469 ( .A(n31287), .B(n31286), .Z(n31275) );
  AND U32470 ( .A(y[8007]), .B(x[483]), .Z(n32171) );
  NAND U32471 ( .A(y[8009]), .B(x[481]), .Z(n31226) );
  XNOR U32472 ( .A(n32171), .B(n31226), .Z(n31300) );
  AND U32473 ( .A(x[482]), .B(y[8008]), .Z(n31299) );
  XOR U32474 ( .A(n31300), .B(n31299), .Z(n31274) );
  XOR U32475 ( .A(n31275), .B(n31274), .Z(n31277) );
  XOR U32476 ( .A(n31276), .B(n31277), .Z(n31268) );
  XOR U32477 ( .A(n31269), .B(n31268), .Z(n31270) );
  XNOR U32478 ( .A(n31271), .B(n31270), .Z(n31254) );
  NAND U32479 ( .A(n31228), .B(n31227), .Z(n31232) );
  NAND U32480 ( .A(n31230), .B(n31229), .Z(n31231) );
  AND U32481 ( .A(n31232), .B(n31231), .Z(n31265) );
  NAND U32482 ( .A(n31234), .B(n31233), .Z(n31238) );
  NAND U32483 ( .A(n31236), .B(n31235), .Z(n31237) );
  AND U32484 ( .A(n31238), .B(n31237), .Z(n31262) );
  NAND U32485 ( .A(n31240), .B(n31239), .Z(n31242) );
  ANDN U32486 ( .B(n31858), .A(n31563), .Z(n31241) );
  ANDN U32487 ( .B(n31242), .A(n31241), .Z(n31263) );
  XOR U32488 ( .A(n31262), .B(n31263), .Z(n31264) );
  XOR U32489 ( .A(n31265), .B(n31264), .Z(n31253) );
  XOR U32490 ( .A(n31254), .B(n31253), .Z(n31255) );
  XOR U32491 ( .A(n31256), .B(n31255), .Z(n31261) );
  NANDN U32492 ( .A(n31244), .B(n31243), .Z(n31248) );
  NAND U32493 ( .A(n31246), .B(n31245), .Z(n31247) );
  NAND U32494 ( .A(n31248), .B(n31247), .Z(n31259) );
  XOR U32495 ( .A(n31259), .B(n31260), .Z(n31252) );
  XNOR U32496 ( .A(n31261), .B(n31252), .Z(N683) );
  NAND U32497 ( .A(n31254), .B(n31253), .Z(n31258) );
  NAND U32498 ( .A(n31256), .B(n31255), .Z(n31257) );
  NAND U32499 ( .A(n31258), .B(n31257), .Z(n31378) );
  IV U32500 ( .A(n31378), .Z(n31376) );
  NAND U32501 ( .A(n31263), .B(n31262), .Z(n31267) );
  NANDN U32502 ( .A(n31265), .B(n31264), .Z(n31266) );
  NAND U32503 ( .A(n31267), .B(n31266), .Z(n31373) );
  NAND U32504 ( .A(n31269), .B(n31268), .Z(n31273) );
  NAND U32505 ( .A(n31271), .B(n31270), .Z(n31272) );
  NAND U32506 ( .A(n31273), .B(n31272), .Z(n31371) );
  NAND U32507 ( .A(n31275), .B(n31274), .Z(n31279) );
  NAND U32508 ( .A(n31277), .B(n31276), .Z(n31278) );
  NAND U32509 ( .A(n31279), .B(n31278), .Z(n31366) );
  AND U32510 ( .A(x[487]), .B(y[8006]), .Z(n31408) );
  AND U32511 ( .A(x[484]), .B(y[8003]), .Z(n31280) );
  NAND U32512 ( .A(n31408), .B(n31280), .Z(n31284) );
  NAND U32513 ( .A(n31282), .B(n31281), .Z(n31283) );
  NAND U32514 ( .A(n31284), .B(n31283), .Z(n31364) );
  AND U32515 ( .A(x[490]), .B(y[8010]), .Z(n31285) );
  NAND U32516 ( .A(n31285), .B(n31603), .Z(n31289) );
  NAND U32517 ( .A(n31287), .B(n31286), .Z(n31288) );
  NAND U32518 ( .A(n31289), .B(n31288), .Z(n31360) );
  AND U32519 ( .A(y[8000]), .B(x[491]), .Z(n31291) );
  NAND U32520 ( .A(y[8011]), .B(x[480]), .Z(n31290) );
  XNOR U32521 ( .A(n31291), .B(n31290), .Z(n31336) );
  AND U32522 ( .A(n31292), .B(o[330]), .Z(n31337) );
  XOR U32523 ( .A(n31336), .B(n31337), .Z(n31359) );
  AND U32524 ( .A(y[8005]), .B(x[486]), .Z(n31294) );
  NAND U32525 ( .A(y[8010]), .B(x[481]), .Z(n31293) );
  XNOR U32526 ( .A(n31294), .B(n31293), .Z(n31327) );
  AND U32527 ( .A(x[490]), .B(y[8001]), .Z(n31345) );
  XOR U32528 ( .A(o[331]), .B(n31345), .Z(n31326) );
  XOR U32529 ( .A(n31327), .B(n31326), .Z(n31358) );
  XOR U32530 ( .A(n31359), .B(n31358), .Z(n31361) );
  XOR U32531 ( .A(n31360), .B(n31361), .Z(n31365) );
  XOR U32532 ( .A(n31364), .B(n31365), .Z(n31367) );
  XNOR U32533 ( .A(n31366), .B(n31367), .Z(n31349) );
  NAND U32534 ( .A(x[483]), .B(y[8008]), .Z(n32336) );
  NAND U32535 ( .A(y[8009]), .B(x[482]), .Z(n31295) );
  XNOR U32536 ( .A(n31296), .B(n31295), .Z(n31322) );
  AND U32537 ( .A(x[484]), .B(y[8007]), .Z(n31321) );
  XNOR U32538 ( .A(n31322), .B(n31321), .Z(n31353) );
  XOR U32539 ( .A(n32336), .B(n31353), .Z(n31354) );
  NAND U32540 ( .A(y[8002]), .B(x[489]), .Z(n31297) );
  XNOR U32541 ( .A(n31298), .B(n31297), .Z(n31341) );
  AND U32542 ( .A(x[488]), .B(y[8003]), .Z(n31342) );
  XOR U32543 ( .A(n31341), .B(n31342), .Z(n31355) );
  AND U32544 ( .A(x[483]), .B(y[8009]), .Z(n31335) );
  IV U32545 ( .A(n31335), .Z(n31403) );
  AND U32546 ( .A(x[481]), .B(y[8007]), .Z(n31598) );
  NANDN U32547 ( .A(n31403), .B(n31598), .Z(n31302) );
  NAND U32548 ( .A(n31300), .B(n31299), .Z(n31301) );
  NAND U32549 ( .A(n31302), .B(n31301), .Z(n31316) );
  NAND U32550 ( .A(n31475), .B(n31303), .Z(n31307) );
  NAND U32551 ( .A(n31305), .B(n31304), .Z(n31306) );
  NAND U32552 ( .A(n31307), .B(n31306), .Z(n31315) );
  XOR U32553 ( .A(n31316), .B(n31315), .Z(n31317) );
  NANDN U32554 ( .A(n31309), .B(n31308), .Z(n31313) );
  NAND U32555 ( .A(n31311), .B(n31310), .Z(n31312) );
  NAND U32556 ( .A(n31313), .B(n31312), .Z(n31347) );
  XOR U32557 ( .A(n31349), .B(n31350), .Z(n31370) );
  XOR U32558 ( .A(n31371), .B(n31370), .Z(n31372) );
  XOR U32559 ( .A(n31373), .B(n31372), .Z(n31379) );
  XNOR U32560 ( .A(n31377), .B(n31379), .Z(n31314) );
  XOR U32561 ( .A(n31376), .B(n31314), .Z(N684) );
  NAND U32562 ( .A(n31316), .B(n31315), .Z(n31320) );
  NANDN U32563 ( .A(n31318), .B(n31317), .Z(n31319) );
  NAND U32564 ( .A(n31320), .B(n31319), .Z(n31439) );
  AND U32565 ( .A(x[485]), .B(y[8009]), .Z(n31849) );
  AND U32566 ( .A(x[482]), .B(y[8006]), .Z(n32025) );
  NAND U32567 ( .A(n31849), .B(n32025), .Z(n31324) );
  NAND U32568 ( .A(n31322), .B(n31321), .Z(n31323) );
  AND U32569 ( .A(n31324), .B(n31323), .Z(n31391) );
  AND U32570 ( .A(x[486]), .B(y[8010]), .Z(n31615) );
  NAND U32571 ( .A(n31615), .B(n31325), .Z(n31329) );
  NAND U32572 ( .A(n31327), .B(n31326), .Z(n31328) );
  NAND U32573 ( .A(n31329), .B(n31328), .Z(n31390) );
  AND U32574 ( .A(x[489]), .B(y[8003]), .Z(n32020) );
  AND U32575 ( .A(y[8002]), .B(x[490]), .Z(n32063) );
  AND U32576 ( .A(y[8008]), .B(x[484]), .Z(n31330) );
  XOR U32577 ( .A(n32063), .B(n31330), .Z(n31430) );
  XOR U32578 ( .A(n32020), .B(n31430), .Z(n31413) );
  NAND U32579 ( .A(x[487]), .B(y[8005]), .Z(n31411) );
  XOR U32580 ( .A(n31412), .B(n31411), .Z(n31414) );
  AND U32581 ( .A(y[8000]), .B(x[492]), .Z(n31332) );
  NAND U32582 ( .A(y[8012]), .B(x[480]), .Z(n31331) );
  XNOR U32583 ( .A(n31332), .B(n31331), .Z(n31426) );
  AND U32584 ( .A(x[491]), .B(y[8001]), .Z(n31406) );
  XOR U32585 ( .A(n31406), .B(o[332]), .Z(n31425) );
  XOR U32586 ( .A(n31426), .B(n31425), .Z(n31397) );
  AND U32587 ( .A(y[8010]), .B(x[482]), .Z(n31334) );
  NAND U32588 ( .A(y[8004]), .B(x[488]), .Z(n31333) );
  XNOR U32589 ( .A(n31334), .B(n31333), .Z(n31402) );
  XOR U32590 ( .A(n31402), .B(n31335), .Z(n31396) );
  XOR U32591 ( .A(n31397), .B(n31396), .Z(n31399) );
  XOR U32592 ( .A(n31398), .B(n31399), .Z(n31392) );
  XOR U32593 ( .A(n31393), .B(n31392), .Z(n31437) );
  AND U32594 ( .A(x[491]), .B(y[8011]), .Z(n32423) );
  NAND U32595 ( .A(n32423), .B(n31603), .Z(n31339) );
  NAND U32596 ( .A(n31337), .B(n31336), .Z(n31338) );
  NAND U32597 ( .A(n31339), .B(n31338), .Z(n31420) );
  AND U32598 ( .A(x[489]), .B(y[8004]), .Z(n31340) );
  AND U32599 ( .A(x[487]), .B(y[8002]), .Z(n31542) );
  NAND U32600 ( .A(n31340), .B(n31542), .Z(n31344) );
  NAND U32601 ( .A(n31342), .B(n31341), .Z(n31343) );
  NAND U32602 ( .A(n31344), .B(n31343), .Z(n31418) );
  AND U32603 ( .A(y[8011]), .B(x[481]), .Z(n32058) );
  XOR U32604 ( .A(n31346), .B(n32058), .Z(n31423) );
  XOR U32605 ( .A(n31424), .B(n31423), .Z(n31417) );
  XOR U32606 ( .A(n31418), .B(n31417), .Z(n31419) );
  XNOR U32607 ( .A(n31420), .B(n31419), .Z(n31438) );
  XNOR U32608 ( .A(n31437), .B(n31438), .Z(n31440) );
  XOR U32609 ( .A(n31439), .B(n31440), .Z(n31447) );
  NANDN U32610 ( .A(n31348), .B(n31347), .Z(n31352) );
  NANDN U32611 ( .A(n31350), .B(n31349), .Z(n31351) );
  NAND U32612 ( .A(n31352), .B(n31351), .Z(n31446) );
  IV U32613 ( .A(n32336), .Z(n32034) );
  NANDN U32614 ( .A(n32034), .B(n31353), .Z(n31357) );
  NANDN U32615 ( .A(n31355), .B(n31354), .Z(n31356) );
  NAND U32616 ( .A(n31357), .B(n31356), .Z(n31384) );
  NAND U32617 ( .A(n31359), .B(n31358), .Z(n31363) );
  NAND U32618 ( .A(n31361), .B(n31360), .Z(n31362) );
  AND U32619 ( .A(n31363), .B(n31362), .Z(n31385) );
  XOR U32620 ( .A(n31384), .B(n31385), .Z(n31387) );
  NAND U32621 ( .A(n31365), .B(n31364), .Z(n31369) );
  NAND U32622 ( .A(n31367), .B(n31366), .Z(n31368) );
  AND U32623 ( .A(n31369), .B(n31368), .Z(n31386) );
  XOR U32624 ( .A(n31387), .B(n31386), .Z(n31448) );
  XOR U32625 ( .A(n31449), .B(n31448), .Z(n31445) );
  NAND U32626 ( .A(n31371), .B(n31370), .Z(n31375) );
  NAND U32627 ( .A(n31373), .B(n31372), .Z(n31374) );
  NAND U32628 ( .A(n31375), .B(n31374), .Z(n31444) );
  NANDN U32629 ( .A(n31376), .B(n31377), .Z(n31382) );
  NOR U32630 ( .A(n31378), .B(n31377), .Z(n31380) );
  OR U32631 ( .A(n31380), .B(n31379), .Z(n31381) );
  AND U32632 ( .A(n31382), .B(n31381), .Z(n31443) );
  XOR U32633 ( .A(n31444), .B(n31443), .Z(n31383) );
  XNOR U32634 ( .A(n31445), .B(n31383), .Z(N685) );
  NAND U32635 ( .A(n31385), .B(n31384), .Z(n31389) );
  NAND U32636 ( .A(n31387), .B(n31386), .Z(n31388) );
  NAND U32637 ( .A(n31389), .B(n31388), .Z(n31517) );
  NANDN U32638 ( .A(n31391), .B(n31390), .Z(n31395) );
  NAND U32639 ( .A(n31393), .B(n31392), .Z(n31394) );
  AND U32640 ( .A(n31395), .B(n31394), .Z(n31454) );
  NAND U32641 ( .A(n31397), .B(n31396), .Z(n31401) );
  NAND U32642 ( .A(n31399), .B(n31398), .Z(n31400) );
  NAND U32643 ( .A(n31401), .B(n31400), .Z(n31461) );
  AND U32644 ( .A(y[8010]), .B(x[488]), .Z(n32679) );
  AND U32645 ( .A(x[482]), .B(y[8004]), .Z(n31552) );
  NAND U32646 ( .A(n32679), .B(n31552), .Z(n31405) );
  NANDN U32647 ( .A(n31403), .B(n31402), .Z(n31404) );
  NAND U32648 ( .A(n31405), .B(n31404), .Z(n31485) );
  AND U32649 ( .A(n31406), .B(o[332]), .Z(n31479) );
  AND U32650 ( .A(y[8012]), .B(x[481]), .Z(n31407) );
  XOR U32651 ( .A(n31408), .B(n31407), .Z(n31478) );
  XOR U32652 ( .A(n31479), .B(n31478), .Z(n31484) );
  AND U32653 ( .A(x[486]), .B(y[8007]), .Z(n32463) );
  AND U32654 ( .A(y[8011]), .B(x[482]), .Z(n31410) );
  NAND U32655 ( .A(y[8004]), .B(x[489]), .Z(n31409) );
  XNOR U32656 ( .A(n31410), .B(n31409), .Z(n31488) );
  XOR U32657 ( .A(n32463), .B(n31488), .Z(n31483) );
  XOR U32658 ( .A(n31484), .B(n31483), .Z(n31486) );
  XOR U32659 ( .A(n31485), .B(n31486), .Z(n31460) );
  NAND U32660 ( .A(n31412), .B(n31411), .Z(n31416) );
  ANDN U32661 ( .B(n31414), .A(n31413), .Z(n31415) );
  ANDN U32662 ( .B(n31416), .A(n31415), .Z(n31459) );
  XOR U32663 ( .A(n31460), .B(n31459), .Z(n31462) );
  XOR U32664 ( .A(n31461), .B(n31462), .Z(n31453) );
  NAND U32665 ( .A(n31418), .B(n31417), .Z(n31422) );
  NAND U32666 ( .A(n31420), .B(n31419), .Z(n31421) );
  NAND U32667 ( .A(n31422), .B(n31421), .Z(n31467) );
  AND U32668 ( .A(x[486]), .B(y[8011]), .Z(n31776) );
  IV U32669 ( .A(n31776), .Z(n31851) );
  AND U32670 ( .A(x[481]), .B(y[8006]), .Z(n31477) );
  AND U32671 ( .A(x[492]), .B(y[8012]), .Z(n32685) );
  AND U32672 ( .A(x[490]), .B(y[8003]), .Z(n32348) );
  AND U32673 ( .A(y[8002]), .B(x[491]), .Z(n32309) );
  AND U32674 ( .A(y[8005]), .B(x[488]), .Z(n31427) );
  XOR U32675 ( .A(n32309), .B(n31427), .Z(n31476) );
  XOR U32676 ( .A(n32348), .B(n31476), .Z(n31472) );
  XOR U32677 ( .A(n31471), .B(n31472), .Z(n31474) );
  XOR U32678 ( .A(n31473), .B(n31474), .Z(n31465) );
  AND U32679 ( .A(x[490]), .B(y[8008]), .Z(n31429) );
  AND U32680 ( .A(x[484]), .B(y[8002]), .Z(n31428) );
  NAND U32681 ( .A(n31429), .B(n31428), .Z(n31432) );
  NAND U32682 ( .A(n32020), .B(n31430), .Z(n31431) );
  NAND U32683 ( .A(n31432), .B(n31431), .Z(n31504) );
  AND U32684 ( .A(y[8000]), .B(x[493]), .Z(n31434) );
  NAND U32685 ( .A(y[8013]), .B(x[480]), .Z(n31433) );
  XNOR U32686 ( .A(n31434), .B(n31433), .Z(n31499) );
  AND U32687 ( .A(x[492]), .B(y[8001]), .Z(n31491) );
  XOR U32688 ( .A(n31491), .B(o[333]), .Z(n31498) );
  XOR U32689 ( .A(n31499), .B(n31498), .Z(n31503) );
  AND U32690 ( .A(y[8008]), .B(x[485]), .Z(n31436) );
  NAND U32691 ( .A(y[8010]), .B(x[483]), .Z(n31435) );
  XNOR U32692 ( .A(n31436), .B(n31435), .Z(n31497) );
  AND U32693 ( .A(x[484]), .B(y[8009]), .Z(n31496) );
  XOR U32694 ( .A(n31497), .B(n31496), .Z(n31502) );
  XOR U32695 ( .A(n31503), .B(n31502), .Z(n31505) );
  XOR U32696 ( .A(n31504), .B(n31505), .Z(n31466) );
  XOR U32697 ( .A(n31465), .B(n31466), .Z(n31468) );
  XOR U32698 ( .A(n31467), .B(n31468), .Z(n31455) );
  XOR U32699 ( .A(n31456), .B(n31455), .Z(n31516) );
  NANDN U32700 ( .A(n31438), .B(n31437), .Z(n31442) );
  NAND U32701 ( .A(n31440), .B(n31439), .Z(n31441) );
  AND U32702 ( .A(n31442), .B(n31441), .Z(n31515) );
  XOR U32703 ( .A(n31517), .B(n31518), .Z(n31511) );
  NANDN U32704 ( .A(n31447), .B(n31446), .Z(n31451) );
  NAND U32705 ( .A(n31449), .B(n31448), .Z(n31450) );
  AND U32706 ( .A(n31451), .B(n31450), .Z(n31509) );
  IV U32707 ( .A(n31509), .Z(n31508) );
  XOR U32708 ( .A(n31510), .B(n31508), .Z(n31452) );
  XNOR U32709 ( .A(n31511), .B(n31452), .Z(N686) );
  NANDN U32710 ( .A(n31454), .B(n31453), .Z(n31458) );
  NAND U32711 ( .A(n31456), .B(n31455), .Z(n31457) );
  AND U32712 ( .A(n31458), .B(n31457), .Z(n31592) );
  NAND U32713 ( .A(n31460), .B(n31459), .Z(n31464) );
  NAND U32714 ( .A(n31462), .B(n31461), .Z(n31463) );
  NAND U32715 ( .A(n31464), .B(n31463), .Z(n31591) );
  NAND U32716 ( .A(n31466), .B(n31465), .Z(n31470) );
  NAND U32717 ( .A(n31468), .B(n31467), .Z(n31469) );
  NAND U32718 ( .A(n31470), .B(n31469), .Z(n31524) );
  AND U32719 ( .A(x[491]), .B(y[8005]), .Z(n31627) );
  NAND U32720 ( .A(x[487]), .B(y[8012]), .Z(n32036) );
  XOR U32721 ( .A(n31574), .B(n31575), .Z(n31577) );
  AND U32722 ( .A(x[484]), .B(y[8010]), .Z(n31956) );
  AND U32723 ( .A(y[8011]), .B(x[483]), .Z(n31481) );
  NAND U32724 ( .A(y[8006]), .B(x[488]), .Z(n31480) );
  XNOR U32725 ( .A(n31481), .B(n31480), .Z(n31564) );
  XOR U32726 ( .A(n31849), .B(n31564), .Z(n31571) );
  XOR U32727 ( .A(n31956), .B(n31571), .Z(n31573) );
  AND U32728 ( .A(x[489]), .B(y[8005]), .Z(n32148) );
  AND U32729 ( .A(y[8012]), .B(x[482]), .Z(n31482) );
  AND U32730 ( .A(y[8004]), .B(x[490]), .Z(n32166) );
  XOR U32731 ( .A(n31482), .B(n32166), .Z(n31553) );
  XOR U32732 ( .A(n32148), .B(n31553), .Z(n31572) );
  XOR U32733 ( .A(n31573), .B(n31572), .Z(n31576) );
  XOR U32734 ( .A(n31577), .B(n31576), .Z(n31529) );
  XOR U32735 ( .A(n31529), .B(n31528), .Z(n31531) );
  XOR U32736 ( .A(n31530), .B(n31531), .Z(n31523) );
  AND U32737 ( .A(x[489]), .B(y[8011]), .Z(n31487) );
  NAND U32738 ( .A(n31487), .B(n31552), .Z(n31490) );
  NAND U32739 ( .A(n32463), .B(n31488), .Z(n31489) );
  NAND U32740 ( .A(n31490), .B(n31489), .Z(n31540) );
  AND U32741 ( .A(n31491), .B(o[333]), .Z(n31562) );
  AND U32742 ( .A(y[8000]), .B(x[494]), .Z(n31493) );
  AND U32743 ( .A(y[8014]), .B(x[480]), .Z(n31492) );
  XOR U32744 ( .A(n31493), .B(n31492), .Z(n31561) );
  XOR U32745 ( .A(n31562), .B(n31561), .Z(n31539) );
  NAND U32746 ( .A(y[8002]), .B(x[492]), .Z(n31494) );
  XNOR U32747 ( .A(n31495), .B(n31494), .Z(n31544) );
  AND U32748 ( .A(x[493]), .B(y[8001]), .Z(n31551) );
  XOR U32749 ( .A(o[334]), .B(n31551), .Z(n31543) );
  XOR U32750 ( .A(n31544), .B(n31543), .Z(n31538) );
  XOR U32751 ( .A(n31539), .B(n31538), .Z(n31541) );
  XNOR U32752 ( .A(n31540), .B(n31541), .Z(n31579) );
  NAND U32753 ( .A(x[485]), .B(y[8010]), .Z(n31616) );
  AND U32754 ( .A(x[493]), .B(y[8013]), .Z(n33069) );
  NAND U32755 ( .A(y[8003]), .B(x[491]), .Z(n31500) );
  XNOR U32756 ( .A(n31501), .B(n31500), .Z(n31558) );
  AND U32757 ( .A(x[481]), .B(y[8013]), .Z(n31557) );
  XOR U32758 ( .A(n31558), .B(n31557), .Z(n31534) );
  XNOR U32759 ( .A(n31535), .B(n31534), .Z(n31537) );
  XOR U32760 ( .A(n31536), .B(n31537), .Z(n31578) );
  XOR U32761 ( .A(n31579), .B(n31578), .Z(n31581) );
  NAND U32762 ( .A(n31503), .B(n31502), .Z(n31507) );
  NAND U32763 ( .A(n31505), .B(n31504), .Z(n31506) );
  AND U32764 ( .A(n31507), .B(n31506), .Z(n31580) );
  XNOR U32765 ( .A(n31581), .B(n31580), .Z(n31522) );
  XOR U32766 ( .A(n31523), .B(n31522), .Z(n31525) );
  XOR U32767 ( .A(n31524), .B(n31525), .Z(n31593) );
  XNOR U32768 ( .A(n31594), .B(n31593), .Z(n31587) );
  OR U32769 ( .A(n31510), .B(n31508), .Z(n31514) );
  ANDN U32770 ( .B(n31510), .A(n31509), .Z(n31512) );
  OR U32771 ( .A(n31512), .B(n31511), .Z(n31513) );
  AND U32772 ( .A(n31514), .B(n31513), .Z(n31586) );
  NANDN U32773 ( .A(n31516), .B(n31515), .Z(n31520) );
  NAND U32774 ( .A(n31518), .B(n31517), .Z(n31519) );
  AND U32775 ( .A(n31520), .B(n31519), .Z(n31585) );
  IV U32776 ( .A(n31585), .Z(n31584) );
  XOR U32777 ( .A(n31586), .B(n31584), .Z(n31521) );
  XNOR U32778 ( .A(n31587), .B(n31521), .Z(N687) );
  NAND U32779 ( .A(n31523), .B(n31522), .Z(n31527) );
  NAND U32780 ( .A(n31525), .B(n31524), .Z(n31526) );
  NAND U32781 ( .A(n31527), .B(n31526), .Z(n31685) );
  NANDN U32782 ( .A(n31529), .B(n31528), .Z(n31533) );
  NANDN U32783 ( .A(n31531), .B(n31530), .Z(n31532) );
  NAND U32784 ( .A(n31533), .B(n31532), .Z(n31656) );
  AND U32785 ( .A(x[492]), .B(y[8007]), .Z(n32026) );
  NAND U32786 ( .A(n32026), .B(n31542), .Z(n31546) );
  NAND U32787 ( .A(n31544), .B(n31543), .Z(n31545) );
  AND U32788 ( .A(n31546), .B(n31545), .Z(n31636) );
  AND U32789 ( .A(y[8004]), .B(x[491]), .Z(n31548) );
  NAND U32790 ( .A(y[8002]), .B(x[493]), .Z(n31547) );
  XNOR U32791 ( .A(n31548), .B(n31547), .Z(n31640) );
  AND U32792 ( .A(x[492]), .B(y[8003]), .Z(n31641) );
  XNOR U32793 ( .A(n31640), .B(n31641), .Z(n31635) );
  AND U32794 ( .A(y[8000]), .B(x[495]), .Z(n31550) );
  NAND U32795 ( .A(y[8015]), .B(x[480]), .Z(n31549) );
  XNOR U32796 ( .A(n31550), .B(n31549), .Z(n31605) );
  AND U32797 ( .A(o[334]), .B(n31551), .Z(n31604) );
  XNOR U32798 ( .A(n31605), .B(n31604), .Z(n31634) );
  XNOR U32799 ( .A(n31635), .B(n31634), .Z(n31637) );
  XNOR U32800 ( .A(n31636), .B(n31637), .Z(n31667) );
  NAND U32801 ( .A(x[490]), .B(y[8012]), .Z(n32465) );
  NANDN U32802 ( .A(n32465), .B(n31552), .Z(n31555) );
  NAND U32803 ( .A(n32148), .B(n31553), .Z(n31554) );
  NAND U32804 ( .A(n31555), .B(n31554), .Z(n31665) );
  AND U32805 ( .A(x[491]), .B(y[8008]), .Z(n31955) );
  NAND U32806 ( .A(n31955), .B(n31556), .Z(n31560) );
  NAND U32807 ( .A(n31558), .B(n31557), .Z(n31559) );
  NAND U32808 ( .A(n31560), .B(n31559), .Z(n31664) );
  XOR U32809 ( .A(n31665), .B(n31664), .Z(n31666) );
  XOR U32810 ( .A(n31658), .B(n31659), .Z(n31661) );
  XOR U32811 ( .A(n31660), .B(n31661), .Z(n31655) );
  AND U32812 ( .A(x[494]), .B(y[8014]), .Z(n33338) );
  XOR U32813 ( .A(n31629), .B(n31628), .Z(n31630) );
  AND U32814 ( .A(y[8005]), .B(x[490]), .Z(n31566) );
  NAND U32815 ( .A(y[8011]), .B(x[484]), .Z(n31565) );
  XNOR U32816 ( .A(n31566), .B(n31565), .Z(n31610) );
  AND U32817 ( .A(x[487]), .B(y[8008]), .Z(n31611) );
  XNOR U32818 ( .A(n31610), .B(n31611), .Z(n31618) );
  NAND U32819 ( .A(x[486]), .B(y[8009]), .Z(n31726) );
  XOR U32820 ( .A(n31726), .B(n31616), .Z(n31617) );
  XOR U32821 ( .A(n31618), .B(n31617), .Z(n31651) );
  AND U32822 ( .A(y[8013]), .B(x[482]), .Z(n31568) );
  NAND U32823 ( .A(y[8006]), .B(x[489]), .Z(n31567) );
  XNOR U32824 ( .A(n31568), .B(n31567), .Z(n31620) );
  AND U32825 ( .A(x[483]), .B(y[8012]), .Z(n31619) );
  XOR U32826 ( .A(n31620), .B(n31619), .Z(n31649) );
  AND U32827 ( .A(y[8014]), .B(x[481]), .Z(n31570) );
  NAND U32828 ( .A(y[8007]), .B(x[488]), .Z(n31569) );
  XNOR U32829 ( .A(n31570), .B(n31569), .Z(n31600) );
  AND U32830 ( .A(x[494]), .B(y[8001]), .Z(n31625) );
  XOR U32831 ( .A(o[335]), .B(n31625), .Z(n31599) );
  XOR U32832 ( .A(n31600), .B(n31599), .Z(n31648) );
  XOR U32833 ( .A(n31649), .B(n31648), .Z(n31650) );
  XNOR U32834 ( .A(n31630), .B(n31631), .Z(n31671) );
  XOR U32835 ( .A(n31673), .B(n31672), .Z(n31654) );
  XNOR U32836 ( .A(n31655), .B(n31654), .Z(n31657) );
  XNOR U32837 ( .A(n31656), .B(n31657), .Z(n31684) );
  NAND U32838 ( .A(n31579), .B(n31578), .Z(n31583) );
  NAND U32839 ( .A(n31581), .B(n31580), .Z(n31582) );
  AND U32840 ( .A(n31583), .B(n31582), .Z(n31683) );
  XNOR U32841 ( .A(n31684), .B(n31683), .Z(n31686) );
  XOR U32842 ( .A(n31685), .B(n31686), .Z(n31679) );
  OR U32843 ( .A(n31586), .B(n31584), .Z(n31590) );
  ANDN U32844 ( .B(n31586), .A(n31585), .Z(n31588) );
  OR U32845 ( .A(n31588), .B(n31587), .Z(n31589) );
  AND U32846 ( .A(n31590), .B(n31589), .Z(n31678) );
  NANDN U32847 ( .A(n31592), .B(n31591), .Z(n31596) );
  NAND U32848 ( .A(n31594), .B(n31593), .Z(n31595) );
  NAND U32849 ( .A(n31596), .B(n31595), .Z(n31677) );
  IV U32850 ( .A(n31677), .Z(n31676) );
  XOR U32851 ( .A(n31678), .B(n31676), .Z(n31597) );
  XNOR U32852 ( .A(n31679), .B(n31597), .Z(N688) );
  AND U32853 ( .A(x[488]), .B(y[8014]), .Z(n31957) );
  NAND U32854 ( .A(n31957), .B(n31598), .Z(n31602) );
  NAND U32855 ( .A(n31600), .B(n31599), .Z(n31601) );
  NAND U32856 ( .A(n31602), .B(n31601), .Z(n31756) );
  AND U32857 ( .A(x[495]), .B(y[8015]), .Z(n33744) );
  NAND U32858 ( .A(n33744), .B(n31603), .Z(n31607) );
  NAND U32859 ( .A(n31605), .B(n31604), .Z(n31606) );
  NAND U32860 ( .A(n31607), .B(n31606), .Z(n31755) );
  XOR U32861 ( .A(n31756), .B(n31755), .Z(n31758) );
  AND U32862 ( .A(x[490]), .B(y[8011]), .Z(n31609) );
  NAND U32863 ( .A(n31609), .B(n31608), .Z(n31613) );
  NAND U32864 ( .A(n31611), .B(n31610), .Z(n31612) );
  NAND U32865 ( .A(n31613), .B(n31612), .Z(n31713) );
  AND U32866 ( .A(x[480]), .B(y[8016]), .Z(n31735) );
  AND U32867 ( .A(x[496]), .B(y[8000]), .Z(n31736) );
  XOR U32868 ( .A(n31735), .B(n31736), .Z(n31738) );
  AND U32869 ( .A(x[495]), .B(y[8001]), .Z(n31723) );
  XOR U32870 ( .A(o[336]), .B(n31723), .Z(n31737) );
  XOR U32871 ( .A(n31738), .B(n31737), .Z(n31712) );
  NAND U32872 ( .A(y[8009]), .B(x[487]), .Z(n31614) );
  XNOR U32873 ( .A(n31615), .B(n31614), .Z(n31728) );
  AND U32874 ( .A(x[490]), .B(y[8006]), .Z(n31727) );
  XOR U32875 ( .A(n31728), .B(n31727), .Z(n31711) );
  XOR U32876 ( .A(n31712), .B(n31711), .Z(n31714) );
  XOR U32877 ( .A(n31713), .B(n31714), .Z(n31757) );
  XOR U32878 ( .A(n31758), .B(n31757), .Z(n31708) );
  AND U32879 ( .A(x[489]), .B(y[8013]), .Z(n32445) );
  NAND U32880 ( .A(n32445), .B(n32025), .Z(n31622) );
  NAND U32881 ( .A(n31620), .B(n31619), .Z(n31621) );
  NAND U32882 ( .A(n31622), .B(n31621), .Z(n31745) );
  AND U32883 ( .A(y[8015]), .B(x[481]), .Z(n31624) );
  NAND U32884 ( .A(y[8008]), .B(x[488]), .Z(n31623) );
  XNOR U32885 ( .A(n31624), .B(n31623), .Z(n31732) );
  AND U32886 ( .A(o[335]), .B(n31625), .Z(n31731) );
  XOR U32887 ( .A(n31732), .B(n31731), .Z(n31744) );
  NAND U32888 ( .A(y[8002]), .B(x[494]), .Z(n31626) );
  XNOR U32889 ( .A(n31627), .B(n31626), .Z(n31767) );
  AND U32890 ( .A(x[484]), .B(y[8012]), .Z(n31768) );
  XOR U32891 ( .A(n31767), .B(n31768), .Z(n31743) );
  XOR U32892 ( .A(n31744), .B(n31743), .Z(n31746) );
  XNOR U32893 ( .A(n31745), .B(n31746), .Z(n31705) );
  XOR U32894 ( .A(n31706), .B(n31705), .Z(n31707) );
  NAND U32895 ( .A(n31629), .B(n31628), .Z(n31633) );
  NANDN U32896 ( .A(n31631), .B(n31630), .Z(n31632) );
  AND U32897 ( .A(n31633), .B(n31632), .Z(n31749) );
  XOR U32898 ( .A(n31750), .B(n31749), .Z(n31751) );
  NAND U32899 ( .A(n31635), .B(n31634), .Z(n31639) );
  NANDN U32900 ( .A(n31637), .B(n31636), .Z(n31638) );
  NAND U32901 ( .A(n31639), .B(n31638), .Z(n31781) );
  AND U32902 ( .A(x[493]), .B(y[8004]), .Z(n31778) );
  NAND U32903 ( .A(n32309), .B(n31778), .Z(n31643) );
  NAND U32904 ( .A(n31641), .B(n31640), .Z(n31642) );
  NAND U32905 ( .A(n31643), .B(n31642), .Z(n31764) );
  AND U32906 ( .A(y[8014]), .B(x[482]), .Z(n31645) );
  NAND U32907 ( .A(y[8007]), .B(x[489]), .Z(n31644) );
  XNOR U32908 ( .A(n31645), .B(n31644), .Z(n31771) );
  AND U32909 ( .A(x[483]), .B(y[8013]), .Z(n31772) );
  XOR U32910 ( .A(n31771), .B(n31772), .Z(n31762) );
  AND U32911 ( .A(x[492]), .B(y[8004]), .Z(n32434) );
  AND U32912 ( .A(y[8011]), .B(x[485]), .Z(n31647) );
  NAND U32913 ( .A(y[8003]), .B(x[493]), .Z(n31646) );
  XNOR U32914 ( .A(n31647), .B(n31646), .Z(n31718) );
  XOR U32915 ( .A(n32434), .B(n31718), .Z(n31761) );
  XOR U32916 ( .A(n31762), .B(n31761), .Z(n31763) );
  XOR U32917 ( .A(n31764), .B(n31763), .Z(n31780) );
  NAND U32918 ( .A(n31649), .B(n31648), .Z(n31653) );
  NANDN U32919 ( .A(n31651), .B(n31650), .Z(n31652) );
  AND U32920 ( .A(n31653), .B(n31652), .Z(n31779) );
  XOR U32921 ( .A(n31781), .B(n31782), .Z(n31752) );
  XNOR U32922 ( .A(n31751), .B(n31752), .Z(n31691) );
  XNOR U32923 ( .A(n31691), .B(n31690), .Z(n31693) );
  NAND U32924 ( .A(n31659), .B(n31658), .Z(n31663) );
  NAND U32925 ( .A(n31661), .B(n31660), .Z(n31662) );
  NAND U32926 ( .A(n31663), .B(n31662), .Z(n31701) );
  NAND U32927 ( .A(n31665), .B(n31664), .Z(n31669) );
  NANDN U32928 ( .A(n31667), .B(n31666), .Z(n31668) );
  NAND U32929 ( .A(n31669), .B(n31668), .Z(n31699) );
  NANDN U32930 ( .A(n31671), .B(n31670), .Z(n31675) );
  NAND U32931 ( .A(n31673), .B(n31672), .Z(n31674) );
  AND U32932 ( .A(n31675), .B(n31674), .Z(n31700) );
  XOR U32933 ( .A(n31699), .B(n31700), .Z(n31702) );
  XOR U32934 ( .A(n31701), .B(n31702), .Z(n31692) );
  XNOR U32935 ( .A(n31693), .B(n31692), .Z(n31698) );
  OR U32936 ( .A(n31678), .B(n31676), .Z(n31682) );
  ANDN U32937 ( .B(n31678), .A(n31677), .Z(n31680) );
  OR U32938 ( .A(n31680), .B(n31679), .Z(n31681) );
  AND U32939 ( .A(n31682), .B(n31681), .Z(n31697) );
  NAND U32940 ( .A(n31684), .B(n31683), .Z(n31688) );
  NANDN U32941 ( .A(n31686), .B(n31685), .Z(n31687) );
  NAND U32942 ( .A(n31688), .B(n31687), .Z(n31696) );
  XNOR U32943 ( .A(n31697), .B(n31696), .Z(n31689) );
  XNOR U32944 ( .A(n31698), .B(n31689), .Z(N689) );
  NANDN U32945 ( .A(n31691), .B(n31690), .Z(n31695) );
  NAND U32946 ( .A(n31693), .B(n31692), .Z(n31694) );
  AND U32947 ( .A(n31695), .B(n31694), .Z(n31793) );
  NAND U32948 ( .A(n31700), .B(n31699), .Z(n31704) );
  NAND U32949 ( .A(n31702), .B(n31701), .Z(n31703) );
  NAND U32950 ( .A(n31704), .B(n31703), .Z(n31788) );
  NAND U32951 ( .A(n31706), .B(n31705), .Z(n31710) );
  NANDN U32952 ( .A(n31708), .B(n31707), .Z(n31709) );
  NAND U32953 ( .A(n31710), .B(n31709), .Z(n31803) );
  NAND U32954 ( .A(n31712), .B(n31711), .Z(n31716) );
  NAND U32955 ( .A(n31714), .B(n31713), .Z(n31715) );
  NAND U32956 ( .A(n31716), .B(n31715), .Z(n31886) );
  AND U32957 ( .A(x[493]), .B(y[8011]), .Z(n32693) );
  NAND U32958 ( .A(n32693), .B(n31717), .Z(n31720) );
  NAND U32959 ( .A(n31718), .B(n32434), .Z(n31719) );
  NAND U32960 ( .A(n31720), .B(n31719), .Z(n31834) );
  AND U32961 ( .A(y[8016]), .B(x[481]), .Z(n31722) );
  NAND U32962 ( .A(y[8008]), .B(x[489]), .Z(n31721) );
  XNOR U32963 ( .A(n31722), .B(n31721), .Z(n31855) );
  AND U32964 ( .A(o[336]), .B(n31723), .Z(n31854) );
  XOR U32965 ( .A(n31855), .B(n31854), .Z(n31832) );
  AND U32966 ( .A(y[8002]), .B(x[495]), .Z(n31725) );
  NAND U32967 ( .A(y[8005]), .B(x[492]), .Z(n31724) );
  XNOR U32968 ( .A(n31725), .B(n31724), .Z(n31808) );
  AND U32969 ( .A(x[494]), .B(y[8003]), .Z(n31807) );
  XOR U32970 ( .A(n31808), .B(n31807), .Z(n31831) );
  XOR U32971 ( .A(n31832), .B(n31831), .Z(n31833) );
  XOR U32972 ( .A(n31834), .B(n31833), .Z(n31884) );
  AND U32973 ( .A(x[487]), .B(y[8010]), .Z(n31866) );
  NANDN U32974 ( .A(n31726), .B(n31866), .Z(n31730) );
  NAND U32975 ( .A(n31728), .B(n31727), .Z(n31729) );
  NAND U32976 ( .A(n31730), .B(n31729), .Z(n31844) );
  NAND U32977 ( .A(x[488]), .B(y[8015]), .Z(n32588) );
  AND U32978 ( .A(x[481]), .B(y[8008]), .Z(n31935) );
  NANDN U32979 ( .A(n32588), .B(n31935), .Z(n31734) );
  NAND U32980 ( .A(n31732), .B(n31731), .Z(n31733) );
  NAND U32981 ( .A(n31734), .B(n31733), .Z(n31843) );
  XOR U32982 ( .A(n31844), .B(n31843), .Z(n31846) );
  NAND U32983 ( .A(n31736), .B(n31735), .Z(n31740) );
  NAND U32984 ( .A(n31738), .B(n31737), .Z(n31739) );
  NAND U32985 ( .A(n31740), .B(n31739), .Z(n31840) );
  AND U32986 ( .A(x[480]), .B(y[8017]), .Z(n31822) );
  AND U32987 ( .A(x[497]), .B(y[8000]), .Z(n31821) );
  XOR U32988 ( .A(n31822), .B(n31821), .Z(n31824) );
  AND U32989 ( .A(x[496]), .B(y[8001]), .Z(n31818) );
  XOR U32990 ( .A(n31818), .B(o[337]), .Z(n31823) );
  XOR U32991 ( .A(n31824), .B(n31823), .Z(n31838) );
  AND U32992 ( .A(y[8015]), .B(x[482]), .Z(n31742) );
  NAND U32993 ( .A(y[8007]), .B(x[490]), .Z(n31741) );
  XNOR U32994 ( .A(n31742), .B(n31741), .Z(n31859) );
  AND U32995 ( .A(x[483]), .B(y[8014]), .Z(n31860) );
  XOR U32996 ( .A(n31859), .B(n31860), .Z(n31837) );
  XOR U32997 ( .A(n31838), .B(n31837), .Z(n31839) );
  XOR U32998 ( .A(n31840), .B(n31839), .Z(n31845) );
  XOR U32999 ( .A(n31846), .B(n31845), .Z(n31883) );
  XOR U33000 ( .A(n31884), .B(n31883), .Z(n31885) );
  XOR U33001 ( .A(n31886), .B(n31885), .Z(n31802) );
  NAND U33002 ( .A(n31744), .B(n31743), .Z(n31748) );
  NAND U33003 ( .A(n31746), .B(n31745), .Z(n31747) );
  AND U33004 ( .A(n31748), .B(n31747), .Z(n31801) );
  XOR U33005 ( .A(n31803), .B(n31804), .Z(n31787) );
  NAND U33006 ( .A(n31750), .B(n31749), .Z(n31754) );
  NANDN U33007 ( .A(n31752), .B(n31751), .Z(n31753) );
  NAND U33008 ( .A(n31754), .B(n31753), .Z(n31797) );
  NAND U33009 ( .A(n31756), .B(n31755), .Z(n31760) );
  NAND U33010 ( .A(n31758), .B(n31757), .Z(n31759) );
  NAND U33011 ( .A(n31760), .B(n31759), .Z(n31880) );
  NAND U33012 ( .A(n31762), .B(n31761), .Z(n31766) );
  NAND U33013 ( .A(n31764), .B(n31763), .Z(n31765) );
  NAND U33014 ( .A(n31766), .B(n31765), .Z(n31878) );
  AND U33015 ( .A(x[494]), .B(y[8005]), .Z(n32059) );
  NAND U33016 ( .A(n32309), .B(n32059), .Z(n31770) );
  NAND U33017 ( .A(n31768), .B(n31767), .Z(n31769) );
  NAND U33018 ( .A(n31770), .B(n31769), .Z(n31872) );
  AND U33019 ( .A(x[489]), .B(y[8014]), .Z(n32674) );
  NANDN U33020 ( .A(n31858), .B(n32674), .Z(n31774) );
  NAND U33021 ( .A(n31772), .B(n31771), .Z(n31773) );
  NAND U33022 ( .A(n31774), .B(n31773), .Z(n31871) );
  XOR U33023 ( .A(n31872), .B(n31871), .Z(n31874) );
  AND U33024 ( .A(y[8012]), .B(x[485]), .Z(n31918) );
  NAND U33025 ( .A(y[8009]), .B(x[488]), .Z(n31775) );
  XNOR U33026 ( .A(n31918), .B(n31775), .Z(n31850) );
  XOR U33027 ( .A(n31850), .B(n31776), .Z(n31865) );
  XOR U33028 ( .A(n31866), .B(n31865), .Z(n31868) );
  NAND U33029 ( .A(y[8013]), .B(x[484]), .Z(n31777) );
  XNOR U33030 ( .A(n31778), .B(n31777), .Z(n31812) );
  AND U33031 ( .A(x[491]), .B(y[8006]), .Z(n31813) );
  XOR U33032 ( .A(n31812), .B(n31813), .Z(n31867) );
  XOR U33033 ( .A(n31868), .B(n31867), .Z(n31873) );
  XOR U33034 ( .A(n31874), .B(n31873), .Z(n31877) );
  XOR U33035 ( .A(n31878), .B(n31877), .Z(n31879) );
  XOR U33036 ( .A(n31880), .B(n31879), .Z(n31796) );
  NANDN U33037 ( .A(n31780), .B(n31779), .Z(n31784) );
  NANDN U33038 ( .A(n31782), .B(n31781), .Z(n31783) );
  NAND U33039 ( .A(n31784), .B(n31783), .Z(n31795) );
  XOR U33040 ( .A(n31797), .B(n31798), .Z(n31786) );
  XOR U33041 ( .A(n31788), .B(n31789), .Z(n31794) );
  XOR U33042 ( .A(n31792), .B(n31794), .Z(n31785) );
  XOR U33043 ( .A(n31793), .B(n31785), .Z(N690) );
  NANDN U33044 ( .A(n31787), .B(n31786), .Z(n31791) );
  NAND U33045 ( .A(n31789), .B(n31788), .Z(n31790) );
  AND U33046 ( .A(n31791), .B(n31790), .Z(n31896) );
  NANDN U33047 ( .A(n31796), .B(n31795), .Z(n31800) );
  NANDN U33048 ( .A(n31798), .B(n31797), .Z(n31799) );
  AND U33049 ( .A(n31800), .B(n31799), .Z(n31893) );
  NANDN U33050 ( .A(n31802), .B(n31801), .Z(n31806) );
  NAND U33051 ( .A(n31804), .B(n31803), .Z(n31805) );
  AND U33052 ( .A(n31806), .B(n31805), .Z(n31891) );
  AND U33053 ( .A(x[492]), .B(y[8002]), .Z(n32138) );
  AND U33054 ( .A(x[495]), .B(y[8005]), .Z(n32033) );
  NAND U33055 ( .A(n32138), .B(n32033), .Z(n31810) );
  NAND U33056 ( .A(n31808), .B(n31807), .Z(n31809) );
  NAND U33057 ( .A(n31810), .B(n31809), .Z(n31983) );
  NAND U33058 ( .A(n33069), .B(n31811), .Z(n31815) );
  NAND U33059 ( .A(n31813), .B(n31812), .Z(n31814) );
  NAND U33060 ( .A(n31815), .B(n31814), .Z(n31974) );
  AND U33061 ( .A(y[8017]), .B(x[481]), .Z(n31817) );
  NAND U33062 ( .A(y[8008]), .B(x[490]), .Z(n31816) );
  XNOR U33063 ( .A(n31817), .B(n31816), .Z(n31936) );
  AND U33064 ( .A(n31818), .B(o[337]), .Z(n31937) );
  XOR U33065 ( .A(n31936), .B(n31937), .Z(n31972) );
  AND U33066 ( .A(y[8003]), .B(x[495]), .Z(n31820) );
  NAND U33067 ( .A(y[8009]), .B(x[489]), .Z(n31819) );
  XNOR U33068 ( .A(n31820), .B(n31819), .Z(n31927) );
  AND U33069 ( .A(x[494]), .B(y[8004]), .Z(n31928) );
  XOR U33070 ( .A(n31927), .B(n31928), .Z(n31971) );
  XOR U33071 ( .A(n31972), .B(n31971), .Z(n31973) );
  XOR U33072 ( .A(n31974), .B(n31973), .Z(n31984) );
  XOR U33073 ( .A(n31983), .B(n31984), .Z(n31986) );
  NAND U33074 ( .A(n31822), .B(n31821), .Z(n31826) );
  NAND U33075 ( .A(n31824), .B(n31823), .Z(n31825) );
  NAND U33076 ( .A(n31826), .B(n31825), .Z(n31995) );
  AND U33077 ( .A(y[8002]), .B(x[496]), .Z(n31828) );
  NAND U33078 ( .A(y[8007]), .B(x[491]), .Z(n31827) );
  XNOR U33079 ( .A(n31828), .B(n31827), .Z(n31923) );
  AND U33080 ( .A(x[482]), .B(y[8016]), .Z(n31924) );
  XOR U33081 ( .A(n31923), .B(n31924), .Z(n31996) );
  XOR U33082 ( .A(n31995), .B(n31996), .Z(n31998) );
  AND U33083 ( .A(y[8013]), .B(x[485]), .Z(n32042) );
  NAND U33084 ( .A(y[8012]), .B(x[486]), .Z(n31829) );
  XNOR U33085 ( .A(n32042), .B(n31829), .Z(n31920) );
  NAND U33086 ( .A(y[8014]), .B(x[484]), .Z(n31830) );
  XNOR U33087 ( .A(n32679), .B(n31830), .Z(n31959) );
  AND U33088 ( .A(x[487]), .B(y[8011]), .Z(n31958) );
  XOR U33089 ( .A(n31959), .B(n31958), .Z(n31919) );
  XOR U33090 ( .A(n31920), .B(n31919), .Z(n31997) );
  XOR U33091 ( .A(n31998), .B(n31997), .Z(n31985) );
  XNOR U33092 ( .A(n31986), .B(n31985), .Z(n31906) );
  NAND U33093 ( .A(n31832), .B(n31831), .Z(n31836) );
  NAND U33094 ( .A(n31834), .B(n31833), .Z(n31835) );
  AND U33095 ( .A(n31836), .B(n31835), .Z(n31978) );
  NAND U33096 ( .A(n31838), .B(n31837), .Z(n31842) );
  NAND U33097 ( .A(n31840), .B(n31839), .Z(n31841) );
  AND U33098 ( .A(n31842), .B(n31841), .Z(n31977) );
  XOR U33099 ( .A(n31978), .B(n31977), .Z(n31980) );
  NAND U33100 ( .A(n31844), .B(n31843), .Z(n31848) );
  NAND U33101 ( .A(n31846), .B(n31845), .Z(n31847) );
  AND U33102 ( .A(n31848), .B(n31847), .Z(n31979) );
  XOR U33103 ( .A(n31980), .B(n31979), .Z(n31905) );
  XOR U33104 ( .A(n31906), .B(n31905), .Z(n31908) );
  AND U33105 ( .A(x[488]), .B(y[8012]), .Z(n32172) );
  NAND U33106 ( .A(n32172), .B(n31849), .Z(n31853) );
  NANDN U33107 ( .A(n31851), .B(n31850), .Z(n31852) );
  NAND U33108 ( .A(n31853), .B(n31852), .Z(n31990) );
  NAND U33109 ( .A(x[489]), .B(y[8016]), .Z(n32812) );
  NANDN U33110 ( .A(n32812), .B(n31935), .Z(n31857) );
  NAND U33111 ( .A(n31855), .B(n31854), .Z(n31856) );
  NAND U33112 ( .A(n31857), .B(n31856), .Z(n31989) );
  XOR U33113 ( .A(n31990), .B(n31989), .Z(n31992) );
  NAND U33114 ( .A(x[490]), .B(y[8015]), .Z(n32702) );
  IV U33115 ( .A(n32702), .Z(n32813) );
  NANDN U33116 ( .A(n31858), .B(n32813), .Z(n31862) );
  NAND U33117 ( .A(n31860), .B(n31859), .Z(n31861) );
  NAND U33118 ( .A(n31862), .B(n31861), .Z(n31968) );
  AND U33119 ( .A(x[480]), .B(y[8018]), .Z(n31940) );
  AND U33120 ( .A(x[498]), .B(y[8000]), .Z(n31941) );
  XOR U33121 ( .A(n31940), .B(n31941), .Z(n31943) );
  AND U33122 ( .A(x[497]), .B(y[8001]), .Z(n31962) );
  XOR U33123 ( .A(o[338]), .B(n31962), .Z(n31942) );
  XOR U33124 ( .A(n31943), .B(n31942), .Z(n31966) );
  AND U33125 ( .A(y[8005]), .B(x[493]), .Z(n31864) );
  NAND U33126 ( .A(y[8015]), .B(x[483]), .Z(n31863) );
  XNOR U33127 ( .A(n31864), .B(n31863), .Z(n31948) );
  AND U33128 ( .A(x[492]), .B(y[8006]), .Z(n31949) );
  XOR U33129 ( .A(n31948), .B(n31949), .Z(n31965) );
  XOR U33130 ( .A(n31966), .B(n31965), .Z(n31967) );
  XOR U33131 ( .A(n31968), .B(n31967), .Z(n31991) );
  XNOR U33132 ( .A(n31992), .B(n31991), .Z(n31912) );
  NAND U33133 ( .A(n31866), .B(n31865), .Z(n31870) );
  NAND U33134 ( .A(n31868), .B(n31867), .Z(n31869) );
  AND U33135 ( .A(n31870), .B(n31869), .Z(n31911) );
  XOR U33136 ( .A(n31912), .B(n31911), .Z(n31913) );
  NAND U33137 ( .A(n31872), .B(n31871), .Z(n31876) );
  NAND U33138 ( .A(n31874), .B(n31873), .Z(n31875) );
  AND U33139 ( .A(n31876), .B(n31875), .Z(n31914) );
  XOR U33140 ( .A(n31913), .B(n31914), .Z(n31907) );
  XNOR U33141 ( .A(n31908), .B(n31907), .Z(n31902) );
  NAND U33142 ( .A(n31878), .B(n31877), .Z(n31882) );
  NAND U33143 ( .A(n31880), .B(n31879), .Z(n31881) );
  NAND U33144 ( .A(n31882), .B(n31881), .Z(n31900) );
  NAND U33145 ( .A(n31884), .B(n31883), .Z(n31888) );
  NAND U33146 ( .A(n31886), .B(n31885), .Z(n31887) );
  NAND U33147 ( .A(n31888), .B(n31887), .Z(n31899) );
  XOR U33148 ( .A(n31900), .B(n31899), .Z(n31901) );
  XOR U33149 ( .A(n31902), .B(n31901), .Z(n31890) );
  XOR U33150 ( .A(n31891), .B(n31890), .Z(n31892) );
  XOR U33151 ( .A(n31893), .B(n31892), .Z(n31898) );
  XNOR U33152 ( .A(n31897), .B(n31898), .Z(n31889) );
  XOR U33153 ( .A(n31896), .B(n31889), .Z(N691) );
  NAND U33154 ( .A(n31891), .B(n31890), .Z(n31895) );
  NAND U33155 ( .A(n31893), .B(n31892), .Z(n31894) );
  AND U33156 ( .A(n31895), .B(n31894), .Z(n32116) );
  NAND U33157 ( .A(n31900), .B(n31899), .Z(n31904) );
  NAND U33158 ( .A(n31902), .B(n31901), .Z(n31903) );
  NAND U33159 ( .A(n31904), .B(n31903), .Z(n32113) );
  NAND U33160 ( .A(n31906), .B(n31905), .Z(n31910) );
  NAND U33161 ( .A(n31908), .B(n31907), .Z(n31909) );
  AND U33162 ( .A(n31910), .B(n31909), .Z(n32111) );
  NAND U33163 ( .A(n31912), .B(n31911), .Z(n31916) );
  NAND U33164 ( .A(n31914), .B(n31913), .Z(n31915) );
  NAND U33165 ( .A(n31916), .B(n31915), .Z(n32005) );
  AND U33166 ( .A(x[486]), .B(y[8013]), .Z(n31917) );
  NAND U33167 ( .A(n31918), .B(n31917), .Z(n31922) );
  NAND U33168 ( .A(n31920), .B(n31919), .Z(n31921) );
  NAND U33169 ( .A(n31922), .B(n31921), .Z(n32095) );
  AND U33170 ( .A(x[496]), .B(y[8007]), .Z(n32450) );
  NAND U33171 ( .A(n32450), .B(n32309), .Z(n31926) );
  NAND U33172 ( .A(n31924), .B(n31923), .Z(n31925) );
  NAND U33173 ( .A(n31926), .B(n31925), .Z(n32093) );
  AND U33174 ( .A(x[495]), .B(y[8009]), .Z(n32707) );
  NAND U33175 ( .A(n32707), .B(n32020), .Z(n31930) );
  NAND U33176 ( .A(n31928), .B(n31927), .Z(n31929) );
  NAND U33177 ( .A(n31930), .B(n31929), .Z(n32010) );
  AND U33178 ( .A(y[8018]), .B(x[481]), .Z(n31932) );
  NAND U33179 ( .A(y[8011]), .B(x[488]), .Z(n31931) );
  XNOR U33180 ( .A(n31932), .B(n31931), .Z(n32060) );
  XOR U33181 ( .A(n32059), .B(n32060), .Z(n32009) );
  AND U33182 ( .A(y[8006]), .B(x[493]), .Z(n31934) );
  NAND U33183 ( .A(y[8017]), .B(x[482]), .Z(n31933) );
  XNOR U33184 ( .A(n31934), .B(n31933), .Z(n32027) );
  XOR U33185 ( .A(n32027), .B(n32026), .Z(n32008) );
  XOR U33186 ( .A(n32009), .B(n32008), .Z(n32011) );
  XOR U33187 ( .A(n32010), .B(n32011), .Z(n32092) );
  XOR U33188 ( .A(n32093), .B(n32092), .Z(n32094) );
  XNOR U33189 ( .A(n32095), .B(n32094), .Z(n32003) );
  AND U33190 ( .A(x[490]), .B(y[8017]), .Z(n33161) );
  IV U33191 ( .A(n33161), .Z(n33022) );
  NANDN U33192 ( .A(n33022), .B(n31935), .Z(n31939) );
  NAND U33193 ( .A(n31937), .B(n31936), .Z(n31938) );
  NAND U33194 ( .A(n31939), .B(n31938), .Z(n32070) );
  NAND U33195 ( .A(n31941), .B(n31940), .Z(n31945) );
  NAND U33196 ( .A(n31943), .B(n31942), .Z(n31944) );
  NAND U33197 ( .A(n31945), .B(n31944), .Z(n32068) );
  AND U33198 ( .A(y[8003]), .B(x[496]), .Z(n32758) );
  NAND U33199 ( .A(y[8010]), .B(x[489]), .Z(n31946) );
  XNOR U33200 ( .A(n32758), .B(n31946), .Z(n32022) );
  AND U33201 ( .A(x[495]), .B(y[8004]), .Z(n32021) );
  XOR U33202 ( .A(n32022), .B(n32021), .Z(n32069) );
  XOR U33203 ( .A(n32068), .B(n32069), .Z(n32071) );
  XNOR U33204 ( .A(n32070), .B(n32071), .Z(n32088) );
  AND U33205 ( .A(x[493]), .B(y[8015]), .Z(n33366) );
  NANDN U33206 ( .A(n31947), .B(n33366), .Z(n31951) );
  NAND U33207 ( .A(n31949), .B(n31948), .Z(n31950) );
  NAND U33208 ( .A(n31951), .B(n31950), .Z(n32076) );
  AND U33209 ( .A(y[8009]), .B(x[490]), .Z(n31953) );
  NAND U33210 ( .A(y[8002]), .B(x[497]), .Z(n31952) );
  XNOR U33211 ( .A(n31953), .B(n31952), .Z(n32065) );
  AND U33212 ( .A(x[498]), .B(y[8001]), .Z(n32041) );
  XOR U33213 ( .A(o[339]), .B(n32041), .Z(n32064) );
  XOR U33214 ( .A(n32065), .B(n32064), .Z(n32075) );
  NAND U33215 ( .A(y[8016]), .B(x[483]), .Z(n31954) );
  XNOR U33216 ( .A(n31955), .B(n31954), .Z(n32035) );
  XOR U33217 ( .A(n32075), .B(n32074), .Z(n32077) );
  XNOR U33218 ( .A(n32076), .B(n32077), .Z(n32087) );
  NAND U33219 ( .A(n31957), .B(n31956), .Z(n31961) );
  NAND U33220 ( .A(n31959), .B(n31958), .Z(n31960) );
  NAND U33221 ( .A(n31961), .B(n31960), .Z(n32016) );
  AND U33222 ( .A(o[338]), .B(n31962), .Z(n32049) );
  AND U33223 ( .A(x[480]), .B(y[8019]), .Z(n32046) );
  AND U33224 ( .A(x[499]), .B(y[8000]), .Z(n32047) );
  XOR U33225 ( .A(n32046), .B(n32047), .Z(n32048) );
  XOR U33226 ( .A(n32049), .B(n32048), .Z(n32015) );
  AND U33227 ( .A(x[484]), .B(y[8015]), .Z(n32186) );
  AND U33228 ( .A(y[8014]), .B(x[485]), .Z(n31964) );
  NAND U33229 ( .A(y[8013]), .B(x[486]), .Z(n31963) );
  XNOR U33230 ( .A(n31964), .B(n31963), .Z(n32043) );
  XOR U33231 ( .A(n32186), .B(n32043), .Z(n32014) );
  XOR U33232 ( .A(n32015), .B(n32014), .Z(n32017) );
  XNOR U33233 ( .A(n32016), .B(n32017), .Z(n32086) );
  XOR U33234 ( .A(n32087), .B(n32086), .Z(n32089) );
  XNOR U33235 ( .A(n32088), .B(n32089), .Z(n32082) );
  NAND U33236 ( .A(n31966), .B(n31965), .Z(n31970) );
  NAND U33237 ( .A(n31968), .B(n31967), .Z(n31969) );
  NAND U33238 ( .A(n31970), .B(n31969), .Z(n32081) );
  NAND U33239 ( .A(n31972), .B(n31971), .Z(n31976) );
  NAND U33240 ( .A(n31974), .B(n31973), .Z(n31975) );
  NAND U33241 ( .A(n31976), .B(n31975), .Z(n32080) );
  XOR U33242 ( .A(n32081), .B(n32080), .Z(n32083) );
  XNOR U33243 ( .A(n32082), .B(n32083), .Z(n32002) );
  XOR U33244 ( .A(n32003), .B(n32002), .Z(n32004) );
  XOR U33245 ( .A(n32005), .B(n32004), .Z(n32107) );
  NAND U33246 ( .A(n31978), .B(n31977), .Z(n31982) );
  NAND U33247 ( .A(n31980), .B(n31979), .Z(n31981) );
  AND U33248 ( .A(n31982), .B(n31981), .Z(n32104) );
  NAND U33249 ( .A(n31984), .B(n31983), .Z(n31988) );
  NAND U33250 ( .A(n31986), .B(n31985), .Z(n31987) );
  NAND U33251 ( .A(n31988), .B(n31987), .Z(n32100) );
  NAND U33252 ( .A(n31990), .B(n31989), .Z(n31994) );
  NAND U33253 ( .A(n31992), .B(n31991), .Z(n31993) );
  NAND U33254 ( .A(n31994), .B(n31993), .Z(n32099) );
  NAND U33255 ( .A(n31996), .B(n31995), .Z(n32000) );
  NAND U33256 ( .A(n31998), .B(n31997), .Z(n31999) );
  NAND U33257 ( .A(n32000), .B(n31999), .Z(n32098) );
  XNOR U33258 ( .A(n32099), .B(n32098), .Z(n32101) );
  XNOR U33259 ( .A(n32104), .B(n32105), .Z(n32106) );
  XOR U33260 ( .A(n32111), .B(n32110), .Z(n32112) );
  XOR U33261 ( .A(n32113), .B(n32112), .Z(n32118) );
  XNOR U33262 ( .A(n32117), .B(n32118), .Z(n32001) );
  XOR U33263 ( .A(n32116), .B(n32001), .Z(N692) );
  NAND U33264 ( .A(n32003), .B(n32002), .Z(n32007) );
  NAND U33265 ( .A(n32005), .B(n32004), .Z(n32006) );
  AND U33266 ( .A(n32007), .B(n32006), .Z(n32224) );
  NAND U33267 ( .A(n32009), .B(n32008), .Z(n32013) );
  NAND U33268 ( .A(n32011), .B(n32010), .Z(n32012) );
  NAND U33269 ( .A(n32013), .B(n32012), .Z(n32121) );
  NAND U33270 ( .A(n32015), .B(n32014), .Z(n32019) );
  NAND U33271 ( .A(n32017), .B(n32016), .Z(n32018) );
  NAND U33272 ( .A(n32019), .B(n32018), .Z(n32120) );
  XOR U33273 ( .A(n32121), .B(n32120), .Z(n32123) );
  AND U33274 ( .A(x[496]), .B(y[8010]), .Z(n32980) );
  NAND U33275 ( .A(n32980), .B(n32020), .Z(n32024) );
  NAND U33276 ( .A(n32022), .B(n32021), .Z(n32023) );
  NAND U33277 ( .A(n32024), .B(n32023), .Z(n32161) );
  AND U33278 ( .A(x[493]), .B(y[8017]), .Z(n33604) );
  NAND U33279 ( .A(n33604), .B(n32025), .Z(n32029) );
  NAND U33280 ( .A(n32027), .B(n32026), .Z(n32028) );
  NAND U33281 ( .A(n32029), .B(n32028), .Z(n32206) );
  AND U33282 ( .A(y[8004]), .B(x[496]), .Z(n32031) );
  NAND U33283 ( .A(y[8010]), .B(x[490]), .Z(n32030) );
  XNOR U33284 ( .A(n32031), .B(n32030), .Z(n32167) );
  AND U33285 ( .A(x[482]), .B(y[8018]), .Z(n32168) );
  XOR U33286 ( .A(n32167), .B(n32168), .Z(n32204) );
  NAND U33287 ( .A(y[8011]), .B(x[489]), .Z(n32032) );
  XNOR U33288 ( .A(n32033), .B(n32032), .Z(n32149) );
  AND U33289 ( .A(x[494]), .B(y[8006]), .Z(n32150) );
  XOR U33290 ( .A(n32149), .B(n32150), .Z(n32203) );
  XOR U33291 ( .A(n32204), .B(n32203), .Z(n32205) );
  XOR U33292 ( .A(n32206), .B(n32205), .Z(n32160) );
  XOR U33293 ( .A(n32161), .B(n32160), .Z(n32163) );
  NAND U33294 ( .A(x[491]), .B(y[8016]), .Z(n33162) );
  NANDN U33295 ( .A(n33162), .B(n32034), .Z(n32038) );
  NANDN U33296 ( .A(n32036), .B(n32035), .Z(n32037) );
  NAND U33297 ( .A(n32038), .B(n32037), .Z(n32212) );
  AND U33298 ( .A(y[8009]), .B(x[491]), .Z(n32040) );
  NAND U33299 ( .A(y[8019]), .B(x[481]), .Z(n32039) );
  XNOR U33300 ( .A(n32040), .B(n32039), .Z(n32145) );
  NAND U33301 ( .A(x[499]), .B(y[8001]), .Z(n32153) );
  XOR U33302 ( .A(n32145), .B(n32144), .Z(n32210) );
  AND U33303 ( .A(x[480]), .B(y[8020]), .Z(n32191) );
  AND U33304 ( .A(x[500]), .B(y[8000]), .Z(n32192) );
  XOR U33305 ( .A(n32191), .B(n32192), .Z(n32194) );
  AND U33306 ( .A(o[339]), .B(n32041), .Z(n32193) );
  XOR U33307 ( .A(n32194), .B(n32193), .Z(n32209) );
  XOR U33308 ( .A(n32210), .B(n32209), .Z(n32211) );
  XOR U33309 ( .A(n32212), .B(n32211), .Z(n32162) );
  XOR U33310 ( .A(n32163), .B(n32162), .Z(n32122) );
  XOR U33311 ( .A(n32123), .B(n32122), .Z(n32218) );
  NAND U33312 ( .A(x[486]), .B(y[8014]), .Z(n32155) );
  NANDN U33313 ( .A(n32155), .B(n32042), .Z(n32045) );
  NAND U33314 ( .A(n32043), .B(n32186), .Z(n32044) );
  NAND U33315 ( .A(n32045), .B(n32044), .Z(n32135) );
  NAND U33316 ( .A(n32047), .B(n32046), .Z(n32051) );
  NAND U33317 ( .A(n32049), .B(n32048), .Z(n32050) );
  NAND U33318 ( .A(n32051), .B(n32050), .Z(n32133) );
  AND U33319 ( .A(y[8002]), .B(x[498]), .Z(n32053) );
  NAND U33320 ( .A(y[8008]), .B(x[492]), .Z(n32052) );
  XNOR U33321 ( .A(n32053), .B(n32052), .Z(n32139) );
  AND U33322 ( .A(x[497]), .B(y[8003]), .Z(n32140) );
  XOR U33323 ( .A(n32139), .B(n32140), .Z(n32132) );
  XOR U33324 ( .A(n32133), .B(n32132), .Z(n32134) );
  XOR U33325 ( .A(n32135), .B(n32134), .Z(n32127) );
  AND U33326 ( .A(y[8007]), .B(x[493]), .Z(n32055) );
  NAND U33327 ( .A(y[8017]), .B(x[483]), .Z(n32054) );
  XNOR U33328 ( .A(n32055), .B(n32054), .Z(n32173) );
  XNOR U33329 ( .A(n32173), .B(n32172), .Z(n32157) );
  AND U33330 ( .A(y[8015]), .B(x[485]), .Z(n32057) );
  NAND U33331 ( .A(y[8016]), .B(x[484]), .Z(n32056) );
  XNOR U33332 ( .A(n32057), .B(n32056), .Z(n32188) );
  AND U33333 ( .A(x[487]), .B(y[8013]), .Z(n32187) );
  XNOR U33334 ( .A(n32188), .B(n32187), .Z(n32154) );
  XOR U33335 ( .A(n32155), .B(n32154), .Z(n32156) );
  XNOR U33336 ( .A(n32157), .B(n32156), .Z(n32199) );
  AND U33337 ( .A(x[488]), .B(y[8018]), .Z(n33318) );
  NAND U33338 ( .A(n33318), .B(n32058), .Z(n32062) );
  NAND U33339 ( .A(n32060), .B(n32059), .Z(n32061) );
  NAND U33340 ( .A(n32062), .B(n32061), .Z(n32198) );
  NAND U33341 ( .A(x[497]), .B(y[8009]), .Z(n32989) );
  NANDN U33342 ( .A(n32989), .B(n32063), .Z(n32067) );
  NAND U33343 ( .A(n32065), .B(n32064), .Z(n32066) );
  NAND U33344 ( .A(n32067), .B(n32066), .Z(n32197) );
  XOR U33345 ( .A(n32198), .B(n32197), .Z(n32200) );
  XNOR U33346 ( .A(n32199), .B(n32200), .Z(n32126) );
  NAND U33347 ( .A(n32069), .B(n32068), .Z(n32073) );
  NAND U33348 ( .A(n32071), .B(n32070), .Z(n32072) );
  AND U33349 ( .A(n32073), .B(n32072), .Z(n32128) );
  XOR U33350 ( .A(n32129), .B(n32128), .Z(n32216) );
  NAND U33351 ( .A(n32075), .B(n32074), .Z(n32079) );
  NAND U33352 ( .A(n32077), .B(n32076), .Z(n32078) );
  AND U33353 ( .A(n32079), .B(n32078), .Z(n32215) );
  XOR U33354 ( .A(n32216), .B(n32215), .Z(n32217) );
  NAND U33355 ( .A(n32081), .B(n32080), .Z(n32085) );
  NAND U33356 ( .A(n32083), .B(n32082), .Z(n32084) );
  AND U33357 ( .A(n32085), .B(n32084), .Z(n32230) );
  NAND U33358 ( .A(n32087), .B(n32086), .Z(n32091) );
  NAND U33359 ( .A(n32089), .B(n32088), .Z(n32090) );
  AND U33360 ( .A(n32091), .B(n32090), .Z(n32228) );
  NAND U33361 ( .A(n32093), .B(n32092), .Z(n32097) );
  NAND U33362 ( .A(n32095), .B(n32094), .Z(n32096) );
  AND U33363 ( .A(n32097), .B(n32096), .Z(n32227) );
  XNOR U33364 ( .A(n32230), .B(n32229), .Z(n32221) );
  XOR U33365 ( .A(n32222), .B(n32221), .Z(n32223) );
  XOR U33366 ( .A(n32224), .B(n32223), .Z(n32239) );
  NAND U33367 ( .A(n32099), .B(n32098), .Z(n32103) );
  NANDN U33368 ( .A(n32101), .B(n32100), .Z(n32102) );
  AND U33369 ( .A(n32103), .B(n32102), .Z(n32237) );
  NANDN U33370 ( .A(n32105), .B(n32104), .Z(n32109) );
  NANDN U33371 ( .A(n32107), .B(n32106), .Z(n32108) );
  AND U33372 ( .A(n32109), .B(n32108), .Z(n32236) );
  XOR U33373 ( .A(n32237), .B(n32236), .Z(n32238) );
  NAND U33374 ( .A(n32111), .B(n32110), .Z(n32115) );
  NAND U33375 ( .A(n32113), .B(n32112), .Z(n32114) );
  NAND U33376 ( .A(n32115), .B(n32114), .Z(n32234) );
  XOR U33377 ( .A(n32234), .B(n32233), .Z(n32119) );
  XNOR U33378 ( .A(n32235), .B(n32119), .Z(N693) );
  NAND U33379 ( .A(n32121), .B(n32120), .Z(n32125) );
  NAND U33380 ( .A(n32123), .B(n32122), .Z(n32124) );
  NAND U33381 ( .A(n32125), .B(n32124), .Z(n32251) );
  NANDN U33382 ( .A(n32127), .B(n32126), .Z(n32131) );
  NAND U33383 ( .A(n32129), .B(n32128), .Z(n32130) );
  AND U33384 ( .A(n32131), .B(n32130), .Z(n32249) );
  NAND U33385 ( .A(n32133), .B(n32132), .Z(n32137) );
  NAND U33386 ( .A(n32135), .B(n32134), .Z(n32136) );
  NAND U33387 ( .A(n32137), .B(n32136), .Z(n32270) );
  AND U33388 ( .A(x[498]), .B(y[8008]), .Z(n32987) );
  NAND U33389 ( .A(n32987), .B(n32138), .Z(n32142) );
  NAND U33390 ( .A(n32140), .B(n32139), .Z(n32141) );
  AND U33391 ( .A(n32142), .B(n32141), .Z(n32274) );
  AND U33392 ( .A(x[491]), .B(y[8019]), .Z(n33677) );
  AND U33393 ( .A(x[481]), .B(y[8009]), .Z(n32143) );
  NAND U33394 ( .A(n33677), .B(n32143), .Z(n32147) );
  NAND U33395 ( .A(n32145), .B(n32144), .Z(n32146) );
  NAND U33396 ( .A(n32147), .B(n32146), .Z(n32273) );
  AND U33397 ( .A(x[495]), .B(y[8011]), .Z(n32975) );
  NAND U33398 ( .A(n32975), .B(n32148), .Z(n32152) );
  NAND U33399 ( .A(n32150), .B(n32149), .Z(n32151) );
  NAND U33400 ( .A(n32152), .B(n32151), .Z(n32322) );
  AND U33401 ( .A(x[480]), .B(y[8021]), .Z(n32342) );
  NAND U33402 ( .A(x[501]), .B(y[8000]), .Z(n32343) );
  ANDN U33403 ( .B(o[340]), .A(n32153), .Z(n32344) );
  XOR U33404 ( .A(n32345), .B(n32344), .Z(n32321) );
  AND U33405 ( .A(x[485]), .B(y[8016]), .Z(n32327) );
  AND U33406 ( .A(x[496]), .B(y[8005]), .Z(n32326) );
  XOR U33407 ( .A(n32327), .B(n32326), .Z(n32329) );
  AND U33408 ( .A(x[495]), .B(y[8006]), .Z(n32328) );
  XOR U33409 ( .A(n32329), .B(n32328), .Z(n32320) );
  XOR U33410 ( .A(n32321), .B(n32320), .Z(n32323) );
  XOR U33411 ( .A(n32322), .B(n32323), .Z(n32275) );
  XOR U33412 ( .A(n32276), .B(n32275), .Z(n32267) );
  NAND U33413 ( .A(n32155), .B(n32154), .Z(n32159) );
  NAND U33414 ( .A(n32157), .B(n32156), .Z(n32158) );
  AND U33415 ( .A(n32159), .B(n32158), .Z(n32268) );
  XOR U33416 ( .A(n32267), .B(n32268), .Z(n32269) );
  XNOR U33417 ( .A(n32270), .B(n32269), .Z(n32250) );
  XNOR U33418 ( .A(n32249), .B(n32250), .Z(n32252) );
  XNOR U33419 ( .A(n32251), .B(n32252), .Z(n32245) );
  NAND U33420 ( .A(n32161), .B(n32160), .Z(n32165) );
  NAND U33421 ( .A(n32163), .B(n32162), .Z(n32164) );
  NAND U33422 ( .A(n32165), .B(n32164), .Z(n32258) );
  NAND U33423 ( .A(n32980), .B(n32166), .Z(n32170) );
  NAND U33424 ( .A(n32168), .B(n32167), .Z(n32169) );
  NAND U33425 ( .A(n32170), .B(n32169), .Z(n32292) );
  NAND U33426 ( .A(n33604), .B(n32171), .Z(n32175) );
  NAND U33427 ( .A(n32173), .B(n32172), .Z(n32174) );
  NAND U33428 ( .A(n32175), .B(n32174), .Z(n32288) );
  AND U33429 ( .A(y[8002]), .B(x[499]), .Z(n32177) );
  NAND U33430 ( .A(y[8010]), .B(x[491]), .Z(n32176) );
  XNOR U33431 ( .A(n32177), .B(n32176), .Z(n32311) );
  AND U33432 ( .A(x[500]), .B(y[8001]), .Z(n32341) );
  XOR U33433 ( .A(n32341), .B(o[341]), .Z(n32310) );
  XOR U33434 ( .A(n32311), .B(n32310), .Z(n32286) );
  AND U33435 ( .A(y[8003]), .B(x[498]), .Z(n32179) );
  NAND U33436 ( .A(y[8011]), .B(x[490]), .Z(n32178) );
  XNOR U33437 ( .A(n32179), .B(n32178), .Z(n32349) );
  NAND U33438 ( .A(x[481]), .B(y[8020]), .Z(n32350) );
  XOR U33439 ( .A(n32286), .B(n32285), .Z(n32287) );
  XOR U33440 ( .A(n32288), .B(n32287), .Z(n32291) );
  XOR U33441 ( .A(n32292), .B(n32291), .Z(n32294) );
  AND U33442 ( .A(x[487]), .B(y[8014]), .Z(n32586) );
  AND U33443 ( .A(y[8015]), .B(x[486]), .Z(n32181) );
  NAND U33444 ( .A(y[8007]), .B(x[494]), .Z(n32180) );
  XOR U33445 ( .A(n32181), .B(n32180), .Z(n32353) );
  NAND U33446 ( .A(x[489]), .B(y[8012]), .Z(n32298) );
  NAND U33447 ( .A(x[488]), .B(y[8013]), .Z(n32297) );
  XOR U33448 ( .A(n32298), .B(n32297), .Z(n32299) );
  AND U33449 ( .A(y[8009]), .B(x[492]), .Z(n32183) );
  NAND U33450 ( .A(y[8004]), .B(x[497]), .Z(n32182) );
  XNOR U33451 ( .A(n32183), .B(n32182), .Z(n32303) );
  NAND U33452 ( .A(x[482]), .B(y[8019]), .Z(n32304) );
  AND U33453 ( .A(y[8008]), .B(x[493]), .Z(n32185) );
  NAND U33454 ( .A(y[8018]), .B(x[483]), .Z(n32184) );
  XNOR U33455 ( .A(n32185), .B(n32184), .Z(n32338) );
  AND U33456 ( .A(x[484]), .B(y[8017]), .Z(n32337) );
  XOR U33457 ( .A(n32338), .B(n32337), .Z(n32314) );
  XOR U33458 ( .A(n32315), .B(n32314), .Z(n32316) );
  NAND U33459 ( .A(n32327), .B(n32186), .Z(n32190) );
  NAND U33460 ( .A(n32188), .B(n32187), .Z(n32189) );
  NAND U33461 ( .A(n32190), .B(n32189), .Z(n32280) );
  NAND U33462 ( .A(n32192), .B(n32191), .Z(n32196) );
  NAND U33463 ( .A(n32194), .B(n32193), .Z(n32195) );
  NAND U33464 ( .A(n32196), .B(n32195), .Z(n32279) );
  XOR U33465 ( .A(n32280), .B(n32279), .Z(n32281) );
  XOR U33466 ( .A(n32282), .B(n32281), .Z(n32293) );
  XOR U33467 ( .A(n32294), .B(n32293), .Z(n32256) );
  NAND U33468 ( .A(n32198), .B(n32197), .Z(n32202) );
  NAND U33469 ( .A(n32200), .B(n32199), .Z(n32201) );
  NAND U33470 ( .A(n32202), .B(n32201), .Z(n32263) );
  NAND U33471 ( .A(n32204), .B(n32203), .Z(n32208) );
  NAND U33472 ( .A(n32206), .B(n32205), .Z(n32207) );
  NAND U33473 ( .A(n32208), .B(n32207), .Z(n32262) );
  NAND U33474 ( .A(n32210), .B(n32209), .Z(n32214) );
  NAND U33475 ( .A(n32212), .B(n32211), .Z(n32213) );
  NAND U33476 ( .A(n32214), .B(n32213), .Z(n32261) );
  XOR U33477 ( .A(n32262), .B(n32261), .Z(n32264) );
  XOR U33478 ( .A(n32263), .B(n32264), .Z(n32255) );
  XOR U33479 ( .A(n32256), .B(n32255), .Z(n32257) );
  XOR U33480 ( .A(n32258), .B(n32257), .Z(n32244) );
  NAND U33481 ( .A(n32216), .B(n32215), .Z(n32220) );
  NANDN U33482 ( .A(n32218), .B(n32217), .Z(n32219) );
  NAND U33483 ( .A(n32220), .B(n32219), .Z(n32243) );
  XOR U33484 ( .A(n32245), .B(n32246), .Z(n32367) );
  NAND U33485 ( .A(n32222), .B(n32221), .Z(n32226) );
  NAND U33486 ( .A(n32224), .B(n32223), .Z(n32225) );
  NAND U33487 ( .A(n32226), .B(n32225), .Z(n32366) );
  NANDN U33488 ( .A(n32228), .B(n32227), .Z(n32232) );
  NAND U33489 ( .A(n32230), .B(n32229), .Z(n32231) );
  AND U33490 ( .A(n32232), .B(n32231), .Z(n32365) );
  XOR U33491 ( .A(n32366), .B(n32365), .Z(n32368) );
  XNOR U33492 ( .A(n32367), .B(n32368), .Z(n32361) );
  NAND U33493 ( .A(n32237), .B(n32236), .Z(n32241) );
  NANDN U33494 ( .A(n32239), .B(n32238), .Z(n32240) );
  AND U33495 ( .A(n32241), .B(n32240), .Z(n32359) );
  IV U33496 ( .A(n32359), .Z(n32358) );
  XOR U33497 ( .A(n32360), .B(n32358), .Z(n32242) );
  XNOR U33498 ( .A(n32361), .B(n32242), .Z(N694) );
  NANDN U33499 ( .A(n32244), .B(n32243), .Z(n32248) );
  NANDN U33500 ( .A(n32246), .B(n32245), .Z(n32247) );
  AND U33501 ( .A(n32248), .B(n32247), .Z(n32501) );
  NANDN U33502 ( .A(n32250), .B(n32249), .Z(n32254) );
  NAND U33503 ( .A(n32252), .B(n32251), .Z(n32253) );
  NAND U33504 ( .A(n32254), .B(n32253), .Z(n32499) );
  NAND U33505 ( .A(n32256), .B(n32255), .Z(n32260) );
  NAND U33506 ( .A(n32258), .B(n32257), .Z(n32259) );
  NAND U33507 ( .A(n32260), .B(n32259), .Z(n32373) );
  NAND U33508 ( .A(n32262), .B(n32261), .Z(n32266) );
  NAND U33509 ( .A(n32264), .B(n32263), .Z(n32265) );
  NAND U33510 ( .A(n32266), .B(n32265), .Z(n32372) );
  XOR U33511 ( .A(n32373), .B(n32372), .Z(n32375) );
  NAND U33512 ( .A(n32268), .B(n32267), .Z(n32272) );
  NAND U33513 ( .A(n32270), .B(n32269), .Z(n32271) );
  NAND U33514 ( .A(n32272), .B(n32271), .Z(n32379) );
  NANDN U33515 ( .A(n32274), .B(n32273), .Z(n32278) );
  NAND U33516 ( .A(n32276), .B(n32275), .Z(n32277) );
  AND U33517 ( .A(n32278), .B(n32277), .Z(n32387) );
  NAND U33518 ( .A(n32280), .B(n32279), .Z(n32284) );
  NAND U33519 ( .A(n32282), .B(n32281), .Z(n32283) );
  AND U33520 ( .A(n32284), .B(n32283), .Z(n32385) );
  NAND U33521 ( .A(n32286), .B(n32285), .Z(n32290) );
  NAND U33522 ( .A(n32288), .B(n32287), .Z(n32289) );
  NAND U33523 ( .A(n32290), .B(n32289), .Z(n32384) );
  XOR U33524 ( .A(n32379), .B(n32378), .Z(n32381) );
  NAND U33525 ( .A(n32292), .B(n32291), .Z(n32296) );
  NAND U33526 ( .A(n32294), .B(n32293), .Z(n32295) );
  AND U33527 ( .A(n32296), .B(n32295), .Z(n32489) );
  NAND U33528 ( .A(n32298), .B(n32297), .Z(n32302) );
  NANDN U33529 ( .A(n32300), .B(n32299), .Z(n32301) );
  AND U33530 ( .A(n32302), .B(n32301), .Z(n32483) );
  NANDN U33531 ( .A(n32989), .B(n32434), .Z(n32306) );
  NANDN U33532 ( .A(n32304), .B(n32303), .Z(n32305) );
  AND U33533 ( .A(n32306), .B(n32305), .Z(n32411) );
  AND U33534 ( .A(x[485]), .B(y[8017]), .Z(n32456) );
  NAND U33535 ( .A(x[497]), .B(y[8005]), .Z(n32457) );
  NAND U33536 ( .A(x[496]), .B(y[8006]), .Z(n32459) );
  AND U33537 ( .A(y[8004]), .B(x[498]), .Z(n32308) );
  NAND U33538 ( .A(y[8010]), .B(x[492]), .Z(n32307) );
  XNOR U33539 ( .A(n32308), .B(n32307), .Z(n32435) );
  NAND U33540 ( .A(x[484]), .B(y[8018]), .Z(n32436) );
  XOR U33541 ( .A(n32409), .B(n32408), .Z(n32410) );
  NAND U33542 ( .A(x[499]), .B(y[8010]), .Z(n33499) );
  NANDN U33543 ( .A(n33499), .B(n32309), .Z(n32313) );
  NAND U33544 ( .A(n32311), .B(n32310), .Z(n32312) );
  AND U33545 ( .A(n32313), .B(n32312), .Z(n32481) );
  XOR U33546 ( .A(n32480), .B(n32481), .Z(n32482) );
  NAND U33547 ( .A(n32315), .B(n32314), .Z(n32319) );
  NANDN U33548 ( .A(n32317), .B(n32316), .Z(n32318) );
  AND U33549 ( .A(n32319), .B(n32318), .Z(n32469) );
  NAND U33550 ( .A(n32321), .B(n32320), .Z(n32325) );
  NAND U33551 ( .A(n32323), .B(n32322), .Z(n32324) );
  NAND U33552 ( .A(n32325), .B(n32324), .Z(n32468) );
  NAND U33553 ( .A(n32327), .B(n32326), .Z(n32331) );
  AND U33554 ( .A(n32329), .B(n32328), .Z(n32330) );
  ANDN U33555 ( .B(n32331), .A(n32330), .Z(n32431) );
  AND U33556 ( .A(y[8009]), .B(x[493]), .Z(n32333) );
  NAND U33557 ( .A(y[8002]), .B(x[500]), .Z(n32332) );
  XNOR U33558 ( .A(n32333), .B(n32332), .Z(n32452) );
  NAND U33559 ( .A(x[482]), .B(y[8020]), .Z(n32453) );
  AND U33560 ( .A(y[8016]), .B(x[486]), .Z(n32335) );
  NAND U33561 ( .A(y[8007]), .B(x[495]), .Z(n32334) );
  XNOR U33562 ( .A(n32335), .B(n32334), .Z(n32464) );
  XOR U33563 ( .A(n32429), .B(n32428), .Z(n32430) );
  AND U33564 ( .A(x[493]), .B(y[8018]), .Z(n33786) );
  NANDN U33565 ( .A(n32336), .B(n33786), .Z(n32340) );
  NAND U33566 ( .A(n32338), .B(n32337), .Z(n32339) );
  AND U33567 ( .A(n32340), .B(n32339), .Z(n32399) );
  AND U33568 ( .A(x[481]), .B(y[8021]), .Z(n32422) );
  XOR U33569 ( .A(n32423), .B(n32422), .Z(n32421) );
  AND U33570 ( .A(n32341), .B(o[341]), .Z(n32420) );
  XOR U33571 ( .A(n32421), .B(n32420), .Z(n32397) );
  AND U33572 ( .A(x[494]), .B(y[8008]), .Z(n32414) );
  AND U33573 ( .A(x[483]), .B(y[8019]), .Z(n32415) );
  XOR U33574 ( .A(n32414), .B(n32415), .Z(n32416) );
  AND U33575 ( .A(x[499]), .B(y[8003]), .Z(n32417) );
  XOR U33576 ( .A(n32416), .B(n32417), .Z(n32396) );
  XOR U33577 ( .A(n32397), .B(n32396), .Z(n32398) );
  XOR U33578 ( .A(n32475), .B(n32474), .Z(n32477) );
  NANDN U33579 ( .A(n32343), .B(n32342), .Z(n32347) );
  NAND U33580 ( .A(n32345), .B(n32344), .Z(n32346) );
  AND U33581 ( .A(n32347), .B(n32346), .Z(n32391) );
  AND U33582 ( .A(x[498]), .B(y[8011]), .Z(n33501) );
  NAND U33583 ( .A(n33501), .B(n32348), .Z(n32352) );
  NANDN U33584 ( .A(n32350), .B(n32349), .Z(n32351) );
  NAND U33585 ( .A(n32352), .B(n32351), .Z(n32390) );
  AND U33586 ( .A(x[494]), .B(y[8015]), .Z(n33535) );
  NAND U33587 ( .A(n33535), .B(n32463), .Z(n32355) );
  NANDN U33588 ( .A(n32353), .B(n32586), .Z(n32354) );
  NAND U33589 ( .A(n32355), .B(n32354), .Z(n32404) );
  AND U33590 ( .A(x[480]), .B(y[8022]), .Z(n32439) );
  NAND U33591 ( .A(x[502]), .B(y[8000]), .Z(n32440) );
  AND U33592 ( .A(x[501]), .B(y[8001]), .Z(n32462) );
  XOR U33593 ( .A(o[342]), .B(n32462), .Z(n32441) );
  XOR U33594 ( .A(n32442), .B(n32441), .Z(n32403) );
  AND U33595 ( .A(y[8015]), .B(x[487]), .Z(n32357) );
  NAND U33596 ( .A(y[8014]), .B(x[488]), .Z(n32356) );
  XNOR U33597 ( .A(n32357), .B(n32356), .Z(n32446) );
  XOR U33598 ( .A(n32446), .B(n32445), .Z(n32402) );
  XOR U33599 ( .A(n32403), .B(n32402), .Z(n32405) );
  XOR U33600 ( .A(n32404), .B(n32405), .Z(n32392) );
  XOR U33601 ( .A(n32393), .B(n32392), .Z(n32476) );
  XOR U33602 ( .A(n32477), .B(n32476), .Z(n32470) );
  XOR U33603 ( .A(n32471), .B(n32470), .Z(n32487) );
  XOR U33604 ( .A(n32486), .B(n32487), .Z(n32488) );
  XOR U33605 ( .A(n32381), .B(n32380), .Z(n32374) );
  XOR U33606 ( .A(n32375), .B(n32374), .Z(n32500) );
  XNOR U33607 ( .A(n32499), .B(n32500), .Z(n32502) );
  OR U33608 ( .A(n32360), .B(n32358), .Z(n32364) );
  ANDN U33609 ( .B(n32360), .A(n32359), .Z(n32362) );
  OR U33610 ( .A(n32362), .B(n32361), .Z(n32363) );
  AND U33611 ( .A(n32364), .B(n32363), .Z(n32493) );
  NAND U33612 ( .A(n32366), .B(n32365), .Z(n32370) );
  NAND U33613 ( .A(n32368), .B(n32367), .Z(n32369) );
  AND U33614 ( .A(n32370), .B(n32369), .Z(n32494) );
  IV U33615 ( .A(n32494), .Z(n32492) );
  XOR U33616 ( .A(n32493), .B(n32492), .Z(n32371) );
  XNOR U33617 ( .A(n32495), .B(n32371), .Z(N695) );
  NAND U33618 ( .A(n32373), .B(n32372), .Z(n32377) );
  NAND U33619 ( .A(n32375), .B(n32374), .Z(n32376) );
  AND U33620 ( .A(n32377), .B(n32376), .Z(n32643) );
  NAND U33621 ( .A(n32379), .B(n32378), .Z(n32383) );
  NAND U33622 ( .A(n32381), .B(n32380), .Z(n32382) );
  AND U33623 ( .A(n32383), .B(n32382), .Z(n32641) );
  NANDN U33624 ( .A(n32385), .B(n32384), .Z(n32389) );
  NANDN U33625 ( .A(n32387), .B(n32386), .Z(n32388) );
  AND U33626 ( .A(n32389), .B(n32388), .Z(n32622) );
  NANDN U33627 ( .A(n32391), .B(n32390), .Z(n32395) );
  NAND U33628 ( .A(n32393), .B(n32392), .Z(n32394) );
  NAND U33629 ( .A(n32395), .B(n32394), .Z(n32568) );
  NAND U33630 ( .A(n32397), .B(n32396), .Z(n32401) );
  NANDN U33631 ( .A(n32399), .B(n32398), .Z(n32400) );
  NAND U33632 ( .A(n32401), .B(n32400), .Z(n32567) );
  NAND U33633 ( .A(n32403), .B(n32402), .Z(n32407) );
  NAND U33634 ( .A(n32405), .B(n32404), .Z(n32406) );
  NAND U33635 ( .A(n32407), .B(n32406), .Z(n32566) );
  XOR U33636 ( .A(n32567), .B(n32566), .Z(n32569) );
  XOR U33637 ( .A(n32568), .B(n32569), .Z(n32633) );
  NAND U33638 ( .A(n32409), .B(n32408), .Z(n32413) );
  NANDN U33639 ( .A(n32411), .B(n32410), .Z(n32412) );
  NAND U33640 ( .A(n32413), .B(n32412), .Z(n32631) );
  NAND U33641 ( .A(n32415), .B(n32414), .Z(n32419) );
  NAND U33642 ( .A(n32417), .B(n32416), .Z(n32418) );
  NAND U33643 ( .A(n32419), .B(n32418), .Z(n32513) );
  AND U33644 ( .A(n32421), .B(n32420), .Z(n32425) );
  NAND U33645 ( .A(n32423), .B(n32422), .Z(n32424) );
  NANDN U33646 ( .A(n32425), .B(n32424), .Z(n32512) );
  XOR U33647 ( .A(n32513), .B(n32512), .Z(n32515) );
  AND U33648 ( .A(y[8016]), .B(x[487]), .Z(n32427) );
  NAND U33649 ( .A(y[8014]), .B(x[489]), .Z(n32426) );
  XNOR U33650 ( .A(n32427), .B(n32426), .Z(n32587) );
  AND U33651 ( .A(x[490]), .B(y[8013]), .Z(n32519) );
  XOR U33652 ( .A(n32518), .B(n32519), .Z(n32521) );
  AND U33653 ( .A(x[486]), .B(y[8017]), .Z(n32578) );
  AND U33654 ( .A(x[495]), .B(y[8008]), .Z(n32579) );
  XOR U33655 ( .A(n32578), .B(n32579), .Z(n32580) );
  AND U33656 ( .A(x[491]), .B(y[8012]), .Z(n32581) );
  XOR U33657 ( .A(n32580), .B(n32581), .Z(n32520) );
  XOR U33658 ( .A(n32521), .B(n32520), .Z(n32514) );
  XOR U33659 ( .A(n32515), .B(n32514), .Z(n32632) );
  XNOR U33660 ( .A(n32631), .B(n32632), .Z(n32634) );
  NAND U33661 ( .A(n32429), .B(n32428), .Z(n32433) );
  NANDN U33662 ( .A(n32431), .B(n32430), .Z(n32432) );
  AND U33663 ( .A(n32433), .B(n32432), .Z(n32614) );
  AND U33664 ( .A(x[498]), .B(y[8010]), .Z(n33348) );
  NAND U33665 ( .A(n33348), .B(n32434), .Z(n32438) );
  NANDN U33666 ( .A(n32436), .B(n32435), .Z(n32437) );
  NAND U33667 ( .A(n32438), .B(n32437), .Z(n32543) );
  NANDN U33668 ( .A(n32440), .B(n32439), .Z(n32444) );
  NAND U33669 ( .A(n32442), .B(n32441), .Z(n32443) );
  NAND U33670 ( .A(n32444), .B(n32443), .Z(n32542) );
  XOR U33671 ( .A(n32543), .B(n32542), .Z(n32544) );
  NANDN U33672 ( .A(n32588), .B(n32586), .Z(n32448) );
  NAND U33673 ( .A(n32446), .B(n32445), .Z(n32447) );
  NAND U33674 ( .A(n32448), .B(n32447), .Z(n32556) );
  AND U33675 ( .A(x[480]), .B(y[8023]), .Z(n32597) );
  AND U33676 ( .A(x[503]), .B(y[8000]), .Z(n32598) );
  XOR U33677 ( .A(n32597), .B(n32598), .Z(n32600) );
  AND U33678 ( .A(x[502]), .B(y[8001]), .Z(n32577) );
  XOR U33679 ( .A(o[343]), .B(n32577), .Z(n32599) );
  XOR U33680 ( .A(n32600), .B(n32599), .Z(n32555) );
  NAND U33681 ( .A(y[8003]), .B(x[500]), .Z(n32449) );
  XNOR U33682 ( .A(n32450), .B(n32449), .Z(n32573) );
  AND U33683 ( .A(x[499]), .B(y[8004]), .Z(n32574) );
  XOR U33684 ( .A(n32573), .B(n32574), .Z(n32554) );
  XOR U33685 ( .A(n32555), .B(n32554), .Z(n32557) );
  XNOR U33686 ( .A(n32556), .B(n32557), .Z(n32545) );
  NAND U33687 ( .A(x[500]), .B(y[8009]), .Z(n33547) );
  AND U33688 ( .A(x[493]), .B(y[8002]), .Z(n32451) );
  NANDN U33689 ( .A(n33547), .B(n32451), .Z(n32455) );
  NANDN U33690 ( .A(n32453), .B(n32452), .Z(n32454) );
  AND U33691 ( .A(n32455), .B(n32454), .Z(n32608) );
  NANDN U33692 ( .A(n32457), .B(n32456), .Z(n32461) );
  NANDN U33693 ( .A(n32459), .B(n32458), .Z(n32460) );
  NAND U33694 ( .A(n32461), .B(n32460), .Z(n32562) );
  AND U33695 ( .A(x[493]), .B(y[8010]), .Z(n32536) );
  AND U33696 ( .A(x[482]), .B(y[8021]), .Z(n32537) );
  XOR U33697 ( .A(n32536), .B(n32537), .Z(n32538) );
  AND U33698 ( .A(x[501]), .B(y[8002]), .Z(n32539) );
  XOR U33699 ( .A(n32538), .B(n32539), .Z(n32561) );
  AND U33700 ( .A(x[492]), .B(y[8011]), .Z(n32591) );
  AND U33701 ( .A(x[481]), .B(y[8022]), .Z(n32592) );
  XOR U33702 ( .A(n32591), .B(n32592), .Z(n32594) );
  AND U33703 ( .A(o[342]), .B(n32462), .Z(n32593) );
  XOR U33704 ( .A(n32594), .B(n32593), .Z(n32560) );
  XOR U33705 ( .A(n32561), .B(n32560), .Z(n32563) );
  XOR U33706 ( .A(n32562), .B(n32563), .Z(n32607) );
  AND U33707 ( .A(x[495]), .B(y[8016]), .Z(n33774) );
  NAND U33708 ( .A(n33774), .B(n32463), .Z(n32467) );
  NANDN U33709 ( .A(n32465), .B(n32464), .Z(n32466) );
  NAND U33710 ( .A(n32467), .B(n32466), .Z(n32550) );
  AND U33711 ( .A(x[494]), .B(y[8009]), .Z(n32530) );
  AND U33712 ( .A(x[483]), .B(y[8020]), .Z(n32531) );
  XOR U33713 ( .A(n32530), .B(n32531), .Z(n32532) );
  AND U33714 ( .A(x[484]), .B(y[8019]), .Z(n32533) );
  XOR U33715 ( .A(n32532), .B(n32533), .Z(n32549) );
  AND U33716 ( .A(x[485]), .B(y[8018]), .Z(n32524) );
  AND U33717 ( .A(x[498]), .B(y[8005]), .Z(n32525) );
  XOR U33718 ( .A(n32524), .B(n32525), .Z(n32527) );
  AND U33719 ( .A(x[497]), .B(y[8006]), .Z(n32526) );
  XOR U33720 ( .A(n32527), .B(n32526), .Z(n32548) );
  XOR U33721 ( .A(n32549), .B(n32548), .Z(n32551) );
  XOR U33722 ( .A(n32550), .B(n32551), .Z(n32609) );
  XOR U33723 ( .A(n32610), .B(n32609), .Z(n32615) );
  XOR U33724 ( .A(n32616), .B(n32615), .Z(n32619) );
  XOR U33725 ( .A(n32620), .B(n32619), .Z(n32621) );
  NANDN U33726 ( .A(n32469), .B(n32468), .Z(n32473) );
  NAND U33727 ( .A(n32471), .B(n32470), .Z(n32472) );
  AND U33728 ( .A(n32473), .B(n32472), .Z(n32628) );
  NAND U33729 ( .A(n32475), .B(n32474), .Z(n32479) );
  NAND U33730 ( .A(n32477), .B(n32476), .Z(n32478) );
  AND U33731 ( .A(n32479), .B(n32478), .Z(n32626) );
  NAND U33732 ( .A(n32481), .B(n32480), .Z(n32485) );
  NANDN U33733 ( .A(n32483), .B(n32482), .Z(n32484) );
  AND U33734 ( .A(n32485), .B(n32484), .Z(n32625) );
  NAND U33735 ( .A(n32487), .B(n32486), .Z(n32491) );
  NANDN U33736 ( .A(n32489), .B(n32488), .Z(n32490) );
  AND U33737 ( .A(n32491), .B(n32490), .Z(n32507) );
  XOR U33738 ( .A(n32506), .B(n32507), .Z(n32509) );
  XOR U33739 ( .A(n32508), .B(n32509), .Z(n32640) );
  XOR U33740 ( .A(n32641), .B(n32640), .Z(n32642) );
  XNOR U33741 ( .A(n32643), .B(n32642), .Z(n32639) );
  NANDN U33742 ( .A(n32492), .B(n32493), .Z(n32498) );
  NOR U33743 ( .A(n32494), .B(n32493), .Z(n32496) );
  OR U33744 ( .A(n32496), .B(n32495), .Z(n32497) );
  AND U33745 ( .A(n32498), .B(n32497), .Z(n32638) );
  NAND U33746 ( .A(n32500), .B(n32499), .Z(n32504) );
  NANDN U33747 ( .A(n32502), .B(n32501), .Z(n32503) );
  AND U33748 ( .A(n32504), .B(n32503), .Z(n32637) );
  XOR U33749 ( .A(n32638), .B(n32637), .Z(n32505) );
  XNOR U33750 ( .A(n32639), .B(n32505), .Z(N696) );
  NAND U33751 ( .A(n32507), .B(n32506), .Z(n32511) );
  NAND U33752 ( .A(n32509), .B(n32508), .Z(n32510) );
  AND U33753 ( .A(n32511), .B(n32510), .Z(n32650) );
  NAND U33754 ( .A(n32513), .B(n32512), .Z(n32517) );
  NAND U33755 ( .A(n32515), .B(n32514), .Z(n32516) );
  NAND U33756 ( .A(n32517), .B(n32516), .Z(n32731) );
  NAND U33757 ( .A(n32519), .B(n32518), .Z(n32523) );
  NAND U33758 ( .A(n32521), .B(n32520), .Z(n32522) );
  NAND U33759 ( .A(n32523), .B(n32522), .Z(n32729) );
  NAND U33760 ( .A(n32525), .B(n32524), .Z(n32529) );
  NAND U33761 ( .A(n32527), .B(n32526), .Z(n32528) );
  NAND U33762 ( .A(n32529), .B(n32528), .Z(n32755) );
  AND U33763 ( .A(x[480]), .B(y[8024]), .Z(n32711) );
  AND U33764 ( .A(x[504]), .B(y[8000]), .Z(n32710) );
  XOR U33765 ( .A(n32711), .B(n32710), .Z(n32713) );
  AND U33766 ( .A(x[503]), .B(y[8001]), .Z(n32703) );
  XOR U33767 ( .A(n32703), .B(o[344]), .Z(n32712) );
  XOR U33768 ( .A(n32713), .B(n32712), .Z(n32753) );
  AND U33769 ( .A(x[487]), .B(y[8017]), .Z(n32696) );
  AND U33770 ( .A(x[498]), .B(y[8006]), .Z(n32697) );
  XOR U33771 ( .A(n32696), .B(n32697), .Z(n32698) );
  AND U33772 ( .A(x[497]), .B(y[8007]), .Z(n32699) );
  XOR U33773 ( .A(n32698), .B(n32699), .Z(n32752) );
  XOR U33774 ( .A(n32753), .B(n32752), .Z(n32754) );
  XOR U33775 ( .A(n32755), .B(n32754), .Z(n32743) );
  NAND U33776 ( .A(n32531), .B(n32530), .Z(n32535) );
  NAND U33777 ( .A(n32533), .B(n32532), .Z(n32534) );
  NAND U33778 ( .A(n32535), .B(n32534), .Z(n32741) );
  NAND U33779 ( .A(n32537), .B(n32536), .Z(n32541) );
  NAND U33780 ( .A(n32539), .B(n32538), .Z(n32540) );
  NAND U33781 ( .A(n32541), .B(n32540), .Z(n32740) );
  XOR U33782 ( .A(n32741), .B(n32740), .Z(n32742) );
  XOR U33783 ( .A(n32743), .B(n32742), .Z(n32728) );
  XOR U33784 ( .A(n32729), .B(n32728), .Z(n32730) );
  XNOR U33785 ( .A(n32731), .B(n32730), .Z(n32736) );
  NAND U33786 ( .A(n32543), .B(n32542), .Z(n32547) );
  NANDN U33787 ( .A(n32545), .B(n32544), .Z(n32546) );
  AND U33788 ( .A(n32547), .B(n32546), .Z(n32784) );
  NAND U33789 ( .A(n32549), .B(n32548), .Z(n32553) );
  NAND U33790 ( .A(n32551), .B(n32550), .Z(n32552) );
  AND U33791 ( .A(n32553), .B(n32552), .Z(n32782) );
  NAND U33792 ( .A(n32555), .B(n32554), .Z(n32559) );
  NAND U33793 ( .A(n32557), .B(n32556), .Z(n32558) );
  AND U33794 ( .A(n32559), .B(n32558), .Z(n32781) );
  XOR U33795 ( .A(n32782), .B(n32781), .Z(n32783) );
  XOR U33796 ( .A(n32784), .B(n32783), .Z(n32734) );
  NAND U33797 ( .A(n32561), .B(n32560), .Z(n32565) );
  NAND U33798 ( .A(n32563), .B(n32562), .Z(n32564) );
  NAND U33799 ( .A(n32565), .B(n32564), .Z(n32735) );
  XOR U33800 ( .A(n32736), .B(n32737), .Z(n32663) );
  NAND U33801 ( .A(n32567), .B(n32566), .Z(n32571) );
  NAND U33802 ( .A(n32569), .B(n32568), .Z(n32570) );
  AND U33803 ( .A(n32571), .B(n32570), .Z(n32662) );
  XOR U33804 ( .A(n32663), .B(n32662), .Z(n32665) );
  AND U33805 ( .A(x[500]), .B(y[8007]), .Z(n32572) );
  NAND U33806 ( .A(n32572), .B(n32758), .Z(n32576) );
  NAND U33807 ( .A(n32574), .B(n32573), .Z(n32575) );
  NAND U33808 ( .A(n32576), .B(n32575), .Z(n32778) );
  AND U33809 ( .A(x[502]), .B(y[8002]), .Z(n32684) );
  XOR U33810 ( .A(n32685), .B(n32684), .Z(n32686) );
  AND U33811 ( .A(x[482]), .B(y[8022]), .Z(n32687) );
  XOR U33812 ( .A(n32686), .B(n32687), .Z(n32776) );
  AND U33813 ( .A(x[481]), .B(y[8023]), .Z(n32692) );
  XOR U33814 ( .A(n32693), .B(n32692), .Z(n32691) );
  AND U33815 ( .A(o[343]), .B(n32577), .Z(n32690) );
  XOR U33816 ( .A(n32691), .B(n32690), .Z(n32775) );
  XOR U33817 ( .A(n32776), .B(n32775), .Z(n32777) );
  XOR U33818 ( .A(n32778), .B(n32777), .Z(n32723) );
  NAND U33819 ( .A(n32579), .B(n32578), .Z(n32583) );
  NAND U33820 ( .A(n32581), .B(n32580), .Z(n32582) );
  NAND U33821 ( .A(n32583), .B(n32582), .Z(n32772) );
  AND U33822 ( .A(y[8008]), .B(x[496]), .Z(n32585) );
  NAND U33823 ( .A(y[8003]), .B(x[501]), .Z(n32584) );
  XNOR U33824 ( .A(n32585), .B(n32584), .Z(n32759) );
  AND U33825 ( .A(x[485]), .B(y[8019]), .Z(n32760) );
  XOR U33826 ( .A(n32759), .B(n32760), .Z(n32770) );
  AND U33827 ( .A(x[486]), .B(y[8018]), .Z(n33080) );
  AND U33828 ( .A(x[500]), .B(y[8004]), .Z(n32887) );
  XOR U33829 ( .A(n33080), .B(n32887), .Z(n32765) );
  AND U33830 ( .A(x[499]), .B(y[8005]), .Z(n32766) );
  XOR U33831 ( .A(n32765), .B(n32766), .Z(n32769) );
  XOR U33832 ( .A(n32770), .B(n32769), .Z(n32771) );
  XOR U33833 ( .A(n32772), .B(n32771), .Z(n32749) );
  NANDN U33834 ( .A(n32812), .B(n32586), .Z(n32590) );
  NANDN U33835 ( .A(n32588), .B(n32587), .Z(n32589) );
  NAND U33836 ( .A(n32590), .B(n32589), .Z(n32747) );
  NAND U33837 ( .A(n32592), .B(n32591), .Z(n32596) );
  NAND U33838 ( .A(n32594), .B(n32593), .Z(n32595) );
  NAND U33839 ( .A(n32596), .B(n32595), .Z(n32746) );
  XOR U33840 ( .A(n32747), .B(n32746), .Z(n32748) );
  XOR U33841 ( .A(n32749), .B(n32748), .Z(n32722) );
  XOR U33842 ( .A(n32723), .B(n32722), .Z(n32725) );
  NAND U33843 ( .A(n32598), .B(n32597), .Z(n32602) );
  NAND U33844 ( .A(n32600), .B(n32599), .Z(n32601) );
  NAND U33845 ( .A(n32602), .B(n32601), .Z(n32717) );
  AND U33846 ( .A(x[483]), .B(y[8021]), .Z(n32706) );
  XOR U33847 ( .A(n32707), .B(n32706), .Z(n32705) );
  AND U33848 ( .A(x[484]), .B(y[8020]), .Z(n32704) );
  XOR U33849 ( .A(n32705), .B(n32704), .Z(n32716) );
  XOR U33850 ( .A(n32717), .B(n32716), .Z(n32719) );
  AND U33851 ( .A(y[8015]), .B(x[489]), .Z(n32604) );
  NAND U33852 ( .A(y[8014]), .B(x[490]), .Z(n32603) );
  XNOR U33853 ( .A(n32604), .B(n32603), .Z(n32676) );
  AND U33854 ( .A(y[8010]), .B(x[494]), .Z(n32606) );
  NAND U33855 ( .A(y[8016]), .B(x[488]), .Z(n32605) );
  XNOR U33856 ( .A(n32606), .B(n32605), .Z(n32680) );
  NAND U33857 ( .A(x[491]), .B(y[8013]), .Z(n32681) );
  XOR U33858 ( .A(n32676), .B(n32675), .Z(n32718) );
  XOR U33859 ( .A(n32719), .B(n32718), .Z(n32724) );
  XOR U33860 ( .A(n32725), .B(n32724), .Z(n32669) );
  NANDN U33861 ( .A(n32608), .B(n32607), .Z(n32612) );
  NAND U33862 ( .A(n32610), .B(n32609), .Z(n32611) );
  AND U33863 ( .A(n32612), .B(n32611), .Z(n32668) );
  NANDN U33864 ( .A(n32614), .B(n32613), .Z(n32618) );
  NAND U33865 ( .A(n32616), .B(n32615), .Z(n32617) );
  NAND U33866 ( .A(n32618), .B(n32617), .Z(n32671) );
  XOR U33867 ( .A(n32665), .B(n32664), .Z(n32648) );
  NAND U33868 ( .A(n32620), .B(n32619), .Z(n32624) );
  NANDN U33869 ( .A(n32622), .B(n32621), .Z(n32623) );
  NAND U33870 ( .A(n32624), .B(n32623), .Z(n32658) );
  NANDN U33871 ( .A(n32626), .B(n32625), .Z(n32630) );
  NANDN U33872 ( .A(n32628), .B(n32627), .Z(n32629) );
  NAND U33873 ( .A(n32630), .B(n32629), .Z(n32657) );
  NAND U33874 ( .A(n32632), .B(n32631), .Z(n32636) );
  NANDN U33875 ( .A(n32634), .B(n32633), .Z(n32635) );
  NAND U33876 ( .A(n32636), .B(n32635), .Z(n32656) );
  XOR U33877 ( .A(n32657), .B(n32656), .Z(n32659) );
  XOR U33878 ( .A(n32658), .B(n32659), .Z(n32647) );
  XNOR U33879 ( .A(n32650), .B(n32649), .Z(n32655) );
  NAND U33880 ( .A(n32641), .B(n32640), .Z(n32645) );
  NAND U33881 ( .A(n32643), .B(n32642), .Z(n32644) );
  AND U33882 ( .A(n32645), .B(n32644), .Z(n32654) );
  XOR U33883 ( .A(n32653), .B(n32654), .Z(n32646) );
  XNOR U33884 ( .A(n32655), .B(n32646), .Z(N697) );
  NANDN U33885 ( .A(n32648), .B(n32647), .Z(n32652) );
  NAND U33886 ( .A(n32650), .B(n32649), .Z(n32651) );
  NAND U33887 ( .A(n32652), .B(n32651), .Z(n32930) );
  IV U33888 ( .A(n32930), .Z(n32929) );
  NAND U33889 ( .A(n32657), .B(n32656), .Z(n32661) );
  NAND U33890 ( .A(n32659), .B(n32658), .Z(n32660) );
  AND U33891 ( .A(n32661), .B(n32660), .Z(n32938) );
  NAND U33892 ( .A(n32663), .B(n32662), .Z(n32667) );
  NAND U33893 ( .A(n32665), .B(n32664), .Z(n32666) );
  NAND U33894 ( .A(n32667), .B(n32666), .Z(n32936) );
  NANDN U33895 ( .A(n32669), .B(n32668), .Z(n32673) );
  NANDN U33896 ( .A(n32671), .B(n32670), .Z(n32672) );
  AND U33897 ( .A(n32673), .B(n32672), .Z(n32789) );
  NANDN U33898 ( .A(n32702), .B(n32674), .Z(n32678) );
  NAND U33899 ( .A(n32676), .B(n32675), .Z(n32677) );
  NAND U33900 ( .A(n32678), .B(n32677), .Z(n32837) );
  AND U33901 ( .A(x[494]), .B(y[8016]), .Z(n33699) );
  NAND U33902 ( .A(n33699), .B(n32679), .Z(n32683) );
  NANDN U33903 ( .A(n32681), .B(n32680), .Z(n32682) );
  NAND U33904 ( .A(n32683), .B(n32682), .Z(n32864) );
  NAND U33905 ( .A(x[491]), .B(y[8014]), .Z(n32883) );
  NAND U33906 ( .A(x[492]), .B(y[8013]), .Z(n32882) );
  NAND U33907 ( .A(x[487]), .B(y[8018]), .Z(n32881) );
  XOR U33908 ( .A(n32882), .B(n32881), .Z(n32884) );
  XOR U33909 ( .A(n32883), .B(n32884), .Z(n32863) );
  AND U33910 ( .A(x[504]), .B(y[8001]), .Z(n32880) );
  XOR U33911 ( .A(o[345]), .B(n32880), .Z(n32851) );
  AND U33912 ( .A(x[481]), .B(y[8024]), .Z(n32850) );
  XOR U33913 ( .A(n32851), .B(n32850), .Z(n32853) );
  AND U33914 ( .A(x[493]), .B(y[8012]), .Z(n32852) );
  XOR U33915 ( .A(n32853), .B(n32852), .Z(n32862) );
  XOR U33916 ( .A(n32864), .B(n32865), .Z(n32836) );
  XOR U33917 ( .A(n32837), .B(n32836), .Z(n32839) );
  AND U33918 ( .A(n32685), .B(n32684), .Z(n32689) );
  NAND U33919 ( .A(n32687), .B(n32686), .Z(n32688) );
  NANDN U33920 ( .A(n32689), .B(n32688), .Z(n32825) );
  AND U33921 ( .A(n32691), .B(n32690), .Z(n32695) );
  NAND U33922 ( .A(n32693), .B(n32692), .Z(n32694) );
  NANDN U33923 ( .A(n32695), .B(n32694), .Z(n32824) );
  XOR U33924 ( .A(n32825), .B(n32824), .Z(n32826) );
  NAND U33925 ( .A(n32697), .B(n32696), .Z(n32701) );
  NAND U33926 ( .A(n32699), .B(n32698), .Z(n32700) );
  NAND U33927 ( .A(n32701), .B(n32700), .Z(n32820) );
  NAND U33928 ( .A(x[488]), .B(y[8017]), .Z(n32814) );
  XOR U33929 ( .A(n32812), .B(n32702), .Z(n32815) );
  XNOR U33930 ( .A(n32814), .B(n32815), .Z(n32819) );
  NAND U33931 ( .A(n32703), .B(o[344]), .Z(n32808) );
  NAND U33932 ( .A(x[505]), .B(y[8000]), .Z(n32807) );
  NAND U33933 ( .A(x[480]), .B(y[8025]), .Z(n32806) );
  XOR U33934 ( .A(n32807), .B(n32806), .Z(n32809) );
  XNOR U33935 ( .A(n32808), .B(n32809), .Z(n32818) );
  XNOR U33936 ( .A(n32819), .B(n32818), .Z(n32821) );
  XOR U33937 ( .A(n32820), .B(n32821), .Z(n32827) );
  XNOR U33938 ( .A(n32826), .B(n32827), .Z(n32838) );
  XNOR U33939 ( .A(n32839), .B(n32838), .Z(n32926) );
  AND U33940 ( .A(n32705), .B(n32704), .Z(n32709) );
  NAND U33941 ( .A(n32707), .B(n32706), .Z(n32708) );
  NANDN U33942 ( .A(n32709), .B(n32708), .Z(n32902) );
  NAND U33943 ( .A(n32711), .B(n32710), .Z(n32715) );
  NAND U33944 ( .A(n32713), .B(n32712), .Z(n32714) );
  NAND U33945 ( .A(n32715), .B(n32714), .Z(n32900) );
  AND U33946 ( .A(x[494]), .B(y[8011]), .Z(n32857) );
  AND U33947 ( .A(x[482]), .B(y[8023]), .Z(n32856) );
  XOR U33948 ( .A(n32857), .B(n32856), .Z(n32859) );
  AND U33949 ( .A(x[483]), .B(y[8022]), .Z(n32858) );
  XOR U33950 ( .A(n32859), .B(n32858), .Z(n32899) );
  XOR U33951 ( .A(n32900), .B(n32899), .Z(n32901) );
  XNOR U33952 ( .A(n32902), .B(n32901), .Z(n32924) );
  NAND U33953 ( .A(n32717), .B(n32716), .Z(n32721) );
  NAND U33954 ( .A(n32719), .B(n32718), .Z(n32720) );
  AND U33955 ( .A(n32721), .B(n32720), .Z(n32923) );
  XOR U33956 ( .A(n32924), .B(n32923), .Z(n32925) );
  XOR U33957 ( .A(n32926), .B(n32925), .Z(n32917) );
  NAND U33958 ( .A(n32723), .B(n32722), .Z(n32727) );
  NAND U33959 ( .A(n32725), .B(n32724), .Z(n32726) );
  AND U33960 ( .A(n32727), .B(n32726), .Z(n32918) );
  XOR U33961 ( .A(n32917), .B(n32918), .Z(n32919) );
  NAND U33962 ( .A(n32729), .B(n32728), .Z(n32733) );
  NAND U33963 ( .A(n32731), .B(n32730), .Z(n32732) );
  AND U33964 ( .A(n32733), .B(n32732), .Z(n32920) );
  XOR U33965 ( .A(n32919), .B(n32920), .Z(n32788) );
  NANDN U33966 ( .A(n32735), .B(n32734), .Z(n32739) );
  NAND U33967 ( .A(n32737), .B(n32736), .Z(n32738) );
  NAND U33968 ( .A(n32739), .B(n32738), .Z(n32796) );
  NAND U33969 ( .A(n32741), .B(n32740), .Z(n32745) );
  NAND U33970 ( .A(n32743), .B(n32742), .Z(n32744) );
  NAND U33971 ( .A(n32745), .B(n32744), .Z(n32801) );
  NAND U33972 ( .A(n32747), .B(n32746), .Z(n32751) );
  NAND U33973 ( .A(n32749), .B(n32748), .Z(n32750) );
  NAND U33974 ( .A(n32751), .B(n32750), .Z(n32800) );
  XOR U33975 ( .A(n32801), .B(n32800), .Z(n32803) );
  NAND U33976 ( .A(n32753), .B(n32752), .Z(n32757) );
  NAND U33977 ( .A(n32755), .B(n32754), .Z(n32756) );
  AND U33978 ( .A(n32757), .B(n32756), .Z(n32833) );
  NAND U33979 ( .A(x[501]), .B(y[8008]), .Z(n33704) );
  NANDN U33980 ( .A(n33704), .B(n32758), .Z(n32762) );
  NAND U33981 ( .A(n32760), .B(n32759), .Z(n32761) );
  NAND U33982 ( .A(n32762), .B(n32761), .Z(n32907) );
  NAND U33983 ( .A(x[502]), .B(y[8003]), .Z(n32876) );
  NAND U33984 ( .A(x[485]), .B(y[8020]), .Z(n32875) );
  NAND U33985 ( .A(x[497]), .B(y[8008]), .Z(n32874) );
  XOR U33986 ( .A(n32875), .B(n32874), .Z(n32877) );
  XNOR U33987 ( .A(n32876), .B(n32877), .Z(n32906) );
  AND U33988 ( .A(y[8005]), .B(x[500]), .Z(n32764) );
  NAND U33989 ( .A(y[8004]), .B(x[501]), .Z(n32763) );
  XNOR U33990 ( .A(n32764), .B(n32763), .Z(n32889) );
  AND U33991 ( .A(x[499]), .B(y[8006]), .Z(n32888) );
  XOR U33992 ( .A(n32889), .B(n32888), .Z(n32905) );
  XNOR U33993 ( .A(n32906), .B(n32905), .Z(n32908) );
  XOR U33994 ( .A(n32907), .B(n32908), .Z(n32831) );
  NAND U33995 ( .A(n32887), .B(n33080), .Z(n32768) );
  NAND U33996 ( .A(n32766), .B(n32765), .Z(n32767) );
  NAND U33997 ( .A(n32768), .B(n32767), .Z(n32913) );
  NAND U33998 ( .A(x[495]), .B(y[8010]), .Z(n32895) );
  NAND U33999 ( .A(x[498]), .B(y[8007]), .Z(n32894) );
  NAND U34000 ( .A(x[486]), .B(y[8019]), .Z(n32893) );
  XOR U34001 ( .A(n32894), .B(n32893), .Z(n32896) );
  XNOR U34002 ( .A(n32895), .B(n32896), .Z(n32912) );
  NAND U34003 ( .A(x[503]), .B(y[8002]), .Z(n32870) );
  NAND U34004 ( .A(x[484]), .B(y[8021]), .Z(n32869) );
  NAND U34005 ( .A(x[496]), .B(y[8009]), .Z(n32868) );
  XOR U34006 ( .A(n32869), .B(n32868), .Z(n32871) );
  XNOR U34007 ( .A(n32870), .B(n32871), .Z(n32911) );
  XNOR U34008 ( .A(n32912), .B(n32911), .Z(n32914) );
  XOR U34009 ( .A(n32913), .B(n32914), .Z(n32830) );
  XOR U34010 ( .A(n32831), .B(n32830), .Z(n32832) );
  XNOR U34011 ( .A(n32833), .B(n32832), .Z(n32845) );
  NAND U34012 ( .A(n32770), .B(n32769), .Z(n32774) );
  NAND U34013 ( .A(n32772), .B(n32771), .Z(n32773) );
  NAND U34014 ( .A(n32774), .B(n32773), .Z(n32843) );
  NAND U34015 ( .A(n32776), .B(n32775), .Z(n32780) );
  NAND U34016 ( .A(n32778), .B(n32777), .Z(n32779) );
  NAND U34017 ( .A(n32780), .B(n32779), .Z(n32842) );
  XOR U34018 ( .A(n32843), .B(n32842), .Z(n32844) );
  XOR U34019 ( .A(n32845), .B(n32844), .Z(n32802) );
  XOR U34020 ( .A(n32803), .B(n32802), .Z(n32795) );
  NAND U34021 ( .A(n32782), .B(n32781), .Z(n32786) );
  NAND U34022 ( .A(n32784), .B(n32783), .Z(n32785) );
  NAND U34023 ( .A(n32786), .B(n32785), .Z(n32794) );
  XOR U34024 ( .A(n32796), .B(n32797), .Z(n32790) );
  XOR U34025 ( .A(n32791), .B(n32790), .Z(n32937) );
  XNOR U34026 ( .A(n32936), .B(n32937), .Z(n32939) );
  XNOR U34027 ( .A(n32931), .B(n32932), .Z(n32787) );
  XOR U34028 ( .A(n32929), .B(n32787), .Z(N698) );
  NANDN U34029 ( .A(n32789), .B(n32788), .Z(n32793) );
  NAND U34030 ( .A(n32791), .B(n32790), .Z(n32792) );
  AND U34031 ( .A(n32793), .B(n32792), .Z(n32943) );
  NANDN U34032 ( .A(n32795), .B(n32794), .Z(n32799) );
  NAND U34033 ( .A(n32797), .B(n32796), .Z(n32798) );
  NAND U34034 ( .A(n32799), .B(n32798), .Z(n32944) );
  NAND U34035 ( .A(n32801), .B(n32800), .Z(n32805) );
  NAND U34036 ( .A(n32803), .B(n32802), .Z(n32804) );
  NAND U34037 ( .A(n32805), .B(n32804), .Z(n33101) );
  AND U34038 ( .A(x[482]), .B(y[8024]), .Z(n32974) );
  XOR U34039 ( .A(n32975), .B(n32974), .Z(n32977) );
  AND U34040 ( .A(x[504]), .B(y[8002]), .Z(n32976) );
  XOR U34041 ( .A(n32977), .B(n32976), .Z(n33011) );
  NAND U34042 ( .A(n32807), .B(n32806), .Z(n32811) );
  NAND U34043 ( .A(n32809), .B(n32808), .Z(n32810) );
  AND U34044 ( .A(n32811), .B(n32810), .Z(n33010) );
  XOR U34045 ( .A(n33011), .B(n33010), .Z(n33013) );
  NANDN U34046 ( .A(n32813), .B(n32812), .Z(n32817) );
  NAND U34047 ( .A(n32815), .B(n32814), .Z(n32816) );
  AND U34048 ( .A(n32817), .B(n32816), .Z(n33012) );
  XNOR U34049 ( .A(n33013), .B(n33012), .Z(n33049) );
  NAND U34050 ( .A(n32819), .B(n32818), .Z(n32823) );
  NANDN U34051 ( .A(n32821), .B(n32820), .Z(n32822) );
  AND U34052 ( .A(n32823), .B(n32822), .Z(n33048) );
  XOR U34053 ( .A(n33049), .B(n33048), .Z(n33051) );
  NAND U34054 ( .A(n32825), .B(n32824), .Z(n32829) );
  NANDN U34055 ( .A(n32827), .B(n32826), .Z(n32828) );
  AND U34056 ( .A(n32829), .B(n32828), .Z(n33050) );
  XOR U34057 ( .A(n33051), .B(n33050), .Z(n33095) );
  NAND U34058 ( .A(n32831), .B(n32830), .Z(n32835) );
  NAND U34059 ( .A(n32833), .B(n32832), .Z(n32834) );
  NAND U34060 ( .A(n32835), .B(n32834), .Z(n33093) );
  NAND U34061 ( .A(n32837), .B(n32836), .Z(n32841) );
  NAND U34062 ( .A(n32839), .B(n32838), .Z(n32840) );
  AND U34063 ( .A(n32841), .B(n32840), .Z(n33092) );
  XOR U34064 ( .A(n33093), .B(n33092), .Z(n33094) );
  XNOR U34065 ( .A(n33095), .B(n33094), .Z(n33099) );
  NAND U34066 ( .A(n32843), .B(n32842), .Z(n32847) );
  NAND U34067 ( .A(n32845), .B(n32844), .Z(n32846) );
  NAND U34068 ( .A(n32847), .B(n32846), .Z(n33045) );
  AND U34069 ( .A(y[8020]), .B(x[486]), .Z(n32849) );
  NAND U34070 ( .A(y[8018]), .B(x[488]), .Z(n32848) );
  XNOR U34071 ( .A(n32849), .B(n32848), .Z(n33082) );
  AND U34072 ( .A(x[489]), .B(y[8017]), .Z(n33081) );
  XOR U34073 ( .A(n33082), .B(n33081), .Z(n33054) );
  AND U34074 ( .A(x[487]), .B(y[8019]), .Z(n33055) );
  XOR U34075 ( .A(n33054), .B(n33055), .Z(n33057) );
  AND U34076 ( .A(x[492]), .B(y[8014]), .Z(n33172) );
  AND U34077 ( .A(x[485]), .B(y[8021]), .Z(n33025) );
  XOR U34078 ( .A(n33172), .B(n33025), .Z(n33027) );
  AND U34079 ( .A(x[490]), .B(y[8016]), .Z(n33026) );
  XOR U34080 ( .A(n33027), .B(n33026), .Z(n33056) );
  XOR U34081 ( .A(n33057), .B(n33056), .Z(n33001) );
  NAND U34082 ( .A(n32851), .B(n32850), .Z(n32855) );
  NAND U34083 ( .A(n32853), .B(n32852), .Z(n32854) );
  NAND U34084 ( .A(n32855), .B(n32854), .Z(n32999) );
  NAND U34085 ( .A(n32857), .B(n32856), .Z(n32861) );
  NAND U34086 ( .A(n32859), .B(n32858), .Z(n32860) );
  NAND U34087 ( .A(n32861), .B(n32860), .Z(n32998) );
  XOR U34088 ( .A(n32999), .B(n32998), .Z(n33000) );
  XNOR U34089 ( .A(n33001), .B(n33000), .Z(n33037) );
  NANDN U34090 ( .A(n32863), .B(n32862), .Z(n32867) );
  NAND U34091 ( .A(n32865), .B(n32864), .Z(n32866) );
  AND U34092 ( .A(n32867), .B(n32866), .Z(n33036) );
  XOR U34093 ( .A(n33037), .B(n33036), .Z(n33039) );
  NAND U34094 ( .A(n32869), .B(n32868), .Z(n32873) );
  NAND U34095 ( .A(n32871), .B(n32870), .Z(n32872) );
  AND U34096 ( .A(n32873), .B(n32872), .Z(n32962) );
  NAND U34097 ( .A(n32875), .B(n32874), .Z(n32879) );
  NAND U34098 ( .A(n32877), .B(n32876), .Z(n32878) );
  AND U34099 ( .A(n32879), .B(n32878), .Z(n32963) );
  XOR U34100 ( .A(n32962), .B(n32963), .Z(n32965) );
  AND U34101 ( .A(n32880), .B(o[345]), .Z(n33074) );
  AND U34102 ( .A(x[494]), .B(y[8012]), .Z(n33075) );
  XOR U34103 ( .A(n33074), .B(n33075), .Z(n33076) );
  AND U34104 ( .A(x[481]), .B(y[8025]), .Z(n33077) );
  XOR U34105 ( .A(n33076), .B(n33077), .Z(n33017) );
  AND U34106 ( .A(x[505]), .B(y[8001]), .Z(n33085) );
  XOR U34107 ( .A(o[346]), .B(n33085), .Z(n33031) );
  AND U34108 ( .A(x[506]), .B(y[8000]), .Z(n33030) );
  XOR U34109 ( .A(n33031), .B(n33030), .Z(n33033) );
  AND U34110 ( .A(x[480]), .B(y[8026]), .Z(n33032) );
  XOR U34111 ( .A(n33033), .B(n33032), .Z(n33016) );
  XOR U34112 ( .A(n33017), .B(n33016), .Z(n33019) );
  NAND U34113 ( .A(n32882), .B(n32881), .Z(n32886) );
  NAND U34114 ( .A(n32884), .B(n32883), .Z(n32885) );
  AND U34115 ( .A(n32886), .B(n32885), .Z(n33018) );
  XOR U34116 ( .A(n33019), .B(n33018), .Z(n32964) );
  XNOR U34117 ( .A(n32965), .B(n32964), .Z(n33007) );
  AND U34118 ( .A(x[501]), .B(y[8005]), .Z(n32892) );
  IV U34119 ( .A(n32892), .Z(n33068) );
  NANDN U34120 ( .A(n33068), .B(n32887), .Z(n32891) );
  NAND U34121 ( .A(n32889), .B(n32888), .Z(n32890) );
  NAND U34122 ( .A(n32891), .B(n32890), .Z(n32995) );
  XOR U34123 ( .A(n33069), .B(n32892), .Z(n33070) );
  AND U34124 ( .A(x[500]), .B(y[8006]), .Z(n33071) );
  XOR U34125 ( .A(n33070), .B(n33071), .Z(n32993) );
  AND U34126 ( .A(x[503]), .B(y[8003]), .Z(n32981) );
  XOR U34127 ( .A(n32980), .B(n32981), .Z(n32982) );
  AND U34128 ( .A(x[502]), .B(y[8004]), .Z(n32983) );
  XOR U34129 ( .A(n32982), .B(n32983), .Z(n32992) );
  XOR U34130 ( .A(n32993), .B(n32992), .Z(n32994) );
  XNOR U34131 ( .A(n32995), .B(n32994), .Z(n33005) );
  AND U34132 ( .A(x[484]), .B(y[8022]), .Z(n32986) );
  XOR U34133 ( .A(n32987), .B(n32986), .Z(n32988) );
  XNOR U34134 ( .A(n32988), .B(n32989), .Z(n32969) );
  AND U34135 ( .A(x[483]), .B(y[8023]), .Z(n33060) );
  AND U34136 ( .A(x[491]), .B(y[8015]), .Z(n33061) );
  XOR U34137 ( .A(n33060), .B(n33061), .Z(n33062) );
  AND U34138 ( .A(x[499]), .B(y[8007]), .Z(n33063) );
  XOR U34139 ( .A(n33062), .B(n33063), .Z(n32968) );
  XOR U34140 ( .A(n32969), .B(n32968), .Z(n32971) );
  NAND U34141 ( .A(n32894), .B(n32893), .Z(n32898) );
  NAND U34142 ( .A(n32896), .B(n32895), .Z(n32897) );
  AND U34143 ( .A(n32898), .B(n32897), .Z(n32970) );
  XNOR U34144 ( .A(n32971), .B(n32970), .Z(n33004) );
  XOR U34145 ( .A(n33005), .B(n33004), .Z(n33006) );
  XOR U34146 ( .A(n33007), .B(n33006), .Z(n33038) );
  XNOR U34147 ( .A(n33039), .B(n33038), .Z(n33043) );
  NAND U34148 ( .A(n32900), .B(n32899), .Z(n32904) );
  NAND U34149 ( .A(n32902), .B(n32901), .Z(n32903) );
  NAND U34150 ( .A(n32904), .B(n32903), .Z(n33089) );
  NAND U34151 ( .A(n32906), .B(n32905), .Z(n32910) );
  NANDN U34152 ( .A(n32908), .B(n32907), .Z(n32909) );
  NAND U34153 ( .A(n32910), .B(n32909), .Z(n33087) );
  NAND U34154 ( .A(n32912), .B(n32911), .Z(n32916) );
  NANDN U34155 ( .A(n32914), .B(n32913), .Z(n32915) );
  NAND U34156 ( .A(n32916), .B(n32915), .Z(n33086) );
  XOR U34157 ( .A(n33087), .B(n33086), .Z(n33088) );
  XOR U34158 ( .A(n33089), .B(n33088), .Z(n33042) );
  XOR U34159 ( .A(n33043), .B(n33042), .Z(n33044) );
  XOR U34160 ( .A(n33045), .B(n33044), .Z(n33098) );
  XOR U34161 ( .A(n33099), .B(n33098), .Z(n33100) );
  XOR U34162 ( .A(n33101), .B(n33100), .Z(n32959) );
  NAND U34163 ( .A(n32918), .B(n32917), .Z(n32922) );
  NAND U34164 ( .A(n32920), .B(n32919), .Z(n32921) );
  AND U34165 ( .A(n32922), .B(n32921), .Z(n32956) );
  NAND U34166 ( .A(n32924), .B(n32923), .Z(n32928) );
  NAND U34167 ( .A(n32926), .B(n32925), .Z(n32927) );
  AND U34168 ( .A(n32928), .B(n32927), .Z(n32957) );
  XOR U34169 ( .A(n32956), .B(n32957), .Z(n32958) );
  XOR U34170 ( .A(n32959), .B(n32958), .Z(n32945) );
  XNOR U34171 ( .A(n32946), .B(n32945), .Z(n32952) );
  OR U34172 ( .A(n32931), .B(n32929), .Z(n32935) );
  ANDN U34173 ( .B(n32931), .A(n32930), .Z(n32933) );
  OR U34174 ( .A(n32933), .B(n32932), .Z(n32934) );
  AND U34175 ( .A(n32935), .B(n32934), .Z(n32951) );
  NAND U34176 ( .A(n32937), .B(n32936), .Z(n32941) );
  NANDN U34177 ( .A(n32939), .B(n32938), .Z(n32940) );
  AND U34178 ( .A(n32941), .B(n32940), .Z(n32950) );
  IV U34179 ( .A(n32950), .Z(n32949) );
  XOR U34180 ( .A(n32951), .B(n32949), .Z(n32942) );
  XNOR U34181 ( .A(n32952), .B(n32942), .Z(N699) );
  NANDN U34182 ( .A(n32944), .B(n32943), .Z(n32948) );
  NAND U34183 ( .A(n32946), .B(n32945), .Z(n32947) );
  NAND U34184 ( .A(n32948), .B(n32947), .Z(n33112) );
  IV U34185 ( .A(n33112), .Z(n33111) );
  OR U34186 ( .A(n32951), .B(n32949), .Z(n32955) );
  ANDN U34187 ( .B(n32951), .A(n32950), .Z(n32953) );
  OR U34188 ( .A(n32953), .B(n32952), .Z(n32954) );
  AND U34189 ( .A(n32955), .B(n32954), .Z(n33113) );
  NAND U34190 ( .A(n32957), .B(n32956), .Z(n32961) );
  NAND U34191 ( .A(n32959), .B(n32958), .Z(n32960) );
  AND U34192 ( .A(n32961), .B(n32960), .Z(n33108) );
  NAND U34193 ( .A(n32963), .B(n32962), .Z(n32967) );
  NAND U34194 ( .A(n32965), .B(n32964), .Z(n32966) );
  NAND U34195 ( .A(n32967), .B(n32966), .Z(n33247) );
  NAND U34196 ( .A(n32969), .B(n32968), .Z(n32973) );
  NAND U34197 ( .A(n32971), .B(n32970), .Z(n32972) );
  NAND U34198 ( .A(n32973), .B(n32972), .Z(n33245) );
  AND U34199 ( .A(n32975), .B(n32974), .Z(n32979) );
  NAND U34200 ( .A(n32977), .B(n32976), .Z(n32978) );
  NANDN U34201 ( .A(n32979), .B(n32978), .Z(n33143) );
  NAND U34202 ( .A(n32981), .B(n32980), .Z(n32985) );
  NAND U34203 ( .A(n32983), .B(n32982), .Z(n32984) );
  NAND U34204 ( .A(n32985), .B(n32984), .Z(n33142) );
  XOR U34205 ( .A(n33143), .B(n33142), .Z(n33144) );
  AND U34206 ( .A(n32987), .B(n32986), .Z(n32991) );
  NANDN U34207 ( .A(n32989), .B(n32988), .Z(n32990) );
  NANDN U34208 ( .A(n32991), .B(n32990), .Z(n33156) );
  AND U34209 ( .A(x[480]), .B(y[8027]), .Z(n33234) );
  AND U34210 ( .A(x[507]), .B(y[8000]), .Z(n33233) );
  XOR U34211 ( .A(n33234), .B(n33233), .Z(n33236) );
  AND U34212 ( .A(x[506]), .B(y[8001]), .Z(n33224) );
  XOR U34213 ( .A(n33224), .B(o[347]), .Z(n33235) );
  XOR U34214 ( .A(n33236), .B(n33235), .Z(n33155) );
  AND U34215 ( .A(x[489]), .B(y[8018]), .Z(n33219) );
  AND U34216 ( .A(x[501]), .B(y[8006]), .Z(n33218) );
  XOR U34217 ( .A(n33219), .B(n33218), .Z(n33221) );
  AND U34218 ( .A(x[498]), .B(y[8009]), .Z(n33220) );
  XOR U34219 ( .A(n33221), .B(n33220), .Z(n33154) );
  XOR U34220 ( .A(n33155), .B(n33154), .Z(n33157) );
  XNOR U34221 ( .A(n33156), .B(n33157), .Z(n33145) );
  XOR U34222 ( .A(n33245), .B(n33246), .Z(n33248) );
  XOR U34223 ( .A(n33247), .B(n33248), .Z(n33266) );
  NAND U34224 ( .A(n32993), .B(n32992), .Z(n32997) );
  NAND U34225 ( .A(n32995), .B(n32994), .Z(n32996) );
  AND U34226 ( .A(n32997), .B(n32996), .Z(n33264) );
  NAND U34227 ( .A(n32999), .B(n32998), .Z(n33003) );
  NAND U34228 ( .A(n33001), .B(n33000), .Z(n33002) );
  AND U34229 ( .A(n33003), .B(n33002), .Z(n33263) );
  XOR U34230 ( .A(n33264), .B(n33263), .Z(n33265) );
  NAND U34231 ( .A(n33005), .B(n33004), .Z(n33009) );
  NAND U34232 ( .A(n33007), .B(n33006), .Z(n33008) );
  AND U34233 ( .A(n33009), .B(n33008), .Z(n33251) );
  NAND U34234 ( .A(n33011), .B(n33010), .Z(n33015) );
  NAND U34235 ( .A(n33013), .B(n33012), .Z(n33014) );
  NAND U34236 ( .A(n33015), .B(n33014), .Z(n33241) );
  NAND U34237 ( .A(n33017), .B(n33016), .Z(n33021) );
  NAND U34238 ( .A(n33019), .B(n33018), .Z(n33020) );
  NAND U34239 ( .A(n33021), .B(n33020), .Z(n33239) );
  AND U34240 ( .A(x[499]), .B(y[8008]), .Z(n33213) );
  AND U34241 ( .A(x[505]), .B(y[8002]), .Z(n33212) );
  XOR U34242 ( .A(n33213), .B(n33212), .Z(n33215) );
  AND U34243 ( .A(x[486]), .B(y[8021]), .Z(n33214) );
  XOR U34244 ( .A(n33215), .B(n33214), .Z(n33202) );
  AND U34245 ( .A(x[495]), .B(y[8012]), .Z(n33178) );
  AND U34246 ( .A(x[482]), .B(y[8025]), .Z(n33177) );
  XOR U34247 ( .A(n33178), .B(n33177), .Z(n33180) );
  AND U34248 ( .A(x[483]), .B(y[8024]), .Z(n33179) );
  XOR U34249 ( .A(n33180), .B(n33179), .Z(n33201) );
  XOR U34250 ( .A(n33202), .B(n33201), .Z(n33203) );
  NAND U34251 ( .A(x[496]), .B(y[8011]), .Z(n33160) );
  XOR U34252 ( .A(n33160), .B(n33022), .Z(n33163) );
  XOR U34253 ( .A(n33162), .B(n33163), .Z(n33174) );
  AND U34254 ( .A(y[8014]), .B(x[493]), .Z(n33024) );
  AND U34255 ( .A(y[8015]), .B(x[492]), .Z(n33023) );
  XOR U34256 ( .A(n33024), .B(n33023), .Z(n33173) );
  XNOR U34257 ( .A(n33203), .B(n33204), .Z(n33139) );
  AND U34258 ( .A(n33172), .B(n33025), .Z(n33029) );
  NAND U34259 ( .A(n33027), .B(n33026), .Z(n33028) );
  NANDN U34260 ( .A(n33029), .B(n33028), .Z(n33137) );
  NAND U34261 ( .A(n33031), .B(n33030), .Z(n33035) );
  NAND U34262 ( .A(n33033), .B(n33032), .Z(n33034) );
  NAND U34263 ( .A(n33035), .B(n33034), .Z(n33136) );
  XOR U34264 ( .A(n33137), .B(n33136), .Z(n33138) );
  XOR U34265 ( .A(n33139), .B(n33138), .Z(n33240) );
  XNOR U34266 ( .A(n33239), .B(n33240), .Z(n33242) );
  XNOR U34267 ( .A(n33251), .B(n33252), .Z(n33254) );
  NAND U34268 ( .A(n33037), .B(n33036), .Z(n33041) );
  NAND U34269 ( .A(n33039), .B(n33038), .Z(n33040) );
  AND U34270 ( .A(n33041), .B(n33040), .Z(n33253) );
  XOR U34271 ( .A(n33254), .B(n33253), .Z(n33124) );
  NAND U34272 ( .A(n33043), .B(n33042), .Z(n33047) );
  NAND U34273 ( .A(n33045), .B(n33044), .Z(n33046) );
  NAND U34274 ( .A(n33047), .B(n33046), .Z(n33126) );
  XOR U34275 ( .A(n33127), .B(n33126), .Z(n33121) );
  NAND U34276 ( .A(n33049), .B(n33048), .Z(n33053) );
  NAND U34277 ( .A(n33051), .B(n33050), .Z(n33052) );
  NAND U34278 ( .A(n33053), .B(n33052), .Z(n33130) );
  NAND U34279 ( .A(n33055), .B(n33054), .Z(n33059) );
  NAND U34280 ( .A(n33057), .B(n33056), .Z(n33058) );
  AND U34281 ( .A(n33059), .B(n33058), .Z(n33259) );
  NAND U34282 ( .A(n33061), .B(n33060), .Z(n33065) );
  NAND U34283 ( .A(n33063), .B(n33062), .Z(n33064) );
  NAND U34284 ( .A(n33065), .B(n33064), .Z(n33197) );
  AND U34285 ( .A(y[8003]), .B(x[504]), .Z(n33067) );
  NAND U34286 ( .A(y[8007]), .B(x[500]), .Z(n33066) );
  XNOR U34287 ( .A(n33067), .B(n33066), .Z(n33209) );
  AND U34288 ( .A(x[487]), .B(y[8020]), .Z(n33208) );
  XOR U34289 ( .A(n33209), .B(n33208), .Z(n33196) );
  AND U34290 ( .A(x[488]), .B(y[8019]), .Z(n33167) );
  AND U34291 ( .A(x[503]), .B(y[8004]), .Z(n33166) );
  XOR U34292 ( .A(n33167), .B(n33166), .Z(n33169) );
  AND U34293 ( .A(x[502]), .B(y[8005]), .Z(n33168) );
  XOR U34294 ( .A(n33169), .B(n33168), .Z(n33195) );
  XOR U34295 ( .A(n33196), .B(n33195), .Z(n33198) );
  XOR U34296 ( .A(n33197), .B(n33198), .Z(n33258) );
  ANDN U34297 ( .B(n33069), .A(n33068), .Z(n33073) );
  NAND U34298 ( .A(n33071), .B(n33070), .Z(n33072) );
  NANDN U34299 ( .A(n33073), .B(n33072), .Z(n33190) );
  NAND U34300 ( .A(n33075), .B(n33074), .Z(n33079) );
  NAND U34301 ( .A(n33077), .B(n33076), .Z(n33078) );
  NAND U34302 ( .A(n33079), .B(n33078), .Z(n33189) );
  XOR U34303 ( .A(n33190), .B(n33189), .Z(n33191) );
  AND U34304 ( .A(y[8020]), .B(x[488]), .Z(n33226) );
  NAND U34305 ( .A(n33080), .B(n33226), .Z(n33084) );
  NAND U34306 ( .A(n33082), .B(n33081), .Z(n33083) );
  NAND U34307 ( .A(n33084), .B(n33083), .Z(n33150) );
  AND U34308 ( .A(x[494]), .B(y[8013]), .Z(n33184) );
  AND U34309 ( .A(x[481]), .B(y[8026]), .Z(n33183) );
  XOR U34310 ( .A(n33184), .B(n33183), .Z(n33186) );
  AND U34311 ( .A(o[346]), .B(n33085), .Z(n33185) );
  XOR U34312 ( .A(n33186), .B(n33185), .Z(n33149) );
  AND U34313 ( .A(x[497]), .B(y[8010]), .Z(n33228) );
  AND U34314 ( .A(x[484]), .B(y[8023]), .Z(n33227) );
  XOR U34315 ( .A(n33228), .B(n33227), .Z(n33230) );
  AND U34316 ( .A(x[485]), .B(y[8022]), .Z(n33229) );
  XOR U34317 ( .A(n33230), .B(n33229), .Z(n33148) );
  XOR U34318 ( .A(n33149), .B(n33148), .Z(n33151) );
  XOR U34319 ( .A(n33150), .B(n33151), .Z(n33192) );
  XNOR U34320 ( .A(n33191), .B(n33192), .Z(n33257) );
  XNOR U34321 ( .A(n33259), .B(n33260), .Z(n33131) );
  XOR U34322 ( .A(n33130), .B(n33131), .Z(n33133) );
  NAND U34323 ( .A(n33087), .B(n33086), .Z(n33091) );
  NAND U34324 ( .A(n33089), .B(n33088), .Z(n33090) );
  AND U34325 ( .A(n33091), .B(n33090), .Z(n33132) );
  XNOR U34326 ( .A(n33133), .B(n33132), .Z(n33119) );
  NAND U34327 ( .A(n33093), .B(n33092), .Z(n33097) );
  NAND U34328 ( .A(n33095), .B(n33094), .Z(n33096) );
  AND U34329 ( .A(n33097), .B(n33096), .Z(n33118) );
  XOR U34330 ( .A(n33119), .B(n33118), .Z(n33120) );
  XNOR U34331 ( .A(n33121), .B(n33120), .Z(n33106) );
  NAND U34332 ( .A(n33099), .B(n33098), .Z(n33103) );
  NAND U34333 ( .A(n33101), .B(n33100), .Z(n33102) );
  AND U34334 ( .A(n33103), .B(n33102), .Z(n33105) );
  XOR U34335 ( .A(n33106), .B(n33105), .Z(n33107) );
  XOR U34336 ( .A(n33108), .B(n33107), .Z(n33114) );
  XNOR U34337 ( .A(n33113), .B(n33114), .Z(n33104) );
  XOR U34338 ( .A(n33111), .B(n33104), .Z(N700) );
  NAND U34339 ( .A(n33106), .B(n33105), .Z(n33110) );
  NAND U34340 ( .A(n33108), .B(n33107), .Z(n33109) );
  NAND U34341 ( .A(n33110), .B(n33109), .Z(n33435) );
  IV U34342 ( .A(n33435), .Z(n33433) );
  OR U34343 ( .A(n33113), .B(n33111), .Z(n33117) );
  ANDN U34344 ( .B(n33113), .A(n33112), .Z(n33115) );
  OR U34345 ( .A(n33115), .B(n33114), .Z(n33116) );
  AND U34346 ( .A(n33117), .B(n33116), .Z(n33434) );
  NAND U34347 ( .A(n33119), .B(n33118), .Z(n33123) );
  NAND U34348 ( .A(n33121), .B(n33120), .Z(n33122) );
  NAND U34349 ( .A(n33123), .B(n33122), .Z(n33428) );
  NANDN U34350 ( .A(n33125), .B(n33124), .Z(n33129) );
  NAND U34351 ( .A(n33127), .B(n33126), .Z(n33128) );
  NAND U34352 ( .A(n33129), .B(n33128), .Z(n33427) );
  XOR U34353 ( .A(n33428), .B(n33427), .Z(n33430) );
  NAND U34354 ( .A(n33131), .B(n33130), .Z(n33135) );
  NAND U34355 ( .A(n33133), .B(n33132), .Z(n33134) );
  AND U34356 ( .A(n33135), .B(n33134), .Z(n33270) );
  NAND U34357 ( .A(n33137), .B(n33136), .Z(n33141) );
  NAND U34358 ( .A(n33139), .B(n33138), .Z(n33140) );
  NAND U34359 ( .A(n33141), .B(n33140), .Z(n33294) );
  NAND U34360 ( .A(n33143), .B(n33142), .Z(n33147) );
  NANDN U34361 ( .A(n33145), .B(n33144), .Z(n33146) );
  NAND U34362 ( .A(n33147), .B(n33146), .Z(n33399) );
  NAND U34363 ( .A(n33149), .B(n33148), .Z(n33153) );
  NAND U34364 ( .A(n33151), .B(n33150), .Z(n33152) );
  NAND U34365 ( .A(n33153), .B(n33152), .Z(n33398) );
  NAND U34366 ( .A(n33155), .B(n33154), .Z(n33159) );
  NAND U34367 ( .A(n33157), .B(n33156), .Z(n33158) );
  NAND U34368 ( .A(n33159), .B(n33158), .Z(n33397) );
  XOR U34369 ( .A(n33398), .B(n33397), .Z(n33400) );
  XOR U34370 ( .A(n33399), .B(n33400), .Z(n33295) );
  XOR U34371 ( .A(n33294), .B(n33295), .Z(n33297) );
  AND U34372 ( .A(x[495]), .B(y[8013]), .Z(n33374) );
  AND U34373 ( .A(x[507]), .B(y[8001]), .Z(n33358) );
  XOR U34374 ( .A(o[348]), .B(n33358), .Z(n33372) );
  AND U34375 ( .A(x[506]), .B(y[8002]), .Z(n33371) );
  XOR U34376 ( .A(n33372), .B(n33371), .Z(n33373) );
  XOR U34377 ( .A(n33374), .B(n33373), .Z(n33360) );
  AND U34378 ( .A(x[487]), .B(y[8021]), .Z(n33342) );
  AND U34379 ( .A(x[492]), .B(y[8016]), .Z(n33341) );
  XOR U34380 ( .A(n33342), .B(n33341), .Z(n33344) );
  AND U34381 ( .A(x[491]), .B(y[8017]), .Z(n33343) );
  XNOR U34382 ( .A(n33344), .B(n33343), .Z(n33359) );
  NANDN U34383 ( .A(n33161), .B(n33160), .Z(n33165) );
  NAND U34384 ( .A(n33163), .B(n33162), .Z(n33164) );
  NAND U34385 ( .A(n33165), .B(n33164), .Z(n33361) );
  XOR U34386 ( .A(n33362), .B(n33361), .Z(n33404) );
  AND U34387 ( .A(x[497]), .B(y[8011]), .Z(n33307) );
  AND U34388 ( .A(x[502]), .B(y[8006]), .Z(n33306) );
  XOR U34389 ( .A(n33307), .B(n33306), .Z(n33309) );
  AND U34390 ( .A(x[484]), .B(y[8024]), .Z(n33308) );
  XOR U34391 ( .A(n33309), .B(n33308), .Z(n33380) );
  AND U34392 ( .A(x[486]), .B(y[8022]), .Z(n33521) );
  AND U34393 ( .A(x[499]), .B(y[8009]), .Z(n33347) );
  XOR U34394 ( .A(n33521), .B(n33347), .Z(n33349) );
  XOR U34395 ( .A(n33349), .B(n33348), .Z(n33379) );
  XOR U34396 ( .A(n33380), .B(n33379), .Z(n33382) );
  NAND U34397 ( .A(n33167), .B(n33166), .Z(n33171) );
  NAND U34398 ( .A(n33169), .B(n33168), .Z(n33170) );
  NAND U34399 ( .A(n33171), .B(n33170), .Z(n33381) );
  XOR U34400 ( .A(n33382), .B(n33381), .Z(n33403) );
  NAND U34401 ( .A(n33366), .B(n33172), .Z(n33176) );
  NANDN U34402 ( .A(n33174), .B(n33173), .Z(n33175) );
  NAND U34403 ( .A(n33176), .B(n33175), .Z(n33325) );
  NAND U34404 ( .A(n33178), .B(n33177), .Z(n33182) );
  NAND U34405 ( .A(n33180), .B(n33179), .Z(n33181) );
  NAND U34406 ( .A(n33182), .B(n33181), .Z(n33324) );
  NAND U34407 ( .A(n33184), .B(n33183), .Z(n33188) );
  NAND U34408 ( .A(n33186), .B(n33185), .Z(n33187) );
  NAND U34409 ( .A(n33188), .B(n33187), .Z(n33323) );
  XOR U34410 ( .A(n33324), .B(n33323), .Z(n33326) );
  XOR U34411 ( .A(n33325), .B(n33326), .Z(n33405) );
  XOR U34412 ( .A(n33406), .B(n33405), .Z(n33296) );
  XNOR U34413 ( .A(n33297), .B(n33296), .Z(n33291) );
  NAND U34414 ( .A(n33190), .B(n33189), .Z(n33194) );
  NAND U34415 ( .A(n33192), .B(n33191), .Z(n33193) );
  NAND U34416 ( .A(n33194), .B(n33193), .Z(n33387) );
  NAND U34417 ( .A(n33196), .B(n33195), .Z(n33200) );
  NAND U34418 ( .A(n33198), .B(n33197), .Z(n33199) );
  NAND U34419 ( .A(n33200), .B(n33199), .Z(n33386) );
  NAND U34420 ( .A(n33202), .B(n33201), .Z(n33206) );
  NANDN U34421 ( .A(n33204), .B(n33203), .Z(n33205) );
  NAND U34422 ( .A(n33206), .B(n33205), .Z(n33385) );
  XOR U34423 ( .A(n33386), .B(n33385), .Z(n33388) );
  XOR U34424 ( .A(n33387), .B(n33388), .Z(n33289) );
  AND U34425 ( .A(x[504]), .B(y[8007]), .Z(n33764) );
  AND U34426 ( .A(x[500]), .B(y[8003]), .Z(n33207) );
  NAND U34427 ( .A(n33764), .B(n33207), .Z(n33211) );
  NAND U34428 ( .A(n33209), .B(n33208), .Z(n33210) );
  NAND U34429 ( .A(n33211), .B(n33210), .Z(n33423) );
  AND U34430 ( .A(x[505]), .B(y[8003]), .Z(n33337) );
  XOR U34431 ( .A(n33338), .B(n33337), .Z(n33336) );
  AND U34432 ( .A(x[481]), .B(y[8027]), .Z(n33335) );
  XOR U34433 ( .A(n33336), .B(n33335), .Z(n33422) );
  AND U34434 ( .A(x[496]), .B(y[8012]), .Z(n33330) );
  AND U34435 ( .A(x[504]), .B(y[8004]), .Z(n33329) );
  XOR U34436 ( .A(n33330), .B(n33329), .Z(n33332) );
  AND U34437 ( .A(x[482]), .B(y[8026]), .Z(n33331) );
  XOR U34438 ( .A(n33332), .B(n33331), .Z(n33421) );
  XOR U34439 ( .A(n33422), .B(n33421), .Z(n33424) );
  XOR U34440 ( .A(n33423), .B(n33424), .Z(n33394) );
  NAND U34441 ( .A(n33213), .B(n33212), .Z(n33217) );
  NAND U34442 ( .A(n33215), .B(n33214), .Z(n33216) );
  NAND U34443 ( .A(n33217), .B(n33216), .Z(n33417) );
  AND U34444 ( .A(x[483]), .B(y[8025]), .Z(n33365) );
  XOR U34445 ( .A(n33366), .B(n33365), .Z(n33368) );
  AND U34446 ( .A(x[503]), .B(y[8005]), .Z(n33367) );
  XOR U34447 ( .A(n33368), .B(n33367), .Z(n33416) );
  AND U34448 ( .A(x[485]), .B(y[8023]), .Z(n33353) );
  AND U34449 ( .A(x[501]), .B(y[8007]), .Z(n33352) );
  XOR U34450 ( .A(n33353), .B(n33352), .Z(n33355) );
  AND U34451 ( .A(x[500]), .B(y[8008]), .Z(n33354) );
  XOR U34452 ( .A(n33355), .B(n33354), .Z(n33415) );
  XOR U34453 ( .A(n33416), .B(n33415), .Z(n33418) );
  XOR U34454 ( .A(n33417), .B(n33418), .Z(n33392) );
  NAND U34455 ( .A(n33219), .B(n33218), .Z(n33223) );
  NAND U34456 ( .A(n33221), .B(n33220), .Z(n33222) );
  NAND U34457 ( .A(n33223), .B(n33222), .Z(n33302) );
  AND U34458 ( .A(x[480]), .B(y[8028]), .Z(n33313) );
  AND U34459 ( .A(x[508]), .B(y[8000]), .Z(n33312) );
  XOR U34460 ( .A(n33313), .B(n33312), .Z(n33315) );
  AND U34461 ( .A(n33224), .B(o[347]), .Z(n33314) );
  XOR U34462 ( .A(n33315), .B(n33314), .Z(n33301) );
  NAND U34463 ( .A(y[8018]), .B(x[490]), .Z(n33225) );
  XNOR U34464 ( .A(n33226), .B(n33225), .Z(n33320) );
  AND U34465 ( .A(x[489]), .B(y[8019]), .Z(n33319) );
  XOR U34466 ( .A(n33320), .B(n33319), .Z(n33300) );
  XOR U34467 ( .A(n33301), .B(n33300), .Z(n33303) );
  XOR U34468 ( .A(n33302), .B(n33303), .Z(n33412) );
  NAND U34469 ( .A(n33228), .B(n33227), .Z(n33232) );
  NAND U34470 ( .A(n33230), .B(n33229), .Z(n33231) );
  NAND U34471 ( .A(n33232), .B(n33231), .Z(n33410) );
  NAND U34472 ( .A(n33234), .B(n33233), .Z(n33238) );
  NAND U34473 ( .A(n33236), .B(n33235), .Z(n33237) );
  NAND U34474 ( .A(n33238), .B(n33237), .Z(n33409) );
  XOR U34475 ( .A(n33410), .B(n33409), .Z(n33411) );
  XNOR U34476 ( .A(n33412), .B(n33411), .Z(n33391) );
  XNOR U34477 ( .A(n33291), .B(n33290), .Z(n33284) );
  NAND U34478 ( .A(n33240), .B(n33239), .Z(n33244) );
  NANDN U34479 ( .A(n33242), .B(n33241), .Z(n33243) );
  NAND U34480 ( .A(n33244), .B(n33243), .Z(n33283) );
  NAND U34481 ( .A(n33246), .B(n33245), .Z(n33250) );
  NAND U34482 ( .A(n33248), .B(n33247), .Z(n33249) );
  NAND U34483 ( .A(n33250), .B(n33249), .Z(n33282) );
  XNOR U34484 ( .A(n33283), .B(n33282), .Z(n33285) );
  XNOR U34485 ( .A(n33270), .B(n33271), .Z(n33272) );
  NANDN U34486 ( .A(n33252), .B(n33251), .Z(n33256) );
  NAND U34487 ( .A(n33254), .B(n33253), .Z(n33255) );
  NAND U34488 ( .A(n33256), .B(n33255), .Z(n33278) );
  NANDN U34489 ( .A(n33258), .B(n33257), .Z(n33262) );
  NANDN U34490 ( .A(n33260), .B(n33259), .Z(n33261) );
  AND U34491 ( .A(n33262), .B(n33261), .Z(n33277) );
  NAND U34492 ( .A(n33264), .B(n33263), .Z(n33268) );
  NANDN U34493 ( .A(n33266), .B(n33265), .Z(n33267) );
  AND U34494 ( .A(n33268), .B(n33267), .Z(n33276) );
  XOR U34495 ( .A(n33277), .B(n33276), .Z(n33279) );
  XNOR U34496 ( .A(n33278), .B(n33279), .Z(n33273) );
  XOR U34497 ( .A(n33430), .B(n33429), .Z(n33436) );
  XNOR U34498 ( .A(n33434), .B(n33436), .Z(n33269) );
  XOR U34499 ( .A(n33433), .B(n33269), .Z(N701) );
  NANDN U34500 ( .A(n33271), .B(n33270), .Z(n33275) );
  NANDN U34501 ( .A(n33273), .B(n33272), .Z(n33274) );
  NAND U34502 ( .A(n33275), .B(n33274), .Z(n33446) );
  NAND U34503 ( .A(n33277), .B(n33276), .Z(n33281) );
  NAND U34504 ( .A(n33279), .B(n33278), .Z(n33280) );
  NAND U34505 ( .A(n33281), .B(n33280), .Z(n33444) );
  NAND U34506 ( .A(n33283), .B(n33282), .Z(n33287) );
  NANDN U34507 ( .A(n33285), .B(n33284), .Z(n33286) );
  NAND U34508 ( .A(n33287), .B(n33286), .Z(n33450) );
  NANDN U34509 ( .A(n33289), .B(n33288), .Z(n33293) );
  NAND U34510 ( .A(n33291), .B(n33290), .Z(n33292) );
  AND U34511 ( .A(n33293), .B(n33292), .Z(n33451) );
  XOR U34512 ( .A(n33450), .B(n33451), .Z(n33453) );
  NAND U34513 ( .A(n33295), .B(n33294), .Z(n33299) );
  NAND U34514 ( .A(n33297), .B(n33296), .Z(n33298) );
  NAND U34515 ( .A(n33299), .B(n33298), .Z(n33462) );
  NAND U34516 ( .A(n33301), .B(n33300), .Z(n33305) );
  NAND U34517 ( .A(n33303), .B(n33302), .Z(n33304) );
  AND U34518 ( .A(n33305), .B(n33304), .Z(n33571) );
  NAND U34519 ( .A(n33307), .B(n33306), .Z(n33311) );
  NAND U34520 ( .A(n33309), .B(n33308), .Z(n33310) );
  NAND U34521 ( .A(n33311), .B(n33310), .Z(n33608) );
  NAND U34522 ( .A(n33313), .B(n33312), .Z(n33317) );
  NAND U34523 ( .A(n33315), .B(n33314), .Z(n33316) );
  NAND U34524 ( .A(n33317), .B(n33316), .Z(n33607) );
  XOR U34525 ( .A(n33608), .B(n33607), .Z(n33609) );
  AND U34526 ( .A(y[8020]), .B(x[490]), .Z(n33605) );
  NAND U34527 ( .A(n33318), .B(n33605), .Z(n33322) );
  NAND U34528 ( .A(n33320), .B(n33319), .Z(n33321) );
  NAND U34529 ( .A(n33322), .B(n33321), .Z(n33579) );
  AND U34530 ( .A(x[502]), .B(y[8007]), .Z(n33542) );
  AND U34531 ( .A(x[492]), .B(y[8017]), .Z(n33675) );
  AND U34532 ( .A(x[481]), .B(y[8028]), .Z(n33540) );
  XOR U34533 ( .A(n33675), .B(n33540), .Z(n33541) );
  XOR U34534 ( .A(n33542), .B(n33541), .Z(n33578) );
  AND U34535 ( .A(x[495]), .B(y[8014]), .Z(n33545) );
  XOR U34536 ( .A(n33578), .B(n33577), .Z(n33580) );
  XNOR U34537 ( .A(n33579), .B(n33580), .Z(n33610) );
  NAND U34538 ( .A(n33324), .B(n33323), .Z(n33328) );
  NAND U34539 ( .A(n33326), .B(n33325), .Z(n33327) );
  AND U34540 ( .A(n33328), .B(n33327), .Z(n33573) );
  XOR U34541 ( .A(n33574), .B(n33573), .Z(n33568) );
  NAND U34542 ( .A(n33330), .B(n33329), .Z(n33334) );
  NAND U34543 ( .A(n33332), .B(n33331), .Z(n33333) );
  NAND U34544 ( .A(n33334), .B(n33333), .Z(n33584) );
  AND U34545 ( .A(n33336), .B(n33335), .Z(n33340) );
  NAND U34546 ( .A(n33338), .B(n33337), .Z(n33339) );
  NANDN U34547 ( .A(n33340), .B(n33339), .Z(n33583) );
  XOR U34548 ( .A(n33584), .B(n33583), .Z(n33585) );
  NAND U34549 ( .A(n33342), .B(n33341), .Z(n33346) );
  NAND U34550 ( .A(n33344), .B(n33343), .Z(n33345) );
  NAND U34551 ( .A(n33346), .B(n33345), .Z(n33482) );
  AND U34552 ( .A(x[503]), .B(y[8006]), .Z(n33512) );
  AND U34553 ( .A(x[493]), .B(y[8016]), .Z(n33510) );
  AND U34554 ( .A(x[504]), .B(y[8005]), .Z(n33751) );
  XOR U34555 ( .A(n33510), .B(n33751), .Z(n33511) );
  XOR U34556 ( .A(n33512), .B(n33511), .Z(n33481) );
  AND U34557 ( .A(x[491]), .B(y[8018]), .Z(n33518) );
  AND U34558 ( .A(x[483]), .B(y[8026]), .Z(n33516) );
  AND U34559 ( .A(x[497]), .B(y[8012]), .Z(n33515) );
  XOR U34560 ( .A(n33516), .B(n33515), .Z(n33517) );
  XOR U34561 ( .A(n33518), .B(n33517), .Z(n33480) );
  XOR U34562 ( .A(n33481), .B(n33480), .Z(n33483) );
  XNOR U34563 ( .A(n33482), .B(n33483), .Z(n33586) );
  NAND U34564 ( .A(n33521), .B(n33347), .Z(n33351) );
  NAND U34565 ( .A(n33349), .B(n33348), .Z(n33350) );
  NAND U34566 ( .A(n33351), .B(n33350), .Z(n33592) );
  AND U34567 ( .A(x[505]), .B(y[8004]), .Z(n33537) );
  AND U34568 ( .A(x[506]), .B(y[8003]), .Z(n33534) );
  XOR U34569 ( .A(n33535), .B(n33534), .Z(n33536) );
  XOR U34570 ( .A(n33537), .B(n33536), .Z(n33590) );
  AND U34571 ( .A(x[508]), .B(y[8001]), .Z(n33552) );
  XOR U34572 ( .A(o[349]), .B(n33552), .Z(n33600) );
  AND U34573 ( .A(x[480]), .B(y[8029]), .Z(n33598) );
  AND U34574 ( .A(x[509]), .B(y[8000]), .Z(n33597) );
  XOR U34575 ( .A(n33598), .B(n33597), .Z(n33599) );
  XNOR U34576 ( .A(n33600), .B(n33599), .Z(n33589) );
  XOR U34577 ( .A(n33592), .B(n33591), .Z(n33559) );
  NAND U34578 ( .A(n33353), .B(n33352), .Z(n33357) );
  NAND U34579 ( .A(n33355), .B(n33354), .Z(n33356) );
  NAND U34580 ( .A(n33357), .B(n33356), .Z(n33530) );
  AND U34581 ( .A(o[348]), .B(n33358), .Z(n33489) );
  AND U34582 ( .A(x[496]), .B(y[8013]), .Z(n33487) );
  AND U34583 ( .A(x[507]), .B(y[8002]), .Z(n33486) );
  XOR U34584 ( .A(n33487), .B(n33486), .Z(n33488) );
  XOR U34585 ( .A(n33489), .B(n33488), .Z(n33529) );
  AND U34586 ( .A(x[482]), .B(y[8027]), .Z(n33498) );
  XOR U34587 ( .A(n33501), .B(n33500), .Z(n33528) );
  XOR U34588 ( .A(n33529), .B(n33528), .Z(n33531) );
  XOR U34589 ( .A(n33530), .B(n33531), .Z(n33560) );
  NANDN U34590 ( .A(n33360), .B(n33359), .Z(n33364) );
  NAND U34591 ( .A(n33362), .B(n33361), .Z(n33363) );
  NAND U34592 ( .A(n33364), .B(n33363), .Z(n33474) );
  NAND U34593 ( .A(n33366), .B(n33365), .Z(n33370) );
  NAND U34594 ( .A(n33368), .B(n33367), .Z(n33369) );
  NAND U34595 ( .A(n33370), .B(n33369), .Z(n33505) );
  NAND U34596 ( .A(n33372), .B(n33371), .Z(n33376) );
  NAND U34597 ( .A(n33374), .B(n33373), .Z(n33375) );
  NAND U34598 ( .A(n33376), .B(n33375), .Z(n33504) );
  XOR U34599 ( .A(n33505), .B(n33504), .Z(n33506) );
  AND U34600 ( .A(x[488]), .B(y[8021]), .Z(n33523) );
  AND U34601 ( .A(y[8023]), .B(x[486]), .Z(n33378) );
  NAND U34602 ( .A(y[8022]), .B(x[487]), .Z(n33377) );
  XNOR U34603 ( .A(n33378), .B(n33377), .Z(n33522) );
  XOR U34604 ( .A(n33523), .B(n33522), .Z(n33595) );
  AND U34605 ( .A(x[485]), .B(y[8024]), .Z(n33495) );
  AND U34606 ( .A(x[484]), .B(y[8025]), .Z(n33493) );
  AND U34607 ( .A(x[490]), .B(y[8019]), .Z(n33492) );
  XOR U34608 ( .A(n33493), .B(n33492), .Z(n33494) );
  XOR U34609 ( .A(n33495), .B(n33494), .Z(n33596) );
  AND U34610 ( .A(x[489]), .B(y[8020]), .Z(n33758) );
  XNOR U34611 ( .A(n33476), .B(n33477), .Z(n33566) );
  NAND U34612 ( .A(n33380), .B(n33379), .Z(n33384) );
  NAND U34613 ( .A(n33382), .B(n33381), .Z(n33383) );
  NAND U34614 ( .A(n33384), .B(n33383), .Z(n33565) );
  XOR U34615 ( .A(n33462), .B(n33463), .Z(n33465) );
  NAND U34616 ( .A(n33386), .B(n33385), .Z(n33390) );
  NAND U34617 ( .A(n33388), .B(n33387), .Z(n33389) );
  NAND U34618 ( .A(n33390), .B(n33389), .Z(n33456) );
  NANDN U34619 ( .A(n33392), .B(n33391), .Z(n33396) );
  NANDN U34620 ( .A(n33394), .B(n33393), .Z(n33395) );
  AND U34621 ( .A(n33396), .B(n33395), .Z(n33457) );
  XOR U34622 ( .A(n33456), .B(n33457), .Z(n33459) );
  NAND U34623 ( .A(n33398), .B(n33397), .Z(n33402) );
  NAND U34624 ( .A(n33400), .B(n33399), .Z(n33401) );
  NAND U34625 ( .A(n33402), .B(n33401), .Z(n33470) );
  NANDN U34626 ( .A(n33404), .B(n33403), .Z(n33408) );
  NAND U34627 ( .A(n33406), .B(n33405), .Z(n33407) );
  NAND U34628 ( .A(n33408), .B(n33407), .Z(n33468) );
  NAND U34629 ( .A(n33410), .B(n33409), .Z(n33414) );
  NAND U34630 ( .A(n33412), .B(n33411), .Z(n33413) );
  NAND U34631 ( .A(n33414), .B(n33413), .Z(n33555) );
  NAND U34632 ( .A(n33416), .B(n33415), .Z(n33420) );
  NAND U34633 ( .A(n33418), .B(n33417), .Z(n33419) );
  NAND U34634 ( .A(n33420), .B(n33419), .Z(n33554) );
  NAND U34635 ( .A(n33422), .B(n33421), .Z(n33426) );
  NAND U34636 ( .A(n33424), .B(n33423), .Z(n33425) );
  NAND U34637 ( .A(n33426), .B(n33425), .Z(n33553) );
  XOR U34638 ( .A(n33554), .B(n33553), .Z(n33556) );
  XOR U34639 ( .A(n33555), .B(n33556), .Z(n33469) );
  XOR U34640 ( .A(n33468), .B(n33469), .Z(n33471) );
  XOR U34641 ( .A(n33470), .B(n33471), .Z(n33458) );
  XOR U34642 ( .A(n33459), .B(n33458), .Z(n33464) );
  XOR U34643 ( .A(n33465), .B(n33464), .Z(n33452) );
  XOR U34644 ( .A(n33453), .B(n33452), .Z(n33445) );
  XNOR U34645 ( .A(n33444), .B(n33445), .Z(n33447) );
  XOR U34646 ( .A(n33446), .B(n33447), .Z(n33443) );
  NAND U34647 ( .A(n33428), .B(n33427), .Z(n33432) );
  NAND U34648 ( .A(n33430), .B(n33429), .Z(n33431) );
  NAND U34649 ( .A(n33432), .B(n33431), .Z(n33442) );
  NANDN U34650 ( .A(n33433), .B(n33434), .Z(n33439) );
  NOR U34651 ( .A(n33435), .B(n33434), .Z(n33437) );
  OR U34652 ( .A(n33437), .B(n33436), .Z(n33438) );
  AND U34653 ( .A(n33439), .B(n33438), .Z(n33441) );
  XOR U34654 ( .A(n33442), .B(n33441), .Z(n33440) );
  XNOR U34655 ( .A(n33443), .B(n33440), .Z(N702) );
  NAND U34656 ( .A(n33445), .B(n33444), .Z(n33449) );
  NANDN U34657 ( .A(n33447), .B(n33446), .Z(n33448) );
  NAND U34658 ( .A(n33449), .B(n33448), .Z(n33616) );
  NAND U34659 ( .A(n33451), .B(n33450), .Z(n33455) );
  NAND U34660 ( .A(n33453), .B(n33452), .Z(n33454) );
  NAND U34661 ( .A(n33455), .B(n33454), .Z(n33897) );
  NAND U34662 ( .A(n33457), .B(n33456), .Z(n33461) );
  NAND U34663 ( .A(n33459), .B(n33458), .Z(n33460) );
  AND U34664 ( .A(n33461), .B(n33460), .Z(n33906) );
  NAND U34665 ( .A(n33463), .B(n33462), .Z(n33467) );
  NAND U34666 ( .A(n33465), .B(n33464), .Z(n33466) );
  AND U34667 ( .A(n33467), .B(n33466), .Z(n33905) );
  XOR U34668 ( .A(n33906), .B(n33905), .Z(n33904) );
  NAND U34669 ( .A(n33469), .B(n33468), .Z(n33473) );
  NAND U34670 ( .A(n33471), .B(n33470), .Z(n33472) );
  AND U34671 ( .A(n33473), .B(n33472), .Z(n33903) );
  XNOR U34672 ( .A(n33904), .B(n33903), .Z(n33899) );
  NANDN U34673 ( .A(n33475), .B(n33474), .Z(n33479) );
  NANDN U34674 ( .A(n33477), .B(n33476), .Z(n33478) );
  AND U34675 ( .A(n33479), .B(n33478), .Z(n33619) );
  NAND U34676 ( .A(n33481), .B(n33480), .Z(n33485) );
  NAND U34677 ( .A(n33483), .B(n33482), .Z(n33484) );
  AND U34678 ( .A(n33485), .B(n33484), .Z(n33869) );
  NAND U34679 ( .A(n33487), .B(n33486), .Z(n33491) );
  NAND U34680 ( .A(n33489), .B(n33488), .Z(n33490) );
  NAND U34681 ( .A(n33491), .B(n33490), .Z(n33827) );
  NAND U34682 ( .A(n33493), .B(n33492), .Z(n33497) );
  NAND U34683 ( .A(n33495), .B(n33494), .Z(n33496) );
  NAND U34684 ( .A(n33497), .B(n33496), .Z(n33830) );
  AND U34685 ( .A(x[486]), .B(y[8024]), .Z(n33670) );
  AND U34686 ( .A(x[485]), .B(y[8025]), .Z(n33672) );
  AND U34687 ( .A(x[499]), .B(y[8011]), .Z(n33671) );
  XOR U34688 ( .A(n33672), .B(n33671), .Z(n33669) );
  XNOR U34689 ( .A(n33670), .B(n33669), .Z(n33637) );
  AND U34690 ( .A(x[484]), .B(y[8026]), .Z(n33708) );
  AND U34691 ( .A(x[483]), .B(y[8027]), .Z(n33710) );
  AND U34692 ( .A(x[498]), .B(y[8012]), .Z(n33709) );
  XOR U34693 ( .A(n33710), .B(n33709), .Z(n33707) );
  XOR U34694 ( .A(n33708), .B(n33707), .Z(n33640) );
  NANDN U34695 ( .A(n33499), .B(n33498), .Z(n33503) );
  NAND U34696 ( .A(n33501), .B(n33500), .Z(n33502) );
  AND U34697 ( .A(n33503), .B(n33502), .Z(n33639) );
  XOR U34698 ( .A(n33637), .B(n33638), .Z(n33829) );
  XOR U34699 ( .A(n33830), .B(n33829), .Z(n33828) );
  XOR U34700 ( .A(n33827), .B(n33828), .Z(n33870) );
  NAND U34701 ( .A(n33505), .B(n33504), .Z(n33509) );
  NANDN U34702 ( .A(n33507), .B(n33506), .Z(n33508) );
  AND U34703 ( .A(n33509), .B(n33508), .Z(n33867) );
  XOR U34704 ( .A(n33868), .B(n33867), .Z(n33622) );
  NAND U34705 ( .A(n33510), .B(n33751), .Z(n33514) );
  NAND U34706 ( .A(n33512), .B(n33511), .Z(n33513) );
  NAND U34707 ( .A(n33514), .B(n33513), .Z(n33852) );
  NAND U34708 ( .A(n33516), .B(n33515), .Z(n33520) );
  NAND U34709 ( .A(n33518), .B(n33517), .Z(n33519) );
  AND U34710 ( .A(n33520), .B(n33519), .Z(n33658) );
  AND U34711 ( .A(x[480]), .B(y[8030]), .Z(n33738) );
  AND U34712 ( .A(x[509]), .B(y[8001]), .Z(n33761) );
  XOR U34713 ( .A(o[350]), .B(n33761), .Z(n33740) );
  AND U34714 ( .A(x[510]), .B(y[8000]), .Z(n33739) );
  XOR U34715 ( .A(n33740), .B(n33739), .Z(n33737) );
  XOR U34716 ( .A(n33738), .B(n33737), .Z(n33660) );
  AND U34717 ( .A(x[500]), .B(y[8010]), .Z(n33698) );
  XOR U34718 ( .A(n33699), .B(n33698), .Z(n33697) );
  AND U34719 ( .A(x[488]), .B(y[8022]), .Z(n33696) );
  XNOR U34720 ( .A(n33697), .B(n33696), .Z(n33659) );
  XNOR U34721 ( .A(n33658), .B(n33657), .Z(n33851) );
  XOR U34722 ( .A(n33852), .B(n33851), .Z(n33849) );
  AND U34723 ( .A(x[487]), .B(y[8023]), .Z(n33703) );
  NAND U34724 ( .A(n33521), .B(n33703), .Z(n33525) );
  NAND U34725 ( .A(n33523), .B(n33522), .Z(n33524) );
  AND U34726 ( .A(n33525), .B(n33524), .Z(n33666) );
  AND U34727 ( .A(y[8009]), .B(x[501]), .Z(n33527) );
  AND U34728 ( .A(y[8008]), .B(x[502]), .Z(n33526) );
  XOR U34729 ( .A(n33527), .B(n33526), .Z(n33702) );
  XNOR U34730 ( .A(n33703), .B(n33702), .Z(n33664) );
  AND U34731 ( .A(x[497]), .B(y[8013]), .Z(n33689) );
  AND U34732 ( .A(x[482]), .B(y[8028]), .Z(n33691) );
  AND U34733 ( .A(x[506]), .B(y[8004]), .Z(n33690) );
  XOR U34734 ( .A(n33691), .B(n33690), .Z(n33688) );
  XOR U34735 ( .A(n33689), .B(n33688), .Z(n33663) );
  XNOR U34736 ( .A(n33666), .B(n33665), .Z(n33850) );
  NAND U34737 ( .A(n33529), .B(n33528), .Z(n33533) );
  NAND U34738 ( .A(n33531), .B(n33530), .Z(n33532) );
  NAND U34739 ( .A(n33533), .B(n33532), .Z(n33863) );
  XOR U34740 ( .A(n33864), .B(n33863), .Z(n33862) );
  AND U34741 ( .A(n33535), .B(n33534), .Z(n33539) );
  NAND U34742 ( .A(n33537), .B(n33536), .Z(n33538) );
  NANDN U34743 ( .A(n33539), .B(n33538), .Z(n33821) );
  AND U34744 ( .A(n33675), .B(n33540), .Z(n33544) );
  NAND U34745 ( .A(n33542), .B(n33541), .Z(n33543) );
  NANDN U34746 ( .A(n33544), .B(n33543), .Z(n33824) );
  NANDN U34747 ( .A(n33704), .B(n33545), .Z(n33549) );
  NANDN U34748 ( .A(n33547), .B(n33546), .Z(n33548) );
  AND U34749 ( .A(n33549), .B(n33548), .Z(n33650) );
  AND U34750 ( .A(x[503]), .B(y[8007]), .Z(n33750) );
  AND U34751 ( .A(y[8006]), .B(x[504]), .Z(n33551) );
  AND U34752 ( .A(y[8005]), .B(x[505]), .Z(n33550) );
  XOR U34753 ( .A(n33551), .B(n33550), .Z(n33749) );
  XOR U34754 ( .A(n33750), .B(n33749), .Z(n33652) );
  AND U34755 ( .A(n33552), .B(o[349]), .Z(n33683) );
  AND U34756 ( .A(x[508]), .B(y[8002]), .Z(n33685) );
  AND U34757 ( .A(x[496]), .B(y[8014]), .Z(n33684) );
  XOR U34758 ( .A(n33685), .B(n33684), .Z(n33682) );
  XNOR U34759 ( .A(n33683), .B(n33682), .Z(n33651) );
  XNOR U34760 ( .A(n33650), .B(n33649), .Z(n33823) );
  XOR U34761 ( .A(n33824), .B(n33823), .Z(n33822) );
  XOR U34762 ( .A(n33821), .B(n33822), .Z(n33861) );
  XOR U34763 ( .A(n33862), .B(n33861), .Z(n33621) );
  XOR U34764 ( .A(n33619), .B(n33620), .Z(n33886) );
  NAND U34765 ( .A(n33554), .B(n33553), .Z(n33558) );
  NAND U34766 ( .A(n33556), .B(n33555), .Z(n33557) );
  AND U34767 ( .A(n33558), .B(n33557), .Z(n33888) );
  NANDN U34768 ( .A(n33560), .B(n33559), .Z(n33564) );
  NANDN U34769 ( .A(n33562), .B(n33561), .Z(n33563) );
  NAND U34770 ( .A(n33564), .B(n33563), .Z(n33887) );
  XOR U34771 ( .A(n33888), .B(n33887), .Z(n33885) );
  XNOR U34772 ( .A(n33886), .B(n33885), .Z(n33879) );
  NANDN U34773 ( .A(n33566), .B(n33565), .Z(n33570) );
  NANDN U34774 ( .A(n33568), .B(n33567), .Z(n33569) );
  NAND U34775 ( .A(n33570), .B(n33569), .Z(n33881) );
  NANDN U34776 ( .A(n33572), .B(n33571), .Z(n33576) );
  NAND U34777 ( .A(n33574), .B(n33573), .Z(n33575) );
  AND U34778 ( .A(n33576), .B(n33575), .Z(n33626) );
  NAND U34779 ( .A(n33578), .B(n33577), .Z(n33582) );
  NAND U34780 ( .A(n33580), .B(n33579), .Z(n33581) );
  AND U34781 ( .A(n33582), .B(n33581), .Z(n33634) );
  NAND U34782 ( .A(n33584), .B(n33583), .Z(n33588) );
  NANDN U34783 ( .A(n33586), .B(n33585), .Z(n33587) );
  AND U34784 ( .A(n33588), .B(n33587), .Z(n33633) );
  XOR U34785 ( .A(n33634), .B(n33633), .Z(n33632) );
  NANDN U34786 ( .A(n33590), .B(n33589), .Z(n33594) );
  OR U34787 ( .A(n33592), .B(n33591), .Z(n33593) );
  NAND U34788 ( .A(n33594), .B(n33593), .Z(n33631) );
  XOR U34789 ( .A(n33632), .B(n33631), .Z(n33628) );
  NAND U34790 ( .A(n33598), .B(n33597), .Z(n33602) );
  NAND U34791 ( .A(n33600), .B(n33599), .Z(n33601) );
  NAND U34792 ( .A(n33602), .B(n33601), .Z(n33643) );
  AND U34793 ( .A(y[8018]), .B(x[492]), .Z(n33603) );
  XOR U34794 ( .A(n33604), .B(n33603), .Z(n33676) );
  XOR U34795 ( .A(n33677), .B(n33676), .Z(n33757) );
  AND U34796 ( .A(y[8021]), .B(x[489]), .Z(n33606) );
  XOR U34797 ( .A(n33606), .B(n33605), .Z(n33756) );
  XOR U34798 ( .A(n33757), .B(n33756), .Z(n33646) );
  AND U34799 ( .A(x[507]), .B(y[8003]), .Z(n33746) );
  AND U34800 ( .A(x[481]), .B(y[8029]), .Z(n33745) );
  XOR U34801 ( .A(n33746), .B(n33745), .Z(n33743) );
  XOR U34802 ( .A(n33744), .B(n33743), .Z(n33645) );
  XOR U34803 ( .A(n33646), .B(n33645), .Z(n33644) );
  XOR U34804 ( .A(n33643), .B(n33644), .Z(n33846) );
  NAND U34805 ( .A(n33608), .B(n33607), .Z(n33612) );
  NANDN U34806 ( .A(n33610), .B(n33609), .Z(n33611) );
  AND U34807 ( .A(n33612), .B(n33611), .Z(n33843) );
  XNOR U34808 ( .A(n33844), .B(n33843), .Z(n33627) );
  XOR U34809 ( .A(n33626), .B(n33625), .Z(n33882) );
  XNOR U34810 ( .A(n33881), .B(n33882), .Z(n33880) );
  XOR U34811 ( .A(n33899), .B(n33900), .Z(n33898) );
  XOR U34812 ( .A(n33897), .B(n33898), .Z(n33613) );
  XNOR U34813 ( .A(n33614), .B(n33613), .Z(N703) );
  NAND U34814 ( .A(n33614), .B(n33613), .Z(n33618) );
  NANDN U34815 ( .A(n33616), .B(n33615), .Z(n33617) );
  AND U34816 ( .A(n33618), .B(n33617), .Z(n33914) );
  NANDN U34817 ( .A(n33620), .B(n33619), .Z(n33624) );
  NANDN U34818 ( .A(n33622), .B(n33621), .Z(n33623) );
  AND U34819 ( .A(n33624), .B(n33623), .Z(n33896) );
  NAND U34820 ( .A(n33626), .B(n33625), .Z(n33630) );
  NANDN U34821 ( .A(n33628), .B(n33627), .Z(n33629) );
  AND U34822 ( .A(n33630), .B(n33629), .Z(n33878) );
  NAND U34823 ( .A(n33632), .B(n33631), .Z(n33636) );
  NAND U34824 ( .A(n33634), .B(n33633), .Z(n33635) );
  AND U34825 ( .A(n33636), .B(n33635), .Z(n33860) );
  NANDN U34826 ( .A(n33638), .B(n33637), .Z(n33642) );
  NANDN U34827 ( .A(n33640), .B(n33639), .Z(n33641) );
  AND U34828 ( .A(n33642), .B(n33641), .Z(n33842) );
  NAND U34829 ( .A(n33644), .B(n33643), .Z(n33648) );
  NAND U34830 ( .A(n33646), .B(n33645), .Z(n33647) );
  AND U34831 ( .A(n33648), .B(n33647), .Z(n33656) );
  NAND U34832 ( .A(n33650), .B(n33649), .Z(n33654) );
  NANDN U34833 ( .A(n33652), .B(n33651), .Z(n33653) );
  NAND U34834 ( .A(n33654), .B(n33653), .Z(n33655) );
  XNOR U34835 ( .A(n33656), .B(n33655), .Z(n33840) );
  NAND U34836 ( .A(n33658), .B(n33657), .Z(n33662) );
  NANDN U34837 ( .A(n33660), .B(n33659), .Z(n33661) );
  AND U34838 ( .A(n33662), .B(n33661), .Z(n33838) );
  ANDN U34839 ( .B(n33664), .A(n33663), .Z(n33668) );
  ANDN U34840 ( .B(n33666), .A(n33665), .Z(n33667) );
  NOR U34841 ( .A(n33668), .B(n33667), .Z(n33820) );
  NAND U34842 ( .A(n33670), .B(n33669), .Z(n33674) );
  NAND U34843 ( .A(n33672), .B(n33671), .Z(n33673) );
  AND U34844 ( .A(n33674), .B(n33673), .Z(n33681) );
  NAND U34845 ( .A(n33675), .B(n33786), .Z(n33679) );
  NAND U34846 ( .A(n33677), .B(n33676), .Z(n33678) );
  AND U34847 ( .A(n33679), .B(n33678), .Z(n33680) );
  XNOR U34848 ( .A(n33681), .B(n33680), .Z(n33736) );
  NAND U34849 ( .A(n33683), .B(n33682), .Z(n33687) );
  NAND U34850 ( .A(n33685), .B(n33684), .Z(n33686) );
  AND U34851 ( .A(n33687), .B(n33686), .Z(n33695) );
  NAND U34852 ( .A(n33689), .B(n33688), .Z(n33693) );
  NAND U34853 ( .A(n33691), .B(n33690), .Z(n33692) );
  NAND U34854 ( .A(n33693), .B(n33692), .Z(n33694) );
  XNOR U34855 ( .A(n33695), .B(n33694), .Z(n33734) );
  NAND U34856 ( .A(n33697), .B(n33696), .Z(n33701) );
  NAND U34857 ( .A(n33699), .B(n33698), .Z(n33700) );
  AND U34858 ( .A(n33701), .B(n33700), .Z(n33732) );
  NAND U34859 ( .A(n33703), .B(n33702), .Z(n33706) );
  AND U34860 ( .A(x[502]), .B(y[8009]), .Z(n33763) );
  NANDN U34861 ( .A(n33704), .B(n33763), .Z(n33705) );
  AND U34862 ( .A(n33706), .B(n33705), .Z(n33714) );
  NAND U34863 ( .A(n33708), .B(n33707), .Z(n33712) );
  NAND U34864 ( .A(n33710), .B(n33709), .Z(n33711) );
  NAND U34865 ( .A(n33712), .B(n33711), .Z(n33713) );
  XNOR U34866 ( .A(n33714), .B(n33713), .Z(n33730) );
  AND U34867 ( .A(y[8030]), .B(x[481]), .Z(n33716) );
  NAND U34868 ( .A(y[8031]), .B(x[480]), .Z(n33715) );
  XNOR U34869 ( .A(n33716), .B(n33715), .Z(n33720) );
  AND U34870 ( .A(y[8019]), .B(x[492]), .Z(n33718) );
  NAND U34871 ( .A(y[8003]), .B(x[508]), .Z(n33717) );
  XNOR U34872 ( .A(n33718), .B(n33717), .Z(n33719) );
  XOR U34873 ( .A(n33720), .B(n33719), .Z(n33728) );
  AND U34874 ( .A(y[8004]), .B(x[507]), .Z(n33722) );
  NAND U34875 ( .A(y[8027]), .B(x[484]), .Z(n33721) );
  XNOR U34876 ( .A(n33722), .B(n33721), .Z(n33726) );
  AND U34877 ( .A(y[8000]), .B(x[511]), .Z(n33724) );
  NAND U34878 ( .A(y[8013]), .B(x[498]), .Z(n33723) );
  XNOR U34879 ( .A(n33724), .B(n33723), .Z(n33725) );
  XNOR U34880 ( .A(n33726), .B(n33725), .Z(n33727) );
  XNOR U34881 ( .A(n33728), .B(n33727), .Z(n33729) );
  XNOR U34882 ( .A(n33730), .B(n33729), .Z(n33731) );
  XNOR U34883 ( .A(n33732), .B(n33731), .Z(n33733) );
  XNOR U34884 ( .A(n33734), .B(n33733), .Z(n33735) );
  XNOR U34885 ( .A(n33736), .B(n33735), .Z(n33818) );
  NAND U34886 ( .A(n33738), .B(n33737), .Z(n33742) );
  NAND U34887 ( .A(n33740), .B(n33739), .Z(n33741) );
  AND U34888 ( .A(n33742), .B(n33741), .Z(n33816) );
  NAND U34889 ( .A(n33744), .B(n33743), .Z(n33748) );
  NAND U34890 ( .A(n33746), .B(n33745), .Z(n33747) );
  AND U34891 ( .A(n33748), .B(n33747), .Z(n33755) );
  NAND U34892 ( .A(n33750), .B(n33749), .Z(n33753) );
  AND U34893 ( .A(x[505]), .B(y[8006]), .Z(n33762) );
  NAND U34894 ( .A(n33751), .B(n33762), .Z(n33752) );
  NAND U34895 ( .A(n33753), .B(n33752), .Z(n33754) );
  XNOR U34896 ( .A(n33755), .B(n33754), .Z(n33814) );
  NAND U34897 ( .A(n33757), .B(n33756), .Z(n33760) );
  AND U34898 ( .A(x[490]), .B(y[8021]), .Z(n33785) );
  NAND U34899 ( .A(n33758), .B(n33785), .Z(n33759) );
  AND U34900 ( .A(n33760), .B(n33759), .Z(n33812) );
  AND U34901 ( .A(y[8012]), .B(x[499]), .Z(n33770) );
  AND U34902 ( .A(n33761), .B(o[350]), .Z(n33768) );
  XOR U34903 ( .A(n33762), .B(o[351]), .Z(n33766) );
  XNOR U34904 ( .A(n33764), .B(n33763), .Z(n33765) );
  XNOR U34905 ( .A(n33766), .B(n33765), .Z(n33767) );
  XNOR U34906 ( .A(n33768), .B(n33767), .Z(n33769) );
  XNOR U34907 ( .A(n33770), .B(n33769), .Z(n33810) );
  AND U34908 ( .A(y[8001]), .B(x[510]), .Z(n33776) );
  AND U34909 ( .A(y[8020]), .B(x[491]), .Z(n33772) );
  NAND U34910 ( .A(y[8005]), .B(x[506]), .Z(n33771) );
  XNOR U34911 ( .A(n33772), .B(n33771), .Z(n33773) );
  XNOR U34912 ( .A(n33774), .B(n33773), .Z(n33775) );
  XNOR U34913 ( .A(n33776), .B(n33775), .Z(n33800) );
  AND U34914 ( .A(y[8010]), .B(x[501]), .Z(n33778) );
  NAND U34915 ( .A(y[8023]), .B(x[488]), .Z(n33777) );
  XNOR U34916 ( .A(n33778), .B(n33777), .Z(n33790) );
  AND U34917 ( .A(y[8008]), .B(x[503]), .Z(n33780) );
  NAND U34918 ( .A(y[8014]), .B(x[497]), .Z(n33779) );
  XNOR U34919 ( .A(n33780), .B(n33779), .Z(n33784) );
  AND U34920 ( .A(y[8017]), .B(x[494]), .Z(n33782) );
  NAND U34921 ( .A(y[8029]), .B(x[482]), .Z(n33781) );
  XNOR U34922 ( .A(n33782), .B(n33781), .Z(n33783) );
  XOR U34923 ( .A(n33784), .B(n33783), .Z(n33788) );
  XNOR U34924 ( .A(n33786), .B(n33785), .Z(n33787) );
  XNOR U34925 ( .A(n33788), .B(n33787), .Z(n33789) );
  XOR U34926 ( .A(n33790), .B(n33789), .Z(n33798) );
  AND U34927 ( .A(y[8026]), .B(x[485]), .Z(n33792) );
  NAND U34928 ( .A(y[8024]), .B(x[487]), .Z(n33791) );
  XNOR U34929 ( .A(n33792), .B(n33791), .Z(n33796) );
  AND U34930 ( .A(y[8025]), .B(x[486]), .Z(n33794) );
  NAND U34931 ( .A(y[8028]), .B(x[483]), .Z(n33793) );
  XNOR U34932 ( .A(n33794), .B(n33793), .Z(n33795) );
  XNOR U34933 ( .A(n33796), .B(n33795), .Z(n33797) );
  XNOR U34934 ( .A(n33798), .B(n33797), .Z(n33799) );
  XOR U34935 ( .A(n33800), .B(n33799), .Z(n33808) );
  AND U34936 ( .A(y[8015]), .B(x[496]), .Z(n33802) );
  NAND U34937 ( .A(y[8022]), .B(x[489]), .Z(n33801) );
  XNOR U34938 ( .A(n33802), .B(n33801), .Z(n33806) );
  AND U34939 ( .A(y[8002]), .B(x[509]), .Z(n33804) );
  NAND U34940 ( .A(y[8011]), .B(x[500]), .Z(n33803) );
  XNOR U34941 ( .A(n33804), .B(n33803), .Z(n33805) );
  XNOR U34942 ( .A(n33806), .B(n33805), .Z(n33807) );
  XNOR U34943 ( .A(n33808), .B(n33807), .Z(n33809) );
  XNOR U34944 ( .A(n33810), .B(n33809), .Z(n33811) );
  XNOR U34945 ( .A(n33812), .B(n33811), .Z(n33813) );
  XNOR U34946 ( .A(n33814), .B(n33813), .Z(n33815) );
  XNOR U34947 ( .A(n33816), .B(n33815), .Z(n33817) );
  XOR U34948 ( .A(n33818), .B(n33817), .Z(n33819) );
  XNOR U34949 ( .A(n33820), .B(n33819), .Z(n33836) );
  NAND U34950 ( .A(n33822), .B(n33821), .Z(n33826) );
  NAND U34951 ( .A(n33824), .B(n33823), .Z(n33825) );
  AND U34952 ( .A(n33826), .B(n33825), .Z(n33834) );
  NAND U34953 ( .A(n33828), .B(n33827), .Z(n33832) );
  NAND U34954 ( .A(n33830), .B(n33829), .Z(n33831) );
  NAND U34955 ( .A(n33832), .B(n33831), .Z(n33833) );
  XNOR U34956 ( .A(n33834), .B(n33833), .Z(n33835) );
  XNOR U34957 ( .A(n33836), .B(n33835), .Z(n33837) );
  XNOR U34958 ( .A(n33838), .B(n33837), .Z(n33839) );
  XNOR U34959 ( .A(n33840), .B(n33839), .Z(n33841) );
  XNOR U34960 ( .A(n33842), .B(n33841), .Z(n33858) );
  NAND U34961 ( .A(n33844), .B(n33843), .Z(n33848) );
  NANDN U34962 ( .A(n33846), .B(n33845), .Z(n33847) );
  AND U34963 ( .A(n33848), .B(n33847), .Z(n33856) );
  NANDN U34964 ( .A(n33850), .B(n33849), .Z(n33854) );
  NAND U34965 ( .A(n33852), .B(n33851), .Z(n33853) );
  NAND U34966 ( .A(n33854), .B(n33853), .Z(n33855) );
  XNOR U34967 ( .A(n33856), .B(n33855), .Z(n33857) );
  XNOR U34968 ( .A(n33858), .B(n33857), .Z(n33859) );
  XNOR U34969 ( .A(n33860), .B(n33859), .Z(n33876) );
  NAND U34970 ( .A(n33862), .B(n33861), .Z(n33866) );
  NAND U34971 ( .A(n33864), .B(n33863), .Z(n33865) );
  AND U34972 ( .A(n33866), .B(n33865), .Z(n33874) );
  NAND U34973 ( .A(n33868), .B(n33867), .Z(n33872) );
  NANDN U34974 ( .A(n33870), .B(n33869), .Z(n33871) );
  NAND U34975 ( .A(n33872), .B(n33871), .Z(n33873) );
  XNOR U34976 ( .A(n33874), .B(n33873), .Z(n33875) );
  XNOR U34977 ( .A(n33876), .B(n33875), .Z(n33877) );
  XNOR U34978 ( .A(n33878), .B(n33877), .Z(n33894) );
  NANDN U34979 ( .A(n33880), .B(n33879), .Z(n33884) );
  NAND U34980 ( .A(n33882), .B(n33881), .Z(n33883) );
  AND U34981 ( .A(n33884), .B(n33883), .Z(n33892) );
  NAND U34982 ( .A(n33886), .B(n33885), .Z(n33890) );
  NAND U34983 ( .A(n33888), .B(n33887), .Z(n33889) );
  NAND U34984 ( .A(n33890), .B(n33889), .Z(n33891) );
  XNOR U34985 ( .A(n33892), .B(n33891), .Z(n33893) );
  XNOR U34986 ( .A(n33894), .B(n33893), .Z(n33895) );
  XNOR U34987 ( .A(n33896), .B(n33895), .Z(n33912) );
  NANDN U34988 ( .A(n33898), .B(n33897), .Z(n33902) );
  NANDN U34989 ( .A(n33900), .B(n33899), .Z(n33901) );
  AND U34990 ( .A(n33902), .B(n33901), .Z(n33910) );
  NAND U34991 ( .A(n33904), .B(n33903), .Z(n33908) );
  NAND U34992 ( .A(n33906), .B(n33905), .Z(n33907) );
  NAND U34993 ( .A(n33908), .B(n33907), .Z(n33909) );
  XNOR U34994 ( .A(n33910), .B(n33909), .Z(n33911) );
  XNOR U34995 ( .A(n33912), .B(n33911), .Z(n33913) );
  XNOR U34996 ( .A(n33914), .B(n33913), .Z(N704) );
  AND U34997 ( .A(x[480]), .B(y[8032]), .Z(n34561) );
  XOR U34998 ( .A(n34561), .B(o[352]), .Z(N737) );
  AND U34999 ( .A(x[481]), .B(y[8032]), .Z(n33923) );
  AND U35000 ( .A(x[480]), .B(y[8033]), .Z(n33922) );
  XNOR U35001 ( .A(n33922), .B(o[353]), .Z(n33915) );
  XNOR U35002 ( .A(n33923), .B(n33915), .Z(n33917) );
  NAND U35003 ( .A(n34561), .B(o[352]), .Z(n33916) );
  XNOR U35004 ( .A(n33917), .B(n33916), .Z(N738) );
  NANDN U35005 ( .A(n33923), .B(n33915), .Z(n33919) );
  NAND U35006 ( .A(n33917), .B(n33916), .Z(n33918) );
  AND U35007 ( .A(n33919), .B(n33918), .Z(n33929) );
  AND U35008 ( .A(x[480]), .B(y[8034]), .Z(n33936) );
  XNOR U35009 ( .A(n33936), .B(o[354]), .Z(n33928) );
  XNOR U35010 ( .A(n33929), .B(n33928), .Z(n33931) );
  AND U35011 ( .A(y[8032]), .B(x[482]), .Z(n33921) );
  NAND U35012 ( .A(y[8033]), .B(x[481]), .Z(n33920) );
  XNOR U35013 ( .A(n33921), .B(n33920), .Z(n33925) );
  AND U35014 ( .A(n33922), .B(o[353]), .Z(n33924) );
  XNOR U35015 ( .A(n33925), .B(n33924), .Z(n33930) );
  XNOR U35016 ( .A(n33931), .B(n33930), .Z(N739) );
  AND U35017 ( .A(x[482]), .B(y[8033]), .Z(n33943) );
  NAND U35018 ( .A(n33943), .B(n33923), .Z(n33927) );
  NAND U35019 ( .A(n33925), .B(n33924), .Z(n33926) );
  AND U35020 ( .A(n33927), .B(n33926), .Z(n33946) );
  NANDN U35021 ( .A(n33929), .B(n33928), .Z(n33933) );
  NAND U35022 ( .A(n33931), .B(n33930), .Z(n33932) );
  AND U35023 ( .A(n33933), .B(n33932), .Z(n33945) );
  XNOR U35024 ( .A(n33946), .B(n33945), .Z(n33948) );
  AND U35025 ( .A(x[481]), .B(y[8034]), .Z(n34051) );
  XOR U35026 ( .A(n33943), .B(o[355]), .Z(n33951) );
  XOR U35027 ( .A(n34051), .B(n33951), .Z(n33953) );
  AND U35028 ( .A(y[8032]), .B(x[483]), .Z(n33935) );
  NAND U35029 ( .A(y[8035]), .B(x[480]), .Z(n33934) );
  XNOR U35030 ( .A(n33935), .B(n33934), .Z(n33938) );
  AND U35031 ( .A(n33936), .B(o[354]), .Z(n33937) );
  XOR U35032 ( .A(n33938), .B(n33937), .Z(n33952) );
  XOR U35033 ( .A(n33953), .B(n33952), .Z(n33947) );
  XOR U35034 ( .A(n33948), .B(n33947), .Z(N740) );
  AND U35035 ( .A(x[483]), .B(y[8035]), .Z(n33995) );
  NAND U35036 ( .A(n34561), .B(n33995), .Z(n33940) );
  NAND U35037 ( .A(n33938), .B(n33937), .Z(n33939) );
  AND U35038 ( .A(n33940), .B(n33939), .Z(n33974) );
  AND U35039 ( .A(y[8036]), .B(x[480]), .Z(n33942) );
  NAND U35040 ( .A(y[8032]), .B(x[484]), .Z(n33941) );
  XNOR U35041 ( .A(n33942), .B(n33941), .Z(n33967) );
  AND U35042 ( .A(n33943), .B(o[355]), .Z(n33968) );
  XOR U35043 ( .A(n33967), .B(n33968), .Z(n33972) );
  AND U35044 ( .A(y[8034]), .B(x[482]), .Z(n34106) );
  NAND U35045 ( .A(y[8035]), .B(x[481]), .Z(n33944) );
  XNOR U35046 ( .A(n34106), .B(n33944), .Z(n33964) );
  AND U35047 ( .A(x[483]), .B(y[8033]), .Z(n33959) );
  XOR U35048 ( .A(o[356]), .B(n33959), .Z(n33963) );
  XOR U35049 ( .A(n33964), .B(n33963), .Z(n33971) );
  XOR U35050 ( .A(n33972), .B(n33971), .Z(n33973) );
  XOR U35051 ( .A(n33974), .B(n33973), .Z(n33979) );
  NANDN U35052 ( .A(n33946), .B(n33945), .Z(n33950) );
  NAND U35053 ( .A(n33948), .B(n33947), .Z(n33949) );
  NAND U35054 ( .A(n33950), .B(n33949), .Z(n33977) );
  NAND U35055 ( .A(n34051), .B(n33951), .Z(n33955) );
  NAND U35056 ( .A(n33953), .B(n33952), .Z(n33954) );
  NAND U35057 ( .A(n33955), .B(n33954), .Z(n33978) );
  XOR U35058 ( .A(n33977), .B(n33978), .Z(n33956) );
  XNOR U35059 ( .A(n33979), .B(n33956), .Z(N741) );
  AND U35060 ( .A(y[8032]), .B(x[485]), .Z(n33958) );
  NAND U35061 ( .A(y[8037]), .B(x[480]), .Z(n33957) );
  XNOR U35062 ( .A(n33958), .B(n33957), .Z(n33988) );
  AND U35063 ( .A(o[356]), .B(n33959), .Z(n33987) );
  XOR U35064 ( .A(n33988), .B(n33987), .Z(n33986) );
  NAND U35065 ( .A(x[482]), .B(y[8035]), .Z(n34059) );
  AND U35066 ( .A(y[8034]), .B(x[483]), .Z(n33961) );
  NAND U35067 ( .A(y[8036]), .B(x[481]), .Z(n33960) );
  XNOR U35068 ( .A(n33961), .B(n33960), .Z(n33982) );
  AND U35069 ( .A(x[484]), .B(y[8033]), .Z(n33993) );
  XOR U35070 ( .A(n33993), .B(o[357]), .Z(n33981) );
  XOR U35071 ( .A(n33982), .B(n33981), .Z(n33985) );
  XOR U35072 ( .A(n34059), .B(n33985), .Z(n33962) );
  XNOR U35073 ( .A(n33986), .B(n33962), .Z(n34003) );
  NANDN U35074 ( .A(n34059), .B(n34051), .Z(n33966) );
  NAND U35075 ( .A(n33964), .B(n33963), .Z(n33965) );
  NAND U35076 ( .A(n33966), .B(n33965), .Z(n34001) );
  AND U35077 ( .A(x[484]), .B(y[8036]), .Z(n34763) );
  NAND U35078 ( .A(n34763), .B(n34561), .Z(n33970) );
  NAND U35079 ( .A(n33968), .B(n33967), .Z(n33969) );
  NAND U35080 ( .A(n33970), .B(n33969), .Z(n34000) );
  XOR U35081 ( .A(n34001), .B(n34000), .Z(n34002) );
  XNOR U35082 ( .A(n34003), .B(n34002), .Z(n33999) );
  NAND U35083 ( .A(n33972), .B(n33971), .Z(n33976) );
  NANDN U35084 ( .A(n33974), .B(n33973), .Z(n33975) );
  NAND U35085 ( .A(n33976), .B(n33975), .Z(n33997) );
  XOR U35086 ( .A(n33997), .B(n33998), .Z(n33980) );
  XNOR U35087 ( .A(n33999), .B(n33980), .Z(N742) );
  AND U35088 ( .A(x[483]), .B(y[8036]), .Z(n34060) );
  NAND U35089 ( .A(n34060), .B(n34051), .Z(n33984) );
  NAND U35090 ( .A(n33982), .B(n33981), .Z(n33983) );
  NAND U35091 ( .A(n33984), .B(n33983), .Z(n34032) );
  XOR U35092 ( .A(n34032), .B(n34031), .Z(n34034) );
  AND U35093 ( .A(x[485]), .B(y[8037]), .Z(n34231) );
  NAND U35094 ( .A(n34561), .B(n34231), .Z(n33990) );
  NAND U35095 ( .A(n33988), .B(n33987), .Z(n33989) );
  NAND U35096 ( .A(n33990), .B(n33989), .Z(n34008) );
  AND U35097 ( .A(y[8032]), .B(x[486]), .Z(n33992) );
  NAND U35098 ( .A(y[8038]), .B(x[480]), .Z(n33991) );
  XNOR U35099 ( .A(n33992), .B(n33991), .Z(n34014) );
  AND U35100 ( .A(n33993), .B(o[357]), .Z(n34015) );
  XOR U35101 ( .A(n34014), .B(n34015), .Z(n34007) );
  XOR U35102 ( .A(n34008), .B(n34007), .Z(n34010) );
  NAND U35103 ( .A(y[8036]), .B(x[482]), .Z(n33994) );
  XNOR U35104 ( .A(n33995), .B(n33994), .Z(n34019) );
  AND U35105 ( .A(y[8037]), .B(x[481]), .Z(n34260) );
  NAND U35106 ( .A(y[8034]), .B(x[484]), .Z(n33996) );
  XNOR U35107 ( .A(n34260), .B(n33996), .Z(n34023) );
  AND U35108 ( .A(x[485]), .B(y[8033]), .Z(n34030) );
  XOR U35109 ( .A(o[358]), .B(n34030), .Z(n34022) );
  XOR U35110 ( .A(n34023), .B(n34022), .Z(n34018) );
  XOR U35111 ( .A(n34019), .B(n34018), .Z(n34009) );
  XOR U35112 ( .A(n34010), .B(n34009), .Z(n34033) );
  XOR U35113 ( .A(n34034), .B(n34033), .Z(n34040) );
  NAND U35114 ( .A(n34001), .B(n34000), .Z(n34005) );
  NAND U35115 ( .A(n34003), .B(n34002), .Z(n34004) );
  AND U35116 ( .A(n34005), .B(n34004), .Z(n34039) );
  IV U35117 ( .A(n34039), .Z(n34037) );
  XOR U35118 ( .A(n34038), .B(n34037), .Z(n34006) );
  XNOR U35119 ( .A(n34040), .B(n34006), .Z(N743) );
  NAND U35120 ( .A(n34008), .B(n34007), .Z(n34012) );
  NAND U35121 ( .A(n34010), .B(n34009), .Z(n34011) );
  AND U35122 ( .A(n34012), .B(n34011), .Z(n34082) );
  AND U35123 ( .A(y[8034]), .B(x[485]), .Z(n34142) );
  NAND U35124 ( .A(y[8038]), .B(x[481]), .Z(n34013) );
  XNOR U35125 ( .A(n34142), .B(n34013), .Z(n34053) );
  AND U35126 ( .A(x[486]), .B(y[8033]), .Z(n34056) );
  XOR U35127 ( .A(o[359]), .B(n34056), .Z(n34052) );
  XOR U35128 ( .A(n34053), .B(n34052), .Z(n34071) );
  AND U35129 ( .A(x[486]), .B(y[8038]), .Z(n34280) );
  NAND U35130 ( .A(n34561), .B(n34280), .Z(n34017) );
  NAND U35131 ( .A(n34015), .B(n34014), .Z(n34016) );
  AND U35132 ( .A(n34017), .B(n34016), .Z(n34070) );
  NANDN U35133 ( .A(n34059), .B(n34060), .Z(n34021) );
  NAND U35134 ( .A(n34019), .B(n34018), .Z(n34020) );
  NAND U35135 ( .A(n34021), .B(n34020), .Z(n34073) );
  AND U35136 ( .A(x[484]), .B(y[8037]), .Z(n34566) );
  NAND U35137 ( .A(n34566), .B(n34051), .Z(n34025) );
  NAND U35138 ( .A(n34023), .B(n34022), .Z(n34024) );
  AND U35139 ( .A(n34025), .B(n34024), .Z(n34048) );
  AND U35140 ( .A(y[8037]), .B(x[482]), .Z(n34027) );
  NAND U35141 ( .A(y[8035]), .B(x[484]), .Z(n34026) );
  XNOR U35142 ( .A(n34027), .B(n34026), .Z(n34061) );
  XNOR U35143 ( .A(n34061), .B(n34060), .Z(n34046) );
  AND U35144 ( .A(y[8032]), .B(x[487]), .Z(n34029) );
  NAND U35145 ( .A(y[8039]), .B(x[480]), .Z(n34028) );
  XNOR U35146 ( .A(n34029), .B(n34028), .Z(n34065) );
  AND U35147 ( .A(o[358]), .B(n34030), .Z(n34064) );
  XNOR U35148 ( .A(n34065), .B(n34064), .Z(n34045) );
  XOR U35149 ( .A(n34046), .B(n34045), .Z(n34047) );
  XOR U35150 ( .A(n34048), .B(n34047), .Z(n34079) );
  XOR U35151 ( .A(n34080), .B(n34079), .Z(n34081) );
  XOR U35152 ( .A(n34082), .B(n34081), .Z(n34078) );
  NAND U35153 ( .A(n34032), .B(n34031), .Z(n34036) );
  NAND U35154 ( .A(n34034), .B(n34033), .Z(n34035) );
  NAND U35155 ( .A(n34036), .B(n34035), .Z(n34077) );
  NANDN U35156 ( .A(n34037), .B(n34038), .Z(n34043) );
  NOR U35157 ( .A(n34039), .B(n34038), .Z(n34041) );
  OR U35158 ( .A(n34041), .B(n34040), .Z(n34042) );
  AND U35159 ( .A(n34043), .B(n34042), .Z(n34076) );
  XOR U35160 ( .A(n34077), .B(n34076), .Z(n34044) );
  XNOR U35161 ( .A(n34078), .B(n34044), .Z(N744) );
  NAND U35162 ( .A(n34046), .B(n34045), .Z(n34050) );
  NAND U35163 ( .A(n34048), .B(n34047), .Z(n34049) );
  AND U35164 ( .A(n34050), .B(n34049), .Z(n34119) );
  AND U35165 ( .A(x[485]), .B(y[8038]), .Z(n34222) );
  NAND U35166 ( .A(n34051), .B(n34222), .Z(n34055) );
  NAND U35167 ( .A(n34053), .B(n34052), .Z(n34054) );
  NAND U35168 ( .A(n34055), .B(n34054), .Z(n34117) );
  AND U35169 ( .A(o[359]), .B(n34056), .Z(n34097) );
  AND U35170 ( .A(y[8035]), .B(x[485]), .Z(n34670) );
  NAND U35171 ( .A(y[8039]), .B(x[481]), .Z(n34057) );
  XNOR U35172 ( .A(n34670), .B(n34057), .Z(n34098) );
  XNOR U35173 ( .A(n34097), .B(n34098), .Z(n34102) );
  NAND U35174 ( .A(x[483]), .B(y[8037]), .Z(n34897) );
  AND U35175 ( .A(y[8034]), .B(x[486]), .Z(n34058) );
  AND U35176 ( .A(y[8038]), .B(x[482]), .Z(n34978) );
  XOR U35177 ( .A(n34058), .B(n34978), .Z(n34107) );
  XOR U35178 ( .A(n34763), .B(n34107), .Z(n34101) );
  XOR U35179 ( .A(n34102), .B(n34103), .Z(n34116) );
  XOR U35180 ( .A(n34117), .B(n34116), .Z(n34118) );
  XOR U35181 ( .A(n34119), .B(n34118), .Z(n34125) );
  NANDN U35182 ( .A(n34059), .B(n34566), .Z(n34063) );
  NAND U35183 ( .A(n34061), .B(n34060), .Z(n34062) );
  NAND U35184 ( .A(n34063), .B(n34062), .Z(n34113) );
  AND U35185 ( .A(x[487]), .B(y[8039]), .Z(n34444) );
  NAND U35186 ( .A(n34561), .B(n34444), .Z(n34067) );
  NAND U35187 ( .A(n34065), .B(n34064), .Z(n34066) );
  NAND U35188 ( .A(n34067), .B(n34066), .Z(n34111) );
  AND U35189 ( .A(y[8032]), .B(x[488]), .Z(n34069) );
  NAND U35190 ( .A(y[8040]), .B(x[480]), .Z(n34068) );
  XNOR U35191 ( .A(n34069), .B(n34068), .Z(n34088) );
  AND U35192 ( .A(x[487]), .B(y[8033]), .Z(n34091) );
  XOR U35193 ( .A(o[360]), .B(n34091), .Z(n34087) );
  XOR U35194 ( .A(n34088), .B(n34087), .Z(n34110) );
  XOR U35195 ( .A(n34111), .B(n34110), .Z(n34112) );
  XNOR U35196 ( .A(n34113), .B(n34112), .Z(n34123) );
  NANDN U35197 ( .A(n34071), .B(n34070), .Z(n34075) );
  NANDN U35198 ( .A(n34073), .B(n34072), .Z(n34074) );
  NAND U35199 ( .A(n34075), .B(n34074), .Z(n34122) );
  XOR U35200 ( .A(n34123), .B(n34122), .Z(n34124) );
  XOR U35201 ( .A(n34125), .B(n34124), .Z(n34131) );
  NAND U35202 ( .A(n34080), .B(n34079), .Z(n34084) );
  NAND U35203 ( .A(n34082), .B(n34081), .Z(n34083) );
  NAND U35204 ( .A(n34084), .B(n34083), .Z(n34130) );
  IV U35205 ( .A(n34130), .Z(n34128) );
  XOR U35206 ( .A(n34129), .B(n34128), .Z(n34085) );
  XNOR U35207 ( .A(n34131), .B(n34085), .Z(N745) );
  AND U35208 ( .A(x[488]), .B(y[8040]), .Z(n34086) );
  NAND U35209 ( .A(n34086), .B(n34561), .Z(n34090) );
  NAND U35210 ( .A(n34088), .B(n34087), .Z(n34089) );
  AND U35211 ( .A(n34090), .B(n34089), .Z(n34171) );
  AND U35212 ( .A(o[360]), .B(n34091), .Z(n34144) );
  AND U35213 ( .A(y[8036]), .B(x[485]), .Z(n34093) );
  NAND U35214 ( .A(y[8034]), .B(x[487]), .Z(n34092) );
  XNOR U35215 ( .A(n34093), .B(n34092), .Z(n34143) );
  XNOR U35216 ( .A(n34144), .B(n34143), .Z(n34169) );
  AND U35217 ( .A(y[8032]), .B(x[489]), .Z(n34095) );
  NAND U35218 ( .A(y[8041]), .B(x[480]), .Z(n34094) );
  XNOR U35219 ( .A(n34095), .B(n34094), .Z(n34151) );
  AND U35220 ( .A(x[488]), .B(y[8033]), .Z(n34158) );
  XOR U35221 ( .A(o[361]), .B(n34158), .Z(n34150) );
  XNOR U35222 ( .A(n34151), .B(n34150), .Z(n34168) );
  XOR U35223 ( .A(n34169), .B(n34168), .Z(n34170) );
  XNOR U35224 ( .A(n34171), .B(n34170), .Z(n34165) );
  AND U35225 ( .A(y[8035]), .B(x[486]), .Z(n34509) );
  NAND U35226 ( .A(y[8040]), .B(x[481]), .Z(n34096) );
  XNOR U35227 ( .A(n34509), .B(n34096), .Z(n34155) );
  XNOR U35228 ( .A(n34566), .B(n34155), .Z(n34175) );
  AND U35229 ( .A(x[482]), .B(y[8039]), .Z(n34810) );
  NAND U35230 ( .A(x[483]), .B(y[8038]), .Z(n34517) );
  XNOR U35231 ( .A(n34810), .B(n34517), .Z(n34174) );
  XNOR U35232 ( .A(n34175), .B(n34174), .Z(n34163) );
  NAND U35233 ( .A(x[485]), .B(y[8039]), .Z(n34360) );
  AND U35234 ( .A(x[481]), .B(y[8035]), .Z(n34154) );
  NANDN U35235 ( .A(n34360), .B(n34154), .Z(n34100) );
  NAND U35236 ( .A(n34098), .B(n34097), .Z(n34099) );
  NAND U35237 ( .A(n34100), .B(n34099), .Z(n34162) );
  XOR U35238 ( .A(n34163), .B(n34162), .Z(n34164) );
  XNOR U35239 ( .A(n34165), .B(n34164), .Z(n34138) );
  NANDN U35240 ( .A(n34101), .B(n34897), .Z(n34105) );
  NANDN U35241 ( .A(n34103), .B(n34102), .Z(n34104) );
  NAND U35242 ( .A(n34105), .B(n34104), .Z(n34136) );
  NAND U35243 ( .A(n34280), .B(n34106), .Z(n34109) );
  NAND U35244 ( .A(n34763), .B(n34107), .Z(n34108) );
  AND U35245 ( .A(n34109), .B(n34108), .Z(n34137) );
  XNOR U35246 ( .A(n34136), .B(n34137), .Z(n34139) );
  NAND U35247 ( .A(n34111), .B(n34110), .Z(n34115) );
  NAND U35248 ( .A(n34113), .B(n34112), .Z(n34114) );
  NAND U35249 ( .A(n34115), .B(n34114), .Z(n34179) );
  NAND U35250 ( .A(n34117), .B(n34116), .Z(n34121) );
  NAND U35251 ( .A(n34119), .B(n34118), .Z(n34120) );
  NAND U35252 ( .A(n34121), .B(n34120), .Z(n34178) );
  XOR U35253 ( .A(n34179), .B(n34178), .Z(n34181) );
  XOR U35254 ( .A(n34180), .B(n34181), .Z(n34186) );
  NAND U35255 ( .A(n34123), .B(n34122), .Z(n34127) );
  NANDN U35256 ( .A(n34125), .B(n34124), .Z(n34126) );
  NAND U35257 ( .A(n34127), .B(n34126), .Z(n34184) );
  NANDN U35258 ( .A(n34128), .B(n34129), .Z(n34134) );
  NOR U35259 ( .A(n34130), .B(n34129), .Z(n34132) );
  OR U35260 ( .A(n34132), .B(n34131), .Z(n34133) );
  AND U35261 ( .A(n34134), .B(n34133), .Z(n34185) );
  XOR U35262 ( .A(n34184), .B(n34185), .Z(n34135) );
  XNOR U35263 ( .A(n34186), .B(n34135), .Z(N746) );
  NAND U35264 ( .A(n34137), .B(n34136), .Z(n34141) );
  NANDN U35265 ( .A(n34139), .B(n34138), .Z(n34140) );
  NAND U35266 ( .A(n34141), .B(n34140), .Z(n34245) );
  AND U35267 ( .A(x[487]), .B(y[8036]), .Z(n34224) );
  NAND U35268 ( .A(n34224), .B(n34142), .Z(n34146) );
  NAND U35269 ( .A(n34144), .B(n34143), .Z(n34145) );
  AND U35270 ( .A(n34146), .B(n34145), .Z(n34237) );
  AND U35271 ( .A(y[8035]), .B(x[487]), .Z(n34148) );
  NAND U35272 ( .A(y[8038]), .B(x[484]), .Z(n34147) );
  XNOR U35273 ( .A(n34148), .B(n34147), .Z(n34208) );
  AND U35274 ( .A(x[486]), .B(y[8036]), .Z(n34207) );
  XNOR U35275 ( .A(n34208), .B(n34207), .Z(n34235) );
  AND U35276 ( .A(x[488]), .B(y[8034]), .Z(n34420) );
  AND U35277 ( .A(x[489]), .B(y[8033]), .Z(n34218) );
  XOR U35278 ( .A(o[362]), .B(n34218), .Z(n34229) );
  XOR U35279 ( .A(n34420), .B(n34229), .Z(n34230) );
  XNOR U35280 ( .A(n34231), .B(n34230), .Z(n34234) );
  XOR U35281 ( .A(n34235), .B(n34234), .Z(n34236) );
  XNOR U35282 ( .A(n34237), .B(n34236), .Z(n34197) );
  AND U35283 ( .A(x[489]), .B(y[8041]), .Z(n34149) );
  NAND U35284 ( .A(n34149), .B(n34561), .Z(n34153) );
  NAND U35285 ( .A(n34151), .B(n34150), .Z(n34152) );
  NAND U35286 ( .A(n34153), .B(n34152), .Z(n34195) );
  AND U35287 ( .A(x[486]), .B(y[8040]), .Z(n34454) );
  NAND U35288 ( .A(n34454), .B(n34154), .Z(n34157) );
  NAND U35289 ( .A(n34566), .B(n34155), .Z(n34156) );
  NAND U35290 ( .A(n34157), .B(n34156), .Z(n34203) );
  AND U35291 ( .A(o[361]), .B(n34158), .Z(n34213) );
  AND U35292 ( .A(y[8032]), .B(x[490]), .Z(n34160) );
  AND U35293 ( .A(y[8042]), .B(x[480]), .Z(n34159) );
  XOR U35294 ( .A(n34160), .B(n34159), .Z(n34212) );
  XOR U35295 ( .A(n34213), .B(n34212), .Z(n34201) );
  AND U35296 ( .A(y[8039]), .B(x[483]), .Z(n35129) );
  NAND U35297 ( .A(y[8041]), .B(x[481]), .Z(n34161) );
  XNOR U35298 ( .A(n35129), .B(n34161), .Z(n34225) );
  AND U35299 ( .A(x[482]), .B(y[8040]), .Z(n34226) );
  XOR U35300 ( .A(n34225), .B(n34226), .Z(n34200) );
  XOR U35301 ( .A(n34201), .B(n34200), .Z(n34202) );
  XOR U35302 ( .A(n34203), .B(n34202), .Z(n34194) );
  XOR U35303 ( .A(n34195), .B(n34194), .Z(n34196) );
  XOR U35304 ( .A(n34197), .B(n34196), .Z(n34244) );
  NAND U35305 ( .A(n34163), .B(n34162), .Z(n34167) );
  NAND U35306 ( .A(n34165), .B(n34164), .Z(n34166) );
  AND U35307 ( .A(n34167), .B(n34166), .Z(n34191) );
  NAND U35308 ( .A(n34169), .B(n34168), .Z(n34173) );
  NAND U35309 ( .A(n34171), .B(n34170), .Z(n34172) );
  AND U35310 ( .A(n34173), .B(n34172), .Z(n34188) );
  NAND U35311 ( .A(n34175), .B(n34174), .Z(n34177) );
  ANDN U35312 ( .B(n34517), .A(n34810), .Z(n34176) );
  ANDN U35313 ( .B(n34177), .A(n34176), .Z(n34189) );
  XOR U35314 ( .A(n34188), .B(n34189), .Z(n34190) );
  XOR U35315 ( .A(n34191), .B(n34190), .Z(n34243) );
  XOR U35316 ( .A(n34245), .B(n34246), .Z(n34242) );
  NAND U35317 ( .A(n34179), .B(n34178), .Z(n34183) );
  NAND U35318 ( .A(n34181), .B(n34180), .Z(n34182) );
  NAND U35319 ( .A(n34183), .B(n34182), .Z(n34241) );
  XOR U35320 ( .A(n34241), .B(n34240), .Z(n34187) );
  XNOR U35321 ( .A(n34242), .B(n34187), .Z(N747) );
  NAND U35322 ( .A(n34189), .B(n34188), .Z(n34193) );
  NANDN U35323 ( .A(n34191), .B(n34190), .Z(n34192) );
  AND U35324 ( .A(n34193), .B(n34192), .Z(n34315) );
  NAND U35325 ( .A(n34195), .B(n34194), .Z(n34199) );
  NAND U35326 ( .A(n34197), .B(n34196), .Z(n34198) );
  NAND U35327 ( .A(n34199), .B(n34198), .Z(n34313) );
  NAND U35328 ( .A(n34201), .B(n34200), .Z(n34205) );
  NAND U35329 ( .A(n34203), .B(n34202), .Z(n34204) );
  NAND U35330 ( .A(n34205), .B(n34204), .Z(n34301) );
  AND U35331 ( .A(x[487]), .B(y[8038]), .Z(n34355) );
  AND U35332 ( .A(x[484]), .B(y[8035]), .Z(n34206) );
  NAND U35333 ( .A(n34355), .B(n34206), .Z(n34210) );
  NAND U35334 ( .A(n34208), .B(n34207), .Z(n34209) );
  NAND U35335 ( .A(n34210), .B(n34209), .Z(n34299) );
  AND U35336 ( .A(x[490]), .B(y[8042]), .Z(n34211) );
  NAND U35337 ( .A(n34211), .B(n34561), .Z(n34215) );
  NAND U35338 ( .A(n34213), .B(n34212), .Z(n34214) );
  NAND U35339 ( .A(n34215), .B(n34214), .Z(n34295) );
  AND U35340 ( .A(y[8032]), .B(x[491]), .Z(n34217) );
  NAND U35341 ( .A(y[8043]), .B(x[480]), .Z(n34216) );
  XNOR U35342 ( .A(n34217), .B(n34216), .Z(n34271) );
  AND U35343 ( .A(o[362]), .B(n34218), .Z(n34270) );
  XOR U35344 ( .A(n34271), .B(n34270), .Z(n34294) );
  AND U35345 ( .A(y[8037]), .B(x[486]), .Z(n34220) );
  NAND U35346 ( .A(y[8042]), .B(x[481]), .Z(n34219) );
  XNOR U35347 ( .A(n34220), .B(n34219), .Z(n34262) );
  AND U35348 ( .A(x[490]), .B(y[8033]), .Z(n34281) );
  XOR U35349 ( .A(o[363]), .B(n34281), .Z(n34261) );
  XOR U35350 ( .A(n34262), .B(n34261), .Z(n34293) );
  XOR U35351 ( .A(n34294), .B(n34293), .Z(n34296) );
  XNOR U35352 ( .A(n34295), .B(n34296), .Z(n34300) );
  XOR U35353 ( .A(n34301), .B(n34302), .Z(n34284) );
  AND U35354 ( .A(x[483]), .B(y[8040]), .Z(n35262) );
  NAND U35355 ( .A(y[8041]), .B(x[482]), .Z(n34221) );
  XNOR U35356 ( .A(n34222), .B(n34221), .Z(n34257) );
  AND U35357 ( .A(x[484]), .B(y[8039]), .Z(n34256) );
  XNOR U35358 ( .A(n34257), .B(n34256), .Z(n34288) );
  XNOR U35359 ( .A(n35262), .B(n34288), .Z(n34290) );
  NAND U35360 ( .A(y[8034]), .B(x[489]), .Z(n34223) );
  XNOR U35361 ( .A(n34224), .B(n34223), .Z(n34276) );
  AND U35362 ( .A(x[488]), .B(y[8035]), .Z(n34275) );
  XNOR U35363 ( .A(n34276), .B(n34275), .Z(n34289) );
  XNOR U35364 ( .A(n34290), .B(n34289), .Z(n34253) );
  NAND U35365 ( .A(x[483]), .B(y[8041]), .Z(n34351) );
  AND U35366 ( .A(x[481]), .B(y[8039]), .Z(n34556) );
  NANDN U35367 ( .A(n34351), .B(n34556), .Z(n34228) );
  NAND U35368 ( .A(n34226), .B(n34225), .Z(n34227) );
  NAND U35369 ( .A(n34228), .B(n34227), .Z(n34251) );
  NAND U35370 ( .A(n34420), .B(n34229), .Z(n34233) );
  NAND U35371 ( .A(n34231), .B(n34230), .Z(n34232) );
  NAND U35372 ( .A(n34233), .B(n34232), .Z(n34250) );
  XOR U35373 ( .A(n34251), .B(n34250), .Z(n34252) );
  XNOR U35374 ( .A(n34253), .B(n34252), .Z(n34283) );
  NAND U35375 ( .A(n34235), .B(n34234), .Z(n34239) );
  NAND U35376 ( .A(n34237), .B(n34236), .Z(n34238) );
  NAND U35377 ( .A(n34239), .B(n34238), .Z(n34282) );
  XOR U35378 ( .A(n34283), .B(n34282), .Z(n34285) );
  XNOR U35379 ( .A(n34284), .B(n34285), .Z(n34312) );
  XOR U35380 ( .A(n34313), .B(n34312), .Z(n34314) );
  XOR U35381 ( .A(n34315), .B(n34314), .Z(n34308) );
  NANDN U35382 ( .A(n34244), .B(n34243), .Z(n34248) );
  NAND U35383 ( .A(n34246), .B(n34245), .Z(n34247) );
  AND U35384 ( .A(n34248), .B(n34247), .Z(n34306) );
  IV U35385 ( .A(n34306), .Z(n34305) );
  XOR U35386 ( .A(n34307), .B(n34305), .Z(n34249) );
  XNOR U35387 ( .A(n34308), .B(n34249), .Z(N748) );
  NAND U35388 ( .A(n34251), .B(n34250), .Z(n34255) );
  NAND U35389 ( .A(n34253), .B(n34252), .Z(n34254) );
  NAND U35390 ( .A(n34255), .B(n34254), .Z(n34391) );
  AND U35391 ( .A(x[485]), .B(y[8041]), .Z(n34801) );
  NAND U35392 ( .A(n34978), .B(n34801), .Z(n34259) );
  NAND U35393 ( .A(n34257), .B(n34256), .Z(n34258) );
  NAND U35394 ( .A(n34259), .B(n34258), .Z(n34339) );
  AND U35395 ( .A(x[486]), .B(y[8042]), .Z(n34573) );
  NAND U35396 ( .A(n34573), .B(n34260), .Z(n34264) );
  NAND U35397 ( .A(n34262), .B(n34261), .Z(n34263) );
  NAND U35398 ( .A(n34264), .B(n34263), .Z(n34338) );
  XOR U35399 ( .A(n34339), .B(n34338), .Z(n34341) );
  AND U35400 ( .A(x[489]), .B(y[8035]), .Z(n34973) );
  AND U35401 ( .A(y[8034]), .B(x[490]), .Z(n35027) );
  NAND U35402 ( .A(y[8040]), .B(x[484]), .Z(n34265) );
  XNOR U35403 ( .A(n35027), .B(n34265), .Z(n34382) );
  XOR U35404 ( .A(n34973), .B(n34382), .Z(n34361) );
  NAND U35405 ( .A(x[487]), .B(y[8037]), .Z(n34359) );
  XOR U35406 ( .A(n34360), .B(n34359), .Z(n34362) );
  AND U35407 ( .A(y[8032]), .B(x[492]), .Z(n34267) );
  NAND U35408 ( .A(y[8044]), .B(x[480]), .Z(n34266) );
  XNOR U35409 ( .A(n34267), .B(n34266), .Z(n34375) );
  NAND U35410 ( .A(x[491]), .B(y[8033]), .Z(n34356) );
  XNOR U35411 ( .A(o[364]), .B(n34356), .Z(n34376) );
  XOR U35412 ( .A(n34375), .B(n34376), .Z(n34345) );
  AND U35413 ( .A(y[8042]), .B(x[482]), .Z(n34269) );
  NAND U35414 ( .A(y[8036]), .B(x[488]), .Z(n34268) );
  XNOR U35415 ( .A(n34269), .B(n34268), .Z(n34350) );
  XOR U35416 ( .A(n34345), .B(n34344), .Z(n34347) );
  XOR U35417 ( .A(n34346), .B(n34347), .Z(n34340) );
  XOR U35418 ( .A(n34341), .B(n34340), .Z(n34390) );
  AND U35419 ( .A(x[491]), .B(y[8043]), .Z(n35381) );
  NAND U35420 ( .A(n35381), .B(n34561), .Z(n34273) );
  NAND U35421 ( .A(n34271), .B(n34270), .Z(n34272) );
  NAND U35422 ( .A(n34273), .B(n34272), .Z(n34368) );
  AND U35423 ( .A(x[487]), .B(y[8034]), .Z(n34495) );
  AND U35424 ( .A(x[489]), .B(y[8036]), .Z(n34274) );
  NAND U35425 ( .A(n34495), .B(n34274), .Z(n34278) );
  NAND U35426 ( .A(n34276), .B(n34275), .Z(n34277) );
  NAND U35427 ( .A(n34278), .B(n34277), .Z(n34366) );
  NAND U35428 ( .A(y[8043]), .B(x[481]), .Z(n34279) );
  XNOR U35429 ( .A(n34280), .B(n34279), .Z(n34372) );
  AND U35430 ( .A(o[363]), .B(n34281), .Z(n34371) );
  XOR U35431 ( .A(n34372), .B(n34371), .Z(n34365) );
  XOR U35432 ( .A(n34366), .B(n34365), .Z(n34367) );
  XOR U35433 ( .A(n34368), .B(n34367), .Z(n34389) );
  XOR U35434 ( .A(n34390), .B(n34389), .Z(n34392) );
  XNOR U35435 ( .A(n34391), .B(n34392), .Z(n34320) );
  NAND U35436 ( .A(n34283), .B(n34282), .Z(n34287) );
  NAND U35437 ( .A(n34285), .B(n34284), .Z(n34286) );
  NAND U35438 ( .A(n34287), .B(n34286), .Z(n34319) );
  XOR U35439 ( .A(n34320), .B(n34319), .Z(n34322) );
  NANDN U35440 ( .A(n35262), .B(n34288), .Z(n34292) );
  NAND U35441 ( .A(n34290), .B(n34289), .Z(n34291) );
  NAND U35442 ( .A(n34292), .B(n34291), .Z(n34332) );
  NAND U35443 ( .A(n34294), .B(n34293), .Z(n34298) );
  NAND U35444 ( .A(n34296), .B(n34295), .Z(n34297) );
  AND U35445 ( .A(n34298), .B(n34297), .Z(n34333) );
  XOR U35446 ( .A(n34332), .B(n34333), .Z(n34335) );
  NANDN U35447 ( .A(n34300), .B(n34299), .Z(n34304) );
  NANDN U35448 ( .A(n34302), .B(n34301), .Z(n34303) );
  AND U35449 ( .A(n34304), .B(n34303), .Z(n34334) );
  XOR U35450 ( .A(n34335), .B(n34334), .Z(n34321) );
  XNOR U35451 ( .A(n34322), .B(n34321), .Z(n34328) );
  OR U35452 ( .A(n34307), .B(n34305), .Z(n34311) );
  ANDN U35453 ( .B(n34307), .A(n34306), .Z(n34309) );
  OR U35454 ( .A(n34309), .B(n34308), .Z(n34310) );
  AND U35455 ( .A(n34311), .B(n34310), .Z(n34326) );
  NAND U35456 ( .A(n34313), .B(n34312), .Z(n34317) );
  NANDN U35457 ( .A(n34315), .B(n34314), .Z(n34316) );
  AND U35458 ( .A(n34317), .B(n34316), .Z(n34327) );
  IV U35459 ( .A(n34327), .Z(n34325) );
  XOR U35460 ( .A(n34326), .B(n34325), .Z(n34318) );
  XNOR U35461 ( .A(n34328), .B(n34318), .Z(N749) );
  NAND U35462 ( .A(n34320), .B(n34319), .Z(n34324) );
  NAND U35463 ( .A(n34322), .B(n34321), .Z(n34323) );
  AND U35464 ( .A(n34324), .B(n34323), .Z(n34462) );
  NANDN U35465 ( .A(n34325), .B(n34326), .Z(n34331) );
  NOR U35466 ( .A(n34327), .B(n34326), .Z(n34329) );
  OR U35467 ( .A(n34329), .B(n34328), .Z(n34330) );
  AND U35468 ( .A(n34331), .B(n34330), .Z(n34461) );
  NAND U35469 ( .A(n34333), .B(n34332), .Z(n34337) );
  NAND U35470 ( .A(n34335), .B(n34334), .Z(n34336) );
  NAND U35471 ( .A(n34337), .B(n34336), .Z(n34466) );
  NAND U35472 ( .A(n34339), .B(n34338), .Z(n34343) );
  NAND U35473 ( .A(n34341), .B(n34340), .Z(n34342) );
  NAND U35474 ( .A(n34343), .B(n34342), .Z(n34397) );
  NAND U35475 ( .A(n34345), .B(n34344), .Z(n34349) );
  NAND U35476 ( .A(n34347), .B(n34346), .Z(n34348) );
  NAND U35477 ( .A(n34349), .B(n34348), .Z(n34404) );
  AND U35478 ( .A(y[8042]), .B(x[488]), .Z(n35678) );
  AND U35479 ( .A(x[482]), .B(y[8036]), .Z(n34505) );
  NAND U35480 ( .A(n35678), .B(n34505), .Z(n34353) );
  NANDN U35481 ( .A(n34351), .B(n34350), .Z(n34352) );
  NAND U35482 ( .A(n34353), .B(n34352), .Z(n34433) );
  NAND U35483 ( .A(y[8044]), .B(x[481]), .Z(n34354) );
  XNOR U35484 ( .A(n34355), .B(n34354), .Z(n34426) );
  ANDN U35485 ( .B(o[364]), .A(n34356), .Z(n34425) );
  XOR U35486 ( .A(n34426), .B(n34425), .Z(n34430) );
  AND U35487 ( .A(x[486]), .B(y[8039]), .Z(n35421) );
  AND U35488 ( .A(y[8043]), .B(x[482]), .Z(n34358) );
  NAND U35489 ( .A(y[8036]), .B(x[489]), .Z(n34357) );
  XOR U35490 ( .A(n34358), .B(n34357), .Z(n34437) );
  XNOR U35491 ( .A(n35421), .B(n34437), .Z(n34431) );
  XOR U35492 ( .A(n34430), .B(n34431), .Z(n34432) );
  XOR U35493 ( .A(n34433), .B(n34432), .Z(n34403) );
  NAND U35494 ( .A(n34360), .B(n34359), .Z(n34364) );
  ANDN U35495 ( .B(n34362), .A(n34361), .Z(n34363) );
  ANDN U35496 ( .B(n34364), .A(n34363), .Z(n34402) );
  XOR U35497 ( .A(n34403), .B(n34402), .Z(n34405) );
  XOR U35498 ( .A(n34404), .B(n34405), .Z(n34396) );
  XOR U35499 ( .A(n34397), .B(n34396), .Z(n34399) );
  NAND U35500 ( .A(n34366), .B(n34365), .Z(n34370) );
  NAND U35501 ( .A(n34368), .B(n34367), .Z(n34369) );
  NAND U35502 ( .A(n34370), .B(n34369), .Z(n34411) );
  AND U35503 ( .A(x[486]), .B(y[8043]), .Z(n34802) );
  AND U35504 ( .A(x[481]), .B(y[8038]), .Z(n34424) );
  NAND U35505 ( .A(n34802), .B(n34424), .Z(n34374) );
  NAND U35506 ( .A(n34372), .B(n34371), .Z(n34373) );
  NAND U35507 ( .A(n34374), .B(n34373), .Z(n34417) );
  AND U35508 ( .A(x[492]), .B(y[8044]), .Z(n35684) );
  NAND U35509 ( .A(n35684), .B(n34561), .Z(n34378) );
  NAND U35510 ( .A(n34376), .B(n34375), .Z(n34377) );
  NAND U35511 ( .A(n34378), .B(n34377), .Z(n34415) );
  AND U35512 ( .A(x[490]), .B(y[8035]), .Z(n35274) );
  AND U35513 ( .A(y[8034]), .B(x[491]), .Z(n35223) );
  NAND U35514 ( .A(y[8037]), .B(x[488]), .Z(n34379) );
  XOR U35515 ( .A(n35223), .B(n34379), .Z(n34421) );
  XNOR U35516 ( .A(n35274), .B(n34421), .Z(n34414) );
  XOR U35517 ( .A(n34415), .B(n34414), .Z(n34416) );
  XOR U35518 ( .A(n34417), .B(n34416), .Z(n34409) );
  AND U35519 ( .A(x[490]), .B(y[8040]), .Z(n34381) );
  AND U35520 ( .A(x[484]), .B(y[8034]), .Z(n34380) );
  NAND U35521 ( .A(n34381), .B(n34380), .Z(n34384) );
  NAND U35522 ( .A(n34382), .B(n34973), .Z(n34383) );
  NAND U35523 ( .A(n34384), .B(n34383), .Z(n34458) );
  AND U35524 ( .A(y[8032]), .B(x[493]), .Z(n34386) );
  NAND U35525 ( .A(y[8045]), .B(x[480]), .Z(n34385) );
  XNOR U35526 ( .A(n34386), .B(n34385), .Z(n34449) );
  NAND U35527 ( .A(x[492]), .B(y[8033]), .Z(n34442) );
  XOR U35528 ( .A(o[365]), .B(n34442), .Z(n34450) );
  XNOR U35529 ( .A(n34449), .B(n34450), .Z(n34455) );
  AND U35530 ( .A(y[8040]), .B(x[485]), .Z(n34388) );
  NAND U35531 ( .A(y[8042]), .B(x[483]), .Z(n34387) );
  XNOR U35532 ( .A(n34388), .B(n34387), .Z(n34445) );
  NAND U35533 ( .A(x[484]), .B(y[8041]), .Z(n34446) );
  XNOR U35534 ( .A(n34445), .B(n34446), .Z(n34456) );
  XOR U35535 ( .A(n34455), .B(n34456), .Z(n34457) );
  XOR U35536 ( .A(n34458), .B(n34457), .Z(n34408) );
  XOR U35537 ( .A(n34409), .B(n34408), .Z(n34410) );
  XOR U35538 ( .A(n34411), .B(n34410), .Z(n34398) );
  XOR U35539 ( .A(n34399), .B(n34398), .Z(n34465) );
  NAND U35540 ( .A(n34390), .B(n34389), .Z(n34394) );
  NAND U35541 ( .A(n34392), .B(n34391), .Z(n34393) );
  AND U35542 ( .A(n34394), .B(n34393), .Z(n34464) );
  XOR U35543 ( .A(n34466), .B(n34467), .Z(n34463) );
  XNOR U35544 ( .A(n34461), .B(n34463), .Z(n34395) );
  XOR U35545 ( .A(n34462), .B(n34395), .Z(N750) );
  NAND U35546 ( .A(n34397), .B(n34396), .Z(n34401) );
  NAND U35547 ( .A(n34399), .B(n34398), .Z(n34400) );
  NAND U35548 ( .A(n34401), .B(n34400), .Z(n34550) );
  NAND U35549 ( .A(n34403), .B(n34402), .Z(n34407) );
  NAND U35550 ( .A(n34405), .B(n34404), .Z(n34406) );
  NAND U35551 ( .A(n34407), .B(n34406), .Z(n34549) );
  XOR U35552 ( .A(n34550), .B(n34549), .Z(n34552) );
  NAND U35553 ( .A(n34409), .B(n34408), .Z(n34413) );
  NAND U35554 ( .A(n34411), .B(n34410), .Z(n34412) );
  NAND U35555 ( .A(n34413), .B(n34412), .Z(n34474) );
  NAND U35556 ( .A(n34415), .B(n34414), .Z(n34419) );
  NAND U35557 ( .A(n34417), .B(n34416), .Z(n34418) );
  AND U35558 ( .A(n34419), .B(n34418), .Z(n34480) );
  AND U35559 ( .A(x[491]), .B(y[8037]), .Z(n34587) );
  NAND U35560 ( .A(n34587), .B(n34420), .Z(n34423) );
  NANDN U35561 ( .A(n34421), .B(n35274), .Z(n34422) );
  AND U35562 ( .A(n34423), .B(n34422), .Z(n34531) );
  NAND U35563 ( .A(x[487]), .B(y[8044]), .Z(n34988) );
  XNOR U35564 ( .A(n34531), .B(n34530), .Z(n34533) );
  AND U35565 ( .A(x[484]), .B(y[8042]), .Z(n34906) );
  AND U35566 ( .A(y[8043]), .B(x[483]), .Z(n34428) );
  NAND U35567 ( .A(y[8038]), .B(x[488]), .Z(n34427) );
  XOR U35568 ( .A(n34428), .B(n34427), .Z(n34518) );
  XOR U35569 ( .A(n34801), .B(n34518), .Z(n34527) );
  XNOR U35570 ( .A(n34906), .B(n34527), .Z(n34529) );
  AND U35571 ( .A(x[489]), .B(y[8037]), .Z(n35094) );
  AND U35572 ( .A(y[8044]), .B(x[482]), .Z(n34429) );
  AND U35573 ( .A(y[8036]), .B(x[490]), .Z(n35124) );
  XOR U35574 ( .A(n34429), .B(n35124), .Z(n34506) );
  XOR U35575 ( .A(n35094), .B(n34506), .Z(n34528) );
  XOR U35576 ( .A(n34529), .B(n34528), .Z(n34532) );
  XNOR U35577 ( .A(n34533), .B(n34532), .Z(n34478) );
  NAND U35578 ( .A(n34431), .B(n34430), .Z(n34435) );
  NAND U35579 ( .A(n34433), .B(n34432), .Z(n34434) );
  AND U35580 ( .A(n34435), .B(n34434), .Z(n34477) );
  XOR U35581 ( .A(n34478), .B(n34477), .Z(n34479) );
  XNOR U35582 ( .A(n34480), .B(n34479), .Z(n34472) );
  AND U35583 ( .A(x[489]), .B(y[8043]), .Z(n34436) );
  NAND U35584 ( .A(n34436), .B(n34505), .Z(n34439) );
  NANDN U35585 ( .A(n34437), .B(n35421), .Z(n34438) );
  AND U35586 ( .A(n34439), .B(n34438), .Z(n34491) );
  AND U35587 ( .A(y[8032]), .B(x[494]), .Z(n34441) );
  NAND U35588 ( .A(y[8046]), .B(x[480]), .Z(n34440) );
  XNOR U35589 ( .A(n34441), .B(n34440), .Z(n34515) );
  ANDN U35590 ( .B(o[365]), .A(n34442), .Z(n34514) );
  XOR U35591 ( .A(n34515), .B(n34514), .Z(n34489) );
  NAND U35592 ( .A(y[8034]), .B(x[492]), .Z(n34443) );
  XNOR U35593 ( .A(n34444), .B(n34443), .Z(n34496) );
  NAND U35594 ( .A(x[493]), .B(y[8033]), .Z(n34504) );
  XOR U35595 ( .A(o[366]), .B(n34504), .Z(n34497) );
  XOR U35596 ( .A(n34496), .B(n34497), .Z(n34490) );
  XOR U35597 ( .A(n34489), .B(n34490), .Z(n34492) );
  XNOR U35598 ( .A(n34491), .B(n34492), .Z(n34537) );
  AND U35599 ( .A(x[485]), .B(y[8042]), .Z(n34574) );
  NAND U35600 ( .A(n35262), .B(n34574), .Z(n34448) );
  NANDN U35601 ( .A(n34446), .B(n34445), .Z(n34447) );
  AND U35602 ( .A(n34448), .B(n34447), .Z(n34485) );
  AND U35603 ( .A(x[493]), .B(y[8045]), .Z(n35925) );
  NAND U35604 ( .A(n35925), .B(n34561), .Z(n34452) );
  NANDN U35605 ( .A(n34450), .B(n34449), .Z(n34451) );
  AND U35606 ( .A(n34452), .B(n34451), .Z(n34484) );
  NAND U35607 ( .A(y[8035]), .B(x[491]), .Z(n34453) );
  XNOR U35608 ( .A(n34454), .B(n34453), .Z(n34510) );
  NAND U35609 ( .A(x[481]), .B(y[8045]), .Z(n34511) );
  XNOR U35610 ( .A(n34510), .B(n34511), .Z(n34483) );
  XOR U35611 ( .A(n34484), .B(n34483), .Z(n34486) );
  XNOR U35612 ( .A(n34485), .B(n34486), .Z(n34536) );
  XOR U35613 ( .A(n34537), .B(n34536), .Z(n34539) );
  NAND U35614 ( .A(n34456), .B(n34455), .Z(n34460) );
  NAND U35615 ( .A(n34458), .B(n34457), .Z(n34459) );
  AND U35616 ( .A(n34460), .B(n34459), .Z(n34538) );
  XNOR U35617 ( .A(n34539), .B(n34538), .Z(n34471) );
  XOR U35618 ( .A(n34472), .B(n34471), .Z(n34473) );
  XOR U35619 ( .A(n34474), .B(n34473), .Z(n34551) );
  XNOR U35620 ( .A(n34552), .B(n34551), .Z(n34545) );
  NANDN U35621 ( .A(n34465), .B(n34464), .Z(n34469) );
  NAND U35622 ( .A(n34467), .B(n34466), .Z(n34468) );
  AND U35623 ( .A(n34469), .B(n34468), .Z(n34543) );
  IV U35624 ( .A(n34543), .Z(n34542) );
  XOR U35625 ( .A(n34544), .B(n34542), .Z(n34470) );
  XNOR U35626 ( .A(n34545), .B(n34470), .Z(N751) );
  NAND U35627 ( .A(n34472), .B(n34471), .Z(n34476) );
  NAND U35628 ( .A(n34474), .B(n34473), .Z(n34475) );
  NAND U35629 ( .A(n34476), .B(n34475), .Z(n34641) );
  NAND U35630 ( .A(n34478), .B(n34477), .Z(n34482) );
  NAND U35631 ( .A(n34480), .B(n34479), .Z(n34481) );
  NAND U35632 ( .A(n34482), .B(n34481), .Z(n34616) );
  NANDN U35633 ( .A(n34484), .B(n34483), .Z(n34488) );
  OR U35634 ( .A(n34486), .B(n34485), .Z(n34487) );
  AND U35635 ( .A(n34488), .B(n34487), .Z(n34623) );
  NANDN U35636 ( .A(n34490), .B(n34489), .Z(n34494) );
  OR U35637 ( .A(n34492), .B(n34491), .Z(n34493) );
  AND U35638 ( .A(n34494), .B(n34493), .Z(n34621) );
  NAND U35639 ( .A(x[492]), .B(y[8039]), .Z(n34980) );
  NANDN U35640 ( .A(n34980), .B(n34495), .Z(n34499) );
  NANDN U35641 ( .A(n34497), .B(n34496), .Z(n34498) );
  AND U35642 ( .A(n34499), .B(n34498), .Z(n34597) );
  AND U35643 ( .A(y[8036]), .B(x[491]), .Z(n34501) );
  NAND U35644 ( .A(y[8034]), .B(x[493]), .Z(n34500) );
  XNOR U35645 ( .A(n34501), .B(n34500), .Z(n34601) );
  AND U35646 ( .A(x[492]), .B(y[8035]), .Z(n34600) );
  XOR U35647 ( .A(n34601), .B(n34600), .Z(n34595) );
  AND U35648 ( .A(y[8032]), .B(x[495]), .Z(n34503) );
  NAND U35649 ( .A(y[8047]), .B(x[480]), .Z(n34502) );
  XNOR U35650 ( .A(n34503), .B(n34502), .Z(n34563) );
  ANDN U35651 ( .B(o[366]), .A(n34504), .Z(n34562) );
  XNOR U35652 ( .A(n34563), .B(n34562), .Z(n34594) );
  XNOR U35653 ( .A(n34595), .B(n34594), .Z(n34596) );
  XOR U35654 ( .A(n34597), .B(n34596), .Z(n34629) );
  NAND U35655 ( .A(x[490]), .B(y[8044]), .Z(n35423) );
  NANDN U35656 ( .A(n35423), .B(n34505), .Z(n34508) );
  NAND U35657 ( .A(n35094), .B(n34506), .Z(n34507) );
  AND U35658 ( .A(n34508), .B(n34507), .Z(n34627) );
  AND U35659 ( .A(x[491]), .B(y[8040]), .Z(n34905) );
  NAND U35660 ( .A(n34905), .B(n34509), .Z(n34513) );
  NANDN U35661 ( .A(n34511), .B(n34510), .Z(n34512) );
  NAND U35662 ( .A(n34513), .B(n34512), .Z(n34626) );
  XNOR U35663 ( .A(n34627), .B(n34626), .Z(n34628) );
  XNOR U35664 ( .A(n34629), .B(n34628), .Z(n34620) );
  XNOR U35665 ( .A(n34621), .B(n34620), .Z(n34622) );
  XOR U35666 ( .A(n34623), .B(n34622), .Z(n34614) );
  AND U35667 ( .A(x[494]), .B(y[8046]), .Z(n36240) );
  AND U35668 ( .A(x[488]), .B(y[8043]), .Z(n34516) );
  NANDN U35669 ( .A(n34517), .B(n34516), .Z(n34520) );
  NANDN U35670 ( .A(n34518), .B(n34801), .Z(n34519) );
  NAND U35671 ( .A(n34520), .B(n34519), .Z(n34588) );
  XNOR U35672 ( .A(n34589), .B(n34588), .Z(n34591) );
  AND U35673 ( .A(y[8037]), .B(x[490]), .Z(n34522) );
  NAND U35674 ( .A(y[8043]), .B(x[484]), .Z(n34521) );
  XNOR U35675 ( .A(n34522), .B(n34521), .Z(n34569) );
  AND U35676 ( .A(x[487]), .B(y[8040]), .Z(n34568) );
  XOR U35677 ( .A(n34569), .B(n34568), .Z(n34576) );
  NAND U35678 ( .A(x[486]), .B(y[8041]), .Z(n34679) );
  XNOR U35679 ( .A(n34679), .B(n34574), .Z(n34575) );
  XOR U35680 ( .A(n34576), .B(n34575), .Z(n34610) );
  AND U35681 ( .A(y[8045]), .B(x[482]), .Z(n34524) );
  NAND U35682 ( .A(y[8038]), .B(x[489]), .Z(n34523) );
  XNOR U35683 ( .A(n34524), .B(n34523), .Z(n34579) );
  NAND U35684 ( .A(x[483]), .B(y[8044]), .Z(n34580) );
  XNOR U35685 ( .A(n34579), .B(n34580), .Z(n34608) );
  AND U35686 ( .A(y[8046]), .B(x[481]), .Z(n34526) );
  NAND U35687 ( .A(y[8039]), .B(x[488]), .Z(n34525) );
  XNOR U35688 ( .A(n34526), .B(n34525), .Z(n34557) );
  NAND U35689 ( .A(x[494]), .B(y[8033]), .Z(n34585) );
  XOR U35690 ( .A(o[367]), .B(n34585), .Z(n34558) );
  XOR U35691 ( .A(n34557), .B(n34558), .Z(n34609) );
  XOR U35692 ( .A(n34610), .B(n34611), .Z(n34590) );
  XOR U35693 ( .A(n34591), .B(n34590), .Z(n34633) );
  XNOR U35694 ( .A(n34633), .B(n34632), .Z(n34635) );
  NANDN U35695 ( .A(n34531), .B(n34530), .Z(n34535) );
  NAND U35696 ( .A(n34533), .B(n34532), .Z(n34534) );
  AND U35697 ( .A(n34535), .B(n34534), .Z(n34634) );
  XOR U35698 ( .A(n34635), .B(n34634), .Z(n34615) );
  XOR U35699 ( .A(n34614), .B(n34615), .Z(n34617) );
  XNOR U35700 ( .A(n34616), .B(n34617), .Z(n34638) );
  NAND U35701 ( .A(n34537), .B(n34536), .Z(n34541) );
  NAND U35702 ( .A(n34539), .B(n34538), .Z(n34540) );
  AND U35703 ( .A(n34541), .B(n34540), .Z(n34639) );
  XOR U35704 ( .A(n34638), .B(n34639), .Z(n34640) );
  XOR U35705 ( .A(n34641), .B(n34640), .Z(n34647) );
  OR U35706 ( .A(n34544), .B(n34542), .Z(n34548) );
  ANDN U35707 ( .B(n34544), .A(n34543), .Z(n34546) );
  OR U35708 ( .A(n34546), .B(n34545), .Z(n34547) );
  AND U35709 ( .A(n34548), .B(n34547), .Z(n34645) );
  NAND U35710 ( .A(n34550), .B(n34549), .Z(n34554) );
  NAND U35711 ( .A(n34552), .B(n34551), .Z(n34553) );
  AND U35712 ( .A(n34554), .B(n34553), .Z(n34646) );
  IV U35713 ( .A(n34646), .Z(n34644) );
  XOR U35714 ( .A(n34645), .B(n34644), .Z(n34555) );
  XNOR U35715 ( .A(n34647), .B(n34555), .Z(N752) );
  AND U35716 ( .A(x[488]), .B(y[8046]), .Z(n34907) );
  NAND U35717 ( .A(n34907), .B(n34556), .Z(n34560) );
  NANDN U35718 ( .A(n34558), .B(n34557), .Z(n34559) );
  NAND U35719 ( .A(n34560), .B(n34559), .Z(n34709) );
  AND U35720 ( .A(x[495]), .B(y[8047]), .Z(n36616) );
  NAND U35721 ( .A(n36616), .B(n34561), .Z(n34565) );
  NAND U35722 ( .A(n34563), .B(n34562), .Z(n34564) );
  NAND U35723 ( .A(n34565), .B(n34564), .Z(n34708) );
  XOR U35724 ( .A(n34709), .B(n34708), .Z(n34711) );
  AND U35725 ( .A(x[490]), .B(y[8043]), .Z(n34567) );
  NAND U35726 ( .A(n34567), .B(n34566), .Z(n34571) );
  NAND U35727 ( .A(n34569), .B(n34568), .Z(n34570) );
  NAND U35728 ( .A(n34571), .B(n34570), .Z(n34666) );
  AND U35729 ( .A(x[480]), .B(y[8048]), .Z(n34688) );
  AND U35730 ( .A(x[496]), .B(y[8032]), .Z(n34689) );
  XOR U35731 ( .A(n34688), .B(n34689), .Z(n34690) );
  NAND U35732 ( .A(x[495]), .B(y[8033]), .Z(n34676) );
  XNOR U35733 ( .A(o[368]), .B(n34676), .Z(n34691) );
  XOR U35734 ( .A(n34690), .B(n34691), .Z(n34665) );
  NAND U35735 ( .A(y[8041]), .B(x[487]), .Z(n34572) );
  XNOR U35736 ( .A(n34573), .B(n34572), .Z(n34681) );
  AND U35737 ( .A(x[490]), .B(y[8038]), .Z(n34680) );
  XOR U35738 ( .A(n34681), .B(n34680), .Z(n34664) );
  XOR U35739 ( .A(n34665), .B(n34664), .Z(n34667) );
  XOR U35740 ( .A(n34666), .B(n34667), .Z(n34710) );
  XOR U35741 ( .A(n34711), .B(n34710), .Z(n34661) );
  NANDN U35742 ( .A(n34574), .B(n34679), .Z(n34578) );
  NANDN U35743 ( .A(n34576), .B(n34575), .Z(n34577) );
  AND U35744 ( .A(n34578), .B(n34577), .Z(n34659) );
  NAND U35745 ( .A(x[489]), .B(y[8045]), .Z(n35393) );
  NANDN U35746 ( .A(n35393), .B(n34978), .Z(n34582) );
  NANDN U35747 ( .A(n34580), .B(n34579), .Z(n34581) );
  AND U35748 ( .A(n34582), .B(n34581), .Z(n34699) );
  AND U35749 ( .A(y[8047]), .B(x[481]), .Z(n34584) );
  NAND U35750 ( .A(y[8040]), .B(x[488]), .Z(n34583) );
  XNOR U35751 ( .A(n34584), .B(n34583), .Z(n34685) );
  ANDN U35752 ( .B(o[367]), .A(n34585), .Z(n34684) );
  XOR U35753 ( .A(n34685), .B(n34684), .Z(n34696) );
  NAND U35754 ( .A(y[8034]), .B(x[494]), .Z(n34586) );
  XNOR U35755 ( .A(n34587), .B(n34586), .Z(n34720) );
  NAND U35756 ( .A(x[484]), .B(y[8044]), .Z(n34721) );
  XOR U35757 ( .A(n34720), .B(n34721), .Z(n34697) );
  XOR U35758 ( .A(n34699), .B(n34698), .Z(n34658) );
  XNOR U35759 ( .A(n34659), .B(n34658), .Z(n34660) );
  XNOR U35760 ( .A(n34661), .B(n34660), .Z(n34702) );
  NANDN U35761 ( .A(n34589), .B(n34588), .Z(n34593) );
  NAND U35762 ( .A(n34591), .B(n34590), .Z(n34592) );
  NAND U35763 ( .A(n34593), .B(n34592), .Z(n34703) );
  XNOR U35764 ( .A(n34702), .B(n34703), .Z(n34704) );
  NANDN U35765 ( .A(n34595), .B(n34594), .Z(n34599) );
  NAND U35766 ( .A(n34597), .B(n34596), .Z(n34598) );
  AND U35767 ( .A(n34599), .B(n34598), .Z(n34734) );
  AND U35768 ( .A(x[493]), .B(y[8036]), .Z(n34730) );
  NAND U35769 ( .A(n35223), .B(n34730), .Z(n34603) );
  NAND U35770 ( .A(n34601), .B(n34600), .Z(n34602) );
  NAND U35771 ( .A(n34603), .B(n34602), .Z(n34717) );
  AND U35772 ( .A(y[8046]), .B(x[482]), .Z(n34605) );
  NAND U35773 ( .A(y[8039]), .B(x[489]), .Z(n34604) );
  XNOR U35774 ( .A(n34605), .B(n34604), .Z(n34724) );
  NAND U35775 ( .A(x[483]), .B(y[8045]), .Z(n34725) );
  XNOR U35776 ( .A(n34724), .B(n34725), .Z(n34714) );
  AND U35777 ( .A(x[492]), .B(y[8036]), .Z(n35398) );
  AND U35778 ( .A(y[8043]), .B(x[485]), .Z(n34607) );
  NAND U35779 ( .A(y[8035]), .B(x[493]), .Z(n34606) );
  XOR U35780 ( .A(n34607), .B(n34606), .Z(n34671) );
  XNOR U35781 ( .A(n35398), .B(n34671), .Z(n34715) );
  XOR U35782 ( .A(n34714), .B(n34715), .Z(n34716) );
  XNOR U35783 ( .A(n34717), .B(n34716), .Z(n34731) );
  NANDN U35784 ( .A(n34609), .B(n34608), .Z(n34613) );
  NAND U35785 ( .A(n34611), .B(n34610), .Z(n34612) );
  AND U35786 ( .A(n34613), .B(n34612), .Z(n34732) );
  XOR U35787 ( .A(n34731), .B(n34732), .Z(n34733) );
  XOR U35788 ( .A(n34704), .B(n34705), .Z(n34741) );
  NAND U35789 ( .A(n34615), .B(n34614), .Z(n34619) );
  NAND U35790 ( .A(n34617), .B(n34616), .Z(n34618) );
  AND U35791 ( .A(n34619), .B(n34618), .Z(n34740) );
  XOR U35792 ( .A(n34741), .B(n34740), .Z(n34743) );
  NANDN U35793 ( .A(n34621), .B(n34620), .Z(n34625) );
  NANDN U35794 ( .A(n34623), .B(n34622), .Z(n34624) );
  AND U35795 ( .A(n34625), .B(n34624), .Z(n34655) );
  NANDN U35796 ( .A(n34627), .B(n34626), .Z(n34631) );
  NANDN U35797 ( .A(n34629), .B(n34628), .Z(n34630) );
  AND U35798 ( .A(n34631), .B(n34630), .Z(n34653) );
  NANDN U35799 ( .A(n34633), .B(n34632), .Z(n34637) );
  NAND U35800 ( .A(n34635), .B(n34634), .Z(n34636) );
  AND U35801 ( .A(n34637), .B(n34636), .Z(n34652) );
  XNOR U35802 ( .A(n34653), .B(n34652), .Z(n34654) );
  XNOR U35803 ( .A(n34655), .B(n34654), .Z(n34742) );
  XNOR U35804 ( .A(n34743), .B(n34742), .Z(n34739) );
  NAND U35805 ( .A(n34639), .B(n34638), .Z(n34643) );
  NAND U35806 ( .A(n34641), .B(n34640), .Z(n34642) );
  NAND U35807 ( .A(n34643), .B(n34642), .Z(n34738) );
  NANDN U35808 ( .A(n34644), .B(n34645), .Z(n34650) );
  NOR U35809 ( .A(n34646), .B(n34645), .Z(n34648) );
  OR U35810 ( .A(n34648), .B(n34647), .Z(n34649) );
  AND U35811 ( .A(n34650), .B(n34649), .Z(n34737) );
  XOR U35812 ( .A(n34738), .B(n34737), .Z(n34651) );
  XNOR U35813 ( .A(n34739), .B(n34651), .Z(N753) );
  NANDN U35814 ( .A(n34653), .B(n34652), .Z(n34657) );
  NANDN U35815 ( .A(n34655), .B(n34654), .Z(n34656) );
  AND U35816 ( .A(n34657), .B(n34656), .Z(n34847) );
  NANDN U35817 ( .A(n34659), .B(n34658), .Z(n34663) );
  NANDN U35818 ( .A(n34661), .B(n34660), .Z(n34662) );
  AND U35819 ( .A(n34663), .B(n34662), .Z(n34756) );
  NAND U35820 ( .A(n34665), .B(n34664), .Z(n34669) );
  NAND U35821 ( .A(n34667), .B(n34666), .Z(n34668) );
  NAND U35822 ( .A(n34669), .B(n34668), .Z(n34838) );
  AND U35823 ( .A(x[493]), .B(y[8043]), .Z(n35692) );
  NAND U35824 ( .A(n35692), .B(n34670), .Z(n34673) );
  NANDN U35825 ( .A(n34671), .B(n35398), .Z(n34672) );
  NAND U35826 ( .A(n34673), .B(n34672), .Z(n34786) );
  AND U35827 ( .A(y[8048]), .B(x[481]), .Z(n34675) );
  NAND U35828 ( .A(y[8040]), .B(x[489]), .Z(n34674) );
  XNOR U35829 ( .A(n34675), .B(n34674), .Z(n34806) );
  NANDN U35830 ( .A(n34676), .B(o[368]), .Z(n34807) );
  XNOR U35831 ( .A(n34806), .B(n34807), .Z(n34784) );
  AND U35832 ( .A(y[8034]), .B(x[495]), .Z(n34678) );
  NAND U35833 ( .A(y[8037]), .B(x[492]), .Z(n34677) );
  XNOR U35834 ( .A(n34678), .B(n34677), .Z(n34759) );
  NAND U35835 ( .A(x[494]), .B(y[8035]), .Z(n34760) );
  XOR U35836 ( .A(n34784), .B(n34783), .Z(n34785) );
  XOR U35837 ( .A(n34786), .B(n34785), .Z(n34836) );
  AND U35838 ( .A(x[487]), .B(y[8042]), .Z(n34818) );
  NANDN U35839 ( .A(n34679), .B(n34818), .Z(n34683) );
  NAND U35840 ( .A(n34681), .B(n34680), .Z(n34682) );
  NAND U35841 ( .A(n34683), .B(n34682), .Z(n34796) );
  NAND U35842 ( .A(x[488]), .B(y[8047]), .Z(n35482) );
  AND U35843 ( .A(x[481]), .B(y[8040]), .Z(n34887) );
  NANDN U35844 ( .A(n35482), .B(n34887), .Z(n34687) );
  NAND U35845 ( .A(n34685), .B(n34684), .Z(n34686) );
  NAND U35846 ( .A(n34687), .B(n34686), .Z(n34795) );
  XOR U35847 ( .A(n34796), .B(n34795), .Z(n34798) );
  NAND U35848 ( .A(n34689), .B(n34688), .Z(n34693) );
  NAND U35849 ( .A(n34691), .B(n34690), .Z(n34692) );
  NAND U35850 ( .A(n34693), .B(n34692), .Z(n34792) );
  AND U35851 ( .A(x[480]), .B(y[8049]), .Z(n34773) );
  NAND U35852 ( .A(x[497]), .B(y[8032]), .Z(n34774) );
  NAND U35853 ( .A(x[496]), .B(y[8033]), .Z(n34770) );
  XOR U35854 ( .A(o[369]), .B(n34770), .Z(n34776) );
  AND U35855 ( .A(y[8047]), .B(x[482]), .Z(n34695) );
  NAND U35856 ( .A(y[8039]), .B(x[490]), .Z(n34694) );
  XNOR U35857 ( .A(n34695), .B(n34694), .Z(n34811) );
  NAND U35858 ( .A(x[483]), .B(y[8046]), .Z(n34812) );
  XNOR U35859 ( .A(n34811), .B(n34812), .Z(n34790) );
  XOR U35860 ( .A(n34789), .B(n34790), .Z(n34791) );
  XOR U35861 ( .A(n34792), .B(n34791), .Z(n34797) );
  XOR U35862 ( .A(n34798), .B(n34797), .Z(n34835) );
  XOR U35863 ( .A(n34836), .B(n34835), .Z(n34837) );
  XNOR U35864 ( .A(n34838), .B(n34837), .Z(n34753) );
  NANDN U35865 ( .A(n34697), .B(n34696), .Z(n34701) );
  NANDN U35866 ( .A(n34699), .B(n34698), .Z(n34700) );
  AND U35867 ( .A(n34701), .B(n34700), .Z(n34754) );
  XOR U35868 ( .A(n34753), .B(n34754), .Z(n34755) );
  NANDN U35869 ( .A(n34703), .B(n34702), .Z(n34707) );
  NANDN U35870 ( .A(n34705), .B(n34704), .Z(n34706) );
  AND U35871 ( .A(n34707), .B(n34706), .Z(n34750) );
  NAND U35872 ( .A(n34709), .B(n34708), .Z(n34713) );
  NAND U35873 ( .A(n34711), .B(n34710), .Z(n34712) );
  NAND U35874 ( .A(n34713), .B(n34712), .Z(n34832) );
  NAND U35875 ( .A(n34715), .B(n34714), .Z(n34719) );
  NAND U35876 ( .A(n34717), .B(n34716), .Z(n34718) );
  NAND U35877 ( .A(n34719), .B(n34718), .Z(n34830) );
  NAND U35878 ( .A(x[494]), .B(y[8037]), .Z(n35024) );
  NANDN U35879 ( .A(n35024), .B(n35223), .Z(n34723) );
  NANDN U35880 ( .A(n34721), .B(n34720), .Z(n34722) );
  AND U35881 ( .A(n34723), .B(n34722), .Z(n34824) );
  AND U35882 ( .A(x[489]), .B(y[8046]), .Z(n35673) );
  NAND U35883 ( .A(n34810), .B(n35673), .Z(n34727) );
  NANDN U35884 ( .A(n34725), .B(n34724), .Z(n34726) );
  NAND U35885 ( .A(n34727), .B(n34726), .Z(n34823) );
  XNOR U35886 ( .A(n34824), .B(n34823), .Z(n34825) );
  AND U35887 ( .A(x[485]), .B(y[8044]), .Z(n34869) );
  NAND U35888 ( .A(y[8041]), .B(x[488]), .Z(n34728) );
  XNOR U35889 ( .A(n34869), .B(n34728), .Z(n34803) );
  XOR U35890 ( .A(n34803), .B(n34802), .Z(n34817) );
  XOR U35891 ( .A(n34817), .B(n34818), .Z(n34819) );
  NAND U35892 ( .A(y[8045]), .B(x[484]), .Z(n34729) );
  XNOR U35893 ( .A(n34730), .B(n34729), .Z(n34764) );
  NAND U35894 ( .A(x[491]), .B(y[8038]), .Z(n34765) );
  XOR U35895 ( .A(n34764), .B(n34765), .Z(n34820) );
  XOR U35896 ( .A(n34819), .B(n34820), .Z(n34826) );
  XNOR U35897 ( .A(n34825), .B(n34826), .Z(n34829) );
  XOR U35898 ( .A(n34830), .B(n34829), .Z(n34831) );
  XNOR U35899 ( .A(n34832), .B(n34831), .Z(n34748) );
  NAND U35900 ( .A(n34732), .B(n34731), .Z(n34736) );
  NANDN U35901 ( .A(n34734), .B(n34733), .Z(n34735) );
  NAND U35902 ( .A(n34736), .B(n34735), .Z(n34747) );
  XOR U35903 ( .A(n34748), .B(n34747), .Z(n34749) );
  XOR U35904 ( .A(n34750), .B(n34749), .Z(n34844) );
  XOR U35905 ( .A(n34845), .B(n34844), .Z(n34846) );
  XOR U35906 ( .A(n34847), .B(n34846), .Z(n34843) );
  NAND U35907 ( .A(n34741), .B(n34740), .Z(n34745) );
  NAND U35908 ( .A(n34743), .B(n34742), .Z(n34744) );
  NAND U35909 ( .A(n34745), .B(n34744), .Z(n34841) );
  XNOR U35910 ( .A(n34842), .B(n34841), .Z(n34746) );
  XNOR U35911 ( .A(n34843), .B(n34746), .Z(N754) );
  NAND U35912 ( .A(n34748), .B(n34747), .Z(n34752) );
  NANDN U35913 ( .A(n34750), .B(n34749), .Z(n34751) );
  AND U35914 ( .A(n34752), .B(n34751), .Z(n34954) );
  NAND U35915 ( .A(n34754), .B(n34753), .Z(n34758) );
  NANDN U35916 ( .A(n34756), .B(n34755), .Z(n34757) );
  AND U35917 ( .A(n34758), .B(n34757), .Z(n34952) );
  AND U35918 ( .A(x[495]), .B(y[8037]), .Z(n34986) );
  AND U35919 ( .A(x[492]), .B(y[8034]), .Z(n35084) );
  NAND U35920 ( .A(n34986), .B(n35084), .Z(n34762) );
  NANDN U35921 ( .A(n34760), .B(n34759), .Z(n34761) );
  NAND U35922 ( .A(n34762), .B(n34761), .Z(n34934) );
  NAND U35923 ( .A(n35925), .B(n34763), .Z(n34767) );
  NANDN U35924 ( .A(n34765), .B(n34764), .Z(n34766) );
  AND U35925 ( .A(n34767), .B(n34766), .Z(n34924) );
  AND U35926 ( .A(y[8049]), .B(x[481]), .Z(n34769) );
  NAND U35927 ( .A(y[8040]), .B(x[490]), .Z(n34768) );
  XNOR U35928 ( .A(n34769), .B(n34768), .Z(n34889) );
  ANDN U35929 ( .B(o[369]), .A(n34770), .Z(n34888) );
  XOR U35930 ( .A(n34889), .B(n34888), .Z(n34921) );
  AND U35931 ( .A(y[8035]), .B(x[495]), .Z(n34772) );
  NAND U35932 ( .A(y[8041]), .B(x[489]), .Z(n34771) );
  XNOR U35933 ( .A(n34772), .B(n34771), .Z(n34879) );
  NAND U35934 ( .A(x[494]), .B(y[8036]), .Z(n34880) );
  XOR U35935 ( .A(n34879), .B(n34880), .Z(n34922) );
  XNOR U35936 ( .A(n34921), .B(n34922), .Z(n34923) );
  XNOR U35937 ( .A(n34924), .B(n34923), .Z(n34933) );
  XOR U35938 ( .A(n34934), .B(n34933), .Z(n34936) );
  NANDN U35939 ( .A(n34774), .B(n34773), .Z(n34778) );
  NANDN U35940 ( .A(n34776), .B(n34775), .Z(n34777) );
  AND U35941 ( .A(n34778), .B(n34777), .Z(n34946) );
  AND U35942 ( .A(y[8034]), .B(x[496]), .Z(n34780) );
  NAND U35943 ( .A(y[8039]), .B(x[491]), .Z(n34779) );
  XNOR U35944 ( .A(n34780), .B(n34779), .Z(n34875) );
  NAND U35945 ( .A(x[482]), .B(y[8048]), .Z(n34876) );
  XNOR U35946 ( .A(n34875), .B(n34876), .Z(n34945) );
  AND U35947 ( .A(y[8045]), .B(x[485]), .Z(n35006) );
  NAND U35948 ( .A(y[8044]), .B(x[486]), .Z(n34781) );
  XNOR U35949 ( .A(n35006), .B(n34781), .Z(n34871) );
  NAND U35950 ( .A(y[8046]), .B(x[484]), .Z(n34782) );
  XNOR U35951 ( .A(n35678), .B(n34782), .Z(n34908) );
  AND U35952 ( .A(x[487]), .B(y[8043]), .Z(n34909) );
  XNOR U35953 ( .A(n34908), .B(n34909), .Z(n34872) );
  XNOR U35954 ( .A(n34871), .B(n34872), .Z(n34947) );
  XOR U35955 ( .A(n34948), .B(n34947), .Z(n34935) );
  XNOR U35956 ( .A(n34936), .B(n34935), .Z(n34858) );
  NAND U35957 ( .A(n34784), .B(n34783), .Z(n34788) );
  NAND U35958 ( .A(n34786), .B(n34785), .Z(n34787) );
  AND U35959 ( .A(n34788), .B(n34787), .Z(n34927) );
  NAND U35960 ( .A(n34790), .B(n34789), .Z(n34794) );
  NAND U35961 ( .A(n34792), .B(n34791), .Z(n34793) );
  AND U35962 ( .A(n34794), .B(n34793), .Z(n34928) );
  XOR U35963 ( .A(n34927), .B(n34928), .Z(n34929) );
  NAND U35964 ( .A(n34796), .B(n34795), .Z(n34800) );
  NAND U35965 ( .A(n34798), .B(n34797), .Z(n34799) );
  AND U35966 ( .A(n34800), .B(n34799), .Z(n34930) );
  XOR U35967 ( .A(n34929), .B(n34930), .Z(n34857) );
  XOR U35968 ( .A(n34858), .B(n34857), .Z(n34860) );
  AND U35969 ( .A(x[488]), .B(y[8044]), .Z(n35130) );
  NAND U35970 ( .A(n35130), .B(n34801), .Z(n34805) );
  NAND U35971 ( .A(n34803), .B(n34802), .Z(n34804) );
  NAND U35972 ( .A(n34805), .B(n34804), .Z(n34940) );
  AND U35973 ( .A(x[489]), .B(y[8048]), .Z(n35784) );
  NAND U35974 ( .A(n35784), .B(n34887), .Z(n34809) );
  NANDN U35975 ( .A(n34807), .B(n34806), .Z(n34808) );
  NAND U35976 ( .A(n34809), .B(n34808), .Z(n34939) );
  XOR U35977 ( .A(n34940), .B(n34939), .Z(n34942) );
  AND U35978 ( .A(x[490]), .B(y[8047]), .Z(n35701) );
  IV U35979 ( .A(n35701), .Z(n35783) );
  NANDN U35980 ( .A(n35783), .B(n34810), .Z(n34814) );
  NANDN U35981 ( .A(n34812), .B(n34811), .Z(n34813) );
  AND U35982 ( .A(n34814), .B(n34813), .Z(n34918) );
  AND U35983 ( .A(x[480]), .B(y[8050]), .Z(n34890) );
  NAND U35984 ( .A(x[498]), .B(y[8032]), .Z(n34891) );
  XNOR U35985 ( .A(n34890), .B(n34891), .Z(n34892) );
  NAND U35986 ( .A(x[497]), .B(y[8033]), .Z(n34912) );
  XOR U35987 ( .A(o[370]), .B(n34912), .Z(n34893) );
  XNOR U35988 ( .A(n34892), .B(n34893), .Z(n34915) );
  AND U35989 ( .A(y[8037]), .B(x[493]), .Z(n34816) );
  NAND U35990 ( .A(y[8047]), .B(x[483]), .Z(n34815) );
  XNOR U35991 ( .A(n34816), .B(n34815), .Z(n34898) );
  NAND U35992 ( .A(x[492]), .B(y[8038]), .Z(n34899) );
  XOR U35993 ( .A(n34898), .B(n34899), .Z(n34916) );
  XNOR U35994 ( .A(n34915), .B(n34916), .Z(n34917) );
  XNOR U35995 ( .A(n34918), .B(n34917), .Z(n34941) );
  XOR U35996 ( .A(n34942), .B(n34941), .Z(n34864) );
  NAND U35997 ( .A(n34818), .B(n34817), .Z(n34822) );
  NANDN U35998 ( .A(n34820), .B(n34819), .Z(n34821) );
  AND U35999 ( .A(n34822), .B(n34821), .Z(n34863) );
  XNOR U36000 ( .A(n34864), .B(n34863), .Z(n34865) );
  NANDN U36001 ( .A(n34824), .B(n34823), .Z(n34828) );
  NANDN U36002 ( .A(n34826), .B(n34825), .Z(n34827) );
  NAND U36003 ( .A(n34828), .B(n34827), .Z(n34866) );
  XNOR U36004 ( .A(n34865), .B(n34866), .Z(n34859) );
  XNOR U36005 ( .A(n34860), .B(n34859), .Z(n34854) );
  NAND U36006 ( .A(n34830), .B(n34829), .Z(n34834) );
  NAND U36007 ( .A(n34832), .B(n34831), .Z(n34833) );
  NAND U36008 ( .A(n34834), .B(n34833), .Z(n34852) );
  NAND U36009 ( .A(n34836), .B(n34835), .Z(n34840) );
  NAND U36010 ( .A(n34838), .B(n34837), .Z(n34839) );
  NAND U36011 ( .A(n34840), .B(n34839), .Z(n34851) );
  XOR U36012 ( .A(n34852), .B(n34851), .Z(n34853) );
  XOR U36013 ( .A(n34854), .B(n34853), .Z(n34951) );
  XOR U36014 ( .A(n34952), .B(n34951), .Z(n34953) );
  XNOR U36015 ( .A(n34954), .B(n34953), .Z(n34959) );
  NAND U36016 ( .A(n34845), .B(n34844), .Z(n34849) );
  NANDN U36017 ( .A(n34847), .B(n34846), .Z(n34848) );
  NAND U36018 ( .A(n34849), .B(n34848), .Z(n34957) );
  XOR U36019 ( .A(n34958), .B(n34957), .Z(n34850) );
  XNOR U36020 ( .A(n34959), .B(n34850), .Z(N755) );
  NAND U36021 ( .A(n34852), .B(n34851), .Z(n34856) );
  NAND U36022 ( .A(n34854), .B(n34853), .Z(n34855) );
  AND U36023 ( .A(n34856), .B(n34855), .Z(n35074) );
  NAND U36024 ( .A(n34858), .B(n34857), .Z(n34862) );
  NAND U36025 ( .A(n34860), .B(n34859), .Z(n34861) );
  AND U36026 ( .A(n34862), .B(n34861), .Z(n35072) );
  NANDN U36027 ( .A(n34864), .B(n34863), .Z(n34868) );
  NANDN U36028 ( .A(n34866), .B(n34865), .Z(n34867) );
  AND U36029 ( .A(n34868), .B(n34867), .Z(n35052) );
  AND U36030 ( .A(x[486]), .B(y[8045]), .Z(n34870) );
  NAND U36031 ( .A(n34870), .B(n34869), .Z(n34874) );
  NANDN U36032 ( .A(n34872), .B(n34871), .Z(n34873) );
  AND U36033 ( .A(n34874), .B(n34873), .Z(n35046) );
  AND U36034 ( .A(x[496]), .B(y[8039]), .Z(n35397) );
  NAND U36035 ( .A(n35397), .B(n35223), .Z(n34878) );
  NANDN U36036 ( .A(n34876), .B(n34875), .Z(n34877) );
  AND U36037 ( .A(n34878), .B(n34877), .Z(n35045) );
  AND U36038 ( .A(x[495]), .B(y[8041]), .Z(n35712) );
  NAND U36039 ( .A(n35712), .B(n34973), .Z(n34882) );
  NANDN U36040 ( .A(n34880), .B(n34879), .Z(n34881) );
  NAND U36041 ( .A(n34882), .B(n34881), .Z(n34964) );
  AND U36042 ( .A(y[8050]), .B(x[481]), .Z(n34884) );
  NAND U36043 ( .A(y[8043]), .B(x[488]), .Z(n34883) );
  XNOR U36044 ( .A(n34884), .B(n34883), .Z(n35023) );
  AND U36045 ( .A(y[8038]), .B(x[493]), .Z(n34886) );
  NAND U36046 ( .A(y[8049]), .B(x[482]), .Z(n34885) );
  XNOR U36047 ( .A(n34886), .B(n34885), .Z(n34979) );
  XOR U36048 ( .A(n34962), .B(n34961), .Z(n34963) );
  XOR U36049 ( .A(n34964), .B(n34963), .Z(n35044) );
  XOR U36050 ( .A(n35045), .B(n35044), .Z(n35047) );
  XOR U36051 ( .A(n35046), .B(n35047), .Z(n35051) );
  NAND U36052 ( .A(x[490]), .B(y[8049]), .Z(n36093) );
  NANDN U36053 ( .A(n34891), .B(n34890), .Z(n34895) );
  NANDN U36054 ( .A(n34893), .B(n34892), .Z(n34894) );
  NAND U36055 ( .A(n34895), .B(n34894), .Z(n35001) );
  AND U36056 ( .A(y[8035]), .B(x[496]), .Z(n35644) );
  NAND U36057 ( .A(y[8042]), .B(x[489]), .Z(n34896) );
  XNOR U36058 ( .A(n35644), .B(n34896), .Z(n34974) );
  AND U36059 ( .A(x[495]), .B(y[8036]), .Z(n34975) );
  XOR U36060 ( .A(n34974), .B(n34975), .Z(n35000) );
  XOR U36061 ( .A(n35001), .B(n35000), .Z(n35002) );
  XNOR U36062 ( .A(n35003), .B(n35002), .Z(n35040) );
  AND U36063 ( .A(x[493]), .B(y[8047]), .Z(n36264) );
  NANDN U36064 ( .A(n34897), .B(n36264), .Z(n34901) );
  NANDN U36065 ( .A(n34899), .B(n34898), .Z(n34900) );
  NAND U36066 ( .A(n34901), .B(n34900), .Z(n34997) );
  AND U36067 ( .A(y[8041]), .B(x[490]), .Z(n34903) );
  NAND U36068 ( .A(y[8034]), .B(x[497]), .Z(n34902) );
  XNOR U36069 ( .A(n34903), .B(n34902), .Z(n35029) );
  AND U36070 ( .A(x[498]), .B(y[8033]), .Z(n34993) );
  XOR U36071 ( .A(o[371]), .B(n34993), .Z(n35028) );
  XOR U36072 ( .A(n35029), .B(n35028), .Z(n34995) );
  NAND U36073 ( .A(y[8048]), .B(x[483]), .Z(n34904) );
  XNOR U36074 ( .A(n34905), .B(n34904), .Z(n34987) );
  XOR U36075 ( .A(n34995), .B(n34994), .Z(n34996) );
  XNOR U36076 ( .A(n34997), .B(n34996), .Z(n35039) );
  NAND U36077 ( .A(n34907), .B(n34906), .Z(n34911) );
  NAND U36078 ( .A(n34909), .B(n34908), .Z(n34910) );
  AND U36079 ( .A(n34911), .B(n34910), .Z(n34970) );
  AND U36080 ( .A(x[480]), .B(y[8051]), .Z(n35010) );
  AND U36081 ( .A(x[499]), .B(y[8032]), .Z(n35011) );
  XOR U36082 ( .A(n35010), .B(n35011), .Z(n35013) );
  ANDN U36083 ( .B(o[370]), .A(n34912), .Z(n35012) );
  XOR U36084 ( .A(n35013), .B(n35012), .Z(n34968) );
  AND U36085 ( .A(x[484]), .B(y[8047]), .Z(n35144) );
  AND U36086 ( .A(y[8046]), .B(x[485]), .Z(n34914) );
  NAND U36087 ( .A(y[8045]), .B(x[486]), .Z(n34913) );
  XNOR U36088 ( .A(n34914), .B(n34913), .Z(n35007) );
  XOR U36089 ( .A(n35144), .B(n35007), .Z(n34967) );
  XOR U36090 ( .A(n34968), .B(n34967), .Z(n34969) );
  XOR U36091 ( .A(n34970), .B(n34969), .Z(n35038) );
  XNOR U36092 ( .A(n35039), .B(n35038), .Z(n35041) );
  XOR U36093 ( .A(n35040), .B(n35041), .Z(n35034) );
  NANDN U36094 ( .A(n34916), .B(n34915), .Z(n34920) );
  NANDN U36095 ( .A(n34918), .B(n34917), .Z(n34919) );
  AND U36096 ( .A(n34920), .B(n34919), .Z(n35033) );
  NANDN U36097 ( .A(n34922), .B(n34921), .Z(n34926) );
  NANDN U36098 ( .A(n34924), .B(n34923), .Z(n34925) );
  NAND U36099 ( .A(n34926), .B(n34925), .Z(n35032) );
  XOR U36100 ( .A(n35033), .B(n35032), .Z(n35035) );
  XOR U36101 ( .A(n35034), .B(n35035), .Z(n35050) );
  XOR U36102 ( .A(n35051), .B(n35050), .Z(n35053) );
  XNOR U36103 ( .A(n35052), .B(n35053), .Z(n35065) );
  NAND U36104 ( .A(n34928), .B(n34927), .Z(n34932) );
  NAND U36105 ( .A(n34930), .B(n34929), .Z(n34931) );
  AND U36106 ( .A(n34932), .B(n34931), .Z(n35063) );
  NAND U36107 ( .A(n34934), .B(n34933), .Z(n34938) );
  NAND U36108 ( .A(n34936), .B(n34935), .Z(n34937) );
  AND U36109 ( .A(n34938), .B(n34937), .Z(n35059) );
  NAND U36110 ( .A(n34940), .B(n34939), .Z(n34944) );
  NAND U36111 ( .A(n34942), .B(n34941), .Z(n34943) );
  AND U36112 ( .A(n34944), .B(n34943), .Z(n35057) );
  NANDN U36113 ( .A(n34946), .B(n34945), .Z(n34950) );
  NAND U36114 ( .A(n34948), .B(n34947), .Z(n34949) );
  NAND U36115 ( .A(n34950), .B(n34949), .Z(n35056) );
  XOR U36116 ( .A(n35063), .B(n35062), .Z(n35064) );
  XOR U36117 ( .A(n35065), .B(n35064), .Z(n35071) );
  XOR U36118 ( .A(n35072), .B(n35071), .Z(n35073) );
  XOR U36119 ( .A(n35074), .B(n35073), .Z(n35070) );
  NAND U36120 ( .A(n34952), .B(n34951), .Z(n34956) );
  NAND U36121 ( .A(n34954), .B(n34953), .Z(n34955) );
  NAND U36122 ( .A(n34956), .B(n34955), .Z(n35068) );
  XOR U36123 ( .A(n35068), .B(n35069), .Z(n34960) );
  XNOR U36124 ( .A(n35070), .B(n34960), .Z(N756) );
  NAND U36125 ( .A(n34962), .B(n34961), .Z(n34966) );
  NAND U36126 ( .A(n34964), .B(n34963), .Z(n34965) );
  NAND U36127 ( .A(n34966), .B(n34965), .Z(n35079) );
  NAND U36128 ( .A(n34968), .B(n34967), .Z(n34972) );
  NANDN U36129 ( .A(n34970), .B(n34969), .Z(n34971) );
  NAND U36130 ( .A(n34972), .B(n34971), .Z(n35078) );
  XOR U36131 ( .A(n35079), .B(n35078), .Z(n35081) );
  AND U36132 ( .A(x[496]), .B(y[8042]), .Z(n36006) );
  NAND U36133 ( .A(n36006), .B(n34973), .Z(n34977) );
  NAND U36134 ( .A(n34975), .B(n34974), .Z(n34976) );
  NAND U36135 ( .A(n34977), .B(n34976), .Z(n35119) );
  AND U36136 ( .A(x[493]), .B(y[8049]), .Z(n36482) );
  NAND U36137 ( .A(n36482), .B(n34978), .Z(n34982) );
  NANDN U36138 ( .A(n34980), .B(n34979), .Z(n34981) );
  NAND U36139 ( .A(n34982), .B(n34981), .Z(n35164) );
  AND U36140 ( .A(y[8036]), .B(x[496]), .Z(n34984) );
  NAND U36141 ( .A(y[8042]), .B(x[490]), .Z(n34983) );
  XNOR U36142 ( .A(n34984), .B(n34983), .Z(n35125) );
  AND U36143 ( .A(x[482]), .B(y[8050]), .Z(n35126) );
  XOR U36144 ( .A(n35125), .B(n35126), .Z(n35162) );
  NAND U36145 ( .A(y[8043]), .B(x[489]), .Z(n34985) );
  XNOR U36146 ( .A(n34986), .B(n34985), .Z(n35095) );
  AND U36147 ( .A(x[494]), .B(y[8038]), .Z(n35096) );
  XOR U36148 ( .A(n35095), .B(n35096), .Z(n35161) );
  XOR U36149 ( .A(n35162), .B(n35161), .Z(n35163) );
  XOR U36150 ( .A(n35164), .B(n35163), .Z(n35118) );
  XOR U36151 ( .A(n35119), .B(n35118), .Z(n35121) );
  NAND U36152 ( .A(x[491]), .B(y[8048]), .Z(n36094) );
  NANDN U36153 ( .A(n36094), .B(n35262), .Z(n34990) );
  NANDN U36154 ( .A(n34988), .B(n34987), .Z(n34989) );
  NAND U36155 ( .A(n34990), .B(n34989), .Z(n35170) );
  AND U36156 ( .A(y[8041]), .B(x[491]), .Z(n34992) );
  NAND U36157 ( .A(y[8051]), .B(x[481]), .Z(n34991) );
  XNOR U36158 ( .A(n34992), .B(n34991), .Z(n35091) );
  AND U36159 ( .A(x[499]), .B(y[8033]), .Z(n35099) );
  XOR U36160 ( .A(o[372]), .B(n35099), .Z(n35090) );
  XOR U36161 ( .A(n35091), .B(n35090), .Z(n35168) );
  AND U36162 ( .A(x[480]), .B(y[8052]), .Z(n35149) );
  AND U36163 ( .A(x[500]), .B(y[8032]), .Z(n35150) );
  XOR U36164 ( .A(n35149), .B(n35150), .Z(n35152) );
  AND U36165 ( .A(o[371]), .B(n34993), .Z(n35151) );
  XOR U36166 ( .A(n35152), .B(n35151), .Z(n35167) );
  XOR U36167 ( .A(n35168), .B(n35167), .Z(n35169) );
  XOR U36168 ( .A(n35170), .B(n35169), .Z(n35120) );
  XOR U36169 ( .A(n35121), .B(n35120), .Z(n35080) );
  XNOR U36170 ( .A(n35081), .B(n35080), .Z(n35176) );
  NAND U36171 ( .A(n34995), .B(n34994), .Z(n34999) );
  NAND U36172 ( .A(n34997), .B(n34996), .Z(n34998) );
  AND U36173 ( .A(n34999), .B(n34998), .Z(n35174) );
  NAND U36174 ( .A(n35001), .B(n35000), .Z(n35005) );
  NAND U36175 ( .A(n35003), .B(n35002), .Z(n35004) );
  AND U36176 ( .A(n35005), .B(n35004), .Z(n35115) );
  NAND U36177 ( .A(x[486]), .B(y[8046]), .Z(n35101) );
  NANDN U36178 ( .A(n35101), .B(n35006), .Z(n35009) );
  NAND U36179 ( .A(n35007), .B(n35144), .Z(n35008) );
  NAND U36180 ( .A(n35009), .B(n35008), .Z(n35109) );
  NAND U36181 ( .A(n35011), .B(n35010), .Z(n35015) );
  NAND U36182 ( .A(n35013), .B(n35012), .Z(n35014) );
  NAND U36183 ( .A(n35015), .B(n35014), .Z(n35107) );
  AND U36184 ( .A(y[8034]), .B(x[498]), .Z(n35017) );
  NAND U36185 ( .A(y[8040]), .B(x[492]), .Z(n35016) );
  XNOR U36186 ( .A(n35017), .B(n35016), .Z(n35085) );
  AND U36187 ( .A(x[497]), .B(y[8035]), .Z(n35086) );
  XOR U36188 ( .A(n35085), .B(n35086), .Z(n35106) );
  XOR U36189 ( .A(n35107), .B(n35106), .Z(n35108) );
  XNOR U36190 ( .A(n35109), .B(n35108), .Z(n35113) );
  AND U36191 ( .A(y[8039]), .B(x[493]), .Z(n35019) );
  NAND U36192 ( .A(y[8049]), .B(x[483]), .Z(n35018) );
  XNOR U36193 ( .A(n35019), .B(n35018), .Z(n35131) );
  XNOR U36194 ( .A(n35131), .B(n35130), .Z(n35103) );
  AND U36195 ( .A(y[8047]), .B(x[485]), .Z(n35021) );
  NAND U36196 ( .A(y[8048]), .B(x[484]), .Z(n35020) );
  XNOR U36197 ( .A(n35021), .B(n35020), .Z(n35146) );
  AND U36198 ( .A(x[487]), .B(y[8045]), .Z(n35145) );
  XNOR U36199 ( .A(n35146), .B(n35145), .Z(n35100) );
  XOR U36200 ( .A(n35101), .B(n35100), .Z(n35102) );
  XNOR U36201 ( .A(n35103), .B(n35102), .Z(n35157) );
  AND U36202 ( .A(x[488]), .B(y[8050]), .Z(n36224) );
  AND U36203 ( .A(x[481]), .B(y[8043]), .Z(n35022) );
  NAND U36204 ( .A(n36224), .B(n35022), .Z(n35026) );
  NANDN U36205 ( .A(n35024), .B(n35023), .Z(n35025) );
  NAND U36206 ( .A(n35026), .B(n35025), .Z(n35156) );
  AND U36207 ( .A(x[497]), .B(y[8041]), .Z(n35863) );
  IV U36208 ( .A(n35863), .Z(n36015) );
  NANDN U36209 ( .A(n36015), .B(n35027), .Z(n35031) );
  NAND U36210 ( .A(n35029), .B(n35028), .Z(n35030) );
  NAND U36211 ( .A(n35031), .B(n35030), .Z(n35155) );
  XOR U36212 ( .A(n35156), .B(n35155), .Z(n35158) );
  XNOR U36213 ( .A(n35157), .B(n35158), .Z(n35112) );
  XOR U36214 ( .A(n35113), .B(n35112), .Z(n35114) );
  XOR U36215 ( .A(n35115), .B(n35114), .Z(n35173) );
  XOR U36216 ( .A(n35174), .B(n35173), .Z(n35175) );
  XNOR U36217 ( .A(n35176), .B(n35175), .Z(n35180) );
  NANDN U36218 ( .A(n35033), .B(n35032), .Z(n35037) );
  NANDN U36219 ( .A(n35035), .B(n35034), .Z(n35036) );
  AND U36220 ( .A(n35037), .B(n35036), .Z(n35188) );
  NAND U36221 ( .A(n35039), .B(n35038), .Z(n35043) );
  NANDN U36222 ( .A(n35041), .B(n35040), .Z(n35042) );
  AND U36223 ( .A(n35043), .B(n35042), .Z(n35186) );
  NANDN U36224 ( .A(n35045), .B(n35044), .Z(n35049) );
  OR U36225 ( .A(n35047), .B(n35046), .Z(n35048) );
  AND U36226 ( .A(n35049), .B(n35048), .Z(n35185) );
  XNOR U36227 ( .A(n35186), .B(n35185), .Z(n35187) );
  XNOR U36228 ( .A(n35188), .B(n35187), .Z(n35179) );
  XOR U36229 ( .A(n35180), .B(n35179), .Z(n35182) );
  NANDN U36230 ( .A(n35051), .B(n35050), .Z(n35055) );
  OR U36231 ( .A(n35053), .B(n35052), .Z(n35054) );
  AND U36232 ( .A(n35055), .B(n35054), .Z(n35181) );
  XOR U36233 ( .A(n35182), .B(n35181), .Z(n35201) );
  NANDN U36234 ( .A(n35057), .B(n35056), .Z(n35061) );
  NANDN U36235 ( .A(n35059), .B(n35058), .Z(n35060) );
  AND U36236 ( .A(n35061), .B(n35060), .Z(n35198) );
  NAND U36237 ( .A(n35063), .B(n35062), .Z(n35067) );
  NAND U36238 ( .A(n35065), .B(n35064), .Z(n35066) );
  AND U36239 ( .A(n35067), .B(n35066), .Z(n35199) );
  XOR U36240 ( .A(n35198), .B(n35199), .Z(n35200) );
  XOR U36241 ( .A(n35201), .B(n35200), .Z(n35194) );
  NAND U36242 ( .A(n35072), .B(n35071), .Z(n35076) );
  NANDN U36243 ( .A(n35074), .B(n35073), .Z(n35075) );
  AND U36244 ( .A(n35076), .B(n35075), .Z(n35193) );
  IV U36245 ( .A(n35193), .Z(n35191) );
  XOR U36246 ( .A(n35192), .B(n35191), .Z(n35077) );
  XNOR U36247 ( .A(n35194), .B(n35077), .Z(N757) );
  NAND U36248 ( .A(n35079), .B(n35078), .Z(n35083) );
  NAND U36249 ( .A(n35081), .B(n35080), .Z(n35082) );
  NAND U36250 ( .A(n35083), .B(n35082), .Z(n35214) );
  AND U36251 ( .A(x[498]), .B(y[8040]), .Z(n36013) );
  NAND U36252 ( .A(n36013), .B(n35084), .Z(n35088) );
  NAND U36253 ( .A(n35086), .B(n35085), .Z(n35087) );
  NAND U36254 ( .A(n35088), .B(n35087), .Z(n35291) );
  AND U36255 ( .A(x[491]), .B(y[8051]), .Z(n36612) );
  AND U36256 ( .A(x[481]), .B(y[8041]), .Z(n35089) );
  NAND U36257 ( .A(n36612), .B(n35089), .Z(n35093) );
  NAND U36258 ( .A(n35091), .B(n35090), .Z(n35092) );
  NAND U36259 ( .A(n35093), .B(n35092), .Z(n35290) );
  XOR U36260 ( .A(n35291), .B(n35290), .Z(n35293) );
  AND U36261 ( .A(x[495]), .B(y[8043]), .Z(n36001) );
  NAND U36262 ( .A(n36001), .B(n35094), .Z(n35098) );
  NAND U36263 ( .A(n35096), .B(n35095), .Z(n35097) );
  NAND U36264 ( .A(n35098), .B(n35097), .Z(n35249) );
  AND U36265 ( .A(x[480]), .B(y[8053]), .Z(n35268) );
  AND U36266 ( .A(x[501]), .B(y[8032]), .Z(n35269) );
  XOR U36267 ( .A(n35268), .B(n35269), .Z(n35271) );
  AND U36268 ( .A(o[372]), .B(n35099), .Z(n35270) );
  XOR U36269 ( .A(n35271), .B(n35270), .Z(n35247) );
  AND U36270 ( .A(x[485]), .B(y[8048]), .Z(n35255) );
  AND U36271 ( .A(x[496]), .B(y[8037]), .Z(n35254) );
  XOR U36272 ( .A(n35255), .B(n35254), .Z(n35253) );
  AND U36273 ( .A(x[495]), .B(y[8038]), .Z(n35252) );
  XOR U36274 ( .A(n35253), .B(n35252), .Z(n35246) );
  XOR U36275 ( .A(n35247), .B(n35246), .Z(n35248) );
  XOR U36276 ( .A(n35249), .B(n35248), .Z(n35292) );
  XNOR U36277 ( .A(n35293), .B(n35292), .Z(n35285) );
  NAND U36278 ( .A(n35101), .B(n35100), .Z(n35105) );
  NAND U36279 ( .A(n35103), .B(n35102), .Z(n35104) );
  NAND U36280 ( .A(n35105), .B(n35104), .Z(n35284) );
  XOR U36281 ( .A(n35285), .B(n35284), .Z(n35287) );
  NAND U36282 ( .A(n35107), .B(n35106), .Z(n35111) );
  NAND U36283 ( .A(n35109), .B(n35108), .Z(n35110) );
  AND U36284 ( .A(n35111), .B(n35110), .Z(n35286) );
  XNOR U36285 ( .A(n35287), .B(n35286), .Z(n35212) );
  NAND U36286 ( .A(n35113), .B(n35112), .Z(n35117) );
  NAND U36287 ( .A(n35115), .B(n35114), .Z(n35116) );
  AND U36288 ( .A(n35117), .B(n35116), .Z(n35211) );
  XOR U36289 ( .A(n35212), .B(n35211), .Z(n35213) );
  XNOR U36290 ( .A(n35214), .B(n35213), .Z(n35207) );
  NAND U36291 ( .A(n35119), .B(n35118), .Z(n35123) );
  NAND U36292 ( .A(n35121), .B(n35120), .Z(n35122) );
  NAND U36293 ( .A(n35123), .B(n35122), .Z(n35311) );
  NAND U36294 ( .A(n36006), .B(n35124), .Z(n35128) );
  NAND U36295 ( .A(n35126), .B(n35125), .Z(n35127) );
  NAND U36296 ( .A(n35128), .B(n35127), .Z(n35218) );
  NAND U36297 ( .A(n35129), .B(n36482), .Z(n35133) );
  NAND U36298 ( .A(n35131), .B(n35130), .Z(n35132) );
  NAND U36299 ( .A(n35133), .B(n35132), .Z(n35305) );
  AND U36300 ( .A(y[8035]), .B(x[498]), .Z(n35135) );
  NAND U36301 ( .A(y[8043]), .B(x[490]), .Z(n35134) );
  XNOR U36302 ( .A(n35135), .B(n35134), .Z(n35275) );
  AND U36303 ( .A(x[481]), .B(y[8052]), .Z(n35276) );
  XOR U36304 ( .A(n35275), .B(n35276), .Z(n35303) );
  AND U36305 ( .A(y[8034]), .B(x[499]), .Z(n35137) );
  NAND U36306 ( .A(y[8042]), .B(x[491]), .Z(n35136) );
  XNOR U36307 ( .A(n35137), .B(n35136), .Z(n35225) );
  AND U36308 ( .A(x[500]), .B(y[8033]), .Z(n35267) );
  XOR U36309 ( .A(o[373]), .B(n35267), .Z(n35224) );
  XOR U36310 ( .A(n35225), .B(n35224), .Z(n35302) );
  XOR U36311 ( .A(n35303), .B(n35302), .Z(n35304) );
  XOR U36312 ( .A(n35305), .B(n35304), .Z(n35217) );
  XOR U36313 ( .A(n35218), .B(n35217), .Z(n35220) );
  AND U36314 ( .A(x[487]), .B(y[8046]), .Z(n35480) );
  AND U36315 ( .A(y[8047]), .B(x[486]), .Z(n35139) );
  NAND U36316 ( .A(y[8039]), .B(x[494]), .Z(n35138) );
  XNOR U36317 ( .A(n35139), .B(n35138), .Z(n35279) );
  XNOR U36318 ( .A(n35480), .B(n35279), .Z(n35237) );
  NAND U36319 ( .A(x[489]), .B(y[8044]), .Z(n35235) );
  NAND U36320 ( .A(x[488]), .B(y[8045]), .Z(n35234) );
  XOR U36321 ( .A(n35235), .B(n35234), .Z(n35236) );
  XNOR U36322 ( .A(n35237), .B(n35236), .Z(n35242) );
  AND U36323 ( .A(y[8041]), .B(x[492]), .Z(n35141) );
  NAND U36324 ( .A(y[8036]), .B(x[497]), .Z(n35140) );
  XNOR U36325 ( .A(n35141), .B(n35140), .Z(n35228) );
  AND U36326 ( .A(x[482]), .B(y[8051]), .Z(n35229) );
  XOR U36327 ( .A(n35228), .B(n35229), .Z(n35241) );
  AND U36328 ( .A(y[8040]), .B(x[493]), .Z(n35143) );
  NAND U36329 ( .A(y[8050]), .B(x[483]), .Z(n35142) );
  XNOR U36330 ( .A(n35143), .B(n35142), .Z(n35263) );
  AND U36331 ( .A(x[484]), .B(y[8049]), .Z(n35264) );
  XOR U36332 ( .A(n35263), .B(n35264), .Z(n35240) );
  XOR U36333 ( .A(n35241), .B(n35240), .Z(n35243) );
  XOR U36334 ( .A(n35242), .B(n35243), .Z(n35299) );
  NAND U36335 ( .A(n35255), .B(n35144), .Z(n35148) );
  NAND U36336 ( .A(n35146), .B(n35145), .Z(n35147) );
  NAND U36337 ( .A(n35148), .B(n35147), .Z(n35297) );
  NAND U36338 ( .A(n35150), .B(n35149), .Z(n35154) );
  NAND U36339 ( .A(n35152), .B(n35151), .Z(n35153) );
  NAND U36340 ( .A(n35154), .B(n35153), .Z(n35296) );
  XOR U36341 ( .A(n35297), .B(n35296), .Z(n35298) );
  XOR U36342 ( .A(n35299), .B(n35298), .Z(n35219) );
  XOR U36343 ( .A(n35220), .B(n35219), .Z(n35309) );
  NAND U36344 ( .A(n35156), .B(n35155), .Z(n35160) );
  NAND U36345 ( .A(n35158), .B(n35157), .Z(n35159) );
  NAND U36346 ( .A(n35160), .B(n35159), .Z(n35316) );
  NAND U36347 ( .A(n35162), .B(n35161), .Z(n35166) );
  NAND U36348 ( .A(n35164), .B(n35163), .Z(n35165) );
  NAND U36349 ( .A(n35166), .B(n35165), .Z(n35315) );
  NAND U36350 ( .A(n35168), .B(n35167), .Z(n35172) );
  NAND U36351 ( .A(n35170), .B(n35169), .Z(n35171) );
  NAND U36352 ( .A(n35172), .B(n35171), .Z(n35314) );
  XOR U36353 ( .A(n35315), .B(n35314), .Z(n35317) );
  XOR U36354 ( .A(n35316), .B(n35317), .Z(n35308) );
  XOR U36355 ( .A(n35309), .B(n35308), .Z(n35310) );
  XNOR U36356 ( .A(n35311), .B(n35310), .Z(n35206) );
  NAND U36357 ( .A(n35174), .B(n35173), .Z(n35178) );
  NAND U36358 ( .A(n35176), .B(n35175), .Z(n35177) );
  NAND U36359 ( .A(n35178), .B(n35177), .Z(n35205) );
  XOR U36360 ( .A(n35206), .B(n35205), .Z(n35208) );
  XNOR U36361 ( .A(n35207), .B(n35208), .Z(n35325) );
  NAND U36362 ( .A(n35180), .B(n35179), .Z(n35184) );
  NAND U36363 ( .A(n35182), .B(n35181), .Z(n35183) );
  AND U36364 ( .A(n35184), .B(n35183), .Z(n35324) );
  NANDN U36365 ( .A(n35186), .B(n35185), .Z(n35190) );
  NAND U36366 ( .A(n35188), .B(n35187), .Z(n35189) );
  AND U36367 ( .A(n35190), .B(n35189), .Z(n35323) );
  XOR U36368 ( .A(n35324), .B(n35323), .Z(n35326) );
  XOR U36369 ( .A(n35325), .B(n35326), .Z(n35322) );
  NANDN U36370 ( .A(n35191), .B(n35192), .Z(n35197) );
  NOR U36371 ( .A(n35193), .B(n35192), .Z(n35195) );
  OR U36372 ( .A(n35195), .B(n35194), .Z(n35196) );
  AND U36373 ( .A(n35197), .B(n35196), .Z(n35320) );
  NAND U36374 ( .A(n35199), .B(n35198), .Z(n35203) );
  NANDN U36375 ( .A(n35201), .B(n35200), .Z(n35202) );
  AND U36376 ( .A(n35203), .B(n35202), .Z(n35321) );
  XOR U36377 ( .A(n35320), .B(n35321), .Z(n35204) );
  XNOR U36378 ( .A(n35322), .B(n35204), .Z(N758) );
  NAND U36379 ( .A(n35206), .B(n35205), .Z(n35210) );
  NAND U36380 ( .A(n35208), .B(n35207), .Z(n35209) );
  AND U36381 ( .A(n35210), .B(n35209), .Z(n35456) );
  NAND U36382 ( .A(n35212), .B(n35211), .Z(n35216) );
  NAND U36383 ( .A(n35214), .B(n35213), .Z(n35215) );
  NAND U36384 ( .A(n35216), .B(n35215), .Z(n35454) );
  NAND U36385 ( .A(n35218), .B(n35217), .Z(n35222) );
  NAND U36386 ( .A(n35220), .B(n35219), .Z(n35221) );
  AND U36387 ( .A(n35222), .B(n35221), .Z(n35447) );
  AND U36388 ( .A(x[499]), .B(y[8042]), .Z(n36381) );
  NAND U36389 ( .A(n36381), .B(n35223), .Z(n35227) );
  NAND U36390 ( .A(n35225), .B(n35224), .Z(n35226) );
  NAND U36391 ( .A(n35227), .B(n35226), .Z(n35439) );
  NANDN U36392 ( .A(n36015), .B(n35398), .Z(n35231) );
  NAND U36393 ( .A(n35229), .B(n35228), .Z(n35230) );
  NAND U36394 ( .A(n35231), .B(n35230), .Z(n35368) );
  AND U36395 ( .A(x[485]), .B(y[8049]), .Z(n35414) );
  AND U36396 ( .A(x[497]), .B(y[8037]), .Z(n35415) );
  XOR U36397 ( .A(n35414), .B(n35415), .Z(n35416) );
  AND U36398 ( .A(x[496]), .B(y[8038]), .Z(n35417) );
  XOR U36399 ( .A(n35416), .B(n35417), .Z(n35367) );
  AND U36400 ( .A(y[8036]), .B(x[498]), .Z(n35233) );
  NAND U36401 ( .A(y[8042]), .B(x[492]), .Z(n35232) );
  XNOR U36402 ( .A(n35233), .B(n35232), .Z(n35400) );
  AND U36403 ( .A(x[484]), .B(y[8050]), .Z(n35399) );
  XOR U36404 ( .A(n35400), .B(n35399), .Z(n35366) );
  XOR U36405 ( .A(n35367), .B(n35366), .Z(n35369) );
  XOR U36406 ( .A(n35368), .B(n35369), .Z(n35438) );
  XOR U36407 ( .A(n35439), .B(n35438), .Z(n35441) );
  NAND U36408 ( .A(n35235), .B(n35234), .Z(n35239) );
  NAND U36409 ( .A(n35237), .B(n35236), .Z(n35238) );
  AND U36410 ( .A(n35239), .B(n35238), .Z(n35440) );
  XOR U36411 ( .A(n35441), .B(n35440), .Z(n35445) );
  NAND U36412 ( .A(n35241), .B(n35240), .Z(n35245) );
  NAND U36413 ( .A(n35243), .B(n35242), .Z(n35244) );
  NAND U36414 ( .A(n35245), .B(n35244), .Z(n35427) );
  NAND U36415 ( .A(n35247), .B(n35246), .Z(n35251) );
  NAND U36416 ( .A(n35249), .B(n35248), .Z(n35250) );
  NAND U36417 ( .A(n35251), .B(n35250), .Z(n35426) );
  XOR U36418 ( .A(n35427), .B(n35426), .Z(n35429) );
  AND U36419 ( .A(n35253), .B(n35252), .Z(n35257) );
  NAND U36420 ( .A(n35255), .B(n35254), .Z(n35256) );
  NANDN U36421 ( .A(n35257), .B(n35256), .Z(n35389) );
  AND U36422 ( .A(y[8041]), .B(x[493]), .Z(n35259) );
  NAND U36423 ( .A(y[8034]), .B(x[500]), .Z(n35258) );
  XNOR U36424 ( .A(n35259), .B(n35258), .Z(n35410) );
  AND U36425 ( .A(x[482]), .B(y[8052]), .Z(n35411) );
  XOR U36426 ( .A(n35410), .B(n35411), .Z(n35387) );
  AND U36427 ( .A(y[8048]), .B(x[486]), .Z(n35261) );
  NAND U36428 ( .A(y[8039]), .B(x[495]), .Z(n35260) );
  XNOR U36429 ( .A(n35261), .B(n35260), .Z(n35422) );
  XOR U36430 ( .A(n35387), .B(n35386), .Z(n35388) );
  XOR U36431 ( .A(n35389), .B(n35388), .Z(n35433) );
  AND U36432 ( .A(x[493]), .B(y[8050]), .Z(n36614) );
  NAND U36433 ( .A(n35262), .B(n36614), .Z(n35266) );
  NAND U36434 ( .A(n35264), .B(n35263), .Z(n35265) );
  NAND U36435 ( .A(n35266), .B(n35265), .Z(n35357) );
  AND U36436 ( .A(x[481]), .B(y[8053]), .Z(n35380) );
  XOR U36437 ( .A(n35381), .B(n35380), .Z(n35379) );
  AND U36438 ( .A(o[373]), .B(n35267), .Z(n35378) );
  XOR U36439 ( .A(n35379), .B(n35378), .Z(n35355) );
  AND U36440 ( .A(x[494]), .B(y[8040]), .Z(n35372) );
  AND U36441 ( .A(x[483]), .B(y[8051]), .Z(n35373) );
  XOR U36442 ( .A(n35372), .B(n35373), .Z(n35374) );
  AND U36443 ( .A(x[499]), .B(y[8035]), .Z(n35375) );
  XOR U36444 ( .A(n35374), .B(n35375), .Z(n35354) );
  XOR U36445 ( .A(n35355), .B(n35354), .Z(n35356) );
  XOR U36446 ( .A(n35357), .B(n35356), .Z(n35432) );
  XOR U36447 ( .A(n35433), .B(n35432), .Z(n35435) );
  NAND U36448 ( .A(n35269), .B(n35268), .Z(n35273) );
  NAND U36449 ( .A(n35271), .B(n35270), .Z(n35272) );
  NAND U36450 ( .A(n35273), .B(n35272), .Z(n35349) );
  AND U36451 ( .A(x[498]), .B(y[8043]), .Z(n36383) );
  NAND U36452 ( .A(n36383), .B(n35274), .Z(n35278) );
  NAND U36453 ( .A(n35276), .B(n35275), .Z(n35277) );
  NAND U36454 ( .A(n35278), .B(n35277), .Z(n35348) );
  XOR U36455 ( .A(n35349), .B(n35348), .Z(n35351) );
  AND U36456 ( .A(x[494]), .B(y[8047]), .Z(n36418) );
  NAND U36457 ( .A(n35421), .B(n36418), .Z(n35281) );
  NAND U36458 ( .A(n35480), .B(n35279), .Z(n35280) );
  NAND U36459 ( .A(n35281), .B(n35280), .Z(n35363) );
  AND U36460 ( .A(x[480]), .B(y[8054]), .Z(n35403) );
  AND U36461 ( .A(x[502]), .B(y[8032]), .Z(n35404) );
  XOR U36462 ( .A(n35403), .B(n35404), .Z(n35406) );
  AND U36463 ( .A(x[501]), .B(y[8033]), .Z(n35420) );
  XOR U36464 ( .A(o[374]), .B(n35420), .Z(n35405) );
  XOR U36465 ( .A(n35406), .B(n35405), .Z(n35361) );
  AND U36466 ( .A(y[8047]), .B(x[487]), .Z(n35283) );
  NAND U36467 ( .A(y[8046]), .B(x[488]), .Z(n35282) );
  XNOR U36468 ( .A(n35283), .B(n35282), .Z(n35392) );
  XOR U36469 ( .A(n35361), .B(n35360), .Z(n35362) );
  XOR U36470 ( .A(n35363), .B(n35362), .Z(n35350) );
  XOR U36471 ( .A(n35351), .B(n35350), .Z(n35434) );
  XOR U36472 ( .A(n35435), .B(n35434), .Z(n35428) );
  XNOR U36473 ( .A(n35429), .B(n35428), .Z(n35444) );
  XOR U36474 ( .A(n35447), .B(n35446), .Z(n35339) );
  NAND U36475 ( .A(n35285), .B(n35284), .Z(n35289) );
  NAND U36476 ( .A(n35287), .B(n35286), .Z(n35288) );
  NAND U36477 ( .A(n35289), .B(n35288), .Z(n35337) );
  NAND U36478 ( .A(n35291), .B(n35290), .Z(n35295) );
  NAND U36479 ( .A(n35293), .B(n35292), .Z(n35294) );
  AND U36480 ( .A(n35295), .B(n35294), .Z(n35345) );
  NAND U36481 ( .A(n35297), .B(n35296), .Z(n35301) );
  NAND U36482 ( .A(n35299), .B(n35298), .Z(n35300) );
  NAND U36483 ( .A(n35301), .B(n35300), .Z(n35343) );
  NAND U36484 ( .A(n35303), .B(n35302), .Z(n35307) );
  NAND U36485 ( .A(n35305), .B(n35304), .Z(n35306) );
  NAND U36486 ( .A(n35307), .B(n35306), .Z(n35342) );
  XOR U36487 ( .A(n35343), .B(n35342), .Z(n35344) );
  XOR U36488 ( .A(n35345), .B(n35344), .Z(n35336) );
  XOR U36489 ( .A(n35337), .B(n35336), .Z(n35338) );
  XNOR U36490 ( .A(n35339), .B(n35338), .Z(n35333) );
  NAND U36491 ( .A(n35309), .B(n35308), .Z(n35313) );
  NAND U36492 ( .A(n35311), .B(n35310), .Z(n35312) );
  NAND U36493 ( .A(n35313), .B(n35312), .Z(n35331) );
  NAND U36494 ( .A(n35315), .B(n35314), .Z(n35319) );
  NAND U36495 ( .A(n35317), .B(n35316), .Z(n35318) );
  NAND U36496 ( .A(n35319), .B(n35318), .Z(n35330) );
  XOR U36497 ( .A(n35331), .B(n35330), .Z(n35332) );
  XOR U36498 ( .A(n35333), .B(n35332), .Z(n35453) );
  XOR U36499 ( .A(n35454), .B(n35453), .Z(n35455) );
  XNOR U36500 ( .A(n35456), .B(n35455), .Z(n35450) );
  NANDN U36501 ( .A(n35324), .B(n35323), .Z(n35328) );
  NANDN U36502 ( .A(n35326), .B(n35325), .Z(n35327) );
  AND U36503 ( .A(n35328), .B(n35327), .Z(n35452) );
  XOR U36504 ( .A(n35451), .B(n35452), .Z(n35329) );
  XNOR U36505 ( .A(n35450), .B(n35329), .Z(N759) );
  NAND U36506 ( .A(n35331), .B(n35330), .Z(n35335) );
  NAND U36507 ( .A(n35333), .B(n35332), .Z(n35334) );
  AND U36508 ( .A(n35335), .B(n35334), .Z(n35601) );
  NAND U36509 ( .A(n35337), .B(n35336), .Z(n35341) );
  NAND U36510 ( .A(n35339), .B(n35338), .Z(n35340) );
  NAND U36511 ( .A(n35341), .B(n35340), .Z(n35599) );
  NAND U36512 ( .A(n35343), .B(n35342), .Z(n35347) );
  NANDN U36513 ( .A(n35345), .B(n35344), .Z(n35346) );
  NAND U36514 ( .A(n35347), .B(n35346), .Z(n35576) );
  NAND U36515 ( .A(n35349), .B(n35348), .Z(n35353) );
  NAND U36516 ( .A(n35351), .B(n35350), .Z(n35352) );
  NAND U36517 ( .A(n35353), .B(n35352), .Z(n35570) );
  NAND U36518 ( .A(n35355), .B(n35354), .Z(n35359) );
  NAND U36519 ( .A(n35357), .B(n35356), .Z(n35358) );
  NAND U36520 ( .A(n35359), .B(n35358), .Z(n35568) );
  NAND U36521 ( .A(n35361), .B(n35360), .Z(n35365) );
  NAND U36522 ( .A(n35363), .B(n35362), .Z(n35364) );
  NAND U36523 ( .A(n35365), .B(n35364), .Z(n35567) );
  XOR U36524 ( .A(n35568), .B(n35567), .Z(n35569) );
  XOR U36525 ( .A(n35570), .B(n35569), .Z(n35588) );
  NAND U36526 ( .A(n35367), .B(n35366), .Z(n35371) );
  NAND U36527 ( .A(n35369), .B(n35368), .Z(n35370) );
  NAND U36528 ( .A(n35371), .B(n35370), .Z(n35586) );
  NAND U36529 ( .A(n35373), .B(n35372), .Z(n35377) );
  NAND U36530 ( .A(n35375), .B(n35374), .Z(n35376) );
  NAND U36531 ( .A(n35377), .B(n35376), .Z(n35514) );
  AND U36532 ( .A(n35379), .B(n35378), .Z(n35383) );
  NAND U36533 ( .A(n35381), .B(n35380), .Z(n35382) );
  NANDN U36534 ( .A(n35383), .B(n35382), .Z(n35513) );
  XOR U36535 ( .A(n35514), .B(n35513), .Z(n35516) );
  AND U36536 ( .A(y[8048]), .B(x[487]), .Z(n35385) );
  NAND U36537 ( .A(y[8046]), .B(x[489]), .Z(n35384) );
  XNOR U36538 ( .A(n35385), .B(n35384), .Z(n35481) );
  AND U36539 ( .A(x[490]), .B(y[8045]), .Z(n35520) );
  XOR U36540 ( .A(n35519), .B(n35520), .Z(n35522) );
  AND U36541 ( .A(x[486]), .B(y[8049]), .Z(n35472) );
  AND U36542 ( .A(x[495]), .B(y[8040]), .Z(n35473) );
  XOR U36543 ( .A(n35472), .B(n35473), .Z(n35474) );
  AND U36544 ( .A(x[491]), .B(y[8044]), .Z(n35475) );
  XOR U36545 ( .A(n35474), .B(n35475), .Z(n35521) );
  XOR U36546 ( .A(n35522), .B(n35521), .Z(n35515) );
  XOR U36547 ( .A(n35516), .B(n35515), .Z(n35585) );
  XOR U36548 ( .A(n35586), .B(n35585), .Z(n35587) );
  XOR U36549 ( .A(n35588), .B(n35587), .Z(n35574) );
  NAND U36550 ( .A(n35387), .B(n35386), .Z(n35391) );
  NAND U36551 ( .A(n35389), .B(n35388), .Z(n35390) );
  NAND U36552 ( .A(n35391), .B(n35390), .Z(n35508) );
  NANDN U36553 ( .A(n35482), .B(n35480), .Z(n35395) );
  NANDN U36554 ( .A(n35393), .B(n35392), .Z(n35394) );
  AND U36555 ( .A(n35395), .B(n35394), .Z(n35558) );
  AND U36556 ( .A(x[480]), .B(y[8055]), .Z(n35491) );
  AND U36557 ( .A(x[503]), .B(y[8032]), .Z(n35492) );
  XOR U36558 ( .A(n35491), .B(n35492), .Z(n35494) );
  AND U36559 ( .A(x[502]), .B(y[8033]), .Z(n35471) );
  XOR U36560 ( .A(o[375]), .B(n35471), .Z(n35493) );
  XOR U36561 ( .A(n35494), .B(n35493), .Z(n35556) );
  NAND U36562 ( .A(y[8035]), .B(x[500]), .Z(n35396) );
  XNOR U36563 ( .A(n35397), .B(n35396), .Z(n35467) );
  AND U36564 ( .A(x[499]), .B(y[8036]), .Z(n35468) );
  XOR U36565 ( .A(n35467), .B(n35468), .Z(n35555) );
  XOR U36566 ( .A(n35556), .B(n35555), .Z(n35557) );
  AND U36567 ( .A(x[498]), .B(y[8042]), .Z(n36253) );
  NAND U36568 ( .A(n36253), .B(n35398), .Z(n35402) );
  NAND U36569 ( .A(n35400), .B(n35399), .Z(n35401) );
  AND U36570 ( .A(n35402), .B(n35401), .Z(n35544) );
  NAND U36571 ( .A(n35404), .B(n35403), .Z(n35408) );
  NAND U36572 ( .A(n35406), .B(n35405), .Z(n35407) );
  NAND U36573 ( .A(n35408), .B(n35407), .Z(n35543) );
  XOR U36574 ( .A(n35546), .B(n35545), .Z(n35507) );
  XOR U36575 ( .A(n35508), .B(n35507), .Z(n35510) );
  AND U36576 ( .A(x[500]), .B(y[8041]), .Z(n36428) );
  AND U36577 ( .A(x[493]), .B(y[8034]), .Z(n35409) );
  NAND U36578 ( .A(n36428), .B(n35409), .Z(n35413) );
  NAND U36579 ( .A(n35411), .B(n35410), .Z(n35412) );
  NAND U36580 ( .A(n35413), .B(n35412), .Z(n35502) );
  NAND U36581 ( .A(n35415), .B(n35414), .Z(n35419) );
  NAND U36582 ( .A(n35417), .B(n35416), .Z(n35418) );
  AND U36583 ( .A(n35419), .B(n35418), .Z(n35564) );
  AND U36584 ( .A(x[493]), .B(y[8042]), .Z(n35537) );
  AND U36585 ( .A(x[482]), .B(y[8053]), .Z(n35538) );
  XOR U36586 ( .A(n35537), .B(n35538), .Z(n35539) );
  AND U36587 ( .A(x[501]), .B(y[8034]), .Z(n35540) );
  XOR U36588 ( .A(n35539), .B(n35540), .Z(n35562) );
  AND U36589 ( .A(x[492]), .B(y[8043]), .Z(n35485) );
  AND U36590 ( .A(x[481]), .B(y[8054]), .Z(n35486) );
  XOR U36591 ( .A(n35485), .B(n35486), .Z(n35488) );
  AND U36592 ( .A(o[374]), .B(n35420), .Z(n35487) );
  XOR U36593 ( .A(n35488), .B(n35487), .Z(n35561) );
  XOR U36594 ( .A(n35562), .B(n35561), .Z(n35563) );
  XOR U36595 ( .A(n35502), .B(n35501), .Z(n35504) );
  AND U36596 ( .A(x[495]), .B(y[8048]), .Z(n36561) );
  NAND U36597 ( .A(n36561), .B(n35421), .Z(n35425) );
  NANDN U36598 ( .A(n35423), .B(n35422), .Z(n35424) );
  AND U36599 ( .A(n35425), .B(n35424), .Z(n35552) );
  AND U36600 ( .A(x[494]), .B(y[8041]), .Z(n35531) );
  AND U36601 ( .A(x[483]), .B(y[8052]), .Z(n35532) );
  XOR U36602 ( .A(n35531), .B(n35532), .Z(n35533) );
  AND U36603 ( .A(x[484]), .B(y[8051]), .Z(n35534) );
  XOR U36604 ( .A(n35533), .B(n35534), .Z(n35550) );
  AND U36605 ( .A(x[485]), .B(y[8050]), .Z(n35525) );
  AND U36606 ( .A(x[498]), .B(y[8037]), .Z(n35526) );
  XOR U36607 ( .A(n35525), .B(n35526), .Z(n35527) );
  AND U36608 ( .A(x[497]), .B(y[8038]), .Z(n35528) );
  XOR U36609 ( .A(n35527), .B(n35528), .Z(n35549) );
  XOR U36610 ( .A(n35550), .B(n35549), .Z(n35551) );
  XOR U36611 ( .A(n35504), .B(n35503), .Z(n35509) );
  XOR U36612 ( .A(n35510), .B(n35509), .Z(n35573) );
  XOR U36613 ( .A(n35574), .B(n35573), .Z(n35575) );
  XNOR U36614 ( .A(n35576), .B(n35575), .Z(n35462) );
  NAND U36615 ( .A(n35427), .B(n35426), .Z(n35431) );
  NAND U36616 ( .A(n35429), .B(n35428), .Z(n35430) );
  NAND U36617 ( .A(n35431), .B(n35430), .Z(n35582) );
  NAND U36618 ( .A(n35433), .B(n35432), .Z(n35437) );
  NAND U36619 ( .A(n35435), .B(n35434), .Z(n35436) );
  NAND U36620 ( .A(n35437), .B(n35436), .Z(n35580) );
  NAND U36621 ( .A(n35439), .B(n35438), .Z(n35443) );
  NAND U36622 ( .A(n35441), .B(n35440), .Z(n35442) );
  NAND U36623 ( .A(n35443), .B(n35442), .Z(n35579) );
  XOR U36624 ( .A(n35580), .B(n35579), .Z(n35581) );
  XNOR U36625 ( .A(n35582), .B(n35581), .Z(n35461) );
  NANDN U36626 ( .A(n35445), .B(n35444), .Z(n35449) );
  NAND U36627 ( .A(n35447), .B(n35446), .Z(n35448) );
  NAND U36628 ( .A(n35449), .B(n35448), .Z(n35460) );
  XOR U36629 ( .A(n35461), .B(n35460), .Z(n35463) );
  XOR U36630 ( .A(n35462), .B(n35463), .Z(n35598) );
  XOR U36631 ( .A(n35599), .B(n35598), .Z(n35600) );
  XNOR U36632 ( .A(n35601), .B(n35600), .Z(n35594) );
  NAND U36633 ( .A(n35454), .B(n35453), .Z(n35458) );
  NAND U36634 ( .A(n35456), .B(n35455), .Z(n35457) );
  AND U36635 ( .A(n35458), .B(n35457), .Z(n35593) );
  IV U36636 ( .A(n35593), .Z(n35591) );
  XOR U36637 ( .A(n35592), .B(n35591), .Z(n35459) );
  XNOR U36638 ( .A(n35594), .B(n35459), .Z(N760) );
  NAND U36639 ( .A(n35461), .B(n35460), .Z(n35465) );
  NAND U36640 ( .A(n35463), .B(n35462), .Z(n35464) );
  AND U36641 ( .A(n35465), .B(n35464), .Z(n35608) );
  AND U36642 ( .A(x[500]), .B(y[8039]), .Z(n35466) );
  NAND U36643 ( .A(n35644), .B(n35466), .Z(n35470) );
  NAND U36644 ( .A(n35468), .B(n35467), .Z(n35469) );
  NAND U36645 ( .A(n35470), .B(n35469), .Z(n35664) );
  AND U36646 ( .A(x[502]), .B(y[8034]), .Z(n35683) );
  XOR U36647 ( .A(n35684), .B(n35683), .Z(n35686) );
  AND U36648 ( .A(x[482]), .B(y[8054]), .Z(n35685) );
  XOR U36649 ( .A(n35686), .B(n35685), .Z(n35662) );
  AND U36650 ( .A(x[481]), .B(y[8055]), .Z(n35691) );
  XOR U36651 ( .A(n35692), .B(n35691), .Z(n35690) );
  AND U36652 ( .A(o[375]), .B(n35471), .Z(n35689) );
  XOR U36653 ( .A(n35690), .B(n35689), .Z(n35661) );
  XOR U36654 ( .A(n35662), .B(n35661), .Z(n35663) );
  XOR U36655 ( .A(n35664), .B(n35663), .Z(n35722) );
  NAND U36656 ( .A(n35473), .B(n35472), .Z(n35477) );
  NAND U36657 ( .A(n35475), .B(n35474), .Z(n35476) );
  NAND U36658 ( .A(n35477), .B(n35476), .Z(n35658) );
  AND U36659 ( .A(y[8040]), .B(x[496]), .Z(n35479) );
  NAND U36660 ( .A(y[8035]), .B(x[501]), .Z(n35478) );
  XNOR U36661 ( .A(n35479), .B(n35478), .Z(n35645) );
  AND U36662 ( .A(x[485]), .B(y[8051]), .Z(n35646) );
  XOR U36663 ( .A(n35645), .B(n35646), .Z(n35656) );
  AND U36664 ( .A(x[500]), .B(y[8036]), .Z(n35858) );
  AND U36665 ( .A(x[486]), .B(y[8050]), .Z(n35935) );
  XOR U36666 ( .A(n35858), .B(n35935), .Z(n35651) );
  AND U36667 ( .A(x[499]), .B(y[8037]), .Z(n35652) );
  XOR U36668 ( .A(n35651), .B(n35652), .Z(n35655) );
  XOR U36669 ( .A(n35656), .B(n35655), .Z(n35657) );
  XOR U36670 ( .A(n35658), .B(n35657), .Z(n35635) );
  NAND U36671 ( .A(n35784), .B(n35480), .Z(n35484) );
  NANDN U36672 ( .A(n35482), .B(n35481), .Z(n35483) );
  NAND U36673 ( .A(n35484), .B(n35483), .Z(n35633) );
  NAND U36674 ( .A(n35486), .B(n35485), .Z(n35490) );
  NAND U36675 ( .A(n35488), .B(n35487), .Z(n35489) );
  NAND U36676 ( .A(n35490), .B(n35489), .Z(n35632) );
  XOR U36677 ( .A(n35633), .B(n35632), .Z(n35634) );
  XOR U36678 ( .A(n35635), .B(n35634), .Z(n35721) );
  XOR U36679 ( .A(n35722), .B(n35721), .Z(n35724) );
  NAND U36680 ( .A(n35492), .B(n35491), .Z(n35496) );
  NAND U36681 ( .A(n35494), .B(n35493), .Z(n35495) );
  AND U36682 ( .A(n35496), .B(n35495), .Z(n35704) );
  AND U36683 ( .A(x[483]), .B(y[8053]), .Z(n35711) );
  XOR U36684 ( .A(n35712), .B(n35711), .Z(n35710) );
  AND U36685 ( .A(x[484]), .B(y[8052]), .Z(n35709) );
  XOR U36686 ( .A(n35710), .B(n35709), .Z(n35703) );
  AND U36687 ( .A(y[8047]), .B(x[489]), .Z(n35498) );
  NAND U36688 ( .A(y[8046]), .B(x[490]), .Z(n35497) );
  XNOR U36689 ( .A(n35498), .B(n35497), .Z(n35675) );
  AND U36690 ( .A(y[8042]), .B(x[494]), .Z(n35500) );
  NAND U36691 ( .A(y[8048]), .B(x[488]), .Z(n35499) );
  XNOR U36692 ( .A(n35500), .B(n35499), .Z(n35679) );
  NAND U36693 ( .A(x[491]), .B(y[8045]), .Z(n35680) );
  XOR U36694 ( .A(n35675), .B(n35674), .Z(n35705) );
  XOR U36695 ( .A(n35706), .B(n35705), .Z(n35723) );
  XNOR U36696 ( .A(n35724), .B(n35723), .Z(n35734) );
  NAND U36697 ( .A(n35502), .B(n35501), .Z(n35506) );
  NAND U36698 ( .A(n35504), .B(n35503), .Z(n35505) );
  AND U36699 ( .A(n35506), .B(n35505), .Z(n35733) );
  XOR U36700 ( .A(n35734), .B(n35733), .Z(n35735) );
  NAND U36701 ( .A(n35508), .B(n35507), .Z(n35512) );
  NAND U36702 ( .A(n35510), .B(n35509), .Z(n35511) );
  AND U36703 ( .A(n35512), .B(n35511), .Z(n35736) );
  XOR U36704 ( .A(n35735), .B(n35736), .Z(n35742) );
  NAND U36705 ( .A(n35514), .B(n35513), .Z(n35518) );
  NAND U36706 ( .A(n35516), .B(n35515), .Z(n35517) );
  NAND U36707 ( .A(n35518), .B(n35517), .Z(n35730) );
  NAND U36708 ( .A(n35520), .B(n35519), .Z(n35524) );
  NAND U36709 ( .A(n35522), .B(n35521), .Z(n35523) );
  NAND U36710 ( .A(n35524), .B(n35523), .Z(n35728) );
  NAND U36711 ( .A(n35526), .B(n35525), .Z(n35530) );
  NAND U36712 ( .A(n35528), .B(n35527), .Z(n35529) );
  NAND U36713 ( .A(n35530), .B(n35529), .Z(n35641) );
  AND U36714 ( .A(x[480]), .B(y[8056]), .Z(n35715) );
  NAND U36715 ( .A(x[504]), .B(y[8032]), .Z(n35716) );
  NAND U36716 ( .A(x[503]), .B(y[8033]), .Z(n35702) );
  XOR U36717 ( .A(o[376]), .B(n35702), .Z(n35718) );
  AND U36718 ( .A(x[487]), .B(y[8049]), .Z(n35696) );
  AND U36719 ( .A(x[498]), .B(y[8038]), .Z(n35695) );
  XOR U36720 ( .A(n35696), .B(n35695), .Z(n35698) );
  AND U36721 ( .A(x[497]), .B(y[8039]), .Z(n35697) );
  XOR U36722 ( .A(n35698), .B(n35697), .Z(n35638) );
  XOR U36723 ( .A(n35639), .B(n35638), .Z(n35640) );
  XOR U36724 ( .A(n35641), .B(n35640), .Z(n35629) );
  NAND U36725 ( .A(n35532), .B(n35531), .Z(n35536) );
  NAND U36726 ( .A(n35534), .B(n35533), .Z(n35535) );
  NAND U36727 ( .A(n35536), .B(n35535), .Z(n35627) );
  NAND U36728 ( .A(n35538), .B(n35537), .Z(n35542) );
  NAND U36729 ( .A(n35540), .B(n35539), .Z(n35541) );
  NAND U36730 ( .A(n35542), .B(n35541), .Z(n35626) );
  XOR U36731 ( .A(n35627), .B(n35626), .Z(n35628) );
  XOR U36732 ( .A(n35629), .B(n35628), .Z(n35727) );
  XOR U36733 ( .A(n35728), .B(n35727), .Z(n35729) );
  XNOR U36734 ( .A(n35730), .B(n35729), .Z(n35669) );
  NANDN U36735 ( .A(n35544), .B(n35543), .Z(n35548) );
  NAND U36736 ( .A(n35546), .B(n35545), .Z(n35547) );
  AND U36737 ( .A(n35548), .B(n35547), .Z(n35623) );
  NAND U36738 ( .A(n35550), .B(n35549), .Z(n35554) );
  NANDN U36739 ( .A(n35552), .B(n35551), .Z(n35553) );
  AND U36740 ( .A(n35554), .B(n35553), .Z(n35620) );
  NAND U36741 ( .A(n35556), .B(n35555), .Z(n35560) );
  NANDN U36742 ( .A(n35558), .B(n35557), .Z(n35559) );
  AND U36743 ( .A(n35560), .B(n35559), .Z(n35621) );
  XOR U36744 ( .A(n35620), .B(n35621), .Z(n35622) );
  XOR U36745 ( .A(n35623), .B(n35622), .Z(n35667) );
  NAND U36746 ( .A(n35562), .B(n35561), .Z(n35566) );
  NANDN U36747 ( .A(n35564), .B(n35563), .Z(n35565) );
  AND U36748 ( .A(n35566), .B(n35565), .Z(n35668) );
  XOR U36749 ( .A(n35667), .B(n35668), .Z(n35670) );
  XOR U36750 ( .A(n35669), .B(n35670), .Z(n35739) );
  NAND U36751 ( .A(n35568), .B(n35567), .Z(n35572) );
  NAND U36752 ( .A(n35570), .B(n35569), .Z(n35571) );
  AND U36753 ( .A(n35572), .B(n35571), .Z(n35740) );
  XOR U36754 ( .A(n35739), .B(n35740), .Z(n35741) );
  XOR U36755 ( .A(n35742), .B(n35741), .Z(n35606) );
  NAND U36756 ( .A(n35574), .B(n35573), .Z(n35578) );
  NAND U36757 ( .A(n35576), .B(n35575), .Z(n35577) );
  NAND U36758 ( .A(n35578), .B(n35577), .Z(n35617) );
  NAND U36759 ( .A(n35580), .B(n35579), .Z(n35584) );
  NAND U36760 ( .A(n35582), .B(n35581), .Z(n35583) );
  NAND U36761 ( .A(n35584), .B(n35583), .Z(n35615) );
  NAND U36762 ( .A(n35586), .B(n35585), .Z(n35590) );
  NAND U36763 ( .A(n35588), .B(n35587), .Z(n35589) );
  NAND U36764 ( .A(n35590), .B(n35589), .Z(n35614) );
  XOR U36765 ( .A(n35615), .B(n35614), .Z(n35616) );
  XOR U36766 ( .A(n35617), .B(n35616), .Z(n35605) );
  XNOR U36767 ( .A(n35608), .B(n35607), .Z(n35613) );
  NANDN U36768 ( .A(n35591), .B(n35592), .Z(n35597) );
  NOR U36769 ( .A(n35593), .B(n35592), .Z(n35595) );
  OR U36770 ( .A(n35595), .B(n35594), .Z(n35596) );
  AND U36771 ( .A(n35597), .B(n35596), .Z(n35611) );
  NAND U36772 ( .A(n35599), .B(n35598), .Z(n35603) );
  NAND U36773 ( .A(n35601), .B(n35600), .Z(n35602) );
  AND U36774 ( .A(n35603), .B(n35602), .Z(n35612) );
  XOR U36775 ( .A(n35611), .B(n35612), .Z(n35604) );
  XNOR U36776 ( .A(n35613), .B(n35604), .Z(N761) );
  NANDN U36777 ( .A(n35606), .B(n35605), .Z(n35610) );
  NAND U36778 ( .A(n35608), .B(n35607), .Z(n35609) );
  NAND U36779 ( .A(n35610), .B(n35609), .Z(n35753) );
  IV U36780 ( .A(n35753), .Z(n35752) );
  NAND U36781 ( .A(n35615), .B(n35614), .Z(n35619) );
  NAND U36782 ( .A(n35617), .B(n35616), .Z(n35618) );
  AND U36783 ( .A(n35619), .B(n35618), .Z(n35749) );
  NAND U36784 ( .A(n35621), .B(n35620), .Z(n35625) );
  NAND U36785 ( .A(n35623), .B(n35622), .Z(n35624) );
  AND U36786 ( .A(n35625), .B(n35624), .Z(n35766) );
  NAND U36787 ( .A(n35627), .B(n35626), .Z(n35631) );
  NAND U36788 ( .A(n35629), .B(n35628), .Z(n35630) );
  NAND U36789 ( .A(n35631), .B(n35630), .Z(n35772) );
  NAND U36790 ( .A(n35633), .B(n35632), .Z(n35637) );
  NAND U36791 ( .A(n35635), .B(n35634), .Z(n35636) );
  NAND U36792 ( .A(n35637), .B(n35636), .Z(n35771) );
  XOR U36793 ( .A(n35772), .B(n35771), .Z(n35774) );
  NAND U36794 ( .A(n35639), .B(n35638), .Z(n35643) );
  NAND U36795 ( .A(n35641), .B(n35640), .Z(n35642) );
  AND U36796 ( .A(n35643), .B(n35642), .Z(n35804) );
  AND U36797 ( .A(x[501]), .B(y[8040]), .Z(n36656) );
  NAND U36798 ( .A(n36656), .B(n35644), .Z(n35648) );
  NAND U36799 ( .A(n35646), .B(n35645), .Z(n35647) );
  AND U36800 ( .A(n35648), .B(n35647), .Z(n35879) );
  AND U36801 ( .A(x[502]), .B(y[8035]), .Z(n35847) );
  AND U36802 ( .A(x[485]), .B(y[8052]), .Z(n35846) );
  NAND U36803 ( .A(x[497]), .B(y[8040]), .Z(n35845) );
  XOR U36804 ( .A(n35846), .B(n35845), .Z(n35848) );
  XOR U36805 ( .A(n35847), .B(n35848), .Z(n35877) );
  AND U36806 ( .A(y[8037]), .B(x[500]), .Z(n35650) );
  NAND U36807 ( .A(y[8036]), .B(x[501]), .Z(n35649) );
  XNOR U36808 ( .A(n35650), .B(n35649), .Z(n35859) );
  NAND U36809 ( .A(x[499]), .B(y[8038]), .Z(n35860) );
  NAND U36810 ( .A(n35935), .B(n35858), .Z(n35654) );
  NAND U36811 ( .A(n35652), .B(n35651), .Z(n35653) );
  AND U36812 ( .A(n35654), .B(n35653), .Z(n35885) );
  AND U36813 ( .A(x[495]), .B(y[8042]), .Z(n35866) );
  AND U36814 ( .A(x[498]), .B(y[8039]), .Z(n35865) );
  NAND U36815 ( .A(x[486]), .B(y[8051]), .Z(n35864) );
  XOR U36816 ( .A(n35865), .B(n35864), .Z(n35867) );
  XOR U36817 ( .A(n35866), .B(n35867), .Z(n35883) );
  AND U36818 ( .A(x[503]), .B(y[8034]), .Z(n35841) );
  AND U36819 ( .A(x[484]), .B(y[8053]), .Z(n35840) );
  NAND U36820 ( .A(x[496]), .B(y[8041]), .Z(n35839) );
  XOR U36821 ( .A(n35840), .B(n35839), .Z(n35842) );
  XNOR U36822 ( .A(n35841), .B(n35842), .Z(n35882) );
  XOR U36823 ( .A(n35885), .B(n35884), .Z(n35801) );
  XOR U36824 ( .A(n35802), .B(n35801), .Z(n35803) );
  XNOR U36825 ( .A(n35804), .B(n35803), .Z(n35816) );
  NAND U36826 ( .A(n35656), .B(n35655), .Z(n35660) );
  NAND U36827 ( .A(n35658), .B(n35657), .Z(n35659) );
  NAND U36828 ( .A(n35660), .B(n35659), .Z(n35814) );
  NAND U36829 ( .A(n35662), .B(n35661), .Z(n35666) );
  NAND U36830 ( .A(n35664), .B(n35663), .Z(n35665) );
  NAND U36831 ( .A(n35666), .B(n35665), .Z(n35813) );
  XOR U36832 ( .A(n35814), .B(n35813), .Z(n35815) );
  XOR U36833 ( .A(n35816), .B(n35815), .Z(n35773) );
  XNOR U36834 ( .A(n35774), .B(n35773), .Z(n35765) );
  NAND U36835 ( .A(n35668), .B(n35667), .Z(n35672) );
  NAND U36836 ( .A(n35670), .B(n35669), .Z(n35671) );
  NAND U36837 ( .A(n35672), .B(n35671), .Z(n35767) );
  XNOR U36838 ( .A(n35768), .B(n35767), .Z(n35762) );
  NANDN U36839 ( .A(n35783), .B(n35673), .Z(n35677) );
  NAND U36840 ( .A(n35675), .B(n35674), .Z(n35676) );
  NAND U36841 ( .A(n35677), .B(n35676), .Z(n35808) );
  AND U36842 ( .A(x[494]), .B(y[8048]), .Z(n36648) );
  NAND U36843 ( .A(n36648), .B(n35678), .Z(n35682) );
  NANDN U36844 ( .A(n35680), .B(n35679), .Z(n35681) );
  AND U36845 ( .A(n35682), .B(n35681), .Z(n35836) );
  AND U36846 ( .A(x[491]), .B(y[8046]), .Z(n35854) );
  AND U36847 ( .A(x[492]), .B(y[8045]), .Z(n35853) );
  NAND U36848 ( .A(x[487]), .B(y[8050]), .Z(n35852) );
  XOR U36849 ( .A(n35853), .B(n35852), .Z(n35855) );
  XOR U36850 ( .A(n35854), .B(n35855), .Z(n35834) );
  NAND U36851 ( .A(x[504]), .B(y[8033]), .Z(n35851) );
  XNOR U36852 ( .A(o[377]), .B(n35851), .Z(n35821) );
  NAND U36853 ( .A(x[481]), .B(y[8056]), .Z(n35822) );
  NAND U36854 ( .A(x[493]), .B(y[8044]), .Z(n35824) );
  XOR U36855 ( .A(n35808), .B(n35807), .Z(n35810) );
  NAND U36856 ( .A(n35684), .B(n35683), .Z(n35688) );
  AND U36857 ( .A(n35686), .B(n35685), .Z(n35687) );
  ANDN U36858 ( .B(n35688), .A(n35687), .Z(n35796) );
  AND U36859 ( .A(n35690), .B(n35689), .Z(n35694) );
  NAND U36860 ( .A(n35692), .B(n35691), .Z(n35693) );
  NANDN U36861 ( .A(n35694), .B(n35693), .Z(n35795) );
  NAND U36862 ( .A(n35696), .B(n35695), .Z(n35700) );
  NAND U36863 ( .A(n35698), .B(n35697), .Z(n35699) );
  AND U36864 ( .A(n35700), .B(n35699), .Z(n35792) );
  AND U36865 ( .A(x[488]), .B(y[8049]), .Z(n35786) );
  XOR U36866 ( .A(n35784), .B(n35701), .Z(n35785) );
  XOR U36867 ( .A(n35786), .B(n35785), .Z(n35790) );
  ANDN U36868 ( .B(o[376]), .A(n35702), .Z(n35779) );
  AND U36869 ( .A(x[505]), .B(y[8032]), .Z(n35778) );
  NAND U36870 ( .A(x[480]), .B(y[8057]), .Z(n35777) );
  XOR U36871 ( .A(n35778), .B(n35777), .Z(n35780) );
  XNOR U36872 ( .A(n35779), .B(n35780), .Z(n35789) );
  XOR U36873 ( .A(n35790), .B(n35789), .Z(n35791) );
  XOR U36874 ( .A(n35798), .B(n35797), .Z(n35809) );
  XOR U36875 ( .A(n35810), .B(n35809), .Z(n35891) );
  NANDN U36876 ( .A(n35704), .B(n35703), .Z(n35708) );
  NAND U36877 ( .A(n35706), .B(n35705), .Z(n35707) );
  AND U36878 ( .A(n35708), .B(n35707), .Z(n35889) );
  AND U36879 ( .A(n35710), .B(n35709), .Z(n35714) );
  NAND U36880 ( .A(n35712), .B(n35711), .Z(n35713) );
  NANDN U36881 ( .A(n35714), .B(n35713), .Z(n35873) );
  NANDN U36882 ( .A(n35716), .B(n35715), .Z(n35720) );
  NANDN U36883 ( .A(n35718), .B(n35717), .Z(n35719) );
  NAND U36884 ( .A(n35720), .B(n35719), .Z(n35871) );
  AND U36885 ( .A(x[494]), .B(y[8043]), .Z(n35827) );
  NAND U36886 ( .A(x[482]), .B(y[8055]), .Z(n35828) );
  NAND U36887 ( .A(x[483]), .B(y[8054]), .Z(n35830) );
  XOR U36888 ( .A(n35871), .B(n35870), .Z(n35872) );
  XNOR U36889 ( .A(n35873), .B(n35872), .Z(n35888) );
  XOR U36890 ( .A(n35889), .B(n35888), .Z(n35890) );
  NAND U36891 ( .A(n35722), .B(n35721), .Z(n35726) );
  NAND U36892 ( .A(n35724), .B(n35723), .Z(n35725) );
  AND U36893 ( .A(n35726), .B(n35725), .Z(n35895) );
  XOR U36894 ( .A(n35894), .B(n35895), .Z(n35897) );
  NAND U36895 ( .A(n35728), .B(n35727), .Z(n35732) );
  NAND U36896 ( .A(n35730), .B(n35729), .Z(n35731) );
  AND U36897 ( .A(n35732), .B(n35731), .Z(n35896) );
  XNOR U36898 ( .A(n35897), .B(n35896), .Z(n35760) );
  NAND U36899 ( .A(n35734), .B(n35733), .Z(n35738) );
  NAND U36900 ( .A(n35736), .B(n35735), .Z(n35737) );
  AND U36901 ( .A(n35738), .B(n35737), .Z(n35759) );
  XOR U36902 ( .A(n35760), .B(n35759), .Z(n35761) );
  XNOR U36903 ( .A(n35762), .B(n35761), .Z(n35747) );
  NAND U36904 ( .A(n35740), .B(n35739), .Z(n35744) );
  NAND U36905 ( .A(n35742), .B(n35741), .Z(n35743) );
  NAND U36906 ( .A(n35744), .B(n35743), .Z(n35746) );
  XOR U36907 ( .A(n35747), .B(n35746), .Z(n35748) );
  XOR U36908 ( .A(n35749), .B(n35748), .Z(n35755) );
  XNOR U36909 ( .A(n35754), .B(n35755), .Z(n35745) );
  XOR U36910 ( .A(n35752), .B(n35745), .Z(N762) );
  NAND U36911 ( .A(n35747), .B(n35746), .Z(n35751) );
  NAND U36912 ( .A(n35749), .B(n35748), .Z(n35750) );
  NAND U36913 ( .A(n35751), .B(n35750), .Z(n36044) );
  IV U36914 ( .A(n36044), .Z(n36042) );
  OR U36915 ( .A(n35754), .B(n35752), .Z(n35758) );
  ANDN U36916 ( .B(n35754), .A(n35753), .Z(n35756) );
  OR U36917 ( .A(n35756), .B(n35755), .Z(n35757) );
  AND U36918 ( .A(n35758), .B(n35757), .Z(n36043) );
  NAND U36919 ( .A(n35760), .B(n35759), .Z(n35764) );
  NAND U36920 ( .A(n35762), .B(n35761), .Z(n35763) );
  NAND U36921 ( .A(n35764), .B(n35763), .Z(n36037) );
  NANDN U36922 ( .A(n35766), .B(n35765), .Z(n35770) );
  NAND U36923 ( .A(n35768), .B(n35767), .Z(n35769) );
  AND U36924 ( .A(n35770), .B(n35769), .Z(n36036) );
  XOR U36925 ( .A(n36037), .B(n36036), .Z(n36039) );
  NAND U36926 ( .A(n35772), .B(n35771), .Z(n35776) );
  NAND U36927 ( .A(n35774), .B(n35773), .Z(n35775) );
  NAND U36928 ( .A(n35776), .B(n35775), .Z(n36033) );
  AND U36929 ( .A(x[482]), .B(y[8056]), .Z(n36000) );
  XOR U36930 ( .A(n36001), .B(n36000), .Z(n36002) );
  AND U36931 ( .A(x[504]), .B(y[8034]), .Z(n36003) );
  XOR U36932 ( .A(n36002), .B(n36003), .Z(n35965) );
  NANDN U36933 ( .A(n35778), .B(n35777), .Z(n35782) );
  OR U36934 ( .A(n35780), .B(n35779), .Z(n35781) );
  NAND U36935 ( .A(n35782), .B(n35781), .Z(n35966) );
  XNOR U36936 ( .A(n35965), .B(n35966), .Z(n35968) );
  NANDN U36937 ( .A(n35784), .B(n35783), .Z(n35788) );
  NANDN U36938 ( .A(n35786), .B(n35785), .Z(n35787) );
  AND U36939 ( .A(n35788), .B(n35787), .Z(n35967) );
  XOR U36940 ( .A(n35968), .B(n35967), .Z(n35914) );
  NAND U36941 ( .A(n35790), .B(n35789), .Z(n35794) );
  NANDN U36942 ( .A(n35792), .B(n35791), .Z(n35793) );
  AND U36943 ( .A(n35794), .B(n35793), .Z(n35913) );
  NANDN U36944 ( .A(n35796), .B(n35795), .Z(n35800) );
  NAND U36945 ( .A(n35798), .B(n35797), .Z(n35799) );
  NAND U36946 ( .A(n35800), .B(n35799), .Z(n35916) );
  NAND U36947 ( .A(n35802), .B(n35801), .Z(n35806) );
  NAND U36948 ( .A(n35804), .B(n35803), .Z(n35805) );
  NAND U36949 ( .A(n35806), .B(n35805), .Z(n35908) );
  NAND U36950 ( .A(n35808), .B(n35807), .Z(n35812) );
  NAND U36951 ( .A(n35810), .B(n35809), .Z(n35811) );
  AND U36952 ( .A(n35812), .B(n35811), .Z(n35907) );
  XOR U36953 ( .A(n35908), .B(n35907), .Z(n35909) );
  XNOR U36954 ( .A(n35910), .B(n35909), .Z(n36031) );
  NAND U36955 ( .A(n35814), .B(n35813), .Z(n35818) );
  NAND U36956 ( .A(n35816), .B(n35815), .Z(n35817) );
  NAND U36957 ( .A(n35818), .B(n35817), .Z(n35956) );
  AND U36958 ( .A(x[492]), .B(y[8046]), .Z(n36100) );
  AND U36959 ( .A(x[485]), .B(y[8053]), .Z(n35977) );
  XOR U36960 ( .A(n36100), .B(n35977), .Z(n35979) );
  AND U36961 ( .A(x[490]), .B(y[8048]), .Z(n35978) );
  XOR U36962 ( .A(n35979), .B(n35978), .Z(n35922) );
  AND U36963 ( .A(y[8052]), .B(x[486]), .Z(n35820) );
  NAND U36964 ( .A(y[8050]), .B(x[488]), .Z(n35819) );
  XNOR U36965 ( .A(n35820), .B(n35819), .Z(n35937) );
  AND U36966 ( .A(x[489]), .B(y[8049]), .Z(n35936) );
  XOR U36967 ( .A(n35937), .B(n35936), .Z(n35920) );
  AND U36968 ( .A(x[487]), .B(y[8051]), .Z(n35919) );
  XOR U36969 ( .A(n35920), .B(n35919), .Z(n35921) );
  XOR U36970 ( .A(n35922), .B(n35921), .Z(n36027) );
  NANDN U36971 ( .A(n35822), .B(n35821), .Z(n35826) );
  NANDN U36972 ( .A(n35824), .B(n35823), .Z(n35825) );
  AND U36973 ( .A(n35826), .B(n35825), .Z(n36025) );
  NANDN U36974 ( .A(n35828), .B(n35827), .Z(n35832) );
  NANDN U36975 ( .A(n35830), .B(n35829), .Z(n35831) );
  NAND U36976 ( .A(n35832), .B(n35831), .Z(n36024) );
  XOR U36977 ( .A(n36027), .B(n36026), .Z(n35985) );
  NANDN U36978 ( .A(n35834), .B(n35833), .Z(n35838) );
  NANDN U36979 ( .A(n35836), .B(n35835), .Z(n35837) );
  AND U36980 ( .A(n35838), .B(n35837), .Z(n35984) );
  NANDN U36981 ( .A(n35840), .B(n35839), .Z(n35844) );
  OR U36982 ( .A(n35842), .B(n35841), .Z(n35843) );
  AND U36983 ( .A(n35844), .B(n35843), .Z(n35990) );
  NANDN U36984 ( .A(n35846), .B(n35845), .Z(n35850) );
  OR U36985 ( .A(n35848), .B(n35847), .Z(n35849) );
  NAND U36986 ( .A(n35850), .B(n35849), .Z(n35991) );
  XNOR U36987 ( .A(n35990), .B(n35991), .Z(n35993) );
  ANDN U36988 ( .B(o[377]), .A(n35851), .Z(n35930) );
  AND U36989 ( .A(x[494]), .B(y[8044]), .Z(n35929) );
  XOR U36990 ( .A(n35930), .B(n35929), .Z(n35932) );
  AND U36991 ( .A(x[481]), .B(y[8057]), .Z(n35931) );
  XOR U36992 ( .A(n35932), .B(n35931), .Z(n35972) );
  AND U36993 ( .A(x[505]), .B(y[8033]), .Z(n35938) );
  XOR U36994 ( .A(o[378]), .B(n35938), .Z(n35981) );
  AND U36995 ( .A(x[506]), .B(y[8032]), .Z(n35980) );
  XOR U36996 ( .A(n35981), .B(n35980), .Z(n35983) );
  AND U36997 ( .A(x[480]), .B(y[8058]), .Z(n35982) );
  XOR U36998 ( .A(n35983), .B(n35982), .Z(n35971) );
  XOR U36999 ( .A(n35972), .B(n35971), .Z(n35974) );
  NANDN U37000 ( .A(n35853), .B(n35852), .Z(n35857) );
  OR U37001 ( .A(n35855), .B(n35854), .Z(n35856) );
  AND U37002 ( .A(n35857), .B(n35856), .Z(n35973) );
  XOR U37003 ( .A(n35974), .B(n35973), .Z(n35992) );
  XOR U37004 ( .A(n35993), .B(n35992), .Z(n35962) );
  AND U37005 ( .A(x[501]), .B(y[8037]), .Z(n35926) );
  NAND U37006 ( .A(n35926), .B(n35858), .Z(n35862) );
  NANDN U37007 ( .A(n35860), .B(n35859), .Z(n35861) );
  AND U37008 ( .A(n35862), .B(n35861), .Z(n36021) );
  XOR U37009 ( .A(n35926), .B(n35925), .Z(n35928) );
  AND U37010 ( .A(x[500]), .B(y[8038]), .Z(n35927) );
  XOR U37011 ( .A(n35928), .B(n35927), .Z(n36018) );
  NAND U37012 ( .A(x[503]), .B(y[8035]), .Z(n36007) );
  XNOR U37013 ( .A(n36006), .B(n36007), .Z(n36008) );
  NAND U37014 ( .A(x[502]), .B(y[8036]), .Z(n36009) );
  XOR U37015 ( .A(n36008), .B(n36009), .Z(n36019) );
  AND U37016 ( .A(x[484]), .B(y[8054]), .Z(n36012) );
  XOR U37017 ( .A(n36013), .B(n36012), .Z(n36014) );
  XOR U37018 ( .A(n36014), .B(n35863), .Z(n35997) );
  AND U37019 ( .A(x[491]), .B(y[8047]), .Z(n35940) );
  AND U37020 ( .A(x[483]), .B(y[8055]), .Z(n35939) );
  XOR U37021 ( .A(n35940), .B(n35939), .Z(n35942) );
  AND U37022 ( .A(x[499]), .B(y[8039]), .Z(n35941) );
  XOR U37023 ( .A(n35942), .B(n35941), .Z(n35996) );
  XOR U37024 ( .A(n35997), .B(n35996), .Z(n35999) );
  NANDN U37025 ( .A(n35865), .B(n35864), .Z(n35869) );
  OR U37026 ( .A(n35867), .B(n35866), .Z(n35868) );
  AND U37027 ( .A(n35869), .B(n35868), .Z(n35998) );
  XNOR U37028 ( .A(n35999), .B(n35998), .Z(n35959) );
  XOR U37029 ( .A(n35960), .B(n35959), .Z(n35961) );
  XNOR U37030 ( .A(n35987), .B(n35986), .Z(n35954) );
  NAND U37031 ( .A(n35871), .B(n35870), .Z(n35875) );
  NAND U37032 ( .A(n35873), .B(n35872), .Z(n35874) );
  NAND U37033 ( .A(n35875), .B(n35874), .Z(n35949) );
  NANDN U37034 ( .A(n35877), .B(n35876), .Z(n35881) );
  NANDN U37035 ( .A(n35879), .B(n35878), .Z(n35880) );
  NAND U37036 ( .A(n35881), .B(n35880), .Z(n35948) );
  NANDN U37037 ( .A(n35883), .B(n35882), .Z(n35887) );
  NANDN U37038 ( .A(n35885), .B(n35884), .Z(n35886) );
  NAND U37039 ( .A(n35887), .B(n35886), .Z(n35947) );
  XOR U37040 ( .A(n35948), .B(n35947), .Z(n35950) );
  XOR U37041 ( .A(n35949), .B(n35950), .Z(n35953) );
  XOR U37042 ( .A(n35954), .B(n35953), .Z(n35955) );
  XOR U37043 ( .A(n35956), .B(n35955), .Z(n36030) );
  XOR U37044 ( .A(n36031), .B(n36030), .Z(n36032) );
  XOR U37045 ( .A(n36033), .B(n36032), .Z(n35904) );
  NAND U37046 ( .A(n35889), .B(n35888), .Z(n35893) );
  NANDN U37047 ( .A(n35891), .B(n35890), .Z(n35892) );
  AND U37048 ( .A(n35893), .B(n35892), .Z(n35901) );
  NAND U37049 ( .A(n35895), .B(n35894), .Z(n35899) );
  NAND U37050 ( .A(n35897), .B(n35896), .Z(n35898) );
  AND U37051 ( .A(n35899), .B(n35898), .Z(n35902) );
  XOR U37052 ( .A(n35901), .B(n35902), .Z(n35903) );
  XOR U37053 ( .A(n35904), .B(n35903), .Z(n36038) );
  XOR U37054 ( .A(n36039), .B(n36038), .Z(n36045) );
  XNOR U37055 ( .A(n36043), .B(n36045), .Z(n35900) );
  XOR U37056 ( .A(n36042), .B(n35900), .Z(N763) );
  NAND U37057 ( .A(n35902), .B(n35901), .Z(n35906) );
  NAND U37058 ( .A(n35904), .B(n35903), .Z(n35905) );
  AND U37059 ( .A(n35906), .B(n35905), .Z(n36180) );
  NAND U37060 ( .A(n35908), .B(n35907), .Z(n35912) );
  NAND U37061 ( .A(n35910), .B(n35909), .Z(n35911) );
  NAND U37062 ( .A(n35912), .B(n35911), .Z(n36057) );
  NANDN U37063 ( .A(n35914), .B(n35913), .Z(n35918) );
  NANDN U37064 ( .A(n35916), .B(n35915), .Z(n35917) );
  NAND U37065 ( .A(n35918), .B(n35917), .Z(n36063) );
  NAND U37066 ( .A(n35920), .B(n35919), .Z(n35924) );
  NAND U37067 ( .A(n35922), .B(n35921), .Z(n35923) );
  NAND U37068 ( .A(n35924), .B(n35923), .Z(n36164) );
  NAND U37069 ( .A(n35930), .B(n35929), .Z(n35934) );
  NAND U37070 ( .A(n35932), .B(n35931), .Z(n35933) );
  NAND U37071 ( .A(n35934), .B(n35933), .Z(n36114) );
  XOR U37072 ( .A(n36113), .B(n36114), .Z(n36115) );
  AND U37073 ( .A(x[488]), .B(y[8052]), .Z(n36139) );
  AND U37074 ( .A(x[494]), .B(y[8045]), .Z(n36110) );
  AND U37075 ( .A(x[481]), .B(y[8058]), .Z(n36109) );
  XOR U37076 ( .A(n36110), .B(n36109), .Z(n36111) );
  XOR U37077 ( .A(n36112), .B(n36111), .Z(n36081) );
  AND U37078 ( .A(x[497]), .B(y[8042]), .Z(n36141) );
  AND U37079 ( .A(x[484]), .B(y[8055]), .Z(n36140) );
  XOR U37080 ( .A(n36141), .B(n36140), .Z(n36143) );
  AND U37081 ( .A(x[485]), .B(y[8054]), .Z(n36142) );
  XOR U37082 ( .A(n36143), .B(n36142), .Z(n36080) );
  XNOR U37083 ( .A(n36081), .B(n36080), .Z(n36083) );
  XOR U37084 ( .A(n36082), .B(n36083), .Z(n36116) );
  XNOR U37085 ( .A(n36115), .B(n36116), .Z(n36163) );
  NAND U37086 ( .A(n35940), .B(n35939), .Z(n35944) );
  NAND U37087 ( .A(n35942), .B(n35941), .Z(n35943) );
  NAND U37088 ( .A(n35944), .B(n35943), .Z(n36119) );
  AND U37089 ( .A(y[8035]), .B(x[504]), .Z(n35946) );
  NAND U37090 ( .A(y[8039]), .B(x[500]), .Z(n35945) );
  XNOR U37091 ( .A(n35946), .B(n35945), .Z(n36128) );
  AND U37092 ( .A(x[487]), .B(y[8052]), .Z(n36127) );
  XOR U37093 ( .A(n36128), .B(n36127), .Z(n36118) );
  AND U37094 ( .A(x[488]), .B(y[8051]), .Z(n36097) );
  AND U37095 ( .A(x[503]), .B(y[8036]), .Z(n36096) );
  XOR U37096 ( .A(n36097), .B(n36096), .Z(n36099) );
  AND U37097 ( .A(x[502]), .B(y[8037]), .Z(n36098) );
  XOR U37098 ( .A(n36099), .B(n36098), .Z(n36117) );
  XOR U37099 ( .A(n36118), .B(n36117), .Z(n36120) );
  XOR U37100 ( .A(n36119), .B(n36120), .Z(n36162) );
  XOR U37101 ( .A(n36163), .B(n36162), .Z(n36165) );
  XNOR U37102 ( .A(n36164), .B(n36165), .Z(n36062) );
  XOR U37103 ( .A(n36063), .B(n36062), .Z(n36065) );
  NAND U37104 ( .A(n35948), .B(n35947), .Z(n35952) );
  NAND U37105 ( .A(n35950), .B(n35949), .Z(n35951) );
  AND U37106 ( .A(n35952), .B(n35951), .Z(n36064) );
  XOR U37107 ( .A(n36065), .B(n36064), .Z(n36056) );
  XOR U37108 ( .A(n36057), .B(n36056), .Z(n36059) );
  NAND U37109 ( .A(n35954), .B(n35953), .Z(n35958) );
  NAND U37110 ( .A(n35956), .B(n35955), .Z(n35957) );
  AND U37111 ( .A(n35958), .B(n35957), .Z(n36053) );
  NAND U37112 ( .A(n35960), .B(n35959), .Z(n35964) );
  NANDN U37113 ( .A(n35962), .B(n35961), .Z(n35963) );
  AND U37114 ( .A(n35964), .B(n35963), .Z(n36156) );
  NANDN U37115 ( .A(n35966), .B(n35965), .Z(n35970) );
  NAND U37116 ( .A(n35968), .B(n35967), .Z(n35969) );
  NAND U37117 ( .A(n35970), .B(n35969), .Z(n36150) );
  AND U37118 ( .A(x[495]), .B(y[8044]), .Z(n36106) );
  AND U37119 ( .A(x[482]), .B(y[8057]), .Z(n36105) );
  XOR U37120 ( .A(n36106), .B(n36105), .Z(n36108) );
  AND U37121 ( .A(x[483]), .B(y[8056]), .Z(n36107) );
  XOR U37122 ( .A(n36108), .B(n36107), .Z(n36122) );
  AND U37123 ( .A(x[499]), .B(y[8040]), .Z(n36130) );
  AND U37124 ( .A(x[505]), .B(y[8034]), .Z(n36129) );
  XOR U37125 ( .A(n36130), .B(n36129), .Z(n36132) );
  AND U37126 ( .A(x[486]), .B(y[8053]), .Z(n36131) );
  XOR U37127 ( .A(n36132), .B(n36131), .Z(n36121) );
  XOR U37128 ( .A(n36122), .B(n36121), .Z(n36123) );
  NAND U37129 ( .A(x[496]), .B(y[8043]), .Z(n36092) );
  XOR U37130 ( .A(n36092), .B(n36093), .Z(n36095) );
  XOR U37131 ( .A(n36094), .B(n36095), .Z(n36102) );
  AND U37132 ( .A(y[8046]), .B(x[493]), .Z(n35976) );
  AND U37133 ( .A(y[8047]), .B(x[492]), .Z(n35975) );
  XOR U37134 ( .A(n35976), .B(n35975), .Z(n36101) );
  XNOR U37135 ( .A(n36102), .B(n36101), .Z(n36124) );
  XOR U37136 ( .A(n36123), .B(n36124), .Z(n36071) );
  XOR U37137 ( .A(n36069), .B(n36068), .Z(n36070) );
  XOR U37138 ( .A(n36071), .B(n36070), .Z(n36148) );
  XNOR U37139 ( .A(n36149), .B(n36148), .Z(n36151) );
  XOR U37140 ( .A(n36150), .B(n36151), .Z(n36157) );
  NANDN U37141 ( .A(n35985), .B(n35984), .Z(n35989) );
  NAND U37142 ( .A(n35987), .B(n35986), .Z(n35988) );
  AND U37143 ( .A(n35989), .B(n35988), .Z(n36158) );
  XOR U37144 ( .A(n36159), .B(n36158), .Z(n36051) );
  NANDN U37145 ( .A(n35991), .B(n35990), .Z(n35995) );
  NAND U37146 ( .A(n35993), .B(n35992), .Z(n35994) );
  NAND U37147 ( .A(n35995), .B(n35994), .Z(n36154) );
  AND U37148 ( .A(n36001), .B(n36000), .Z(n36005) );
  NAND U37149 ( .A(n36003), .B(n36002), .Z(n36004) );
  NANDN U37150 ( .A(n36005), .B(n36004), .Z(n36075) );
  NANDN U37151 ( .A(n36007), .B(n36006), .Z(n36011) );
  NANDN U37152 ( .A(n36009), .B(n36008), .Z(n36010) );
  NAND U37153 ( .A(n36011), .B(n36010), .Z(n36074) );
  XOR U37154 ( .A(n36075), .B(n36074), .Z(n36076) );
  AND U37155 ( .A(n36013), .B(n36012), .Z(n36017) );
  NANDN U37156 ( .A(n36015), .B(n36014), .Z(n36016) );
  NANDN U37157 ( .A(n36017), .B(n36016), .Z(n36088) );
  AND U37158 ( .A(x[480]), .B(y[8059]), .Z(n36145) );
  AND U37159 ( .A(x[507]), .B(y[8032]), .Z(n36144) );
  XOR U37160 ( .A(n36145), .B(n36144), .Z(n36147) );
  AND U37161 ( .A(x[506]), .B(y[8033]), .Z(n36137) );
  XOR U37162 ( .A(n36137), .B(o[379]), .Z(n36146) );
  XOR U37163 ( .A(n36147), .B(n36146), .Z(n36087) );
  AND U37164 ( .A(x[489]), .B(y[8050]), .Z(n36134) );
  AND U37165 ( .A(x[501]), .B(y[8038]), .Z(n36133) );
  XOR U37166 ( .A(n36134), .B(n36133), .Z(n36136) );
  AND U37167 ( .A(x[498]), .B(y[8041]), .Z(n36135) );
  XOR U37168 ( .A(n36136), .B(n36135), .Z(n36086) );
  XOR U37169 ( .A(n36087), .B(n36086), .Z(n36089) );
  XOR U37170 ( .A(n36088), .B(n36089), .Z(n36077) );
  XOR U37171 ( .A(n36076), .B(n36077), .Z(n36153) );
  XOR U37172 ( .A(n36152), .B(n36153), .Z(n36155) );
  XOR U37173 ( .A(n36154), .B(n36155), .Z(n36171) );
  NANDN U37174 ( .A(n36019), .B(n36018), .Z(n36023) );
  NANDN U37175 ( .A(n36021), .B(n36020), .Z(n36022) );
  AND U37176 ( .A(n36023), .B(n36022), .Z(n36169) );
  NANDN U37177 ( .A(n36025), .B(n36024), .Z(n36029) );
  NAND U37178 ( .A(n36027), .B(n36026), .Z(n36028) );
  AND U37179 ( .A(n36029), .B(n36028), .Z(n36168) );
  XOR U37180 ( .A(n36169), .B(n36168), .Z(n36170) );
  XOR U37181 ( .A(n36053), .B(n36052), .Z(n36058) );
  XNOR U37182 ( .A(n36059), .B(n36058), .Z(n36178) );
  NAND U37183 ( .A(n36031), .B(n36030), .Z(n36035) );
  NAND U37184 ( .A(n36033), .B(n36032), .Z(n36034) );
  NAND U37185 ( .A(n36035), .B(n36034), .Z(n36177) );
  XOR U37186 ( .A(n36178), .B(n36177), .Z(n36179) );
  XOR U37187 ( .A(n36180), .B(n36179), .Z(n36176) );
  NAND U37188 ( .A(n36037), .B(n36036), .Z(n36041) );
  NAND U37189 ( .A(n36039), .B(n36038), .Z(n36040) );
  NAND U37190 ( .A(n36041), .B(n36040), .Z(n36175) );
  NANDN U37191 ( .A(n36042), .B(n36043), .Z(n36048) );
  NOR U37192 ( .A(n36044), .B(n36043), .Z(n36046) );
  OR U37193 ( .A(n36046), .B(n36045), .Z(n36047) );
  AND U37194 ( .A(n36048), .B(n36047), .Z(n36174) );
  XOR U37195 ( .A(n36175), .B(n36174), .Z(n36049) );
  XNOR U37196 ( .A(n36176), .B(n36049), .Z(N764) );
  NANDN U37197 ( .A(n36051), .B(n36050), .Z(n36055) );
  NAND U37198 ( .A(n36053), .B(n36052), .Z(n36054) );
  AND U37199 ( .A(n36055), .B(n36054), .Z(n36311) );
  NAND U37200 ( .A(n36057), .B(n36056), .Z(n36061) );
  NAND U37201 ( .A(n36059), .B(n36058), .Z(n36060) );
  AND U37202 ( .A(n36061), .B(n36060), .Z(n36312) );
  XOR U37203 ( .A(n36311), .B(n36312), .Z(n36314) );
  NAND U37204 ( .A(n36063), .B(n36062), .Z(n36067) );
  NAND U37205 ( .A(n36065), .B(n36064), .Z(n36066) );
  AND U37206 ( .A(n36067), .B(n36066), .Z(n36185) );
  NAND U37207 ( .A(n36069), .B(n36068), .Z(n36073) );
  NAND U37208 ( .A(n36071), .B(n36070), .Z(n36072) );
  NAND U37209 ( .A(n36073), .B(n36072), .Z(n36206) );
  NAND U37210 ( .A(n36075), .B(n36074), .Z(n36079) );
  NAND U37211 ( .A(n36077), .B(n36076), .Z(n36078) );
  NAND U37212 ( .A(n36079), .B(n36078), .Z(n36289) );
  NAND U37213 ( .A(n36081), .B(n36080), .Z(n36085) );
  NANDN U37214 ( .A(n36083), .B(n36082), .Z(n36084) );
  NAND U37215 ( .A(n36085), .B(n36084), .Z(n36288) );
  NAND U37216 ( .A(n36087), .B(n36086), .Z(n36091) );
  NAND U37217 ( .A(n36089), .B(n36088), .Z(n36090) );
  NAND U37218 ( .A(n36091), .B(n36090), .Z(n36287) );
  XOR U37219 ( .A(n36288), .B(n36287), .Z(n36290) );
  XOR U37220 ( .A(n36289), .B(n36290), .Z(n36207) );
  XOR U37221 ( .A(n36206), .B(n36207), .Z(n36209) );
  AND U37222 ( .A(x[487]), .B(y[8053]), .Z(n36242) );
  AND U37223 ( .A(x[492]), .B(y[8048]), .Z(n36241) );
  XOR U37224 ( .A(n36242), .B(n36241), .Z(n36244) );
  AND U37225 ( .A(x[491]), .B(y[8049]), .Z(n36243) );
  XOR U37226 ( .A(n36244), .B(n36243), .Z(n36268) );
  AND U37227 ( .A(x[507]), .B(y[8033]), .Z(n36251) );
  XOR U37228 ( .A(o[380]), .B(n36251), .Z(n36260) );
  AND U37229 ( .A(x[506]), .B(y[8034]), .Z(n36259) );
  XOR U37230 ( .A(n36260), .B(n36259), .Z(n36262) );
  AND U37231 ( .A(x[495]), .B(y[8045]), .Z(n36261) );
  XNOR U37232 ( .A(n36262), .B(n36261), .Z(n36267) );
  XNOR U37233 ( .A(n36268), .B(n36267), .Z(n36270) );
  XOR U37234 ( .A(n36269), .B(n36270), .Z(n36294) );
  AND U37235 ( .A(x[497]), .B(y[8043]), .Z(n36217) );
  AND U37236 ( .A(x[502]), .B(y[8038]), .Z(n36216) );
  XOR U37237 ( .A(n36217), .B(n36216), .Z(n36219) );
  AND U37238 ( .A(x[484]), .B(y[8056]), .Z(n36218) );
  XOR U37239 ( .A(n36219), .B(n36218), .Z(n36272) );
  AND U37240 ( .A(x[486]), .B(y[8054]), .Z(n36403) );
  AND U37241 ( .A(x[499]), .B(y[8041]), .Z(n36252) );
  XOR U37242 ( .A(n36403), .B(n36252), .Z(n36254) );
  XOR U37243 ( .A(n36254), .B(n36253), .Z(n36271) );
  XOR U37244 ( .A(n36272), .B(n36271), .Z(n36274) );
  XOR U37245 ( .A(n36273), .B(n36274), .Z(n36293) );
  NAND U37246 ( .A(n36264), .B(n36100), .Z(n36104) );
  NANDN U37247 ( .A(n36102), .B(n36101), .Z(n36103) );
  NAND U37248 ( .A(n36104), .B(n36103), .Z(n36214) );
  XOR U37249 ( .A(n36212), .B(n36213), .Z(n36215) );
  XOR U37250 ( .A(n36214), .B(n36215), .Z(n36295) );
  XOR U37251 ( .A(n36296), .B(n36295), .Z(n36208) );
  XNOR U37252 ( .A(n36209), .B(n36208), .Z(n36203) );
  NAND U37253 ( .A(n36122), .B(n36121), .Z(n36126) );
  NAND U37254 ( .A(n36124), .B(n36123), .Z(n36125) );
  NAND U37255 ( .A(n36126), .B(n36125), .Z(n36275) );
  XOR U37256 ( .A(n36276), .B(n36275), .Z(n36278) );
  XNOR U37257 ( .A(n36277), .B(n36278), .Z(n36201) );
  AND U37258 ( .A(x[504]), .B(y[8039]), .Z(n36556) );
  AND U37259 ( .A(x[505]), .B(y[8035]), .Z(n36239) );
  XOR U37260 ( .A(n36240), .B(n36239), .Z(n36238) );
  AND U37261 ( .A(x[481]), .B(y[8059]), .Z(n36237) );
  XOR U37262 ( .A(n36238), .B(n36237), .Z(n36308) );
  AND U37263 ( .A(x[496]), .B(y[8044]), .Z(n36234) );
  AND U37264 ( .A(x[504]), .B(y[8036]), .Z(n36233) );
  XOR U37265 ( .A(n36234), .B(n36233), .Z(n36236) );
  AND U37266 ( .A(x[482]), .B(y[8058]), .Z(n36235) );
  XOR U37267 ( .A(n36236), .B(n36235), .Z(n36307) );
  XOR U37268 ( .A(n36308), .B(n36307), .Z(n36310) );
  XOR U37269 ( .A(n36309), .B(n36310), .Z(n36284) );
  AND U37270 ( .A(x[483]), .B(y[8057]), .Z(n36263) );
  XOR U37271 ( .A(n36264), .B(n36263), .Z(n36266) );
  AND U37272 ( .A(x[503]), .B(y[8037]), .Z(n36265) );
  XOR U37273 ( .A(n36266), .B(n36265), .Z(n36304) );
  AND U37274 ( .A(x[485]), .B(y[8055]), .Z(n36248) );
  AND U37275 ( .A(x[501]), .B(y[8039]), .Z(n36247) );
  XOR U37276 ( .A(n36248), .B(n36247), .Z(n36250) );
  AND U37277 ( .A(x[500]), .B(y[8040]), .Z(n36249) );
  XOR U37278 ( .A(n36250), .B(n36249), .Z(n36303) );
  XOR U37279 ( .A(n36304), .B(n36303), .Z(n36306) );
  XOR U37280 ( .A(n36305), .B(n36306), .Z(n36282) );
  AND U37281 ( .A(n36137), .B(o[379]), .Z(n36223) );
  AND U37282 ( .A(x[480]), .B(y[8060]), .Z(n36221) );
  AND U37283 ( .A(x[508]), .B(y[8032]), .Z(n36220) );
  XOR U37284 ( .A(n36221), .B(n36220), .Z(n36222) );
  XOR U37285 ( .A(n36223), .B(n36222), .Z(n36230) );
  NAND U37286 ( .A(y[8050]), .B(x[490]), .Z(n36138) );
  XNOR U37287 ( .A(n36139), .B(n36138), .Z(n36226) );
  AND U37288 ( .A(x[489]), .B(y[8051]), .Z(n36225) );
  XOR U37289 ( .A(n36226), .B(n36225), .Z(n36229) );
  XOR U37290 ( .A(n36230), .B(n36229), .Z(n36232) );
  XOR U37291 ( .A(n36231), .B(n36232), .Z(n36302) );
  XOR U37292 ( .A(n36299), .B(n36300), .Z(n36301) );
  XNOR U37293 ( .A(n36302), .B(n36301), .Z(n36281) );
  XOR U37294 ( .A(n36201), .B(n36200), .Z(n36202) );
  XOR U37295 ( .A(n36203), .B(n36202), .Z(n36198) );
  XNOR U37296 ( .A(n36196), .B(n36197), .Z(n36199) );
  XOR U37297 ( .A(n36198), .B(n36199), .Z(n36184) );
  XOR U37298 ( .A(n36185), .B(n36184), .Z(n36186) );
  NANDN U37299 ( .A(n36157), .B(n36156), .Z(n36161) );
  NAND U37300 ( .A(n36159), .B(n36158), .Z(n36160) );
  NAND U37301 ( .A(n36161), .B(n36160), .Z(n36192) );
  NAND U37302 ( .A(n36163), .B(n36162), .Z(n36167) );
  NAND U37303 ( .A(n36165), .B(n36164), .Z(n36166) );
  NAND U37304 ( .A(n36167), .B(n36166), .Z(n36190) );
  NAND U37305 ( .A(n36169), .B(n36168), .Z(n36173) );
  NANDN U37306 ( .A(n36171), .B(n36170), .Z(n36172) );
  AND U37307 ( .A(n36173), .B(n36172), .Z(n36191) );
  XNOR U37308 ( .A(n36190), .B(n36191), .Z(n36193) );
  XNOR U37309 ( .A(n36186), .B(n36187), .Z(n36313) );
  XOR U37310 ( .A(n36314), .B(n36313), .Z(n36320) );
  NAND U37311 ( .A(n36178), .B(n36177), .Z(n36182) );
  NANDN U37312 ( .A(n36180), .B(n36179), .Z(n36181) );
  AND U37313 ( .A(n36182), .B(n36181), .Z(n36319) );
  IV U37314 ( .A(n36319), .Z(n36317) );
  XOR U37315 ( .A(n36318), .B(n36317), .Z(n36183) );
  XNOR U37316 ( .A(n36320), .B(n36183), .Z(N765) );
  NAND U37317 ( .A(n36185), .B(n36184), .Z(n36189) );
  NANDN U37318 ( .A(n36187), .B(n36186), .Z(n36188) );
  NAND U37319 ( .A(n36189), .B(n36188), .Z(n36330) );
  NAND U37320 ( .A(n36191), .B(n36190), .Z(n36195) );
  NANDN U37321 ( .A(n36193), .B(n36192), .Z(n36194) );
  NAND U37322 ( .A(n36195), .B(n36194), .Z(n36329) );
  NAND U37323 ( .A(n36201), .B(n36200), .Z(n36205) );
  NAND U37324 ( .A(n36203), .B(n36202), .Z(n36204) );
  NAND U37325 ( .A(n36205), .B(n36204), .Z(n36334) );
  XOR U37326 ( .A(n36335), .B(n36334), .Z(n36336) );
  NAND U37327 ( .A(n36207), .B(n36206), .Z(n36211) );
  NAND U37328 ( .A(n36209), .B(n36208), .Z(n36210) );
  NAND U37329 ( .A(n36211), .B(n36210), .Z(n36350) );
  XOR U37330 ( .A(n36469), .B(n36470), .Z(n36471) );
  AND U37331 ( .A(x[490]), .B(y[8052]), .Z(n36483) );
  NAND U37332 ( .A(n36224), .B(n36483), .Z(n36228) );
  NAND U37333 ( .A(n36226), .B(n36225), .Z(n36227) );
  NAND U37334 ( .A(n36228), .B(n36227), .Z(n36459) );
  AND U37335 ( .A(x[492]), .B(y[8049]), .Z(n36613) );
  AND U37336 ( .A(x[481]), .B(y[8060]), .Z(n36423) );
  XOR U37337 ( .A(n36613), .B(n36423), .Z(n36425) );
  AND U37338 ( .A(x[502]), .B(y[8039]), .Z(n36424) );
  XOR U37339 ( .A(n36425), .B(n36424), .Z(n36458) );
  AND U37340 ( .A(x[495]), .B(y[8046]), .Z(n36426) );
  XOR U37341 ( .A(n36656), .B(n36426), .Z(n36427) );
  XOR U37342 ( .A(n36428), .B(n36427), .Z(n36457) );
  XOR U37343 ( .A(n36458), .B(n36457), .Z(n36460) );
  XNOR U37344 ( .A(n36459), .B(n36460), .Z(n36472) );
  XOR U37345 ( .A(n36471), .B(n36472), .Z(n36448) );
  XNOR U37346 ( .A(n36448), .B(n36447), .Z(n36450) );
  XOR U37347 ( .A(n36449), .B(n36450), .Z(n36445) );
  XOR U37348 ( .A(n36464), .B(n36463), .Z(n36465) );
  NAND U37349 ( .A(n36242), .B(n36241), .Z(n36246) );
  NAND U37350 ( .A(n36244), .B(n36243), .Z(n36245) );
  NAND U37351 ( .A(n36246), .B(n36245), .Z(n36364) );
  AND U37352 ( .A(x[503]), .B(y[8038]), .Z(n36394) );
  AND U37353 ( .A(x[493]), .B(y[8048]), .Z(n36392) );
  AND U37354 ( .A(x[504]), .B(y[8037]), .Z(n36538) );
  XOR U37355 ( .A(n36392), .B(n36538), .Z(n36393) );
  XOR U37356 ( .A(n36394), .B(n36393), .Z(n36363) );
  AND U37357 ( .A(x[491]), .B(y[8050]), .Z(n36400) );
  AND U37358 ( .A(x[483]), .B(y[8058]), .Z(n36398) );
  AND U37359 ( .A(x[497]), .B(y[8044]), .Z(n36397) );
  XOR U37360 ( .A(n36398), .B(n36397), .Z(n36399) );
  XOR U37361 ( .A(n36400), .B(n36399), .Z(n36362) );
  XOR U37362 ( .A(n36363), .B(n36362), .Z(n36365) );
  XNOR U37363 ( .A(n36364), .B(n36365), .Z(n36466) );
  AND U37364 ( .A(n36251), .B(o[380]), .Z(n36371) );
  AND U37365 ( .A(x[496]), .B(y[8045]), .Z(n36369) );
  AND U37366 ( .A(x[507]), .B(y[8034]), .Z(n36368) );
  XOR U37367 ( .A(n36369), .B(n36368), .Z(n36370) );
  XOR U37368 ( .A(n36371), .B(n36370), .Z(n36412) );
  AND U37369 ( .A(x[482]), .B(y[8059]), .Z(n36380) );
  XOR U37370 ( .A(n36381), .B(n36380), .Z(n36382) );
  XOR U37371 ( .A(n36383), .B(n36382), .Z(n36411) );
  XOR U37372 ( .A(n36412), .B(n36411), .Z(n36414) );
  XOR U37373 ( .A(n36413), .B(n36414), .Z(n36434) );
  AND U37374 ( .A(x[505]), .B(y[8036]), .Z(n36420) );
  AND U37375 ( .A(x[506]), .B(y[8035]), .Z(n36417) );
  XOR U37376 ( .A(n36418), .B(n36417), .Z(n36419) );
  XOR U37377 ( .A(n36420), .B(n36419), .Z(n36452) );
  IV U37378 ( .A(n36452), .Z(n36255) );
  AND U37379 ( .A(x[508]), .B(y[8033]), .Z(n36431) );
  XOR U37380 ( .A(o[381]), .B(n36431), .Z(n36478) );
  AND U37381 ( .A(x[480]), .B(y[8061]), .Z(n36476) );
  AND U37382 ( .A(x[509]), .B(y[8032]), .Z(n36475) );
  XOR U37383 ( .A(n36476), .B(n36475), .Z(n36477) );
  XNOR U37384 ( .A(n36478), .B(n36477), .Z(n36451) );
  XNOR U37385 ( .A(n36255), .B(n36451), .Z(n36453) );
  XOR U37386 ( .A(n36454), .B(n36453), .Z(n36433) );
  AND U37387 ( .A(y[8055]), .B(x[486]), .Z(n36257) );
  NAND U37388 ( .A(y[8054]), .B(x[487]), .Z(n36256) );
  XNOR U37389 ( .A(n36257), .B(n36256), .Z(n36405) );
  AND U37390 ( .A(x[488]), .B(y[8053]), .Z(n36404) );
  XOR U37391 ( .A(n36405), .B(n36404), .Z(n36473) );
  NAND U37392 ( .A(x[489]), .B(y[8052]), .Z(n36535) );
  AND U37393 ( .A(x[484]), .B(y[8057]), .Z(n36375) );
  AND U37394 ( .A(x[490]), .B(y[8051]), .Z(n36374) );
  XOR U37395 ( .A(n36375), .B(n36374), .Z(n36377) );
  AND U37396 ( .A(x[485]), .B(y[8056]), .Z(n36376) );
  XNOR U37397 ( .A(n36377), .B(n36376), .Z(n36474) );
  XOR U37398 ( .A(n36535), .B(n36474), .Z(n36258) );
  XOR U37399 ( .A(n36473), .B(n36258), .Z(n36388) );
  XOR U37400 ( .A(n36387), .B(n36386), .Z(n36389) );
  XOR U37401 ( .A(n36388), .B(n36389), .Z(n36357) );
  XOR U37402 ( .A(n36357), .B(n36356), .Z(n36359) );
  XOR U37403 ( .A(n36358), .B(n36359), .Z(n36443) );
  XOR U37404 ( .A(n36443), .B(n36444), .Z(n36446) );
  XOR U37405 ( .A(n36445), .B(n36446), .Z(n36351) );
  XOR U37406 ( .A(n36350), .B(n36351), .Z(n36353) );
  NAND U37407 ( .A(n36276), .B(n36275), .Z(n36280) );
  NAND U37408 ( .A(n36278), .B(n36277), .Z(n36279) );
  NAND U37409 ( .A(n36280), .B(n36279), .Z(n36344) );
  NANDN U37410 ( .A(n36282), .B(n36281), .Z(n36286) );
  NANDN U37411 ( .A(n36284), .B(n36283), .Z(n36285) );
  AND U37412 ( .A(n36286), .B(n36285), .Z(n36345) );
  XOR U37413 ( .A(n36344), .B(n36345), .Z(n36347) );
  NAND U37414 ( .A(n36288), .B(n36287), .Z(n36292) );
  NAND U37415 ( .A(n36290), .B(n36289), .Z(n36291) );
  NAND U37416 ( .A(n36292), .B(n36291), .Z(n36340) );
  NANDN U37417 ( .A(n36294), .B(n36293), .Z(n36298) );
  NAND U37418 ( .A(n36296), .B(n36295), .Z(n36297) );
  NAND U37419 ( .A(n36298), .B(n36297), .Z(n36338) );
  XOR U37420 ( .A(n36439), .B(n36440), .Z(n36442) );
  XOR U37421 ( .A(n36441), .B(n36442), .Z(n36339) );
  XOR U37422 ( .A(n36338), .B(n36339), .Z(n36341) );
  XOR U37423 ( .A(n36340), .B(n36341), .Z(n36346) );
  XOR U37424 ( .A(n36347), .B(n36346), .Z(n36352) );
  XOR U37425 ( .A(n36353), .B(n36352), .Z(n36337) );
  XOR U37426 ( .A(n36336), .B(n36337), .Z(n36328) );
  XNOR U37427 ( .A(n36329), .B(n36328), .Z(n36331) );
  XOR U37428 ( .A(n36330), .B(n36331), .Z(n36327) );
  NAND U37429 ( .A(n36312), .B(n36311), .Z(n36316) );
  NAND U37430 ( .A(n36314), .B(n36313), .Z(n36315) );
  NAND U37431 ( .A(n36316), .B(n36315), .Z(n36326) );
  NANDN U37432 ( .A(n36317), .B(n36318), .Z(n36323) );
  NOR U37433 ( .A(n36319), .B(n36318), .Z(n36321) );
  OR U37434 ( .A(n36321), .B(n36320), .Z(n36322) );
  AND U37435 ( .A(n36323), .B(n36322), .Z(n36325) );
  XOR U37436 ( .A(n36326), .B(n36325), .Z(n36324) );
  XNOR U37437 ( .A(n36327), .B(n36324), .Z(N766) );
  NAND U37438 ( .A(n36329), .B(n36328), .Z(n36333) );
  NANDN U37439 ( .A(n36331), .B(n36330), .Z(n36332) );
  NAND U37440 ( .A(n36333), .B(n36332), .Z(n36746) );
  NAND U37441 ( .A(n36339), .B(n36338), .Z(n36343) );
  NAND U37442 ( .A(n36341), .B(n36340), .Z(n36342) );
  AND U37443 ( .A(n36343), .B(n36342), .Z(n36732) );
  NAND U37444 ( .A(n36345), .B(n36344), .Z(n36349) );
  NAND U37445 ( .A(n36347), .B(n36346), .Z(n36348) );
  AND U37446 ( .A(n36349), .B(n36348), .Z(n36734) );
  NAND U37447 ( .A(n36351), .B(n36350), .Z(n36355) );
  NAND U37448 ( .A(n36353), .B(n36352), .Z(n36354) );
  AND U37449 ( .A(n36355), .B(n36354), .Z(n36733) );
  XOR U37450 ( .A(n36734), .B(n36733), .Z(n36731) );
  XOR U37451 ( .A(n36732), .B(n36731), .Z(n36728) );
  NANDN U37452 ( .A(n36357), .B(n36356), .Z(n36361) );
  NANDN U37453 ( .A(n36359), .B(n36358), .Z(n36360) );
  AND U37454 ( .A(n36361), .B(n36360), .Z(n36485) );
  NAND U37455 ( .A(n36363), .B(n36362), .Z(n36367) );
  NAND U37456 ( .A(n36365), .B(n36364), .Z(n36366) );
  AND U37457 ( .A(n36367), .B(n36366), .Z(n36493) );
  NAND U37458 ( .A(n36369), .B(n36368), .Z(n36373) );
  NAND U37459 ( .A(n36371), .B(n36370), .Z(n36372) );
  NAND U37460 ( .A(n36373), .B(n36372), .Z(n36503) );
  NAND U37461 ( .A(n36375), .B(n36374), .Z(n36379) );
  NAND U37462 ( .A(n36377), .B(n36376), .Z(n36378) );
  NAND U37463 ( .A(n36379), .B(n36378), .Z(n36506) );
  AND U37464 ( .A(x[486]), .B(y[8056]), .Z(n36542) );
  AND U37465 ( .A(x[485]), .B(y[8057]), .Z(n36544) );
  AND U37466 ( .A(x[499]), .B(y[8043]), .Z(n36543) );
  XOR U37467 ( .A(n36544), .B(n36543), .Z(n36541) );
  XNOR U37468 ( .A(n36542), .B(n36541), .Z(n36509) );
  AND U37469 ( .A(x[484]), .B(y[8058]), .Z(n36660) );
  AND U37470 ( .A(x[483]), .B(y[8059]), .Z(n36662) );
  AND U37471 ( .A(x[498]), .B(y[8044]), .Z(n36661) );
  XOR U37472 ( .A(n36662), .B(n36661), .Z(n36659) );
  XOR U37473 ( .A(n36660), .B(n36659), .Z(n36512) );
  NAND U37474 ( .A(n36381), .B(n36380), .Z(n36385) );
  NAND U37475 ( .A(n36383), .B(n36382), .Z(n36384) );
  AND U37476 ( .A(n36385), .B(n36384), .Z(n36511) );
  XOR U37477 ( .A(n36509), .B(n36510), .Z(n36505) );
  XOR U37478 ( .A(n36506), .B(n36505), .Z(n36504) );
  XOR U37479 ( .A(n36503), .B(n36504), .Z(n36494) );
  NAND U37480 ( .A(n36387), .B(n36386), .Z(n36391) );
  NAND U37481 ( .A(n36389), .B(n36388), .Z(n36390) );
  AND U37482 ( .A(n36391), .B(n36390), .Z(n36491) );
  XOR U37483 ( .A(n36492), .B(n36491), .Z(n36488) );
  IV U37484 ( .A(n36488), .Z(n36432) );
  NAND U37485 ( .A(n36392), .B(n36538), .Z(n36396) );
  NAND U37486 ( .A(n36394), .B(n36393), .Z(n36395) );
  NAND U37487 ( .A(n36396), .B(n36395), .Z(n36500) );
  NAND U37488 ( .A(n36398), .B(n36397), .Z(n36402) );
  NAND U37489 ( .A(n36400), .B(n36399), .Z(n36401) );
  AND U37490 ( .A(n36402), .B(n36401), .Z(n36522) );
  AND U37491 ( .A(x[480]), .B(y[8062]), .Z(n36550) );
  AND U37492 ( .A(x[509]), .B(y[8033]), .Z(n36555) );
  XOR U37493 ( .A(o[382]), .B(n36555), .Z(n36552) );
  AND U37494 ( .A(x[510]), .B(y[8032]), .Z(n36551) );
  XOR U37495 ( .A(n36552), .B(n36551), .Z(n36549) );
  XOR U37496 ( .A(n36550), .B(n36549), .Z(n36524) );
  AND U37497 ( .A(x[500]), .B(y[8042]), .Z(n36647) );
  XOR U37498 ( .A(n36648), .B(n36647), .Z(n36646) );
  AND U37499 ( .A(x[488]), .B(y[8054]), .Z(n36645) );
  XNOR U37500 ( .A(n36646), .B(n36645), .Z(n36523) );
  XNOR U37501 ( .A(n36522), .B(n36521), .Z(n36499) );
  XOR U37502 ( .A(n36500), .B(n36499), .Z(n36497) );
  AND U37503 ( .A(x[487]), .B(y[8055]), .Z(n36654) );
  NAND U37504 ( .A(n36403), .B(n36654), .Z(n36407) );
  NAND U37505 ( .A(n36405), .B(n36404), .Z(n36406) );
  AND U37506 ( .A(n36407), .B(n36406), .Z(n36515) );
  AND U37507 ( .A(y[8041]), .B(x[501]), .Z(n36409) );
  AND U37508 ( .A(y[8040]), .B(x[502]), .Z(n36408) );
  XOR U37509 ( .A(n36409), .B(n36408), .Z(n36653) );
  XOR U37510 ( .A(n36654), .B(n36653), .Z(n36518) );
  AND U37511 ( .A(x[497]), .B(y[8045]), .Z(n36606) );
  AND U37512 ( .A(x[482]), .B(y[8060]), .Z(n36608) );
  AND U37513 ( .A(x[506]), .B(y[8036]), .Z(n36607) );
  XOR U37514 ( .A(n36608), .B(n36607), .Z(n36605) );
  XNOR U37515 ( .A(n36606), .B(n36605), .Z(n36517) );
  XNOR U37516 ( .A(n36515), .B(n36516), .Z(n36498) );
  IV U37517 ( .A(n36498), .Z(n36410) );
  XOR U37518 ( .A(n36497), .B(n36410), .Z(n36698) );
  NAND U37519 ( .A(n36412), .B(n36411), .Z(n36416) );
  NAND U37520 ( .A(n36414), .B(n36413), .Z(n36415) );
  NAND U37521 ( .A(n36416), .B(n36415), .Z(n36697) );
  XOR U37522 ( .A(n36698), .B(n36697), .Z(n36696) );
  AND U37523 ( .A(n36418), .B(n36417), .Z(n36422) );
  NAND U37524 ( .A(n36420), .B(n36419), .Z(n36421) );
  NANDN U37525 ( .A(n36422), .B(n36421), .Z(n36529) );
  AND U37526 ( .A(x[503]), .B(y[8039]), .Z(n36537) );
  AND U37527 ( .A(y[8038]), .B(x[504]), .Z(n36430) );
  AND U37528 ( .A(y[8037]), .B(x[505]), .Z(n36429) );
  XOR U37529 ( .A(n36430), .B(n36429), .Z(n36536) );
  XOR U37530 ( .A(n36537), .B(n36536), .Z(n36634) );
  AND U37531 ( .A(n36431), .B(o[381]), .Z(n36640) );
  AND U37532 ( .A(x[508]), .B(y[8034]), .Z(n36642) );
  AND U37533 ( .A(x[496]), .B(y[8046]), .Z(n36641) );
  XOR U37534 ( .A(n36642), .B(n36641), .Z(n36639) );
  XNOR U37535 ( .A(n36640), .B(n36639), .Z(n36633) );
  XNOR U37536 ( .A(n36632), .B(n36631), .Z(n36531) );
  XOR U37537 ( .A(n36532), .B(n36531), .Z(n36530) );
  XOR U37538 ( .A(n36529), .B(n36530), .Z(n36695) );
  XOR U37539 ( .A(n36696), .B(n36695), .Z(n36487) );
  XNOR U37540 ( .A(n36432), .B(n36487), .Z(n36486) );
  XOR U37541 ( .A(n36485), .B(n36486), .Z(n36713) );
  NANDN U37542 ( .A(n36434), .B(n36433), .Z(n36438) );
  NANDN U37543 ( .A(n36436), .B(n36435), .Z(n36437) );
  NAND U37544 ( .A(n36438), .B(n36437), .Z(n36715) );
  XOR U37545 ( .A(n36715), .B(n36716), .Z(n36714) );
  XOR U37546 ( .A(n36713), .B(n36714), .Z(n36708) );
  NANDN U37547 ( .A(n36452), .B(n36451), .Z(n36456) );
  OR U37548 ( .A(n36454), .B(n36453), .Z(n36455) );
  NAND U37549 ( .A(n36456), .B(n36455), .Z(n36677) );
  NAND U37550 ( .A(n36458), .B(n36457), .Z(n36462) );
  NAND U37551 ( .A(n36460), .B(n36459), .Z(n36461) );
  AND U37552 ( .A(n36462), .B(n36461), .Z(n36680) );
  NAND U37553 ( .A(n36464), .B(n36463), .Z(n36468) );
  NANDN U37554 ( .A(n36466), .B(n36465), .Z(n36467) );
  AND U37555 ( .A(n36468), .B(n36467), .Z(n36679) );
  XOR U37556 ( .A(n36680), .B(n36679), .Z(n36678) );
  XOR U37557 ( .A(n36677), .B(n36678), .Z(n36692) );
  NAND U37558 ( .A(n36476), .B(n36475), .Z(n36480) );
  NAND U37559 ( .A(n36478), .B(n36477), .Z(n36479) );
  NAND U37560 ( .A(n36480), .B(n36479), .Z(n36625) );
  AND U37561 ( .A(x[507]), .B(y[8035]), .Z(n36618) );
  AND U37562 ( .A(x[481]), .B(y[8061]), .Z(n36617) );
  XOR U37563 ( .A(n36618), .B(n36617), .Z(n36615) );
  XOR U37564 ( .A(n36616), .B(n36615), .Z(n36627) );
  AND U37565 ( .A(y[8050]), .B(x[492]), .Z(n36481) );
  XOR U37566 ( .A(n36482), .B(n36481), .Z(n36611) );
  XOR U37567 ( .A(n36612), .B(n36611), .Z(n36534) );
  AND U37568 ( .A(x[489]), .B(y[8053]), .Z(n36484) );
  XOR U37569 ( .A(n36484), .B(n36483), .Z(n36533) );
  XOR U37570 ( .A(n36534), .B(n36533), .Z(n36628) );
  XOR U37571 ( .A(n36625), .B(n36626), .Z(n36673) );
  XOR U37572 ( .A(n36674), .B(n36673), .Z(n36672) );
  XNOR U37573 ( .A(n36671), .B(n36672), .Z(n36691) );
  XNOR U37574 ( .A(n36689), .B(n36690), .Z(n36710) );
  XOR U37575 ( .A(n36709), .B(n36710), .Z(n36707) );
  XNOR U37576 ( .A(n36708), .B(n36707), .Z(n36727) );
  XNOR U37577 ( .A(n36726), .B(n36725), .Z(n36743) );
  XNOR U37578 ( .A(n36744), .B(n36743), .Z(N767) );
  NANDN U37579 ( .A(n36486), .B(n36485), .Z(n36490) );
  NANDN U37580 ( .A(n36488), .B(n36487), .Z(n36489) );
  AND U37581 ( .A(n36490), .B(n36489), .Z(n36742) );
  NAND U37582 ( .A(n36492), .B(n36491), .Z(n36496) );
  NANDN U37583 ( .A(n36494), .B(n36493), .Z(n36495) );
  AND U37584 ( .A(n36496), .B(n36495), .Z(n36724) );
  NANDN U37585 ( .A(n36498), .B(n36497), .Z(n36502) );
  NAND U37586 ( .A(n36500), .B(n36499), .Z(n36501) );
  AND U37587 ( .A(n36502), .B(n36501), .Z(n36706) );
  NAND U37588 ( .A(n36504), .B(n36503), .Z(n36508) );
  NAND U37589 ( .A(n36506), .B(n36505), .Z(n36507) );
  AND U37590 ( .A(n36508), .B(n36507), .Z(n36688) );
  NANDN U37591 ( .A(n36510), .B(n36509), .Z(n36514) );
  NANDN U37592 ( .A(n36512), .B(n36511), .Z(n36513) );
  AND U37593 ( .A(n36514), .B(n36513), .Z(n36670) );
  NANDN U37594 ( .A(n36516), .B(n36515), .Z(n36520) );
  NANDN U37595 ( .A(n36518), .B(n36517), .Z(n36519) );
  AND U37596 ( .A(n36520), .B(n36519), .Z(n36528) );
  NAND U37597 ( .A(n36522), .B(n36521), .Z(n36526) );
  NANDN U37598 ( .A(n36524), .B(n36523), .Z(n36525) );
  NAND U37599 ( .A(n36526), .B(n36525), .Z(n36527) );
  XNOR U37600 ( .A(n36528), .B(n36527), .Z(n36668) );
  AND U37601 ( .A(x[490]), .B(y[8053]), .Z(n36569) );
  NAND U37602 ( .A(n36537), .B(n36536), .Z(n36540) );
  AND U37603 ( .A(x[505]), .B(y[8038]), .Z(n36574) );
  NAND U37604 ( .A(n36538), .B(n36574), .Z(n36539) );
  AND U37605 ( .A(n36540), .B(n36539), .Z(n36548) );
  NAND U37606 ( .A(n36542), .B(n36541), .Z(n36546) );
  NAND U37607 ( .A(n36544), .B(n36543), .Z(n36545) );
  NAND U37608 ( .A(n36546), .B(n36545), .Z(n36547) );
  NAND U37609 ( .A(n36550), .B(n36549), .Z(n36554) );
  NAND U37610 ( .A(n36552), .B(n36551), .Z(n36553) );
  AND U37611 ( .A(n36554), .B(n36553), .Z(n36604) );
  AND U37612 ( .A(n36555), .B(o[382]), .Z(n36560) );
  AND U37613 ( .A(y[8042]), .B(x[501]), .Z(n36558) );
  XNOR U37614 ( .A(n36556), .B(o[383]), .Z(n36557) );
  XNOR U37615 ( .A(n36558), .B(n36557), .Z(n36559) );
  XOR U37616 ( .A(n36560), .B(n36559), .Z(n36563) );
  XNOR U37617 ( .A(n36561), .B(n36614), .Z(n36562) );
  XNOR U37618 ( .A(n36563), .B(n36562), .Z(n36602) );
  AND U37619 ( .A(y[8052]), .B(x[491]), .Z(n36565) );
  NAND U37620 ( .A(y[8051]), .B(x[492]), .Z(n36564) );
  XNOR U37621 ( .A(n36565), .B(n36564), .Z(n36573) );
  AND U37622 ( .A(y[8037]), .B(x[506]), .Z(n36571) );
  AND U37623 ( .A(y[8032]), .B(x[511]), .Z(n36567) );
  NAND U37624 ( .A(y[8045]), .B(x[498]), .Z(n36566) );
  XNOR U37625 ( .A(n36567), .B(n36566), .Z(n36568) );
  XNOR U37626 ( .A(n36569), .B(n36568), .Z(n36570) );
  XNOR U37627 ( .A(n36571), .B(n36570), .Z(n36572) );
  XOR U37628 ( .A(n36573), .B(n36572), .Z(n36576) );
  AND U37629 ( .A(x[502]), .B(y[8041]), .Z(n36655) );
  XNOR U37630 ( .A(n36655), .B(n36574), .Z(n36575) );
  XNOR U37631 ( .A(n36576), .B(n36575), .Z(n36592) );
  AND U37632 ( .A(y[8061]), .B(x[482]), .Z(n36578) );
  NAND U37633 ( .A(y[8046]), .B(x[497]), .Z(n36577) );
  XNOR U37634 ( .A(n36578), .B(n36577), .Z(n36582) );
  AND U37635 ( .A(y[8047]), .B(x[496]), .Z(n36580) );
  NAND U37636 ( .A(y[8043]), .B(x[500]), .Z(n36579) );
  XNOR U37637 ( .A(n36580), .B(n36579), .Z(n36581) );
  XOR U37638 ( .A(n36582), .B(n36581), .Z(n36590) );
  AND U37639 ( .A(y[8058]), .B(x[485]), .Z(n36584) );
  NAND U37640 ( .A(y[8059]), .B(x[484]), .Z(n36583) );
  XNOR U37641 ( .A(n36584), .B(n36583), .Z(n36588) );
  AND U37642 ( .A(y[8036]), .B(x[507]), .Z(n36586) );
  NAND U37643 ( .A(y[8040]), .B(x[503]), .Z(n36585) );
  XNOR U37644 ( .A(n36586), .B(n36585), .Z(n36587) );
  XNOR U37645 ( .A(n36588), .B(n36587), .Z(n36589) );
  XNOR U37646 ( .A(n36590), .B(n36589), .Z(n36591) );
  XOR U37647 ( .A(n36592), .B(n36591), .Z(n36600) );
  AND U37648 ( .A(y[8044]), .B(x[499]), .Z(n36594) );
  NAND U37649 ( .A(y[8055]), .B(x[488]), .Z(n36593) );
  XNOR U37650 ( .A(n36594), .B(n36593), .Z(n36598) );
  AND U37651 ( .A(y[8056]), .B(x[487]), .Z(n36596) );
  NAND U37652 ( .A(y[8060]), .B(x[483]), .Z(n36595) );
  XNOR U37653 ( .A(n36596), .B(n36595), .Z(n36597) );
  XNOR U37654 ( .A(n36598), .B(n36597), .Z(n36599) );
  XNOR U37655 ( .A(n36600), .B(n36599), .Z(n36601) );
  XNOR U37656 ( .A(n36602), .B(n36601), .Z(n36603) );
  NAND U37657 ( .A(n36606), .B(n36605), .Z(n36610) );
  NAND U37658 ( .A(n36608), .B(n36607), .Z(n36609) );
  AND U37659 ( .A(n36610), .B(n36609), .Z(n36624) );
  AND U37660 ( .A(y[8035]), .B(x[508]), .Z(n36620) );
  NAND U37661 ( .A(y[8063]), .B(x[480]), .Z(n36619) );
  AND U37662 ( .A(y[8057]), .B(x[486]), .Z(n36622) );
  NAND U37663 ( .A(y[8062]), .B(x[481]), .Z(n36621) );
  NANDN U37664 ( .A(n36626), .B(n36625), .Z(n36630) );
  NAND U37665 ( .A(n36628), .B(n36627), .Z(n36629) );
  AND U37666 ( .A(n36630), .B(n36629), .Z(n36638) );
  NAND U37667 ( .A(n36632), .B(n36631), .Z(n36636) );
  NANDN U37668 ( .A(n36634), .B(n36633), .Z(n36635) );
  NAND U37669 ( .A(n36636), .B(n36635), .Z(n36637) );
  NAND U37670 ( .A(n36640), .B(n36639), .Z(n36644) );
  NAND U37671 ( .A(n36642), .B(n36641), .Z(n36643) );
  AND U37672 ( .A(n36644), .B(n36643), .Z(n36652) );
  NAND U37673 ( .A(n36646), .B(n36645), .Z(n36650) );
  NAND U37674 ( .A(n36648), .B(n36647), .Z(n36649) );
  NAND U37675 ( .A(n36650), .B(n36649), .Z(n36651) );
  NAND U37676 ( .A(n36654), .B(n36653), .Z(n36658) );
  NAND U37677 ( .A(n36656), .B(n36655), .Z(n36657) );
  AND U37678 ( .A(n36658), .B(n36657), .Z(n36666) );
  NAND U37679 ( .A(n36660), .B(n36659), .Z(n36664) );
  NAND U37680 ( .A(n36662), .B(n36661), .Z(n36663) );
  NAND U37681 ( .A(n36664), .B(n36663), .Z(n36665) );
  XNOR U37682 ( .A(n36668), .B(n36667), .Z(n36669) );
  XNOR U37683 ( .A(n36670), .B(n36669), .Z(n36686) );
  NAND U37684 ( .A(n36672), .B(n36671), .Z(n36676) );
  NAND U37685 ( .A(n36674), .B(n36673), .Z(n36675) );
  AND U37686 ( .A(n36676), .B(n36675), .Z(n36684) );
  NAND U37687 ( .A(n36680), .B(n36679), .Z(n36681) );
  NAND U37688 ( .A(n36682), .B(n36681), .Z(n36683) );
  XNOR U37689 ( .A(n36684), .B(n36683), .Z(n36685) );
  XNOR U37690 ( .A(n36686), .B(n36685), .Z(n36687) );
  XNOR U37691 ( .A(n36688), .B(n36687), .Z(n36704) );
  NANDN U37692 ( .A(n36690), .B(n36689), .Z(n36694) );
  NANDN U37693 ( .A(n36692), .B(n36691), .Z(n36693) );
  AND U37694 ( .A(n36694), .B(n36693), .Z(n36702) );
  NAND U37695 ( .A(n36696), .B(n36695), .Z(n36700) );
  NAND U37696 ( .A(n36698), .B(n36697), .Z(n36699) );
  NAND U37697 ( .A(n36700), .B(n36699), .Z(n36701) );
  XNOR U37698 ( .A(n36702), .B(n36701), .Z(n36703) );
  XNOR U37699 ( .A(n36704), .B(n36703), .Z(n36705) );
  XNOR U37700 ( .A(n36706), .B(n36705), .Z(n36722) );
  NANDN U37701 ( .A(n36708), .B(n36707), .Z(n36712) );
  NAND U37702 ( .A(n36710), .B(n36709), .Z(n36711) );
  AND U37703 ( .A(n36712), .B(n36711), .Z(n36720) );
  NAND U37704 ( .A(n36714), .B(n36713), .Z(n36718) );
  NAND U37705 ( .A(n36716), .B(n36715), .Z(n36717) );
  NAND U37706 ( .A(n36718), .B(n36717), .Z(n36719) );
  XNOR U37707 ( .A(n36720), .B(n36719), .Z(n36721) );
  XNOR U37708 ( .A(n36722), .B(n36721), .Z(n36723) );
  XNOR U37709 ( .A(n36724), .B(n36723), .Z(n36740) );
  NAND U37710 ( .A(n36726), .B(n36725), .Z(n36730) );
  NANDN U37711 ( .A(n36728), .B(n36727), .Z(n36729) );
  AND U37712 ( .A(n36730), .B(n36729), .Z(n36738) );
  NAND U37713 ( .A(n36732), .B(n36731), .Z(n36736) );
  NAND U37714 ( .A(n36734), .B(n36733), .Z(n36735) );
  NAND U37715 ( .A(n36736), .B(n36735), .Z(n36737) );
  XNOR U37716 ( .A(n36738), .B(n36737), .Z(n36739) );
  XNOR U37717 ( .A(n36740), .B(n36739), .Z(n36741) );
  XNOR U37718 ( .A(n36742), .B(n36741), .Z(n36750) );
  NAND U37719 ( .A(n36744), .B(n36743), .Z(n36748) );
  NANDN U37720 ( .A(n36746), .B(n36745), .Z(n36747) );
  NAND U37721 ( .A(n36748), .B(n36747), .Z(n36749) );
  XNOR U37722 ( .A(n36750), .B(n36749), .Z(N768) );
  AND U37723 ( .A(x[480]), .B(y[8064]), .Z(n37397) );
  XOR U37724 ( .A(n37397), .B(o[384]), .Z(N801) );
  AND U37725 ( .A(x[481]), .B(y[8064]), .Z(n36759) );
  AND U37726 ( .A(x[480]), .B(y[8065]), .Z(n36758) );
  XNOR U37727 ( .A(n36758), .B(o[385]), .Z(n36751) );
  XNOR U37728 ( .A(n36759), .B(n36751), .Z(n36753) );
  NAND U37729 ( .A(n37397), .B(o[384]), .Z(n36752) );
  XNOR U37730 ( .A(n36753), .B(n36752), .Z(N802) );
  NANDN U37731 ( .A(n36759), .B(n36751), .Z(n36755) );
  NAND U37732 ( .A(n36753), .B(n36752), .Z(n36754) );
  AND U37733 ( .A(n36755), .B(n36754), .Z(n36765) );
  AND U37734 ( .A(x[480]), .B(y[8066]), .Z(n36772) );
  XNOR U37735 ( .A(n36772), .B(o[386]), .Z(n36764) );
  XNOR U37736 ( .A(n36765), .B(n36764), .Z(n36767) );
  AND U37737 ( .A(y[8064]), .B(x[482]), .Z(n36757) );
  NAND U37738 ( .A(y[8065]), .B(x[481]), .Z(n36756) );
  XNOR U37739 ( .A(n36757), .B(n36756), .Z(n36761) );
  AND U37740 ( .A(n36758), .B(o[385]), .Z(n36760) );
  XNOR U37741 ( .A(n36761), .B(n36760), .Z(n36766) );
  XNOR U37742 ( .A(n36767), .B(n36766), .Z(N803) );
  AND U37743 ( .A(x[482]), .B(y[8065]), .Z(n36779) );
  NAND U37744 ( .A(n36779), .B(n36759), .Z(n36763) );
  NAND U37745 ( .A(n36761), .B(n36760), .Z(n36762) );
  AND U37746 ( .A(n36763), .B(n36762), .Z(n36785) );
  NANDN U37747 ( .A(n36765), .B(n36764), .Z(n36769) );
  NAND U37748 ( .A(n36767), .B(n36766), .Z(n36768) );
  AND U37749 ( .A(n36769), .B(n36768), .Z(n36784) );
  XNOR U37750 ( .A(n36785), .B(n36784), .Z(n36787) );
  AND U37751 ( .A(x[481]), .B(y[8066]), .Z(n36881) );
  XOR U37752 ( .A(o[387]), .B(n36779), .Z(n36781) );
  XOR U37753 ( .A(n36881), .B(n36781), .Z(n36783) );
  AND U37754 ( .A(y[8064]), .B(x[483]), .Z(n36771) );
  NAND U37755 ( .A(y[8067]), .B(x[480]), .Z(n36770) );
  XNOR U37756 ( .A(n36771), .B(n36770), .Z(n36774) );
  AND U37757 ( .A(n36772), .B(o[386]), .Z(n36773) );
  XOR U37758 ( .A(n36774), .B(n36773), .Z(n36782) );
  XOR U37759 ( .A(n36783), .B(n36782), .Z(n36786) );
  XOR U37760 ( .A(n36787), .B(n36786), .Z(N804) );
  AND U37761 ( .A(x[483]), .B(y[8067]), .Z(n36829) );
  NAND U37762 ( .A(n37397), .B(n36829), .Z(n36776) );
  NAND U37763 ( .A(n36774), .B(n36773), .Z(n36775) );
  NAND U37764 ( .A(n36776), .B(n36775), .Z(n36807) );
  AND U37765 ( .A(y[8068]), .B(x[480]), .Z(n36778) );
  NAND U37766 ( .A(y[8064]), .B(x[484]), .Z(n36777) );
  XNOR U37767 ( .A(n36778), .B(n36777), .Z(n36802) );
  AND U37768 ( .A(n36779), .B(o[387]), .Z(n36801) );
  XOR U37769 ( .A(n36802), .B(n36801), .Z(n36806) );
  AND U37770 ( .A(y[8066]), .B(x[482]), .Z(n36929) );
  NAND U37771 ( .A(y[8067]), .B(x[481]), .Z(n36780) );
  XNOR U37772 ( .A(n36929), .B(n36780), .Z(n36798) );
  AND U37773 ( .A(x[483]), .B(y[8065]), .Z(n36793) );
  XOR U37774 ( .A(n36793), .B(o[388]), .Z(n36797) );
  XOR U37775 ( .A(n36798), .B(n36797), .Z(n36805) );
  XOR U37776 ( .A(n36806), .B(n36805), .Z(n36808) );
  XNOR U37777 ( .A(n36807), .B(n36808), .Z(n36813) );
  NANDN U37778 ( .A(n36785), .B(n36784), .Z(n36789) );
  NAND U37779 ( .A(n36787), .B(n36786), .Z(n36788) );
  NAND U37780 ( .A(n36789), .B(n36788), .Z(n36812) );
  XOR U37781 ( .A(n36811), .B(n36812), .Z(n36790) );
  XNOR U37782 ( .A(n36813), .B(n36790), .Z(N805) );
  AND U37783 ( .A(y[8064]), .B(x[485]), .Z(n36792) );
  NAND U37784 ( .A(y[8069]), .B(x[480]), .Z(n36791) );
  XNOR U37785 ( .A(n36792), .B(n36791), .Z(n36822) );
  AND U37786 ( .A(n36793), .B(o[388]), .Z(n36821) );
  XOR U37787 ( .A(n36822), .B(n36821), .Z(n36820) );
  NAND U37788 ( .A(x[482]), .B(y[8067]), .Z(n36889) );
  AND U37789 ( .A(y[8066]), .B(x[483]), .Z(n36795) );
  NAND U37790 ( .A(y[8068]), .B(x[481]), .Z(n36794) );
  XNOR U37791 ( .A(n36795), .B(n36794), .Z(n36816) );
  AND U37792 ( .A(x[484]), .B(y[8065]), .Z(n36827) );
  XOR U37793 ( .A(n36827), .B(o[389]), .Z(n36815) );
  XOR U37794 ( .A(n36816), .B(n36815), .Z(n36819) );
  XOR U37795 ( .A(n36889), .B(n36819), .Z(n36796) );
  XNOR U37796 ( .A(n36820), .B(n36796), .Z(n36836) );
  NANDN U37797 ( .A(n36889), .B(n36881), .Z(n36800) );
  NAND U37798 ( .A(n36798), .B(n36797), .Z(n36799) );
  NAND U37799 ( .A(n36800), .B(n36799), .Z(n36835) );
  AND U37800 ( .A(x[484]), .B(y[8068]), .Z(n37595) );
  NAND U37801 ( .A(n37595), .B(n37397), .Z(n36804) );
  NAND U37802 ( .A(n36802), .B(n36801), .Z(n36803) );
  NAND U37803 ( .A(n36804), .B(n36803), .Z(n36834) );
  XNOR U37804 ( .A(n36835), .B(n36834), .Z(n36837) );
  NAND U37805 ( .A(n36806), .B(n36805), .Z(n36810) );
  NAND U37806 ( .A(n36808), .B(n36807), .Z(n36809) );
  AND U37807 ( .A(n36810), .B(n36809), .Z(n36832) );
  XNOR U37808 ( .A(n36832), .B(n36831), .Z(n36814) );
  XNOR U37809 ( .A(n36833), .B(n36814), .Z(N806) );
  AND U37810 ( .A(x[483]), .B(y[8068]), .Z(n36890) );
  NAND U37811 ( .A(n36890), .B(n36881), .Z(n36818) );
  NAND U37812 ( .A(n36816), .B(n36815), .Z(n36817) );
  NAND U37813 ( .A(n36818), .B(n36817), .Z(n36866) );
  XOR U37814 ( .A(n36866), .B(n36865), .Z(n36868) );
  AND U37815 ( .A(x[485]), .B(y[8069]), .Z(n37064) );
  NAND U37816 ( .A(n37397), .B(n37064), .Z(n36824) );
  NAND U37817 ( .A(n36822), .B(n36821), .Z(n36823) );
  NAND U37818 ( .A(n36824), .B(n36823), .Z(n36841) );
  AND U37819 ( .A(y[8064]), .B(x[486]), .Z(n36826) );
  NAND U37820 ( .A(y[8070]), .B(x[480]), .Z(n36825) );
  XNOR U37821 ( .A(n36826), .B(n36825), .Z(n36848) );
  AND U37822 ( .A(n36827), .B(o[389]), .Z(n36849) );
  XOR U37823 ( .A(n36848), .B(n36849), .Z(n36842) );
  XOR U37824 ( .A(n36841), .B(n36842), .Z(n36844) );
  NAND U37825 ( .A(y[8068]), .B(x[482]), .Z(n36828) );
  XNOR U37826 ( .A(n36829), .B(n36828), .Z(n36853) );
  AND U37827 ( .A(y[8069]), .B(x[481]), .Z(n37111) );
  NAND U37828 ( .A(y[8066]), .B(x[484]), .Z(n36830) );
  XNOR U37829 ( .A(n37111), .B(n36830), .Z(n36857) );
  AND U37830 ( .A(x[485]), .B(y[8065]), .Z(n36864) );
  XOR U37831 ( .A(o[390]), .B(n36864), .Z(n36856) );
  XOR U37832 ( .A(n36857), .B(n36856), .Z(n36852) );
  XOR U37833 ( .A(n36853), .B(n36852), .Z(n36843) );
  XOR U37834 ( .A(n36844), .B(n36843), .Z(n36867) );
  XOR U37835 ( .A(n36868), .B(n36867), .Z(n36873) );
  NAND U37836 ( .A(n36835), .B(n36834), .Z(n36839) );
  NANDN U37837 ( .A(n36837), .B(n36836), .Z(n36838) );
  AND U37838 ( .A(n36839), .B(n36838), .Z(n36871) );
  XOR U37839 ( .A(n36872), .B(n36871), .Z(n36840) );
  XNOR U37840 ( .A(n36873), .B(n36840), .Z(N807) );
  NAND U37841 ( .A(n36842), .B(n36841), .Z(n36846) );
  NAND U37842 ( .A(n36844), .B(n36843), .Z(n36845) );
  AND U37843 ( .A(n36846), .B(n36845), .Z(n36912) );
  AND U37844 ( .A(y[8066]), .B(x[485]), .Z(n36972) );
  NAND U37845 ( .A(y[8070]), .B(x[481]), .Z(n36847) );
  XNOR U37846 ( .A(n36972), .B(n36847), .Z(n36883) );
  AND U37847 ( .A(x[486]), .B(y[8065]), .Z(n36886) );
  XOR U37848 ( .A(o[391]), .B(n36886), .Z(n36882) );
  XNOR U37849 ( .A(n36883), .B(n36882), .Z(n36901) );
  AND U37850 ( .A(x[486]), .B(y[8070]), .Z(n37131) );
  NAND U37851 ( .A(n37397), .B(n37131), .Z(n36851) );
  NAND U37852 ( .A(n36849), .B(n36848), .Z(n36850) );
  AND U37853 ( .A(n36851), .B(n36850), .Z(n36900) );
  XOR U37854 ( .A(n36901), .B(n36900), .Z(n36902) );
  NANDN U37855 ( .A(n36889), .B(n36890), .Z(n36855) );
  NAND U37856 ( .A(n36853), .B(n36852), .Z(n36854) );
  AND U37857 ( .A(n36855), .B(n36854), .Z(n36903) );
  XOR U37858 ( .A(n36902), .B(n36903), .Z(n36910) );
  AND U37859 ( .A(x[484]), .B(y[8069]), .Z(n37402) );
  NAND U37860 ( .A(n37402), .B(n36881), .Z(n36859) );
  NAND U37861 ( .A(n36857), .B(n36856), .Z(n36858) );
  AND U37862 ( .A(n36859), .B(n36858), .Z(n36878) );
  AND U37863 ( .A(y[8069]), .B(x[482]), .Z(n36861) );
  NAND U37864 ( .A(y[8067]), .B(x[484]), .Z(n36860) );
  XNOR U37865 ( .A(n36861), .B(n36860), .Z(n36891) );
  XNOR U37866 ( .A(n36891), .B(n36890), .Z(n36876) );
  AND U37867 ( .A(y[8064]), .B(x[487]), .Z(n36863) );
  NAND U37868 ( .A(y[8071]), .B(x[480]), .Z(n36862) );
  XNOR U37869 ( .A(n36863), .B(n36862), .Z(n36895) );
  AND U37870 ( .A(o[390]), .B(n36864), .Z(n36894) );
  XNOR U37871 ( .A(n36895), .B(n36894), .Z(n36875) );
  XOR U37872 ( .A(n36876), .B(n36875), .Z(n36877) );
  XOR U37873 ( .A(n36878), .B(n36877), .Z(n36909) );
  XOR U37874 ( .A(n36910), .B(n36909), .Z(n36911) );
  XOR U37875 ( .A(n36912), .B(n36911), .Z(n36908) );
  NAND U37876 ( .A(n36866), .B(n36865), .Z(n36870) );
  NAND U37877 ( .A(n36868), .B(n36867), .Z(n36869) );
  NAND U37878 ( .A(n36870), .B(n36869), .Z(n36907) );
  XOR U37879 ( .A(n36907), .B(n36906), .Z(n36874) );
  XNOR U37880 ( .A(n36908), .B(n36874), .Z(N808) );
  NAND U37881 ( .A(n36876), .B(n36875), .Z(n36880) );
  NAND U37882 ( .A(n36878), .B(n36877), .Z(n36879) );
  AND U37883 ( .A(n36880), .B(n36879), .Z(n36962) );
  AND U37884 ( .A(x[485]), .B(y[8070]), .Z(n37056) );
  NAND U37885 ( .A(n37056), .B(n36881), .Z(n36885) );
  NAND U37886 ( .A(n36883), .B(n36882), .Z(n36884) );
  NAND U37887 ( .A(n36885), .B(n36884), .Z(n36960) );
  AND U37888 ( .A(o[391]), .B(n36886), .Z(n36949) );
  AND U37889 ( .A(y[8067]), .B(x[485]), .Z(n37503) );
  NAND U37890 ( .A(y[8071]), .B(x[481]), .Z(n36887) );
  XNOR U37891 ( .A(n37503), .B(n36887), .Z(n36950) );
  XNOR U37892 ( .A(n36949), .B(n36950), .Z(n36934) );
  NAND U37893 ( .A(x[483]), .B(y[8069]), .Z(n37721) );
  AND U37894 ( .A(x[486]), .B(y[8066]), .Z(n36888) );
  AND U37895 ( .A(y[8070]), .B(x[482]), .Z(n37800) );
  XOR U37896 ( .A(n36888), .B(n37800), .Z(n36930) );
  XOR U37897 ( .A(n37595), .B(n36930), .Z(n36933) );
  XOR U37898 ( .A(n36934), .B(n36935), .Z(n36959) );
  XOR U37899 ( .A(n36960), .B(n36959), .Z(n36961) );
  XNOR U37900 ( .A(n36962), .B(n36961), .Z(n36919) );
  NANDN U37901 ( .A(n36889), .B(n37402), .Z(n36893) );
  NAND U37902 ( .A(n36891), .B(n36890), .Z(n36892) );
  NAND U37903 ( .A(n36893), .B(n36892), .Z(n36956) );
  AND U37904 ( .A(x[487]), .B(y[8071]), .Z(n37280) );
  NAND U37905 ( .A(n37397), .B(n37280), .Z(n36897) );
  NAND U37906 ( .A(n36895), .B(n36894), .Z(n36896) );
  NAND U37907 ( .A(n36897), .B(n36896), .Z(n36954) );
  AND U37908 ( .A(y[8064]), .B(x[488]), .Z(n36899) );
  NAND U37909 ( .A(y[8072]), .B(x[480]), .Z(n36898) );
  XNOR U37910 ( .A(n36899), .B(n36898), .Z(n36940) );
  AND U37911 ( .A(x[487]), .B(y[8065]), .Z(n36943) );
  XOR U37912 ( .A(o[392]), .B(n36943), .Z(n36939) );
  XOR U37913 ( .A(n36940), .B(n36939), .Z(n36953) );
  XOR U37914 ( .A(n36954), .B(n36953), .Z(n36955) );
  XNOR U37915 ( .A(n36956), .B(n36955), .Z(n36917) );
  NAND U37916 ( .A(n36901), .B(n36900), .Z(n36905) );
  NAND U37917 ( .A(n36903), .B(n36902), .Z(n36904) );
  NAND U37918 ( .A(n36905), .B(n36904), .Z(n36916) );
  XOR U37919 ( .A(n36917), .B(n36916), .Z(n36918) );
  XOR U37920 ( .A(n36919), .B(n36918), .Z(n36925) );
  NAND U37921 ( .A(n36910), .B(n36909), .Z(n36914) );
  NAND U37922 ( .A(n36912), .B(n36911), .Z(n36913) );
  AND U37923 ( .A(n36914), .B(n36913), .Z(n36923) );
  IV U37924 ( .A(n36923), .Z(n36922) );
  XOR U37925 ( .A(n36924), .B(n36922), .Z(n36915) );
  XNOR U37926 ( .A(n36925), .B(n36915), .Z(N809) );
  NAND U37927 ( .A(n36917), .B(n36916), .Z(n36921) );
  NAND U37928 ( .A(n36919), .B(n36918), .Z(n36920) );
  NAND U37929 ( .A(n36921), .B(n36920), .Z(n37016) );
  IV U37930 ( .A(n37016), .Z(n37014) );
  OR U37931 ( .A(n36924), .B(n36922), .Z(n36928) );
  ANDN U37932 ( .B(n36924), .A(n36923), .Z(n36926) );
  OR U37933 ( .A(n36926), .B(n36925), .Z(n36927) );
  AND U37934 ( .A(n36928), .B(n36927), .Z(n37015) );
  NAND U37935 ( .A(n37131), .B(n36929), .Z(n36932) );
  NAND U37936 ( .A(n37595), .B(n36930), .Z(n36931) );
  NAND U37937 ( .A(n36932), .B(n36931), .Z(n36966) );
  NANDN U37938 ( .A(n36933), .B(n37721), .Z(n36937) );
  NANDN U37939 ( .A(n36935), .B(n36934), .Z(n36936) );
  AND U37940 ( .A(n36937), .B(n36936), .Z(n36967) );
  XOR U37941 ( .A(n36966), .B(n36967), .Z(n36968) );
  AND U37942 ( .A(x[488]), .B(y[8072]), .Z(n36938) );
  NAND U37943 ( .A(n36938), .B(n37397), .Z(n36942) );
  NAND U37944 ( .A(n36940), .B(n36939), .Z(n36941) );
  AND U37945 ( .A(n36942), .B(n36941), .Z(n37001) );
  AND U37946 ( .A(o[392]), .B(n36943), .Z(n36974) );
  AND U37947 ( .A(y[8068]), .B(x[485]), .Z(n36945) );
  NAND U37948 ( .A(y[8066]), .B(x[487]), .Z(n36944) );
  XNOR U37949 ( .A(n36945), .B(n36944), .Z(n36973) );
  XNOR U37950 ( .A(n36974), .B(n36973), .Z(n36999) );
  AND U37951 ( .A(y[8064]), .B(x[489]), .Z(n36947) );
  NAND U37952 ( .A(y[8073]), .B(x[480]), .Z(n36946) );
  XNOR U37953 ( .A(n36947), .B(n36946), .Z(n36981) );
  AND U37954 ( .A(x[488]), .B(y[8065]), .Z(n36990) );
  XOR U37955 ( .A(o[393]), .B(n36990), .Z(n36980) );
  XNOR U37956 ( .A(n36981), .B(n36980), .Z(n36998) );
  XOR U37957 ( .A(n36999), .B(n36998), .Z(n37000) );
  XNOR U37958 ( .A(n37001), .B(n37000), .Z(n36995) );
  AND U37959 ( .A(y[8067]), .B(x[486]), .Z(n37345) );
  NAND U37960 ( .A(y[8072]), .B(x[481]), .Z(n36948) );
  XNOR U37961 ( .A(n37345), .B(n36948), .Z(n36985) );
  XNOR U37962 ( .A(n37402), .B(n36985), .Z(n37005) );
  NAND U37963 ( .A(x[482]), .B(y[8071]), .Z(n37634) );
  AND U37964 ( .A(x[483]), .B(y[8070]), .Z(n37355) );
  XNOR U37965 ( .A(n37634), .B(n37355), .Z(n37004) );
  XNOR U37966 ( .A(n37005), .B(n37004), .Z(n36993) );
  NAND U37967 ( .A(x[485]), .B(y[8071]), .Z(n37194) );
  AND U37968 ( .A(x[481]), .B(y[8067]), .Z(n36984) );
  NANDN U37969 ( .A(n37194), .B(n36984), .Z(n36952) );
  NAND U37970 ( .A(n36950), .B(n36949), .Z(n36951) );
  NAND U37971 ( .A(n36952), .B(n36951), .Z(n36992) );
  XOR U37972 ( .A(n36993), .B(n36992), .Z(n36994) );
  XNOR U37973 ( .A(n36995), .B(n36994), .Z(n36969) );
  XNOR U37974 ( .A(n36968), .B(n36969), .Z(n37011) );
  NAND U37975 ( .A(n36954), .B(n36953), .Z(n36958) );
  NAND U37976 ( .A(n36956), .B(n36955), .Z(n36957) );
  NAND U37977 ( .A(n36958), .B(n36957), .Z(n37009) );
  NAND U37978 ( .A(n36960), .B(n36959), .Z(n36964) );
  NAND U37979 ( .A(n36962), .B(n36961), .Z(n36963) );
  NAND U37980 ( .A(n36964), .B(n36963), .Z(n37008) );
  XOR U37981 ( .A(n37009), .B(n37008), .Z(n37010) );
  XOR U37982 ( .A(n37011), .B(n37010), .Z(n37017) );
  XNOR U37983 ( .A(n37015), .B(n37017), .Z(n36965) );
  XOR U37984 ( .A(n37014), .B(n36965), .Z(N810) );
  NAND U37985 ( .A(n36967), .B(n36966), .Z(n36971) );
  NANDN U37986 ( .A(n36969), .B(n36968), .Z(n36970) );
  AND U37987 ( .A(n36971), .B(n36970), .Z(n37079) );
  AND U37988 ( .A(x[487]), .B(y[8068]), .Z(n37058) );
  NAND U37989 ( .A(n37058), .B(n36972), .Z(n36976) );
  NAND U37990 ( .A(n36974), .B(n36973), .Z(n36975) );
  AND U37991 ( .A(n36976), .B(n36975), .Z(n37071) );
  AND U37992 ( .A(y[8067]), .B(x[487]), .Z(n36978) );
  NAND U37993 ( .A(y[8070]), .B(x[484]), .Z(n36977) );
  XNOR U37994 ( .A(n36978), .B(n36977), .Z(n37042) );
  AND U37995 ( .A(x[486]), .B(y[8068]), .Z(n37041) );
  XNOR U37996 ( .A(n37042), .B(n37041), .Z(n37069) );
  AND U37997 ( .A(x[488]), .B(y[8066]), .Z(n37254) );
  AND U37998 ( .A(x[489]), .B(y[8065]), .Z(n37052) );
  XOR U37999 ( .A(o[394]), .B(n37052), .Z(n37063) );
  XOR U38000 ( .A(n37254), .B(n37063), .Z(n37065) );
  XNOR U38001 ( .A(n37065), .B(n37064), .Z(n37068) );
  XOR U38002 ( .A(n37069), .B(n37068), .Z(n37070) );
  XNOR U38003 ( .A(n37071), .B(n37070), .Z(n37031) );
  AND U38004 ( .A(x[489]), .B(y[8073]), .Z(n36979) );
  NAND U38005 ( .A(n36979), .B(n37397), .Z(n36983) );
  NAND U38006 ( .A(n36981), .B(n36980), .Z(n36982) );
  NAND U38007 ( .A(n36983), .B(n36982), .Z(n37029) );
  AND U38008 ( .A(x[486]), .B(y[8072]), .Z(n37290) );
  NAND U38009 ( .A(n37290), .B(n36984), .Z(n36987) );
  NAND U38010 ( .A(n37402), .B(n36985), .Z(n36986) );
  NAND U38011 ( .A(n36987), .B(n36986), .Z(n37037) );
  AND U38012 ( .A(y[8064]), .B(x[490]), .Z(n36989) );
  NAND U38013 ( .A(y[8074]), .B(x[480]), .Z(n36988) );
  XNOR U38014 ( .A(n36989), .B(n36988), .Z(n37047) );
  AND U38015 ( .A(o[393]), .B(n36990), .Z(n37046) );
  XOR U38016 ( .A(n37047), .B(n37046), .Z(n37035) );
  AND U38017 ( .A(y[8071]), .B(x[483]), .Z(n37943) );
  NAND U38018 ( .A(y[8073]), .B(x[481]), .Z(n36991) );
  XNOR U38019 ( .A(n37943), .B(n36991), .Z(n37059) );
  AND U38020 ( .A(x[482]), .B(y[8072]), .Z(n37060) );
  XOR U38021 ( .A(n37059), .B(n37060), .Z(n37034) );
  XOR U38022 ( .A(n37035), .B(n37034), .Z(n37036) );
  XOR U38023 ( .A(n37037), .B(n37036), .Z(n37028) );
  XOR U38024 ( .A(n37029), .B(n37028), .Z(n37030) );
  XOR U38025 ( .A(n37031), .B(n37030), .Z(n37078) );
  NAND U38026 ( .A(n36993), .B(n36992), .Z(n36997) );
  NAND U38027 ( .A(n36995), .B(n36994), .Z(n36996) );
  NAND U38028 ( .A(n36997), .B(n36996), .Z(n37025) );
  NAND U38029 ( .A(n36999), .B(n36998), .Z(n37003) );
  NAND U38030 ( .A(n37001), .B(n37000), .Z(n37002) );
  AND U38031 ( .A(n37003), .B(n37002), .Z(n37022) );
  NAND U38032 ( .A(n37005), .B(n37004), .Z(n37007) );
  ANDN U38033 ( .B(n37634), .A(n37355), .Z(n37006) );
  ANDN U38034 ( .B(n37007), .A(n37006), .Z(n37023) );
  XOR U38035 ( .A(n37022), .B(n37023), .Z(n37024) );
  XNOR U38036 ( .A(n37025), .B(n37024), .Z(n37077) );
  XNOR U38037 ( .A(n37079), .B(n37080), .Z(n37076) );
  NAND U38038 ( .A(n37009), .B(n37008), .Z(n37013) );
  NAND U38039 ( .A(n37011), .B(n37010), .Z(n37012) );
  NAND U38040 ( .A(n37013), .B(n37012), .Z(n37075) );
  NANDN U38041 ( .A(n37014), .B(n37015), .Z(n37020) );
  NOR U38042 ( .A(n37016), .B(n37015), .Z(n37018) );
  OR U38043 ( .A(n37018), .B(n37017), .Z(n37019) );
  AND U38044 ( .A(n37020), .B(n37019), .Z(n37074) );
  XOR U38045 ( .A(n37075), .B(n37074), .Z(n37021) );
  XNOR U38046 ( .A(n37076), .B(n37021), .Z(N811) );
  NAND U38047 ( .A(n37023), .B(n37022), .Z(n37027) );
  NAND U38048 ( .A(n37025), .B(n37024), .Z(n37026) );
  AND U38049 ( .A(n37027), .B(n37026), .Z(n37149) );
  NAND U38050 ( .A(n37029), .B(n37028), .Z(n37033) );
  NAND U38051 ( .A(n37031), .B(n37030), .Z(n37032) );
  NAND U38052 ( .A(n37033), .B(n37032), .Z(n37147) );
  NAND U38053 ( .A(n37035), .B(n37034), .Z(n37039) );
  NAND U38054 ( .A(n37037), .B(n37036), .Z(n37038) );
  NAND U38055 ( .A(n37039), .B(n37038), .Z(n37097) );
  AND U38056 ( .A(x[487]), .B(y[8070]), .Z(n37189) );
  AND U38057 ( .A(x[484]), .B(y[8067]), .Z(n37040) );
  NAND U38058 ( .A(n37189), .B(n37040), .Z(n37044) );
  NAND U38059 ( .A(n37042), .B(n37041), .Z(n37043) );
  NAND U38060 ( .A(n37044), .B(n37043), .Z(n37095) );
  AND U38061 ( .A(x[490]), .B(y[8074]), .Z(n37045) );
  NAND U38062 ( .A(n37045), .B(n37397), .Z(n37049) );
  NAND U38063 ( .A(n37047), .B(n37046), .Z(n37048) );
  NAND U38064 ( .A(n37049), .B(n37048), .Z(n37091) );
  AND U38065 ( .A(y[8064]), .B(x[491]), .Z(n37051) );
  NAND U38066 ( .A(y[8075]), .B(x[480]), .Z(n37050) );
  XNOR U38067 ( .A(n37051), .B(n37050), .Z(n37122) );
  AND U38068 ( .A(o[394]), .B(n37052), .Z(n37121) );
  XOR U38069 ( .A(n37122), .B(n37121), .Z(n37090) );
  AND U38070 ( .A(y[8069]), .B(x[486]), .Z(n37054) );
  NAND U38071 ( .A(y[8074]), .B(x[481]), .Z(n37053) );
  XNOR U38072 ( .A(n37054), .B(n37053), .Z(n37113) );
  AND U38073 ( .A(x[490]), .B(y[8065]), .Z(n37132) );
  XOR U38074 ( .A(o[395]), .B(n37132), .Z(n37112) );
  XOR U38075 ( .A(n37113), .B(n37112), .Z(n37089) );
  XOR U38076 ( .A(n37090), .B(n37089), .Z(n37092) );
  XOR U38077 ( .A(n37091), .B(n37092), .Z(n37096) );
  XNOR U38078 ( .A(n37095), .B(n37096), .Z(n37098) );
  XOR U38079 ( .A(n37097), .B(n37098), .Z(n37135) );
  AND U38080 ( .A(x[483]), .B(y[8072]), .Z(n38084) );
  NAND U38081 ( .A(y[8073]), .B(x[482]), .Z(n37055) );
  XNOR U38082 ( .A(n37056), .B(n37055), .Z(n37108) );
  AND U38083 ( .A(x[484]), .B(y[8071]), .Z(n37107) );
  XNOR U38084 ( .A(n37108), .B(n37107), .Z(n37084) );
  XNOR U38085 ( .A(n38084), .B(n37084), .Z(n37086) );
  NAND U38086 ( .A(y[8066]), .B(x[489]), .Z(n37057) );
  XNOR U38087 ( .A(n37058), .B(n37057), .Z(n37127) );
  AND U38088 ( .A(x[488]), .B(y[8067]), .Z(n37126) );
  XNOR U38089 ( .A(n37127), .B(n37126), .Z(n37085) );
  XNOR U38090 ( .A(n37086), .B(n37085), .Z(n37104) );
  NAND U38091 ( .A(x[483]), .B(y[8073]), .Z(n37185) );
  AND U38092 ( .A(x[481]), .B(y[8071]), .Z(n37392) );
  NANDN U38093 ( .A(n37185), .B(n37392), .Z(n37062) );
  NAND U38094 ( .A(n37060), .B(n37059), .Z(n37061) );
  NAND U38095 ( .A(n37062), .B(n37061), .Z(n37102) );
  NAND U38096 ( .A(n37254), .B(n37063), .Z(n37067) );
  NAND U38097 ( .A(n37065), .B(n37064), .Z(n37066) );
  NAND U38098 ( .A(n37067), .B(n37066), .Z(n37101) );
  XOR U38099 ( .A(n37102), .B(n37101), .Z(n37103) );
  XNOR U38100 ( .A(n37104), .B(n37103), .Z(n37134) );
  NAND U38101 ( .A(n37069), .B(n37068), .Z(n37073) );
  NAND U38102 ( .A(n37071), .B(n37070), .Z(n37072) );
  NAND U38103 ( .A(n37073), .B(n37072), .Z(n37133) );
  XOR U38104 ( .A(n37134), .B(n37133), .Z(n37136) );
  XNOR U38105 ( .A(n37135), .B(n37136), .Z(n37146) );
  XOR U38106 ( .A(n37147), .B(n37146), .Z(n37148) );
  XOR U38107 ( .A(n37149), .B(n37148), .Z(n37142) );
  NANDN U38108 ( .A(n37078), .B(n37077), .Z(n37082) );
  NANDN U38109 ( .A(n37080), .B(n37079), .Z(n37081) );
  AND U38110 ( .A(n37082), .B(n37081), .Z(n37140) );
  IV U38111 ( .A(n37140), .Z(n37139) );
  XOR U38112 ( .A(n37141), .B(n37139), .Z(n37083) );
  XNOR U38113 ( .A(n37142), .B(n37083), .Z(N812) );
  NANDN U38114 ( .A(n38084), .B(n37084), .Z(n37088) );
  NAND U38115 ( .A(n37086), .B(n37085), .Z(n37087) );
  NAND U38116 ( .A(n37088), .B(n37087), .Z(n37166) );
  NAND U38117 ( .A(n37090), .B(n37089), .Z(n37094) );
  NAND U38118 ( .A(n37092), .B(n37091), .Z(n37093) );
  AND U38119 ( .A(n37094), .B(n37093), .Z(n37167) );
  XOR U38120 ( .A(n37166), .B(n37167), .Z(n37169) );
  NAND U38121 ( .A(n37096), .B(n37095), .Z(n37100) );
  NANDN U38122 ( .A(n37098), .B(n37097), .Z(n37099) );
  AND U38123 ( .A(n37100), .B(n37099), .Z(n37168) );
  XOR U38124 ( .A(n37169), .B(n37168), .Z(n37156) );
  NAND U38125 ( .A(n37102), .B(n37101), .Z(n37106) );
  NAND U38126 ( .A(n37104), .B(n37103), .Z(n37105) );
  NAND U38127 ( .A(n37106), .B(n37105), .Z(n37225) );
  AND U38128 ( .A(x[485]), .B(y[8073]), .Z(n37625) );
  NAND U38129 ( .A(n37800), .B(n37625), .Z(n37110) );
  NAND U38130 ( .A(n37108), .B(n37107), .Z(n37109) );
  NAND U38131 ( .A(n37110), .B(n37109), .Z(n37173) );
  AND U38132 ( .A(x[486]), .B(y[8074]), .Z(n37409) );
  NAND U38133 ( .A(n37409), .B(n37111), .Z(n37115) );
  NAND U38134 ( .A(n37113), .B(n37112), .Z(n37114) );
  NAND U38135 ( .A(n37115), .B(n37114), .Z(n37172) );
  XOR U38136 ( .A(n37173), .B(n37172), .Z(n37175) );
  AND U38137 ( .A(x[489]), .B(y[8067]), .Z(n37795) );
  AND U38138 ( .A(y[8066]), .B(x[490]), .Z(n37837) );
  NAND U38139 ( .A(y[8072]), .B(x[484]), .Z(n37116) );
  XNOR U38140 ( .A(n37837), .B(n37116), .Z(n37216) );
  XOR U38141 ( .A(n37795), .B(n37216), .Z(n37195) );
  NAND U38142 ( .A(x[487]), .B(y[8069]), .Z(n37193) );
  XOR U38143 ( .A(n37194), .B(n37193), .Z(n37196) );
  AND U38144 ( .A(y[8064]), .B(x[492]), .Z(n37118) );
  NAND U38145 ( .A(y[8076]), .B(x[480]), .Z(n37117) );
  XNOR U38146 ( .A(n37118), .B(n37117), .Z(n37210) );
  AND U38147 ( .A(x[491]), .B(y[8065]), .Z(n37190) );
  XOR U38148 ( .A(o[396]), .B(n37190), .Z(n37209) );
  XOR U38149 ( .A(n37210), .B(n37209), .Z(n37179) );
  AND U38150 ( .A(y[8074]), .B(x[482]), .Z(n37120) );
  NAND U38151 ( .A(y[8068]), .B(x[488]), .Z(n37119) );
  XNOR U38152 ( .A(n37120), .B(n37119), .Z(n37184) );
  XOR U38153 ( .A(n37179), .B(n37178), .Z(n37181) );
  XOR U38154 ( .A(n37180), .B(n37181), .Z(n37174) );
  XOR U38155 ( .A(n37175), .B(n37174), .Z(n37224) );
  AND U38156 ( .A(x[491]), .B(y[8075]), .Z(n38191) );
  NAND U38157 ( .A(n38191), .B(n37397), .Z(n37124) );
  NAND U38158 ( .A(n37122), .B(n37121), .Z(n37123) );
  NAND U38159 ( .A(n37124), .B(n37123), .Z(n37202) );
  AND U38160 ( .A(x[487]), .B(y[8066]), .Z(n37331) );
  AND U38161 ( .A(x[489]), .B(y[8068]), .Z(n37125) );
  NAND U38162 ( .A(n37331), .B(n37125), .Z(n37129) );
  NAND U38163 ( .A(n37127), .B(n37126), .Z(n37128) );
  NAND U38164 ( .A(n37129), .B(n37128), .Z(n37200) );
  NAND U38165 ( .A(y[8075]), .B(x[481]), .Z(n37130) );
  XNOR U38166 ( .A(n37131), .B(n37130), .Z(n37206) );
  AND U38167 ( .A(o[395]), .B(n37132), .Z(n37205) );
  XOR U38168 ( .A(n37206), .B(n37205), .Z(n37199) );
  XOR U38169 ( .A(n37200), .B(n37199), .Z(n37201) );
  XOR U38170 ( .A(n37202), .B(n37201), .Z(n37223) );
  XOR U38171 ( .A(n37224), .B(n37223), .Z(n37226) );
  XNOR U38172 ( .A(n37225), .B(n37226), .Z(n37154) );
  NAND U38173 ( .A(n37134), .B(n37133), .Z(n37138) );
  NAND U38174 ( .A(n37136), .B(n37135), .Z(n37137) );
  NAND U38175 ( .A(n37138), .B(n37137), .Z(n37153) );
  XOR U38176 ( .A(n37154), .B(n37153), .Z(n37155) );
  XNOR U38177 ( .A(n37156), .B(n37155), .Z(n37163) );
  OR U38178 ( .A(n37141), .B(n37139), .Z(n37145) );
  ANDN U38179 ( .B(n37141), .A(n37140), .Z(n37143) );
  OR U38180 ( .A(n37143), .B(n37142), .Z(n37144) );
  AND U38181 ( .A(n37145), .B(n37144), .Z(n37160) );
  NAND U38182 ( .A(n37147), .B(n37146), .Z(n37151) );
  NANDN U38183 ( .A(n37149), .B(n37148), .Z(n37150) );
  AND U38184 ( .A(n37151), .B(n37150), .Z(n37161) );
  IV U38185 ( .A(n37161), .Z(n37159) );
  XOR U38186 ( .A(n37160), .B(n37159), .Z(n37152) );
  XNOR U38187 ( .A(n37163), .B(n37152), .Z(N813) );
  NAND U38188 ( .A(n37154), .B(n37153), .Z(n37158) );
  NAND U38189 ( .A(n37156), .B(n37155), .Z(n37157) );
  AND U38190 ( .A(n37158), .B(n37157), .Z(n37304) );
  NANDN U38191 ( .A(n37159), .B(n37160), .Z(n37165) );
  NOR U38192 ( .A(n37161), .B(n37160), .Z(n37162) );
  OR U38193 ( .A(n37163), .B(n37162), .Z(n37164) );
  AND U38194 ( .A(n37165), .B(n37164), .Z(n37303) );
  NAND U38195 ( .A(n37167), .B(n37166), .Z(n37171) );
  NAND U38196 ( .A(n37169), .B(n37168), .Z(n37170) );
  NAND U38197 ( .A(n37171), .B(n37170), .Z(n37299) );
  NAND U38198 ( .A(n37173), .B(n37172), .Z(n37177) );
  NAND U38199 ( .A(n37175), .B(n37174), .Z(n37176) );
  AND U38200 ( .A(n37177), .B(n37176), .Z(n37231) );
  NAND U38201 ( .A(n37179), .B(n37178), .Z(n37183) );
  NAND U38202 ( .A(n37181), .B(n37180), .Z(n37182) );
  NAND U38203 ( .A(n37183), .B(n37182), .Z(n37238) );
  AND U38204 ( .A(y[8074]), .B(x[488]), .Z(n38477) );
  AND U38205 ( .A(x[482]), .B(y[8068]), .Z(n37341) );
  NAND U38206 ( .A(n38477), .B(n37341), .Z(n37187) );
  NANDN U38207 ( .A(n37185), .B(n37184), .Z(n37186) );
  NAND U38208 ( .A(n37187), .B(n37186), .Z(n37269) );
  NAND U38209 ( .A(y[8076]), .B(x[481]), .Z(n37188) );
  XNOR U38210 ( .A(n37189), .B(n37188), .Z(n37260) );
  AND U38211 ( .A(o[396]), .B(n37190), .Z(n37259) );
  XOR U38212 ( .A(n37260), .B(n37259), .Z(n37267) );
  AND U38213 ( .A(x[486]), .B(y[8071]), .Z(n38231) );
  AND U38214 ( .A(y[8075]), .B(x[482]), .Z(n37192) );
  NAND U38215 ( .A(y[8068]), .B(x[489]), .Z(n37191) );
  XNOR U38216 ( .A(n37192), .B(n37191), .Z(n37273) );
  XOR U38217 ( .A(n38231), .B(n37273), .Z(n37266) );
  XOR U38218 ( .A(n37267), .B(n37266), .Z(n37268) );
  XOR U38219 ( .A(n37269), .B(n37268), .Z(n37237) );
  NAND U38220 ( .A(n37194), .B(n37193), .Z(n37198) );
  ANDN U38221 ( .B(n37196), .A(n37195), .Z(n37197) );
  ANDN U38222 ( .B(n37198), .A(n37197), .Z(n37236) );
  XOR U38223 ( .A(n37237), .B(n37236), .Z(n37239) );
  XOR U38224 ( .A(n37238), .B(n37239), .Z(n37230) );
  NAND U38225 ( .A(n37200), .B(n37199), .Z(n37204) );
  NAND U38226 ( .A(n37202), .B(n37201), .Z(n37203) );
  NAND U38227 ( .A(n37204), .B(n37203), .Z(n37245) );
  AND U38228 ( .A(x[486]), .B(y[8075]), .Z(n37556) );
  IV U38229 ( .A(n37556), .Z(n37627) );
  AND U38230 ( .A(x[481]), .B(y[8070]), .Z(n37258) );
  NANDN U38231 ( .A(n37627), .B(n37258), .Z(n37208) );
  NAND U38232 ( .A(n37206), .B(n37205), .Z(n37207) );
  NAND U38233 ( .A(n37208), .B(n37207), .Z(n37251) );
  AND U38234 ( .A(x[492]), .B(y[8076]), .Z(n38483) );
  NAND U38235 ( .A(n38483), .B(n37397), .Z(n37212) );
  NAND U38236 ( .A(n37210), .B(n37209), .Z(n37211) );
  NAND U38237 ( .A(n37212), .B(n37211), .Z(n37249) );
  AND U38238 ( .A(x[490]), .B(y[8067]), .Z(n38096) );
  AND U38239 ( .A(y[8066]), .B(x[491]), .Z(n38045) );
  NAND U38240 ( .A(y[8069]), .B(x[488]), .Z(n37213) );
  XNOR U38241 ( .A(n38045), .B(n37213), .Z(n37255) );
  XOR U38242 ( .A(n38096), .B(n37255), .Z(n37248) );
  XOR U38243 ( .A(n37249), .B(n37248), .Z(n37250) );
  XOR U38244 ( .A(n37251), .B(n37250), .Z(n37243) );
  AND U38245 ( .A(x[490]), .B(y[8072]), .Z(n37215) );
  AND U38246 ( .A(x[484]), .B(y[8066]), .Z(n37214) );
  NAND U38247 ( .A(n37215), .B(n37214), .Z(n37218) );
  NAND U38248 ( .A(n37216), .B(n37795), .Z(n37217) );
  NAND U38249 ( .A(n37218), .B(n37217), .Z(n37294) );
  AND U38250 ( .A(y[8064]), .B(x[493]), .Z(n37220) );
  NAND U38251 ( .A(y[8077]), .B(x[480]), .Z(n37219) );
  XNOR U38252 ( .A(n37220), .B(n37219), .Z(n37286) );
  AND U38253 ( .A(x[492]), .B(y[8065]), .Z(n37278) );
  XOR U38254 ( .A(o[397]), .B(n37278), .Z(n37285) );
  XOR U38255 ( .A(n37286), .B(n37285), .Z(n37292) );
  AND U38256 ( .A(y[8072]), .B(x[485]), .Z(n37222) );
  NAND U38257 ( .A(y[8074]), .B(x[483]), .Z(n37221) );
  XNOR U38258 ( .A(n37222), .B(n37221), .Z(n37281) );
  AND U38259 ( .A(x[484]), .B(y[8073]), .Z(n37282) );
  XOR U38260 ( .A(n37281), .B(n37282), .Z(n37291) );
  XOR U38261 ( .A(n37292), .B(n37291), .Z(n37293) );
  XOR U38262 ( .A(n37294), .B(n37293), .Z(n37242) );
  XOR U38263 ( .A(n37243), .B(n37242), .Z(n37244) );
  XOR U38264 ( .A(n37245), .B(n37244), .Z(n37232) );
  XNOR U38265 ( .A(n37233), .B(n37232), .Z(n37298) );
  NAND U38266 ( .A(n37224), .B(n37223), .Z(n37228) );
  NAND U38267 ( .A(n37226), .B(n37225), .Z(n37227) );
  AND U38268 ( .A(n37228), .B(n37227), .Z(n37297) );
  XOR U38269 ( .A(n37298), .B(n37297), .Z(n37300) );
  XOR U38270 ( .A(n37299), .B(n37300), .Z(n37305) );
  XNOR U38271 ( .A(n37303), .B(n37305), .Z(n37229) );
  XOR U38272 ( .A(n37304), .B(n37229), .Z(N814) );
  NANDN U38273 ( .A(n37231), .B(n37230), .Z(n37235) );
  NAND U38274 ( .A(n37233), .B(n37232), .Z(n37234) );
  AND U38275 ( .A(n37235), .B(n37234), .Z(n37383) );
  NAND U38276 ( .A(n37237), .B(n37236), .Z(n37241) );
  NAND U38277 ( .A(n37239), .B(n37238), .Z(n37240) );
  NAND U38278 ( .A(n37241), .B(n37240), .Z(n37382) );
  NAND U38279 ( .A(n37243), .B(n37242), .Z(n37247) );
  NAND U38280 ( .A(n37245), .B(n37244), .Z(n37246) );
  NAND U38281 ( .A(n37247), .B(n37246), .Z(n37310) );
  NAND U38282 ( .A(n37249), .B(n37248), .Z(n37253) );
  NAND U38283 ( .A(n37251), .B(n37250), .Z(n37252) );
  AND U38284 ( .A(n37253), .B(n37252), .Z(n37316) );
  AND U38285 ( .A(x[491]), .B(y[8069]), .Z(n37424) );
  NAND U38286 ( .A(n37424), .B(n37254), .Z(n37257) );
  NAND U38287 ( .A(n37255), .B(n38096), .Z(n37256) );
  NAND U38288 ( .A(n37257), .B(n37256), .Z(n37371) );
  NAND U38289 ( .A(x[487]), .B(y[8076]), .Z(n37810) );
  NANDN U38290 ( .A(n37810), .B(n37258), .Z(n37262) );
  NAND U38291 ( .A(n37260), .B(n37259), .Z(n37261) );
  NAND U38292 ( .A(n37262), .B(n37261), .Z(n37370) );
  XOR U38293 ( .A(n37371), .B(n37370), .Z(n37373) );
  AND U38294 ( .A(x[484]), .B(y[8074]), .Z(n37730) );
  AND U38295 ( .A(y[8075]), .B(x[483]), .Z(n37264) );
  NAND U38296 ( .A(y[8070]), .B(x[488]), .Z(n37263) );
  XNOR U38297 ( .A(n37264), .B(n37263), .Z(n37356) );
  XOR U38298 ( .A(n37625), .B(n37356), .Z(n37365) );
  XOR U38299 ( .A(n37730), .B(n37365), .Z(n37367) );
  AND U38300 ( .A(x[489]), .B(y[8069]), .Z(n37914) );
  AND U38301 ( .A(y[8076]), .B(x[482]), .Z(n37265) );
  AND U38302 ( .A(y[8068]), .B(x[490]), .Z(n37938) );
  XOR U38303 ( .A(n37265), .B(n37938), .Z(n37342) );
  XOR U38304 ( .A(n37914), .B(n37342), .Z(n37366) );
  XOR U38305 ( .A(n37367), .B(n37366), .Z(n37372) );
  XNOR U38306 ( .A(n37373), .B(n37372), .Z(n37314) );
  NAND U38307 ( .A(n37267), .B(n37266), .Z(n37271) );
  NAND U38308 ( .A(n37269), .B(n37268), .Z(n37270) );
  AND U38309 ( .A(n37271), .B(n37270), .Z(n37313) );
  XOR U38310 ( .A(n37314), .B(n37313), .Z(n37315) );
  XNOR U38311 ( .A(n37316), .B(n37315), .Z(n37308) );
  AND U38312 ( .A(x[489]), .B(y[8075]), .Z(n37272) );
  NAND U38313 ( .A(n37272), .B(n37341), .Z(n37275) );
  NAND U38314 ( .A(n37273), .B(n38231), .Z(n37274) );
  NAND U38315 ( .A(n37275), .B(n37274), .Z(n37328) );
  AND U38316 ( .A(y[8064]), .B(x[494]), .Z(n37277) );
  NAND U38317 ( .A(y[8078]), .B(x[480]), .Z(n37276) );
  XNOR U38318 ( .A(n37277), .B(n37276), .Z(n37351) );
  AND U38319 ( .A(o[397]), .B(n37278), .Z(n37350) );
  XOR U38320 ( .A(n37351), .B(n37350), .Z(n37326) );
  NAND U38321 ( .A(y[8066]), .B(x[492]), .Z(n37279) );
  XNOR U38322 ( .A(n37280), .B(n37279), .Z(n37333) );
  AND U38323 ( .A(x[493]), .B(y[8065]), .Z(n37340) );
  XOR U38324 ( .A(n37340), .B(o[398]), .Z(n37332) );
  XOR U38325 ( .A(n37333), .B(n37332), .Z(n37325) );
  XOR U38326 ( .A(n37326), .B(n37325), .Z(n37327) );
  XNOR U38327 ( .A(n37328), .B(n37327), .Z(n37377) );
  NAND U38328 ( .A(x[485]), .B(y[8074]), .Z(n37411) );
  NANDN U38329 ( .A(n37411), .B(n38084), .Z(n37284) );
  NAND U38330 ( .A(n37282), .B(n37281), .Z(n37283) );
  AND U38331 ( .A(n37284), .B(n37283), .Z(n37322) );
  AND U38332 ( .A(x[493]), .B(y[8077]), .Z(n38822) );
  NAND U38333 ( .A(n38822), .B(n37397), .Z(n37288) );
  NAND U38334 ( .A(n37286), .B(n37285), .Z(n37287) );
  NAND U38335 ( .A(n37288), .B(n37287), .Z(n37320) );
  NAND U38336 ( .A(y[8067]), .B(x[491]), .Z(n37289) );
  XNOR U38337 ( .A(n37290), .B(n37289), .Z(n37347) );
  AND U38338 ( .A(x[481]), .B(y[8077]), .Z(n37346) );
  XOR U38339 ( .A(n37347), .B(n37346), .Z(n37319) );
  XOR U38340 ( .A(n37320), .B(n37319), .Z(n37321) );
  XOR U38341 ( .A(n37322), .B(n37321), .Z(n37376) );
  XOR U38342 ( .A(n37377), .B(n37376), .Z(n37379) );
  NAND U38343 ( .A(n37292), .B(n37291), .Z(n37296) );
  NAND U38344 ( .A(n37294), .B(n37293), .Z(n37295) );
  AND U38345 ( .A(n37296), .B(n37295), .Z(n37378) );
  XNOR U38346 ( .A(n37379), .B(n37378), .Z(n37307) );
  XOR U38347 ( .A(n37308), .B(n37307), .Z(n37309) );
  XOR U38348 ( .A(n37310), .B(n37309), .Z(n37384) );
  XNOR U38349 ( .A(n37385), .B(n37384), .Z(n37390) );
  NAND U38350 ( .A(n37298), .B(n37297), .Z(n37302) );
  NAND U38351 ( .A(n37300), .B(n37299), .Z(n37301) );
  AND U38352 ( .A(n37302), .B(n37301), .Z(n37388) );
  XNOR U38353 ( .A(n37388), .B(n37389), .Z(n37306) );
  XNOR U38354 ( .A(n37390), .B(n37306), .Z(N815) );
  NAND U38355 ( .A(n37308), .B(n37307), .Z(n37312) );
  NAND U38356 ( .A(n37310), .B(n37309), .Z(n37311) );
  AND U38357 ( .A(n37312), .B(n37311), .Z(n37481) );
  NAND U38358 ( .A(n37314), .B(n37313), .Z(n37318) );
  NAND U38359 ( .A(n37316), .B(n37315), .Z(n37317) );
  NAND U38360 ( .A(n37318), .B(n37317), .Z(n37454) );
  NAND U38361 ( .A(n37320), .B(n37319), .Z(n37324) );
  NANDN U38362 ( .A(n37322), .B(n37321), .Z(n37323) );
  NAND U38363 ( .A(n37324), .B(n37323), .Z(n37459) );
  NAND U38364 ( .A(n37326), .B(n37325), .Z(n37330) );
  NAND U38365 ( .A(n37328), .B(n37327), .Z(n37329) );
  NAND U38366 ( .A(n37330), .B(n37329), .Z(n37457) );
  NAND U38367 ( .A(x[492]), .B(y[8071]), .Z(n37802) );
  NANDN U38368 ( .A(n37802), .B(n37331), .Z(n37335) );
  NAND U38369 ( .A(n37333), .B(n37332), .Z(n37334) );
  AND U38370 ( .A(n37335), .B(n37334), .Z(n37433) );
  AND U38371 ( .A(y[8068]), .B(x[491]), .Z(n37337) );
  NAND U38372 ( .A(y[8066]), .B(x[493]), .Z(n37336) );
  XNOR U38373 ( .A(n37337), .B(n37336), .Z(n37438) );
  AND U38374 ( .A(x[492]), .B(y[8067]), .Z(n37437) );
  XNOR U38375 ( .A(n37438), .B(n37437), .Z(n37432) );
  AND U38376 ( .A(y[8064]), .B(x[495]), .Z(n37339) );
  NAND U38377 ( .A(y[8079]), .B(x[480]), .Z(n37338) );
  XNOR U38378 ( .A(n37339), .B(n37338), .Z(n37399) );
  AND U38379 ( .A(n37340), .B(o[398]), .Z(n37398) );
  XNOR U38380 ( .A(n37399), .B(n37398), .Z(n37431) );
  XNOR U38381 ( .A(n37432), .B(n37431), .Z(n37434) );
  XOR U38382 ( .A(n37433), .B(n37434), .Z(n37465) );
  NAND U38383 ( .A(x[490]), .B(y[8076]), .Z(n38233) );
  NANDN U38384 ( .A(n38233), .B(n37341), .Z(n37344) );
  NAND U38385 ( .A(n37914), .B(n37342), .Z(n37343) );
  NAND U38386 ( .A(n37344), .B(n37343), .Z(n37464) );
  AND U38387 ( .A(x[491]), .B(y[8072]), .Z(n37729) );
  NAND U38388 ( .A(n37729), .B(n37345), .Z(n37349) );
  NAND U38389 ( .A(n37347), .B(n37346), .Z(n37348) );
  NAND U38390 ( .A(n37349), .B(n37348), .Z(n37463) );
  XNOR U38391 ( .A(n37464), .B(n37463), .Z(n37466) );
  XOR U38392 ( .A(n37457), .B(n37458), .Z(n37460) );
  XOR U38393 ( .A(n37459), .B(n37460), .Z(n37451) );
  AND U38394 ( .A(x[494]), .B(y[8078]), .Z(n39076) );
  NAND U38395 ( .A(n39076), .B(n37397), .Z(n37353) );
  NAND U38396 ( .A(n37351), .B(n37350), .Z(n37352) );
  NAND U38397 ( .A(n37353), .B(n37352), .Z(n37426) );
  AND U38398 ( .A(x[488]), .B(y[8075]), .Z(n37354) );
  NAND U38399 ( .A(n37355), .B(n37354), .Z(n37358) );
  NAND U38400 ( .A(n37356), .B(n37625), .Z(n37357) );
  NAND U38401 ( .A(n37358), .B(n37357), .Z(n37425) );
  XOR U38402 ( .A(n37426), .B(n37425), .Z(n37427) );
  AND U38403 ( .A(y[8069]), .B(x[490]), .Z(n37360) );
  NAND U38404 ( .A(y[8075]), .B(x[484]), .Z(n37359) );
  XNOR U38405 ( .A(n37360), .B(n37359), .Z(n37405) );
  AND U38406 ( .A(x[487]), .B(y[8072]), .Z(n37404) );
  XNOR U38407 ( .A(n37405), .B(n37404), .Z(n37413) );
  NAND U38408 ( .A(x[486]), .B(y[8073]), .Z(n37410) );
  XOR U38409 ( .A(n37410), .B(n37411), .Z(n37412) );
  XNOR U38410 ( .A(n37413), .B(n37412), .Z(n37448) );
  AND U38411 ( .A(y[8077]), .B(x[482]), .Z(n37362) );
  NAND U38412 ( .A(y[8070]), .B(x[489]), .Z(n37361) );
  XNOR U38413 ( .A(n37362), .B(n37361), .Z(n37417) );
  AND U38414 ( .A(x[483]), .B(y[8076]), .Z(n37416) );
  XOR U38415 ( .A(n37417), .B(n37416), .Z(n37446) );
  AND U38416 ( .A(y[8078]), .B(x[481]), .Z(n37364) );
  NAND U38417 ( .A(y[8071]), .B(x[488]), .Z(n37363) );
  XNOR U38418 ( .A(n37364), .B(n37363), .Z(n37394) );
  AND U38419 ( .A(x[494]), .B(y[8065]), .Z(n37422) );
  XOR U38420 ( .A(n37422), .B(o[399]), .Z(n37393) );
  XOR U38421 ( .A(n37394), .B(n37393), .Z(n37445) );
  XOR U38422 ( .A(n37446), .B(n37445), .Z(n37447) );
  XNOR U38423 ( .A(n37448), .B(n37447), .Z(n37428) );
  XNOR U38424 ( .A(n37427), .B(n37428), .Z(n37470) );
  NAND U38425 ( .A(n37730), .B(n37365), .Z(n37369) );
  NAND U38426 ( .A(n37367), .B(n37366), .Z(n37368) );
  AND U38427 ( .A(n37369), .B(n37368), .Z(n37469) );
  NAND U38428 ( .A(n37371), .B(n37370), .Z(n37375) );
  NAND U38429 ( .A(n37373), .B(n37372), .Z(n37374) );
  AND U38430 ( .A(n37375), .B(n37374), .Z(n37471) );
  XOR U38431 ( .A(n37472), .B(n37471), .Z(n37452) );
  XOR U38432 ( .A(n37451), .B(n37452), .Z(n37453) );
  XNOR U38433 ( .A(n37454), .B(n37453), .Z(n37478) );
  NAND U38434 ( .A(n37377), .B(n37376), .Z(n37381) );
  NAND U38435 ( .A(n37379), .B(n37378), .Z(n37380) );
  AND U38436 ( .A(n37381), .B(n37380), .Z(n37479) );
  XOR U38437 ( .A(n37478), .B(n37479), .Z(n37480) );
  XOR U38438 ( .A(n37481), .B(n37480), .Z(n37477) );
  NANDN U38439 ( .A(n37383), .B(n37382), .Z(n37387) );
  NAND U38440 ( .A(n37385), .B(n37384), .Z(n37386) );
  NAND U38441 ( .A(n37387), .B(n37386), .Z(n37475) );
  XOR U38442 ( .A(n37475), .B(n37476), .Z(n37391) );
  XNOR U38443 ( .A(n37477), .B(n37391), .Z(N816) );
  AND U38444 ( .A(x[488]), .B(y[8078]), .Z(n37731) );
  NAND U38445 ( .A(n37731), .B(n37392), .Z(n37396) );
  NAND U38446 ( .A(n37394), .B(n37393), .Z(n37395) );
  NAND U38447 ( .A(n37396), .B(n37395), .Z(n37536) );
  AND U38448 ( .A(x[495]), .B(y[8079]), .Z(n39430) );
  NAND U38449 ( .A(n39430), .B(n37397), .Z(n37401) );
  NAND U38450 ( .A(n37399), .B(n37398), .Z(n37400) );
  NAND U38451 ( .A(n37401), .B(n37400), .Z(n37535) );
  XOR U38452 ( .A(n37536), .B(n37535), .Z(n37537) );
  AND U38453 ( .A(x[490]), .B(y[8075]), .Z(n37403) );
  NAND U38454 ( .A(n37403), .B(n37402), .Z(n37407) );
  NAND U38455 ( .A(n37405), .B(n37404), .Z(n37406) );
  NAND U38456 ( .A(n37407), .B(n37406), .Z(n37499) );
  AND U38457 ( .A(x[480]), .B(y[8080]), .Z(n37518) );
  AND U38458 ( .A(x[496]), .B(y[8064]), .Z(n37517) );
  XOR U38459 ( .A(n37518), .B(n37517), .Z(n37520) );
  AND U38460 ( .A(x[495]), .B(y[8065]), .Z(n37509) );
  XOR U38461 ( .A(n37509), .B(o[400]), .Z(n37519) );
  XOR U38462 ( .A(n37520), .B(n37519), .Z(n37498) );
  NAND U38463 ( .A(y[8073]), .B(x[487]), .Z(n37408) );
  XNOR U38464 ( .A(n37409), .B(n37408), .Z(n37514) );
  AND U38465 ( .A(x[490]), .B(y[8070]), .Z(n37513) );
  XOR U38466 ( .A(n37514), .B(n37513), .Z(n37497) );
  XOR U38467 ( .A(n37498), .B(n37497), .Z(n37500) );
  XNOR U38468 ( .A(n37499), .B(n37500), .Z(n37538) );
  IV U38469 ( .A(n37410), .Z(n37512) );
  NANDN U38470 ( .A(n37512), .B(n37411), .Z(n37415) );
  NAND U38471 ( .A(n37413), .B(n37412), .Z(n37414) );
  NAND U38472 ( .A(n37415), .B(n37414), .Z(n37492) );
  AND U38473 ( .A(x[489]), .B(y[8077]), .Z(n38213) );
  NAND U38474 ( .A(n38213), .B(n37800), .Z(n37419) );
  NAND U38475 ( .A(n37417), .B(n37416), .Z(n37418) );
  NAND U38476 ( .A(n37419), .B(n37418), .Z(n37525) );
  AND U38477 ( .A(y[8079]), .B(x[481]), .Z(n37421) );
  NAND U38478 ( .A(y[8072]), .B(x[488]), .Z(n37420) );
  XNOR U38479 ( .A(n37421), .B(n37420), .Z(n37516) );
  AND U38480 ( .A(n37422), .B(o[399]), .Z(n37515) );
  XOR U38481 ( .A(n37516), .B(n37515), .Z(n37524) );
  NAND U38482 ( .A(y[8066]), .B(x[494]), .Z(n37423) );
  XNOR U38483 ( .A(n37424), .B(n37423), .Z(n37547) );
  NAND U38484 ( .A(x[484]), .B(y[8076]), .Z(n37548) );
  XNOR U38485 ( .A(n37547), .B(n37548), .Z(n37523) );
  XOR U38486 ( .A(n37524), .B(n37523), .Z(n37526) );
  XNOR U38487 ( .A(n37525), .B(n37526), .Z(n37491) );
  XOR U38488 ( .A(n37492), .B(n37491), .Z(n37493) );
  XOR U38489 ( .A(n37494), .B(n37493), .Z(n37530) );
  NAND U38490 ( .A(n37426), .B(n37425), .Z(n37430) );
  NANDN U38491 ( .A(n37428), .B(n37427), .Z(n37429) );
  AND U38492 ( .A(n37430), .B(n37429), .Z(n37529) );
  XOR U38493 ( .A(n37530), .B(n37529), .Z(n37532) );
  NAND U38494 ( .A(n37432), .B(n37431), .Z(n37436) );
  NANDN U38495 ( .A(n37434), .B(n37433), .Z(n37435) );
  NAND U38496 ( .A(n37436), .B(n37435), .Z(n37561) );
  AND U38497 ( .A(x[493]), .B(y[8068]), .Z(n37558) );
  NAND U38498 ( .A(n38045), .B(n37558), .Z(n37440) );
  NAND U38499 ( .A(n37438), .B(n37437), .Z(n37439) );
  NAND U38500 ( .A(n37440), .B(n37439), .Z(n37543) );
  AND U38501 ( .A(y[8078]), .B(x[482]), .Z(n37442) );
  NAND U38502 ( .A(y[8071]), .B(x[489]), .Z(n37441) );
  XNOR U38503 ( .A(n37442), .B(n37441), .Z(n37551) );
  NAND U38504 ( .A(x[483]), .B(y[8077]), .Z(n37552) );
  XNOR U38505 ( .A(n37551), .B(n37552), .Z(n37542) );
  AND U38506 ( .A(x[492]), .B(y[8068]), .Z(n38202) );
  AND U38507 ( .A(y[8075]), .B(x[485]), .Z(n37444) );
  NAND U38508 ( .A(y[8067]), .B(x[493]), .Z(n37443) );
  XNOR U38509 ( .A(n37444), .B(n37443), .Z(n37504) );
  XOR U38510 ( .A(n38202), .B(n37504), .Z(n37541) );
  XOR U38511 ( .A(n37542), .B(n37541), .Z(n37544) );
  XNOR U38512 ( .A(n37543), .B(n37544), .Z(n37560) );
  NAND U38513 ( .A(n37446), .B(n37445), .Z(n37450) );
  NAND U38514 ( .A(n37448), .B(n37447), .Z(n37449) );
  AND U38515 ( .A(n37450), .B(n37449), .Z(n37559) );
  XOR U38516 ( .A(n37560), .B(n37559), .Z(n37562) );
  XOR U38517 ( .A(n37561), .B(n37562), .Z(n37531) );
  XNOR U38518 ( .A(n37532), .B(n37531), .Z(n37566) );
  NAND U38519 ( .A(n37452), .B(n37451), .Z(n37456) );
  NAND U38520 ( .A(n37454), .B(n37453), .Z(n37455) );
  AND U38521 ( .A(n37456), .B(n37455), .Z(n37565) );
  XOR U38522 ( .A(n37566), .B(n37565), .Z(n37568) );
  NANDN U38523 ( .A(n37458), .B(n37457), .Z(n37462) );
  NANDN U38524 ( .A(n37460), .B(n37459), .Z(n37461) );
  NAND U38525 ( .A(n37462), .B(n37461), .Z(n37487) );
  NAND U38526 ( .A(n37464), .B(n37463), .Z(n37468) );
  NANDN U38527 ( .A(n37466), .B(n37465), .Z(n37467) );
  NAND U38528 ( .A(n37468), .B(n37467), .Z(n37485) );
  NANDN U38529 ( .A(n37470), .B(n37469), .Z(n37474) );
  NAND U38530 ( .A(n37472), .B(n37471), .Z(n37473) );
  AND U38531 ( .A(n37474), .B(n37473), .Z(n37486) );
  XOR U38532 ( .A(n37485), .B(n37486), .Z(n37488) );
  XOR U38533 ( .A(n37487), .B(n37488), .Z(n37567) );
  XOR U38534 ( .A(n37568), .B(n37567), .Z(n37574) );
  NAND U38535 ( .A(n37479), .B(n37478), .Z(n37483) );
  NANDN U38536 ( .A(n37481), .B(n37480), .Z(n37482) );
  AND U38537 ( .A(n37483), .B(n37482), .Z(n37573) );
  IV U38538 ( .A(n37573), .Z(n37571) );
  XOR U38539 ( .A(n37572), .B(n37571), .Z(n37484) );
  XNOR U38540 ( .A(n37574), .B(n37484), .Z(N817) );
  NAND U38541 ( .A(n37486), .B(n37485), .Z(n37490) );
  NAND U38542 ( .A(n37488), .B(n37487), .Z(n37489) );
  NAND U38543 ( .A(n37490), .B(n37489), .Z(n37665) );
  NAND U38544 ( .A(n37492), .B(n37491), .Z(n37496) );
  NAND U38545 ( .A(n37494), .B(n37493), .Z(n37495) );
  NAND U38546 ( .A(n37496), .B(n37495), .Z(n37587) );
  NAND U38547 ( .A(n37498), .B(n37497), .Z(n37502) );
  NAND U38548 ( .A(n37500), .B(n37499), .Z(n37501) );
  NAND U38549 ( .A(n37502), .B(n37501), .Z(n37659) );
  AND U38550 ( .A(x[493]), .B(y[8075]), .Z(n38491) );
  NAND U38551 ( .A(n38491), .B(n37503), .Z(n37506) );
  NAND U38552 ( .A(n38202), .B(n37504), .Z(n37505) );
  NAND U38553 ( .A(n37506), .B(n37505), .Z(n37615) );
  AND U38554 ( .A(y[8080]), .B(x[481]), .Z(n37508) );
  NAND U38555 ( .A(y[8072]), .B(x[489]), .Z(n37507) );
  XNOR U38556 ( .A(n37508), .B(n37507), .Z(n37630) );
  NAND U38557 ( .A(n37509), .B(o[400]), .Z(n37631) );
  XNOR U38558 ( .A(n37630), .B(n37631), .Z(n37614) );
  AND U38559 ( .A(y[8066]), .B(x[495]), .Z(n37511) );
  NAND U38560 ( .A(y[8069]), .B(x[492]), .Z(n37510) );
  XNOR U38561 ( .A(n37511), .B(n37510), .Z(n37592) );
  AND U38562 ( .A(x[494]), .B(y[8067]), .Z(n37591) );
  XOR U38563 ( .A(n37592), .B(n37591), .Z(n37613) );
  XOR U38564 ( .A(n37614), .B(n37613), .Z(n37616) );
  XOR U38565 ( .A(n37615), .B(n37616), .Z(n37658) );
  NAND U38566 ( .A(x[487]), .B(y[8074]), .Z(n37640) );
  NAND U38567 ( .A(x[488]), .B(y[8079]), .Z(n38296) );
  AND U38568 ( .A(x[481]), .B(y[8072]), .Z(n37709) );
  XOR U38569 ( .A(n37621), .B(n37622), .Z(n37624) );
  AND U38570 ( .A(x[480]), .B(y[8081]), .Z(n37606) );
  AND U38571 ( .A(x[497]), .B(y[8064]), .Z(n37605) );
  XOR U38572 ( .A(n37606), .B(n37605), .Z(n37608) );
  AND U38573 ( .A(x[496]), .B(y[8065]), .Z(n37602) );
  XOR U38574 ( .A(n37602), .B(o[401]), .Z(n37607) );
  XOR U38575 ( .A(n37608), .B(n37607), .Z(n37618) );
  AND U38576 ( .A(y[8079]), .B(x[482]), .Z(n37522) );
  NAND U38577 ( .A(y[8071]), .B(x[490]), .Z(n37521) );
  XNOR U38578 ( .A(n37522), .B(n37521), .Z(n37636) );
  AND U38579 ( .A(x[483]), .B(y[8078]), .Z(n37635) );
  XOR U38580 ( .A(n37636), .B(n37635), .Z(n37617) );
  XOR U38581 ( .A(n37618), .B(n37617), .Z(n37620) );
  XOR U38582 ( .A(n37619), .B(n37620), .Z(n37623) );
  XOR U38583 ( .A(n37624), .B(n37623), .Z(n37657) );
  XOR U38584 ( .A(n37658), .B(n37657), .Z(n37660) );
  XNOR U38585 ( .A(n37659), .B(n37660), .Z(n37586) );
  NAND U38586 ( .A(n37524), .B(n37523), .Z(n37528) );
  NAND U38587 ( .A(n37526), .B(n37525), .Z(n37527) );
  AND U38588 ( .A(n37528), .B(n37527), .Z(n37585) );
  XOR U38589 ( .A(n37586), .B(n37585), .Z(n37588) );
  XOR U38590 ( .A(n37587), .B(n37588), .Z(n37664) );
  NAND U38591 ( .A(n37530), .B(n37529), .Z(n37534) );
  NAND U38592 ( .A(n37532), .B(n37531), .Z(n37533) );
  NAND U38593 ( .A(n37534), .B(n37533), .Z(n37581) );
  NAND U38594 ( .A(n37536), .B(n37535), .Z(n37540) );
  NANDN U38595 ( .A(n37538), .B(n37537), .Z(n37539) );
  NAND U38596 ( .A(n37540), .B(n37539), .Z(n37653) );
  NAND U38597 ( .A(n37542), .B(n37541), .Z(n37546) );
  NAND U38598 ( .A(n37544), .B(n37543), .Z(n37545) );
  NAND U38599 ( .A(n37546), .B(n37545), .Z(n37651) );
  NAND U38600 ( .A(x[494]), .B(y[8069]), .Z(n37834) );
  NANDN U38601 ( .A(n37834), .B(n38045), .Z(n37550) );
  NANDN U38602 ( .A(n37548), .B(n37547), .Z(n37549) );
  AND U38603 ( .A(n37550), .B(n37549), .Z(n37646) );
  AND U38604 ( .A(x[489]), .B(y[8078]), .Z(n38472) );
  NANDN U38605 ( .A(n37634), .B(n38472), .Z(n37554) );
  NANDN U38606 ( .A(n37552), .B(n37551), .Z(n37553) );
  NAND U38607 ( .A(n37554), .B(n37553), .Z(n37645) );
  XNOR U38608 ( .A(n37646), .B(n37645), .Z(n37647) );
  AND U38609 ( .A(x[485]), .B(y[8076]), .Z(n37691) );
  NAND U38610 ( .A(y[8073]), .B(x[488]), .Z(n37555) );
  XNOR U38611 ( .A(n37691), .B(n37555), .Z(n37626) );
  XOR U38612 ( .A(n37626), .B(n37556), .Z(n37639) );
  XNOR U38613 ( .A(n37639), .B(n37640), .Z(n37641) );
  NAND U38614 ( .A(y[8077]), .B(x[484]), .Z(n37557) );
  XNOR U38615 ( .A(n37558), .B(n37557), .Z(n37596) );
  NAND U38616 ( .A(x[491]), .B(y[8070]), .Z(n37597) );
  XOR U38617 ( .A(n37596), .B(n37597), .Z(n37642) );
  XOR U38618 ( .A(n37641), .B(n37642), .Z(n37648) );
  XNOR U38619 ( .A(n37647), .B(n37648), .Z(n37652) );
  XOR U38620 ( .A(n37651), .B(n37652), .Z(n37654) );
  XNOR U38621 ( .A(n37653), .B(n37654), .Z(n37580) );
  NAND U38622 ( .A(n37560), .B(n37559), .Z(n37564) );
  NAND U38623 ( .A(n37562), .B(n37561), .Z(n37563) );
  NAND U38624 ( .A(n37564), .B(n37563), .Z(n37579) );
  XOR U38625 ( .A(n37580), .B(n37579), .Z(n37582) );
  XNOR U38626 ( .A(n37581), .B(n37582), .Z(n37663) );
  XOR U38627 ( .A(n37665), .B(n37666), .Z(n37671) );
  NAND U38628 ( .A(n37566), .B(n37565), .Z(n37570) );
  NAND U38629 ( .A(n37568), .B(n37567), .Z(n37569) );
  NAND U38630 ( .A(n37570), .B(n37569), .Z(n37670) );
  NANDN U38631 ( .A(n37571), .B(n37572), .Z(n37577) );
  NOR U38632 ( .A(n37573), .B(n37572), .Z(n37575) );
  OR U38633 ( .A(n37575), .B(n37574), .Z(n37576) );
  AND U38634 ( .A(n37577), .B(n37576), .Z(n37669) );
  XOR U38635 ( .A(n37670), .B(n37669), .Z(n37578) );
  XNOR U38636 ( .A(n37671), .B(n37578), .Z(N818) );
  NAND U38637 ( .A(n37580), .B(n37579), .Z(n37584) );
  NAND U38638 ( .A(n37582), .B(n37581), .Z(n37583) );
  AND U38639 ( .A(n37584), .B(n37583), .Z(n37773) );
  NAND U38640 ( .A(n37586), .B(n37585), .Z(n37590) );
  NAND U38641 ( .A(n37588), .B(n37587), .Z(n37589) );
  AND U38642 ( .A(n37590), .B(n37589), .Z(n37771) );
  AND U38643 ( .A(x[492]), .B(y[8066]), .Z(n37904) );
  AND U38644 ( .A(x[495]), .B(y[8069]), .Z(n37808) );
  NAND U38645 ( .A(n37904), .B(n37808), .Z(n37594) );
  NAND U38646 ( .A(n37592), .B(n37591), .Z(n37593) );
  NAND U38647 ( .A(n37594), .B(n37593), .Z(n37755) );
  NAND U38648 ( .A(n38822), .B(n37595), .Z(n37599) );
  NANDN U38649 ( .A(n37597), .B(n37596), .Z(n37598) );
  AND U38650 ( .A(n37599), .B(n37598), .Z(n37748) );
  AND U38651 ( .A(y[8081]), .B(x[481]), .Z(n37601) );
  NAND U38652 ( .A(y[8072]), .B(x[490]), .Z(n37600) );
  XNOR U38653 ( .A(n37601), .B(n37600), .Z(n37710) );
  AND U38654 ( .A(n37602), .B(o[401]), .Z(n37711) );
  XOR U38655 ( .A(n37710), .B(n37711), .Z(n37746) );
  AND U38656 ( .A(y[8067]), .B(x[495]), .Z(n37604) );
  NAND U38657 ( .A(y[8073]), .B(x[489]), .Z(n37603) );
  XNOR U38658 ( .A(n37604), .B(n37603), .Z(n37701) );
  AND U38659 ( .A(x[494]), .B(y[8068]), .Z(n37702) );
  XOR U38660 ( .A(n37701), .B(n37702), .Z(n37745) );
  XOR U38661 ( .A(n37746), .B(n37745), .Z(n37747) );
  XOR U38662 ( .A(n37755), .B(n37756), .Z(n37758) );
  AND U38663 ( .A(y[8066]), .B(x[496]), .Z(n37610) );
  NAND U38664 ( .A(y[8071]), .B(x[491]), .Z(n37609) );
  XNOR U38665 ( .A(n37610), .B(n37609), .Z(n37697) );
  NAND U38666 ( .A(x[482]), .B(y[8080]), .Z(n37698) );
  XOR U38667 ( .A(n37763), .B(n37764), .Z(n37766) );
  AND U38668 ( .A(y[8077]), .B(x[485]), .Z(n37816) );
  NAND U38669 ( .A(y[8076]), .B(x[486]), .Z(n37611) );
  XNOR U38670 ( .A(n37816), .B(n37611), .Z(n37694) );
  NAND U38671 ( .A(y[8078]), .B(x[484]), .Z(n37612) );
  XNOR U38672 ( .A(n38477), .B(n37612), .Z(n37732) );
  AND U38673 ( .A(x[487]), .B(y[8075]), .Z(n37733) );
  XOR U38674 ( .A(n37732), .B(n37733), .Z(n37693) );
  XOR U38675 ( .A(n37694), .B(n37693), .Z(n37765) );
  XOR U38676 ( .A(n37766), .B(n37765), .Z(n37757) );
  XOR U38677 ( .A(n37758), .B(n37757), .Z(n37680) );
  XOR U38678 ( .A(n37752), .B(n37751), .Z(n37754) );
  XOR U38679 ( .A(n37754), .B(n37753), .Z(n37679) );
  AND U38680 ( .A(x[488]), .B(y[8076]), .Z(n37944) );
  NAND U38681 ( .A(n37944), .B(n37625), .Z(n37629) );
  NANDN U38682 ( .A(n37627), .B(n37626), .Z(n37628) );
  NAND U38683 ( .A(n37629), .B(n37628), .Z(n37759) );
  NAND U38684 ( .A(x[489]), .B(y[8080]), .Z(n38584) );
  NANDN U38685 ( .A(n38584), .B(n37709), .Z(n37633) );
  NANDN U38686 ( .A(n37631), .B(n37630), .Z(n37632) );
  NAND U38687 ( .A(n37633), .B(n37632), .Z(n37760) );
  XOR U38688 ( .A(n37759), .B(n37760), .Z(n37762) );
  NAND U38689 ( .A(x[490]), .B(y[8079]), .Z(n38583) );
  AND U38690 ( .A(x[480]), .B(y[8082]), .Z(n37714) );
  AND U38691 ( .A(x[498]), .B(y[8064]), .Z(n37715) );
  XOR U38692 ( .A(n37714), .B(n37715), .Z(n37717) );
  AND U38693 ( .A(x[497]), .B(y[8065]), .Z(n37736) );
  XOR U38694 ( .A(o[402]), .B(n37736), .Z(n37716) );
  XOR U38695 ( .A(n37717), .B(n37716), .Z(n37740) );
  AND U38696 ( .A(y[8069]), .B(x[493]), .Z(n37638) );
  NAND U38697 ( .A(y[8079]), .B(x[483]), .Z(n37637) );
  XNOR U38698 ( .A(n37638), .B(n37637), .Z(n37722) );
  AND U38699 ( .A(x[492]), .B(y[8070]), .Z(n37723) );
  XOR U38700 ( .A(n37722), .B(n37723), .Z(n37739) );
  XOR U38701 ( .A(n37740), .B(n37739), .Z(n37741) );
  XOR U38702 ( .A(n37762), .B(n37761), .Z(n37686) );
  NANDN U38703 ( .A(n37640), .B(n37639), .Z(n37644) );
  NANDN U38704 ( .A(n37642), .B(n37641), .Z(n37643) );
  AND U38705 ( .A(n37644), .B(n37643), .Z(n37685) );
  XNOR U38706 ( .A(n37686), .B(n37685), .Z(n37688) );
  NANDN U38707 ( .A(n37646), .B(n37645), .Z(n37650) );
  NANDN U38708 ( .A(n37648), .B(n37647), .Z(n37649) );
  AND U38709 ( .A(n37650), .B(n37649), .Z(n37687) );
  XOR U38710 ( .A(n37688), .B(n37687), .Z(n37681) );
  XOR U38711 ( .A(n37682), .B(n37681), .Z(n37676) );
  NAND U38712 ( .A(n37652), .B(n37651), .Z(n37656) );
  NAND U38713 ( .A(n37654), .B(n37653), .Z(n37655) );
  NAND U38714 ( .A(n37656), .B(n37655), .Z(n37674) );
  NAND U38715 ( .A(n37658), .B(n37657), .Z(n37662) );
  NAND U38716 ( .A(n37660), .B(n37659), .Z(n37661) );
  NAND U38717 ( .A(n37662), .B(n37661), .Z(n37673) );
  XOR U38718 ( .A(n37674), .B(n37673), .Z(n37675) );
  XOR U38719 ( .A(n37771), .B(n37770), .Z(n37772) );
  XOR U38720 ( .A(n37773), .B(n37772), .Z(n37769) );
  NANDN U38721 ( .A(n37664), .B(n37663), .Z(n37668) );
  NANDN U38722 ( .A(n37666), .B(n37665), .Z(n37667) );
  AND U38723 ( .A(n37668), .B(n37667), .Z(n37768) );
  XNOR U38724 ( .A(n37768), .B(n37767), .Z(n37672) );
  XNOR U38725 ( .A(n37769), .B(n37672), .Z(N819) );
  NAND U38726 ( .A(n37674), .B(n37673), .Z(n37678) );
  NANDN U38727 ( .A(n37676), .B(n37675), .Z(n37677) );
  NAND U38728 ( .A(n37678), .B(n37677), .Z(n37884) );
  NANDN U38729 ( .A(n37680), .B(n37679), .Z(n37684) );
  NAND U38730 ( .A(n37682), .B(n37681), .Z(n37683) );
  AND U38731 ( .A(n37684), .B(n37683), .Z(n37883) );
  NANDN U38732 ( .A(n37686), .B(n37685), .Z(n37690) );
  NAND U38733 ( .A(n37688), .B(n37687), .Z(n37689) );
  AND U38734 ( .A(n37690), .B(n37689), .Z(n37780) );
  AND U38735 ( .A(x[486]), .B(y[8077]), .Z(n37692) );
  NAND U38736 ( .A(n37692), .B(n37691), .Z(n37696) );
  NAND U38737 ( .A(n37694), .B(n37693), .Z(n37695) );
  AND U38738 ( .A(n37696), .B(n37695), .Z(n37869) );
  AND U38739 ( .A(x[496]), .B(y[8071]), .Z(n38218) );
  NAND U38740 ( .A(n38218), .B(n38045), .Z(n37700) );
  NANDN U38741 ( .A(n37698), .B(n37697), .Z(n37699) );
  AND U38742 ( .A(n37700), .B(n37699), .Z(n37867) );
  AND U38743 ( .A(x[495]), .B(y[8073]), .Z(n38504) );
  NAND U38744 ( .A(n38504), .B(n37795), .Z(n37704) );
  NAND U38745 ( .A(n37702), .B(n37701), .Z(n37703) );
  NAND U38746 ( .A(n37704), .B(n37703), .Z(n37786) );
  AND U38747 ( .A(y[8082]), .B(x[481]), .Z(n37706) );
  NAND U38748 ( .A(y[8075]), .B(x[488]), .Z(n37705) );
  XNOR U38749 ( .A(n37706), .B(n37705), .Z(n37833) );
  AND U38750 ( .A(y[8070]), .B(x[493]), .Z(n37708) );
  NAND U38751 ( .A(y[8081]), .B(x[482]), .Z(n37707) );
  XNOR U38752 ( .A(n37708), .B(n37707), .Z(n37801) );
  XOR U38753 ( .A(n37784), .B(n37783), .Z(n37785) );
  XOR U38754 ( .A(n37786), .B(n37785), .Z(n37866) );
  AND U38755 ( .A(x[490]), .B(y[8081]), .Z(n38928) );
  IV U38756 ( .A(n38928), .Z(n38795) );
  NANDN U38757 ( .A(n38795), .B(n37709), .Z(n37713) );
  NAND U38758 ( .A(n37711), .B(n37710), .Z(n37712) );
  NAND U38759 ( .A(n37713), .B(n37712), .Z(n37845) );
  NAND U38760 ( .A(n37715), .B(n37714), .Z(n37719) );
  NAND U38761 ( .A(n37717), .B(n37716), .Z(n37718) );
  NAND U38762 ( .A(n37719), .B(n37718), .Z(n37843) );
  AND U38763 ( .A(y[8067]), .B(x[496]), .Z(n38443) );
  NAND U38764 ( .A(y[8074]), .B(x[489]), .Z(n37720) );
  XNOR U38765 ( .A(n38443), .B(n37720), .Z(n37796) );
  NAND U38766 ( .A(x[495]), .B(y[8068]), .Z(n37797) );
  XOR U38767 ( .A(n37843), .B(n37842), .Z(n37844) );
  XNOR U38768 ( .A(n37845), .B(n37844), .Z(n37862) );
  AND U38769 ( .A(x[493]), .B(y[8079]), .Z(n39094) );
  NANDN U38770 ( .A(n37721), .B(n39094), .Z(n37725) );
  NAND U38771 ( .A(n37723), .B(n37722), .Z(n37724) );
  NAND U38772 ( .A(n37725), .B(n37724), .Z(n37851) );
  AND U38773 ( .A(y[8073]), .B(x[490]), .Z(n37727) );
  NAND U38774 ( .A(y[8066]), .B(x[497]), .Z(n37726) );
  XNOR U38775 ( .A(n37727), .B(n37726), .Z(n37839) );
  AND U38776 ( .A(x[498]), .B(y[8065]), .Z(n37815) );
  XOR U38777 ( .A(o[403]), .B(n37815), .Z(n37838) );
  XOR U38778 ( .A(n37839), .B(n37838), .Z(n37849) );
  NAND U38779 ( .A(y[8080]), .B(x[483]), .Z(n37728) );
  XNOR U38780 ( .A(n37729), .B(n37728), .Z(n37809) );
  XOR U38781 ( .A(n37849), .B(n37848), .Z(n37850) );
  XNOR U38782 ( .A(n37851), .B(n37850), .Z(n37861) );
  NAND U38783 ( .A(n37731), .B(n37730), .Z(n37735) );
  NAND U38784 ( .A(n37733), .B(n37732), .Z(n37734) );
  AND U38785 ( .A(n37735), .B(n37734), .Z(n37792) );
  AND U38786 ( .A(x[480]), .B(y[8083]), .Z(n37820) );
  AND U38787 ( .A(x[499]), .B(y[8064]), .Z(n37821) );
  XOR U38788 ( .A(n37820), .B(n37821), .Z(n37823) );
  AND U38789 ( .A(o[402]), .B(n37736), .Z(n37822) );
  XOR U38790 ( .A(n37823), .B(n37822), .Z(n37790) );
  AND U38791 ( .A(x[484]), .B(y[8079]), .Z(n37958) );
  AND U38792 ( .A(y[8078]), .B(x[485]), .Z(n37738) );
  NAND U38793 ( .A(y[8077]), .B(x[486]), .Z(n37737) );
  XNOR U38794 ( .A(n37738), .B(n37737), .Z(n37817) );
  XOR U38795 ( .A(n37958), .B(n37817), .Z(n37789) );
  XOR U38796 ( .A(n37790), .B(n37789), .Z(n37791) );
  XOR U38797 ( .A(n37792), .B(n37791), .Z(n37860) );
  XOR U38798 ( .A(n37861), .B(n37860), .Z(n37863) );
  XNOR U38799 ( .A(n37862), .B(n37863), .Z(n37856) );
  NAND U38800 ( .A(n37740), .B(n37739), .Z(n37744) );
  NANDN U38801 ( .A(n37742), .B(n37741), .Z(n37743) );
  AND U38802 ( .A(n37744), .B(n37743), .Z(n37855) );
  NAND U38803 ( .A(n37746), .B(n37745), .Z(n37750) );
  NANDN U38804 ( .A(n37748), .B(n37747), .Z(n37749) );
  NAND U38805 ( .A(n37750), .B(n37749), .Z(n37854) );
  XNOR U38806 ( .A(n37856), .B(n37857), .Z(n37777) );
  XOR U38807 ( .A(n37778), .B(n37777), .Z(n37779) );
  XNOR U38808 ( .A(n37872), .B(n37873), .Z(n37875) );
  XOR U38809 ( .A(n37874), .B(n37875), .Z(n37877) );
  XNOR U38810 ( .A(n37876), .B(n37877), .Z(n37878) );
  XNOR U38811 ( .A(n37879), .B(n37878), .Z(n37882) );
  XOR U38812 ( .A(n37883), .B(n37882), .Z(n37885) );
  XNOR U38813 ( .A(n37884), .B(n37885), .Z(n37890) );
  NAND U38814 ( .A(n37771), .B(n37770), .Z(n37775) );
  NAND U38815 ( .A(n37773), .B(n37772), .Z(n37774) );
  NAND U38816 ( .A(n37775), .B(n37774), .Z(n37889) );
  XOR U38817 ( .A(n37888), .B(n37889), .Z(n37776) );
  XNOR U38818 ( .A(n37890), .B(n37776), .Z(N820) );
  NAND U38819 ( .A(n37778), .B(n37777), .Z(n37782) );
  NANDN U38820 ( .A(n37780), .B(n37779), .Z(n37781) );
  AND U38821 ( .A(n37782), .B(n37781), .Z(n37996) );
  NAND U38822 ( .A(n37784), .B(n37783), .Z(n37788) );
  NAND U38823 ( .A(n37786), .B(n37785), .Z(n37787) );
  NAND U38824 ( .A(n37788), .B(n37787), .Z(n37893) );
  NAND U38825 ( .A(n37790), .B(n37789), .Z(n37794) );
  NANDN U38826 ( .A(n37792), .B(n37791), .Z(n37793) );
  NAND U38827 ( .A(n37794), .B(n37793), .Z(n37892) );
  XOR U38828 ( .A(n37893), .B(n37892), .Z(n37895) );
  AND U38829 ( .A(x[496]), .B(y[8074]), .Z(n38747) );
  NAND U38830 ( .A(n38747), .B(n37795), .Z(n37799) );
  NANDN U38831 ( .A(n37797), .B(n37796), .Z(n37798) );
  AND U38832 ( .A(n37799), .B(n37798), .Z(n37933) );
  AND U38833 ( .A(x[493]), .B(y[8081]), .Z(n39303) );
  NAND U38834 ( .A(n39303), .B(n37800), .Z(n37804) );
  NANDN U38835 ( .A(n37802), .B(n37801), .Z(n37803) );
  AND U38836 ( .A(n37804), .B(n37803), .Z(n37978) );
  AND U38837 ( .A(y[8068]), .B(x[496]), .Z(n37806) );
  NAND U38838 ( .A(y[8074]), .B(x[490]), .Z(n37805) );
  XNOR U38839 ( .A(n37806), .B(n37805), .Z(n37939) );
  AND U38840 ( .A(x[482]), .B(y[8082]), .Z(n37940) );
  XOR U38841 ( .A(n37939), .B(n37940), .Z(n37976) );
  NAND U38842 ( .A(y[8075]), .B(x[489]), .Z(n37807) );
  XNOR U38843 ( .A(n37808), .B(n37807), .Z(n37915) );
  AND U38844 ( .A(x[494]), .B(y[8070]), .Z(n37916) );
  XOR U38845 ( .A(n37915), .B(n37916), .Z(n37975) );
  XOR U38846 ( .A(n37976), .B(n37975), .Z(n37977) );
  NAND U38847 ( .A(x[491]), .B(y[8080]), .Z(n38929) );
  NANDN U38848 ( .A(n38929), .B(n38084), .Z(n37812) );
  NANDN U38849 ( .A(n37810), .B(n37809), .Z(n37811) );
  AND U38850 ( .A(n37812), .B(n37811), .Z(n37984) );
  AND U38851 ( .A(y[8073]), .B(x[491]), .Z(n37814) );
  NAND U38852 ( .A(y[8083]), .B(x[481]), .Z(n37813) );
  XNOR U38853 ( .A(n37814), .B(n37813), .Z(n37911) );
  AND U38854 ( .A(x[499]), .B(y[8065]), .Z(n37919) );
  XOR U38855 ( .A(o[404]), .B(n37919), .Z(n37910) );
  XOR U38856 ( .A(n37911), .B(n37910), .Z(n37982) );
  AND U38857 ( .A(x[480]), .B(y[8084]), .Z(n37963) );
  AND U38858 ( .A(x[500]), .B(y[8064]), .Z(n37964) );
  XOR U38859 ( .A(n37963), .B(n37964), .Z(n37966) );
  AND U38860 ( .A(o[403]), .B(n37815), .Z(n37965) );
  XOR U38861 ( .A(n37966), .B(n37965), .Z(n37981) );
  XOR U38862 ( .A(n37982), .B(n37981), .Z(n37983) );
  XOR U38863 ( .A(n37935), .B(n37934), .Z(n37894) );
  XNOR U38864 ( .A(n37895), .B(n37894), .Z(n37990) );
  NAND U38865 ( .A(x[486]), .B(y[8078]), .Z(n37899) );
  NANDN U38866 ( .A(n37899), .B(n37816), .Z(n37819) );
  NAND U38867 ( .A(n37817), .B(n37958), .Z(n37818) );
  NAND U38868 ( .A(n37819), .B(n37818), .Z(n37923) );
  NAND U38869 ( .A(n37821), .B(n37820), .Z(n37825) );
  NAND U38870 ( .A(n37823), .B(n37822), .Z(n37824) );
  NAND U38871 ( .A(n37825), .B(n37824), .Z(n37921) );
  AND U38872 ( .A(y[8066]), .B(x[498]), .Z(n37827) );
  NAND U38873 ( .A(y[8072]), .B(x[492]), .Z(n37826) );
  XNOR U38874 ( .A(n37827), .B(n37826), .Z(n37905) );
  AND U38875 ( .A(x[497]), .B(y[8067]), .Z(n37906) );
  XOR U38876 ( .A(n37905), .B(n37906), .Z(n37920) );
  XOR U38877 ( .A(n37921), .B(n37920), .Z(n37922) );
  XNOR U38878 ( .A(n37923), .B(n37922), .Z(n37927) );
  AND U38879 ( .A(y[8071]), .B(x[493]), .Z(n37829) );
  NAND U38880 ( .A(y[8081]), .B(x[483]), .Z(n37828) );
  XNOR U38881 ( .A(n37829), .B(n37828), .Z(n37945) );
  XNOR U38882 ( .A(n37945), .B(n37944), .Z(n37901) );
  AND U38883 ( .A(y[8079]), .B(x[485]), .Z(n37831) );
  NAND U38884 ( .A(y[8080]), .B(x[484]), .Z(n37830) );
  XNOR U38885 ( .A(n37831), .B(n37830), .Z(n37960) );
  AND U38886 ( .A(x[487]), .B(y[8077]), .Z(n37959) );
  XNOR U38887 ( .A(n37960), .B(n37959), .Z(n37898) );
  XOR U38888 ( .A(n37899), .B(n37898), .Z(n37900) );
  XNOR U38889 ( .A(n37901), .B(n37900), .Z(n37971) );
  AND U38890 ( .A(x[488]), .B(y[8082]), .Z(n39060) );
  AND U38891 ( .A(x[481]), .B(y[8075]), .Z(n37832) );
  NAND U38892 ( .A(n39060), .B(n37832), .Z(n37836) );
  NANDN U38893 ( .A(n37834), .B(n37833), .Z(n37835) );
  AND U38894 ( .A(n37836), .B(n37835), .Z(n37970) );
  NAND U38895 ( .A(x[497]), .B(y[8073]), .Z(n38756) );
  NANDN U38896 ( .A(n38756), .B(n37837), .Z(n37841) );
  NAND U38897 ( .A(n37839), .B(n37838), .Z(n37840) );
  NAND U38898 ( .A(n37841), .B(n37840), .Z(n37969) );
  XNOR U38899 ( .A(n37971), .B(n37972), .Z(n37926) );
  XOR U38900 ( .A(n37927), .B(n37926), .Z(n37928) );
  NAND U38901 ( .A(n37843), .B(n37842), .Z(n37847) );
  NAND U38902 ( .A(n37845), .B(n37844), .Z(n37846) );
  AND U38903 ( .A(n37847), .B(n37846), .Z(n37929) );
  XOR U38904 ( .A(n37928), .B(n37929), .Z(n37987) );
  NAND U38905 ( .A(n37849), .B(n37848), .Z(n37853) );
  NAND U38906 ( .A(n37851), .B(n37850), .Z(n37852) );
  AND U38907 ( .A(n37853), .B(n37852), .Z(n37988) );
  XOR U38908 ( .A(n37987), .B(n37988), .Z(n37989) );
  XNOR U38909 ( .A(n37990), .B(n37989), .Z(n37994) );
  NANDN U38910 ( .A(n37855), .B(n37854), .Z(n37859) );
  NAND U38911 ( .A(n37857), .B(n37856), .Z(n37858) );
  AND U38912 ( .A(n37859), .B(n37858), .Z(n38002) );
  NAND U38913 ( .A(n37861), .B(n37860), .Z(n37865) );
  NAND U38914 ( .A(n37863), .B(n37862), .Z(n37864) );
  AND U38915 ( .A(n37865), .B(n37864), .Z(n38000) );
  NANDN U38916 ( .A(n37867), .B(n37866), .Z(n37871) );
  NANDN U38917 ( .A(n37869), .B(n37868), .Z(n37870) );
  AND U38918 ( .A(n37871), .B(n37870), .Z(n37999) );
  XNOR U38919 ( .A(n38002), .B(n38001), .Z(n37993) );
  XOR U38920 ( .A(n37994), .B(n37993), .Z(n37995) );
  XOR U38921 ( .A(n37996), .B(n37995), .Z(n38011) );
  NANDN U38922 ( .A(n37877), .B(n37876), .Z(n37881) );
  NANDN U38923 ( .A(n37879), .B(n37878), .Z(n37880) );
  AND U38924 ( .A(n37881), .B(n37880), .Z(n38008) );
  XOR U38925 ( .A(n38009), .B(n38008), .Z(n38010) );
  XOR U38926 ( .A(n38011), .B(n38010), .Z(n38007) );
  NAND U38927 ( .A(n37883), .B(n37882), .Z(n37887) );
  NAND U38928 ( .A(n37885), .B(n37884), .Z(n37886) );
  AND U38929 ( .A(n37887), .B(n37886), .Z(n38006) );
  XNOR U38930 ( .A(n38006), .B(n38005), .Z(n37891) );
  XNOR U38931 ( .A(n38007), .B(n37891), .Z(N821) );
  NAND U38932 ( .A(n37893), .B(n37892), .Z(n37897) );
  NAND U38933 ( .A(n37895), .B(n37894), .Z(n37896) );
  NAND U38934 ( .A(n37897), .B(n37896), .Z(n38024) );
  NAND U38935 ( .A(n37899), .B(n37898), .Z(n37903) );
  NAND U38936 ( .A(n37901), .B(n37900), .Z(n37902) );
  AND U38937 ( .A(n37903), .B(n37902), .Z(n38125) );
  AND U38938 ( .A(x[498]), .B(y[8072]), .Z(n38754) );
  NAND U38939 ( .A(n38754), .B(n37904), .Z(n37908) );
  NAND U38940 ( .A(n37906), .B(n37905), .Z(n37907) );
  NAND U38941 ( .A(n37908), .B(n37907), .Z(n38107) );
  AND U38942 ( .A(x[491]), .B(y[8083]), .Z(n39479) );
  AND U38943 ( .A(x[481]), .B(y[8073]), .Z(n37909) );
  NAND U38944 ( .A(n39479), .B(n37909), .Z(n37913) );
  NAND U38945 ( .A(n37911), .B(n37910), .Z(n37912) );
  NAND U38946 ( .A(n37913), .B(n37912), .Z(n38106) );
  XOR U38947 ( .A(n38107), .B(n38106), .Z(n38109) );
  AND U38948 ( .A(x[495]), .B(y[8075]), .Z(n38742) );
  NAND U38949 ( .A(n38742), .B(n37914), .Z(n37918) );
  NAND U38950 ( .A(n37916), .B(n37915), .Z(n37917) );
  NAND U38951 ( .A(n37918), .B(n37917), .Z(n38070) );
  AND U38952 ( .A(x[480]), .B(y[8085]), .Z(n38090) );
  AND U38953 ( .A(x[501]), .B(y[8064]), .Z(n38091) );
  XOR U38954 ( .A(n38090), .B(n38091), .Z(n38093) );
  AND U38955 ( .A(o[404]), .B(n37919), .Z(n38092) );
  XOR U38956 ( .A(n38093), .B(n38092), .Z(n38069) );
  AND U38957 ( .A(x[485]), .B(y[8080]), .Z(n38077) );
  AND U38958 ( .A(x[496]), .B(y[8069]), .Z(n38076) );
  XOR U38959 ( .A(n38077), .B(n38076), .Z(n38075) );
  AND U38960 ( .A(x[495]), .B(y[8070]), .Z(n38074) );
  XOR U38961 ( .A(n38075), .B(n38074), .Z(n38068) );
  XOR U38962 ( .A(n38069), .B(n38068), .Z(n38071) );
  XOR U38963 ( .A(n38070), .B(n38071), .Z(n38108) );
  XNOR U38964 ( .A(n38109), .B(n38108), .Z(n38124) );
  NAND U38965 ( .A(n37921), .B(n37920), .Z(n37925) );
  NAND U38966 ( .A(n37923), .B(n37922), .Z(n37924) );
  AND U38967 ( .A(n37925), .B(n37924), .Z(n38126) );
  XNOR U38968 ( .A(n38127), .B(n38126), .Z(n38022) );
  NAND U38969 ( .A(n37927), .B(n37926), .Z(n37931) );
  NAND U38970 ( .A(n37929), .B(n37928), .Z(n37930) );
  AND U38971 ( .A(n37931), .B(n37930), .Z(n38021) );
  XOR U38972 ( .A(n38022), .B(n38021), .Z(n38023) );
  XNOR U38973 ( .A(n38024), .B(n38023), .Z(n38017) );
  NANDN U38974 ( .A(n37933), .B(n37932), .Z(n37937) );
  NAND U38975 ( .A(n37935), .B(n37934), .Z(n37936) );
  NAND U38976 ( .A(n37937), .B(n37936), .Z(n38030) );
  NAND U38977 ( .A(n38747), .B(n37938), .Z(n37942) );
  NAND U38978 ( .A(n37940), .B(n37939), .Z(n37941) );
  NAND U38979 ( .A(n37942), .B(n37941), .Z(n38040) );
  NAND U38980 ( .A(n39303), .B(n37943), .Z(n37947) );
  NAND U38981 ( .A(n37945), .B(n37944), .Z(n37946) );
  NAND U38982 ( .A(n37947), .B(n37946), .Z(n38121) );
  AND U38983 ( .A(y[8066]), .B(x[499]), .Z(n37949) );
  NAND U38984 ( .A(y[8074]), .B(x[491]), .Z(n37948) );
  XNOR U38985 ( .A(n37949), .B(n37948), .Z(n38047) );
  AND U38986 ( .A(x[500]), .B(y[8065]), .Z(n38089) );
  XOR U38987 ( .A(n38089), .B(o[405]), .Z(n38046) );
  XOR U38988 ( .A(n38047), .B(n38046), .Z(n38119) );
  AND U38989 ( .A(y[8067]), .B(x[498]), .Z(n37951) );
  NAND U38990 ( .A(y[8075]), .B(x[490]), .Z(n37950) );
  XNOR U38991 ( .A(n37951), .B(n37950), .Z(n38097) );
  AND U38992 ( .A(x[481]), .B(y[8084]), .Z(n38098) );
  XOR U38993 ( .A(n38097), .B(n38098), .Z(n38118) );
  XOR U38994 ( .A(n38119), .B(n38118), .Z(n38120) );
  XOR U38995 ( .A(n38121), .B(n38120), .Z(n38039) );
  XOR U38996 ( .A(n38040), .B(n38039), .Z(n38042) );
  AND U38997 ( .A(x[487]), .B(y[8078]), .Z(n38294) );
  AND U38998 ( .A(y[8079]), .B(x[486]), .Z(n37953) );
  NAND U38999 ( .A(y[8071]), .B(x[494]), .Z(n37952) );
  XNOR U39000 ( .A(n37953), .B(n37952), .Z(n38101) );
  XOR U39001 ( .A(n38294), .B(n38101), .Z(n38059) );
  NAND U39002 ( .A(x[489]), .B(y[8076]), .Z(n38057) );
  NAND U39003 ( .A(x[488]), .B(y[8077]), .Z(n38056) );
  XOR U39004 ( .A(n38057), .B(n38056), .Z(n38058) );
  AND U39005 ( .A(y[8073]), .B(x[492]), .Z(n37955) );
  NAND U39006 ( .A(y[8068]), .B(x[497]), .Z(n37954) );
  XNOR U39007 ( .A(n37955), .B(n37954), .Z(n38050) );
  AND U39008 ( .A(x[482]), .B(y[8083]), .Z(n38051) );
  XOR U39009 ( .A(n38050), .B(n38051), .Z(n38063) );
  AND U39010 ( .A(y[8072]), .B(x[493]), .Z(n37957) );
  NAND U39011 ( .A(y[8082]), .B(x[483]), .Z(n37956) );
  XNOR U39012 ( .A(n37957), .B(n37956), .Z(n38086) );
  AND U39013 ( .A(x[484]), .B(y[8081]), .Z(n38085) );
  XOR U39014 ( .A(n38086), .B(n38085), .Z(n38062) );
  XOR U39015 ( .A(n38063), .B(n38062), .Z(n38064) );
  NAND U39016 ( .A(n38077), .B(n37958), .Z(n37962) );
  NAND U39017 ( .A(n37960), .B(n37959), .Z(n37961) );
  NAND U39018 ( .A(n37962), .B(n37961), .Z(n38113) );
  NAND U39019 ( .A(n37964), .B(n37963), .Z(n37968) );
  NAND U39020 ( .A(n37966), .B(n37965), .Z(n37967) );
  NAND U39021 ( .A(n37968), .B(n37967), .Z(n38112) );
  XOR U39022 ( .A(n38113), .B(n38112), .Z(n38114) );
  XOR U39023 ( .A(n38115), .B(n38114), .Z(n38041) );
  XOR U39024 ( .A(n38042), .B(n38041), .Z(n38028) );
  NANDN U39025 ( .A(n37970), .B(n37969), .Z(n37974) );
  NAND U39026 ( .A(n37972), .B(n37971), .Z(n37973) );
  NAND U39027 ( .A(n37974), .B(n37973), .Z(n38035) );
  NAND U39028 ( .A(n37976), .B(n37975), .Z(n37980) );
  NANDN U39029 ( .A(n37978), .B(n37977), .Z(n37979) );
  NAND U39030 ( .A(n37980), .B(n37979), .Z(n38034) );
  NAND U39031 ( .A(n37982), .B(n37981), .Z(n37986) );
  NANDN U39032 ( .A(n37984), .B(n37983), .Z(n37985) );
  NAND U39033 ( .A(n37986), .B(n37985), .Z(n38033) );
  XOR U39034 ( .A(n38034), .B(n38033), .Z(n38036) );
  XOR U39035 ( .A(n38035), .B(n38036), .Z(n38027) );
  XOR U39036 ( .A(n38028), .B(n38027), .Z(n38029) );
  XNOR U39037 ( .A(n38030), .B(n38029), .Z(n38016) );
  NAND U39038 ( .A(n37988), .B(n37987), .Z(n37992) );
  NAND U39039 ( .A(n37990), .B(n37989), .Z(n37991) );
  NAND U39040 ( .A(n37992), .B(n37991), .Z(n38015) );
  XOR U39041 ( .A(n38016), .B(n38015), .Z(n38018) );
  XNOR U39042 ( .A(n38017), .B(n38018), .Z(n38135) );
  NAND U39043 ( .A(n37994), .B(n37993), .Z(n37998) );
  NAND U39044 ( .A(n37996), .B(n37995), .Z(n37997) );
  AND U39045 ( .A(n37998), .B(n37997), .Z(n38134) );
  NANDN U39046 ( .A(n38000), .B(n37999), .Z(n38004) );
  NAND U39047 ( .A(n38002), .B(n38001), .Z(n38003) );
  AND U39048 ( .A(n38004), .B(n38003), .Z(n38133) );
  XNOR U39049 ( .A(n38135), .B(n38136), .Z(n38132) );
  NAND U39050 ( .A(n38009), .B(n38008), .Z(n38013) );
  NANDN U39051 ( .A(n38011), .B(n38010), .Z(n38012) );
  AND U39052 ( .A(n38013), .B(n38012), .Z(n38131) );
  XOR U39053 ( .A(n38130), .B(n38131), .Z(n38014) );
  XNOR U39054 ( .A(n38132), .B(n38014), .Z(N822) );
  NAND U39055 ( .A(n38016), .B(n38015), .Z(n38020) );
  NAND U39056 ( .A(n38018), .B(n38017), .Z(n38019) );
  AND U39057 ( .A(n38020), .B(n38019), .Z(n38270) );
  NAND U39058 ( .A(n38022), .B(n38021), .Z(n38026) );
  NAND U39059 ( .A(n38024), .B(n38023), .Z(n38025) );
  NAND U39060 ( .A(n38026), .B(n38025), .Z(n38268) );
  NAND U39061 ( .A(n38028), .B(n38027), .Z(n38032) );
  NAND U39062 ( .A(n38030), .B(n38029), .Z(n38031) );
  AND U39063 ( .A(n38032), .B(n38031), .Z(n38141) );
  NAND U39064 ( .A(n38034), .B(n38033), .Z(n38038) );
  NAND U39065 ( .A(n38036), .B(n38035), .Z(n38037) );
  NAND U39066 ( .A(n38038), .B(n38037), .Z(n38140) );
  NAND U39067 ( .A(n38040), .B(n38039), .Z(n38044) );
  NAND U39068 ( .A(n38042), .B(n38041), .Z(n38043) );
  AND U39069 ( .A(n38044), .B(n38043), .Z(n38257) );
  AND U39070 ( .A(x[499]), .B(y[8074]), .Z(n39210) );
  NAND U39071 ( .A(n39210), .B(n38045), .Z(n38049) );
  NAND U39072 ( .A(n38047), .B(n38046), .Z(n38048) );
  NAND U39073 ( .A(n38049), .B(n38048), .Z(n38249) );
  NANDN U39074 ( .A(n38756), .B(n38202), .Z(n38053) );
  NAND U39075 ( .A(n38051), .B(n38050), .Z(n38052) );
  NAND U39076 ( .A(n38053), .B(n38052), .Z(n38179) );
  AND U39077 ( .A(x[485]), .B(y[8081]), .Z(n38224) );
  AND U39078 ( .A(x[497]), .B(y[8069]), .Z(n38225) );
  XOR U39079 ( .A(n38224), .B(n38225), .Z(n38226) );
  AND U39080 ( .A(x[496]), .B(y[8070]), .Z(n38227) );
  XOR U39081 ( .A(n38226), .B(n38227), .Z(n38177) );
  AND U39082 ( .A(y[8068]), .B(x[498]), .Z(n38055) );
  NAND U39083 ( .A(y[8074]), .B(x[492]), .Z(n38054) );
  XNOR U39084 ( .A(n38055), .B(n38054), .Z(n38203) );
  AND U39085 ( .A(x[484]), .B(y[8082]), .Z(n38204) );
  XOR U39086 ( .A(n38203), .B(n38204), .Z(n38176) );
  XOR U39087 ( .A(n38177), .B(n38176), .Z(n38178) );
  XOR U39088 ( .A(n38179), .B(n38178), .Z(n38248) );
  XOR U39089 ( .A(n38249), .B(n38248), .Z(n38251) );
  NAND U39090 ( .A(n38057), .B(n38056), .Z(n38061) );
  NANDN U39091 ( .A(n38059), .B(n38058), .Z(n38060) );
  AND U39092 ( .A(n38061), .B(n38060), .Z(n38250) );
  XNOR U39093 ( .A(n38251), .B(n38250), .Z(n38255) );
  NAND U39094 ( .A(n38063), .B(n38062), .Z(n38067) );
  NANDN U39095 ( .A(n38065), .B(n38064), .Z(n38066) );
  NAND U39096 ( .A(n38067), .B(n38066), .Z(n38237) );
  NAND U39097 ( .A(n38069), .B(n38068), .Z(n38073) );
  NAND U39098 ( .A(n38071), .B(n38070), .Z(n38072) );
  NAND U39099 ( .A(n38073), .B(n38072), .Z(n38236) );
  XOR U39100 ( .A(n38237), .B(n38236), .Z(n38239) );
  AND U39101 ( .A(n38075), .B(n38074), .Z(n38079) );
  NAND U39102 ( .A(n38077), .B(n38076), .Z(n38078) );
  NANDN U39103 ( .A(n38079), .B(n38078), .Z(n38199) );
  AND U39104 ( .A(y[8073]), .B(x[493]), .Z(n38081) );
  NAND U39105 ( .A(y[8066]), .B(x[500]), .Z(n38080) );
  XNOR U39106 ( .A(n38081), .B(n38080), .Z(n38220) );
  AND U39107 ( .A(x[482]), .B(y[8084]), .Z(n38221) );
  XOR U39108 ( .A(n38220), .B(n38221), .Z(n38197) );
  AND U39109 ( .A(y[8080]), .B(x[486]), .Z(n38083) );
  NAND U39110 ( .A(y[8071]), .B(x[495]), .Z(n38082) );
  XNOR U39111 ( .A(n38083), .B(n38082), .Z(n38232) );
  XOR U39112 ( .A(n38197), .B(n38196), .Z(n38198) );
  XOR U39113 ( .A(n38199), .B(n38198), .Z(n38243) );
  AND U39114 ( .A(x[493]), .B(y[8082]), .Z(n39480) );
  NAND U39115 ( .A(n38084), .B(n39480), .Z(n38088) );
  NAND U39116 ( .A(n38086), .B(n38085), .Z(n38087) );
  NAND U39117 ( .A(n38088), .B(n38087), .Z(n38167) );
  AND U39118 ( .A(x[481]), .B(y[8085]), .Z(n38190) );
  XOR U39119 ( .A(n38191), .B(n38190), .Z(n38189) );
  AND U39120 ( .A(n38089), .B(o[405]), .Z(n38188) );
  XOR U39121 ( .A(n38189), .B(n38188), .Z(n38165) );
  AND U39122 ( .A(x[494]), .B(y[8072]), .Z(n38182) );
  AND U39123 ( .A(x[483]), .B(y[8083]), .Z(n38183) );
  XOR U39124 ( .A(n38182), .B(n38183), .Z(n38184) );
  AND U39125 ( .A(x[499]), .B(y[8067]), .Z(n38185) );
  XOR U39126 ( .A(n38184), .B(n38185), .Z(n38164) );
  XOR U39127 ( .A(n38165), .B(n38164), .Z(n38166) );
  XOR U39128 ( .A(n38167), .B(n38166), .Z(n38242) );
  XOR U39129 ( .A(n38243), .B(n38242), .Z(n38245) );
  NAND U39130 ( .A(n38091), .B(n38090), .Z(n38095) );
  NAND U39131 ( .A(n38093), .B(n38092), .Z(n38094) );
  NAND U39132 ( .A(n38095), .B(n38094), .Z(n38159) );
  AND U39133 ( .A(x[498]), .B(y[8075]), .Z(n39213) );
  NAND U39134 ( .A(n39213), .B(n38096), .Z(n38100) );
  NAND U39135 ( .A(n38098), .B(n38097), .Z(n38099) );
  NAND U39136 ( .A(n38100), .B(n38099), .Z(n38158) );
  XOR U39137 ( .A(n38159), .B(n38158), .Z(n38161) );
  AND U39138 ( .A(x[494]), .B(y[8079]), .Z(n39249) );
  NAND U39139 ( .A(n39249), .B(n38231), .Z(n38103) );
  NAND U39140 ( .A(n38101), .B(n38294), .Z(n38102) );
  NAND U39141 ( .A(n38103), .B(n38102), .Z(n38172) );
  AND U39142 ( .A(x[480]), .B(y[8086]), .Z(n38207) );
  AND U39143 ( .A(x[502]), .B(y[8064]), .Z(n38208) );
  XOR U39144 ( .A(n38207), .B(n38208), .Z(n38210) );
  AND U39145 ( .A(x[501]), .B(y[8065]), .Z(n38230) );
  XOR U39146 ( .A(o[406]), .B(n38230), .Z(n38209) );
  XOR U39147 ( .A(n38210), .B(n38209), .Z(n38171) );
  AND U39148 ( .A(y[8079]), .B(x[487]), .Z(n38105) );
  NAND U39149 ( .A(y[8078]), .B(x[488]), .Z(n38104) );
  XNOR U39150 ( .A(n38105), .B(n38104), .Z(n38214) );
  XOR U39151 ( .A(n38214), .B(n38213), .Z(n38170) );
  XOR U39152 ( .A(n38171), .B(n38170), .Z(n38173) );
  XOR U39153 ( .A(n38172), .B(n38173), .Z(n38160) );
  XOR U39154 ( .A(n38161), .B(n38160), .Z(n38244) );
  XOR U39155 ( .A(n38245), .B(n38244), .Z(n38238) );
  XNOR U39156 ( .A(n38239), .B(n38238), .Z(n38254) );
  XOR U39157 ( .A(n38255), .B(n38254), .Z(n38256) );
  XOR U39158 ( .A(n38257), .B(n38256), .Z(n38149) );
  NAND U39159 ( .A(n38107), .B(n38106), .Z(n38111) );
  NAND U39160 ( .A(n38109), .B(n38108), .Z(n38110) );
  NAND U39161 ( .A(n38111), .B(n38110), .Z(n38155) );
  NAND U39162 ( .A(n38113), .B(n38112), .Z(n38117) );
  NAND U39163 ( .A(n38115), .B(n38114), .Z(n38116) );
  NAND U39164 ( .A(n38117), .B(n38116), .Z(n38153) );
  NAND U39165 ( .A(n38119), .B(n38118), .Z(n38123) );
  NAND U39166 ( .A(n38121), .B(n38120), .Z(n38122) );
  NAND U39167 ( .A(n38123), .B(n38122), .Z(n38152) );
  XOR U39168 ( .A(n38153), .B(n38152), .Z(n38154) );
  XOR U39169 ( .A(n38155), .B(n38154), .Z(n38146) );
  NANDN U39170 ( .A(n38125), .B(n38124), .Z(n38129) );
  NAND U39171 ( .A(n38127), .B(n38126), .Z(n38128) );
  NAND U39172 ( .A(n38129), .B(n38128), .Z(n38147) );
  XOR U39173 ( .A(n38143), .B(n38142), .Z(n38267) );
  XOR U39174 ( .A(n38268), .B(n38267), .Z(n38269) );
  XNOR U39175 ( .A(n38270), .B(n38269), .Z(n38263) );
  NANDN U39176 ( .A(n38134), .B(n38133), .Z(n38138) );
  NAND U39177 ( .A(n38136), .B(n38135), .Z(n38137) );
  NAND U39178 ( .A(n38138), .B(n38137), .Z(n38261) );
  IV U39179 ( .A(n38261), .Z(n38260) );
  XOR U39180 ( .A(n38262), .B(n38260), .Z(n38139) );
  XNOR U39181 ( .A(n38263), .B(n38139), .Z(N823) );
  NANDN U39182 ( .A(n38141), .B(n38140), .Z(n38145) );
  NAND U39183 ( .A(n38143), .B(n38142), .Z(n38144) );
  AND U39184 ( .A(n38145), .B(n38144), .Z(n38408) );
  NANDN U39185 ( .A(n38147), .B(n38146), .Z(n38151) );
  NANDN U39186 ( .A(n38149), .B(n38148), .Z(n38150) );
  AND U39187 ( .A(n38151), .B(n38150), .Z(n38406) );
  NAND U39188 ( .A(n38153), .B(n38152), .Z(n38157) );
  NAND U39189 ( .A(n38155), .B(n38154), .Z(n38156) );
  NAND U39190 ( .A(n38157), .B(n38156), .Z(n38390) );
  NAND U39191 ( .A(n38159), .B(n38158), .Z(n38163) );
  NAND U39192 ( .A(n38161), .B(n38160), .Z(n38162) );
  NAND U39193 ( .A(n38163), .B(n38162), .Z(n38383) );
  NAND U39194 ( .A(n38165), .B(n38164), .Z(n38169) );
  NAND U39195 ( .A(n38167), .B(n38166), .Z(n38168) );
  NAND U39196 ( .A(n38169), .B(n38168), .Z(n38382) );
  NAND U39197 ( .A(n38171), .B(n38170), .Z(n38175) );
  NAND U39198 ( .A(n38173), .B(n38172), .Z(n38174) );
  NAND U39199 ( .A(n38175), .B(n38174), .Z(n38381) );
  XOR U39200 ( .A(n38382), .B(n38381), .Z(n38384) );
  XOR U39201 ( .A(n38383), .B(n38384), .Z(n38401) );
  NAND U39202 ( .A(n38177), .B(n38176), .Z(n38181) );
  NAND U39203 ( .A(n38179), .B(n38178), .Z(n38180) );
  NAND U39204 ( .A(n38181), .B(n38180), .Z(n38399) );
  NAND U39205 ( .A(n38183), .B(n38182), .Z(n38187) );
  NAND U39206 ( .A(n38185), .B(n38184), .Z(n38186) );
  NAND U39207 ( .A(n38187), .B(n38186), .Z(n38328) );
  AND U39208 ( .A(n38189), .B(n38188), .Z(n38193) );
  NAND U39209 ( .A(n38191), .B(n38190), .Z(n38192) );
  NANDN U39210 ( .A(n38193), .B(n38192), .Z(n38327) );
  XOR U39211 ( .A(n38328), .B(n38327), .Z(n38330) );
  AND U39212 ( .A(y[8080]), .B(x[487]), .Z(n38195) );
  NAND U39213 ( .A(y[8078]), .B(x[489]), .Z(n38194) );
  XNOR U39214 ( .A(n38195), .B(n38194), .Z(n38295) );
  AND U39215 ( .A(x[490]), .B(y[8077]), .Z(n38334) );
  XOR U39216 ( .A(n38333), .B(n38334), .Z(n38336) );
  AND U39217 ( .A(x[486]), .B(y[8081]), .Z(n38286) );
  AND U39218 ( .A(x[495]), .B(y[8072]), .Z(n38287) );
  XOR U39219 ( .A(n38286), .B(n38287), .Z(n38288) );
  AND U39220 ( .A(x[491]), .B(y[8076]), .Z(n38289) );
  XOR U39221 ( .A(n38288), .B(n38289), .Z(n38335) );
  XOR U39222 ( .A(n38336), .B(n38335), .Z(n38329) );
  XOR U39223 ( .A(n38330), .B(n38329), .Z(n38400) );
  XNOR U39224 ( .A(n38399), .B(n38400), .Z(n38402) );
  NAND U39225 ( .A(n38197), .B(n38196), .Z(n38201) );
  NAND U39226 ( .A(n38199), .B(n38198), .Z(n38200) );
  NAND U39227 ( .A(n38201), .B(n38200), .Z(n38322) );
  AND U39228 ( .A(x[498]), .B(y[8074]), .Z(n39082) );
  NAND U39229 ( .A(n39082), .B(n38202), .Z(n38206) );
  NAND U39230 ( .A(n38204), .B(n38203), .Z(n38205) );
  AND U39231 ( .A(n38206), .B(n38205), .Z(n38370) );
  NAND U39232 ( .A(n38208), .B(n38207), .Z(n38212) );
  NAND U39233 ( .A(n38210), .B(n38209), .Z(n38211) );
  NAND U39234 ( .A(n38212), .B(n38211), .Z(n38369) );
  NANDN U39235 ( .A(n38296), .B(n38294), .Z(n38216) );
  NAND U39236 ( .A(n38214), .B(n38213), .Z(n38215) );
  AND U39237 ( .A(n38216), .B(n38215), .Z(n38366) );
  AND U39238 ( .A(x[480]), .B(y[8087]), .Z(n38305) );
  AND U39239 ( .A(x[503]), .B(y[8064]), .Z(n38306) );
  XOR U39240 ( .A(n38305), .B(n38306), .Z(n38308) );
  AND U39241 ( .A(x[502]), .B(y[8065]), .Z(n38285) );
  XOR U39242 ( .A(o[407]), .B(n38285), .Z(n38307) );
  XOR U39243 ( .A(n38308), .B(n38307), .Z(n38364) );
  NAND U39244 ( .A(y[8067]), .B(x[500]), .Z(n38217) );
  XNOR U39245 ( .A(n38218), .B(n38217), .Z(n38281) );
  AND U39246 ( .A(x[499]), .B(y[8068]), .Z(n38282) );
  XOR U39247 ( .A(n38281), .B(n38282), .Z(n38363) );
  XOR U39248 ( .A(n38364), .B(n38363), .Z(n38365) );
  XOR U39249 ( .A(n38372), .B(n38371), .Z(n38321) );
  XOR U39250 ( .A(n38322), .B(n38321), .Z(n38324) );
  NAND U39251 ( .A(x[500]), .B(y[8073]), .Z(n39258) );
  AND U39252 ( .A(x[493]), .B(y[8066]), .Z(n38219) );
  NANDN U39253 ( .A(n39258), .B(n38219), .Z(n38223) );
  NAND U39254 ( .A(n38221), .B(n38220), .Z(n38222) );
  NAND U39255 ( .A(n38223), .B(n38222), .Z(n38316) );
  NAND U39256 ( .A(n38225), .B(n38224), .Z(n38229) );
  NAND U39257 ( .A(n38227), .B(n38226), .Z(n38228) );
  AND U39258 ( .A(n38229), .B(n38228), .Z(n38378) );
  AND U39259 ( .A(x[493]), .B(y[8074]), .Z(n38351) );
  AND U39260 ( .A(x[482]), .B(y[8085]), .Z(n38352) );
  XOR U39261 ( .A(n38351), .B(n38352), .Z(n38353) );
  AND U39262 ( .A(x[501]), .B(y[8066]), .Z(n38354) );
  XOR U39263 ( .A(n38353), .B(n38354), .Z(n38376) );
  AND U39264 ( .A(x[492]), .B(y[8075]), .Z(n38299) );
  AND U39265 ( .A(x[481]), .B(y[8086]), .Z(n38300) );
  XOR U39266 ( .A(n38299), .B(n38300), .Z(n38302) );
  AND U39267 ( .A(o[406]), .B(n38230), .Z(n38301) );
  XOR U39268 ( .A(n38302), .B(n38301), .Z(n38375) );
  XOR U39269 ( .A(n38376), .B(n38375), .Z(n38377) );
  XOR U39270 ( .A(n38316), .B(n38315), .Z(n38318) );
  AND U39271 ( .A(x[495]), .B(y[8080]), .Z(n39383) );
  NAND U39272 ( .A(n39383), .B(n38231), .Z(n38235) );
  NANDN U39273 ( .A(n38233), .B(n38232), .Z(n38234) );
  AND U39274 ( .A(n38235), .B(n38234), .Z(n38360) );
  AND U39275 ( .A(x[494]), .B(y[8073]), .Z(n38345) );
  AND U39276 ( .A(x[483]), .B(y[8084]), .Z(n38346) );
  XOR U39277 ( .A(n38345), .B(n38346), .Z(n38347) );
  AND U39278 ( .A(x[484]), .B(y[8083]), .Z(n38348) );
  XOR U39279 ( .A(n38347), .B(n38348), .Z(n38358) );
  AND U39280 ( .A(x[485]), .B(y[8082]), .Z(n38339) );
  AND U39281 ( .A(x[498]), .B(y[8069]), .Z(n38340) );
  XOR U39282 ( .A(n38339), .B(n38340), .Z(n38341) );
  AND U39283 ( .A(x[497]), .B(y[8070]), .Z(n38342) );
  XOR U39284 ( .A(n38341), .B(n38342), .Z(n38357) );
  XOR U39285 ( .A(n38358), .B(n38357), .Z(n38359) );
  XOR U39286 ( .A(n38318), .B(n38317), .Z(n38323) );
  XOR U39287 ( .A(n38324), .B(n38323), .Z(n38387) );
  XOR U39288 ( .A(n38388), .B(n38387), .Z(n38389) );
  XNOR U39289 ( .A(n38390), .B(n38389), .Z(n38276) );
  NAND U39290 ( .A(n38237), .B(n38236), .Z(n38241) );
  NAND U39291 ( .A(n38239), .B(n38238), .Z(n38240) );
  NAND U39292 ( .A(n38241), .B(n38240), .Z(n38396) );
  NAND U39293 ( .A(n38243), .B(n38242), .Z(n38247) );
  NAND U39294 ( .A(n38245), .B(n38244), .Z(n38246) );
  NAND U39295 ( .A(n38247), .B(n38246), .Z(n38394) );
  NAND U39296 ( .A(n38249), .B(n38248), .Z(n38253) );
  NAND U39297 ( .A(n38251), .B(n38250), .Z(n38252) );
  NAND U39298 ( .A(n38253), .B(n38252), .Z(n38393) );
  XOR U39299 ( .A(n38394), .B(n38393), .Z(n38395) );
  XNOR U39300 ( .A(n38396), .B(n38395), .Z(n38275) );
  NAND U39301 ( .A(n38255), .B(n38254), .Z(n38259) );
  NAND U39302 ( .A(n38257), .B(n38256), .Z(n38258) );
  NAND U39303 ( .A(n38259), .B(n38258), .Z(n38274) );
  XOR U39304 ( .A(n38275), .B(n38274), .Z(n38277) );
  XOR U39305 ( .A(n38276), .B(n38277), .Z(n38405) );
  XOR U39306 ( .A(n38406), .B(n38405), .Z(n38407) );
  XNOR U39307 ( .A(n38408), .B(n38407), .Z(n38414) );
  OR U39308 ( .A(n38262), .B(n38260), .Z(n38266) );
  ANDN U39309 ( .B(n38262), .A(n38261), .Z(n38264) );
  OR U39310 ( .A(n38264), .B(n38263), .Z(n38265) );
  AND U39311 ( .A(n38266), .B(n38265), .Z(n38412) );
  NAND U39312 ( .A(n38268), .B(n38267), .Z(n38272) );
  NAND U39313 ( .A(n38270), .B(n38269), .Z(n38271) );
  AND U39314 ( .A(n38272), .B(n38271), .Z(n38413) );
  IV U39315 ( .A(n38413), .Z(n38411) );
  XOR U39316 ( .A(n38412), .B(n38411), .Z(n38273) );
  XNOR U39317 ( .A(n38414), .B(n38273), .Z(N824) );
  NAND U39318 ( .A(n38275), .B(n38274), .Z(n38279) );
  NAND U39319 ( .A(n38277), .B(n38276), .Z(n38278) );
  AND U39320 ( .A(n38279), .B(n38278), .Z(n38552) );
  AND U39321 ( .A(x[500]), .B(y[8071]), .Z(n38280) );
  NAND U39322 ( .A(n38280), .B(n38443), .Z(n38284) );
  NAND U39323 ( .A(n38282), .B(n38281), .Z(n38283) );
  NAND U39324 ( .A(n38284), .B(n38283), .Z(n38463) );
  AND U39325 ( .A(x[502]), .B(y[8066]), .Z(n38482) );
  XOR U39326 ( .A(n38483), .B(n38482), .Z(n38484) );
  AND U39327 ( .A(x[482]), .B(y[8086]), .Z(n38485) );
  XOR U39328 ( .A(n38484), .B(n38485), .Z(n38461) );
  AND U39329 ( .A(x[481]), .B(y[8087]), .Z(n38490) );
  XOR U39330 ( .A(n38491), .B(n38490), .Z(n38489) );
  AND U39331 ( .A(o[407]), .B(n38285), .Z(n38488) );
  XOR U39332 ( .A(n38489), .B(n38488), .Z(n38460) );
  XOR U39333 ( .A(n38461), .B(n38460), .Z(n38462) );
  XOR U39334 ( .A(n38463), .B(n38462), .Z(n38520) );
  NAND U39335 ( .A(n38287), .B(n38286), .Z(n38291) );
  NAND U39336 ( .A(n38289), .B(n38288), .Z(n38290) );
  NAND U39337 ( .A(n38291), .B(n38290), .Z(n38457) );
  AND U39338 ( .A(y[8072]), .B(x[496]), .Z(n38293) );
  NAND U39339 ( .A(y[8067]), .B(x[501]), .Z(n38292) );
  XNOR U39340 ( .A(n38293), .B(n38292), .Z(n38444) );
  AND U39341 ( .A(x[485]), .B(y[8083]), .Z(n38445) );
  XOR U39342 ( .A(n38444), .B(n38445), .Z(n38455) );
  AND U39343 ( .A(x[486]), .B(y[8082]), .Z(n38833) );
  AND U39344 ( .A(x[500]), .B(y[8068]), .Z(n38658) );
  XOR U39345 ( .A(n38833), .B(n38658), .Z(n38450) );
  AND U39346 ( .A(x[499]), .B(y[8069]), .Z(n38451) );
  XOR U39347 ( .A(n38450), .B(n38451), .Z(n38454) );
  XOR U39348 ( .A(n38455), .B(n38454), .Z(n38456) );
  XOR U39349 ( .A(n38457), .B(n38456), .Z(n38434) );
  NANDN U39350 ( .A(n38584), .B(n38294), .Z(n38298) );
  NANDN U39351 ( .A(n38296), .B(n38295), .Z(n38297) );
  NAND U39352 ( .A(n38298), .B(n38297), .Z(n38432) );
  NAND U39353 ( .A(n38300), .B(n38299), .Z(n38304) );
  NAND U39354 ( .A(n38302), .B(n38301), .Z(n38303) );
  NAND U39355 ( .A(n38304), .B(n38303), .Z(n38431) );
  XOR U39356 ( .A(n38432), .B(n38431), .Z(n38433) );
  XOR U39357 ( .A(n38434), .B(n38433), .Z(n38519) );
  XOR U39358 ( .A(n38520), .B(n38519), .Z(n38522) );
  NAND U39359 ( .A(n38306), .B(n38305), .Z(n38310) );
  NAND U39360 ( .A(n38308), .B(n38307), .Z(n38309) );
  AND U39361 ( .A(n38310), .B(n38309), .Z(n38514) );
  AND U39362 ( .A(x[483]), .B(y[8085]), .Z(n38503) );
  XOR U39363 ( .A(n38504), .B(n38503), .Z(n38502) );
  AND U39364 ( .A(x[484]), .B(y[8084]), .Z(n38501) );
  XOR U39365 ( .A(n38502), .B(n38501), .Z(n38513) );
  AND U39366 ( .A(y[8079]), .B(x[489]), .Z(n38312) );
  NAND U39367 ( .A(y[8078]), .B(x[490]), .Z(n38311) );
  XNOR U39368 ( .A(n38312), .B(n38311), .Z(n38474) );
  AND U39369 ( .A(y[8074]), .B(x[494]), .Z(n38314) );
  NAND U39370 ( .A(y[8080]), .B(x[488]), .Z(n38313) );
  XNOR U39371 ( .A(n38314), .B(n38313), .Z(n38478) );
  NAND U39372 ( .A(x[491]), .B(y[8077]), .Z(n38479) );
  XOR U39373 ( .A(n38474), .B(n38473), .Z(n38515) );
  XOR U39374 ( .A(n38516), .B(n38515), .Z(n38521) );
  XOR U39375 ( .A(n38522), .B(n38521), .Z(n38532) );
  NAND U39376 ( .A(n38316), .B(n38315), .Z(n38320) );
  NAND U39377 ( .A(n38318), .B(n38317), .Z(n38319) );
  AND U39378 ( .A(n38320), .B(n38319), .Z(n38531) );
  NAND U39379 ( .A(n38322), .B(n38321), .Z(n38326) );
  NAND U39380 ( .A(n38324), .B(n38323), .Z(n38325) );
  NAND U39381 ( .A(n38326), .B(n38325), .Z(n38534) );
  NAND U39382 ( .A(n38328), .B(n38327), .Z(n38332) );
  NAND U39383 ( .A(n38330), .B(n38329), .Z(n38331) );
  NAND U39384 ( .A(n38332), .B(n38331), .Z(n38528) );
  NAND U39385 ( .A(n38334), .B(n38333), .Z(n38338) );
  NAND U39386 ( .A(n38336), .B(n38335), .Z(n38337) );
  NAND U39387 ( .A(n38338), .B(n38337), .Z(n38526) );
  NAND U39388 ( .A(n38340), .B(n38339), .Z(n38344) );
  NAND U39389 ( .A(n38342), .B(n38341), .Z(n38343) );
  NAND U39390 ( .A(n38344), .B(n38343), .Z(n38440) );
  AND U39391 ( .A(x[480]), .B(y[8088]), .Z(n38508) );
  AND U39392 ( .A(x[504]), .B(y[8064]), .Z(n38507) );
  XOR U39393 ( .A(n38508), .B(n38507), .Z(n38510) );
  AND U39394 ( .A(x[503]), .B(y[8065]), .Z(n38500) );
  XOR U39395 ( .A(n38500), .B(o[408]), .Z(n38509) );
  XOR U39396 ( .A(n38510), .B(n38509), .Z(n38438) );
  AND U39397 ( .A(x[487]), .B(y[8081]), .Z(n38494) );
  AND U39398 ( .A(x[498]), .B(y[8070]), .Z(n38495) );
  XOR U39399 ( .A(n38494), .B(n38495), .Z(n38496) );
  AND U39400 ( .A(x[497]), .B(y[8071]), .Z(n38497) );
  XOR U39401 ( .A(n38496), .B(n38497), .Z(n38437) );
  XOR U39402 ( .A(n38438), .B(n38437), .Z(n38439) );
  XOR U39403 ( .A(n38440), .B(n38439), .Z(n38428) );
  NAND U39404 ( .A(n38346), .B(n38345), .Z(n38350) );
  NAND U39405 ( .A(n38348), .B(n38347), .Z(n38349) );
  NAND U39406 ( .A(n38350), .B(n38349), .Z(n38426) );
  NAND U39407 ( .A(n38352), .B(n38351), .Z(n38356) );
  NAND U39408 ( .A(n38354), .B(n38353), .Z(n38355) );
  NAND U39409 ( .A(n38356), .B(n38355), .Z(n38425) );
  XOR U39410 ( .A(n38426), .B(n38425), .Z(n38427) );
  XOR U39411 ( .A(n38428), .B(n38427), .Z(n38525) );
  XOR U39412 ( .A(n38526), .B(n38525), .Z(n38527) );
  XNOR U39413 ( .A(n38528), .B(n38527), .Z(n38421) );
  NAND U39414 ( .A(n38358), .B(n38357), .Z(n38362) );
  NANDN U39415 ( .A(n38360), .B(n38359), .Z(n38361) );
  AND U39416 ( .A(n38362), .B(n38361), .Z(n38466) );
  NAND U39417 ( .A(n38364), .B(n38363), .Z(n38368) );
  NANDN U39418 ( .A(n38366), .B(n38365), .Z(n38367) );
  NAND U39419 ( .A(n38368), .B(n38367), .Z(n38467) );
  NANDN U39420 ( .A(n38370), .B(n38369), .Z(n38374) );
  NAND U39421 ( .A(n38372), .B(n38371), .Z(n38373) );
  NAND U39422 ( .A(n38374), .B(n38373), .Z(n38469) );
  NAND U39423 ( .A(n38376), .B(n38375), .Z(n38380) );
  NANDN U39424 ( .A(n38378), .B(n38377), .Z(n38379) );
  NAND U39425 ( .A(n38380), .B(n38379), .Z(n38420) );
  XOR U39426 ( .A(n38421), .B(n38422), .Z(n38538) );
  NAND U39427 ( .A(n38382), .B(n38381), .Z(n38386) );
  NAND U39428 ( .A(n38384), .B(n38383), .Z(n38385) );
  AND U39429 ( .A(n38386), .B(n38385), .Z(n38537) );
  XOR U39430 ( .A(n38538), .B(n38537), .Z(n38539) );
  XNOR U39431 ( .A(n38540), .B(n38539), .Z(n38550) );
  NAND U39432 ( .A(n38388), .B(n38387), .Z(n38392) );
  NAND U39433 ( .A(n38390), .B(n38389), .Z(n38391) );
  NAND U39434 ( .A(n38392), .B(n38391), .Z(n38545) );
  NAND U39435 ( .A(n38394), .B(n38393), .Z(n38398) );
  NAND U39436 ( .A(n38396), .B(n38395), .Z(n38397) );
  NAND U39437 ( .A(n38398), .B(n38397), .Z(n38544) );
  NAND U39438 ( .A(n38400), .B(n38399), .Z(n38404) );
  NANDN U39439 ( .A(n38402), .B(n38401), .Z(n38403) );
  NAND U39440 ( .A(n38404), .B(n38403), .Z(n38543) );
  XOR U39441 ( .A(n38544), .B(n38543), .Z(n38546) );
  XOR U39442 ( .A(n38545), .B(n38546), .Z(n38549) );
  XOR U39443 ( .A(n38550), .B(n38549), .Z(n38551) );
  XOR U39444 ( .A(n38552), .B(n38551), .Z(n38557) );
  NAND U39445 ( .A(n38406), .B(n38405), .Z(n38410) );
  NAND U39446 ( .A(n38408), .B(n38407), .Z(n38409) );
  NAND U39447 ( .A(n38410), .B(n38409), .Z(n38555) );
  NANDN U39448 ( .A(n38411), .B(n38412), .Z(n38417) );
  NOR U39449 ( .A(n38413), .B(n38412), .Z(n38415) );
  OR U39450 ( .A(n38415), .B(n38414), .Z(n38416) );
  AND U39451 ( .A(n38417), .B(n38416), .Z(n38556) );
  XOR U39452 ( .A(n38555), .B(n38556), .Z(n38418) );
  XNOR U39453 ( .A(n38557), .B(n38418), .Z(N825) );
  NANDN U39454 ( .A(n38420), .B(n38419), .Z(n38424) );
  NAND U39455 ( .A(n38422), .B(n38421), .Z(n38423) );
  AND U39456 ( .A(n38424), .B(n38423), .Z(n38568) );
  NAND U39457 ( .A(n38426), .B(n38425), .Z(n38430) );
  NAND U39458 ( .A(n38428), .B(n38427), .Z(n38429) );
  NAND U39459 ( .A(n38430), .B(n38429), .Z(n38572) );
  NAND U39460 ( .A(n38432), .B(n38431), .Z(n38436) );
  NAND U39461 ( .A(n38434), .B(n38433), .Z(n38435) );
  NAND U39462 ( .A(n38436), .B(n38435), .Z(n38571) );
  XOR U39463 ( .A(n38572), .B(n38571), .Z(n38574) );
  NAND U39464 ( .A(n38438), .B(n38437), .Z(n38442) );
  NAND U39465 ( .A(n38440), .B(n38439), .Z(n38441) );
  AND U39466 ( .A(n38442), .B(n38441), .Z(n38604) );
  AND U39467 ( .A(x[501]), .B(y[8072]), .Z(n39487) );
  NAND U39468 ( .A(n39487), .B(n38443), .Z(n38447) );
  NAND U39469 ( .A(n38445), .B(n38444), .Z(n38446) );
  NAND U39470 ( .A(n38447), .B(n38446), .Z(n38678) );
  NAND U39471 ( .A(x[502]), .B(y[8067]), .Z(n38647) );
  NAND U39472 ( .A(x[485]), .B(y[8084]), .Z(n38646) );
  NAND U39473 ( .A(x[497]), .B(y[8072]), .Z(n38645) );
  XOR U39474 ( .A(n38646), .B(n38645), .Z(n38648) );
  XNOR U39475 ( .A(n38647), .B(n38648), .Z(n38677) );
  AND U39476 ( .A(y[8069]), .B(x[500]), .Z(n38449) );
  NAND U39477 ( .A(y[8068]), .B(x[501]), .Z(n38448) );
  XNOR U39478 ( .A(n38449), .B(n38448), .Z(n38660) );
  AND U39479 ( .A(x[499]), .B(y[8070]), .Z(n38659) );
  XOR U39480 ( .A(n38660), .B(n38659), .Z(n38676) );
  XNOR U39481 ( .A(n38677), .B(n38676), .Z(n38679) );
  XOR U39482 ( .A(n38678), .B(n38679), .Z(n38602) );
  NAND U39483 ( .A(n38658), .B(n38833), .Z(n38453) );
  NAND U39484 ( .A(n38451), .B(n38450), .Z(n38452) );
  NAND U39485 ( .A(n38453), .B(n38452), .Z(n38684) );
  NAND U39486 ( .A(x[495]), .B(y[8074]), .Z(n38666) );
  NAND U39487 ( .A(x[498]), .B(y[8071]), .Z(n38665) );
  NAND U39488 ( .A(x[486]), .B(y[8083]), .Z(n38664) );
  XOR U39489 ( .A(n38665), .B(n38664), .Z(n38667) );
  XNOR U39490 ( .A(n38666), .B(n38667), .Z(n38683) );
  NAND U39491 ( .A(x[503]), .B(y[8066]), .Z(n38641) );
  NAND U39492 ( .A(x[484]), .B(y[8085]), .Z(n38640) );
  NAND U39493 ( .A(x[496]), .B(y[8073]), .Z(n38639) );
  XOR U39494 ( .A(n38640), .B(n38639), .Z(n38642) );
  XNOR U39495 ( .A(n38641), .B(n38642), .Z(n38682) );
  XNOR U39496 ( .A(n38683), .B(n38682), .Z(n38685) );
  XOR U39497 ( .A(n38684), .B(n38685), .Z(n38601) );
  XOR U39498 ( .A(n38602), .B(n38601), .Z(n38603) );
  XNOR U39499 ( .A(n38604), .B(n38603), .Z(n38616) );
  NAND U39500 ( .A(n38455), .B(n38454), .Z(n38459) );
  NAND U39501 ( .A(n38457), .B(n38456), .Z(n38458) );
  NAND U39502 ( .A(n38459), .B(n38458), .Z(n38614) );
  NAND U39503 ( .A(n38461), .B(n38460), .Z(n38465) );
  NAND U39504 ( .A(n38463), .B(n38462), .Z(n38464) );
  NAND U39505 ( .A(n38465), .B(n38464), .Z(n38613) );
  XOR U39506 ( .A(n38614), .B(n38613), .Z(n38615) );
  XOR U39507 ( .A(n38616), .B(n38615), .Z(n38573) );
  XOR U39508 ( .A(n38574), .B(n38573), .Z(n38566) );
  NANDN U39509 ( .A(n38467), .B(n38466), .Z(n38471) );
  NANDN U39510 ( .A(n38469), .B(n38468), .Z(n38470) );
  NAND U39511 ( .A(n38471), .B(n38470), .Z(n38565) );
  NANDN U39512 ( .A(n38583), .B(n38472), .Z(n38476) );
  NAND U39513 ( .A(n38474), .B(n38473), .Z(n38475) );
  NAND U39514 ( .A(n38476), .B(n38475), .Z(n38608) );
  NAND U39515 ( .A(x[494]), .B(y[8080]), .Z(n39501) );
  NANDN U39516 ( .A(n39501), .B(n38477), .Z(n38481) );
  NANDN U39517 ( .A(n38479), .B(n38478), .Z(n38480) );
  NAND U39518 ( .A(n38481), .B(n38480), .Z(n38635) );
  NAND U39519 ( .A(x[491]), .B(y[8078]), .Z(n38654) );
  NAND U39520 ( .A(x[492]), .B(y[8077]), .Z(n38653) );
  NAND U39521 ( .A(x[487]), .B(y[8082]), .Z(n38652) );
  XOR U39522 ( .A(n38653), .B(n38652), .Z(n38655) );
  XOR U39523 ( .A(n38654), .B(n38655), .Z(n38634) );
  AND U39524 ( .A(x[504]), .B(y[8065]), .Z(n38651) );
  XOR U39525 ( .A(o[409]), .B(n38651), .Z(n38622) );
  AND U39526 ( .A(x[481]), .B(y[8088]), .Z(n38621) );
  XOR U39527 ( .A(n38622), .B(n38621), .Z(n38624) );
  AND U39528 ( .A(x[493]), .B(y[8076]), .Z(n38623) );
  XOR U39529 ( .A(n38624), .B(n38623), .Z(n38633) );
  XOR U39530 ( .A(n38635), .B(n38636), .Z(n38607) );
  XOR U39531 ( .A(n38608), .B(n38607), .Z(n38610) );
  AND U39532 ( .A(n38483), .B(n38482), .Z(n38487) );
  NAND U39533 ( .A(n38485), .B(n38484), .Z(n38486) );
  NANDN U39534 ( .A(n38487), .B(n38486), .Z(n38596) );
  AND U39535 ( .A(n38489), .B(n38488), .Z(n38493) );
  NAND U39536 ( .A(n38491), .B(n38490), .Z(n38492) );
  NANDN U39537 ( .A(n38493), .B(n38492), .Z(n38595) );
  XOR U39538 ( .A(n38596), .B(n38595), .Z(n38597) );
  NAND U39539 ( .A(n38495), .B(n38494), .Z(n38499) );
  NAND U39540 ( .A(n38497), .B(n38496), .Z(n38498) );
  NAND U39541 ( .A(n38499), .B(n38498), .Z(n38591) );
  NAND U39542 ( .A(x[488]), .B(y[8081]), .Z(n38585) );
  XOR U39543 ( .A(n38584), .B(n38583), .Z(n38586) );
  XNOR U39544 ( .A(n38585), .B(n38586), .Z(n38590) );
  NAND U39545 ( .A(n38500), .B(o[408]), .Z(n38579) );
  NAND U39546 ( .A(x[505]), .B(y[8064]), .Z(n38578) );
  NAND U39547 ( .A(x[480]), .B(y[8089]), .Z(n38577) );
  XOR U39548 ( .A(n38578), .B(n38577), .Z(n38580) );
  XNOR U39549 ( .A(n38579), .B(n38580), .Z(n38589) );
  XNOR U39550 ( .A(n38590), .B(n38589), .Z(n38592) );
  XOR U39551 ( .A(n38591), .B(n38592), .Z(n38598) );
  XNOR U39552 ( .A(n38597), .B(n38598), .Z(n38609) );
  XOR U39553 ( .A(n38610), .B(n38609), .Z(n38691) );
  AND U39554 ( .A(n38502), .B(n38501), .Z(n38506) );
  NAND U39555 ( .A(n38504), .B(n38503), .Z(n38505) );
  NANDN U39556 ( .A(n38506), .B(n38505), .Z(n38673) );
  NAND U39557 ( .A(n38508), .B(n38507), .Z(n38512) );
  NAND U39558 ( .A(n38510), .B(n38509), .Z(n38511) );
  NAND U39559 ( .A(n38512), .B(n38511), .Z(n38671) );
  AND U39560 ( .A(x[494]), .B(y[8075]), .Z(n38628) );
  AND U39561 ( .A(x[482]), .B(y[8087]), .Z(n38627) );
  XOR U39562 ( .A(n38628), .B(n38627), .Z(n38630) );
  AND U39563 ( .A(x[483]), .B(y[8086]), .Z(n38629) );
  XOR U39564 ( .A(n38630), .B(n38629), .Z(n38670) );
  XOR U39565 ( .A(n38671), .B(n38670), .Z(n38672) );
  XNOR U39566 ( .A(n38673), .B(n38672), .Z(n38688) );
  NANDN U39567 ( .A(n38514), .B(n38513), .Z(n38518) );
  NAND U39568 ( .A(n38516), .B(n38515), .Z(n38517) );
  AND U39569 ( .A(n38518), .B(n38517), .Z(n38689) );
  XOR U39570 ( .A(n38688), .B(n38689), .Z(n38690) );
  NAND U39571 ( .A(n38520), .B(n38519), .Z(n38524) );
  NAND U39572 ( .A(n38522), .B(n38521), .Z(n38523) );
  AND U39573 ( .A(n38524), .B(n38523), .Z(n38695) );
  XOR U39574 ( .A(n38694), .B(n38695), .Z(n38697) );
  NAND U39575 ( .A(n38526), .B(n38525), .Z(n38530) );
  NAND U39576 ( .A(n38528), .B(n38527), .Z(n38529) );
  AND U39577 ( .A(n38530), .B(n38529), .Z(n38696) );
  XOR U39578 ( .A(n38697), .B(n38696), .Z(n38560) );
  NANDN U39579 ( .A(n38532), .B(n38531), .Z(n38536) );
  NANDN U39580 ( .A(n38534), .B(n38533), .Z(n38535) );
  AND U39581 ( .A(n38536), .B(n38535), .Z(n38559) );
  XOR U39582 ( .A(n38561), .B(n38562), .Z(n38704) );
  NAND U39583 ( .A(n38538), .B(n38537), .Z(n38542) );
  NAND U39584 ( .A(n38540), .B(n38539), .Z(n38541) );
  NAND U39585 ( .A(n38542), .B(n38541), .Z(n38703) );
  NAND U39586 ( .A(n38544), .B(n38543), .Z(n38548) );
  NAND U39587 ( .A(n38546), .B(n38545), .Z(n38547) );
  AND U39588 ( .A(n38548), .B(n38547), .Z(n38705) );
  XOR U39589 ( .A(n38706), .B(n38705), .Z(n38702) );
  NAND U39590 ( .A(n38550), .B(n38549), .Z(n38554) );
  NAND U39591 ( .A(n38552), .B(n38551), .Z(n38553) );
  NAND U39592 ( .A(n38554), .B(n38553), .Z(n38701) );
  XOR U39593 ( .A(n38701), .B(n38700), .Z(n38558) );
  XNOR U39594 ( .A(n38702), .B(n38558), .Z(N826) );
  NANDN U39595 ( .A(n38560), .B(n38559), .Z(n38564) );
  NAND U39596 ( .A(n38562), .B(n38561), .Z(n38563) );
  AND U39597 ( .A(n38564), .B(n38563), .Z(n38711) );
  NANDN U39598 ( .A(n38566), .B(n38565), .Z(n38570) );
  NANDN U39599 ( .A(n38568), .B(n38567), .Z(n38569) );
  AND U39600 ( .A(n38570), .B(n38569), .Z(n38710) );
  NAND U39601 ( .A(n38572), .B(n38571), .Z(n38576) );
  NAND U39602 ( .A(n38574), .B(n38573), .Z(n38575) );
  NAND U39603 ( .A(n38576), .B(n38575), .Z(n38868) );
  AND U39604 ( .A(x[482]), .B(y[8088]), .Z(n38741) );
  XOR U39605 ( .A(n38742), .B(n38741), .Z(n38744) );
  AND U39606 ( .A(x[504]), .B(y[8066]), .Z(n38743) );
  XOR U39607 ( .A(n38744), .B(n38743), .Z(n38784) );
  NAND U39608 ( .A(n38578), .B(n38577), .Z(n38582) );
  NAND U39609 ( .A(n38580), .B(n38579), .Z(n38581) );
  AND U39610 ( .A(n38582), .B(n38581), .Z(n38783) );
  XOR U39611 ( .A(n38784), .B(n38783), .Z(n38786) );
  NAND U39612 ( .A(n38584), .B(n38583), .Z(n38588) );
  NAND U39613 ( .A(n38586), .B(n38585), .Z(n38587) );
  AND U39614 ( .A(n38588), .B(n38587), .Z(n38785) );
  XNOR U39615 ( .A(n38786), .B(n38785), .Z(n38848) );
  NAND U39616 ( .A(n38590), .B(n38589), .Z(n38594) );
  NANDN U39617 ( .A(n38592), .B(n38591), .Z(n38593) );
  AND U39618 ( .A(n38594), .B(n38593), .Z(n38847) );
  XOR U39619 ( .A(n38848), .B(n38847), .Z(n38850) );
  NAND U39620 ( .A(n38596), .B(n38595), .Z(n38600) );
  NANDN U39621 ( .A(n38598), .B(n38597), .Z(n38599) );
  AND U39622 ( .A(n38600), .B(n38599), .Z(n38849) );
  XOR U39623 ( .A(n38850), .B(n38849), .Z(n38862) );
  NAND U39624 ( .A(n38602), .B(n38601), .Z(n38606) );
  NAND U39625 ( .A(n38604), .B(n38603), .Z(n38605) );
  NAND U39626 ( .A(n38606), .B(n38605), .Z(n38860) );
  NAND U39627 ( .A(n38608), .B(n38607), .Z(n38612) );
  NAND U39628 ( .A(n38610), .B(n38609), .Z(n38611) );
  AND U39629 ( .A(n38612), .B(n38611), .Z(n38859) );
  XOR U39630 ( .A(n38860), .B(n38859), .Z(n38861) );
  XNOR U39631 ( .A(n38862), .B(n38861), .Z(n38866) );
  NAND U39632 ( .A(n38614), .B(n38613), .Z(n38618) );
  NAND U39633 ( .A(n38616), .B(n38615), .Z(n38617) );
  NAND U39634 ( .A(n38618), .B(n38617), .Z(n38812) );
  AND U39635 ( .A(y[8084]), .B(x[486]), .Z(n38620) );
  NAND U39636 ( .A(y[8082]), .B(x[488]), .Z(n38619) );
  XNOR U39637 ( .A(n38620), .B(n38619), .Z(n38835) );
  AND U39638 ( .A(x[489]), .B(y[8081]), .Z(n38834) );
  XOR U39639 ( .A(n38835), .B(n38834), .Z(n38815) );
  AND U39640 ( .A(x[487]), .B(y[8083]), .Z(n38816) );
  XOR U39641 ( .A(n38815), .B(n38816), .Z(n38818) );
  AND U39642 ( .A(x[492]), .B(y[8078]), .Z(n38935) );
  AND U39643 ( .A(x[485]), .B(y[8085]), .Z(n38798) );
  XOR U39644 ( .A(n38935), .B(n38798), .Z(n38800) );
  AND U39645 ( .A(x[490]), .B(y[8080]), .Z(n38799) );
  XOR U39646 ( .A(n38800), .B(n38799), .Z(n38817) );
  XOR U39647 ( .A(n38818), .B(n38817), .Z(n38768) );
  NAND U39648 ( .A(n38622), .B(n38621), .Z(n38626) );
  NAND U39649 ( .A(n38624), .B(n38623), .Z(n38625) );
  NAND U39650 ( .A(n38626), .B(n38625), .Z(n38766) );
  NAND U39651 ( .A(n38628), .B(n38627), .Z(n38632) );
  NAND U39652 ( .A(n38630), .B(n38629), .Z(n38631) );
  NAND U39653 ( .A(n38632), .B(n38631), .Z(n38765) );
  XOR U39654 ( .A(n38766), .B(n38765), .Z(n38767) );
  XNOR U39655 ( .A(n38768), .B(n38767), .Z(n38772) );
  NANDN U39656 ( .A(n38634), .B(n38633), .Z(n38638) );
  NAND U39657 ( .A(n38636), .B(n38635), .Z(n38637) );
  AND U39658 ( .A(n38638), .B(n38637), .Z(n38771) );
  XOR U39659 ( .A(n38772), .B(n38771), .Z(n38774) );
  NAND U39660 ( .A(n38640), .B(n38639), .Z(n38644) );
  NAND U39661 ( .A(n38642), .B(n38641), .Z(n38643) );
  AND U39662 ( .A(n38644), .B(n38643), .Z(n38729) );
  NAND U39663 ( .A(n38646), .B(n38645), .Z(n38650) );
  NAND U39664 ( .A(n38648), .B(n38647), .Z(n38649) );
  AND U39665 ( .A(n38650), .B(n38649), .Z(n38730) );
  XOR U39666 ( .A(n38729), .B(n38730), .Z(n38732) );
  AND U39667 ( .A(n38651), .B(o[409]), .Z(n38827) );
  AND U39668 ( .A(x[494]), .B(y[8076]), .Z(n38828) );
  XOR U39669 ( .A(n38827), .B(n38828), .Z(n38829) );
  AND U39670 ( .A(x[481]), .B(y[8089]), .Z(n38830) );
  XOR U39671 ( .A(n38829), .B(n38830), .Z(n38790) );
  NAND U39672 ( .A(x[505]), .B(y[8065]), .Z(n38838) );
  XNOR U39673 ( .A(o[410]), .B(n38838), .Z(n38804) );
  AND U39674 ( .A(x[506]), .B(y[8064]), .Z(n38803) );
  XOR U39675 ( .A(n38804), .B(n38803), .Z(n38806) );
  AND U39676 ( .A(x[480]), .B(y[8090]), .Z(n38805) );
  XOR U39677 ( .A(n38806), .B(n38805), .Z(n38789) );
  XOR U39678 ( .A(n38790), .B(n38789), .Z(n38792) );
  NAND U39679 ( .A(n38653), .B(n38652), .Z(n38657) );
  NAND U39680 ( .A(n38655), .B(n38654), .Z(n38656) );
  AND U39681 ( .A(n38657), .B(n38656), .Z(n38791) );
  XOR U39682 ( .A(n38792), .B(n38791), .Z(n38731) );
  XOR U39683 ( .A(n38732), .B(n38731), .Z(n38780) );
  AND U39684 ( .A(x[501]), .B(y[8069]), .Z(n38663) );
  IV U39685 ( .A(n38663), .Z(n38821) );
  NANDN U39686 ( .A(n38821), .B(n38658), .Z(n38662) );
  NAND U39687 ( .A(n38660), .B(n38659), .Z(n38661) );
  NAND U39688 ( .A(n38662), .B(n38661), .Z(n38762) );
  XOR U39689 ( .A(n38822), .B(n38663), .Z(n38823) );
  AND U39690 ( .A(x[500]), .B(y[8070]), .Z(n38824) );
  XOR U39691 ( .A(n38823), .B(n38824), .Z(n38760) );
  AND U39692 ( .A(x[503]), .B(y[8067]), .Z(n38748) );
  XOR U39693 ( .A(n38747), .B(n38748), .Z(n38749) );
  AND U39694 ( .A(x[502]), .B(y[8068]), .Z(n38750) );
  XOR U39695 ( .A(n38749), .B(n38750), .Z(n38759) );
  XOR U39696 ( .A(n38760), .B(n38759), .Z(n38761) );
  XOR U39697 ( .A(n38762), .B(n38761), .Z(n38778) );
  AND U39698 ( .A(x[484]), .B(y[8086]), .Z(n38753) );
  XOR U39699 ( .A(n38754), .B(n38753), .Z(n38755) );
  XNOR U39700 ( .A(n38755), .B(n38756), .Z(n38736) );
  AND U39701 ( .A(x[499]), .B(y[8071]), .Z(n38839) );
  AND U39702 ( .A(x[483]), .B(y[8087]), .Z(n38840) );
  XOR U39703 ( .A(n38839), .B(n38840), .Z(n38841) );
  AND U39704 ( .A(x[491]), .B(y[8079]), .Z(n38842) );
  XOR U39705 ( .A(n38841), .B(n38842), .Z(n38735) );
  XOR U39706 ( .A(n38736), .B(n38735), .Z(n38738) );
  NAND U39707 ( .A(n38665), .B(n38664), .Z(n38669) );
  NAND U39708 ( .A(n38667), .B(n38666), .Z(n38668) );
  AND U39709 ( .A(n38669), .B(n38668), .Z(n38737) );
  XNOR U39710 ( .A(n38738), .B(n38737), .Z(n38777) );
  XNOR U39711 ( .A(n38774), .B(n38773), .Z(n38810) );
  NAND U39712 ( .A(n38671), .B(n38670), .Z(n38675) );
  NAND U39713 ( .A(n38673), .B(n38672), .Z(n38674) );
  NAND U39714 ( .A(n38675), .B(n38674), .Z(n38856) );
  NAND U39715 ( .A(n38677), .B(n38676), .Z(n38681) );
  NANDN U39716 ( .A(n38679), .B(n38678), .Z(n38680) );
  NAND U39717 ( .A(n38681), .B(n38680), .Z(n38854) );
  NAND U39718 ( .A(n38683), .B(n38682), .Z(n38687) );
  NANDN U39719 ( .A(n38685), .B(n38684), .Z(n38686) );
  NAND U39720 ( .A(n38687), .B(n38686), .Z(n38853) );
  XOR U39721 ( .A(n38854), .B(n38853), .Z(n38855) );
  XOR U39722 ( .A(n38856), .B(n38855), .Z(n38809) );
  XOR U39723 ( .A(n38810), .B(n38809), .Z(n38811) );
  XOR U39724 ( .A(n38812), .B(n38811), .Z(n38865) );
  XOR U39725 ( .A(n38866), .B(n38865), .Z(n38867) );
  XOR U39726 ( .A(n38868), .B(n38867), .Z(n38726) );
  NAND U39727 ( .A(n38689), .B(n38688), .Z(n38693) );
  NANDN U39728 ( .A(n38691), .B(n38690), .Z(n38692) );
  AND U39729 ( .A(n38693), .B(n38692), .Z(n38723) );
  NAND U39730 ( .A(n38695), .B(n38694), .Z(n38699) );
  NAND U39731 ( .A(n38697), .B(n38696), .Z(n38698) );
  AND U39732 ( .A(n38699), .B(n38698), .Z(n38724) );
  XOR U39733 ( .A(n38723), .B(n38724), .Z(n38725) );
  XOR U39734 ( .A(n38726), .B(n38725), .Z(n38712) );
  XNOR U39735 ( .A(n38713), .B(n38712), .Z(n38719) );
  NANDN U39736 ( .A(n38704), .B(n38703), .Z(n38708) );
  NAND U39737 ( .A(n38706), .B(n38705), .Z(n38707) );
  AND U39738 ( .A(n38708), .B(n38707), .Z(n38717) );
  IV U39739 ( .A(n38717), .Z(n38716) );
  XOR U39740 ( .A(n38718), .B(n38716), .Z(n38709) );
  XNOR U39741 ( .A(n38719), .B(n38709), .Z(N827) );
  NANDN U39742 ( .A(n38711), .B(n38710), .Z(n38715) );
  NAND U39743 ( .A(n38713), .B(n38712), .Z(n38714) );
  NAND U39744 ( .A(n38715), .B(n38714), .Z(n38879) );
  IV U39745 ( .A(n38879), .Z(n38878) );
  OR U39746 ( .A(n38718), .B(n38716), .Z(n38722) );
  ANDN U39747 ( .B(n38718), .A(n38717), .Z(n38720) );
  OR U39748 ( .A(n38720), .B(n38719), .Z(n38721) );
  AND U39749 ( .A(n38722), .B(n38721), .Z(n38880) );
  NAND U39750 ( .A(n38724), .B(n38723), .Z(n38728) );
  NAND U39751 ( .A(n38726), .B(n38725), .Z(n38727) );
  AND U39752 ( .A(n38728), .B(n38727), .Z(n38875) );
  NAND U39753 ( .A(n38730), .B(n38729), .Z(n38734) );
  NAND U39754 ( .A(n38732), .B(n38731), .Z(n38733) );
  NAND U39755 ( .A(n38734), .B(n38733), .Z(n38995) );
  NAND U39756 ( .A(n38736), .B(n38735), .Z(n38740) );
  NAND U39757 ( .A(n38738), .B(n38737), .Z(n38739) );
  NAND U39758 ( .A(n38740), .B(n38739), .Z(n38993) );
  AND U39759 ( .A(n38742), .B(n38741), .Z(n38746) );
  NAND U39760 ( .A(n38744), .B(n38743), .Z(n38745) );
  NANDN U39761 ( .A(n38746), .B(n38745), .Z(n38910) );
  NAND U39762 ( .A(n38748), .B(n38747), .Z(n38752) );
  NAND U39763 ( .A(n38750), .B(n38749), .Z(n38751) );
  NAND U39764 ( .A(n38752), .B(n38751), .Z(n38909) );
  XOR U39765 ( .A(n38910), .B(n38909), .Z(n38911) );
  AND U39766 ( .A(n38754), .B(n38753), .Z(n38758) );
  NANDN U39767 ( .A(n38756), .B(n38755), .Z(n38757) );
  NANDN U39768 ( .A(n38758), .B(n38757), .Z(n38923) );
  AND U39769 ( .A(x[480]), .B(y[8091]), .Z(n38977) );
  AND U39770 ( .A(x[507]), .B(y[8064]), .Z(n38976) );
  XOR U39771 ( .A(n38977), .B(n38976), .Z(n38979) );
  AND U39772 ( .A(x[506]), .B(y[8065]), .Z(n38984) );
  XOR U39773 ( .A(n38984), .B(o[411]), .Z(n38978) );
  XOR U39774 ( .A(n38979), .B(n38978), .Z(n38922) );
  AND U39775 ( .A(x[489]), .B(y[8082]), .Z(n38981) );
  AND U39776 ( .A(x[501]), .B(y[8070]), .Z(n38980) );
  XOR U39777 ( .A(n38981), .B(n38980), .Z(n38983) );
  AND U39778 ( .A(x[498]), .B(y[8073]), .Z(n38982) );
  XOR U39779 ( .A(n38983), .B(n38982), .Z(n38921) );
  XOR U39780 ( .A(n38922), .B(n38921), .Z(n38924) );
  XNOR U39781 ( .A(n38923), .B(n38924), .Z(n38912) );
  XOR U39782 ( .A(n38993), .B(n38994), .Z(n38996) );
  XOR U39783 ( .A(n38995), .B(n38996), .Z(n39014) );
  NAND U39784 ( .A(n38760), .B(n38759), .Z(n38764) );
  NAND U39785 ( .A(n38762), .B(n38761), .Z(n38763) );
  AND U39786 ( .A(n38764), .B(n38763), .Z(n39012) );
  NAND U39787 ( .A(n38766), .B(n38765), .Z(n38770) );
  NAND U39788 ( .A(n38768), .B(n38767), .Z(n38769) );
  AND U39789 ( .A(n38770), .B(n38769), .Z(n39011) );
  XOR U39790 ( .A(n39012), .B(n39011), .Z(n39013) );
  NAND U39791 ( .A(n38772), .B(n38771), .Z(n38776) );
  NAND U39792 ( .A(n38774), .B(n38773), .Z(n38775) );
  AND U39793 ( .A(n38776), .B(n38775), .Z(n39002) );
  NANDN U39794 ( .A(n38778), .B(n38777), .Z(n38782) );
  NANDN U39795 ( .A(n38780), .B(n38779), .Z(n38781) );
  AND U39796 ( .A(n38782), .B(n38781), .Z(n39000) );
  NAND U39797 ( .A(n38784), .B(n38783), .Z(n38788) );
  NAND U39798 ( .A(n38786), .B(n38785), .Z(n38787) );
  NAND U39799 ( .A(n38788), .B(n38787), .Z(n38989) );
  NAND U39800 ( .A(n38790), .B(n38789), .Z(n38794) );
  NAND U39801 ( .A(n38792), .B(n38791), .Z(n38793) );
  NAND U39802 ( .A(n38794), .B(n38793), .Z(n38987) );
  AND U39803 ( .A(x[499]), .B(y[8072]), .Z(n38969) );
  AND U39804 ( .A(x[505]), .B(y[8066]), .Z(n38968) );
  XOR U39805 ( .A(n38969), .B(n38968), .Z(n38971) );
  AND U39806 ( .A(x[486]), .B(y[8085]), .Z(n38970) );
  XOR U39807 ( .A(n38971), .B(n38970), .Z(n38961) );
  AND U39808 ( .A(x[495]), .B(y[8076]), .Z(n38941) );
  AND U39809 ( .A(x[482]), .B(y[8089]), .Z(n38940) );
  XOR U39810 ( .A(n38941), .B(n38940), .Z(n38943) );
  AND U39811 ( .A(x[483]), .B(y[8088]), .Z(n38942) );
  XOR U39812 ( .A(n38943), .B(n38942), .Z(n38960) );
  XOR U39813 ( .A(n38961), .B(n38960), .Z(n38962) );
  NAND U39814 ( .A(x[496]), .B(y[8075]), .Z(n38927) );
  XOR U39815 ( .A(n38927), .B(n38795), .Z(n38930) );
  XOR U39816 ( .A(n38929), .B(n38930), .Z(n38937) );
  AND U39817 ( .A(y[8078]), .B(x[493]), .Z(n38797) );
  AND U39818 ( .A(y[8079]), .B(x[492]), .Z(n38796) );
  XOR U39819 ( .A(n38797), .B(n38796), .Z(n38936) );
  XOR U39820 ( .A(n38937), .B(n38936), .Z(n38963) );
  AND U39821 ( .A(n38935), .B(n38798), .Z(n38802) );
  NAND U39822 ( .A(n38800), .B(n38799), .Z(n38801) );
  NANDN U39823 ( .A(n38802), .B(n38801), .Z(n38904) );
  NAND U39824 ( .A(n38804), .B(n38803), .Z(n38808) );
  NAND U39825 ( .A(n38806), .B(n38805), .Z(n38807) );
  NAND U39826 ( .A(n38808), .B(n38807), .Z(n38903) );
  XNOR U39827 ( .A(n38904), .B(n38903), .Z(n38906) );
  XOR U39828 ( .A(n38987), .B(n38988), .Z(n38990) );
  XOR U39829 ( .A(n38989), .B(n38990), .Z(n38999) );
  XOR U39830 ( .A(n39000), .B(n38999), .Z(n39001) );
  XOR U39831 ( .A(n39002), .B(n39001), .Z(n38891) );
  NAND U39832 ( .A(n38810), .B(n38809), .Z(n38814) );
  NAND U39833 ( .A(n38812), .B(n38811), .Z(n38813) );
  NAND U39834 ( .A(n38814), .B(n38813), .Z(n38893) );
  XOR U39835 ( .A(n38894), .B(n38893), .Z(n38888) );
  NAND U39836 ( .A(n38816), .B(n38815), .Z(n38820) );
  NAND U39837 ( .A(n38818), .B(n38817), .Z(n38819) );
  NAND U39838 ( .A(n38820), .B(n38819), .Z(n39007) );
  ANDN U39839 ( .B(n38822), .A(n38821), .Z(n38826) );
  NAND U39840 ( .A(n38824), .B(n38823), .Z(n38825) );
  NANDN U39841 ( .A(n38826), .B(n38825), .Z(n38949) );
  NAND U39842 ( .A(n38828), .B(n38827), .Z(n38832) );
  NAND U39843 ( .A(n38830), .B(n38829), .Z(n38831) );
  NAND U39844 ( .A(n38832), .B(n38831), .Z(n38948) );
  XOR U39845 ( .A(n38949), .B(n38948), .Z(n38950) );
  AND U39846 ( .A(x[488]), .B(y[8084]), .Z(n38986) );
  NAND U39847 ( .A(n38833), .B(n38986), .Z(n38837) );
  NAND U39848 ( .A(n38835), .B(n38834), .Z(n38836) );
  NAND U39849 ( .A(n38837), .B(n38836), .Z(n38917) );
  AND U39850 ( .A(x[494]), .B(y[8077]), .Z(n38945) );
  AND U39851 ( .A(x[481]), .B(y[8090]), .Z(n38944) );
  XOR U39852 ( .A(n38945), .B(n38944), .Z(n38947) );
  ANDN U39853 ( .B(o[410]), .A(n38838), .Z(n38946) );
  XOR U39854 ( .A(n38947), .B(n38946), .Z(n38916) );
  AND U39855 ( .A(x[497]), .B(y[8074]), .Z(n38973) );
  AND U39856 ( .A(x[484]), .B(y[8087]), .Z(n38972) );
  XOR U39857 ( .A(n38973), .B(n38972), .Z(n38975) );
  AND U39858 ( .A(x[485]), .B(y[8086]), .Z(n38974) );
  XOR U39859 ( .A(n38975), .B(n38974), .Z(n38915) );
  XOR U39860 ( .A(n38916), .B(n38915), .Z(n38918) );
  XNOR U39861 ( .A(n38917), .B(n38918), .Z(n38951) );
  NAND U39862 ( .A(n38840), .B(n38839), .Z(n38844) );
  NAND U39863 ( .A(n38842), .B(n38841), .Z(n38843) );
  NAND U39864 ( .A(n38844), .B(n38843), .Z(n38956) );
  AND U39865 ( .A(y[8067]), .B(x[504]), .Z(n38846) );
  NAND U39866 ( .A(y[8071]), .B(x[500]), .Z(n38845) );
  XNOR U39867 ( .A(n38846), .B(n38845), .Z(n38967) );
  AND U39868 ( .A(x[487]), .B(y[8084]), .Z(n38966) );
  XOR U39869 ( .A(n38967), .B(n38966), .Z(n38955) );
  AND U39870 ( .A(x[488]), .B(y[8083]), .Z(n38932) );
  AND U39871 ( .A(x[503]), .B(y[8068]), .Z(n38931) );
  XOR U39872 ( .A(n38932), .B(n38931), .Z(n38934) );
  AND U39873 ( .A(x[502]), .B(y[8069]), .Z(n38933) );
  XOR U39874 ( .A(n38934), .B(n38933), .Z(n38954) );
  XOR U39875 ( .A(n38955), .B(n38954), .Z(n38957) );
  XNOR U39876 ( .A(n38956), .B(n38957), .Z(n39006) );
  XOR U39877 ( .A(n39007), .B(n39008), .Z(n38898) );
  NAND U39878 ( .A(n38848), .B(n38847), .Z(n38852) );
  NAND U39879 ( .A(n38850), .B(n38849), .Z(n38851) );
  NAND U39880 ( .A(n38852), .B(n38851), .Z(n38897) );
  NAND U39881 ( .A(n38854), .B(n38853), .Z(n38858) );
  NAND U39882 ( .A(n38856), .B(n38855), .Z(n38857) );
  AND U39883 ( .A(n38858), .B(n38857), .Z(n38899) );
  XNOR U39884 ( .A(n38900), .B(n38899), .Z(n38886) );
  NAND U39885 ( .A(n38860), .B(n38859), .Z(n38864) );
  NAND U39886 ( .A(n38862), .B(n38861), .Z(n38863) );
  AND U39887 ( .A(n38864), .B(n38863), .Z(n38885) );
  XOR U39888 ( .A(n38886), .B(n38885), .Z(n38887) );
  XNOR U39889 ( .A(n38888), .B(n38887), .Z(n38873) );
  NAND U39890 ( .A(n38866), .B(n38865), .Z(n38870) );
  NAND U39891 ( .A(n38868), .B(n38867), .Z(n38869) );
  AND U39892 ( .A(n38870), .B(n38869), .Z(n38872) );
  XOR U39893 ( .A(n38873), .B(n38872), .Z(n38874) );
  XOR U39894 ( .A(n38875), .B(n38874), .Z(n38881) );
  XNOR U39895 ( .A(n38880), .B(n38881), .Z(n38871) );
  XOR U39896 ( .A(n38878), .B(n38871), .Z(N828) );
  NAND U39897 ( .A(n38873), .B(n38872), .Z(n38877) );
  NAND U39898 ( .A(n38875), .B(n38874), .Z(n38876) );
  NAND U39899 ( .A(n38877), .B(n38876), .Z(n39151) );
  IV U39900 ( .A(n39151), .Z(n39149) );
  OR U39901 ( .A(n38880), .B(n38878), .Z(n38884) );
  ANDN U39902 ( .B(n38880), .A(n38879), .Z(n38882) );
  OR U39903 ( .A(n38882), .B(n38881), .Z(n38883) );
  AND U39904 ( .A(n38884), .B(n38883), .Z(n39150) );
  NAND U39905 ( .A(n38886), .B(n38885), .Z(n38890) );
  NAND U39906 ( .A(n38888), .B(n38887), .Z(n38889) );
  NAND U39907 ( .A(n38890), .B(n38889), .Z(n39144) );
  NANDN U39908 ( .A(n38892), .B(n38891), .Z(n38896) );
  NAND U39909 ( .A(n38894), .B(n38893), .Z(n38895) );
  NAND U39910 ( .A(n38896), .B(n38895), .Z(n39143) );
  XOR U39911 ( .A(n39144), .B(n39143), .Z(n39146) );
  NANDN U39912 ( .A(n38898), .B(n38897), .Z(n38902) );
  NAND U39913 ( .A(n38900), .B(n38899), .Z(n38901) );
  AND U39914 ( .A(n38902), .B(n38901), .Z(n39018) );
  NAND U39915 ( .A(n38904), .B(n38903), .Z(n38908) );
  NANDN U39916 ( .A(n38906), .B(n38905), .Z(n38907) );
  NAND U39917 ( .A(n38908), .B(n38907), .Z(n39042) );
  NAND U39918 ( .A(n38910), .B(n38909), .Z(n38914) );
  NANDN U39919 ( .A(n38912), .B(n38911), .Z(n38913) );
  NAND U39920 ( .A(n38914), .B(n38913), .Z(n39121) );
  NAND U39921 ( .A(n38916), .B(n38915), .Z(n38920) );
  NAND U39922 ( .A(n38918), .B(n38917), .Z(n38919) );
  NAND U39923 ( .A(n38920), .B(n38919), .Z(n39120) );
  NAND U39924 ( .A(n38922), .B(n38921), .Z(n38926) );
  NAND U39925 ( .A(n38924), .B(n38923), .Z(n38925) );
  NAND U39926 ( .A(n38926), .B(n38925), .Z(n39119) );
  XOR U39927 ( .A(n39120), .B(n39119), .Z(n39122) );
  XOR U39928 ( .A(n39121), .B(n39122), .Z(n39043) );
  XOR U39929 ( .A(n39042), .B(n39043), .Z(n39045) );
  AND U39930 ( .A(x[495]), .B(y[8077]), .Z(n39100) );
  NAND U39931 ( .A(x[507]), .B(y[8065]), .Z(n39088) );
  XNOR U39932 ( .A(o[412]), .B(n39088), .Z(n39098) );
  AND U39933 ( .A(x[506]), .B(y[8066]), .Z(n39097) );
  XOR U39934 ( .A(n39098), .B(n39097), .Z(n39099) );
  XOR U39935 ( .A(n39100), .B(n39099), .Z(n39090) );
  AND U39936 ( .A(x[487]), .B(y[8085]), .Z(n39078) );
  AND U39937 ( .A(x[492]), .B(y[8080]), .Z(n39077) );
  XOR U39938 ( .A(n39078), .B(n39077), .Z(n39080) );
  AND U39939 ( .A(x[491]), .B(y[8081]), .Z(n39079) );
  XNOR U39940 ( .A(n39080), .B(n39079), .Z(n39089) );
  XNOR U39941 ( .A(n39090), .B(n39089), .Z(n39092) );
  XOR U39942 ( .A(n39092), .B(n39091), .Z(n39126) );
  AND U39943 ( .A(x[497]), .B(y[8075]), .Z(n39053) );
  AND U39944 ( .A(x[502]), .B(y[8070]), .Z(n39052) );
  XOR U39945 ( .A(n39053), .B(n39052), .Z(n39055) );
  AND U39946 ( .A(x[484]), .B(y[8088]), .Z(n39054) );
  XOR U39947 ( .A(n39055), .B(n39054), .Z(n39104) );
  AND U39948 ( .A(x[486]), .B(y[8086]), .Z(n39241) );
  AND U39949 ( .A(x[499]), .B(y[8073]), .Z(n39081) );
  XOR U39950 ( .A(n39241), .B(n39081), .Z(n39083) );
  XOR U39951 ( .A(n39083), .B(n39082), .Z(n39103) );
  XOR U39952 ( .A(n39104), .B(n39103), .Z(n39106) );
  XOR U39953 ( .A(n39106), .B(n39105), .Z(n39125) );
  NAND U39954 ( .A(n39094), .B(n38935), .Z(n38939) );
  NANDN U39955 ( .A(n38937), .B(n38936), .Z(n38938) );
  NAND U39956 ( .A(n38939), .B(n38938), .Z(n39067) );
  XOR U39957 ( .A(n39065), .B(n39066), .Z(n39068) );
  XOR U39958 ( .A(n39067), .B(n39068), .Z(n39127) );
  XOR U39959 ( .A(n39128), .B(n39127), .Z(n39044) );
  XNOR U39960 ( .A(n39045), .B(n39044), .Z(n39039) );
  NAND U39961 ( .A(n38949), .B(n38948), .Z(n38953) );
  NANDN U39962 ( .A(n38951), .B(n38950), .Z(n38952) );
  NAND U39963 ( .A(n38953), .B(n38952), .Z(n39109) );
  NAND U39964 ( .A(n38955), .B(n38954), .Z(n38959) );
  NAND U39965 ( .A(n38957), .B(n38956), .Z(n38958) );
  NAND U39966 ( .A(n38959), .B(n38958), .Z(n39108) );
  NAND U39967 ( .A(n38961), .B(n38960), .Z(n38965) );
  NANDN U39968 ( .A(n38963), .B(n38962), .Z(n38964) );
  NAND U39969 ( .A(n38965), .B(n38964), .Z(n39107) );
  XOR U39970 ( .A(n39108), .B(n39107), .Z(n39110) );
  XOR U39971 ( .A(n39109), .B(n39110), .Z(n39037) );
  AND U39972 ( .A(x[504]), .B(y[8071]), .Z(n39373) );
  AND U39973 ( .A(x[505]), .B(y[8067]), .Z(n39075) );
  XOR U39974 ( .A(n39076), .B(n39075), .Z(n39074) );
  AND U39975 ( .A(x[481]), .B(y[8091]), .Z(n39073) );
  XOR U39976 ( .A(n39074), .B(n39073), .Z(n39140) );
  AND U39977 ( .A(x[496]), .B(y[8076]), .Z(n39070) );
  AND U39978 ( .A(x[504]), .B(y[8068]), .Z(n39069) );
  XOR U39979 ( .A(n39070), .B(n39069), .Z(n39072) );
  AND U39980 ( .A(x[482]), .B(y[8090]), .Z(n39071) );
  XOR U39981 ( .A(n39072), .B(n39071), .Z(n39139) );
  XOR U39982 ( .A(n39140), .B(n39139), .Z(n39142) );
  XOR U39983 ( .A(n39141), .B(n39142), .Z(n39116) );
  AND U39984 ( .A(x[483]), .B(y[8089]), .Z(n39093) );
  XOR U39985 ( .A(n39094), .B(n39093), .Z(n39096) );
  AND U39986 ( .A(x[503]), .B(y[8069]), .Z(n39095) );
  XOR U39987 ( .A(n39096), .B(n39095), .Z(n39136) );
  AND U39988 ( .A(x[485]), .B(y[8087]), .Z(n39085) );
  AND U39989 ( .A(x[501]), .B(y[8071]), .Z(n39084) );
  XOR U39990 ( .A(n39085), .B(n39084), .Z(n39087) );
  AND U39991 ( .A(x[500]), .B(y[8072]), .Z(n39086) );
  XOR U39992 ( .A(n39087), .B(n39086), .Z(n39135) );
  XOR U39993 ( .A(n39136), .B(n39135), .Z(n39138) );
  XOR U39994 ( .A(n39137), .B(n39138), .Z(n39114) );
  XOR U39995 ( .A(n39131), .B(n39132), .Z(n39134) );
  AND U39996 ( .A(n38984), .B(o[411]), .Z(n39059) );
  AND U39997 ( .A(x[480]), .B(y[8092]), .Z(n39057) );
  AND U39998 ( .A(x[508]), .B(y[8064]), .Z(n39056) );
  XOR U39999 ( .A(n39057), .B(n39056), .Z(n39058) );
  XOR U40000 ( .A(n39059), .B(n39058), .Z(n39049) );
  NAND U40001 ( .A(y[8082]), .B(x[490]), .Z(n38985) );
  XNOR U40002 ( .A(n38986), .B(n38985), .Z(n39062) );
  AND U40003 ( .A(x[489]), .B(y[8083]), .Z(n39061) );
  XOR U40004 ( .A(n39062), .B(n39061), .Z(n39048) );
  XOR U40005 ( .A(n39049), .B(n39048), .Z(n39051) );
  XOR U40006 ( .A(n39050), .B(n39051), .Z(n39133) );
  XNOR U40007 ( .A(n39134), .B(n39133), .Z(n39113) );
  XNOR U40008 ( .A(n39039), .B(n39038), .Z(n39032) );
  NAND U40009 ( .A(n38988), .B(n38987), .Z(n38992) );
  NAND U40010 ( .A(n38990), .B(n38989), .Z(n38991) );
  NAND U40011 ( .A(n38992), .B(n38991), .Z(n39031) );
  NAND U40012 ( .A(n38994), .B(n38993), .Z(n38998) );
  NAND U40013 ( .A(n38996), .B(n38995), .Z(n38997) );
  NAND U40014 ( .A(n38998), .B(n38997), .Z(n39030) );
  XNOR U40015 ( .A(n39031), .B(n39030), .Z(n39033) );
  XNOR U40016 ( .A(n39018), .B(n39019), .Z(n39020) );
  NAND U40017 ( .A(n39000), .B(n38999), .Z(n39004) );
  NAND U40018 ( .A(n39002), .B(n39001), .Z(n39003) );
  NAND U40019 ( .A(n39004), .B(n39003), .Z(n39026) );
  NANDN U40020 ( .A(n39006), .B(n39005), .Z(n39010) );
  NAND U40021 ( .A(n39008), .B(n39007), .Z(n39009) );
  NAND U40022 ( .A(n39010), .B(n39009), .Z(n39024) );
  NAND U40023 ( .A(n39012), .B(n39011), .Z(n39016) );
  NANDN U40024 ( .A(n39014), .B(n39013), .Z(n39015) );
  AND U40025 ( .A(n39016), .B(n39015), .Z(n39025) );
  XNOR U40026 ( .A(n39024), .B(n39025), .Z(n39027) );
  XNOR U40027 ( .A(n39020), .B(n39021), .Z(n39145) );
  XOR U40028 ( .A(n39146), .B(n39145), .Z(n39152) );
  XNOR U40029 ( .A(n39150), .B(n39152), .Z(n39017) );
  XOR U40030 ( .A(n39149), .B(n39017), .Z(N829) );
  NANDN U40031 ( .A(n39019), .B(n39018), .Z(n39023) );
  NANDN U40032 ( .A(n39021), .B(n39020), .Z(n39022) );
  NAND U40033 ( .A(n39023), .B(n39022), .Z(n39162) );
  NAND U40034 ( .A(n39025), .B(n39024), .Z(n39029) );
  NANDN U40035 ( .A(n39027), .B(n39026), .Z(n39028) );
  NAND U40036 ( .A(n39029), .B(n39028), .Z(n39160) );
  NAND U40037 ( .A(n39031), .B(n39030), .Z(n39035) );
  NANDN U40038 ( .A(n39033), .B(n39032), .Z(n39034) );
  NAND U40039 ( .A(n39035), .B(n39034), .Z(n39166) );
  NANDN U40040 ( .A(n39037), .B(n39036), .Z(n39041) );
  NAND U40041 ( .A(n39039), .B(n39038), .Z(n39040) );
  AND U40042 ( .A(n39041), .B(n39040), .Z(n39167) );
  XOR U40043 ( .A(n39166), .B(n39167), .Z(n39169) );
  NAND U40044 ( .A(n39043), .B(n39042), .Z(n39047) );
  NAND U40045 ( .A(n39045), .B(n39044), .Z(n39046) );
  NAND U40046 ( .A(n39047), .B(n39046), .Z(n39178) );
  XOR U40047 ( .A(n39306), .B(n39307), .Z(n39308) );
  AND U40048 ( .A(x[490]), .B(y[8084]), .Z(n39304) );
  NAND U40049 ( .A(n39060), .B(n39304), .Z(n39064) );
  NAND U40050 ( .A(n39062), .B(n39061), .Z(n39063) );
  NAND U40051 ( .A(n39064), .B(n39063), .Z(n39279) );
  AND U40052 ( .A(x[492]), .B(y[8081]), .Z(n39481) );
  AND U40053 ( .A(x[481]), .B(y[8092]), .Z(n39252) );
  XOR U40054 ( .A(n39481), .B(n39252), .Z(n39254) );
  AND U40055 ( .A(x[502]), .B(y[8071]), .Z(n39253) );
  XOR U40056 ( .A(n39254), .B(n39253), .Z(n39278) );
  AND U40057 ( .A(x[495]), .B(y[8078]), .Z(n39255) );
  XOR U40058 ( .A(n39487), .B(n39255), .Z(n39257) );
  XOR U40059 ( .A(n39278), .B(n39277), .Z(n39280) );
  XNOR U40060 ( .A(n39279), .B(n39280), .Z(n39309) );
  XOR U40061 ( .A(n39308), .B(n39309), .Z(n39273) );
  XOR U40062 ( .A(n39274), .B(n39273), .Z(n39276) );
  XOR U40063 ( .A(n39276), .B(n39275), .Z(n39272) );
  XOR U40064 ( .A(n39283), .B(n39284), .Z(n39285) );
  AND U40065 ( .A(x[483]), .B(y[8090]), .Z(n39236) );
  AND U40066 ( .A(x[497]), .B(y[8076]), .Z(n39235) );
  XOR U40067 ( .A(n39236), .B(n39235), .Z(n39238) );
  AND U40068 ( .A(x[491]), .B(y[8082]), .Z(n39237) );
  XOR U40069 ( .A(n39238), .B(n39237), .Z(n39201) );
  AND U40070 ( .A(x[493]), .B(y[8080]), .Z(n39230) );
  AND U40071 ( .A(x[504]), .B(y[8069]), .Z(n39354) );
  XOR U40072 ( .A(n39230), .B(n39354), .Z(n39232) );
  AND U40073 ( .A(x[503]), .B(y[8070]), .Z(n39231) );
  XOR U40074 ( .A(n39232), .B(n39231), .Z(n39200) );
  XOR U40075 ( .A(n39201), .B(n39200), .Z(n39202) );
  XNOR U40076 ( .A(n39203), .B(n39202), .Z(n39286) );
  XOR U40077 ( .A(n39285), .B(n39286), .Z(n39192) );
  AND U40078 ( .A(x[506]), .B(y[8067]), .Z(n39248) );
  XOR U40079 ( .A(n39249), .B(n39248), .Z(n39251) );
  AND U40080 ( .A(x[505]), .B(y[8068]), .Z(n39250) );
  XOR U40081 ( .A(n39251), .B(n39250), .Z(n39288) );
  AND U40082 ( .A(x[508]), .B(y[8065]), .Z(n39263) );
  XOR U40083 ( .A(o[413]), .B(n39263), .Z(n39301) );
  AND U40084 ( .A(x[480]), .B(y[8093]), .Z(n39299) );
  AND U40085 ( .A(x[509]), .B(y[8064]), .Z(n39298) );
  XOR U40086 ( .A(n39299), .B(n39298), .Z(n39300) );
  XOR U40087 ( .A(n39301), .B(n39300), .Z(n39287) );
  XOR U40088 ( .A(n39288), .B(n39287), .Z(n39289) );
  XOR U40089 ( .A(n39290), .B(n39289), .Z(n39190) );
  AND U40090 ( .A(x[482]), .B(y[8091]), .Z(n39211) );
  XOR U40091 ( .A(n39211), .B(n39210), .Z(n39212) );
  XOR U40092 ( .A(n39213), .B(n39212), .Z(n39223) );
  ANDN U40093 ( .B(o[412]), .A(n39088), .Z(n39217) );
  AND U40094 ( .A(x[496]), .B(y[8077]), .Z(n39215) );
  AND U40095 ( .A(x[507]), .B(y[8066]), .Z(n39214) );
  XOR U40096 ( .A(n39215), .B(n39214), .Z(n39216) );
  XOR U40097 ( .A(n39217), .B(n39216), .Z(n39222) );
  XOR U40098 ( .A(n39223), .B(n39222), .Z(n39226) );
  XOR U40099 ( .A(n39225), .B(n39226), .Z(n39191) );
  XNOR U40100 ( .A(n39190), .B(n39191), .Z(n39193) );
  XOR U40101 ( .A(n39192), .B(n39193), .Z(n39196) );
  XOR U40102 ( .A(n39218), .B(n39219), .Z(n39221) );
  AND U40103 ( .A(y[8087]), .B(x[486]), .Z(n39102) );
  NAND U40104 ( .A(y[8086]), .B(x[487]), .Z(n39101) );
  XNOR U40105 ( .A(n39102), .B(n39101), .Z(n39243) );
  AND U40106 ( .A(x[488]), .B(y[8085]), .Z(n39242) );
  XOR U40107 ( .A(n39243), .B(n39242), .Z(n39293) );
  AND U40108 ( .A(x[489]), .B(y[8084]), .Z(n39349) );
  XOR U40109 ( .A(n39293), .B(n39349), .Z(n39295) );
  AND U40110 ( .A(x[485]), .B(y[8088]), .Z(n39206) );
  AND U40111 ( .A(x[484]), .B(y[8089]), .Z(n39205) );
  AND U40112 ( .A(x[490]), .B(y[8083]), .Z(n39204) );
  XNOR U40113 ( .A(n39205), .B(n39204), .Z(n39207) );
  XNOR U40114 ( .A(n39206), .B(n39207), .Z(n39294) );
  XOR U40115 ( .A(n39295), .B(n39294), .Z(n39220) );
  XOR U40116 ( .A(n39221), .B(n39220), .Z(n39195) );
  XOR U40117 ( .A(n39194), .B(n39195), .Z(n39197) );
  XOR U40118 ( .A(n39196), .B(n39197), .Z(n39269) );
  XOR U40119 ( .A(n39269), .B(n39270), .Z(n39271) );
  XNOR U40120 ( .A(n39272), .B(n39271), .Z(n39179) );
  XOR U40121 ( .A(n39178), .B(n39179), .Z(n39181) );
  NAND U40122 ( .A(n39108), .B(n39107), .Z(n39112) );
  NAND U40123 ( .A(n39110), .B(n39109), .Z(n39111) );
  NAND U40124 ( .A(n39112), .B(n39111), .Z(n39172) );
  NANDN U40125 ( .A(n39114), .B(n39113), .Z(n39118) );
  NANDN U40126 ( .A(n39116), .B(n39115), .Z(n39117) );
  AND U40127 ( .A(n39118), .B(n39117), .Z(n39173) );
  XOR U40128 ( .A(n39172), .B(n39173), .Z(n39175) );
  NAND U40129 ( .A(n39120), .B(n39119), .Z(n39124) );
  NAND U40130 ( .A(n39122), .B(n39121), .Z(n39123) );
  NAND U40131 ( .A(n39124), .B(n39123), .Z(n39186) );
  NANDN U40132 ( .A(n39126), .B(n39125), .Z(n39130) );
  NAND U40133 ( .A(n39128), .B(n39127), .Z(n39129) );
  NAND U40134 ( .A(n39130), .B(n39129), .Z(n39184) );
  XOR U40135 ( .A(n39265), .B(n39266), .Z(n39268) );
  XOR U40136 ( .A(n39267), .B(n39268), .Z(n39185) );
  XOR U40137 ( .A(n39184), .B(n39185), .Z(n39187) );
  XOR U40138 ( .A(n39186), .B(n39187), .Z(n39174) );
  XOR U40139 ( .A(n39175), .B(n39174), .Z(n39180) );
  XOR U40140 ( .A(n39181), .B(n39180), .Z(n39168) );
  XOR U40141 ( .A(n39169), .B(n39168), .Z(n39161) );
  XNOR U40142 ( .A(n39160), .B(n39161), .Z(n39163) );
  XOR U40143 ( .A(n39162), .B(n39163), .Z(n39159) );
  NAND U40144 ( .A(n39144), .B(n39143), .Z(n39148) );
  NAND U40145 ( .A(n39146), .B(n39145), .Z(n39147) );
  NAND U40146 ( .A(n39148), .B(n39147), .Z(n39158) );
  NANDN U40147 ( .A(n39149), .B(n39150), .Z(n39155) );
  NOR U40148 ( .A(n39151), .B(n39150), .Z(n39153) );
  OR U40149 ( .A(n39153), .B(n39152), .Z(n39154) );
  AND U40150 ( .A(n39155), .B(n39154), .Z(n39157) );
  XOR U40151 ( .A(n39158), .B(n39157), .Z(n39156) );
  XNOR U40152 ( .A(n39159), .B(n39156), .Z(N830) );
  NAND U40153 ( .A(n39161), .B(n39160), .Z(n39165) );
  NANDN U40154 ( .A(n39163), .B(n39162), .Z(n39164) );
  NAND U40155 ( .A(n39165), .B(n39164), .Z(n39574) );
  NAND U40156 ( .A(n39167), .B(n39166), .Z(n39171) );
  NAND U40157 ( .A(n39169), .B(n39168), .Z(n39170) );
  NAND U40158 ( .A(n39171), .B(n39170), .Z(n39579) );
  NAND U40159 ( .A(n39173), .B(n39172), .Z(n39177) );
  NAND U40160 ( .A(n39175), .B(n39174), .Z(n39176) );
  AND U40161 ( .A(n39177), .B(n39176), .Z(n39586) );
  NAND U40162 ( .A(n39179), .B(n39178), .Z(n39183) );
  NAND U40163 ( .A(n39181), .B(n39180), .Z(n39182) );
  AND U40164 ( .A(n39183), .B(n39182), .Z(n39585) );
  XOR U40165 ( .A(n39586), .B(n39585), .Z(n39588) );
  NAND U40166 ( .A(n39185), .B(n39184), .Z(n39189) );
  NAND U40167 ( .A(n39187), .B(n39186), .Z(n39188) );
  AND U40168 ( .A(n39189), .B(n39188), .Z(n39587) );
  XOR U40169 ( .A(n39588), .B(n39587), .Z(n39581) );
  NANDN U40170 ( .A(n39195), .B(n39194), .Z(n39199) );
  NANDN U40171 ( .A(n39197), .B(n39196), .Z(n39198) );
  AND U40172 ( .A(n39199), .B(n39198), .Z(n39550) );
  NAND U40173 ( .A(n39205), .B(n39204), .Z(n39209) );
  NANDN U40174 ( .A(n39207), .B(n39206), .Z(n39208) );
  NAND U40175 ( .A(n39209), .B(n39208), .Z(n39326) );
  AND U40176 ( .A(x[486]), .B(y[8088]), .Z(n39358) );
  AND U40177 ( .A(x[485]), .B(y[8089]), .Z(n39360) );
  AND U40178 ( .A(x[499]), .B(y[8075]), .Z(n39359) );
  XOR U40179 ( .A(n39360), .B(n39359), .Z(n39357) );
  XNOR U40180 ( .A(n39358), .B(n39357), .Z(n39471) );
  AND U40181 ( .A(x[484]), .B(y[8090]), .Z(n39424) );
  AND U40182 ( .A(x[483]), .B(y[8091]), .Z(n39426) );
  AND U40183 ( .A(x[498]), .B(y[8076]), .Z(n39425) );
  XOR U40184 ( .A(n39426), .B(n39425), .Z(n39423) );
  XOR U40185 ( .A(n39424), .B(n39423), .Z(n39468) );
  XOR U40186 ( .A(n39471), .B(n39470), .Z(n39325) );
  XOR U40187 ( .A(n39326), .B(n39325), .Z(n39324) );
  XOR U40188 ( .A(n39324), .B(n39323), .Z(n39314) );
  XOR U40189 ( .A(n39311), .B(n39310), .Z(n39553) );
  IV U40190 ( .A(n39222), .Z(n39224) );
  NANDN U40191 ( .A(n39224), .B(n39223), .Z(n39229) );
  IV U40192 ( .A(n39225), .Z(n39227) );
  NANDN U40193 ( .A(n39227), .B(n39226), .Z(n39228) );
  NAND U40194 ( .A(n39229), .B(n39228), .Z(n39534) );
  NAND U40195 ( .A(n39230), .B(n39354), .Z(n39234) );
  NAND U40196 ( .A(n39232), .B(n39231), .Z(n39233) );
  NAND U40197 ( .A(n39234), .B(n39233), .Z(n39320) );
  NAND U40198 ( .A(n39236), .B(n39235), .Z(n39240) );
  NAND U40199 ( .A(n39238), .B(n39237), .Z(n39239) );
  AND U40200 ( .A(n39240), .B(n39239), .Z(n39330) );
  AND U40201 ( .A(x[480]), .B(y[8094]), .Z(n39366) );
  AND U40202 ( .A(x[509]), .B(y[8065]), .Z(n39371) );
  XOR U40203 ( .A(o[414]), .B(n39371), .Z(n39368) );
  AND U40204 ( .A(x[510]), .B(y[8064]), .Z(n39367) );
  XOR U40205 ( .A(n39368), .B(n39367), .Z(n39365) );
  XOR U40206 ( .A(n39366), .B(n39365), .Z(n39332) );
  AND U40207 ( .A(x[500]), .B(y[8074]), .Z(n39500) );
  AND U40208 ( .A(x[488]), .B(y[8086]), .Z(n39498) );
  XNOR U40209 ( .A(n39499), .B(n39498), .Z(n39331) );
  XNOR U40210 ( .A(n39330), .B(n39329), .Z(n39319) );
  XOR U40211 ( .A(n39320), .B(n39319), .Z(n39317) );
  AND U40212 ( .A(x[487]), .B(y[8087]), .Z(n39485) );
  NAND U40213 ( .A(n39241), .B(n39485), .Z(n39245) );
  NAND U40214 ( .A(n39243), .B(n39242), .Z(n39244) );
  AND U40215 ( .A(n39245), .B(n39244), .Z(n39339) );
  AND U40216 ( .A(y[8073]), .B(x[501]), .Z(n39247) );
  AND U40217 ( .A(y[8072]), .B(x[502]), .Z(n39246) );
  XOR U40218 ( .A(n39247), .B(n39246), .Z(n39484) );
  XOR U40219 ( .A(n39485), .B(n39484), .Z(n39342) );
  AND U40220 ( .A(x[497]), .B(y[8077]), .Z(n39493) );
  AND U40221 ( .A(x[482]), .B(y[8092]), .Z(n39495) );
  AND U40222 ( .A(x[506]), .B(y[8068]), .Z(n39494) );
  XOR U40223 ( .A(n39495), .B(n39494), .Z(n39492) );
  XNOR U40224 ( .A(n39493), .B(n39492), .Z(n39341) );
  XNOR U40225 ( .A(n39339), .B(n39340), .Z(n39318) );
  XNOR U40226 ( .A(n39317), .B(n39318), .Z(n39535) );
  XOR U40227 ( .A(n39534), .B(n39535), .Z(n39533) );
  IV U40228 ( .A(n39255), .Z(n39256) );
  NANDN U40229 ( .A(n39256), .B(n39487), .Z(n39260) );
  NANDN U40230 ( .A(n39258), .B(n39257), .Z(n39259) );
  AND U40231 ( .A(n39260), .B(n39259), .Z(n39336) );
  AND U40232 ( .A(x[503]), .B(y[8071]), .Z(n39353) );
  AND U40233 ( .A(y[8070]), .B(x[504]), .Z(n39262) );
  AND U40234 ( .A(y[8069]), .B(x[505]), .Z(n39261) );
  XOR U40235 ( .A(n39262), .B(n39261), .Z(n39352) );
  XOR U40236 ( .A(n39353), .B(n39352), .Z(n39338) );
  IV U40237 ( .A(n39338), .Z(n39264) );
  AND U40238 ( .A(x[508]), .B(y[8066]), .Z(n39438) );
  AND U40239 ( .A(x[496]), .B(y[8078]), .Z(n39437) );
  XOR U40240 ( .A(n39438), .B(n39437), .Z(n39435) );
  XNOR U40241 ( .A(n39436), .B(n39435), .Z(n39337) );
  XOR U40242 ( .A(n39264), .B(n39337), .Z(n39335) );
  XNOR U40243 ( .A(n39336), .B(n39335), .Z(n39345) );
  XOR U40244 ( .A(n39346), .B(n39345), .Z(n39344) );
  XOR U40245 ( .A(n39343), .B(n39344), .Z(n39532) );
  XOR U40246 ( .A(n39533), .B(n39532), .Z(n39552) );
  XNOR U40247 ( .A(n39550), .B(n39551), .Z(n39565) );
  NAND U40248 ( .A(n39278), .B(n39277), .Z(n39282) );
  NAND U40249 ( .A(n39280), .B(n39279), .Z(n39281) );
  AND U40250 ( .A(n39282), .B(n39281), .Z(n39519) );
  XOR U40251 ( .A(n39519), .B(n39518), .Z(n39517) );
  OR U40252 ( .A(n39288), .B(n39287), .Z(n39292) );
  NAND U40253 ( .A(n39290), .B(n39289), .Z(n39291) );
  NAND U40254 ( .A(n39292), .B(n39291), .Z(n39516) );
  XOR U40255 ( .A(n39517), .B(n39516), .Z(n39529) );
  NAND U40256 ( .A(n39293), .B(n39349), .Z(n39297) );
  NAND U40257 ( .A(n39295), .B(n39294), .Z(n39296) );
  AND U40258 ( .A(n39297), .B(n39296), .Z(n39512) );
  AND U40259 ( .A(y[8082]), .B(x[492]), .Z(n39302) );
  XOR U40260 ( .A(n39303), .B(n39302), .Z(n39478) );
  XOR U40261 ( .A(n39479), .B(n39478), .Z(n39348) );
  AND U40262 ( .A(y[8085]), .B(x[489]), .Z(n39305) );
  XOR U40263 ( .A(n39305), .B(n39304), .Z(n39347) );
  XOR U40264 ( .A(n39348), .B(n39347), .Z(n39465) );
  AND U40265 ( .A(x[507]), .B(y[8067]), .Z(n39432) );
  AND U40266 ( .A(x[481]), .B(y[8093]), .Z(n39431) );
  XOR U40267 ( .A(n39432), .B(n39431), .Z(n39429) );
  XOR U40268 ( .A(n39430), .B(n39429), .Z(n39464) );
  XOR U40269 ( .A(n39465), .B(n39464), .Z(n39462) );
  XOR U40270 ( .A(n39461), .B(n39462), .Z(n39513) );
  XNOR U40271 ( .A(n39510), .B(n39511), .Z(n39528) );
  XNOR U40272 ( .A(n39526), .B(n39527), .Z(n39547) );
  XOR U40273 ( .A(n39546), .B(n39547), .Z(n39544) );
  XOR U40274 ( .A(n39545), .B(n39544), .Z(n39582) );
  XOR U40275 ( .A(n39579), .B(n39580), .Z(n39571) );
  XNOR U40276 ( .A(n39572), .B(n39571), .Z(N831) );
  IV U40277 ( .A(n39310), .Z(n39312) );
  NANDN U40278 ( .A(n39312), .B(n39311), .Z(n39316) );
  NANDN U40279 ( .A(n39314), .B(n39313), .Z(n39315) );
  AND U40280 ( .A(n39316), .B(n39315), .Z(n39561) );
  NANDN U40281 ( .A(n39318), .B(n39317), .Z(n39322) );
  NAND U40282 ( .A(n39320), .B(n39319), .Z(n39321) );
  AND U40283 ( .A(n39322), .B(n39321), .Z(n39543) );
  NAND U40284 ( .A(n39324), .B(n39323), .Z(n39328) );
  NAND U40285 ( .A(n39326), .B(n39325), .Z(n39327) );
  AND U40286 ( .A(n39328), .B(n39327), .Z(n39525) );
  NAND U40287 ( .A(n39330), .B(n39329), .Z(n39334) );
  NANDN U40288 ( .A(n39332), .B(n39331), .Z(n39333) );
  AND U40289 ( .A(n39334), .B(n39333), .Z(n39509) );
  AND U40290 ( .A(x[490]), .B(y[8085]), .Z(n39394) );
  NAND U40291 ( .A(n39349), .B(n39394), .Z(n39350) );
  NAND U40292 ( .A(n39353), .B(n39352), .Z(n39356) );
  AND U40293 ( .A(x[505]), .B(y[8070]), .Z(n39372) );
  NAND U40294 ( .A(n39354), .B(n39372), .Z(n39355) );
  AND U40295 ( .A(n39356), .B(n39355), .Z(n39364) );
  NAND U40296 ( .A(n39358), .B(n39357), .Z(n39362) );
  NAND U40297 ( .A(n39360), .B(n39359), .Z(n39361) );
  NAND U40298 ( .A(n39362), .B(n39361), .Z(n39363) );
  XNOR U40299 ( .A(n39364), .B(n39363), .Z(n39422) );
  NAND U40300 ( .A(n39366), .B(n39365), .Z(n39370) );
  NAND U40301 ( .A(n39368), .B(n39367), .Z(n39369) );
  AND U40302 ( .A(n39370), .B(n39369), .Z(n39420) );
  AND U40303 ( .A(y[8069]), .B(x[506]), .Z(n39379) );
  AND U40304 ( .A(n39371), .B(o[414]), .Z(n39377) );
  XOR U40305 ( .A(n39372), .B(o[415]), .Z(n39375) );
  AND U40306 ( .A(x[502]), .B(y[8073]), .Z(n39486) );
  XNOR U40307 ( .A(n39373), .B(n39486), .Z(n39374) );
  XNOR U40308 ( .A(n39375), .B(n39374), .Z(n39376) );
  XNOR U40309 ( .A(n39377), .B(n39376), .Z(n39378) );
  XNOR U40310 ( .A(n39379), .B(n39378), .Z(n39418) );
  AND U40311 ( .A(y[8064]), .B(x[511]), .Z(n39385) );
  AND U40312 ( .A(y[8068]), .B(x[507]), .Z(n39381) );
  NAND U40313 ( .A(y[8094]), .B(x[481]), .Z(n39380) );
  XNOR U40314 ( .A(n39381), .B(n39380), .Z(n39382) );
  XNOR U40315 ( .A(n39383), .B(n39382), .Z(n39384) );
  XNOR U40316 ( .A(n39385), .B(n39384), .Z(n39408) );
  AND U40317 ( .A(y[8090]), .B(x[485]), .Z(n39387) );
  NAND U40318 ( .A(y[8088]), .B(x[487]), .Z(n39386) );
  XNOR U40319 ( .A(n39387), .B(n39386), .Z(n39398) );
  AND U40320 ( .A(y[8089]), .B(x[486]), .Z(n39389) );
  NAND U40321 ( .A(y[8077]), .B(x[498]), .Z(n39388) );
  XNOR U40322 ( .A(n39389), .B(n39388), .Z(n39393) );
  AND U40323 ( .A(y[8092]), .B(x[483]), .Z(n39391) );
  NAND U40324 ( .A(y[8091]), .B(x[484]), .Z(n39390) );
  XNOR U40325 ( .A(n39391), .B(n39390), .Z(n39392) );
  XOR U40326 ( .A(n39393), .B(n39392), .Z(n39396) );
  XNOR U40327 ( .A(n39480), .B(n39394), .Z(n39395) );
  XNOR U40328 ( .A(n39396), .B(n39395), .Z(n39397) );
  XOR U40329 ( .A(n39398), .B(n39397), .Z(n39406) );
  AND U40330 ( .A(y[8079]), .B(x[496]), .Z(n39400) );
  NAND U40331 ( .A(y[8075]), .B(x[500]), .Z(n39399) );
  XNOR U40332 ( .A(n39400), .B(n39399), .Z(n39404) );
  AND U40333 ( .A(y[8065]), .B(x[510]), .Z(n39402) );
  NAND U40334 ( .A(y[8066]), .B(x[509]), .Z(n39401) );
  XNOR U40335 ( .A(n39402), .B(n39401), .Z(n39403) );
  XNOR U40336 ( .A(n39404), .B(n39403), .Z(n39405) );
  XNOR U40337 ( .A(n39406), .B(n39405), .Z(n39407) );
  XOR U40338 ( .A(n39408), .B(n39407), .Z(n39416) );
  AND U40339 ( .A(y[8081]), .B(x[494]), .Z(n39410) );
  NAND U40340 ( .A(y[8095]), .B(x[480]), .Z(n39409) );
  XNOR U40341 ( .A(n39410), .B(n39409), .Z(n39414) );
  AND U40342 ( .A(y[8086]), .B(x[489]), .Z(n39412) );
  NAND U40343 ( .A(y[8067]), .B(x[508]), .Z(n39411) );
  XNOR U40344 ( .A(n39412), .B(n39411), .Z(n39413) );
  XNOR U40345 ( .A(n39414), .B(n39413), .Z(n39415) );
  XNOR U40346 ( .A(n39416), .B(n39415), .Z(n39417) );
  XNOR U40347 ( .A(n39418), .B(n39417), .Z(n39419) );
  XNOR U40348 ( .A(n39420), .B(n39419), .Z(n39421) );
  NAND U40349 ( .A(n39424), .B(n39423), .Z(n39428) );
  NAND U40350 ( .A(n39426), .B(n39425), .Z(n39427) );
  AND U40351 ( .A(n39428), .B(n39427), .Z(n39460) );
  NAND U40352 ( .A(n39430), .B(n39429), .Z(n39434) );
  NAND U40353 ( .A(n39432), .B(n39431), .Z(n39433) );
  AND U40354 ( .A(n39434), .B(n39433), .Z(n39442) );
  NAND U40355 ( .A(n39436), .B(n39435), .Z(n39440) );
  NAND U40356 ( .A(n39438), .B(n39437), .Z(n39439) );
  NAND U40357 ( .A(n39440), .B(n39439), .Z(n39441) );
  XNOR U40358 ( .A(n39442), .B(n39441), .Z(n39458) );
  AND U40359 ( .A(y[8093]), .B(x[482]), .Z(n39444) );
  NAND U40360 ( .A(y[8074]), .B(x[501]), .Z(n39443) );
  XNOR U40361 ( .A(n39444), .B(n39443), .Z(n39448) );
  AND U40362 ( .A(y[8072]), .B(x[503]), .Z(n39446) );
  NAND U40363 ( .A(y[8078]), .B(x[497]), .Z(n39445) );
  XNOR U40364 ( .A(n39446), .B(n39445), .Z(n39447) );
  XOR U40365 ( .A(n39448), .B(n39447), .Z(n39456) );
  AND U40366 ( .A(y[8076]), .B(x[499]), .Z(n39450) );
  NAND U40367 ( .A(y[8087]), .B(x[488]), .Z(n39449) );
  XNOR U40368 ( .A(n39450), .B(n39449), .Z(n39454) );
  AND U40369 ( .A(y[8084]), .B(x[491]), .Z(n39452) );
  NAND U40370 ( .A(y[8083]), .B(x[492]), .Z(n39451) );
  XNOR U40371 ( .A(n39452), .B(n39451), .Z(n39453) );
  XNOR U40372 ( .A(n39454), .B(n39453), .Z(n39455) );
  XNOR U40373 ( .A(n39456), .B(n39455), .Z(n39457) );
  XNOR U40374 ( .A(n39458), .B(n39457), .Z(n39459) );
  XNOR U40375 ( .A(n39460), .B(n39459), .Z(n39477) );
  IV U40376 ( .A(n39461), .Z(n39463) );
  NANDN U40377 ( .A(n39463), .B(n39462), .Z(n39467) );
  AND U40378 ( .A(n39465), .B(n39464), .Z(n39466) );
  ANDN U40379 ( .B(n39467), .A(n39466), .Z(n39475) );
  ANDN U40380 ( .B(n39469), .A(n39468), .Z(n39473) );
  ANDN U40381 ( .B(n39471), .A(n39470), .Z(n39472) );
  OR U40382 ( .A(n39473), .B(n39472), .Z(n39474) );
  XNOR U40383 ( .A(n39475), .B(n39474), .Z(n39476) );
  NAND U40384 ( .A(n39479), .B(n39478), .Z(n39483) );
  NAND U40385 ( .A(n39481), .B(n39480), .Z(n39482) );
  AND U40386 ( .A(n39483), .B(n39482), .Z(n39491) );
  NAND U40387 ( .A(n39485), .B(n39484), .Z(n39489) );
  NAND U40388 ( .A(n39487), .B(n39486), .Z(n39488) );
  NAND U40389 ( .A(n39489), .B(n39488), .Z(n39490) );
  XNOR U40390 ( .A(n39491), .B(n39490), .Z(n39507) );
  NAND U40391 ( .A(n39493), .B(n39492), .Z(n39497) );
  NAND U40392 ( .A(n39495), .B(n39494), .Z(n39496) );
  AND U40393 ( .A(n39497), .B(n39496), .Z(n39505) );
  NAND U40394 ( .A(n39499), .B(n39498), .Z(n39503) );
  NANDN U40395 ( .A(n39501), .B(n39500), .Z(n39502) );
  NAND U40396 ( .A(n39503), .B(n39502), .Z(n39504) );
  XNOR U40397 ( .A(n39505), .B(n39504), .Z(n39506) );
  XNOR U40398 ( .A(n39509), .B(n39508), .Z(n39523) );
  NAND U40399 ( .A(n39511), .B(n39510), .Z(n39515) );
  NANDN U40400 ( .A(n39513), .B(n39512), .Z(n39514) );
  AND U40401 ( .A(n39515), .B(n39514), .Z(n39521) );
  XNOR U40402 ( .A(n39521), .B(n39520), .Z(n39522) );
  XNOR U40403 ( .A(n39523), .B(n39522), .Z(n39524) );
  XNOR U40404 ( .A(n39525), .B(n39524), .Z(n39541) );
  NANDN U40405 ( .A(n39527), .B(n39526), .Z(n39531) );
  NANDN U40406 ( .A(n39529), .B(n39528), .Z(n39530) );
  AND U40407 ( .A(n39531), .B(n39530), .Z(n39539) );
  NAND U40408 ( .A(n39533), .B(n39532), .Z(n39537) );
  NAND U40409 ( .A(n39535), .B(n39534), .Z(n39536) );
  NAND U40410 ( .A(n39537), .B(n39536), .Z(n39538) );
  XNOR U40411 ( .A(n39539), .B(n39538), .Z(n39540) );
  XNOR U40412 ( .A(n39541), .B(n39540), .Z(n39542) );
  XNOR U40413 ( .A(n39543), .B(n39542), .Z(n39559) );
  NAND U40414 ( .A(n39545), .B(n39544), .Z(n39549) );
  NAND U40415 ( .A(n39547), .B(n39546), .Z(n39548) );
  AND U40416 ( .A(n39549), .B(n39548), .Z(n39557) );
  NANDN U40417 ( .A(n39551), .B(n39550), .Z(n39555) );
  NANDN U40418 ( .A(n39553), .B(n39552), .Z(n39554) );
  NAND U40419 ( .A(n39555), .B(n39554), .Z(n39556) );
  XNOR U40420 ( .A(n39557), .B(n39556), .Z(n39558) );
  XNOR U40421 ( .A(n39559), .B(n39558), .Z(n39560) );
  XNOR U40422 ( .A(n39561), .B(n39560), .Z(n39570) );
  IV U40423 ( .A(n39563), .Z(n39562) );
  OR U40424 ( .A(n39564), .B(n39562), .Z(n39568) );
  ANDN U40425 ( .B(n39564), .A(n39563), .Z(n39566) );
  NANDN U40426 ( .A(n39566), .B(n39565), .Z(n39567) );
  NAND U40427 ( .A(n39568), .B(n39567), .Z(n39569) );
  XNOR U40428 ( .A(n39570), .B(n39569), .Z(n39578) );
  NAND U40429 ( .A(n39572), .B(n39571), .Z(n39576) );
  NANDN U40430 ( .A(n39574), .B(n39573), .Z(n39575) );
  NAND U40431 ( .A(n39576), .B(n39575), .Z(n39577) );
  XNOR U40432 ( .A(n39578), .B(n39577), .Z(n39594) );
  NANDN U40433 ( .A(n39580), .B(n39579), .Z(n39584) );
  ANDN U40434 ( .B(n39582), .A(n39581), .Z(n39583) );
  ANDN U40435 ( .B(n39584), .A(n39583), .Z(n39592) );
  AND U40436 ( .A(n39586), .B(n39585), .Z(n39590) );
  AND U40437 ( .A(n39588), .B(n39587), .Z(n39589) );
  OR U40438 ( .A(n39590), .B(n39589), .Z(n39591) );
  XNOR U40439 ( .A(n39592), .B(n39591), .Z(n39593) );
  XNOR U40440 ( .A(n39594), .B(n39593), .Z(N832) );
  AND U40441 ( .A(x[480]), .B(y[8096]), .Z(n40246) );
  XOR U40442 ( .A(n40246), .B(o[416]), .Z(N865) );
  NAND U40443 ( .A(x[481]), .B(y[8096]), .Z(n39605) );
  AND U40444 ( .A(x[480]), .B(y[8097]), .Z(n39597) );
  XNOR U40445 ( .A(n39597), .B(o[417]), .Z(n39598) );
  XOR U40446 ( .A(n39605), .B(n39598), .Z(n39600) );
  NAND U40447 ( .A(n40246), .B(o[416]), .Z(n39599) );
  XNOR U40448 ( .A(n39600), .B(n39599), .Z(N866) );
  AND U40449 ( .A(y[8096]), .B(x[482]), .Z(n39596) );
  NAND U40450 ( .A(y[8097]), .B(x[481]), .Z(n39595) );
  XNOR U40451 ( .A(n39596), .B(n39595), .Z(n39606) );
  AND U40452 ( .A(n39597), .B(o[417]), .Z(n39607) );
  XOR U40453 ( .A(n39606), .B(n39607), .Z(n39612) );
  AND U40454 ( .A(x[480]), .B(y[8098]), .Z(n39604) );
  XOR U40455 ( .A(o[418]), .B(n39604), .Z(n39611) );
  XOR U40456 ( .A(n39610), .B(n39611), .Z(n39601) );
  XNOR U40457 ( .A(n39612), .B(n39601), .Z(N867) );
  AND U40458 ( .A(x[481]), .B(y[8098]), .Z(n39733) );
  AND U40459 ( .A(x[482]), .B(y[8097]), .Z(n39618) );
  XOR U40460 ( .A(n39618), .B(o[419]), .Z(n39625) );
  XOR U40461 ( .A(n39733), .B(n39625), .Z(n39627) );
  AND U40462 ( .A(y[8096]), .B(x[483]), .Z(n39603) );
  NAND U40463 ( .A(y[8099]), .B(x[480]), .Z(n39602) );
  XNOR U40464 ( .A(n39603), .B(n39602), .Z(n39615) );
  AND U40465 ( .A(n39604), .B(o[418]), .Z(n39614) );
  XOR U40466 ( .A(n39615), .B(n39614), .Z(n39626) );
  XNOR U40467 ( .A(n39627), .B(n39626), .Z(n39624) );
  NANDN U40468 ( .A(n39605), .B(n39618), .Z(n39609) );
  NAND U40469 ( .A(n39607), .B(n39606), .Z(n39608) );
  NAND U40470 ( .A(n39609), .B(n39608), .Z(n39623) );
  XOR U40471 ( .A(n39623), .B(n39622), .Z(n39613) );
  XNOR U40472 ( .A(n39624), .B(n39613), .Z(N868) );
  AND U40473 ( .A(x[483]), .B(y[8099]), .Z(n39680) );
  NAND U40474 ( .A(n40246), .B(n39680), .Z(n39617) );
  NAND U40475 ( .A(n39615), .B(n39614), .Z(n39616) );
  NAND U40476 ( .A(n39617), .B(n39616), .Z(n39652) );
  AND U40477 ( .A(n39618), .B(o[419]), .Z(n39641) );
  AND U40478 ( .A(y[8100]), .B(x[480]), .Z(n39620) );
  AND U40479 ( .A(y[8096]), .B(x[484]), .Z(n39619) );
  XOR U40480 ( .A(n39620), .B(n39619), .Z(n39640) );
  XOR U40481 ( .A(n39641), .B(n39640), .Z(n39651) );
  AND U40482 ( .A(y[8098]), .B(x[482]), .Z(n39760) );
  NAND U40483 ( .A(y[8099]), .B(x[481]), .Z(n39621) );
  XNOR U40484 ( .A(n39760), .B(n39621), .Z(n39637) );
  NAND U40485 ( .A(x[483]), .B(y[8097]), .Z(n39632) );
  XNOR U40486 ( .A(o[420]), .B(n39632), .Z(n39636) );
  XOR U40487 ( .A(n39637), .B(n39636), .Z(n39650) );
  XOR U40488 ( .A(n39651), .B(n39650), .Z(n39653) );
  XOR U40489 ( .A(n39652), .B(n39653), .Z(n39647) );
  NAND U40490 ( .A(n39733), .B(n39625), .Z(n39629) );
  NAND U40491 ( .A(n39627), .B(n39626), .Z(n39628) );
  NAND U40492 ( .A(n39629), .B(n39628), .Z(n39644) );
  XNOR U40493 ( .A(n39645), .B(n39644), .Z(n39646) );
  XOR U40494 ( .A(n39647), .B(n39646), .Z(N869) );
  AND U40495 ( .A(y[8098]), .B(x[483]), .Z(n39631) );
  NAND U40496 ( .A(y[8100]), .B(x[481]), .Z(n39630) );
  XNOR U40497 ( .A(n39631), .B(n39630), .Z(n39667) );
  AND U40498 ( .A(x[484]), .B(y[8097]), .Z(n39676) );
  XOR U40499 ( .A(n39676), .B(o[421]), .Z(n39666) );
  XOR U40500 ( .A(n39667), .B(n39666), .Z(n39670) );
  NAND U40501 ( .A(x[482]), .B(y[8099]), .Z(n39742) );
  ANDN U40502 ( .B(o[420]), .A(n39632), .Z(n39672) );
  AND U40503 ( .A(y[8096]), .B(x[485]), .Z(n39634) );
  NAND U40504 ( .A(y[8101]), .B(x[480]), .Z(n39633) );
  XNOR U40505 ( .A(n39634), .B(n39633), .Z(n39673) );
  XOR U40506 ( .A(n39672), .B(n39673), .Z(n39671) );
  XOR U40507 ( .A(n39742), .B(n39671), .Z(n39635) );
  XNOR U40508 ( .A(n39670), .B(n39635), .Z(n39663) );
  NANDN U40509 ( .A(n39742), .B(n39733), .Z(n39639) );
  NAND U40510 ( .A(n39637), .B(n39636), .Z(n39638) );
  NAND U40511 ( .A(n39639), .B(n39638), .Z(n39661) );
  AND U40512 ( .A(x[484]), .B(y[8100]), .Z(n40432) );
  NAND U40513 ( .A(n40432), .B(n40246), .Z(n39643) );
  NAND U40514 ( .A(n39641), .B(n39640), .Z(n39642) );
  NAND U40515 ( .A(n39643), .B(n39642), .Z(n39660) );
  XOR U40516 ( .A(n39661), .B(n39660), .Z(n39662) );
  XNOR U40517 ( .A(n39663), .B(n39662), .Z(n39659) );
  NANDN U40518 ( .A(n39645), .B(n39644), .Z(n39649) );
  NAND U40519 ( .A(n39647), .B(n39646), .Z(n39648) );
  NAND U40520 ( .A(n39649), .B(n39648), .Z(n39657) );
  NAND U40521 ( .A(n39651), .B(n39650), .Z(n39655) );
  NAND U40522 ( .A(n39653), .B(n39652), .Z(n39654) );
  NAND U40523 ( .A(n39655), .B(n39654), .Z(n39658) );
  XOR U40524 ( .A(n39657), .B(n39658), .Z(n39656) );
  XNOR U40525 ( .A(n39659), .B(n39656), .Z(N870) );
  NAND U40526 ( .A(n39661), .B(n39660), .Z(n39665) );
  NAND U40527 ( .A(n39663), .B(n39662), .Z(n39664) );
  NAND U40528 ( .A(n39665), .B(n39664), .Z(n39707) );
  XNOR U40529 ( .A(n39706), .B(n39707), .Z(n39709) );
  AND U40530 ( .A(x[483]), .B(y[8100]), .Z(n39744) );
  NAND U40531 ( .A(n39733), .B(n39744), .Z(n39669) );
  NAND U40532 ( .A(n39667), .B(n39666), .Z(n39668) );
  NAND U40533 ( .A(n39669), .B(n39668), .Z(n39712) );
  XOR U40534 ( .A(n39712), .B(n39713), .Z(n39715) );
  AND U40535 ( .A(x[485]), .B(y[8101]), .Z(n39902) );
  NAND U40536 ( .A(n40246), .B(n39902), .Z(n39675) );
  NAND U40537 ( .A(n39673), .B(n39672), .Z(n39674) );
  NAND U40538 ( .A(n39675), .B(n39674), .Z(n39683) );
  AND U40539 ( .A(n39676), .B(o[421]), .Z(n39689) );
  AND U40540 ( .A(y[8096]), .B(x[486]), .Z(n39678) );
  NAND U40541 ( .A(y[8102]), .B(x[480]), .Z(n39677) );
  XNOR U40542 ( .A(n39678), .B(n39677), .Z(n39690) );
  XOR U40543 ( .A(n39689), .B(n39690), .Z(n39682) );
  XOR U40544 ( .A(n39683), .B(n39682), .Z(n39685) );
  NAND U40545 ( .A(y[8100]), .B(x[482]), .Z(n39679) );
  XNOR U40546 ( .A(n39680), .B(n39679), .Z(n39694) );
  AND U40547 ( .A(y[8101]), .B(x[481]), .Z(n39936) );
  NAND U40548 ( .A(y[8098]), .B(x[484]), .Z(n39681) );
  XNOR U40549 ( .A(n39936), .B(n39681), .Z(n39698) );
  AND U40550 ( .A(x[485]), .B(y[8097]), .Z(n39703) );
  XOR U40551 ( .A(o[422]), .B(n39703), .Z(n39697) );
  XOR U40552 ( .A(n39698), .B(n39697), .Z(n39693) );
  XOR U40553 ( .A(n39694), .B(n39693), .Z(n39684) );
  XOR U40554 ( .A(n39685), .B(n39684), .Z(n39714) );
  XNOR U40555 ( .A(n39715), .B(n39714), .Z(n39708) );
  XNOR U40556 ( .A(n39709), .B(n39708), .Z(N871) );
  NAND U40557 ( .A(n39683), .B(n39682), .Z(n39687) );
  NAND U40558 ( .A(n39685), .B(n39684), .Z(n39686) );
  AND U40559 ( .A(n39687), .B(n39686), .Z(n39720) );
  AND U40560 ( .A(y[8098]), .B(x[485]), .Z(n39812) );
  NAND U40561 ( .A(y[8102]), .B(x[481]), .Z(n39688) );
  XNOR U40562 ( .A(n39812), .B(n39688), .Z(n39735) );
  AND U40563 ( .A(x[486]), .B(y[8097]), .Z(n39738) );
  XOR U40564 ( .A(o[423]), .B(n39738), .Z(n39734) );
  XOR U40565 ( .A(n39735), .B(n39734), .Z(n39754) );
  AND U40566 ( .A(x[486]), .B(y[8102]), .Z(n39956) );
  NAND U40567 ( .A(n40246), .B(n39956), .Z(n39692) );
  NAND U40568 ( .A(n39690), .B(n39689), .Z(n39691) );
  AND U40569 ( .A(n39692), .B(n39691), .Z(n39753) );
  NANDN U40570 ( .A(n39742), .B(n39744), .Z(n39696) );
  NAND U40571 ( .A(n39694), .B(n39693), .Z(n39695) );
  AND U40572 ( .A(n39696), .B(n39695), .Z(n39755) );
  XOR U40573 ( .A(n39756), .B(n39755), .Z(n39718) );
  AND U40574 ( .A(x[484]), .B(y[8101]), .Z(n40251) );
  NAND U40575 ( .A(n40251), .B(n39733), .Z(n39700) );
  NAND U40576 ( .A(n39698), .B(n39697), .Z(n39699) );
  AND U40577 ( .A(n39700), .B(n39699), .Z(n39730) );
  AND U40578 ( .A(y[8101]), .B(x[482]), .Z(n39702) );
  NAND U40579 ( .A(y[8099]), .B(x[484]), .Z(n39701) );
  XNOR U40580 ( .A(n39702), .B(n39701), .Z(n39743) );
  XNOR U40581 ( .A(n39744), .B(n39743), .Z(n39728) );
  AND U40582 ( .A(o[422]), .B(n39703), .Z(n39748) );
  AND U40583 ( .A(y[8096]), .B(x[487]), .Z(n39705) );
  NAND U40584 ( .A(y[8103]), .B(x[480]), .Z(n39704) );
  XNOR U40585 ( .A(n39705), .B(n39704), .Z(n39747) );
  XNOR U40586 ( .A(n39748), .B(n39747), .Z(n39727) );
  XOR U40587 ( .A(n39728), .B(n39727), .Z(n39729) );
  XOR U40588 ( .A(n39730), .B(n39729), .Z(n39717) );
  XOR U40589 ( .A(n39718), .B(n39717), .Z(n39719) );
  XNOR U40590 ( .A(n39720), .B(n39719), .Z(n39726) );
  NANDN U40591 ( .A(n39707), .B(n39706), .Z(n39711) );
  NAND U40592 ( .A(n39709), .B(n39708), .Z(n39710) );
  NAND U40593 ( .A(n39711), .B(n39710), .Z(n39724) );
  IV U40594 ( .A(n39725), .Z(n39723) );
  XOR U40595 ( .A(n39724), .B(n39723), .Z(n39716) );
  XNOR U40596 ( .A(n39726), .B(n39716), .Z(N872) );
  NAND U40597 ( .A(n39718), .B(n39717), .Z(n39722) );
  NAND U40598 ( .A(n39720), .B(n39719), .Z(n39721) );
  AND U40599 ( .A(n39722), .B(n39721), .Z(n39797) );
  NAND U40600 ( .A(n39728), .B(n39727), .Z(n39732) );
  NAND U40601 ( .A(n39730), .B(n39729), .Z(n39731) );
  AND U40602 ( .A(n39732), .B(n39731), .Z(n39793) );
  AND U40603 ( .A(x[485]), .B(y[8102]), .Z(n39894) );
  NAND U40604 ( .A(n39894), .B(n39733), .Z(n39737) );
  NAND U40605 ( .A(n39735), .B(n39734), .Z(n39736) );
  NAND U40606 ( .A(n39737), .B(n39736), .Z(n39791) );
  AND U40607 ( .A(o[423]), .B(n39738), .Z(n39781) );
  AND U40608 ( .A(y[8099]), .B(x[485]), .Z(n40342) );
  NAND U40609 ( .A(y[8103]), .B(x[481]), .Z(n39739) );
  XNOR U40610 ( .A(n40342), .B(n39739), .Z(n39780) );
  XOR U40611 ( .A(n39781), .B(n39780), .Z(n39766) );
  NAND U40612 ( .A(x[483]), .B(y[8101]), .Z(n40564) );
  AND U40613 ( .A(y[8098]), .B(x[486]), .Z(n39741) );
  NAND U40614 ( .A(y[8102]), .B(x[482]), .Z(n39740) );
  XNOR U40615 ( .A(n39741), .B(n39740), .Z(n39761) );
  XNOR U40616 ( .A(n40432), .B(n39761), .Z(n39764) );
  XOR U40617 ( .A(n40564), .B(n39764), .Z(n39765) );
  XOR U40618 ( .A(n39766), .B(n39765), .Z(n39790) );
  XOR U40619 ( .A(n39791), .B(n39790), .Z(n39792) );
  XOR U40620 ( .A(n39793), .B(n39792), .Z(n39802) );
  NANDN U40621 ( .A(n39742), .B(n40251), .Z(n39746) );
  NAND U40622 ( .A(n39744), .B(n39743), .Z(n39745) );
  NAND U40623 ( .A(n39746), .B(n39745), .Z(n39787) );
  AND U40624 ( .A(x[487]), .B(y[8103]), .Z(n40125) );
  NAND U40625 ( .A(n40246), .B(n40125), .Z(n39750) );
  NAND U40626 ( .A(n39748), .B(n39747), .Z(n39749) );
  NAND U40627 ( .A(n39750), .B(n39749), .Z(n39785) );
  AND U40628 ( .A(y[8096]), .B(x[488]), .Z(n39752) );
  NAND U40629 ( .A(y[8104]), .B(x[480]), .Z(n39751) );
  XNOR U40630 ( .A(n39752), .B(n39751), .Z(n39771) );
  AND U40631 ( .A(x[487]), .B(y[8097]), .Z(n39774) );
  XOR U40632 ( .A(o[424]), .B(n39774), .Z(n39770) );
  XOR U40633 ( .A(n39771), .B(n39770), .Z(n39784) );
  XOR U40634 ( .A(n39785), .B(n39784), .Z(n39786) );
  XOR U40635 ( .A(n39787), .B(n39786), .Z(n39800) );
  NANDN U40636 ( .A(n39754), .B(n39753), .Z(n39758) );
  NAND U40637 ( .A(n39756), .B(n39755), .Z(n39757) );
  NAND U40638 ( .A(n39758), .B(n39757), .Z(n39799) );
  XNOR U40639 ( .A(n39796), .B(n39798), .Z(n39759) );
  XOR U40640 ( .A(n39797), .B(n39759), .Z(N873) );
  NAND U40641 ( .A(n39956), .B(n39760), .Z(n39763) );
  NAND U40642 ( .A(n40432), .B(n39761), .Z(n39762) );
  NAND U40643 ( .A(n39763), .B(n39762), .Z(n39807) );
  NAND U40644 ( .A(n40564), .B(n39764), .Z(n39768) );
  NANDN U40645 ( .A(n39766), .B(n39765), .Z(n39767) );
  AND U40646 ( .A(n39768), .B(n39767), .Z(n39806) );
  XOR U40647 ( .A(n39807), .B(n39806), .Z(n39809) );
  AND U40648 ( .A(x[488]), .B(y[8104]), .Z(n39769) );
  NAND U40649 ( .A(n39769), .B(n40246), .Z(n39773) );
  NAND U40650 ( .A(n39771), .B(n39770), .Z(n39772) );
  AND U40651 ( .A(n39773), .B(n39772), .Z(n39841) );
  AND U40652 ( .A(o[424]), .B(n39774), .Z(n39814) );
  AND U40653 ( .A(y[8100]), .B(x[485]), .Z(n39776) );
  NAND U40654 ( .A(y[8098]), .B(x[487]), .Z(n39775) );
  XNOR U40655 ( .A(n39776), .B(n39775), .Z(n39813) );
  XNOR U40656 ( .A(n39814), .B(n39813), .Z(n39839) );
  AND U40657 ( .A(y[8096]), .B(x[489]), .Z(n39778) );
  NAND U40658 ( .A(y[8105]), .B(x[480]), .Z(n39777) );
  XNOR U40659 ( .A(n39778), .B(n39777), .Z(n39821) );
  AND U40660 ( .A(x[488]), .B(y[8097]), .Z(n39830) );
  XOR U40661 ( .A(o[425]), .B(n39830), .Z(n39820) );
  XNOR U40662 ( .A(n39821), .B(n39820), .Z(n39838) );
  XOR U40663 ( .A(n39839), .B(n39838), .Z(n39840) );
  XNOR U40664 ( .A(n39841), .B(n39840), .Z(n39835) );
  AND U40665 ( .A(y[8099]), .B(x[486]), .Z(n40194) );
  NAND U40666 ( .A(y[8104]), .B(x[481]), .Z(n39779) );
  XNOR U40667 ( .A(n40194), .B(n39779), .Z(n39825) );
  XNOR U40668 ( .A(n40251), .B(n39825), .Z(n39845) );
  AND U40669 ( .A(x[482]), .B(y[8103]), .Z(n40475) );
  NAND U40670 ( .A(x[483]), .B(y[8102]), .Z(n40204) );
  XNOR U40671 ( .A(n40475), .B(n40204), .Z(n39844) );
  XNOR U40672 ( .A(n39845), .B(n39844), .Z(n39833) );
  NAND U40673 ( .A(x[485]), .B(y[8103]), .Z(n40030) );
  AND U40674 ( .A(x[481]), .B(y[8099]), .Z(n39824) );
  NANDN U40675 ( .A(n40030), .B(n39824), .Z(n39783) );
  NAND U40676 ( .A(n39781), .B(n39780), .Z(n39782) );
  NAND U40677 ( .A(n39783), .B(n39782), .Z(n39832) );
  XOR U40678 ( .A(n39833), .B(n39832), .Z(n39834) );
  XOR U40679 ( .A(n39835), .B(n39834), .Z(n39808) );
  XOR U40680 ( .A(n39809), .B(n39808), .Z(n39856) );
  NAND U40681 ( .A(n39785), .B(n39784), .Z(n39789) );
  NAND U40682 ( .A(n39787), .B(n39786), .Z(n39788) );
  NAND U40683 ( .A(n39789), .B(n39788), .Z(n39854) );
  NAND U40684 ( .A(n39791), .B(n39790), .Z(n39795) );
  NAND U40685 ( .A(n39793), .B(n39792), .Z(n39794) );
  NAND U40686 ( .A(n39795), .B(n39794), .Z(n39853) );
  XOR U40687 ( .A(n39854), .B(n39853), .Z(n39855) );
  XNOR U40688 ( .A(n39856), .B(n39855), .Z(n39849) );
  NANDN U40689 ( .A(n39800), .B(n39799), .Z(n39804) );
  NANDN U40690 ( .A(n39802), .B(n39801), .Z(n39803) );
  AND U40691 ( .A(n39804), .B(n39803), .Z(n39847) );
  IV U40692 ( .A(n39847), .Z(n39846) );
  XOR U40693 ( .A(n39848), .B(n39846), .Z(n39805) );
  XNOR U40694 ( .A(n39849), .B(n39805), .Z(N874) );
  NAND U40695 ( .A(n39807), .B(n39806), .Z(n39811) );
  NAND U40696 ( .A(n39809), .B(n39808), .Z(n39810) );
  AND U40697 ( .A(n39811), .B(n39810), .Z(n39922) );
  AND U40698 ( .A(x[487]), .B(y[8100]), .Z(n39896) );
  NAND U40699 ( .A(n39896), .B(n39812), .Z(n39816) );
  NAND U40700 ( .A(n39814), .B(n39813), .Z(n39815) );
  AND U40701 ( .A(n39816), .B(n39815), .Z(n39909) );
  AND U40702 ( .A(y[8099]), .B(x[487]), .Z(n39818) );
  NAND U40703 ( .A(y[8102]), .B(x[484]), .Z(n39817) );
  XNOR U40704 ( .A(n39818), .B(n39817), .Z(n39880) );
  AND U40705 ( .A(x[486]), .B(y[8100]), .Z(n39879) );
  XNOR U40706 ( .A(n39880), .B(n39879), .Z(n39907) );
  AND U40707 ( .A(x[488]), .B(y[8098]), .Z(n40099) );
  AND U40708 ( .A(x[489]), .B(y[8097]), .Z(n39890) );
  XOR U40709 ( .A(o[426]), .B(n39890), .Z(n39901) );
  XOR U40710 ( .A(n40099), .B(n39901), .Z(n39903) );
  XNOR U40711 ( .A(n39903), .B(n39902), .Z(n39906) );
  XOR U40712 ( .A(n39907), .B(n39906), .Z(n39908) );
  XNOR U40713 ( .A(n39909), .B(n39908), .Z(n39869) );
  AND U40714 ( .A(x[489]), .B(y[8105]), .Z(n39819) );
  NAND U40715 ( .A(n39819), .B(n40246), .Z(n39823) );
  NAND U40716 ( .A(n39821), .B(n39820), .Z(n39822) );
  NAND U40717 ( .A(n39823), .B(n39822), .Z(n39867) );
  AND U40718 ( .A(x[486]), .B(y[8104]), .Z(n40135) );
  NAND U40719 ( .A(n40135), .B(n39824), .Z(n39827) );
  NAND U40720 ( .A(n40251), .B(n39825), .Z(n39826) );
  NAND U40721 ( .A(n39827), .B(n39826), .Z(n39875) );
  AND U40722 ( .A(y[8096]), .B(x[490]), .Z(n39829) );
  NAND U40723 ( .A(y[8106]), .B(x[480]), .Z(n39828) );
  XNOR U40724 ( .A(n39829), .B(n39828), .Z(n39885) );
  AND U40725 ( .A(o[425]), .B(n39830), .Z(n39884) );
  XOR U40726 ( .A(n39885), .B(n39884), .Z(n39873) );
  AND U40727 ( .A(y[8103]), .B(x[483]), .Z(n40801) );
  NAND U40728 ( .A(y[8105]), .B(x[481]), .Z(n39831) );
  XNOR U40729 ( .A(n40801), .B(n39831), .Z(n39897) );
  AND U40730 ( .A(x[482]), .B(y[8104]), .Z(n39898) );
  XOR U40731 ( .A(n39897), .B(n39898), .Z(n39872) );
  XOR U40732 ( .A(n39873), .B(n39872), .Z(n39874) );
  XOR U40733 ( .A(n39875), .B(n39874), .Z(n39866) );
  XOR U40734 ( .A(n39867), .B(n39866), .Z(n39868) );
  XNOR U40735 ( .A(n39869), .B(n39868), .Z(n39920) );
  NAND U40736 ( .A(n39833), .B(n39832), .Z(n39837) );
  NAND U40737 ( .A(n39835), .B(n39834), .Z(n39836) );
  AND U40738 ( .A(n39837), .B(n39836), .Z(n39863) );
  NAND U40739 ( .A(n39839), .B(n39838), .Z(n39843) );
  NAND U40740 ( .A(n39841), .B(n39840), .Z(n39842) );
  AND U40741 ( .A(n39843), .B(n39842), .Z(n39860) );
  XOR U40742 ( .A(n39860), .B(n39861), .Z(n39862) );
  XOR U40743 ( .A(n39863), .B(n39862), .Z(n39919) );
  XOR U40744 ( .A(n39920), .B(n39919), .Z(n39921) );
  XNOR U40745 ( .A(n39922), .B(n39921), .Z(n39915) );
  OR U40746 ( .A(n39848), .B(n39846), .Z(n39852) );
  ANDN U40747 ( .B(n39848), .A(n39847), .Z(n39850) );
  OR U40748 ( .A(n39850), .B(n39849), .Z(n39851) );
  AND U40749 ( .A(n39852), .B(n39851), .Z(n39913) );
  NAND U40750 ( .A(n39854), .B(n39853), .Z(n39858) );
  NAND U40751 ( .A(n39856), .B(n39855), .Z(n39857) );
  AND U40752 ( .A(n39858), .B(n39857), .Z(n39914) );
  IV U40753 ( .A(n39914), .Z(n39912) );
  XOR U40754 ( .A(n39913), .B(n39912), .Z(n39859) );
  XNOR U40755 ( .A(n39915), .B(n39859), .Z(N875) );
  NAND U40756 ( .A(n39861), .B(n39860), .Z(n39865) );
  NANDN U40757 ( .A(n39863), .B(n39862), .Z(n39864) );
  AND U40758 ( .A(n39865), .B(n39864), .Z(n39985) );
  NAND U40759 ( .A(n39867), .B(n39866), .Z(n39871) );
  NAND U40760 ( .A(n39869), .B(n39868), .Z(n39870) );
  NAND U40761 ( .A(n39871), .B(n39870), .Z(n39983) );
  NAND U40762 ( .A(n39873), .B(n39872), .Z(n39877) );
  NAND U40763 ( .A(n39875), .B(n39874), .Z(n39876) );
  NAND U40764 ( .A(n39877), .B(n39876), .Z(n39976) );
  AND U40765 ( .A(x[487]), .B(y[8102]), .Z(n40025) );
  AND U40766 ( .A(x[484]), .B(y[8099]), .Z(n39878) );
  NAND U40767 ( .A(n40025), .B(n39878), .Z(n39882) );
  NAND U40768 ( .A(n39880), .B(n39879), .Z(n39881) );
  NAND U40769 ( .A(n39882), .B(n39881), .Z(n39974) );
  AND U40770 ( .A(x[490]), .B(y[8106]), .Z(n39883) );
  NAND U40771 ( .A(n39883), .B(n40246), .Z(n39887) );
  NAND U40772 ( .A(n39885), .B(n39884), .Z(n39886) );
  NAND U40773 ( .A(n39887), .B(n39886), .Z(n39970) );
  AND U40774 ( .A(y[8096]), .B(x[491]), .Z(n39889) );
  NAND U40775 ( .A(y[8107]), .B(x[480]), .Z(n39888) );
  XNOR U40776 ( .A(n39889), .B(n39888), .Z(n39947) );
  AND U40777 ( .A(o[426]), .B(n39890), .Z(n39946) );
  XOR U40778 ( .A(n39947), .B(n39946), .Z(n39968) );
  AND U40779 ( .A(y[8101]), .B(x[486]), .Z(n39892) );
  NAND U40780 ( .A(y[8106]), .B(x[481]), .Z(n39891) );
  XNOR U40781 ( .A(n39892), .B(n39891), .Z(n39938) );
  AND U40782 ( .A(x[490]), .B(y[8097]), .Z(n39957) );
  XOR U40783 ( .A(o[427]), .B(n39957), .Z(n39937) );
  XOR U40784 ( .A(n39938), .B(n39937), .Z(n39967) );
  XOR U40785 ( .A(n39968), .B(n39967), .Z(n39969) );
  XOR U40786 ( .A(n39970), .B(n39969), .Z(n39973) );
  XOR U40787 ( .A(n39974), .B(n39973), .Z(n39975) );
  XNOR U40788 ( .A(n39976), .B(n39975), .Z(n39960) );
  NAND U40789 ( .A(x[483]), .B(y[8104]), .Z(n40930) );
  NAND U40790 ( .A(y[8105]), .B(x[482]), .Z(n39893) );
  XNOR U40791 ( .A(n39894), .B(n39893), .Z(n39933) );
  AND U40792 ( .A(x[484]), .B(y[8103]), .Z(n39932) );
  XNOR U40793 ( .A(n39933), .B(n39932), .Z(n39964) );
  XOR U40794 ( .A(n40930), .B(n39964), .Z(n39966) );
  NAND U40795 ( .A(y[8098]), .B(x[489]), .Z(n39895) );
  XNOR U40796 ( .A(n39896), .B(n39895), .Z(n39952) );
  AND U40797 ( .A(x[488]), .B(y[8099]), .Z(n39951) );
  XNOR U40798 ( .A(n39952), .B(n39951), .Z(n39965) );
  XNOR U40799 ( .A(n39966), .B(n39965), .Z(n39929) );
  NAND U40800 ( .A(x[483]), .B(y[8105]), .Z(n40021) );
  AND U40801 ( .A(x[481]), .B(y[8103]), .Z(n40241) );
  NANDN U40802 ( .A(n40021), .B(n40241), .Z(n39900) );
  NAND U40803 ( .A(n39898), .B(n39897), .Z(n39899) );
  NAND U40804 ( .A(n39900), .B(n39899), .Z(n39927) );
  NAND U40805 ( .A(n40099), .B(n39901), .Z(n39905) );
  NAND U40806 ( .A(n39903), .B(n39902), .Z(n39904) );
  NAND U40807 ( .A(n39905), .B(n39904), .Z(n39926) );
  XOR U40808 ( .A(n39927), .B(n39926), .Z(n39928) );
  XNOR U40809 ( .A(n39929), .B(n39928), .Z(n39959) );
  NAND U40810 ( .A(n39907), .B(n39906), .Z(n39911) );
  NAND U40811 ( .A(n39909), .B(n39908), .Z(n39910) );
  NAND U40812 ( .A(n39911), .B(n39910), .Z(n39958) );
  XOR U40813 ( .A(n39959), .B(n39958), .Z(n39961) );
  XNOR U40814 ( .A(n39960), .B(n39961), .Z(n39982) );
  XOR U40815 ( .A(n39983), .B(n39982), .Z(n39984) );
  XOR U40816 ( .A(n39985), .B(n39984), .Z(n39981) );
  NANDN U40817 ( .A(n39912), .B(n39913), .Z(n39918) );
  NOR U40818 ( .A(n39914), .B(n39913), .Z(n39916) );
  OR U40819 ( .A(n39916), .B(n39915), .Z(n39917) );
  AND U40820 ( .A(n39918), .B(n39917), .Z(n39979) );
  NAND U40821 ( .A(n39920), .B(n39919), .Z(n39924) );
  NAND U40822 ( .A(n39922), .B(n39921), .Z(n39923) );
  AND U40823 ( .A(n39924), .B(n39923), .Z(n39980) );
  XOR U40824 ( .A(n39979), .B(n39980), .Z(n39925) );
  XNOR U40825 ( .A(n39981), .B(n39925), .Z(N876) );
  NAND U40826 ( .A(n39927), .B(n39926), .Z(n39931) );
  NAND U40827 ( .A(n39929), .B(n39928), .Z(n39930) );
  NAND U40828 ( .A(n39931), .B(n39930), .Z(n40062) );
  AND U40829 ( .A(x[482]), .B(y[8102]), .Z(n40658) );
  AND U40830 ( .A(x[485]), .B(y[8105]), .Z(n40466) );
  NAND U40831 ( .A(n40658), .B(n40466), .Z(n39935) );
  NAND U40832 ( .A(n39933), .B(n39932), .Z(n39934) );
  NAND U40833 ( .A(n39935), .B(n39934), .Z(n40009) );
  AND U40834 ( .A(x[486]), .B(y[8106]), .Z(n40258) );
  NAND U40835 ( .A(n40258), .B(n39936), .Z(n39940) );
  NAND U40836 ( .A(n39938), .B(n39937), .Z(n39939) );
  NAND U40837 ( .A(n39940), .B(n39939), .Z(n40008) );
  XOR U40838 ( .A(n40009), .B(n40008), .Z(n40010) );
  AND U40839 ( .A(x[489]), .B(y[8099]), .Z(n40653) );
  AND U40840 ( .A(x[490]), .B(y[8098]), .Z(n40696) );
  AND U40841 ( .A(y[8104]), .B(x[484]), .Z(n39941) );
  XOR U40842 ( .A(n40696), .B(n39941), .Z(n40052) );
  XOR U40843 ( .A(n40653), .B(n40052), .Z(n40031) );
  NAND U40844 ( .A(x[487]), .B(y[8101]), .Z(n40029) );
  XOR U40845 ( .A(n40030), .B(n40029), .Z(n40032) );
  AND U40846 ( .A(y[8096]), .B(x[492]), .Z(n39943) );
  NAND U40847 ( .A(y[8108]), .B(x[480]), .Z(n39942) );
  XNOR U40848 ( .A(n39943), .B(n39942), .Z(n40046) );
  AND U40849 ( .A(x[491]), .B(y[8097]), .Z(n40026) );
  XOR U40850 ( .A(o[428]), .B(n40026), .Z(n40045) );
  XOR U40851 ( .A(n40046), .B(n40045), .Z(n40015) );
  AND U40852 ( .A(y[8106]), .B(x[482]), .Z(n39945) );
  NAND U40853 ( .A(y[8100]), .B(x[488]), .Z(n39944) );
  XNOR U40854 ( .A(n39945), .B(n39944), .Z(n40020) );
  XOR U40855 ( .A(n40015), .B(n40014), .Z(n40016) );
  XNOR U40856 ( .A(n40010), .B(n40011), .Z(n40060) );
  AND U40857 ( .A(x[491]), .B(y[8107]), .Z(n41066) );
  NAND U40858 ( .A(n41066), .B(n40246), .Z(n39949) );
  NAND U40859 ( .A(n39947), .B(n39946), .Z(n39948) );
  NAND U40860 ( .A(n39949), .B(n39948), .Z(n40037) );
  AND U40861 ( .A(x[487]), .B(y[8098]), .Z(n40180) );
  AND U40862 ( .A(x[489]), .B(y[8100]), .Z(n39950) );
  NAND U40863 ( .A(n40180), .B(n39950), .Z(n39954) );
  NAND U40864 ( .A(n39952), .B(n39951), .Z(n39953) );
  NAND U40865 ( .A(n39954), .B(n39953), .Z(n40035) );
  NAND U40866 ( .A(y[8107]), .B(x[481]), .Z(n39955) );
  XNOR U40867 ( .A(n39956), .B(n39955), .Z(n40042) );
  AND U40868 ( .A(o[427]), .B(n39957), .Z(n40041) );
  XOR U40869 ( .A(n40042), .B(n40041), .Z(n40036) );
  XOR U40870 ( .A(n40035), .B(n40036), .Z(n40038) );
  XOR U40871 ( .A(n40037), .B(n40038), .Z(n40059) );
  XOR U40872 ( .A(n40060), .B(n40059), .Z(n40061) );
  XNOR U40873 ( .A(n40062), .B(n40061), .Z(n39990) );
  NAND U40874 ( .A(n39959), .B(n39958), .Z(n39963) );
  NAND U40875 ( .A(n39961), .B(n39960), .Z(n39962) );
  NAND U40876 ( .A(n39963), .B(n39962), .Z(n39989) );
  XOR U40877 ( .A(n39990), .B(n39989), .Z(n39992) );
  NAND U40878 ( .A(n39968), .B(n39967), .Z(n39972) );
  NAND U40879 ( .A(n39970), .B(n39969), .Z(n39971) );
  AND U40880 ( .A(n39972), .B(n39971), .Z(n40002) );
  XOR U40881 ( .A(n40003), .B(n40002), .Z(n40004) );
  NAND U40882 ( .A(n39974), .B(n39973), .Z(n39978) );
  NAND U40883 ( .A(n39976), .B(n39975), .Z(n39977) );
  AND U40884 ( .A(n39978), .B(n39977), .Z(n40005) );
  XOR U40885 ( .A(n40004), .B(n40005), .Z(n39991) );
  XNOR U40886 ( .A(n39992), .B(n39991), .Z(n39998) );
  NAND U40887 ( .A(n39983), .B(n39982), .Z(n39987) );
  NANDN U40888 ( .A(n39985), .B(n39984), .Z(n39986) );
  AND U40889 ( .A(n39987), .B(n39986), .Z(n39997) );
  IV U40890 ( .A(n39997), .Z(n39995) );
  XOR U40891 ( .A(n39996), .B(n39995), .Z(n39988) );
  XNOR U40892 ( .A(n39998), .B(n39988), .Z(N877) );
  NAND U40893 ( .A(n39990), .B(n39989), .Z(n39994) );
  NAND U40894 ( .A(n39992), .B(n39991), .Z(n39993) );
  AND U40895 ( .A(n39994), .B(n39993), .Z(n40073) );
  NANDN U40896 ( .A(n39995), .B(n39996), .Z(n40001) );
  NOR U40897 ( .A(n39997), .B(n39996), .Z(n39999) );
  OR U40898 ( .A(n39999), .B(n39998), .Z(n40000) );
  AND U40899 ( .A(n40001), .B(n40000), .Z(n40072) );
  NAND U40900 ( .A(n40003), .B(n40002), .Z(n40007) );
  NAND U40901 ( .A(n40005), .B(n40004), .Z(n40006) );
  NAND U40902 ( .A(n40007), .B(n40006), .Z(n40069) );
  NAND U40903 ( .A(n40009), .B(n40008), .Z(n40013) );
  NANDN U40904 ( .A(n40011), .B(n40010), .Z(n40012) );
  NAND U40905 ( .A(n40013), .B(n40012), .Z(n40075) );
  NAND U40906 ( .A(n40015), .B(n40014), .Z(n40019) );
  NANDN U40907 ( .A(n40017), .B(n40016), .Z(n40018) );
  NAND U40908 ( .A(n40019), .B(n40018), .Z(n40083) );
  AND U40909 ( .A(y[8106]), .B(x[488]), .Z(n41302) );
  AND U40910 ( .A(x[482]), .B(y[8100]), .Z(n40190) );
  NAND U40911 ( .A(n41302), .B(n40190), .Z(n40023) );
  NANDN U40912 ( .A(n40021), .B(n40020), .Z(n40022) );
  NAND U40913 ( .A(n40023), .B(n40022), .Z(n40114) );
  NAND U40914 ( .A(y[8108]), .B(x[481]), .Z(n40024) );
  XNOR U40915 ( .A(n40025), .B(n40024), .Z(n40105) );
  AND U40916 ( .A(o[428]), .B(n40026), .Z(n40104) );
  XOR U40917 ( .A(n40105), .B(n40104), .Z(n40112) );
  AND U40918 ( .A(x[486]), .B(y[8103]), .Z(n41106) );
  AND U40919 ( .A(y[8107]), .B(x[482]), .Z(n40028) );
  NAND U40920 ( .A(y[8100]), .B(x[489]), .Z(n40027) );
  XNOR U40921 ( .A(n40028), .B(n40027), .Z(n40118) );
  XOR U40922 ( .A(n41106), .B(n40118), .Z(n40111) );
  XOR U40923 ( .A(n40112), .B(n40111), .Z(n40113) );
  XOR U40924 ( .A(n40114), .B(n40113), .Z(n40082) );
  NAND U40925 ( .A(n40030), .B(n40029), .Z(n40034) );
  ANDN U40926 ( .B(n40032), .A(n40031), .Z(n40033) );
  ANDN U40927 ( .B(n40034), .A(n40033), .Z(n40081) );
  XOR U40928 ( .A(n40082), .B(n40081), .Z(n40084) );
  XOR U40929 ( .A(n40083), .B(n40084), .Z(n40076) );
  XOR U40930 ( .A(n40075), .B(n40076), .Z(n40078) );
  NAND U40931 ( .A(n40036), .B(n40035), .Z(n40040) );
  NAND U40932 ( .A(n40038), .B(n40037), .Z(n40039) );
  NAND U40933 ( .A(n40040), .B(n40039), .Z(n40089) );
  AND U40934 ( .A(x[486]), .B(y[8107]), .Z(n40397) );
  IV U40935 ( .A(n40397), .Z(n40468) );
  AND U40936 ( .A(x[481]), .B(y[8102]), .Z(n40103) );
  NANDN U40937 ( .A(n40468), .B(n40103), .Z(n40044) );
  NAND U40938 ( .A(n40042), .B(n40041), .Z(n40043) );
  NAND U40939 ( .A(n40044), .B(n40043), .Z(n40096) );
  AND U40940 ( .A(x[492]), .B(y[8108]), .Z(n41308) );
  NAND U40941 ( .A(n41308), .B(n40246), .Z(n40048) );
  NAND U40942 ( .A(n40046), .B(n40045), .Z(n40047) );
  NAND U40943 ( .A(n40048), .B(n40047), .Z(n40094) );
  AND U40944 ( .A(x[490]), .B(y[8099]), .Z(n40942) );
  AND U40945 ( .A(y[8098]), .B(x[491]), .Z(n40903) );
  NAND U40946 ( .A(y[8101]), .B(x[488]), .Z(n40049) );
  XNOR U40947 ( .A(n40903), .B(n40049), .Z(n40100) );
  XOR U40948 ( .A(n40942), .B(n40100), .Z(n40093) );
  XOR U40949 ( .A(n40094), .B(n40093), .Z(n40095) );
  XOR U40950 ( .A(n40096), .B(n40095), .Z(n40087) );
  AND U40951 ( .A(x[490]), .B(y[8104]), .Z(n40051) );
  AND U40952 ( .A(x[484]), .B(y[8098]), .Z(n40050) );
  NAND U40953 ( .A(n40051), .B(n40050), .Z(n40054) );
  NAND U40954 ( .A(n40653), .B(n40052), .Z(n40053) );
  NAND U40955 ( .A(n40054), .B(n40053), .Z(n40138) );
  AND U40956 ( .A(y[8096]), .B(x[493]), .Z(n40056) );
  NAND U40957 ( .A(y[8109]), .B(x[480]), .Z(n40055) );
  XNOR U40958 ( .A(n40056), .B(n40055), .Z(n40131) );
  AND U40959 ( .A(x[492]), .B(y[8097]), .Z(n40123) );
  XOR U40960 ( .A(o[429]), .B(n40123), .Z(n40130) );
  XOR U40961 ( .A(n40131), .B(n40130), .Z(n40137) );
  AND U40962 ( .A(y[8104]), .B(x[485]), .Z(n40058) );
  NAND U40963 ( .A(y[8106]), .B(x[483]), .Z(n40057) );
  XNOR U40964 ( .A(n40058), .B(n40057), .Z(n40126) );
  AND U40965 ( .A(x[484]), .B(y[8105]), .Z(n40127) );
  XOR U40966 ( .A(n40126), .B(n40127), .Z(n40136) );
  XOR U40967 ( .A(n40137), .B(n40136), .Z(n40139) );
  XNOR U40968 ( .A(n40138), .B(n40139), .Z(n40088) );
  XOR U40969 ( .A(n40089), .B(n40090), .Z(n40077) );
  XNOR U40970 ( .A(n40078), .B(n40077), .Z(n40067) );
  NAND U40971 ( .A(n40060), .B(n40059), .Z(n40064) );
  NAND U40972 ( .A(n40062), .B(n40061), .Z(n40063) );
  AND U40973 ( .A(n40064), .B(n40063), .Z(n40066) );
  XOR U40974 ( .A(n40067), .B(n40066), .Z(n40068) );
  XOR U40975 ( .A(n40069), .B(n40068), .Z(n40074) );
  XNOR U40976 ( .A(n40072), .B(n40074), .Z(n40065) );
  XOR U40977 ( .A(n40073), .B(n40065), .Z(N878) );
  NAND U40978 ( .A(n40067), .B(n40066), .Z(n40071) );
  NAND U40979 ( .A(n40069), .B(n40068), .Z(n40070) );
  NAND U40980 ( .A(n40071), .B(n40070), .Z(n40151) );
  IV U40981 ( .A(n40151), .Z(n40149) );
  NAND U40982 ( .A(n40076), .B(n40075), .Z(n40080) );
  NAND U40983 ( .A(n40078), .B(n40077), .Z(n40079) );
  NAND U40984 ( .A(n40080), .B(n40079), .Z(n40144) );
  NAND U40985 ( .A(n40082), .B(n40081), .Z(n40086) );
  NAND U40986 ( .A(n40084), .B(n40083), .Z(n40085) );
  NAND U40987 ( .A(n40086), .B(n40085), .Z(n40143) );
  XOR U40988 ( .A(n40144), .B(n40143), .Z(n40145) );
  NANDN U40989 ( .A(n40088), .B(n40087), .Z(n40092) );
  NAND U40990 ( .A(n40090), .B(n40089), .Z(n40091) );
  NAND U40991 ( .A(n40092), .B(n40091), .Z(n40158) );
  NAND U40992 ( .A(n40094), .B(n40093), .Z(n40098) );
  NAND U40993 ( .A(n40096), .B(n40095), .Z(n40097) );
  AND U40994 ( .A(n40098), .B(n40097), .Z(n40165) );
  AND U40995 ( .A(x[491]), .B(y[8101]), .Z(n40272) );
  NAND U40996 ( .A(n40272), .B(n40099), .Z(n40102) );
  NAND U40997 ( .A(n40100), .B(n40942), .Z(n40101) );
  NAND U40998 ( .A(n40102), .B(n40101), .Z(n40220) );
  NAND U40999 ( .A(x[487]), .B(y[8108]), .Z(n40668) );
  NANDN U41000 ( .A(n40668), .B(n40103), .Z(n40107) );
  NAND U41001 ( .A(n40105), .B(n40104), .Z(n40106) );
  NAND U41002 ( .A(n40107), .B(n40106), .Z(n40219) );
  XOR U41003 ( .A(n40220), .B(n40219), .Z(n40222) );
  AND U41004 ( .A(x[484]), .B(y[8106]), .Z(n40573) );
  AND U41005 ( .A(y[8107]), .B(x[483]), .Z(n40109) );
  NAND U41006 ( .A(y[8102]), .B(x[488]), .Z(n40108) );
  XNOR U41007 ( .A(n40109), .B(n40108), .Z(n40205) );
  XOR U41008 ( .A(n40466), .B(n40205), .Z(n40214) );
  XOR U41009 ( .A(n40573), .B(n40214), .Z(n40216) );
  AND U41010 ( .A(x[489]), .B(y[8101]), .Z(n40772) );
  AND U41011 ( .A(x[482]), .B(y[8108]), .Z(n40110) );
  AND U41012 ( .A(y[8100]), .B(x[490]), .Z(n40796) );
  XOR U41013 ( .A(n40110), .B(n40796), .Z(n40191) );
  XOR U41014 ( .A(n40772), .B(n40191), .Z(n40215) );
  XOR U41015 ( .A(n40216), .B(n40215), .Z(n40221) );
  XNOR U41016 ( .A(n40222), .B(n40221), .Z(n40163) );
  NAND U41017 ( .A(n40112), .B(n40111), .Z(n40116) );
  NAND U41018 ( .A(n40114), .B(n40113), .Z(n40115) );
  AND U41019 ( .A(n40116), .B(n40115), .Z(n40162) );
  XOR U41020 ( .A(n40163), .B(n40162), .Z(n40164) );
  XOR U41021 ( .A(n40165), .B(n40164), .Z(n40157) );
  AND U41022 ( .A(x[489]), .B(y[8107]), .Z(n40117) );
  NAND U41023 ( .A(n40117), .B(n40190), .Z(n40120) );
  NAND U41024 ( .A(n40118), .B(n41106), .Z(n40119) );
  NAND U41025 ( .A(n40120), .B(n40119), .Z(n40177) );
  AND U41026 ( .A(y[8096]), .B(x[494]), .Z(n40122) );
  NAND U41027 ( .A(y[8110]), .B(x[480]), .Z(n40121) );
  XNOR U41028 ( .A(n40122), .B(n40121), .Z(n40200) );
  AND U41029 ( .A(o[429]), .B(n40123), .Z(n40199) );
  XOR U41030 ( .A(n40200), .B(n40199), .Z(n40175) );
  NAND U41031 ( .A(y[8098]), .B(x[492]), .Z(n40124) );
  XNOR U41032 ( .A(n40125), .B(n40124), .Z(n40181) );
  NAND U41033 ( .A(x[493]), .B(y[8097]), .Z(n40189) );
  XNOR U41034 ( .A(o[430]), .B(n40189), .Z(n40182) );
  XOR U41035 ( .A(n40181), .B(n40182), .Z(n40174) );
  XOR U41036 ( .A(n40175), .B(n40174), .Z(n40176) );
  XOR U41037 ( .A(n40177), .B(n40176), .Z(n40226) );
  AND U41038 ( .A(x[485]), .B(y[8106]), .Z(n40259) );
  NANDN U41039 ( .A(n40930), .B(n40259), .Z(n40129) );
  NAND U41040 ( .A(n40127), .B(n40126), .Z(n40128) );
  AND U41041 ( .A(n40129), .B(n40128), .Z(n40171) );
  AND U41042 ( .A(x[493]), .B(y[8109]), .Z(n41680) );
  NAND U41043 ( .A(n41680), .B(n40246), .Z(n40133) );
  NAND U41044 ( .A(n40131), .B(n40130), .Z(n40132) );
  NAND U41045 ( .A(n40133), .B(n40132), .Z(n40169) );
  NAND U41046 ( .A(y[8099]), .B(x[491]), .Z(n40134) );
  XNOR U41047 ( .A(n40135), .B(n40134), .Z(n40195) );
  AND U41048 ( .A(x[481]), .B(y[8109]), .Z(n40196) );
  XOR U41049 ( .A(n40195), .B(n40196), .Z(n40168) );
  XOR U41050 ( .A(n40169), .B(n40168), .Z(n40170) );
  XOR U41051 ( .A(n40171), .B(n40170), .Z(n40225) );
  NAND U41052 ( .A(n40137), .B(n40136), .Z(n40141) );
  NAND U41053 ( .A(n40139), .B(n40138), .Z(n40140) );
  AND U41054 ( .A(n40141), .B(n40140), .Z(n40227) );
  XNOR U41055 ( .A(n40228), .B(n40227), .Z(n40156) );
  XOR U41056 ( .A(n40158), .B(n40159), .Z(n40146) );
  XNOR U41057 ( .A(n40145), .B(n40146), .Z(n40152) );
  XNOR U41058 ( .A(n40150), .B(n40152), .Z(n40142) );
  XOR U41059 ( .A(n40149), .B(n40142), .Z(N879) );
  NAND U41060 ( .A(n40144), .B(n40143), .Z(n40148) );
  NANDN U41061 ( .A(n40146), .B(n40145), .Z(n40147) );
  AND U41062 ( .A(n40148), .B(n40147), .Z(n40238) );
  NANDN U41063 ( .A(n40149), .B(n40150), .Z(n40155) );
  NOR U41064 ( .A(n40151), .B(n40150), .Z(n40153) );
  OR U41065 ( .A(n40153), .B(n40152), .Z(n40154) );
  AND U41066 ( .A(n40155), .B(n40154), .Z(n40239) );
  NANDN U41067 ( .A(n40157), .B(n40156), .Z(n40161) );
  NANDN U41068 ( .A(n40159), .B(n40158), .Z(n40160) );
  NAND U41069 ( .A(n40161), .B(n40160), .Z(n40234) );
  NAND U41070 ( .A(n40163), .B(n40162), .Z(n40167) );
  NAND U41071 ( .A(n40165), .B(n40164), .Z(n40166) );
  NAND U41072 ( .A(n40167), .B(n40166), .Z(n40302) );
  NAND U41073 ( .A(n40169), .B(n40168), .Z(n40173) );
  NANDN U41074 ( .A(n40171), .B(n40170), .Z(n40172) );
  NAND U41075 ( .A(n40173), .B(n40172), .Z(n40308) );
  NAND U41076 ( .A(n40175), .B(n40174), .Z(n40179) );
  NAND U41077 ( .A(n40177), .B(n40176), .Z(n40178) );
  NAND U41078 ( .A(n40179), .B(n40178), .Z(n40306) );
  NAND U41079 ( .A(x[492]), .B(y[8103]), .Z(n40660) );
  NANDN U41080 ( .A(n40660), .B(n40180), .Z(n40184) );
  NAND U41081 ( .A(n40182), .B(n40181), .Z(n40183) );
  AND U41082 ( .A(n40184), .B(n40183), .Z(n40282) );
  AND U41083 ( .A(y[8100]), .B(x[491]), .Z(n40186) );
  NAND U41084 ( .A(y[8098]), .B(x[493]), .Z(n40185) );
  XNOR U41085 ( .A(n40186), .B(n40185), .Z(n40286) );
  AND U41086 ( .A(x[492]), .B(y[8099]), .Z(n40285) );
  XNOR U41087 ( .A(n40286), .B(n40285), .Z(n40280) );
  AND U41088 ( .A(y[8096]), .B(x[495]), .Z(n40188) );
  NAND U41089 ( .A(y[8111]), .B(x[480]), .Z(n40187) );
  XNOR U41090 ( .A(n40188), .B(n40187), .Z(n40248) );
  ANDN U41091 ( .B(o[430]), .A(n40189), .Z(n40247) );
  XNOR U41092 ( .A(n40248), .B(n40247), .Z(n40279) );
  XOR U41093 ( .A(n40280), .B(n40279), .Z(n40281) );
  XNOR U41094 ( .A(n40282), .B(n40281), .Z(n40314) );
  NAND U41095 ( .A(x[490]), .B(y[8108]), .Z(n41108) );
  NANDN U41096 ( .A(n41108), .B(n40190), .Z(n40193) );
  NAND U41097 ( .A(n40772), .B(n40191), .Z(n40192) );
  NAND U41098 ( .A(n40193), .B(n40192), .Z(n40312) );
  AND U41099 ( .A(y[8104]), .B(x[491]), .Z(n40572) );
  NAND U41100 ( .A(n40572), .B(n40194), .Z(n40198) );
  NAND U41101 ( .A(n40196), .B(n40195), .Z(n40197) );
  NAND U41102 ( .A(n40198), .B(n40197), .Z(n40311) );
  XOR U41103 ( .A(n40312), .B(n40311), .Z(n40313) );
  XOR U41104 ( .A(n40314), .B(n40313), .Z(n40305) );
  XOR U41105 ( .A(n40306), .B(n40305), .Z(n40307) );
  XNOR U41106 ( .A(n40308), .B(n40307), .Z(n40299) );
  AND U41107 ( .A(x[494]), .B(y[8110]), .Z(n41935) );
  NAND U41108 ( .A(n40246), .B(n41935), .Z(n40202) );
  NAND U41109 ( .A(n40200), .B(n40199), .Z(n40201) );
  NAND U41110 ( .A(n40202), .B(n40201), .Z(n40274) );
  AND U41111 ( .A(x[488]), .B(y[8107]), .Z(n40203) );
  NANDN U41112 ( .A(n40204), .B(n40203), .Z(n40207) );
  NAND U41113 ( .A(n40205), .B(n40466), .Z(n40206) );
  NAND U41114 ( .A(n40207), .B(n40206), .Z(n40273) );
  XOR U41115 ( .A(n40274), .B(n40273), .Z(n40276) );
  AND U41116 ( .A(y[8101]), .B(x[490]), .Z(n40209) );
  NAND U41117 ( .A(y[8107]), .B(x[484]), .Z(n40208) );
  XNOR U41118 ( .A(n40209), .B(n40208), .Z(n40254) );
  AND U41119 ( .A(x[487]), .B(y[8104]), .Z(n40253) );
  XNOR U41120 ( .A(n40254), .B(n40253), .Z(n40261) );
  NAND U41121 ( .A(x[486]), .B(y[8105]), .Z(n40351) );
  XNOR U41122 ( .A(n40351), .B(n40259), .Z(n40260) );
  XNOR U41123 ( .A(n40261), .B(n40260), .Z(n40295) );
  AND U41124 ( .A(y[8109]), .B(x[482]), .Z(n40211) );
  NAND U41125 ( .A(y[8102]), .B(x[489]), .Z(n40210) );
  XNOR U41126 ( .A(n40211), .B(n40210), .Z(n40264) );
  AND U41127 ( .A(x[483]), .B(y[8108]), .Z(n40265) );
  XOR U41128 ( .A(n40264), .B(n40265), .Z(n40293) );
  AND U41129 ( .A(y[8110]), .B(x[481]), .Z(n40213) );
  NAND U41130 ( .A(y[8103]), .B(x[488]), .Z(n40212) );
  XNOR U41131 ( .A(n40213), .B(n40212), .Z(n40242) );
  NAND U41132 ( .A(x[494]), .B(y[8097]), .Z(n40270) );
  XOR U41133 ( .A(o[431]), .B(n40270), .Z(n40243) );
  XNOR U41134 ( .A(n40242), .B(n40243), .Z(n40294) );
  XOR U41135 ( .A(n40293), .B(n40294), .Z(n40296) );
  XOR U41136 ( .A(n40295), .B(n40296), .Z(n40275) );
  XNOR U41137 ( .A(n40276), .B(n40275), .Z(n40318) );
  NAND U41138 ( .A(n40573), .B(n40214), .Z(n40218) );
  NAND U41139 ( .A(n40216), .B(n40215), .Z(n40217) );
  AND U41140 ( .A(n40218), .B(n40217), .Z(n40317) );
  XOR U41141 ( .A(n40318), .B(n40317), .Z(n40319) );
  NAND U41142 ( .A(n40220), .B(n40219), .Z(n40224) );
  NAND U41143 ( .A(n40222), .B(n40221), .Z(n40223) );
  AND U41144 ( .A(n40224), .B(n40223), .Z(n40320) );
  XOR U41145 ( .A(n40319), .B(n40320), .Z(n40300) );
  XOR U41146 ( .A(n40299), .B(n40300), .Z(n40301) );
  XOR U41147 ( .A(n40302), .B(n40301), .Z(n40233) );
  NANDN U41148 ( .A(n40226), .B(n40225), .Z(n40230) );
  NAND U41149 ( .A(n40228), .B(n40227), .Z(n40229) );
  AND U41150 ( .A(n40230), .B(n40229), .Z(n40232) );
  XOR U41151 ( .A(n40234), .B(n40235), .Z(n40240) );
  XNOR U41152 ( .A(n40239), .B(n40240), .Z(n40231) );
  XOR U41153 ( .A(n40238), .B(n40231), .Z(N880) );
  NANDN U41154 ( .A(n40233), .B(n40232), .Z(n40237) );
  NAND U41155 ( .A(n40235), .B(n40234), .Z(n40236) );
  AND U41156 ( .A(n40237), .B(n40236), .Z(n40412) );
  AND U41157 ( .A(x[488]), .B(y[8110]), .Z(n40574) );
  NAND U41158 ( .A(n40574), .B(n40241), .Z(n40245) );
  NANDN U41159 ( .A(n40243), .B(n40242), .Z(n40244) );
  AND U41160 ( .A(n40245), .B(n40244), .Z(n40377) );
  AND U41161 ( .A(x[495]), .B(y[8111]), .Z(n42345) );
  NAND U41162 ( .A(n42345), .B(n40246), .Z(n40250) );
  NAND U41163 ( .A(n40248), .B(n40247), .Z(n40249) );
  NAND U41164 ( .A(n40250), .B(n40249), .Z(n40376) );
  XNOR U41165 ( .A(n40377), .B(n40376), .Z(n40379) );
  AND U41166 ( .A(x[490]), .B(y[8107]), .Z(n40252) );
  NAND U41167 ( .A(n40252), .B(n40251), .Z(n40256) );
  NAND U41168 ( .A(n40254), .B(n40253), .Z(n40255) );
  NAND U41169 ( .A(n40256), .B(n40255), .Z(n40338) );
  AND U41170 ( .A(x[480]), .B(y[8112]), .Z(n40356) );
  NAND U41171 ( .A(x[496]), .B(y[8096]), .Z(n40357) );
  XNOR U41172 ( .A(n40356), .B(n40357), .Z(n40358) );
  NAND U41173 ( .A(x[495]), .B(y[8097]), .Z(n40348) );
  XOR U41174 ( .A(o[432]), .B(n40348), .Z(n40359) );
  XNOR U41175 ( .A(n40358), .B(n40359), .Z(n40337) );
  NAND U41176 ( .A(y[8105]), .B(x[487]), .Z(n40257) );
  XNOR U41177 ( .A(n40258), .B(n40257), .Z(n40353) );
  AND U41178 ( .A(x[490]), .B(y[8102]), .Z(n40352) );
  XOR U41179 ( .A(n40353), .B(n40352), .Z(n40336) );
  XOR U41180 ( .A(n40337), .B(n40336), .Z(n40339) );
  XOR U41181 ( .A(n40338), .B(n40339), .Z(n40378) );
  XNOR U41182 ( .A(n40379), .B(n40378), .Z(n40333) );
  NANDN U41183 ( .A(n40259), .B(n40351), .Z(n40263) );
  NAND U41184 ( .A(n40261), .B(n40260), .Z(n40262) );
  NAND U41185 ( .A(n40263), .B(n40262), .Z(n40331) );
  NAND U41186 ( .A(x[489]), .B(y[8109]), .Z(n41089) );
  NANDN U41187 ( .A(n41089), .B(n40658), .Z(n40267) );
  NAND U41188 ( .A(n40265), .B(n40264), .Z(n40266) );
  AND U41189 ( .A(n40267), .B(n40266), .Z(n40367) );
  AND U41190 ( .A(y[8111]), .B(x[481]), .Z(n40269) );
  NAND U41191 ( .A(y[8104]), .B(x[488]), .Z(n40268) );
  XNOR U41192 ( .A(n40269), .B(n40268), .Z(n40355) );
  ANDN U41193 ( .B(o[431]), .A(n40270), .Z(n40354) );
  XOR U41194 ( .A(n40355), .B(n40354), .Z(n40364) );
  NAND U41195 ( .A(y[8098]), .B(x[494]), .Z(n40271) );
  XNOR U41196 ( .A(n40272), .B(n40271), .Z(n40388) );
  NAND U41197 ( .A(x[484]), .B(y[8108]), .Z(n40389) );
  XNOR U41198 ( .A(n40388), .B(n40389), .Z(n40365) );
  XOR U41199 ( .A(n40364), .B(n40365), .Z(n40366) );
  XOR U41200 ( .A(n40367), .B(n40366), .Z(n40330) );
  XOR U41201 ( .A(n40331), .B(n40330), .Z(n40332) );
  XOR U41202 ( .A(n40333), .B(n40332), .Z(n40370) );
  NAND U41203 ( .A(n40274), .B(n40273), .Z(n40278) );
  NAND U41204 ( .A(n40276), .B(n40275), .Z(n40277) );
  AND U41205 ( .A(n40278), .B(n40277), .Z(n40371) );
  XOR U41206 ( .A(n40370), .B(n40371), .Z(n40373) );
  NAND U41207 ( .A(n40280), .B(n40279), .Z(n40284) );
  NAND U41208 ( .A(n40282), .B(n40281), .Z(n40283) );
  NAND U41209 ( .A(n40284), .B(n40283), .Z(n40403) );
  AND U41210 ( .A(x[493]), .B(y[8100]), .Z(n40399) );
  NAND U41211 ( .A(n40903), .B(n40399), .Z(n40288) );
  NAND U41212 ( .A(n40286), .B(n40285), .Z(n40287) );
  AND U41213 ( .A(n40288), .B(n40287), .Z(n40384) );
  AND U41214 ( .A(y[8110]), .B(x[482]), .Z(n40290) );
  NAND U41215 ( .A(y[8103]), .B(x[489]), .Z(n40289) );
  XNOR U41216 ( .A(n40290), .B(n40289), .Z(n40392) );
  NAND U41217 ( .A(x[483]), .B(y[8109]), .Z(n40393) );
  XNOR U41218 ( .A(n40392), .B(n40393), .Z(n40382) );
  AND U41219 ( .A(x[492]), .B(y[8100]), .Z(n41077) );
  AND U41220 ( .A(y[8107]), .B(x[485]), .Z(n40292) );
  NAND U41221 ( .A(y[8099]), .B(x[493]), .Z(n40291) );
  XOR U41222 ( .A(n40292), .B(n40291), .Z(n40343) );
  XOR U41223 ( .A(n41077), .B(n40343), .Z(n40383) );
  XOR U41224 ( .A(n40382), .B(n40383), .Z(n40385) );
  XNOR U41225 ( .A(n40384), .B(n40385), .Z(n40401) );
  NAND U41226 ( .A(n40294), .B(n40293), .Z(n40298) );
  NAND U41227 ( .A(n40296), .B(n40295), .Z(n40297) );
  AND U41228 ( .A(n40298), .B(n40297), .Z(n40400) );
  XOR U41229 ( .A(n40401), .B(n40400), .Z(n40402) );
  XOR U41230 ( .A(n40403), .B(n40402), .Z(n40372) );
  XNOR U41231 ( .A(n40373), .B(n40372), .Z(n40407) );
  NAND U41232 ( .A(n40300), .B(n40299), .Z(n40304) );
  NAND U41233 ( .A(n40302), .B(n40301), .Z(n40303) );
  AND U41234 ( .A(n40304), .B(n40303), .Z(n40406) );
  XOR U41235 ( .A(n40407), .B(n40406), .Z(n40409) );
  NAND U41236 ( .A(n40306), .B(n40305), .Z(n40310) );
  NAND U41237 ( .A(n40308), .B(n40307), .Z(n40309) );
  NAND U41238 ( .A(n40310), .B(n40309), .Z(n40327) );
  NAND U41239 ( .A(n40312), .B(n40311), .Z(n40316) );
  NAND U41240 ( .A(n40314), .B(n40313), .Z(n40315) );
  NAND U41241 ( .A(n40316), .B(n40315), .Z(n40325) );
  NAND U41242 ( .A(n40318), .B(n40317), .Z(n40322) );
  NAND U41243 ( .A(n40320), .B(n40319), .Z(n40321) );
  AND U41244 ( .A(n40322), .B(n40321), .Z(n40324) );
  XOR U41245 ( .A(n40325), .B(n40324), .Z(n40326) );
  XOR U41246 ( .A(n40327), .B(n40326), .Z(n40408) );
  XOR U41247 ( .A(n40409), .B(n40408), .Z(n40414) );
  XNOR U41248 ( .A(n40413), .B(n40414), .Z(n40323) );
  XOR U41249 ( .A(n40412), .B(n40323), .Z(N881) );
  NAND U41250 ( .A(n40325), .B(n40324), .Z(n40329) );
  NAND U41251 ( .A(n40327), .B(n40326), .Z(n40328) );
  AND U41252 ( .A(n40329), .B(n40328), .Z(n40512) );
  NAND U41253 ( .A(n40331), .B(n40330), .Z(n40335) );
  NAND U41254 ( .A(n40333), .B(n40332), .Z(n40334) );
  NAND U41255 ( .A(n40335), .B(n40334), .Z(n40425) );
  NAND U41256 ( .A(n40337), .B(n40336), .Z(n40341) );
  NAND U41257 ( .A(n40339), .B(n40338), .Z(n40340) );
  AND U41258 ( .A(n40341), .B(n40340), .Z(n40502) );
  AND U41259 ( .A(x[493]), .B(y[8107]), .Z(n41316) );
  NAND U41260 ( .A(n41316), .B(n40342), .Z(n40345) );
  NANDN U41261 ( .A(n40343), .B(n41077), .Z(n40344) );
  AND U41262 ( .A(n40345), .B(n40344), .Z(n40455) );
  AND U41263 ( .A(y[8112]), .B(x[481]), .Z(n40347) );
  NAND U41264 ( .A(y[8104]), .B(x[489]), .Z(n40346) );
  XNOR U41265 ( .A(n40347), .B(n40346), .Z(n40472) );
  ANDN U41266 ( .B(o[432]), .A(n40348), .Z(n40471) );
  XOR U41267 ( .A(n40472), .B(n40471), .Z(n40453) );
  AND U41268 ( .A(y[8098]), .B(x[495]), .Z(n40350) );
  NAND U41269 ( .A(y[8101]), .B(x[492]), .Z(n40349) );
  XNOR U41270 ( .A(n40350), .B(n40349), .Z(n40429) );
  AND U41271 ( .A(x[494]), .B(y[8099]), .Z(n40428) );
  XOR U41272 ( .A(n40429), .B(n40428), .Z(n40452) );
  XOR U41273 ( .A(n40453), .B(n40452), .Z(n40454) );
  XNOR U41274 ( .A(n40455), .B(n40454), .Z(n40500) );
  NAND U41275 ( .A(x[487]), .B(y[8106]), .Z(n40483) );
  NAND U41276 ( .A(x[488]), .B(y[8111]), .Z(n41158) );
  AND U41277 ( .A(x[481]), .B(y[8104]), .Z(n40552) );
  XNOR U41278 ( .A(n40461), .B(n40460), .Z(n40462) );
  NANDN U41279 ( .A(n40357), .B(n40356), .Z(n40361) );
  NANDN U41280 ( .A(n40359), .B(n40358), .Z(n40360) );
  AND U41281 ( .A(n40361), .B(n40360), .Z(n40459) );
  AND U41282 ( .A(x[480]), .B(y[8113]), .Z(n40443) );
  AND U41283 ( .A(x[497]), .B(y[8096]), .Z(n40442) );
  XOR U41284 ( .A(n40443), .B(n40442), .Z(n40445) );
  AND U41285 ( .A(x[496]), .B(y[8097]), .Z(n40439) );
  XOR U41286 ( .A(n40439), .B(o[433]), .Z(n40444) );
  XOR U41287 ( .A(n40445), .B(n40444), .Z(n40457) );
  AND U41288 ( .A(y[8111]), .B(x[482]), .Z(n40363) );
  NAND U41289 ( .A(y[8103]), .B(x[490]), .Z(n40362) );
  XNOR U41290 ( .A(n40363), .B(n40362), .Z(n40476) );
  NAND U41291 ( .A(x[483]), .B(y[8110]), .Z(n40477) );
  XOR U41292 ( .A(n40457), .B(n40456), .Z(n40458) );
  XOR U41293 ( .A(n40459), .B(n40458), .Z(n40463) );
  XOR U41294 ( .A(n40462), .B(n40463), .Z(n40501) );
  XOR U41295 ( .A(n40500), .B(n40501), .Z(n40503) );
  XNOR U41296 ( .A(n40502), .B(n40503), .Z(n40423) );
  NAND U41297 ( .A(n40365), .B(n40364), .Z(n40369) );
  NANDN U41298 ( .A(n40367), .B(n40366), .Z(n40368) );
  AND U41299 ( .A(n40369), .B(n40368), .Z(n40422) );
  XOR U41300 ( .A(n40423), .B(n40422), .Z(n40424) );
  XNOR U41301 ( .A(n40425), .B(n40424), .Z(n40510) );
  NAND U41302 ( .A(n40371), .B(n40370), .Z(n40375) );
  NAND U41303 ( .A(n40373), .B(n40372), .Z(n40374) );
  AND U41304 ( .A(n40375), .B(n40374), .Z(n40419) );
  NANDN U41305 ( .A(n40377), .B(n40376), .Z(n40381) );
  NAND U41306 ( .A(n40379), .B(n40378), .Z(n40380) );
  AND U41307 ( .A(n40381), .B(n40380), .Z(n40496) );
  NANDN U41308 ( .A(n40383), .B(n40382), .Z(n40387) );
  OR U41309 ( .A(n40385), .B(n40384), .Z(n40386) );
  AND U41310 ( .A(n40387), .B(n40386), .Z(n40495) );
  NAND U41311 ( .A(x[494]), .B(y[8101]), .Z(n40693) );
  NANDN U41312 ( .A(n40693), .B(n40903), .Z(n40391) );
  NANDN U41313 ( .A(n40389), .B(n40388), .Z(n40390) );
  AND U41314 ( .A(n40391), .B(n40390), .Z(n40489) );
  AND U41315 ( .A(x[489]), .B(y[8110]), .Z(n41297) );
  NAND U41316 ( .A(n40475), .B(n41297), .Z(n40395) );
  NANDN U41317 ( .A(n40393), .B(n40392), .Z(n40394) );
  NAND U41318 ( .A(n40395), .B(n40394), .Z(n40488) );
  XNOR U41319 ( .A(n40489), .B(n40488), .Z(n40490) );
  AND U41320 ( .A(x[485]), .B(y[8108]), .Z(n40534) );
  NAND U41321 ( .A(y[8105]), .B(x[488]), .Z(n40396) );
  XNOR U41322 ( .A(n40534), .B(n40396), .Z(n40467) );
  XOR U41323 ( .A(n40467), .B(n40397), .Z(n40482) );
  XNOR U41324 ( .A(n40482), .B(n40483), .Z(n40484) );
  NAND U41325 ( .A(y[8109]), .B(x[484]), .Z(n40398) );
  XNOR U41326 ( .A(n40399), .B(n40398), .Z(n40433) );
  NAND U41327 ( .A(x[491]), .B(y[8102]), .Z(n40434) );
  XOR U41328 ( .A(n40433), .B(n40434), .Z(n40485) );
  XOR U41329 ( .A(n40484), .B(n40485), .Z(n40491) );
  XNOR U41330 ( .A(n40490), .B(n40491), .Z(n40494) );
  XOR U41331 ( .A(n40495), .B(n40494), .Z(n40497) );
  XNOR U41332 ( .A(n40496), .B(n40497), .Z(n40417) );
  NAND U41333 ( .A(n40401), .B(n40400), .Z(n40405) );
  NAND U41334 ( .A(n40403), .B(n40402), .Z(n40404) );
  NAND U41335 ( .A(n40405), .B(n40404), .Z(n40416) );
  XOR U41336 ( .A(n40417), .B(n40416), .Z(n40418) );
  XOR U41337 ( .A(n40419), .B(n40418), .Z(n40509) );
  XOR U41338 ( .A(n40510), .B(n40509), .Z(n40511) );
  XOR U41339 ( .A(n40512), .B(n40511), .Z(n40508) );
  NAND U41340 ( .A(n40407), .B(n40406), .Z(n40411) );
  NAND U41341 ( .A(n40409), .B(n40408), .Z(n40410) );
  NAND U41342 ( .A(n40411), .B(n40410), .Z(n40507) );
  XOR U41343 ( .A(n40507), .B(n40506), .Z(n40415) );
  XNOR U41344 ( .A(n40508), .B(n40415), .Z(N882) );
  NAND U41345 ( .A(n40417), .B(n40416), .Z(n40421) );
  NANDN U41346 ( .A(n40419), .B(n40418), .Z(n40420) );
  AND U41347 ( .A(n40421), .B(n40420), .Z(n40621) );
  NAND U41348 ( .A(n40423), .B(n40422), .Z(n40427) );
  NAND U41349 ( .A(n40425), .B(n40424), .Z(n40426) );
  AND U41350 ( .A(n40427), .B(n40426), .Z(n40618) );
  AND U41351 ( .A(x[495]), .B(y[8101]), .Z(n40666) );
  AND U41352 ( .A(x[492]), .B(y[8098]), .Z(n40762) );
  NAND U41353 ( .A(n40666), .B(n40762), .Z(n40431) );
  NAND U41354 ( .A(n40429), .B(n40428), .Z(n40430) );
  NAND U41355 ( .A(n40431), .B(n40430), .Z(n40600) );
  NAND U41356 ( .A(n41680), .B(n40432), .Z(n40436) );
  NANDN U41357 ( .A(n40434), .B(n40433), .Z(n40435) );
  AND U41358 ( .A(n40436), .B(n40435), .Z(n40591) );
  AND U41359 ( .A(y[8113]), .B(x[481]), .Z(n40438) );
  NAND U41360 ( .A(y[8104]), .B(x[490]), .Z(n40437) );
  XNOR U41361 ( .A(n40438), .B(n40437), .Z(n40553) );
  NAND U41362 ( .A(n40439), .B(o[433]), .Z(n40554) );
  AND U41363 ( .A(y[8099]), .B(x[495]), .Z(n40441) );
  NAND U41364 ( .A(y[8105]), .B(x[489]), .Z(n40440) );
  XNOR U41365 ( .A(n40441), .B(n40440), .Z(n40544) );
  NAND U41366 ( .A(x[494]), .B(y[8100]), .Z(n40545) );
  XOR U41367 ( .A(n40589), .B(n40588), .Z(n40590) );
  XOR U41368 ( .A(n40600), .B(n40601), .Z(n40603) );
  NAND U41369 ( .A(n40443), .B(n40442), .Z(n40447) );
  NAND U41370 ( .A(n40445), .B(n40444), .Z(n40446) );
  NAND U41371 ( .A(n40447), .B(n40446), .Z(n40612) );
  AND U41372 ( .A(y[8098]), .B(x[496]), .Z(n40449) );
  NAND U41373 ( .A(y[8103]), .B(x[491]), .Z(n40448) );
  XNOR U41374 ( .A(n40449), .B(n40448), .Z(n40540) );
  NAND U41375 ( .A(x[482]), .B(y[8112]), .Z(n40541) );
  XOR U41376 ( .A(n40612), .B(n40613), .Z(n40615) );
  AND U41377 ( .A(x[485]), .B(y[8109]), .Z(n40674) );
  NAND U41378 ( .A(y[8108]), .B(x[486]), .Z(n40450) );
  XNOR U41379 ( .A(n40674), .B(n40450), .Z(n40537) );
  NAND U41380 ( .A(y[8110]), .B(x[484]), .Z(n40451) );
  XNOR U41381 ( .A(n41302), .B(n40451), .Z(n40575) );
  NAND U41382 ( .A(x[487]), .B(y[8107]), .Z(n40576) );
  XOR U41383 ( .A(n40537), .B(n40536), .Z(n40614) );
  XOR U41384 ( .A(n40615), .B(n40614), .Z(n40602) );
  XOR U41385 ( .A(n40603), .B(n40602), .Z(n40523) );
  XOR U41386 ( .A(n40595), .B(n40594), .Z(n40597) );
  NANDN U41387 ( .A(n40461), .B(n40460), .Z(n40465) );
  NANDN U41388 ( .A(n40463), .B(n40462), .Z(n40464) );
  AND U41389 ( .A(n40465), .B(n40464), .Z(n40596) );
  XOR U41390 ( .A(n40597), .B(n40596), .Z(n40522) );
  XNOR U41391 ( .A(n40523), .B(n40522), .Z(n40525) );
  AND U41392 ( .A(x[488]), .B(y[8108]), .Z(n40802) );
  NAND U41393 ( .A(n40802), .B(n40466), .Z(n40470) );
  NANDN U41394 ( .A(n40468), .B(n40467), .Z(n40469) );
  NAND U41395 ( .A(n40470), .B(n40469), .Z(n40607) );
  AND U41396 ( .A(x[489]), .B(y[8112]), .Z(n41443) );
  NAND U41397 ( .A(n41443), .B(n40552), .Z(n40474) );
  NAND U41398 ( .A(n40472), .B(n40471), .Z(n40473) );
  NAND U41399 ( .A(n40474), .B(n40473), .Z(n40606) );
  XOR U41400 ( .A(n40607), .B(n40606), .Z(n40609) );
  AND U41401 ( .A(x[490]), .B(y[8111]), .Z(n41325) );
  IV U41402 ( .A(n41325), .Z(n41442) );
  NANDN U41403 ( .A(n41442), .B(n40475), .Z(n40479) );
  NANDN U41404 ( .A(n40477), .B(n40476), .Z(n40478) );
  AND U41405 ( .A(n40479), .B(n40478), .Z(n40585) );
  AND U41406 ( .A(y[8101]), .B(x[493]), .Z(n40481) );
  NAND U41407 ( .A(y[8111]), .B(x[483]), .Z(n40480) );
  XNOR U41408 ( .A(n40481), .B(n40480), .Z(n40565) );
  NAND U41409 ( .A(x[492]), .B(y[8102]), .Z(n40566) );
  AND U41410 ( .A(x[480]), .B(y[8114]), .Z(n40557) );
  NAND U41411 ( .A(x[498]), .B(y[8096]), .Z(n40558) );
  NAND U41412 ( .A(x[497]), .B(y[8097]), .Z(n40579) );
  XOR U41413 ( .A(n40560), .B(n40559), .Z(n40582) );
  XOR U41414 ( .A(n40583), .B(n40582), .Z(n40584) );
  XOR U41415 ( .A(n40609), .B(n40608), .Z(n40529) );
  NANDN U41416 ( .A(n40483), .B(n40482), .Z(n40487) );
  NANDN U41417 ( .A(n40485), .B(n40484), .Z(n40486) );
  AND U41418 ( .A(n40487), .B(n40486), .Z(n40528) );
  NANDN U41419 ( .A(n40489), .B(n40488), .Z(n40493) );
  NANDN U41420 ( .A(n40491), .B(n40490), .Z(n40492) );
  NAND U41421 ( .A(n40493), .B(n40492), .Z(n40531) );
  XOR U41422 ( .A(n40525), .B(n40524), .Z(n40519) );
  NANDN U41423 ( .A(n40495), .B(n40494), .Z(n40499) );
  OR U41424 ( .A(n40497), .B(n40496), .Z(n40498) );
  AND U41425 ( .A(n40499), .B(n40498), .Z(n40517) );
  NANDN U41426 ( .A(n40501), .B(n40500), .Z(n40505) );
  OR U41427 ( .A(n40503), .B(n40502), .Z(n40504) );
  NAND U41428 ( .A(n40505), .B(n40504), .Z(n40516) );
  XNOR U41429 ( .A(n40517), .B(n40516), .Z(n40518) );
  XNOR U41430 ( .A(n40519), .B(n40518), .Z(n40619) );
  XOR U41431 ( .A(n40618), .B(n40619), .Z(n40620) );
  XOR U41432 ( .A(n40621), .B(n40620), .Z(n40627) );
  NAND U41433 ( .A(n40510), .B(n40509), .Z(n40514) );
  NANDN U41434 ( .A(n40512), .B(n40511), .Z(n40513) );
  AND U41435 ( .A(n40514), .B(n40513), .Z(n40626) );
  IV U41436 ( .A(n40626), .Z(n40624) );
  XOR U41437 ( .A(n40625), .B(n40624), .Z(n40515) );
  XNOR U41438 ( .A(n40627), .B(n40515), .Z(N883) );
  NANDN U41439 ( .A(n40517), .B(n40516), .Z(n40521) );
  NANDN U41440 ( .A(n40519), .B(n40518), .Z(n40520) );
  AND U41441 ( .A(n40521), .B(n40520), .Z(n40635) );
  NANDN U41442 ( .A(n40523), .B(n40522), .Z(n40527) );
  NAND U41443 ( .A(n40525), .B(n40524), .Z(n40526) );
  AND U41444 ( .A(n40527), .B(n40526), .Z(n40632) );
  NANDN U41445 ( .A(n40529), .B(n40528), .Z(n40533) );
  NANDN U41446 ( .A(n40531), .B(n40530), .Z(n40532) );
  AND U41447 ( .A(n40533), .B(n40532), .Z(n40734) );
  AND U41448 ( .A(x[486]), .B(y[8109]), .Z(n40535) );
  NAND U41449 ( .A(n40535), .B(n40534), .Z(n40539) );
  NAND U41450 ( .A(n40537), .B(n40536), .Z(n40538) );
  AND U41451 ( .A(n40539), .B(n40538), .Z(n40728) );
  AND U41452 ( .A(x[496]), .B(y[8103]), .Z(n41093) );
  NAND U41453 ( .A(n41093), .B(n40903), .Z(n40543) );
  NANDN U41454 ( .A(n40541), .B(n40540), .Z(n40542) );
  AND U41455 ( .A(n40543), .B(n40542), .Z(n40726) );
  AND U41456 ( .A(x[495]), .B(y[8105]), .Z(n41328) );
  NAND U41457 ( .A(n41328), .B(n40653), .Z(n40547) );
  NANDN U41458 ( .A(n40545), .B(n40544), .Z(n40546) );
  AND U41459 ( .A(n40547), .B(n40546), .Z(n40644) );
  AND U41460 ( .A(y[8114]), .B(x[481]), .Z(n40549) );
  NAND U41461 ( .A(y[8107]), .B(x[488]), .Z(n40548) );
  XNOR U41462 ( .A(n40549), .B(n40548), .Z(n40692) );
  AND U41463 ( .A(y[8102]), .B(x[493]), .Z(n40551) );
  NAND U41464 ( .A(y[8113]), .B(x[482]), .Z(n40550) );
  XNOR U41465 ( .A(n40551), .B(n40550), .Z(n40659) );
  XOR U41466 ( .A(n40642), .B(n40641), .Z(n40643) );
  AND U41467 ( .A(x[490]), .B(y[8113]), .Z(n41756) );
  NAND U41468 ( .A(n41756), .B(n40552), .Z(n40556) );
  NANDN U41469 ( .A(n40554), .B(n40553), .Z(n40555) );
  AND U41470 ( .A(n40556), .B(n40555), .Z(n40704) );
  NANDN U41471 ( .A(n40558), .B(n40557), .Z(n40562) );
  NAND U41472 ( .A(n40560), .B(n40559), .Z(n40561) );
  AND U41473 ( .A(n40562), .B(n40561), .Z(n40702) );
  AND U41474 ( .A(y[8099]), .B(x[496]), .Z(n41375) );
  NAND U41475 ( .A(y[8106]), .B(x[489]), .Z(n40563) );
  XNOR U41476 ( .A(n41375), .B(n40563), .Z(n40654) );
  NAND U41477 ( .A(x[495]), .B(y[8100]), .Z(n40655) );
  AND U41478 ( .A(x[493]), .B(y[8111]), .Z(n41964) );
  NANDN U41479 ( .A(n40564), .B(n41964), .Z(n40568) );
  NANDN U41480 ( .A(n40566), .B(n40565), .Z(n40567) );
  AND U41481 ( .A(n40568), .B(n40567), .Z(n40710) );
  AND U41482 ( .A(y[8105]), .B(x[490]), .Z(n40570) );
  NAND U41483 ( .A(y[8098]), .B(x[497]), .Z(n40569) );
  XNOR U41484 ( .A(n40570), .B(n40569), .Z(n40698) );
  AND U41485 ( .A(x[498]), .B(y[8097]), .Z(n40673) );
  XOR U41486 ( .A(o[435]), .B(n40673), .Z(n40697) );
  XOR U41487 ( .A(n40698), .B(n40697), .Z(n40708) );
  NAND U41488 ( .A(y[8112]), .B(x[483]), .Z(n40571) );
  XNOR U41489 ( .A(n40572), .B(n40571), .Z(n40667) );
  XOR U41490 ( .A(n40708), .B(n40707), .Z(n40709) );
  NAND U41491 ( .A(n40574), .B(n40573), .Z(n40578) );
  NANDN U41492 ( .A(n40576), .B(n40575), .Z(n40577) );
  AND U41493 ( .A(n40578), .B(n40577), .Z(n40650) );
  AND U41494 ( .A(x[480]), .B(y[8115]), .Z(n40678) );
  NAND U41495 ( .A(x[499]), .B(y[8096]), .Z(n40679) );
  ANDN U41496 ( .B(o[434]), .A(n40579), .Z(n40680) );
  XOR U41497 ( .A(n40681), .B(n40680), .Z(n40648) );
  AND U41498 ( .A(x[484]), .B(y[8111]), .Z(n40816) );
  AND U41499 ( .A(y[8110]), .B(x[485]), .Z(n40581) );
  NAND U41500 ( .A(y[8109]), .B(x[486]), .Z(n40580) );
  XOR U41501 ( .A(n40581), .B(n40580), .Z(n40675) );
  XOR U41502 ( .A(n40648), .B(n40647), .Z(n40649) );
  XOR U41503 ( .A(n40650), .B(n40649), .Z(n40719) );
  XOR U41504 ( .A(n40720), .B(n40719), .Z(n40722) );
  XNOR U41505 ( .A(n40721), .B(n40722), .Z(n40715) );
  NAND U41506 ( .A(n40583), .B(n40582), .Z(n40587) );
  NANDN U41507 ( .A(n40585), .B(n40584), .Z(n40586) );
  AND U41508 ( .A(n40587), .B(n40586), .Z(n40714) );
  NAND U41509 ( .A(n40589), .B(n40588), .Z(n40593) );
  NANDN U41510 ( .A(n40591), .B(n40590), .Z(n40592) );
  NAND U41511 ( .A(n40593), .B(n40592), .Z(n40713) );
  XNOR U41512 ( .A(n40715), .B(n40716), .Z(n40731) );
  XOR U41513 ( .A(n40732), .B(n40731), .Z(n40733) );
  NAND U41514 ( .A(n40595), .B(n40594), .Z(n40599) );
  NAND U41515 ( .A(n40597), .B(n40596), .Z(n40598) );
  AND U41516 ( .A(n40599), .B(n40598), .Z(n40743) );
  NAND U41517 ( .A(n40601), .B(n40600), .Z(n40605) );
  NAND U41518 ( .A(n40603), .B(n40602), .Z(n40604) );
  NAND U41519 ( .A(n40605), .B(n40604), .Z(n40739) );
  NAND U41520 ( .A(n40607), .B(n40606), .Z(n40611) );
  NAND U41521 ( .A(n40609), .B(n40608), .Z(n40610) );
  NAND U41522 ( .A(n40611), .B(n40610), .Z(n40738) );
  NAND U41523 ( .A(n40613), .B(n40612), .Z(n40617) );
  NAND U41524 ( .A(n40615), .B(n40614), .Z(n40616) );
  NAND U41525 ( .A(n40617), .B(n40616), .Z(n40737) );
  XNOR U41526 ( .A(n40738), .B(n40737), .Z(n40740) );
  XNOR U41527 ( .A(n40743), .B(n40744), .Z(n40745) );
  XNOR U41528 ( .A(n40632), .B(n40633), .Z(n40634) );
  XOR U41529 ( .A(n40635), .B(n40634), .Z(n40640) );
  NAND U41530 ( .A(n40619), .B(n40618), .Z(n40623) );
  NAND U41531 ( .A(n40621), .B(n40620), .Z(n40622) );
  NAND U41532 ( .A(n40623), .B(n40622), .Z(n40639) );
  NANDN U41533 ( .A(n40624), .B(n40625), .Z(n40630) );
  NOR U41534 ( .A(n40626), .B(n40625), .Z(n40628) );
  OR U41535 ( .A(n40628), .B(n40627), .Z(n40629) );
  AND U41536 ( .A(n40630), .B(n40629), .Z(n40638) );
  XOR U41537 ( .A(n40639), .B(n40638), .Z(n40631) );
  XNOR U41538 ( .A(n40640), .B(n40631), .Z(N884) );
  NANDN U41539 ( .A(n40633), .B(n40632), .Z(n40637) );
  NANDN U41540 ( .A(n40635), .B(n40634), .Z(n40636) );
  AND U41541 ( .A(n40637), .B(n40636), .Z(n40865) );
  NAND U41542 ( .A(n40642), .B(n40641), .Z(n40646) );
  NANDN U41543 ( .A(n40644), .B(n40643), .Z(n40645) );
  AND U41544 ( .A(n40646), .B(n40645), .Z(n40751) );
  NAND U41545 ( .A(n40648), .B(n40647), .Z(n40652) );
  NANDN U41546 ( .A(n40650), .B(n40649), .Z(n40651) );
  NAND U41547 ( .A(n40652), .B(n40651), .Z(n40750) );
  AND U41548 ( .A(x[496]), .B(y[8106]), .Z(n41644) );
  NAND U41549 ( .A(n41644), .B(n40653), .Z(n40657) );
  NANDN U41550 ( .A(n40655), .B(n40654), .Z(n40656) );
  AND U41551 ( .A(n40657), .B(n40656), .Z(n40791) );
  AND U41552 ( .A(x[493]), .B(y[8113]), .Z(n42186) );
  NAND U41553 ( .A(n42186), .B(n40658), .Z(n40662) );
  NANDN U41554 ( .A(n40660), .B(n40659), .Z(n40661) );
  AND U41555 ( .A(n40662), .B(n40661), .Z(n40836) );
  AND U41556 ( .A(y[8100]), .B(x[496]), .Z(n40664) );
  NAND U41557 ( .A(y[8106]), .B(x[490]), .Z(n40663) );
  XNOR U41558 ( .A(n40664), .B(n40663), .Z(n40797) );
  AND U41559 ( .A(x[482]), .B(y[8114]), .Z(n40798) );
  XOR U41560 ( .A(n40797), .B(n40798), .Z(n40834) );
  NAND U41561 ( .A(y[8107]), .B(x[489]), .Z(n40665) );
  XNOR U41562 ( .A(n40666), .B(n40665), .Z(n40773) );
  AND U41563 ( .A(x[494]), .B(y[8102]), .Z(n40774) );
  XOR U41564 ( .A(n40773), .B(n40774), .Z(n40833) );
  XOR U41565 ( .A(n40834), .B(n40833), .Z(n40835) );
  AND U41566 ( .A(x[491]), .B(y[8112]), .Z(n41757) );
  NANDN U41567 ( .A(n40930), .B(n41757), .Z(n40670) );
  NANDN U41568 ( .A(n40668), .B(n40667), .Z(n40669) );
  AND U41569 ( .A(n40670), .B(n40669), .Z(n40842) );
  AND U41570 ( .A(y[8105]), .B(x[491]), .Z(n40672) );
  NAND U41571 ( .A(y[8115]), .B(x[481]), .Z(n40671) );
  XNOR U41572 ( .A(n40672), .B(n40671), .Z(n40769) );
  AND U41573 ( .A(x[499]), .B(y[8097]), .Z(n40777) );
  XOR U41574 ( .A(o[436]), .B(n40777), .Z(n40768) );
  XOR U41575 ( .A(n40769), .B(n40768), .Z(n40840) );
  AND U41576 ( .A(x[480]), .B(y[8116]), .Z(n40821) );
  AND U41577 ( .A(x[500]), .B(y[8096]), .Z(n40822) );
  XOR U41578 ( .A(n40821), .B(n40822), .Z(n40824) );
  AND U41579 ( .A(o[435]), .B(n40673), .Z(n40823) );
  XOR U41580 ( .A(n40824), .B(n40823), .Z(n40839) );
  XOR U41581 ( .A(n40840), .B(n40839), .Z(n40841) );
  XOR U41582 ( .A(n40793), .B(n40792), .Z(n40752) );
  XOR U41583 ( .A(n40753), .B(n40752), .Z(n40848) );
  AND U41584 ( .A(x[486]), .B(y[8110]), .Z(n40757) );
  IV U41585 ( .A(n40757), .Z(n40690) );
  NANDN U41586 ( .A(n40690), .B(n40674), .Z(n40677) );
  NANDN U41587 ( .A(n40675), .B(n40816), .Z(n40676) );
  AND U41588 ( .A(n40677), .B(n40676), .Z(n40781) );
  NANDN U41589 ( .A(n40679), .B(n40678), .Z(n40683) );
  NAND U41590 ( .A(n40681), .B(n40680), .Z(n40682) );
  AND U41591 ( .A(n40683), .B(n40682), .Z(n40779) );
  AND U41592 ( .A(y[8098]), .B(x[498]), .Z(n40685) );
  NAND U41593 ( .A(y[8104]), .B(x[492]), .Z(n40684) );
  XNOR U41594 ( .A(n40685), .B(n40684), .Z(n40763) );
  AND U41595 ( .A(x[497]), .B(y[8099]), .Z(n40764) );
  XOR U41596 ( .A(n40763), .B(n40764), .Z(n40778) );
  AND U41597 ( .A(y[8103]), .B(x[493]), .Z(n40687) );
  NAND U41598 ( .A(y[8113]), .B(x[483]), .Z(n40686) );
  XNOR U41599 ( .A(n40687), .B(n40686), .Z(n40803) );
  XOR U41600 ( .A(n40803), .B(n40802), .Z(n40759) );
  AND U41601 ( .A(y[8111]), .B(x[485]), .Z(n40689) );
  NAND U41602 ( .A(y[8112]), .B(x[484]), .Z(n40688) );
  XNOR U41603 ( .A(n40689), .B(n40688), .Z(n40818) );
  AND U41604 ( .A(x[487]), .B(y[8109]), .Z(n40817) );
  XNOR U41605 ( .A(n40818), .B(n40817), .Z(n40756) );
  XOR U41606 ( .A(n40690), .B(n40756), .Z(n40758) );
  AND U41607 ( .A(x[488]), .B(y[8114]), .Z(n41915) );
  AND U41608 ( .A(x[481]), .B(y[8107]), .Z(n40691) );
  NAND U41609 ( .A(n41915), .B(n40691), .Z(n40695) );
  NANDN U41610 ( .A(n40693), .B(n40692), .Z(n40694) );
  AND U41611 ( .A(n40695), .B(n40694), .Z(n40828) );
  AND U41612 ( .A(x[497]), .B(y[8105]), .Z(n41653) );
  NAND U41613 ( .A(n41653), .B(n40696), .Z(n40700) );
  NAND U41614 ( .A(n40698), .B(n40697), .Z(n40699) );
  NAND U41615 ( .A(n40700), .B(n40699), .Z(n40827) );
  XNOR U41616 ( .A(n40829), .B(n40830), .Z(n40784) );
  XOR U41617 ( .A(n40785), .B(n40784), .Z(n40786) );
  NANDN U41618 ( .A(n40702), .B(n40701), .Z(n40706) );
  NANDN U41619 ( .A(n40704), .B(n40703), .Z(n40705) );
  NAND U41620 ( .A(n40706), .B(n40705), .Z(n40787) );
  NAND U41621 ( .A(n40708), .B(n40707), .Z(n40712) );
  NANDN U41622 ( .A(n40710), .B(n40709), .Z(n40711) );
  NAND U41623 ( .A(n40712), .B(n40711), .Z(n40846) );
  NANDN U41624 ( .A(n40714), .B(n40713), .Z(n40718) );
  NAND U41625 ( .A(n40716), .B(n40715), .Z(n40717) );
  AND U41626 ( .A(n40718), .B(n40717), .Z(n40860) );
  NAND U41627 ( .A(n40720), .B(n40719), .Z(n40724) );
  NAND U41628 ( .A(n40722), .B(n40721), .Z(n40723) );
  AND U41629 ( .A(n40724), .B(n40723), .Z(n40858) );
  NANDN U41630 ( .A(n40726), .B(n40725), .Z(n40730) );
  NANDN U41631 ( .A(n40728), .B(n40727), .Z(n40729) );
  AND U41632 ( .A(n40730), .B(n40729), .Z(n40857) );
  XNOR U41633 ( .A(n40860), .B(n40859), .Z(n40851) );
  XOR U41634 ( .A(n40852), .B(n40851), .Z(n40853) );
  NAND U41635 ( .A(n40732), .B(n40731), .Z(n40736) );
  NANDN U41636 ( .A(n40734), .B(n40733), .Z(n40735) );
  NAND U41637 ( .A(n40736), .B(n40735), .Z(n40854) );
  NAND U41638 ( .A(n40738), .B(n40737), .Z(n40742) );
  NANDN U41639 ( .A(n40740), .B(n40739), .Z(n40741) );
  AND U41640 ( .A(n40742), .B(n40741), .Z(n40867) );
  NANDN U41641 ( .A(n40744), .B(n40743), .Z(n40748) );
  NANDN U41642 ( .A(n40746), .B(n40745), .Z(n40747) );
  AND U41643 ( .A(n40748), .B(n40747), .Z(n40866) );
  XOR U41644 ( .A(n40867), .B(n40866), .Z(n40868) );
  XNOR U41645 ( .A(n40864), .B(n40863), .Z(n40749) );
  XOR U41646 ( .A(n40865), .B(n40749), .Z(N885) );
  NANDN U41647 ( .A(n40751), .B(n40750), .Z(n40755) );
  NAND U41648 ( .A(n40753), .B(n40752), .Z(n40754) );
  AND U41649 ( .A(n40755), .B(n40754), .Z(n40882) );
  NANDN U41650 ( .A(n40757), .B(n40756), .Z(n40761) );
  NANDN U41651 ( .A(n40759), .B(n40758), .Z(n40760) );
  AND U41652 ( .A(n40761), .B(n40760), .Z(n40971) );
  AND U41653 ( .A(x[498]), .B(y[8104]), .Z(n41651) );
  NAND U41654 ( .A(n41651), .B(n40762), .Z(n40766) );
  NAND U41655 ( .A(n40764), .B(n40763), .Z(n40765) );
  NAND U41656 ( .A(n40766), .B(n40765), .Z(n40953) );
  AND U41657 ( .A(x[491]), .B(y[8115]), .Z(n42407) );
  AND U41658 ( .A(x[481]), .B(y[8105]), .Z(n40767) );
  NAND U41659 ( .A(n42407), .B(n40767), .Z(n40771) );
  NAND U41660 ( .A(n40769), .B(n40768), .Z(n40770) );
  NAND U41661 ( .A(n40771), .B(n40770), .Z(n40952) );
  XOR U41662 ( .A(n40953), .B(n40952), .Z(n40955) );
  AND U41663 ( .A(x[495]), .B(y[8107]), .Z(n41639) );
  NAND U41664 ( .A(n41639), .B(n40772), .Z(n40776) );
  NAND U41665 ( .A(n40774), .B(n40773), .Z(n40775) );
  AND U41666 ( .A(n40776), .B(n40775), .Z(n40917) );
  AND U41667 ( .A(x[480]), .B(y[8117]), .Z(n40936) );
  AND U41668 ( .A(x[501]), .B(y[8096]), .Z(n40937) );
  XOR U41669 ( .A(n40936), .B(n40937), .Z(n40939) );
  AND U41670 ( .A(o[436]), .B(n40777), .Z(n40938) );
  XOR U41671 ( .A(n40939), .B(n40938), .Z(n40915) );
  AND U41672 ( .A(x[485]), .B(y[8112]), .Z(n40923) );
  AND U41673 ( .A(x[496]), .B(y[8101]), .Z(n40922) );
  XOR U41674 ( .A(n40923), .B(n40922), .Z(n40921) );
  AND U41675 ( .A(x[495]), .B(y[8102]), .Z(n40920) );
  XOR U41676 ( .A(n40921), .B(n40920), .Z(n40914) );
  XOR U41677 ( .A(n40915), .B(n40914), .Z(n40916) );
  XNOR U41678 ( .A(n40955), .B(n40954), .Z(n40970) );
  NANDN U41679 ( .A(n40779), .B(n40778), .Z(n40783) );
  NANDN U41680 ( .A(n40781), .B(n40780), .Z(n40782) );
  AND U41681 ( .A(n40783), .B(n40782), .Z(n40972) );
  XOR U41682 ( .A(n40973), .B(n40972), .Z(n40880) );
  NAND U41683 ( .A(n40785), .B(n40784), .Z(n40789) );
  NANDN U41684 ( .A(n40787), .B(n40786), .Z(n40788) );
  AND U41685 ( .A(n40789), .B(n40788), .Z(n40879) );
  NANDN U41686 ( .A(n40791), .B(n40790), .Z(n40795) );
  NAND U41687 ( .A(n40793), .B(n40792), .Z(n40794) );
  AND U41688 ( .A(n40795), .B(n40794), .Z(n40979) );
  NAND U41689 ( .A(n41644), .B(n40796), .Z(n40800) );
  NAND U41690 ( .A(n40798), .B(n40797), .Z(n40799) );
  NAND U41691 ( .A(n40800), .B(n40799), .Z(n40886) );
  NAND U41692 ( .A(n40801), .B(n42186), .Z(n40805) );
  NAND U41693 ( .A(n40803), .B(n40802), .Z(n40804) );
  NAND U41694 ( .A(n40805), .B(n40804), .Z(n40967) );
  AND U41695 ( .A(y[8098]), .B(x[499]), .Z(n40807) );
  NAND U41696 ( .A(y[8106]), .B(x[491]), .Z(n40806) );
  XNOR U41697 ( .A(n40807), .B(n40806), .Z(n40905) );
  AND U41698 ( .A(x[500]), .B(y[8097]), .Z(n40935) );
  XOR U41699 ( .A(o[437]), .B(n40935), .Z(n40904) );
  XOR U41700 ( .A(n40905), .B(n40904), .Z(n40965) );
  AND U41701 ( .A(y[8099]), .B(x[498]), .Z(n40809) );
  NAND U41702 ( .A(y[8107]), .B(x[490]), .Z(n40808) );
  XNOR U41703 ( .A(n40809), .B(n40808), .Z(n40943) );
  AND U41704 ( .A(x[481]), .B(y[8116]), .Z(n40944) );
  XOR U41705 ( .A(n40943), .B(n40944), .Z(n40964) );
  XOR U41706 ( .A(n40965), .B(n40964), .Z(n40966) );
  XOR U41707 ( .A(n40967), .B(n40966), .Z(n40885) );
  XOR U41708 ( .A(n40886), .B(n40885), .Z(n40888) );
  AND U41709 ( .A(x[487]), .B(y[8110]), .Z(n41156) );
  AND U41710 ( .A(y[8111]), .B(x[486]), .Z(n40811) );
  NAND U41711 ( .A(y[8103]), .B(x[494]), .Z(n40810) );
  XNOR U41712 ( .A(n40811), .B(n40810), .Z(n40947) );
  XOR U41713 ( .A(n41156), .B(n40947), .Z(n40894) );
  AND U41714 ( .A(x[489]), .B(y[8108]), .Z(n40892) );
  NAND U41715 ( .A(x[488]), .B(y[8109]), .Z(n40891) );
  AND U41716 ( .A(y[8105]), .B(x[492]), .Z(n40813) );
  NAND U41717 ( .A(y[8100]), .B(x[497]), .Z(n40812) );
  XNOR U41718 ( .A(n40813), .B(n40812), .Z(n40897) );
  AND U41719 ( .A(x[482]), .B(y[8115]), .Z(n40898) );
  XOR U41720 ( .A(n40897), .B(n40898), .Z(n40909) );
  AND U41721 ( .A(y[8104]), .B(x[493]), .Z(n40815) );
  NAND U41722 ( .A(y[8114]), .B(x[483]), .Z(n40814) );
  XNOR U41723 ( .A(n40815), .B(n40814), .Z(n40931) );
  AND U41724 ( .A(x[484]), .B(y[8113]), .Z(n40932) );
  XOR U41725 ( .A(n40931), .B(n40932), .Z(n40908) );
  XOR U41726 ( .A(n40909), .B(n40908), .Z(n40911) );
  XOR U41727 ( .A(n40910), .B(n40911), .Z(n40961) );
  NAND U41728 ( .A(n40923), .B(n40816), .Z(n40820) );
  NAND U41729 ( .A(n40818), .B(n40817), .Z(n40819) );
  NAND U41730 ( .A(n40820), .B(n40819), .Z(n40959) );
  NAND U41731 ( .A(n40822), .B(n40821), .Z(n40826) );
  NAND U41732 ( .A(n40824), .B(n40823), .Z(n40825) );
  NAND U41733 ( .A(n40826), .B(n40825), .Z(n40958) );
  XOR U41734 ( .A(n40959), .B(n40958), .Z(n40960) );
  XOR U41735 ( .A(n40961), .B(n40960), .Z(n40887) );
  XOR U41736 ( .A(n40888), .B(n40887), .Z(n40977) );
  NANDN U41737 ( .A(n40828), .B(n40827), .Z(n40832) );
  NAND U41738 ( .A(n40830), .B(n40829), .Z(n40831) );
  NAND U41739 ( .A(n40832), .B(n40831), .Z(n40984) );
  NAND U41740 ( .A(n40834), .B(n40833), .Z(n40838) );
  NANDN U41741 ( .A(n40836), .B(n40835), .Z(n40837) );
  NAND U41742 ( .A(n40838), .B(n40837), .Z(n40983) );
  NAND U41743 ( .A(n40840), .B(n40839), .Z(n40844) );
  NANDN U41744 ( .A(n40842), .B(n40841), .Z(n40843) );
  NAND U41745 ( .A(n40844), .B(n40843), .Z(n40982) );
  XOR U41746 ( .A(n40983), .B(n40982), .Z(n40985) );
  XOR U41747 ( .A(n40984), .B(n40985), .Z(n40976) );
  XOR U41748 ( .A(n40977), .B(n40976), .Z(n40978) );
  NANDN U41749 ( .A(n40846), .B(n40845), .Z(n40850) );
  NANDN U41750 ( .A(n40848), .B(n40847), .Z(n40849) );
  NAND U41751 ( .A(n40850), .B(n40849), .Z(n40873) );
  XOR U41752 ( .A(n40874), .B(n40873), .Z(n40876) );
  XNOR U41753 ( .A(n40875), .B(n40876), .Z(n40997) );
  NAND U41754 ( .A(n40852), .B(n40851), .Z(n40856) );
  NANDN U41755 ( .A(n40854), .B(n40853), .Z(n40855) );
  AND U41756 ( .A(n40856), .B(n40855), .Z(n40996) );
  NANDN U41757 ( .A(n40858), .B(n40857), .Z(n40862) );
  NAND U41758 ( .A(n40860), .B(n40859), .Z(n40861) );
  AND U41759 ( .A(n40862), .B(n40861), .Z(n40995) );
  XNOR U41760 ( .A(n40997), .B(n40998), .Z(n40991) );
  NAND U41761 ( .A(n40867), .B(n40866), .Z(n40871) );
  NANDN U41762 ( .A(n40869), .B(n40868), .Z(n40870) );
  AND U41763 ( .A(n40871), .B(n40870), .Z(n40989) );
  IV U41764 ( .A(n40989), .Z(n40988) );
  XOR U41765 ( .A(n40990), .B(n40988), .Z(n40872) );
  XNOR U41766 ( .A(n40991), .B(n40872), .Z(N886) );
  NAND U41767 ( .A(n40874), .B(n40873), .Z(n40878) );
  NAND U41768 ( .A(n40876), .B(n40875), .Z(n40877) );
  AND U41769 ( .A(n40878), .B(n40877), .Z(n41005) );
  NANDN U41770 ( .A(n40880), .B(n40879), .Z(n40884) );
  NANDN U41771 ( .A(n40882), .B(n40881), .Z(n40883) );
  AND U41772 ( .A(n40884), .B(n40883), .Z(n41003) );
  NAND U41773 ( .A(n40886), .B(n40885), .Z(n40890) );
  NAND U41774 ( .A(n40888), .B(n40887), .Z(n40889) );
  NAND U41775 ( .A(n40890), .B(n40889), .Z(n41132) );
  NANDN U41776 ( .A(n40892), .B(n40891), .Z(n40896) );
  NANDN U41777 ( .A(n40894), .B(n40893), .Z(n40895) );
  NAND U41778 ( .A(n40896), .B(n40895), .Z(n41126) );
  NAND U41779 ( .A(n41077), .B(n41653), .Z(n40900) );
  NAND U41780 ( .A(n40898), .B(n40897), .Z(n40899) );
  NAND U41781 ( .A(n40900), .B(n40899), .Z(n41053) );
  AND U41782 ( .A(x[485]), .B(y[8113]), .Z(n41099) );
  AND U41783 ( .A(x[497]), .B(y[8101]), .Z(n41100) );
  XOR U41784 ( .A(n41099), .B(n41100), .Z(n41101) );
  AND U41785 ( .A(x[496]), .B(y[8102]), .Z(n41102) );
  XOR U41786 ( .A(n41101), .B(n41102), .Z(n41052) );
  AND U41787 ( .A(y[8100]), .B(x[498]), .Z(n40902) );
  NAND U41788 ( .A(y[8106]), .B(x[492]), .Z(n40901) );
  XNOR U41789 ( .A(n40902), .B(n40901), .Z(n41078) );
  AND U41790 ( .A(x[484]), .B(y[8114]), .Z(n41079) );
  XOR U41791 ( .A(n41078), .B(n41079), .Z(n41051) );
  XOR U41792 ( .A(n41052), .B(n41051), .Z(n41054) );
  XNOR U41793 ( .A(n41053), .B(n41054), .Z(n41123) );
  AND U41794 ( .A(x[499]), .B(y[8106]), .Z(n42071) );
  NAND U41795 ( .A(n42071), .B(n40903), .Z(n40907) );
  NAND U41796 ( .A(n40905), .B(n40904), .Z(n40906) );
  AND U41797 ( .A(n40907), .B(n40906), .Z(n41124) );
  XOR U41798 ( .A(n41123), .B(n41124), .Z(n41125) );
  XNOR U41799 ( .A(n41126), .B(n41125), .Z(n41129) );
  NAND U41800 ( .A(n40909), .B(n40908), .Z(n40913) );
  NAND U41801 ( .A(n40911), .B(n40910), .Z(n40912) );
  NAND U41802 ( .A(n40913), .B(n40912), .Z(n41112) );
  NAND U41803 ( .A(n40915), .B(n40914), .Z(n40919) );
  NANDN U41804 ( .A(n40917), .B(n40916), .Z(n40918) );
  NAND U41805 ( .A(n40919), .B(n40918), .Z(n41111) );
  XOR U41806 ( .A(n41112), .B(n41111), .Z(n41114) );
  AND U41807 ( .A(n40921), .B(n40920), .Z(n40925) );
  NAND U41808 ( .A(n40923), .B(n40922), .Z(n40924) );
  NANDN U41809 ( .A(n40925), .B(n40924), .Z(n41074) );
  AND U41810 ( .A(y[8105]), .B(x[493]), .Z(n40927) );
  NAND U41811 ( .A(y[8098]), .B(x[500]), .Z(n40926) );
  XNOR U41812 ( .A(n40927), .B(n40926), .Z(n41095) );
  AND U41813 ( .A(x[482]), .B(y[8116]), .Z(n41096) );
  XOR U41814 ( .A(n41095), .B(n41096), .Z(n41072) );
  AND U41815 ( .A(y[8112]), .B(x[486]), .Z(n40929) );
  NAND U41816 ( .A(y[8103]), .B(x[495]), .Z(n40928) );
  XNOR U41817 ( .A(n40929), .B(n40928), .Z(n41107) );
  XOR U41818 ( .A(n41072), .B(n41071), .Z(n41073) );
  XOR U41819 ( .A(n41074), .B(n41073), .Z(n41118) );
  AND U41820 ( .A(x[493]), .B(y[8114]), .Z(n42409) );
  NANDN U41821 ( .A(n40930), .B(n42409), .Z(n40934) );
  NAND U41822 ( .A(n40932), .B(n40931), .Z(n40933) );
  NAND U41823 ( .A(n40934), .B(n40933), .Z(n41042) );
  AND U41824 ( .A(x[481]), .B(y[8117]), .Z(n41065) );
  XOR U41825 ( .A(n41066), .B(n41065), .Z(n41064) );
  AND U41826 ( .A(o[437]), .B(n40935), .Z(n41063) );
  XOR U41827 ( .A(n41064), .B(n41063), .Z(n41040) );
  AND U41828 ( .A(x[494]), .B(y[8104]), .Z(n41057) );
  AND U41829 ( .A(x[483]), .B(y[8115]), .Z(n41058) );
  XOR U41830 ( .A(n41057), .B(n41058), .Z(n41059) );
  AND U41831 ( .A(x[499]), .B(y[8099]), .Z(n41060) );
  XOR U41832 ( .A(n41059), .B(n41060), .Z(n41039) );
  XOR U41833 ( .A(n41040), .B(n41039), .Z(n41041) );
  XOR U41834 ( .A(n41042), .B(n41041), .Z(n41117) );
  XOR U41835 ( .A(n41118), .B(n41117), .Z(n41120) );
  NAND U41836 ( .A(n40937), .B(n40936), .Z(n40941) );
  NAND U41837 ( .A(n40939), .B(n40938), .Z(n40940) );
  NAND U41838 ( .A(n40941), .B(n40940), .Z(n41034) );
  AND U41839 ( .A(x[498]), .B(y[8107]), .Z(n42073) );
  NAND U41840 ( .A(n42073), .B(n40942), .Z(n40946) );
  NAND U41841 ( .A(n40944), .B(n40943), .Z(n40945) );
  NAND U41842 ( .A(n40946), .B(n40945), .Z(n41033) );
  XOR U41843 ( .A(n41034), .B(n41033), .Z(n41036) );
  AND U41844 ( .A(x[494]), .B(y[8111]), .Z(n42113) );
  NAND U41845 ( .A(n41106), .B(n42113), .Z(n40949) );
  NAND U41846 ( .A(n41156), .B(n40947), .Z(n40948) );
  NAND U41847 ( .A(n40949), .B(n40948), .Z(n41048) );
  AND U41848 ( .A(x[480]), .B(y[8118]), .Z(n41082) );
  AND U41849 ( .A(x[502]), .B(y[8096]), .Z(n41083) );
  XOR U41850 ( .A(n41082), .B(n41083), .Z(n41085) );
  AND U41851 ( .A(x[501]), .B(y[8097]), .Z(n41105) );
  XOR U41852 ( .A(o[438]), .B(n41105), .Z(n41084) );
  XOR U41853 ( .A(n41085), .B(n41084), .Z(n41046) );
  AND U41854 ( .A(y[8111]), .B(x[487]), .Z(n40951) );
  NAND U41855 ( .A(y[8110]), .B(x[488]), .Z(n40950) );
  XNOR U41856 ( .A(n40951), .B(n40950), .Z(n41088) );
  XOR U41857 ( .A(n41046), .B(n41045), .Z(n41047) );
  XOR U41858 ( .A(n41048), .B(n41047), .Z(n41035) );
  XOR U41859 ( .A(n41036), .B(n41035), .Z(n41119) );
  XOR U41860 ( .A(n41120), .B(n41119), .Z(n41113) );
  XOR U41861 ( .A(n41114), .B(n41113), .Z(n41130) );
  XOR U41862 ( .A(n41129), .B(n41130), .Z(n41131) );
  XOR U41863 ( .A(n41132), .B(n41131), .Z(n41024) );
  NAND U41864 ( .A(n40953), .B(n40952), .Z(n40957) );
  NAND U41865 ( .A(n40955), .B(n40954), .Z(n40956) );
  NAND U41866 ( .A(n40957), .B(n40956), .Z(n41030) );
  NAND U41867 ( .A(n40959), .B(n40958), .Z(n40963) );
  NAND U41868 ( .A(n40961), .B(n40960), .Z(n40962) );
  NAND U41869 ( .A(n40963), .B(n40962), .Z(n41028) );
  NAND U41870 ( .A(n40965), .B(n40964), .Z(n40969) );
  NAND U41871 ( .A(n40967), .B(n40966), .Z(n40968) );
  NAND U41872 ( .A(n40969), .B(n40968), .Z(n41027) );
  XOR U41873 ( .A(n41028), .B(n41027), .Z(n41029) );
  XOR U41874 ( .A(n41030), .B(n41029), .Z(n41022) );
  NANDN U41875 ( .A(n40971), .B(n40970), .Z(n40975) );
  NAND U41876 ( .A(n40973), .B(n40972), .Z(n40974) );
  NAND U41877 ( .A(n40975), .B(n40974), .Z(n41021) );
  NAND U41878 ( .A(n40977), .B(n40976), .Z(n40981) );
  NANDN U41879 ( .A(n40979), .B(n40978), .Z(n40980) );
  NAND U41880 ( .A(n40981), .B(n40980), .Z(n41016) );
  NAND U41881 ( .A(n40983), .B(n40982), .Z(n40987) );
  NAND U41882 ( .A(n40985), .B(n40984), .Z(n40986) );
  NAND U41883 ( .A(n40987), .B(n40986), .Z(n41015) );
  XOR U41884 ( .A(n41016), .B(n41015), .Z(n41017) );
  XNOR U41885 ( .A(n41005), .B(n41004), .Z(n41011) );
  OR U41886 ( .A(n40990), .B(n40988), .Z(n40994) );
  ANDN U41887 ( .B(n40990), .A(n40989), .Z(n40992) );
  OR U41888 ( .A(n40992), .B(n40991), .Z(n40993) );
  AND U41889 ( .A(n40994), .B(n40993), .Z(n41010) );
  NANDN U41890 ( .A(n40996), .B(n40995), .Z(n41000) );
  NAND U41891 ( .A(n40998), .B(n40997), .Z(n40999) );
  NAND U41892 ( .A(n41000), .B(n40999), .Z(n41009) );
  IV U41893 ( .A(n41009), .Z(n41008) );
  XOR U41894 ( .A(n41010), .B(n41008), .Z(n41001) );
  XNOR U41895 ( .A(n41011), .B(n41001), .Z(N887) );
  NANDN U41896 ( .A(n41003), .B(n41002), .Z(n41007) );
  NAND U41897 ( .A(n41005), .B(n41004), .Z(n41006) );
  NAND U41898 ( .A(n41007), .B(n41006), .Z(n41266) );
  IV U41899 ( .A(n41266), .Z(n41265) );
  OR U41900 ( .A(n41010), .B(n41008), .Z(n41014) );
  ANDN U41901 ( .B(n41010), .A(n41009), .Z(n41012) );
  OR U41902 ( .A(n41012), .B(n41011), .Z(n41013) );
  AND U41903 ( .A(n41014), .B(n41013), .Z(n41267) );
  NAND U41904 ( .A(n41016), .B(n41015), .Z(n41020) );
  NANDN U41905 ( .A(n41018), .B(n41017), .Z(n41019) );
  AND U41906 ( .A(n41020), .B(n41019), .Z(n41274) );
  NANDN U41907 ( .A(n41022), .B(n41021), .Z(n41026) );
  NANDN U41908 ( .A(n41024), .B(n41023), .Z(n41025) );
  NAND U41909 ( .A(n41026), .B(n41025), .Z(n41272) );
  NAND U41910 ( .A(n41028), .B(n41027), .Z(n41032) );
  NAND U41911 ( .A(n41030), .B(n41029), .Z(n41031) );
  NAND U41912 ( .A(n41032), .B(n41031), .Z(n41250) );
  NAND U41913 ( .A(n41034), .B(n41033), .Z(n41038) );
  NAND U41914 ( .A(n41036), .B(n41035), .Z(n41037) );
  NAND U41915 ( .A(n41038), .B(n41037), .Z(n41244) );
  NAND U41916 ( .A(n41040), .B(n41039), .Z(n41044) );
  NAND U41917 ( .A(n41042), .B(n41041), .Z(n41043) );
  NAND U41918 ( .A(n41044), .B(n41043), .Z(n41242) );
  NAND U41919 ( .A(n41046), .B(n41045), .Z(n41050) );
  NAND U41920 ( .A(n41048), .B(n41047), .Z(n41049) );
  NAND U41921 ( .A(n41050), .B(n41049), .Z(n41241) );
  XOR U41922 ( .A(n41242), .B(n41241), .Z(n41243) );
  XOR U41923 ( .A(n41244), .B(n41243), .Z(n41262) );
  NAND U41924 ( .A(n41052), .B(n41051), .Z(n41056) );
  NAND U41925 ( .A(n41054), .B(n41053), .Z(n41055) );
  AND U41926 ( .A(n41056), .B(n41055), .Z(n41260) );
  NAND U41927 ( .A(n41058), .B(n41057), .Z(n41062) );
  NAND U41928 ( .A(n41060), .B(n41059), .Z(n41061) );
  NAND U41929 ( .A(n41062), .B(n41061), .Z(n41190) );
  AND U41930 ( .A(n41064), .B(n41063), .Z(n41068) );
  NAND U41931 ( .A(n41066), .B(n41065), .Z(n41067) );
  NANDN U41932 ( .A(n41068), .B(n41067), .Z(n41189) );
  XOR U41933 ( .A(n41190), .B(n41189), .Z(n41192) );
  AND U41934 ( .A(y[8112]), .B(x[487]), .Z(n41070) );
  NAND U41935 ( .A(y[8110]), .B(x[489]), .Z(n41069) );
  XNOR U41936 ( .A(n41070), .B(n41069), .Z(n41157) );
  NAND U41937 ( .A(x[490]), .B(y[8109]), .Z(n41196) );
  AND U41938 ( .A(x[486]), .B(y[8113]), .Z(n41148) );
  NAND U41939 ( .A(x[495]), .B(y[8104]), .Z(n41149) );
  XNOR U41940 ( .A(n41148), .B(n41149), .Z(n41150) );
  NAND U41941 ( .A(x[491]), .B(y[8108]), .Z(n41151) );
  XOR U41942 ( .A(n41150), .B(n41151), .Z(n41198) );
  XOR U41943 ( .A(n41192), .B(n41191), .Z(n41259) );
  XOR U41944 ( .A(n41262), .B(n41261), .Z(n41248) );
  NAND U41945 ( .A(n41072), .B(n41071), .Z(n41076) );
  NAND U41946 ( .A(n41074), .B(n41073), .Z(n41075) );
  NAND U41947 ( .A(n41076), .B(n41075), .Z(n41184) );
  AND U41948 ( .A(x[498]), .B(y[8106]), .Z(n41945) );
  NAND U41949 ( .A(n41945), .B(n41077), .Z(n41081) );
  NAND U41950 ( .A(n41079), .B(n41078), .Z(n41080) );
  NAND U41951 ( .A(n41081), .B(n41080), .Z(n41218) );
  NAND U41952 ( .A(n41083), .B(n41082), .Z(n41087) );
  NAND U41953 ( .A(n41085), .B(n41084), .Z(n41086) );
  NAND U41954 ( .A(n41087), .B(n41086), .Z(n41217) );
  XOR U41955 ( .A(n41218), .B(n41217), .Z(n41219) );
  NANDN U41956 ( .A(n41158), .B(n41156), .Z(n41091) );
  NANDN U41957 ( .A(n41089), .B(n41088), .Z(n41090) );
  NAND U41958 ( .A(n41091), .B(n41090), .Z(n41231) );
  AND U41959 ( .A(x[480]), .B(y[8119]), .Z(n41167) );
  AND U41960 ( .A(x[503]), .B(y[8096]), .Z(n41168) );
  XOR U41961 ( .A(n41167), .B(n41168), .Z(n41169) );
  NAND U41962 ( .A(x[502]), .B(y[8097]), .Z(n41147) );
  XNOR U41963 ( .A(o[439]), .B(n41147), .Z(n41170) );
  XOR U41964 ( .A(n41169), .B(n41170), .Z(n41230) );
  NAND U41965 ( .A(y[8099]), .B(x[500]), .Z(n41092) );
  XNOR U41966 ( .A(n41093), .B(n41092), .Z(n41143) );
  NAND U41967 ( .A(x[499]), .B(y[8100]), .Z(n41144) );
  XNOR U41968 ( .A(n41143), .B(n41144), .Z(n41229) );
  XOR U41969 ( .A(n41230), .B(n41229), .Z(n41232) );
  XNOR U41970 ( .A(n41231), .B(n41232), .Z(n41220) );
  XOR U41971 ( .A(n41184), .B(n41183), .Z(n41186) );
  AND U41972 ( .A(x[500]), .B(y[8105]), .Z(n42124) );
  AND U41973 ( .A(x[493]), .B(y[8098]), .Z(n41094) );
  NAND U41974 ( .A(n42124), .B(n41094), .Z(n41098) );
  NAND U41975 ( .A(n41096), .B(n41095), .Z(n41097) );
  NAND U41976 ( .A(n41098), .B(n41097), .Z(n41178) );
  NAND U41977 ( .A(n41100), .B(n41099), .Z(n41104) );
  NAND U41978 ( .A(n41102), .B(n41101), .Z(n41103) );
  NAND U41979 ( .A(n41104), .B(n41103), .Z(n41237) );
  AND U41980 ( .A(x[493]), .B(y[8106]), .Z(n41212) );
  AND U41981 ( .A(x[482]), .B(y[8117]), .Z(n41211) );
  XOR U41982 ( .A(n41212), .B(n41211), .Z(n41214) );
  AND U41983 ( .A(x[501]), .B(y[8098]), .Z(n41213) );
  XOR U41984 ( .A(n41214), .B(n41213), .Z(n41236) );
  AND U41985 ( .A(o[438]), .B(n41105), .Z(n41164) );
  AND U41986 ( .A(x[492]), .B(y[8107]), .Z(n41162) );
  AND U41987 ( .A(x[481]), .B(y[8118]), .Z(n41161) );
  XOR U41988 ( .A(n41162), .B(n41161), .Z(n41163) );
  XOR U41989 ( .A(n41164), .B(n41163), .Z(n41235) );
  XOR U41990 ( .A(n41236), .B(n41235), .Z(n41238) );
  XOR U41991 ( .A(n41237), .B(n41238), .Z(n41177) );
  XOR U41992 ( .A(n41178), .B(n41177), .Z(n41180) );
  AND U41993 ( .A(x[495]), .B(y[8112]), .Z(n42286) );
  NAND U41994 ( .A(n42286), .B(n41106), .Z(n41110) );
  NANDN U41995 ( .A(n41108), .B(n41107), .Z(n41109) );
  NAND U41996 ( .A(n41110), .B(n41109), .Z(n41225) );
  AND U41997 ( .A(x[494]), .B(y[8105]), .Z(n41206) );
  AND U41998 ( .A(x[483]), .B(y[8116]), .Z(n41205) );
  XOR U41999 ( .A(n41206), .B(n41205), .Z(n41208) );
  AND U42000 ( .A(x[484]), .B(y[8115]), .Z(n41207) );
  XOR U42001 ( .A(n41208), .B(n41207), .Z(n41224) );
  AND U42002 ( .A(x[485]), .B(y[8114]), .Z(n41202) );
  AND U42003 ( .A(x[498]), .B(y[8101]), .Z(n41201) );
  XOR U42004 ( .A(n41202), .B(n41201), .Z(n41204) );
  AND U42005 ( .A(x[497]), .B(y[8102]), .Z(n41203) );
  XOR U42006 ( .A(n41204), .B(n41203), .Z(n41223) );
  XOR U42007 ( .A(n41224), .B(n41223), .Z(n41226) );
  XOR U42008 ( .A(n41225), .B(n41226), .Z(n41179) );
  XOR U42009 ( .A(n41180), .B(n41179), .Z(n41185) );
  XOR U42010 ( .A(n41186), .B(n41185), .Z(n41247) );
  XOR U42011 ( .A(n41248), .B(n41247), .Z(n41249) );
  XNOR U42012 ( .A(n41250), .B(n41249), .Z(n41138) );
  NAND U42013 ( .A(n41112), .B(n41111), .Z(n41116) );
  NAND U42014 ( .A(n41114), .B(n41113), .Z(n41115) );
  NAND U42015 ( .A(n41116), .B(n41115), .Z(n41256) );
  NAND U42016 ( .A(n41118), .B(n41117), .Z(n41122) );
  NAND U42017 ( .A(n41120), .B(n41119), .Z(n41121) );
  NAND U42018 ( .A(n41122), .B(n41121), .Z(n41254) );
  NAND U42019 ( .A(n41124), .B(n41123), .Z(n41128) );
  NAND U42020 ( .A(n41126), .B(n41125), .Z(n41127) );
  AND U42021 ( .A(n41128), .B(n41127), .Z(n41253) );
  XOR U42022 ( .A(n41254), .B(n41253), .Z(n41255) );
  XNOR U42023 ( .A(n41256), .B(n41255), .Z(n41136) );
  NAND U42024 ( .A(n41130), .B(n41129), .Z(n41134) );
  NAND U42025 ( .A(n41132), .B(n41131), .Z(n41133) );
  AND U42026 ( .A(n41134), .B(n41133), .Z(n41137) );
  XOR U42027 ( .A(n41136), .B(n41137), .Z(n41139) );
  XNOR U42028 ( .A(n41138), .B(n41139), .Z(n41273) );
  XNOR U42029 ( .A(n41274), .B(n41275), .Z(n41268) );
  XNOR U42030 ( .A(n41267), .B(n41268), .Z(n41135) );
  XOR U42031 ( .A(n41265), .B(n41135), .Z(N888) );
  NAND U42032 ( .A(n41137), .B(n41136), .Z(n41141) );
  NAND U42033 ( .A(n41139), .B(n41138), .Z(n41140) );
  AND U42034 ( .A(n41141), .B(n41140), .Z(n41414) );
  AND U42035 ( .A(x[500]), .B(y[8103]), .Z(n41142) );
  NAND U42036 ( .A(n41375), .B(n41142), .Z(n41146) );
  NANDN U42037 ( .A(n41144), .B(n41143), .Z(n41145) );
  NAND U42038 ( .A(n41146), .B(n41145), .Z(n41396) );
  AND U42039 ( .A(x[502]), .B(y[8098]), .Z(n41307) );
  XOR U42040 ( .A(n41308), .B(n41307), .Z(n41310) );
  NAND U42041 ( .A(x[482]), .B(y[8118]), .Z(n41309) );
  XNOR U42042 ( .A(n41310), .B(n41309), .Z(n41395) );
  ANDN U42043 ( .B(o[439]), .A(n41147), .Z(n41314) );
  AND U42044 ( .A(x[481]), .B(y[8119]), .Z(n41315) );
  XOR U42045 ( .A(n41316), .B(n41315), .Z(n41313) );
  XOR U42046 ( .A(n41314), .B(n41313), .Z(n41394) );
  XOR U42047 ( .A(n41395), .B(n41394), .Z(n41397) );
  XOR U42048 ( .A(n41396), .B(n41397), .Z(n41346) );
  NANDN U42049 ( .A(n41149), .B(n41148), .Z(n41153) );
  NANDN U42050 ( .A(n41151), .B(n41150), .Z(n41152) );
  NAND U42051 ( .A(n41153), .B(n41152), .Z(n41392) );
  AND U42052 ( .A(y[8104]), .B(x[496]), .Z(n41155) );
  NAND U42053 ( .A(y[8099]), .B(x[501]), .Z(n41154) );
  XNOR U42054 ( .A(n41155), .B(n41154), .Z(n41376) );
  NAND U42055 ( .A(x[485]), .B(y[8115]), .Z(n41377) );
  XNOR U42056 ( .A(n41376), .B(n41377), .Z(n41391) );
  AND U42057 ( .A(x[486]), .B(y[8114]), .Z(n41692) );
  NAND U42058 ( .A(x[500]), .B(y[8100]), .Z(n41511) );
  XNOR U42059 ( .A(n41692), .B(n41511), .Z(n41383) );
  AND U42060 ( .A(x[499]), .B(y[8101]), .Z(n41382) );
  XOR U42061 ( .A(n41383), .B(n41382), .Z(n41390) );
  XOR U42062 ( .A(n41391), .B(n41390), .Z(n41393) );
  XOR U42063 ( .A(n41392), .B(n41393), .Z(n41372) );
  NAND U42064 ( .A(n41443), .B(n41156), .Z(n41160) );
  NANDN U42065 ( .A(n41158), .B(n41157), .Z(n41159) );
  NAND U42066 ( .A(n41160), .B(n41159), .Z(n41370) );
  NAND U42067 ( .A(n41162), .B(n41161), .Z(n41166) );
  NAND U42068 ( .A(n41164), .B(n41163), .Z(n41165) );
  NAND U42069 ( .A(n41166), .B(n41165), .Z(n41369) );
  XOR U42070 ( .A(n41370), .B(n41369), .Z(n41371) );
  XOR U42071 ( .A(n41372), .B(n41371), .Z(n41345) );
  XOR U42072 ( .A(n41346), .B(n41345), .Z(n41348) );
  NAND U42073 ( .A(n41168), .B(n41167), .Z(n41172) );
  NAND U42074 ( .A(n41170), .B(n41169), .Z(n41171) );
  NAND U42075 ( .A(n41172), .B(n41171), .Z(n41339) );
  AND U42076 ( .A(x[483]), .B(y[8117]), .Z(n41327) );
  XOR U42077 ( .A(n41328), .B(n41327), .Z(n41330) );
  NAND U42078 ( .A(x[484]), .B(y[8116]), .Z(n41329) );
  XNOR U42079 ( .A(n41330), .B(n41329), .Z(n41340) );
  XOR U42080 ( .A(n41339), .B(n41340), .Z(n41342) );
  AND U42081 ( .A(y[8111]), .B(x[489]), .Z(n41174) );
  NAND U42082 ( .A(y[8110]), .B(x[490]), .Z(n41173) );
  XNOR U42083 ( .A(n41174), .B(n41173), .Z(n41299) );
  AND U42084 ( .A(y[8106]), .B(x[494]), .Z(n41176) );
  NAND U42085 ( .A(y[8112]), .B(x[488]), .Z(n41175) );
  XNOR U42086 ( .A(n41176), .B(n41175), .Z(n41303) );
  NAND U42087 ( .A(x[491]), .B(y[8109]), .Z(n41304) );
  XNOR U42088 ( .A(n41303), .B(n41304), .Z(n41298) );
  XOR U42089 ( .A(n41299), .B(n41298), .Z(n41341) );
  XOR U42090 ( .A(n41342), .B(n41341), .Z(n41347) );
  XOR U42091 ( .A(n41348), .B(n41347), .Z(n41292) );
  NAND U42092 ( .A(n41178), .B(n41177), .Z(n41182) );
  NAND U42093 ( .A(n41180), .B(n41179), .Z(n41181) );
  AND U42094 ( .A(n41182), .B(n41181), .Z(n41291) );
  NAND U42095 ( .A(n41184), .B(n41183), .Z(n41188) );
  NAND U42096 ( .A(n41186), .B(n41185), .Z(n41187) );
  NAND U42097 ( .A(n41188), .B(n41187), .Z(n41294) );
  NAND U42098 ( .A(n41190), .B(n41189), .Z(n41194) );
  NAND U42099 ( .A(n41192), .B(n41191), .Z(n41193) );
  AND U42100 ( .A(n41194), .B(n41193), .Z(n41354) );
  NANDN U42101 ( .A(n41196), .B(n41195), .Z(n41200) );
  NANDN U42102 ( .A(n41198), .B(n41197), .Z(n41199) );
  AND U42103 ( .A(n41200), .B(n41199), .Z(n41352) );
  AND U42104 ( .A(x[480]), .B(y[8120]), .Z(n41333) );
  NAND U42105 ( .A(x[504]), .B(y[8096]), .Z(n41334) );
  XNOR U42106 ( .A(n41333), .B(n41334), .Z(n41335) );
  NAND U42107 ( .A(x[503]), .B(y[8097]), .Z(n41326) );
  XOR U42108 ( .A(o[440]), .B(n41326), .Z(n41336) );
  XNOR U42109 ( .A(n41335), .B(n41336), .Z(n41387) );
  AND U42110 ( .A(x[487]), .B(y[8113]), .Z(n41319) );
  NAND U42111 ( .A(x[498]), .B(y[8102]), .Z(n41320) );
  XNOR U42112 ( .A(n41319), .B(n41320), .Z(n41322) );
  AND U42113 ( .A(x[497]), .B(y[8103]), .Z(n41321) );
  XOR U42114 ( .A(n41322), .B(n41321), .Z(n41386) );
  XOR U42115 ( .A(n41387), .B(n41386), .Z(n41389) );
  XOR U42116 ( .A(n41388), .B(n41389), .Z(n41365) );
  NAND U42117 ( .A(n41206), .B(n41205), .Z(n41210) );
  NAND U42118 ( .A(n41208), .B(n41207), .Z(n41209) );
  NAND U42119 ( .A(n41210), .B(n41209), .Z(n41364) );
  NAND U42120 ( .A(n41212), .B(n41211), .Z(n41216) );
  NAND U42121 ( .A(n41214), .B(n41213), .Z(n41215) );
  NAND U42122 ( .A(n41216), .B(n41215), .Z(n41363) );
  XNOR U42123 ( .A(n41364), .B(n41363), .Z(n41366) );
  NAND U42124 ( .A(n41218), .B(n41217), .Z(n41222) );
  NANDN U42125 ( .A(n41220), .B(n41219), .Z(n41221) );
  AND U42126 ( .A(n41222), .B(n41221), .Z(n41401) );
  NAND U42127 ( .A(n41224), .B(n41223), .Z(n41228) );
  NAND U42128 ( .A(n41226), .B(n41225), .Z(n41227) );
  AND U42129 ( .A(n41228), .B(n41227), .Z(n41399) );
  NAND U42130 ( .A(n41230), .B(n41229), .Z(n41234) );
  NAND U42131 ( .A(n41232), .B(n41231), .Z(n41233) );
  AND U42132 ( .A(n41234), .B(n41233), .Z(n41398) );
  XOR U42133 ( .A(n41399), .B(n41398), .Z(n41400) );
  XOR U42134 ( .A(n41401), .B(n41400), .Z(n41357) );
  NAND U42135 ( .A(n41236), .B(n41235), .Z(n41240) );
  NAND U42136 ( .A(n41238), .B(n41237), .Z(n41239) );
  NAND U42137 ( .A(n41240), .B(n41239), .Z(n41358) );
  XOR U42138 ( .A(n41359), .B(n41360), .Z(n41285) );
  NAND U42139 ( .A(n41242), .B(n41241), .Z(n41246) );
  NAND U42140 ( .A(n41244), .B(n41243), .Z(n41245) );
  NAND U42141 ( .A(n41246), .B(n41245), .Z(n41286) );
  XNOR U42142 ( .A(n41288), .B(n41287), .Z(n41412) );
  NAND U42143 ( .A(n41248), .B(n41247), .Z(n41252) );
  NAND U42144 ( .A(n41250), .B(n41249), .Z(n41251) );
  AND U42145 ( .A(n41252), .B(n41251), .Z(n41282) );
  NAND U42146 ( .A(n41254), .B(n41253), .Z(n41258) );
  NAND U42147 ( .A(n41256), .B(n41255), .Z(n41257) );
  AND U42148 ( .A(n41258), .B(n41257), .Z(n41280) );
  NANDN U42149 ( .A(n41260), .B(n41259), .Z(n41264) );
  NAND U42150 ( .A(n41262), .B(n41261), .Z(n41263) );
  NAND U42151 ( .A(n41264), .B(n41263), .Z(n41279) );
  XOR U42152 ( .A(n41412), .B(n41411), .Z(n41413) );
  XNOR U42153 ( .A(n41414), .B(n41413), .Z(n41407) );
  OR U42154 ( .A(n41267), .B(n41265), .Z(n41271) );
  ANDN U42155 ( .B(n41267), .A(n41266), .Z(n41269) );
  OR U42156 ( .A(n41269), .B(n41268), .Z(n41270) );
  AND U42157 ( .A(n41271), .B(n41270), .Z(n41406) );
  NANDN U42158 ( .A(n41273), .B(n41272), .Z(n41277) );
  NANDN U42159 ( .A(n41275), .B(n41274), .Z(n41276) );
  AND U42160 ( .A(n41277), .B(n41276), .Z(n41405) );
  IV U42161 ( .A(n41405), .Z(n41404) );
  XOR U42162 ( .A(n41406), .B(n41404), .Z(n41278) );
  XNOR U42163 ( .A(n41407), .B(n41278), .Z(N889) );
  NANDN U42164 ( .A(n41280), .B(n41279), .Z(n41284) );
  NANDN U42165 ( .A(n41282), .B(n41281), .Z(n41283) );
  AND U42166 ( .A(n41284), .B(n41283), .Z(n41555) );
  NANDN U42167 ( .A(n41286), .B(n41285), .Z(n41290) );
  NAND U42168 ( .A(n41288), .B(n41287), .Z(n41289) );
  AND U42169 ( .A(n41290), .B(n41289), .Z(n41553) );
  NANDN U42170 ( .A(n41292), .B(n41291), .Z(n41296) );
  NANDN U42171 ( .A(n41294), .B(n41293), .Z(n41295) );
  NAND U42172 ( .A(n41296), .B(n41295), .Z(n41418) );
  NANDN U42173 ( .A(n41442), .B(n41297), .Z(n41301) );
  NAND U42174 ( .A(n41299), .B(n41298), .Z(n41300) );
  NAND U42175 ( .A(n41301), .B(n41300), .Z(n41464) );
  AND U42176 ( .A(x[494]), .B(y[8112]), .Z(n42415) );
  NAND U42177 ( .A(n42415), .B(n41302), .Z(n41306) );
  NANDN U42178 ( .A(n41304), .B(n41303), .Z(n41305) );
  AND U42179 ( .A(n41306), .B(n41305), .Z(n41489) );
  AND U42180 ( .A(x[491]), .B(y[8110]), .Z(n41507) );
  AND U42181 ( .A(x[492]), .B(y[8109]), .Z(n41506) );
  NAND U42182 ( .A(x[487]), .B(y[8114]), .Z(n41505) );
  XOR U42183 ( .A(n41506), .B(n41505), .Z(n41508) );
  XOR U42184 ( .A(n41507), .B(n41508), .Z(n41487) );
  NAND U42185 ( .A(x[504]), .B(y[8097]), .Z(n41504) );
  XNOR U42186 ( .A(o[441]), .B(n41504), .Z(n41474) );
  NAND U42187 ( .A(x[481]), .B(y[8120]), .Z(n41475) );
  XNOR U42188 ( .A(n41474), .B(n41475), .Z(n41476) );
  NAND U42189 ( .A(x[493]), .B(y[8108]), .Z(n41477) );
  XNOR U42190 ( .A(n41476), .B(n41477), .Z(n41486) );
  XNOR U42191 ( .A(n41487), .B(n41486), .Z(n41488) );
  XNOR U42192 ( .A(n41489), .B(n41488), .Z(n41465) );
  XOR U42193 ( .A(n41464), .B(n41465), .Z(n41467) );
  NAND U42194 ( .A(n41308), .B(n41307), .Z(n41312) );
  ANDN U42195 ( .B(n41310), .A(n41309), .Z(n41311) );
  ANDN U42196 ( .B(n41312), .A(n41311), .Z(n41453) );
  AND U42197 ( .A(n41314), .B(n41313), .Z(n41318) );
  NAND U42198 ( .A(n41316), .B(n41315), .Z(n41317) );
  NANDN U42199 ( .A(n41318), .B(n41317), .Z(n41452) );
  XNOR U42200 ( .A(n41453), .B(n41452), .Z(n41455) );
  NANDN U42201 ( .A(n41320), .B(n41319), .Z(n41324) );
  NAND U42202 ( .A(n41322), .B(n41321), .Z(n41323) );
  AND U42203 ( .A(n41324), .B(n41323), .Z(n41451) );
  AND U42204 ( .A(x[488]), .B(y[8113]), .Z(n41445) );
  XOR U42205 ( .A(n41443), .B(n41325), .Z(n41444) );
  XOR U42206 ( .A(n41445), .B(n41444), .Z(n41448) );
  ANDN U42207 ( .B(o[440]), .A(n41326), .Z(n41438) );
  AND U42208 ( .A(x[505]), .B(y[8096]), .Z(n41437) );
  NAND U42209 ( .A(x[480]), .B(y[8121]), .Z(n41436) );
  XOR U42210 ( .A(n41437), .B(n41436), .Z(n41439) );
  XNOR U42211 ( .A(n41438), .B(n41439), .Z(n41449) );
  XOR U42212 ( .A(n41448), .B(n41449), .Z(n41450) );
  XNOR U42213 ( .A(n41451), .B(n41450), .Z(n41454) );
  XOR U42214 ( .A(n41455), .B(n41454), .Z(n41466) );
  XOR U42215 ( .A(n41467), .B(n41466), .Z(n41549) );
  NAND U42216 ( .A(n41328), .B(n41327), .Z(n41332) );
  ANDN U42217 ( .B(n41330), .A(n41329), .Z(n41331) );
  ANDN U42218 ( .B(n41332), .A(n41331), .Z(n41525) );
  NANDN U42219 ( .A(n41334), .B(n41333), .Z(n41338) );
  NANDN U42220 ( .A(n41336), .B(n41335), .Z(n41337) );
  AND U42221 ( .A(n41338), .B(n41337), .Z(n41523) );
  AND U42222 ( .A(x[494]), .B(y[8107]), .Z(n41480) );
  NAND U42223 ( .A(x[482]), .B(y[8119]), .Z(n41481) );
  XNOR U42224 ( .A(n41480), .B(n41481), .Z(n41482) );
  NAND U42225 ( .A(x[483]), .B(y[8118]), .Z(n41483) );
  XNOR U42226 ( .A(n41482), .B(n41483), .Z(n41522) );
  XNOR U42227 ( .A(n41523), .B(n41522), .Z(n41524) );
  XOR U42228 ( .A(n41525), .B(n41524), .Z(n41546) );
  NAND U42229 ( .A(n41340), .B(n41339), .Z(n41344) );
  NAND U42230 ( .A(n41342), .B(n41341), .Z(n41343) );
  AND U42231 ( .A(n41344), .B(n41343), .Z(n41547) );
  XOR U42232 ( .A(n41546), .B(n41547), .Z(n41548) );
  NAND U42233 ( .A(n41346), .B(n41345), .Z(n41350) );
  NAND U42234 ( .A(n41348), .B(n41347), .Z(n41349) );
  AND U42235 ( .A(n41350), .B(n41349), .Z(n41540) );
  XOR U42236 ( .A(n41541), .B(n41540), .Z(n41543) );
  NANDN U42237 ( .A(n41352), .B(n41351), .Z(n41356) );
  NANDN U42238 ( .A(n41354), .B(n41353), .Z(n41355) );
  AND U42239 ( .A(n41356), .B(n41355), .Z(n41542) );
  XOR U42240 ( .A(n41543), .B(n41542), .Z(n41419) );
  XOR U42241 ( .A(n41418), .B(n41419), .Z(n41420) );
  NANDN U42242 ( .A(n41358), .B(n41357), .Z(n41362) );
  NAND U42243 ( .A(n41360), .B(n41359), .Z(n41361) );
  NAND U42244 ( .A(n41362), .B(n41361), .Z(n41426) );
  NAND U42245 ( .A(n41364), .B(n41363), .Z(n41368) );
  NANDN U42246 ( .A(n41366), .B(n41365), .Z(n41367) );
  NAND U42247 ( .A(n41368), .B(n41367), .Z(n41431) );
  NAND U42248 ( .A(n41370), .B(n41369), .Z(n41374) );
  NAND U42249 ( .A(n41372), .B(n41371), .Z(n41373) );
  NAND U42250 ( .A(n41374), .B(n41373), .Z(n41430) );
  XOR U42251 ( .A(n41431), .B(n41430), .Z(n41433) );
  AND U42252 ( .A(x[501]), .B(y[8104]), .Z(n42268) );
  NAND U42253 ( .A(n41375), .B(n42268), .Z(n41379) );
  NANDN U42254 ( .A(n41377), .B(n41376), .Z(n41378) );
  AND U42255 ( .A(n41379), .B(n41378), .Z(n41531) );
  AND U42256 ( .A(x[502]), .B(y[8099]), .Z(n41500) );
  AND U42257 ( .A(x[485]), .B(y[8116]), .Z(n41499) );
  NAND U42258 ( .A(x[497]), .B(y[8104]), .Z(n41498) );
  XOR U42259 ( .A(n41499), .B(n41498), .Z(n41501) );
  XOR U42260 ( .A(n41500), .B(n41501), .Z(n41529) );
  AND U42261 ( .A(y[8101]), .B(x[500]), .Z(n41381) );
  NAND U42262 ( .A(y[8100]), .B(x[501]), .Z(n41380) );
  XNOR U42263 ( .A(n41381), .B(n41380), .Z(n41512) );
  NAND U42264 ( .A(x[499]), .B(y[8102]), .Z(n41513) );
  XNOR U42265 ( .A(n41512), .B(n41513), .Z(n41528) );
  XNOR U42266 ( .A(n41529), .B(n41528), .Z(n41530) );
  XOR U42267 ( .A(n41531), .B(n41530), .Z(n41459) );
  NANDN U42268 ( .A(n41511), .B(n41692), .Z(n41385) );
  NAND U42269 ( .A(n41383), .B(n41382), .Z(n41384) );
  AND U42270 ( .A(n41385), .B(n41384), .Z(n41536) );
  AND U42271 ( .A(x[495]), .B(y[8106]), .Z(n41518) );
  AND U42272 ( .A(x[498]), .B(y[8103]), .Z(n41517) );
  NAND U42273 ( .A(x[486]), .B(y[8115]), .Z(n41516) );
  XOR U42274 ( .A(n41517), .B(n41516), .Z(n41519) );
  XOR U42275 ( .A(n41518), .B(n41519), .Z(n41535) );
  AND U42276 ( .A(x[503]), .B(y[8098]), .Z(n41494) );
  AND U42277 ( .A(x[484]), .B(y[8117]), .Z(n41493) );
  NAND U42278 ( .A(x[496]), .B(y[8105]), .Z(n41492) );
  XOR U42279 ( .A(n41493), .B(n41492), .Z(n41495) );
  XNOR U42280 ( .A(n41494), .B(n41495), .Z(n41534) );
  XOR U42281 ( .A(n41535), .B(n41534), .Z(n41537) );
  XNOR U42282 ( .A(n41536), .B(n41537), .Z(n41458) );
  XOR U42283 ( .A(n41459), .B(n41458), .Z(n41461) );
  XOR U42284 ( .A(n41461), .B(n41460), .Z(n41470) );
  XNOR U42285 ( .A(n41468), .B(n41469), .Z(n41471) );
  XOR U42286 ( .A(n41470), .B(n41471), .Z(n41432) );
  XOR U42287 ( .A(n41433), .B(n41432), .Z(n41425) );
  NAND U42288 ( .A(n41399), .B(n41398), .Z(n41403) );
  NAND U42289 ( .A(n41401), .B(n41400), .Z(n41402) );
  NAND U42290 ( .A(n41403), .B(n41402), .Z(n41424) );
  XOR U42291 ( .A(n41426), .B(n41427), .Z(n41421) );
  XNOR U42292 ( .A(n41420), .B(n41421), .Z(n41552) );
  XNOR U42293 ( .A(n41555), .B(n41554), .Z(n41561) );
  OR U42294 ( .A(n41406), .B(n41404), .Z(n41410) );
  ANDN U42295 ( .B(n41406), .A(n41405), .Z(n41408) );
  OR U42296 ( .A(n41408), .B(n41407), .Z(n41409) );
  AND U42297 ( .A(n41410), .B(n41409), .Z(n41559) );
  NAND U42298 ( .A(n41412), .B(n41411), .Z(n41416) );
  NAND U42299 ( .A(n41414), .B(n41413), .Z(n41415) );
  AND U42300 ( .A(n41416), .B(n41415), .Z(n41560) );
  IV U42301 ( .A(n41560), .Z(n41558) );
  XOR U42302 ( .A(n41559), .B(n41558), .Z(n41417) );
  XNOR U42303 ( .A(n41561), .B(n41417), .Z(N890) );
  NAND U42304 ( .A(n41419), .B(n41418), .Z(n41423) );
  NANDN U42305 ( .A(n41421), .B(n41420), .Z(n41422) );
  AND U42306 ( .A(n41423), .B(n41422), .Z(n41567) );
  NANDN U42307 ( .A(n41425), .B(n41424), .Z(n41429) );
  NANDN U42308 ( .A(n41427), .B(n41426), .Z(n41428) );
  AND U42309 ( .A(n41429), .B(n41428), .Z(n41566) );
  XOR U42310 ( .A(n41567), .B(n41566), .Z(n41569) );
  NAND U42311 ( .A(n41431), .B(n41430), .Z(n41435) );
  NAND U42312 ( .A(n41433), .B(n41432), .Z(n41434) );
  NAND U42313 ( .A(n41435), .B(n41434), .Z(n41583) );
  AND U42314 ( .A(x[482]), .B(y[8120]), .Z(n41638) );
  XOR U42315 ( .A(n41639), .B(n41638), .Z(n41641) );
  NAND U42316 ( .A(x[504]), .B(y[8098]), .Z(n41640) );
  XNOR U42317 ( .A(n41641), .B(n41640), .Z(n41597) );
  NANDN U42318 ( .A(n41437), .B(n41436), .Z(n41441) );
  OR U42319 ( .A(n41439), .B(n41438), .Z(n41440) );
  NAND U42320 ( .A(n41441), .B(n41440), .Z(n41598) );
  XNOR U42321 ( .A(n41597), .B(n41598), .Z(n41600) );
  NANDN U42322 ( .A(n41443), .B(n41442), .Z(n41447) );
  NANDN U42323 ( .A(n41445), .B(n41444), .Z(n41446) );
  AND U42324 ( .A(n41447), .B(n41446), .Z(n41599) );
  XOR U42325 ( .A(n41600), .B(n41599), .Z(n41669) );
  XNOR U42326 ( .A(n41669), .B(n41668), .Z(n41670) );
  NANDN U42327 ( .A(n41453), .B(n41452), .Z(n41457) );
  NAND U42328 ( .A(n41455), .B(n41454), .Z(n41456) );
  NAND U42329 ( .A(n41457), .B(n41456), .Z(n41671) );
  XNOR U42330 ( .A(n41670), .B(n41671), .Z(n41714) );
  NAND U42331 ( .A(n41459), .B(n41458), .Z(n41463) );
  NAND U42332 ( .A(n41461), .B(n41460), .Z(n41462) );
  NAND U42333 ( .A(n41463), .B(n41462), .Z(n41713) );
  XNOR U42334 ( .A(n41713), .B(n41712), .Z(n41715) );
  XOR U42335 ( .A(n41714), .B(n41715), .Z(n41581) );
  AND U42336 ( .A(x[492]), .B(y[8110]), .Z(n41767) );
  AND U42337 ( .A(x[485]), .B(y[8117]), .Z(n41611) );
  XOR U42338 ( .A(n41767), .B(n41611), .Z(n41613) );
  NAND U42339 ( .A(x[490]), .B(y[8112]), .Z(n41612) );
  XNOR U42340 ( .A(n41613), .B(n41612), .Z(n41677) );
  AND U42341 ( .A(y[8116]), .B(x[486]), .Z(n41473) );
  NAND U42342 ( .A(y[8114]), .B(x[488]), .Z(n41472) );
  XNOR U42343 ( .A(n41473), .B(n41472), .Z(n41693) );
  NAND U42344 ( .A(x[489]), .B(y[8113]), .Z(n41694) );
  XNOR U42345 ( .A(n41693), .B(n41694), .Z(n41675) );
  AND U42346 ( .A(x[487]), .B(y[8115]), .Z(n41674) );
  XOR U42347 ( .A(n41675), .B(n41674), .Z(n41676) );
  XOR U42348 ( .A(n41677), .B(n41676), .Z(n41665) );
  NANDN U42349 ( .A(n41475), .B(n41474), .Z(n41479) );
  NANDN U42350 ( .A(n41477), .B(n41476), .Z(n41478) );
  AND U42351 ( .A(n41479), .B(n41478), .Z(n41663) );
  NANDN U42352 ( .A(n41481), .B(n41480), .Z(n41485) );
  NANDN U42353 ( .A(n41483), .B(n41482), .Z(n41484) );
  NAND U42354 ( .A(n41485), .B(n41484), .Z(n41662) );
  XNOR U42355 ( .A(n41663), .B(n41662), .Z(n41664) );
  XOR U42356 ( .A(n41665), .B(n41664), .Z(n41623) );
  NANDN U42357 ( .A(n41487), .B(n41486), .Z(n41491) );
  NANDN U42358 ( .A(n41489), .B(n41488), .Z(n41490) );
  AND U42359 ( .A(n41491), .B(n41490), .Z(n41622) );
  XNOR U42360 ( .A(n41623), .B(n41622), .Z(n41624) );
  NANDN U42361 ( .A(n41493), .B(n41492), .Z(n41497) );
  OR U42362 ( .A(n41495), .B(n41494), .Z(n41496) );
  AND U42363 ( .A(n41497), .B(n41496), .Z(n41628) );
  NANDN U42364 ( .A(n41499), .B(n41498), .Z(n41503) );
  OR U42365 ( .A(n41501), .B(n41500), .Z(n41502) );
  NAND U42366 ( .A(n41503), .B(n41502), .Z(n41629) );
  XNOR U42367 ( .A(n41628), .B(n41629), .Z(n41631) );
  ANDN U42368 ( .B(o[441]), .A(n41504), .Z(n41686) );
  NAND U42369 ( .A(x[494]), .B(y[8108]), .Z(n41687) );
  XNOR U42370 ( .A(n41686), .B(n41687), .Z(n41688) );
  NAND U42371 ( .A(x[481]), .B(y[8121]), .Z(n41689) );
  XNOR U42372 ( .A(n41688), .B(n41689), .Z(n41603) );
  NAND U42373 ( .A(x[505]), .B(y[8097]), .Z(n41697) );
  XNOR U42374 ( .A(o[442]), .B(n41697), .Z(n41616) );
  NAND U42375 ( .A(x[506]), .B(y[8096]), .Z(n41617) );
  XNOR U42376 ( .A(n41616), .B(n41617), .Z(n41618) );
  NAND U42377 ( .A(x[480]), .B(y[8122]), .Z(n41619) );
  XOR U42378 ( .A(n41618), .B(n41619), .Z(n41604) );
  XNOR U42379 ( .A(n41603), .B(n41604), .Z(n41605) );
  NANDN U42380 ( .A(n41506), .B(n41505), .Z(n41510) );
  OR U42381 ( .A(n41508), .B(n41507), .Z(n41509) );
  NAND U42382 ( .A(n41510), .B(n41509), .Z(n41606) );
  XNOR U42383 ( .A(n41605), .B(n41606), .Z(n41630) );
  XOR U42384 ( .A(n41631), .B(n41630), .Z(n41594) );
  AND U42385 ( .A(x[501]), .B(y[8101]), .Z(n41681) );
  NANDN U42386 ( .A(n41511), .B(n41681), .Z(n41515) );
  NANDN U42387 ( .A(n41513), .B(n41512), .Z(n41514) );
  AND U42388 ( .A(n41515), .B(n41514), .Z(n41658) );
  XOR U42389 ( .A(n41681), .B(n41680), .Z(n41683) );
  NAND U42390 ( .A(x[500]), .B(y[8102]), .Z(n41682) );
  XNOR U42391 ( .A(n41683), .B(n41682), .Z(n41656) );
  NAND U42392 ( .A(x[503]), .B(y[8099]), .Z(n41645) );
  XNOR U42393 ( .A(n41644), .B(n41645), .Z(n41646) );
  NAND U42394 ( .A(x[502]), .B(y[8100]), .Z(n41647) );
  XOR U42395 ( .A(n41646), .B(n41647), .Z(n41657) );
  XOR U42396 ( .A(n41656), .B(n41657), .Z(n41659) );
  XOR U42397 ( .A(n41658), .B(n41659), .Z(n41592) );
  AND U42398 ( .A(x[483]), .B(y[8119]), .Z(n41698) );
  NAND U42399 ( .A(x[499]), .B(y[8103]), .Z(n41699) );
  XNOR U42400 ( .A(n41698), .B(n41699), .Z(n41700) );
  NAND U42401 ( .A(x[491]), .B(y[8111]), .Z(n41701) );
  XNOR U42402 ( .A(n41700), .B(n41701), .Z(n41635) );
  AND U42403 ( .A(x[484]), .B(y[8118]), .Z(n41650) );
  XNOR U42404 ( .A(n41651), .B(n41650), .Z(n41652) );
  XNOR U42405 ( .A(n41653), .B(n41652), .Z(n41634) );
  XOR U42406 ( .A(n41635), .B(n41634), .Z(n41637) );
  NANDN U42407 ( .A(n41517), .B(n41516), .Z(n41521) );
  OR U42408 ( .A(n41519), .B(n41518), .Z(n41520) );
  AND U42409 ( .A(n41521), .B(n41520), .Z(n41636) );
  XNOR U42410 ( .A(n41637), .B(n41636), .Z(n41591) );
  XNOR U42411 ( .A(n41592), .B(n41591), .Z(n41593) );
  XOR U42412 ( .A(n41594), .B(n41593), .Z(n41625) );
  XOR U42413 ( .A(n41624), .B(n41625), .Z(n41587) );
  NANDN U42414 ( .A(n41523), .B(n41522), .Z(n41527) );
  NANDN U42415 ( .A(n41525), .B(n41524), .Z(n41526) );
  AND U42416 ( .A(n41527), .B(n41526), .Z(n41709) );
  NANDN U42417 ( .A(n41529), .B(n41528), .Z(n41533) );
  NANDN U42418 ( .A(n41531), .B(n41530), .Z(n41532) );
  AND U42419 ( .A(n41533), .B(n41532), .Z(n41707) );
  NANDN U42420 ( .A(n41535), .B(n41534), .Z(n41539) );
  OR U42421 ( .A(n41537), .B(n41536), .Z(n41538) );
  NAND U42422 ( .A(n41539), .B(n41538), .Z(n41706) );
  XNOR U42423 ( .A(n41707), .B(n41706), .Z(n41708) );
  XNOR U42424 ( .A(n41709), .B(n41708), .Z(n41588) );
  XOR U42425 ( .A(n41587), .B(n41588), .Z(n41590) );
  XOR U42426 ( .A(n41589), .B(n41590), .Z(n41582) );
  XOR U42427 ( .A(n41581), .B(n41582), .Z(n41584) );
  XOR U42428 ( .A(n41583), .B(n41584), .Z(n41578) );
  NAND U42429 ( .A(n41541), .B(n41540), .Z(n41545) );
  NAND U42430 ( .A(n41543), .B(n41542), .Z(n41544) );
  AND U42431 ( .A(n41545), .B(n41544), .Z(n41576) );
  NAND U42432 ( .A(n41547), .B(n41546), .Z(n41551) );
  NANDN U42433 ( .A(n41549), .B(n41548), .Z(n41550) );
  AND U42434 ( .A(n41551), .B(n41550), .Z(n41575) );
  XOR U42435 ( .A(n41576), .B(n41575), .Z(n41577) );
  XOR U42436 ( .A(n41578), .B(n41577), .Z(n41568) );
  XOR U42437 ( .A(n41569), .B(n41568), .Z(n41574) );
  NANDN U42438 ( .A(n41553), .B(n41552), .Z(n41557) );
  NAND U42439 ( .A(n41555), .B(n41554), .Z(n41556) );
  NAND U42440 ( .A(n41557), .B(n41556), .Z(n41572) );
  NANDN U42441 ( .A(n41558), .B(n41559), .Z(n41564) );
  NOR U42442 ( .A(n41560), .B(n41559), .Z(n41562) );
  OR U42443 ( .A(n41562), .B(n41561), .Z(n41563) );
  AND U42444 ( .A(n41564), .B(n41563), .Z(n41573) );
  XOR U42445 ( .A(n41572), .B(n41573), .Z(n41565) );
  XNOR U42446 ( .A(n41574), .B(n41565), .Z(N891) );
  NAND U42447 ( .A(n41567), .B(n41566), .Z(n41571) );
  NAND U42448 ( .A(n41569), .B(n41568), .Z(n41570) );
  AND U42449 ( .A(n41571), .B(n41570), .Z(n41862) );
  NAND U42450 ( .A(n41576), .B(n41575), .Z(n41580) );
  NAND U42451 ( .A(n41578), .B(n41577), .Z(n41579) );
  NAND U42452 ( .A(n41580), .B(n41579), .Z(n41867) );
  NAND U42453 ( .A(n41582), .B(n41581), .Z(n41586) );
  NAND U42454 ( .A(n41584), .B(n41583), .Z(n41585) );
  NAND U42455 ( .A(n41586), .B(n41585), .Z(n41865) );
  NANDN U42456 ( .A(n41592), .B(n41591), .Z(n41596) );
  NANDN U42457 ( .A(n41594), .B(n41593), .Z(n41595) );
  AND U42458 ( .A(n41596), .B(n41595), .Z(n41844) );
  NANDN U42459 ( .A(n41598), .B(n41597), .Z(n41602) );
  NAND U42460 ( .A(n41600), .B(n41599), .Z(n41601) );
  AND U42461 ( .A(n41602), .B(n41601), .Z(n41835) );
  NANDN U42462 ( .A(n41604), .B(n41603), .Z(n41608) );
  NANDN U42463 ( .A(n41606), .B(n41605), .Z(n41607) );
  AND U42464 ( .A(n41608), .B(n41607), .Z(n41833) );
  AND U42465 ( .A(x[495]), .B(y[8108]), .Z(n41772) );
  NAND U42466 ( .A(x[482]), .B(y[8121]), .Z(n41773) );
  XNOR U42467 ( .A(n41772), .B(n41773), .Z(n41774) );
  NAND U42468 ( .A(x[483]), .B(y[8120]), .Z(n41775) );
  XNOR U42469 ( .A(n41774), .B(n41775), .Z(n41794) );
  AND U42470 ( .A(x[499]), .B(y[8104]), .Z(n41805) );
  NAND U42471 ( .A(x[505]), .B(y[8098]), .Z(n41806) );
  XNOR U42472 ( .A(n41805), .B(n41806), .Z(n41807) );
  NAND U42473 ( .A(x[486]), .B(y[8117]), .Z(n41808) );
  XOR U42474 ( .A(n41807), .B(n41808), .Z(n41795) );
  XNOR U42475 ( .A(n41794), .B(n41795), .Z(n41796) );
  NAND U42476 ( .A(x[496]), .B(y[8107]), .Z(n41755) );
  XOR U42477 ( .A(n41756), .B(n41755), .Z(n41758) );
  XOR U42478 ( .A(n41757), .B(n41758), .Z(n41769) );
  AND U42479 ( .A(y[8110]), .B(x[493]), .Z(n41610) );
  NAND U42480 ( .A(y[8111]), .B(x[492]), .Z(n41609) );
  XNOR U42481 ( .A(n41610), .B(n41609), .Z(n41768) );
  XOR U42482 ( .A(n41769), .B(n41768), .Z(n41797) );
  XNOR U42483 ( .A(n41796), .B(n41797), .Z(n41735) );
  NAND U42484 ( .A(n41767), .B(n41611), .Z(n41615) );
  ANDN U42485 ( .B(n41613), .A(n41612), .Z(n41614) );
  ANDN U42486 ( .B(n41615), .A(n41614), .Z(n41734) );
  NANDN U42487 ( .A(n41617), .B(n41616), .Z(n41621) );
  NANDN U42488 ( .A(n41619), .B(n41618), .Z(n41620) );
  NAND U42489 ( .A(n41621), .B(n41620), .Z(n41733) );
  XOR U42490 ( .A(n41734), .B(n41733), .Z(n41736) );
  XNOR U42491 ( .A(n41735), .B(n41736), .Z(n41832) );
  XNOR U42492 ( .A(n41833), .B(n41832), .Z(n41834) );
  XOR U42493 ( .A(n41835), .B(n41834), .Z(n41845) );
  XNOR U42494 ( .A(n41844), .B(n41845), .Z(n41846) );
  NANDN U42495 ( .A(n41623), .B(n41622), .Z(n41627) );
  NANDN U42496 ( .A(n41625), .B(n41624), .Z(n41626) );
  NAND U42497 ( .A(n41627), .B(n41626), .Z(n41847) );
  XOR U42498 ( .A(n41846), .B(n41847), .Z(n41721) );
  NANDN U42499 ( .A(n41629), .B(n41628), .Z(n41633) );
  NAND U42500 ( .A(n41631), .B(n41630), .Z(n41632) );
  AND U42501 ( .A(n41633), .B(n41632), .Z(n41840) );
  NAND U42502 ( .A(n41639), .B(n41638), .Z(n41643) );
  ANDN U42503 ( .B(n41641), .A(n41640), .Z(n41642) );
  ANDN U42504 ( .B(n41643), .A(n41642), .Z(n41740) );
  NANDN U42505 ( .A(n41645), .B(n41644), .Z(n41649) );
  NANDN U42506 ( .A(n41647), .B(n41646), .Z(n41648) );
  NAND U42507 ( .A(n41649), .B(n41648), .Z(n41739) );
  XNOR U42508 ( .A(n41740), .B(n41739), .Z(n41741) );
  NAND U42509 ( .A(n41651), .B(n41650), .Z(n41655) );
  ANDN U42510 ( .B(n41653), .A(n41652), .Z(n41654) );
  ANDN U42511 ( .B(n41655), .A(n41654), .Z(n41752) );
  AND U42512 ( .A(x[480]), .B(y[8123]), .Z(n41817) );
  NAND U42513 ( .A(x[507]), .B(y[8096]), .Z(n41818) );
  XNOR U42514 ( .A(n41817), .B(n41818), .Z(n41819) );
  NAND U42515 ( .A(x[506]), .B(y[8097]), .Z(n41823) );
  XOR U42516 ( .A(o[443]), .B(n41823), .Z(n41820) );
  XNOR U42517 ( .A(n41819), .B(n41820), .Z(n41749) );
  AND U42518 ( .A(x[489]), .B(y[8114]), .Z(n41826) );
  NAND U42519 ( .A(x[501]), .B(y[8102]), .Z(n41827) );
  XNOR U42520 ( .A(n41826), .B(n41827), .Z(n41828) );
  NAND U42521 ( .A(x[498]), .B(y[8105]), .Z(n41829) );
  XOR U42522 ( .A(n41828), .B(n41829), .Z(n41750) );
  XNOR U42523 ( .A(n41749), .B(n41750), .Z(n41751) );
  XOR U42524 ( .A(n41752), .B(n41751), .Z(n41742) );
  XNOR U42525 ( .A(n41741), .B(n41742), .Z(n41838) );
  XOR U42526 ( .A(n41839), .B(n41838), .Z(n41841) );
  XOR U42527 ( .A(n41840), .B(n41841), .Z(n41858) );
  NANDN U42528 ( .A(n41657), .B(n41656), .Z(n41661) );
  OR U42529 ( .A(n41659), .B(n41658), .Z(n41660) );
  AND U42530 ( .A(n41661), .B(n41660), .Z(n41856) );
  NANDN U42531 ( .A(n41663), .B(n41662), .Z(n41667) );
  NAND U42532 ( .A(n41665), .B(n41664), .Z(n41666) );
  NAND U42533 ( .A(n41667), .B(n41666), .Z(n41857) );
  XOR U42534 ( .A(n41856), .B(n41857), .Z(n41859) );
  XNOR U42535 ( .A(n41858), .B(n41859), .Z(n41722) );
  XOR U42536 ( .A(n41721), .B(n41722), .Z(n41724) );
  XOR U42537 ( .A(n41723), .B(n41724), .Z(n41719) );
  NANDN U42538 ( .A(n41669), .B(n41668), .Z(n41673) );
  NANDN U42539 ( .A(n41671), .B(n41670), .Z(n41672) );
  AND U42540 ( .A(n41673), .B(n41672), .Z(n41728) );
  NAND U42541 ( .A(n41675), .B(n41674), .Z(n41679) );
  NAND U42542 ( .A(n41677), .B(n41676), .Z(n41678) );
  AND U42543 ( .A(n41679), .B(n41678), .Z(n41852) );
  NAND U42544 ( .A(n41681), .B(n41680), .Z(n41685) );
  ANDN U42545 ( .B(n41683), .A(n41682), .Z(n41684) );
  ANDN U42546 ( .B(n41685), .A(n41684), .Z(n41785) );
  NANDN U42547 ( .A(n41687), .B(n41686), .Z(n41691) );
  NANDN U42548 ( .A(n41689), .B(n41688), .Z(n41690) );
  NAND U42549 ( .A(n41691), .B(n41690), .Z(n41784) );
  XNOR U42550 ( .A(n41785), .B(n41784), .Z(n41787) );
  AND U42551 ( .A(x[488]), .B(y[8116]), .Z(n41825) );
  NAND U42552 ( .A(n41692), .B(n41825), .Z(n41696) );
  NANDN U42553 ( .A(n41694), .B(n41693), .Z(n41695) );
  NAND U42554 ( .A(n41696), .B(n41695), .Z(n41747) );
  ANDN U42555 ( .B(o[442]), .A(n41697), .Z(n41780) );
  AND U42556 ( .A(x[494]), .B(y[8109]), .Z(n41778) );
  NAND U42557 ( .A(x[481]), .B(y[8122]), .Z(n41779) );
  XOR U42558 ( .A(n41778), .B(n41779), .Z(n41781) );
  XNOR U42559 ( .A(n41780), .B(n41781), .Z(n41746) );
  AND U42560 ( .A(x[497]), .B(y[8106]), .Z(n41811) );
  NAND U42561 ( .A(x[484]), .B(y[8119]), .Z(n41812) );
  XNOR U42562 ( .A(n41811), .B(n41812), .Z(n41814) );
  AND U42563 ( .A(x[485]), .B(y[8118]), .Z(n41813) );
  XOR U42564 ( .A(n41814), .B(n41813), .Z(n41745) );
  XOR U42565 ( .A(n41746), .B(n41745), .Z(n41748) );
  XOR U42566 ( .A(n41747), .B(n41748), .Z(n41786) );
  XOR U42567 ( .A(n41787), .B(n41786), .Z(n41850) );
  NANDN U42568 ( .A(n41699), .B(n41698), .Z(n41703) );
  NANDN U42569 ( .A(n41701), .B(n41700), .Z(n41702) );
  AND U42570 ( .A(n41703), .B(n41702), .Z(n41791) );
  AND U42571 ( .A(y[8099]), .B(x[504]), .Z(n41705) );
  NAND U42572 ( .A(y[8103]), .B(x[500]), .Z(n41704) );
  XNOR U42573 ( .A(n41705), .B(n41704), .Z(n41801) );
  NAND U42574 ( .A(x[487]), .B(y[8116]), .Z(n41802) );
  XNOR U42575 ( .A(n41801), .B(n41802), .Z(n41788) );
  AND U42576 ( .A(x[488]), .B(y[8115]), .Z(n41761) );
  NAND U42577 ( .A(x[503]), .B(y[8100]), .Z(n41762) );
  XNOR U42578 ( .A(n41761), .B(n41762), .Z(n41763) );
  NAND U42579 ( .A(x[502]), .B(y[8101]), .Z(n41764) );
  XOR U42580 ( .A(n41763), .B(n41764), .Z(n41789) );
  XNOR U42581 ( .A(n41788), .B(n41789), .Z(n41790) );
  XOR U42582 ( .A(n41791), .B(n41790), .Z(n41851) );
  XOR U42583 ( .A(n41850), .B(n41851), .Z(n41853) );
  XNOR U42584 ( .A(n41852), .B(n41853), .Z(n41727) );
  XNOR U42585 ( .A(n41728), .B(n41727), .Z(n41729) );
  NANDN U42586 ( .A(n41707), .B(n41706), .Z(n41711) );
  NANDN U42587 ( .A(n41709), .B(n41708), .Z(n41710) );
  NAND U42588 ( .A(n41711), .B(n41710), .Z(n41730) );
  XOR U42589 ( .A(n41729), .B(n41730), .Z(n41717) );
  XOR U42590 ( .A(n41717), .B(n41718), .Z(n41720) );
  XOR U42591 ( .A(n41719), .B(n41720), .Z(n41866) );
  XOR U42592 ( .A(n41865), .B(n41866), .Z(n41868) );
  XOR U42593 ( .A(n41867), .B(n41868), .Z(n41864) );
  XNOR U42594 ( .A(n41863), .B(n41864), .Z(n41716) );
  XOR U42595 ( .A(n41862), .B(n41716), .Z(N892) );
  NANDN U42596 ( .A(n41722), .B(n41721), .Z(n41726) );
  NANDN U42597 ( .A(n41724), .B(n41723), .Z(n41725) );
  AND U42598 ( .A(n41726), .B(n41725), .Z(n41873) );
  XOR U42599 ( .A(n41872), .B(n41873), .Z(n41875) );
  NANDN U42600 ( .A(n41728), .B(n41727), .Z(n41732) );
  NANDN U42601 ( .A(n41730), .B(n41729), .Z(n41731) );
  AND U42602 ( .A(n41732), .B(n41731), .Z(n41879) );
  NANDN U42603 ( .A(n41734), .B(n41733), .Z(n41738) );
  NANDN U42604 ( .A(n41736), .B(n41735), .Z(n41737) );
  AND U42605 ( .A(n41738), .B(n41737), .Z(n41892) );
  NANDN U42606 ( .A(n41740), .B(n41739), .Z(n41744) );
  NANDN U42607 ( .A(n41742), .B(n41741), .Z(n41743) );
  AND U42608 ( .A(n41744), .B(n41743), .Z(n41997) );
  NANDN U42609 ( .A(n41750), .B(n41749), .Z(n41754) );
  NANDN U42610 ( .A(n41752), .B(n41751), .Z(n41753) );
  NAND U42611 ( .A(n41754), .B(n41753), .Z(n41994) );
  XNOR U42612 ( .A(n41995), .B(n41994), .Z(n41996) );
  XNOR U42613 ( .A(n41997), .B(n41996), .Z(n41891) );
  XNOR U42614 ( .A(n41892), .B(n41891), .Z(n41894) );
  NANDN U42615 ( .A(n41756), .B(n41755), .Z(n41760) );
  OR U42616 ( .A(n41758), .B(n41757), .Z(n41759) );
  AND U42617 ( .A(n41760), .B(n41759), .Z(n41972) );
  AND U42618 ( .A(x[487]), .B(y[8117]), .Z(n41938) );
  AND U42619 ( .A(x[492]), .B(y[8112]), .Z(n41939) );
  XOR U42620 ( .A(n41938), .B(n41939), .Z(n41941) );
  AND U42621 ( .A(x[491]), .B(y[8113]), .Z(n41940) );
  XOR U42622 ( .A(n41941), .B(n41940), .Z(n41971) );
  AND U42623 ( .A(x[507]), .B(y[8097]), .Z(n41955) );
  XOR U42624 ( .A(o[444]), .B(n41955), .Z(n41958) );
  NAND U42625 ( .A(x[506]), .B(y[8098]), .Z(n41959) );
  XNOR U42626 ( .A(n41958), .B(n41959), .Z(n41961) );
  AND U42627 ( .A(x[495]), .B(y[8109]), .Z(n41960) );
  XNOR U42628 ( .A(n41961), .B(n41960), .Z(n41970) );
  XOR U42629 ( .A(n41971), .B(n41970), .Z(n41973) );
  XOR U42630 ( .A(n41972), .B(n41973), .Z(n42019) );
  NANDN U42631 ( .A(n41762), .B(n41761), .Z(n41766) );
  NANDN U42632 ( .A(n41764), .B(n41763), .Z(n41765) );
  AND U42633 ( .A(n41766), .B(n41765), .Z(n41979) );
  AND U42634 ( .A(x[497]), .B(y[8107]), .Z(n41903) );
  NAND U42635 ( .A(x[502]), .B(y[8102]), .Z(n41904) );
  XNOR U42636 ( .A(n41903), .B(n41904), .Z(n41905) );
  NAND U42637 ( .A(x[484]), .B(y[8120]), .Z(n41906) );
  XNOR U42638 ( .A(n41905), .B(n41906), .Z(n41976) );
  AND U42639 ( .A(x[486]), .B(y[8118]), .Z(n42099) );
  NAND U42640 ( .A(x[499]), .B(y[8105]), .Z(n41944) );
  XOR U42641 ( .A(n42099), .B(n41944), .Z(n41946) );
  XOR U42642 ( .A(n41945), .B(n41946), .Z(n41977) );
  XNOR U42643 ( .A(n41976), .B(n41977), .Z(n41978) );
  XNOR U42644 ( .A(n41979), .B(n41978), .Z(n42018) );
  XNOR U42645 ( .A(n42019), .B(n42018), .Z(n42020) );
  NAND U42646 ( .A(n41964), .B(n41767), .Z(n41771) );
  NANDN U42647 ( .A(n41769), .B(n41768), .Z(n41770) );
  AND U42648 ( .A(n41771), .B(n41770), .Z(n41900) );
  NANDN U42649 ( .A(n41773), .B(n41772), .Z(n41777) );
  NANDN U42650 ( .A(n41775), .B(n41774), .Z(n41776) );
  AND U42651 ( .A(n41777), .B(n41776), .Z(n41898) );
  NANDN U42652 ( .A(n41779), .B(n41778), .Z(n41783) );
  NANDN U42653 ( .A(n41781), .B(n41780), .Z(n41782) );
  NAND U42654 ( .A(n41783), .B(n41782), .Z(n41897) );
  XNOR U42655 ( .A(n41898), .B(n41897), .Z(n41899) );
  XOR U42656 ( .A(n41900), .B(n41899), .Z(n42021) );
  XNOR U42657 ( .A(n42020), .B(n42021), .Z(n41893) );
  XOR U42658 ( .A(n41894), .B(n41893), .Z(n42032) );
  NANDN U42659 ( .A(n41789), .B(n41788), .Z(n41793) );
  NANDN U42660 ( .A(n41791), .B(n41790), .Z(n41792) );
  AND U42661 ( .A(n41793), .B(n41792), .Z(n41983) );
  NANDN U42662 ( .A(n41795), .B(n41794), .Z(n41799) );
  NANDN U42663 ( .A(n41797), .B(n41796), .Z(n41798) );
  NAND U42664 ( .A(n41799), .B(n41798), .Z(n41982) );
  XOR U42665 ( .A(n41983), .B(n41982), .Z(n41985) );
  XOR U42666 ( .A(n41984), .B(n41985), .Z(n42031) );
  AND U42667 ( .A(x[500]), .B(y[8099]), .Z(n41800) );
  AND U42668 ( .A(x[504]), .B(y[8103]), .Z(n42285) );
  NAND U42669 ( .A(n41800), .B(n42285), .Z(n41804) );
  NANDN U42670 ( .A(n41802), .B(n41801), .Z(n41803) );
  AND U42671 ( .A(n41804), .B(n41803), .Z(n42014) );
  AND U42672 ( .A(x[505]), .B(y[8099]), .Z(n41934) );
  XOR U42673 ( .A(n41935), .B(n41934), .Z(n41933) );
  NAND U42674 ( .A(x[481]), .B(y[8123]), .Z(n41932) );
  XNOR U42675 ( .A(n41933), .B(n41932), .Z(n42012) );
  AND U42676 ( .A(x[496]), .B(y[8108]), .Z(n41926) );
  NAND U42677 ( .A(x[504]), .B(y[8100]), .Z(n41927) );
  XNOR U42678 ( .A(n41926), .B(n41927), .Z(n41928) );
  NAND U42679 ( .A(x[482]), .B(y[8122]), .Z(n41929) );
  XOR U42680 ( .A(n41928), .B(n41929), .Z(n42013) );
  XOR U42681 ( .A(n42012), .B(n42013), .Z(n42015) );
  XOR U42682 ( .A(n42014), .B(n42015), .Z(n41991) );
  NANDN U42683 ( .A(n41806), .B(n41805), .Z(n41810) );
  NANDN U42684 ( .A(n41808), .B(n41807), .Z(n41809) );
  AND U42685 ( .A(n41810), .B(n41809), .Z(n42008) );
  NAND U42686 ( .A(x[483]), .B(y[8121]), .Z(n41965) );
  XNOR U42687 ( .A(n41964), .B(n41965), .Z(n41966) );
  NAND U42688 ( .A(x[503]), .B(y[8101]), .Z(n41967) );
  XNOR U42689 ( .A(n41966), .B(n41967), .Z(n42006) );
  AND U42690 ( .A(x[485]), .B(y[8119]), .Z(n41949) );
  NAND U42691 ( .A(x[501]), .B(y[8103]), .Z(n41950) );
  XNOR U42692 ( .A(n41949), .B(n41950), .Z(n41951) );
  NAND U42693 ( .A(x[500]), .B(y[8104]), .Z(n41952) );
  XOR U42694 ( .A(n41951), .B(n41952), .Z(n42007) );
  XOR U42695 ( .A(n42006), .B(n42007), .Z(n42009) );
  XOR U42696 ( .A(n42008), .B(n42009), .Z(n41989) );
  NANDN U42697 ( .A(n41812), .B(n41811), .Z(n41816) );
  NAND U42698 ( .A(n41814), .B(n41813), .Z(n41815) );
  AND U42699 ( .A(n41816), .B(n41815), .Z(n42001) );
  NANDN U42700 ( .A(n41818), .B(n41817), .Z(n41822) );
  NANDN U42701 ( .A(n41820), .B(n41819), .Z(n41821) );
  NAND U42702 ( .A(n41822), .B(n41821), .Z(n42000) );
  XNOR U42703 ( .A(n42001), .B(n42000), .Z(n42003) );
  ANDN U42704 ( .B(o[443]), .A(n41823), .Z(n41911) );
  AND U42705 ( .A(x[480]), .B(y[8124]), .Z(n41909) );
  NAND U42706 ( .A(x[508]), .B(y[8096]), .Z(n41910) );
  XOR U42707 ( .A(n41909), .B(n41910), .Z(n41912) );
  XNOR U42708 ( .A(n41911), .B(n41912), .Z(n41920) );
  NAND U42709 ( .A(y[8114]), .B(x[490]), .Z(n41824) );
  XNOR U42710 ( .A(n41825), .B(n41824), .Z(n41916) );
  NAND U42711 ( .A(x[489]), .B(y[8115]), .Z(n41917) );
  XOR U42712 ( .A(n41916), .B(n41917), .Z(n41921) );
  XNOR U42713 ( .A(n41920), .B(n41921), .Z(n41922) );
  NANDN U42714 ( .A(n41827), .B(n41826), .Z(n41831) );
  NANDN U42715 ( .A(n41829), .B(n41828), .Z(n41830) );
  AND U42716 ( .A(n41831), .B(n41830), .Z(n41923) );
  XNOR U42717 ( .A(n41922), .B(n41923), .Z(n42002) );
  XNOR U42718 ( .A(n42003), .B(n42002), .Z(n41988) );
  XNOR U42719 ( .A(n41989), .B(n41988), .Z(n41990) );
  XNOR U42720 ( .A(n41991), .B(n41990), .Z(n42030) );
  XOR U42721 ( .A(n42031), .B(n42030), .Z(n42033) );
  XOR U42722 ( .A(n42032), .B(n42033), .Z(n42027) );
  NANDN U42723 ( .A(n41833), .B(n41832), .Z(n41837) );
  NANDN U42724 ( .A(n41835), .B(n41834), .Z(n41836) );
  AND U42725 ( .A(n41837), .B(n41836), .Z(n42025) );
  NANDN U42726 ( .A(n41839), .B(n41838), .Z(n41843) );
  OR U42727 ( .A(n41841), .B(n41840), .Z(n41842) );
  NAND U42728 ( .A(n41843), .B(n41842), .Z(n42024) );
  XNOR U42729 ( .A(n42025), .B(n42024), .Z(n42026) );
  XOR U42730 ( .A(n42027), .B(n42026), .Z(n41880) );
  XNOR U42731 ( .A(n41879), .B(n41880), .Z(n41881) );
  NANDN U42732 ( .A(n41845), .B(n41844), .Z(n41849) );
  NANDN U42733 ( .A(n41847), .B(n41846), .Z(n41848) );
  AND U42734 ( .A(n41849), .B(n41848), .Z(n41888) );
  NANDN U42735 ( .A(n41851), .B(n41850), .Z(n41855) );
  OR U42736 ( .A(n41853), .B(n41852), .Z(n41854) );
  AND U42737 ( .A(n41855), .B(n41854), .Z(n41886) );
  NANDN U42738 ( .A(n41857), .B(n41856), .Z(n41861) );
  OR U42739 ( .A(n41859), .B(n41858), .Z(n41860) );
  AND U42740 ( .A(n41861), .B(n41860), .Z(n41885) );
  XNOR U42741 ( .A(n41886), .B(n41885), .Z(n41887) );
  XOR U42742 ( .A(n41888), .B(n41887), .Z(n41882) );
  XNOR U42743 ( .A(n41881), .B(n41882), .Z(n41874) );
  XNOR U42744 ( .A(n41875), .B(n41874), .Z(n41878) );
  NAND U42745 ( .A(n41866), .B(n41865), .Z(n41870) );
  NAND U42746 ( .A(n41868), .B(n41867), .Z(n41869) );
  NAND U42747 ( .A(n41870), .B(n41869), .Z(n41876) );
  XOR U42748 ( .A(n41877), .B(n41876), .Z(n41871) );
  XNOR U42749 ( .A(n41878), .B(n41871), .Z(N893) );
  NANDN U42750 ( .A(n41880), .B(n41879), .Z(n41884) );
  NANDN U42751 ( .A(n41882), .B(n41881), .Z(n41883) );
  AND U42752 ( .A(n41884), .B(n41883), .Z(n42043) );
  NANDN U42753 ( .A(n41886), .B(n41885), .Z(n41890) );
  NANDN U42754 ( .A(n41888), .B(n41887), .Z(n41889) );
  AND U42755 ( .A(n41890), .B(n41889), .Z(n42041) );
  NANDN U42756 ( .A(n41892), .B(n41891), .Z(n41896) );
  NAND U42757 ( .A(n41894), .B(n41893), .Z(n41895) );
  AND U42758 ( .A(n41896), .B(n41895), .Z(n42207) );
  NANDN U42759 ( .A(n41898), .B(n41897), .Z(n41902) );
  NANDN U42760 ( .A(n41900), .B(n41899), .Z(n41901) );
  AND U42761 ( .A(n41902), .B(n41901), .Z(n42152) );
  NANDN U42762 ( .A(n41904), .B(n41903), .Z(n41908) );
  NANDN U42763 ( .A(n41906), .B(n41905), .Z(n41907) );
  AND U42764 ( .A(n41908), .B(n41907), .Z(n42174) );
  NANDN U42765 ( .A(n41910), .B(n41909), .Z(n41914) );
  NANDN U42766 ( .A(n41912), .B(n41911), .Z(n41913) );
  NAND U42767 ( .A(n41914), .B(n41913), .Z(n42173) );
  XNOR U42768 ( .A(n42174), .B(n42173), .Z(n42176) );
  AND U42769 ( .A(x[490]), .B(y[8116]), .Z(n42187) );
  NAND U42770 ( .A(n41915), .B(n42187), .Z(n41919) );
  NANDN U42771 ( .A(n41917), .B(n41916), .Z(n41918) );
  AND U42772 ( .A(n41919), .B(n41918), .Z(n42158) );
  AND U42773 ( .A(x[492]), .B(y[8113]), .Z(n42408) );
  AND U42774 ( .A(x[481]), .B(y[8124]), .Z(n42118) );
  XOR U42775 ( .A(n42408), .B(n42118), .Z(n42119) );
  NAND U42776 ( .A(x[502]), .B(y[8103]), .Z(n42120) );
  XNOR U42777 ( .A(n42119), .B(n42120), .Z(n42155) );
  NAND U42778 ( .A(x[495]), .B(y[8110]), .Z(n42123) );
  XOR U42779 ( .A(n42268), .B(n42123), .Z(n42125) );
  XOR U42780 ( .A(n42124), .B(n42125), .Z(n42156) );
  XOR U42781 ( .A(n42176), .B(n42175), .Z(n42150) );
  NANDN U42782 ( .A(n41921), .B(n41920), .Z(n41925) );
  NANDN U42783 ( .A(n41923), .B(n41922), .Z(n41924) );
  AND U42784 ( .A(n41925), .B(n41924), .Z(n42149) );
  XNOR U42785 ( .A(n42150), .B(n42149), .Z(n42151) );
  XOR U42786 ( .A(n42152), .B(n42151), .Z(n42146) );
  NANDN U42787 ( .A(n41927), .B(n41926), .Z(n41931) );
  NANDN U42788 ( .A(n41929), .B(n41928), .Z(n41930) );
  NAND U42789 ( .A(n41931), .B(n41930), .Z(n42162) );
  ANDN U42790 ( .B(n41933), .A(n41932), .Z(n41937) );
  NAND U42791 ( .A(n41935), .B(n41934), .Z(n41936) );
  NANDN U42792 ( .A(n41937), .B(n41936), .Z(n42161) );
  XOR U42793 ( .A(n42162), .B(n42161), .Z(n42163) );
  NAND U42794 ( .A(n41939), .B(n41938), .Z(n41943) );
  NAND U42795 ( .A(n41941), .B(n41940), .Z(n41942) );
  NAND U42796 ( .A(n41943), .B(n41942), .Z(n42061) );
  AND U42797 ( .A(x[504]), .B(y[8101]), .Z(n42401) );
  AND U42798 ( .A(x[493]), .B(y[8112]), .Z(n42088) );
  XOR U42799 ( .A(n42401), .B(n42088), .Z(n42089) );
  NAND U42800 ( .A(x[503]), .B(y[8102]), .Z(n42090) );
  AND U42801 ( .A(x[483]), .B(y[8122]), .Z(n42093) );
  NAND U42802 ( .A(x[497]), .B(y[8108]), .Z(n42094) );
  NAND U42803 ( .A(x[491]), .B(y[8114]), .Z(n42096) );
  XOR U42804 ( .A(n42059), .B(n42058), .Z(n42060) );
  XNOR U42805 ( .A(n42061), .B(n42060), .Z(n42164) );
  XNOR U42806 ( .A(n42163), .B(n42164), .Z(n42134) );
  NANDN U42807 ( .A(n41944), .B(n42099), .Z(n41948) );
  NANDN U42808 ( .A(n41946), .B(n41945), .Z(n41947) );
  AND U42809 ( .A(n41948), .B(n41947), .Z(n42169) );
  AND U42810 ( .A(x[506]), .B(y[8099]), .Z(n42112) );
  XOR U42811 ( .A(n42113), .B(n42112), .Z(n42114) );
  AND U42812 ( .A(x[505]), .B(y[8100]), .Z(n42115) );
  XOR U42813 ( .A(n42114), .B(n42115), .Z(n42168) );
  AND U42814 ( .A(x[508]), .B(y[8097]), .Z(n42130) );
  XOR U42815 ( .A(o[445]), .B(n42130), .Z(n42182) );
  AND U42816 ( .A(x[480]), .B(y[8125]), .Z(n42180) );
  AND U42817 ( .A(x[509]), .B(y[8096]), .Z(n42179) );
  XOR U42818 ( .A(n42180), .B(n42179), .Z(n42181) );
  XNOR U42819 ( .A(n42182), .B(n42181), .Z(n42167) );
  XNOR U42820 ( .A(n42169), .B(n42170), .Z(n42131) );
  NANDN U42821 ( .A(n41950), .B(n41949), .Z(n41954) );
  NANDN U42822 ( .A(n41952), .B(n41951), .Z(n41953) );
  NAND U42823 ( .A(n41954), .B(n41953), .Z(n42109) );
  AND U42824 ( .A(o[444]), .B(n41955), .Z(n42079) );
  AND U42825 ( .A(x[496]), .B(y[8109]), .Z(n42077) );
  AND U42826 ( .A(x[507]), .B(y[8098]), .Z(n42076) );
  XOR U42827 ( .A(n42077), .B(n42076), .Z(n42078) );
  XOR U42828 ( .A(n42079), .B(n42078), .Z(n42107) );
  AND U42829 ( .A(x[482]), .B(y[8123]), .Z(n42070) );
  XOR U42830 ( .A(n42071), .B(n42070), .Z(n42072) );
  XOR U42831 ( .A(n42073), .B(n42072), .Z(n42106) );
  XOR U42832 ( .A(n42107), .B(n42106), .Z(n42108) );
  XOR U42833 ( .A(n42109), .B(n42108), .Z(n42132) );
  AND U42834 ( .A(y[8119]), .B(x[486]), .Z(n41957) );
  NAND U42835 ( .A(y[8118]), .B(x[487]), .Z(n41956) );
  XNOR U42836 ( .A(n41957), .B(n41956), .Z(n42100) );
  NAND U42837 ( .A(x[488]), .B(y[8117]), .Z(n42101) );
  AND U42838 ( .A(x[489]), .B(y[8116]), .Z(n42281) );
  XOR U42839 ( .A(n42189), .B(n42281), .Z(n42191) );
  AND U42840 ( .A(x[484]), .B(y[8121]), .Z(n42064) );
  AND U42841 ( .A(x[490]), .B(y[8115]), .Z(n42065) );
  XOR U42842 ( .A(n42064), .B(n42065), .Z(n42067) );
  AND U42843 ( .A(x[485]), .B(y[8120]), .Z(n42066) );
  XOR U42844 ( .A(n42067), .B(n42066), .Z(n42190) );
  XOR U42845 ( .A(n42191), .B(n42190), .Z(n42085) );
  NANDN U42846 ( .A(n41959), .B(n41958), .Z(n41963) );
  NAND U42847 ( .A(n41961), .B(n41960), .Z(n41962) );
  NAND U42848 ( .A(n41963), .B(n41962), .Z(n42083) );
  NANDN U42849 ( .A(n41965), .B(n41964), .Z(n41969) );
  NANDN U42850 ( .A(n41967), .B(n41966), .Z(n41968) );
  NAND U42851 ( .A(n41969), .B(n41968), .Z(n42082) );
  XOR U42852 ( .A(n42083), .B(n42082), .Z(n42084) );
  XOR U42853 ( .A(n42085), .B(n42084), .Z(n42053) );
  NANDN U42854 ( .A(n41971), .B(n41970), .Z(n41975) );
  OR U42855 ( .A(n41973), .B(n41972), .Z(n41974) );
  NAND U42856 ( .A(n41975), .B(n41974), .Z(n42052) );
  XNOR U42857 ( .A(n42053), .B(n42052), .Z(n42054) );
  XOR U42858 ( .A(n42055), .B(n42054), .Z(n42144) );
  NANDN U42859 ( .A(n41977), .B(n41976), .Z(n41981) );
  NANDN U42860 ( .A(n41979), .B(n41978), .Z(n41980) );
  NAND U42861 ( .A(n41981), .B(n41980), .Z(n42143) );
  XNOR U42862 ( .A(n42144), .B(n42143), .Z(n42145) );
  XNOR U42863 ( .A(n42146), .B(n42145), .Z(n42206) );
  XNOR U42864 ( .A(n42207), .B(n42206), .Z(n42208) );
  NANDN U42865 ( .A(n41983), .B(n41982), .Z(n41987) );
  OR U42866 ( .A(n41985), .B(n41984), .Z(n41986) );
  AND U42867 ( .A(n41987), .B(n41986), .Z(n42201) );
  NANDN U42868 ( .A(n41989), .B(n41988), .Z(n41993) );
  NANDN U42869 ( .A(n41991), .B(n41990), .Z(n41992) );
  AND U42870 ( .A(n41993), .B(n41992), .Z(n42200) );
  XNOR U42871 ( .A(n42201), .B(n42200), .Z(n42202) );
  NANDN U42872 ( .A(n41995), .B(n41994), .Z(n41999) );
  NANDN U42873 ( .A(n41997), .B(n41996), .Z(n41998) );
  AND U42874 ( .A(n41999), .B(n41998), .Z(n42197) );
  NANDN U42875 ( .A(n42001), .B(n42000), .Z(n42005) );
  NAND U42876 ( .A(n42003), .B(n42002), .Z(n42004) );
  AND U42877 ( .A(n42005), .B(n42004), .Z(n42140) );
  NANDN U42878 ( .A(n42007), .B(n42006), .Z(n42011) );
  OR U42879 ( .A(n42009), .B(n42008), .Z(n42010) );
  AND U42880 ( .A(n42011), .B(n42010), .Z(n42138) );
  NANDN U42881 ( .A(n42013), .B(n42012), .Z(n42017) );
  OR U42882 ( .A(n42015), .B(n42014), .Z(n42016) );
  NAND U42883 ( .A(n42017), .B(n42016), .Z(n42137) );
  XNOR U42884 ( .A(n42138), .B(n42137), .Z(n42139) );
  XNOR U42885 ( .A(n42140), .B(n42139), .Z(n42194) );
  NANDN U42886 ( .A(n42019), .B(n42018), .Z(n42023) );
  NANDN U42887 ( .A(n42021), .B(n42020), .Z(n42022) );
  AND U42888 ( .A(n42023), .B(n42022), .Z(n42195) );
  XNOR U42889 ( .A(n42194), .B(n42195), .Z(n42196) );
  XOR U42890 ( .A(n42197), .B(n42196), .Z(n42203) );
  XOR U42891 ( .A(n42202), .B(n42203), .Z(n42209) );
  XNOR U42892 ( .A(n42208), .B(n42209), .Z(n42048) );
  NANDN U42893 ( .A(n42025), .B(n42024), .Z(n42029) );
  NANDN U42894 ( .A(n42027), .B(n42026), .Z(n42028) );
  AND U42895 ( .A(n42029), .B(n42028), .Z(n42047) );
  NANDN U42896 ( .A(n42031), .B(n42030), .Z(n42035) );
  OR U42897 ( .A(n42033), .B(n42032), .Z(n42034) );
  AND U42898 ( .A(n42035), .B(n42034), .Z(n42046) );
  XOR U42899 ( .A(n42047), .B(n42046), .Z(n42049) );
  XNOR U42900 ( .A(n42048), .B(n42049), .Z(n42040) );
  XNOR U42901 ( .A(n42041), .B(n42040), .Z(n42042) );
  XNOR U42902 ( .A(n42043), .B(n42042), .Z(n42039) );
  XOR U42903 ( .A(n42037), .B(n42039), .Z(n42036) );
  XOR U42904 ( .A(n42038), .B(n42036), .Z(N894) );
  NANDN U42905 ( .A(n42041), .B(n42040), .Z(n42045) );
  NANDN U42906 ( .A(n42043), .B(n42042), .Z(n42044) );
  AND U42907 ( .A(n42045), .B(n42044), .Z(n42489) );
  XNOR U42908 ( .A(n42488), .B(n42489), .Z(n42491) );
  NANDN U42909 ( .A(n42047), .B(n42046), .Z(n42051) );
  NANDN U42910 ( .A(n42049), .B(n42048), .Z(n42050) );
  AND U42911 ( .A(n42051), .B(n42050), .Z(n42471) );
  NANDN U42912 ( .A(n42053), .B(n42052), .Z(n42057) );
  NAND U42913 ( .A(n42055), .B(n42054), .Z(n42056) );
  AND U42914 ( .A(n42057), .B(n42056), .Z(n42212) );
  NAND U42915 ( .A(n42059), .B(n42058), .Z(n42063) );
  NAND U42916 ( .A(n42061), .B(n42060), .Z(n42062) );
  AND U42917 ( .A(n42063), .B(n42062), .Z(n42221) );
  NAND U42918 ( .A(n42065), .B(n42064), .Z(n42069) );
  NAND U42919 ( .A(n42067), .B(n42066), .Z(n42068) );
  AND U42920 ( .A(n42069), .B(n42068), .Z(n42232) );
  AND U42921 ( .A(x[486]), .B(y[8120]), .Z(n42351) );
  AND U42922 ( .A(x[485]), .B(y[8121]), .Z(n42353) );
  AND U42923 ( .A(x[499]), .B(y[8107]), .Z(n42352) );
  XOR U42924 ( .A(n42353), .B(n42352), .Z(n42350) );
  XOR U42925 ( .A(n42351), .B(n42350), .Z(n42384) );
  AND U42926 ( .A(x[484]), .B(y[8122]), .Z(n42272) );
  AND U42927 ( .A(x[483]), .B(y[8123]), .Z(n42274) );
  AND U42928 ( .A(x[498]), .B(y[8108]), .Z(n42273) );
  XOR U42929 ( .A(n42274), .B(n42273), .Z(n42271) );
  XNOR U42930 ( .A(n42272), .B(n42271), .Z(n42382) );
  NAND U42931 ( .A(n42071), .B(n42070), .Z(n42075) );
  NAND U42932 ( .A(n42073), .B(n42072), .Z(n42074) );
  AND U42933 ( .A(n42075), .B(n42074), .Z(n42383) );
  XOR U42934 ( .A(n42382), .B(n42383), .Z(n42385) );
  XNOR U42935 ( .A(n42232), .B(n42233), .Z(n42231) );
  NAND U42936 ( .A(n42077), .B(n42076), .Z(n42081) );
  NAND U42937 ( .A(n42079), .B(n42078), .Z(n42080) );
  AND U42938 ( .A(n42081), .B(n42080), .Z(n42230) );
  XOR U42939 ( .A(n42231), .B(n42230), .Z(n42220) );
  XOR U42940 ( .A(n42221), .B(n42220), .Z(n42219) );
  NAND U42941 ( .A(n42083), .B(n42082), .Z(n42087) );
  NAND U42942 ( .A(n42085), .B(n42084), .Z(n42086) );
  AND U42943 ( .A(n42087), .B(n42086), .Z(n42218) );
  XOR U42944 ( .A(n42219), .B(n42218), .Z(n42215) );
  AND U42945 ( .A(n42401), .B(n42088), .Z(n42092) );
  NANDN U42946 ( .A(n42090), .B(n42089), .Z(n42091) );
  NANDN U42947 ( .A(n42092), .B(n42091), .Z(n42227) );
  NANDN U42948 ( .A(n42094), .B(n42093), .Z(n42098) );
  NANDN U42949 ( .A(n42096), .B(n42095), .Z(n42097) );
  AND U42950 ( .A(n42098), .B(n42097), .Z(n42377) );
  AND U42951 ( .A(x[480]), .B(y[8126]), .Z(n42261) );
  AND U42952 ( .A(x[509]), .B(y[8097]), .Z(n42284) );
  XOR U42953 ( .A(o[446]), .B(n42284), .Z(n42263) );
  AND U42954 ( .A(x[510]), .B(y[8096]), .Z(n42262) );
  XOR U42955 ( .A(n42263), .B(n42262), .Z(n42260) );
  XOR U42956 ( .A(n42261), .B(n42260), .Z(n42378) );
  AND U42957 ( .A(x[500]), .B(y[8106]), .Z(n42414) );
  XOR U42958 ( .A(n42415), .B(n42414), .Z(n42413) );
  AND U42959 ( .A(x[488]), .B(y[8118]), .Z(n42412) );
  XNOR U42960 ( .A(n42413), .B(n42412), .Z(n42379) );
  XNOR U42961 ( .A(n42377), .B(n42376), .Z(n42226) );
  XOR U42962 ( .A(n42227), .B(n42226), .Z(n42224) );
  AND U42963 ( .A(x[487]), .B(y[8119]), .Z(n42267) );
  NAND U42964 ( .A(n42099), .B(n42267), .Z(n42103) );
  NANDN U42965 ( .A(n42101), .B(n42100), .Z(n42102) );
  AND U42966 ( .A(n42103), .B(n42102), .Z(n42234) );
  AND U42967 ( .A(y[8105]), .B(x[501]), .Z(n42105) );
  AND U42968 ( .A(y[8104]), .B(x[502]), .Z(n42104) );
  XOR U42969 ( .A(n42105), .B(n42104), .Z(n42266) );
  XOR U42970 ( .A(n42267), .B(n42266), .Z(n42237) );
  AND U42971 ( .A(x[497]), .B(y[8109]), .Z(n42339) );
  AND U42972 ( .A(x[482]), .B(y[8124]), .Z(n42341) );
  AND U42973 ( .A(x[506]), .B(y[8100]), .Z(n42340) );
  XOR U42974 ( .A(n42341), .B(n42340), .Z(n42338) );
  XNOR U42975 ( .A(n42339), .B(n42338), .Z(n42236) );
  XNOR U42976 ( .A(n42234), .B(n42235), .Z(n42225) );
  NAND U42977 ( .A(n42107), .B(n42106), .Z(n42111) );
  NAND U42978 ( .A(n42109), .B(n42108), .Z(n42110) );
  NAND U42979 ( .A(n42111), .B(n42110), .Z(n42448) );
  XOR U42980 ( .A(n42449), .B(n42448), .Z(n42446) );
  AND U42981 ( .A(n42113), .B(n42112), .Z(n42117) );
  NAND U42982 ( .A(n42115), .B(n42114), .Z(n42116) );
  NANDN U42983 ( .A(n42117), .B(n42116), .Z(n42254) );
  AND U42984 ( .A(n42408), .B(n42118), .Z(n42122) );
  NANDN U42985 ( .A(n42120), .B(n42119), .Z(n42121) );
  NANDN U42986 ( .A(n42122), .B(n42121), .Z(n42256) );
  NANDN U42987 ( .A(n42123), .B(n42268), .Z(n42127) );
  NANDN U42988 ( .A(n42125), .B(n42124), .Z(n42126) );
  AND U42989 ( .A(n42127), .B(n42126), .Z(n42246) );
  AND U42990 ( .A(x[503]), .B(y[8103]), .Z(n42399) );
  AND U42991 ( .A(y[8102]), .B(x[504]), .Z(n42129) );
  AND U42992 ( .A(y[8101]), .B(x[505]), .Z(n42128) );
  XOR U42993 ( .A(n42129), .B(n42128), .Z(n42398) );
  XOR U42994 ( .A(n42399), .B(n42398), .Z(n42249) );
  AND U42995 ( .A(o[445]), .B(n42130), .Z(n42393) );
  AND U42996 ( .A(x[508]), .B(y[8098]), .Z(n42395) );
  AND U42997 ( .A(x[496]), .B(y[8110]), .Z(n42394) );
  XOR U42998 ( .A(n42395), .B(n42394), .Z(n42392) );
  XNOR U42999 ( .A(n42393), .B(n42392), .Z(n42248) );
  XNOR U43000 ( .A(n42246), .B(n42247), .Z(n42257) );
  XOR U43001 ( .A(n42254), .B(n42255), .Z(n42447) );
  XNOR U43002 ( .A(n42446), .B(n42447), .Z(n42214) );
  XNOR U43003 ( .A(n42215), .B(n42214), .Z(n42213) );
  XNOR U43004 ( .A(n42212), .B(n42213), .Z(n42458) );
  NANDN U43005 ( .A(n42132), .B(n42131), .Z(n42136) );
  NANDN U43006 ( .A(n42134), .B(n42133), .Z(n42135) );
  NAND U43007 ( .A(n42136), .B(n42135), .Z(n42460) );
  NANDN U43008 ( .A(n42138), .B(n42137), .Z(n42142) );
  NANDN U43009 ( .A(n42140), .B(n42139), .Z(n42141) );
  NAND U43010 ( .A(n42142), .B(n42141), .Z(n42461) );
  XOR U43011 ( .A(n42458), .B(n42459), .Z(n42453) );
  NANDN U43012 ( .A(n42144), .B(n42143), .Z(n42148) );
  NANDN U43013 ( .A(n42146), .B(n42145), .Z(n42147) );
  AND U43014 ( .A(n42148), .B(n42147), .Z(n42455) );
  NANDN U43015 ( .A(n42150), .B(n42149), .Z(n42154) );
  NAND U43016 ( .A(n42152), .B(n42151), .Z(n42153) );
  AND U43017 ( .A(n42154), .B(n42153), .Z(n42443) );
  NANDN U43018 ( .A(n42156), .B(n42155), .Z(n42160) );
  NANDN U43019 ( .A(n42158), .B(n42157), .Z(n42159) );
  AND U43020 ( .A(n42160), .B(n42159), .Z(n42438) );
  NAND U43021 ( .A(n42162), .B(n42161), .Z(n42166) );
  NANDN U43022 ( .A(n42164), .B(n42163), .Z(n42165) );
  NAND U43023 ( .A(n42166), .B(n42165), .Z(n42439) );
  NANDN U43024 ( .A(n42168), .B(n42167), .Z(n42172) );
  NANDN U43025 ( .A(n42170), .B(n42169), .Z(n42171) );
  NAND U43026 ( .A(n42172), .B(n42171), .Z(n42436) );
  XOR U43027 ( .A(n42437), .B(n42436), .Z(n42445) );
  NANDN U43028 ( .A(n42174), .B(n42173), .Z(n42178) );
  NAND U43029 ( .A(n42176), .B(n42175), .Z(n42177) );
  AND U43030 ( .A(n42178), .B(n42177), .Z(n42431) );
  NAND U43031 ( .A(n42180), .B(n42179), .Z(n42184) );
  NAND U43032 ( .A(n42182), .B(n42181), .Z(n42183) );
  AND U43033 ( .A(n42184), .B(n42183), .Z(n42241) );
  AND U43034 ( .A(y[8114]), .B(x[492]), .Z(n42185) );
  XOR U43035 ( .A(n42186), .B(n42185), .Z(n42406) );
  XOR U43036 ( .A(n42407), .B(n42406), .Z(n42280) );
  AND U43037 ( .A(x[489]), .B(y[8117]), .Z(n42188) );
  XOR U43038 ( .A(n42188), .B(n42187), .Z(n42279) );
  XOR U43039 ( .A(n42280), .B(n42279), .Z(n42243) );
  AND U43040 ( .A(x[507]), .B(y[8099]), .Z(n42347) );
  AND U43041 ( .A(x[481]), .B(y[8125]), .Z(n42346) );
  XOR U43042 ( .A(n42347), .B(n42346), .Z(n42344) );
  XOR U43043 ( .A(n42345), .B(n42344), .Z(n42242) );
  XOR U43044 ( .A(n42243), .B(n42242), .Z(n42240) );
  XOR U43045 ( .A(n42241), .B(n42240), .Z(n42432) );
  NAND U43046 ( .A(n42189), .B(n42281), .Z(n42193) );
  NAND U43047 ( .A(n42191), .B(n42190), .Z(n42192) );
  AND U43048 ( .A(n42193), .B(n42192), .Z(n42433) );
  XOR U43049 ( .A(n42432), .B(n42433), .Z(n42430) );
  XNOR U43050 ( .A(n42431), .B(n42430), .Z(n42444) );
  XOR U43051 ( .A(n42443), .B(n42442), .Z(n42454) );
  XOR U43052 ( .A(n42453), .B(n42452), .Z(n42472) );
  NANDN U43053 ( .A(n42195), .B(n42194), .Z(n42199) );
  NANDN U43054 ( .A(n42197), .B(n42196), .Z(n42198) );
  AND U43055 ( .A(n42199), .B(n42198), .Z(n42477) );
  NANDN U43056 ( .A(n42201), .B(n42200), .Z(n42205) );
  NANDN U43057 ( .A(n42203), .B(n42202), .Z(n42204) );
  AND U43058 ( .A(n42205), .B(n42204), .Z(n42478) );
  NANDN U43059 ( .A(n42207), .B(n42206), .Z(n42211) );
  NANDN U43060 ( .A(n42209), .B(n42208), .Z(n42210) );
  NAND U43061 ( .A(n42211), .B(n42210), .Z(n42479) );
  XOR U43062 ( .A(n42477), .B(n42476), .Z(n42473) );
  XOR U43063 ( .A(n42471), .B(n42470), .Z(n42490) );
  XNOR U43064 ( .A(n42491), .B(n42490), .Z(N895) );
  NAND U43065 ( .A(n42213), .B(n42212), .Z(n42217) );
  NANDN U43066 ( .A(n42215), .B(n42214), .Z(n42216) );
  AND U43067 ( .A(n42217), .B(n42216), .Z(n42487) );
  NAND U43068 ( .A(n42219), .B(n42218), .Z(n42223) );
  NAND U43069 ( .A(n42221), .B(n42220), .Z(n42222) );
  AND U43070 ( .A(n42223), .B(n42222), .Z(n42469) );
  NANDN U43071 ( .A(n42225), .B(n42224), .Z(n42229) );
  NAND U43072 ( .A(n42227), .B(n42226), .Z(n42228) );
  AND U43073 ( .A(n42229), .B(n42228), .Z(n42451) );
  NANDN U43074 ( .A(n42235), .B(n42234), .Z(n42239) );
  NANDN U43075 ( .A(n42237), .B(n42236), .Z(n42238) );
  NANDN U43076 ( .A(n42241), .B(n42240), .Z(n42245) );
  NAND U43077 ( .A(n42243), .B(n42242), .Z(n42244) );
  AND U43078 ( .A(n42245), .B(n42244), .Z(n42253) );
  NANDN U43079 ( .A(n42247), .B(n42246), .Z(n42251) );
  NANDN U43080 ( .A(n42249), .B(n42248), .Z(n42250) );
  NAND U43081 ( .A(n42251), .B(n42250), .Z(n42252) );
  XNOR U43082 ( .A(n42253), .B(n42252), .Z(n42429) );
  NANDN U43083 ( .A(n42255), .B(n42254), .Z(n42259) );
  NANDN U43084 ( .A(n42257), .B(n42256), .Z(n42258) );
  AND U43085 ( .A(n42259), .B(n42258), .Z(n42427) );
  NAND U43086 ( .A(n42261), .B(n42260), .Z(n42265) );
  NAND U43087 ( .A(n42263), .B(n42262), .Z(n42264) );
  AND U43088 ( .A(n42265), .B(n42264), .Z(n42337) );
  NAND U43089 ( .A(n42267), .B(n42266), .Z(n42270) );
  AND U43090 ( .A(x[502]), .B(y[8105]), .Z(n42303) );
  NAND U43091 ( .A(n42268), .B(n42303), .Z(n42269) );
  AND U43092 ( .A(n42270), .B(n42269), .Z(n42278) );
  NAND U43093 ( .A(n42272), .B(n42271), .Z(n42276) );
  NAND U43094 ( .A(n42274), .B(n42273), .Z(n42275) );
  NAND U43095 ( .A(n42276), .B(n42275), .Z(n42277) );
  XNOR U43096 ( .A(n42278), .B(n42277), .Z(n42335) );
  NAND U43097 ( .A(n42280), .B(n42279), .Z(n42283) );
  AND U43098 ( .A(x[490]), .B(y[8117]), .Z(n42298) );
  NAND U43099 ( .A(n42281), .B(n42298), .Z(n42282) );
  AND U43100 ( .A(n42283), .B(n42282), .Z(n42333) );
  AND U43101 ( .A(y[8101]), .B(x[506]), .Z(n42292) );
  AND U43102 ( .A(n42284), .B(o[446]), .Z(n42290) );
  XOR U43103 ( .A(n42285), .B(o[447]), .Z(n42288) );
  XNOR U43104 ( .A(n42286), .B(n42409), .Z(n42287) );
  XNOR U43105 ( .A(n42288), .B(n42287), .Z(n42289) );
  XNOR U43106 ( .A(n42290), .B(n42289), .Z(n42291) );
  XNOR U43107 ( .A(n42292), .B(n42291), .Z(n42331) );
  AND U43108 ( .A(y[8106]), .B(x[501]), .Z(n42294) );
  NAND U43109 ( .A(y[8119]), .B(x[488]), .Z(n42293) );
  XNOR U43110 ( .A(n42294), .B(n42293), .Z(n42302) );
  AND U43111 ( .A(y[8108]), .B(x[499]), .Z(n42300) );
  AND U43112 ( .A(y[8126]), .B(x[481]), .Z(n42296) );
  NAND U43113 ( .A(y[8099]), .B(x[508]), .Z(n42295) );
  XNOR U43114 ( .A(n42296), .B(n42295), .Z(n42297) );
  XNOR U43115 ( .A(n42298), .B(n42297), .Z(n42299) );
  XNOR U43116 ( .A(n42300), .B(n42299), .Z(n42301) );
  XOR U43117 ( .A(n42302), .B(n42301), .Z(n42305) );
  AND U43118 ( .A(x[505]), .B(y[8102]), .Z(n42400) );
  XNOR U43119 ( .A(n42303), .B(n42400), .Z(n42304) );
  XNOR U43120 ( .A(n42305), .B(n42304), .Z(n42321) );
  AND U43121 ( .A(y[8096]), .B(x[511]), .Z(n42307) );
  NAND U43122 ( .A(y[8124]), .B(x[483]), .Z(n42306) );
  XNOR U43123 ( .A(n42307), .B(n42306), .Z(n42311) );
  AND U43124 ( .A(y[8122]), .B(x[485]), .Z(n42309) );
  NAND U43125 ( .A(y[8123]), .B(x[484]), .Z(n42308) );
  XNOR U43126 ( .A(n42309), .B(n42308), .Z(n42310) );
  XOR U43127 ( .A(n42311), .B(n42310), .Z(n42319) );
  AND U43128 ( .A(y[8121]), .B(x[486]), .Z(n42313) );
  NAND U43129 ( .A(y[8125]), .B(x[482]), .Z(n42312) );
  XNOR U43130 ( .A(n42313), .B(n42312), .Z(n42317) );
  AND U43131 ( .A(y[8109]), .B(x[498]), .Z(n42315) );
  NAND U43132 ( .A(y[8110]), .B(x[497]), .Z(n42314) );
  XNOR U43133 ( .A(n42315), .B(n42314), .Z(n42316) );
  XNOR U43134 ( .A(n42317), .B(n42316), .Z(n42318) );
  XNOR U43135 ( .A(n42319), .B(n42318), .Z(n42320) );
  XOR U43136 ( .A(n42321), .B(n42320), .Z(n42329) );
  AND U43137 ( .A(y[8120]), .B(x[487]), .Z(n42323) );
  NAND U43138 ( .A(y[8118]), .B(x[489]), .Z(n42322) );
  XNOR U43139 ( .A(n42323), .B(n42322), .Z(n42327) );
  AND U43140 ( .A(y[8100]), .B(x[507]), .Z(n42325) );
  NAND U43141 ( .A(y[8104]), .B(x[503]), .Z(n42324) );
  XNOR U43142 ( .A(n42325), .B(n42324), .Z(n42326) );
  XNOR U43143 ( .A(n42327), .B(n42326), .Z(n42328) );
  XNOR U43144 ( .A(n42329), .B(n42328), .Z(n42330) );
  XNOR U43145 ( .A(n42331), .B(n42330), .Z(n42332) );
  XNOR U43146 ( .A(n42333), .B(n42332), .Z(n42334) );
  XNOR U43147 ( .A(n42335), .B(n42334), .Z(n42336) );
  XNOR U43148 ( .A(n42337), .B(n42336), .Z(n42425) );
  NAND U43149 ( .A(n42339), .B(n42338), .Z(n42343) );
  NAND U43150 ( .A(n42341), .B(n42340), .Z(n42342) );
  AND U43151 ( .A(n42343), .B(n42342), .Z(n42375) );
  NAND U43152 ( .A(n42345), .B(n42344), .Z(n42349) );
  NAND U43153 ( .A(n42347), .B(n42346), .Z(n42348) );
  AND U43154 ( .A(n42349), .B(n42348), .Z(n42357) );
  NAND U43155 ( .A(n42351), .B(n42350), .Z(n42355) );
  NAND U43156 ( .A(n42353), .B(n42352), .Z(n42354) );
  NAND U43157 ( .A(n42355), .B(n42354), .Z(n42356) );
  XNOR U43158 ( .A(n42357), .B(n42356), .Z(n42373) );
  AND U43159 ( .A(y[8116]), .B(x[491]), .Z(n42359) );
  NAND U43160 ( .A(y[8127]), .B(x[480]), .Z(n42358) );
  XNOR U43161 ( .A(n42359), .B(n42358), .Z(n42363) );
  AND U43162 ( .A(y[8111]), .B(x[496]), .Z(n42361) );
  NAND U43163 ( .A(y[8107]), .B(x[500]), .Z(n42360) );
  XNOR U43164 ( .A(n42361), .B(n42360), .Z(n42362) );
  XOR U43165 ( .A(n42363), .B(n42362), .Z(n42371) );
  AND U43166 ( .A(y[8098]), .B(x[509]), .Z(n42365) );
  NAND U43167 ( .A(y[8115]), .B(x[492]), .Z(n42364) );
  XNOR U43168 ( .A(n42365), .B(n42364), .Z(n42369) );
  AND U43169 ( .A(y[8097]), .B(x[510]), .Z(n42367) );
  NAND U43170 ( .A(y[8113]), .B(x[494]), .Z(n42366) );
  XNOR U43171 ( .A(n42367), .B(n42366), .Z(n42368) );
  XNOR U43172 ( .A(n42369), .B(n42368), .Z(n42370) );
  XNOR U43173 ( .A(n42371), .B(n42370), .Z(n42372) );
  XNOR U43174 ( .A(n42373), .B(n42372), .Z(n42374) );
  XNOR U43175 ( .A(n42375), .B(n42374), .Z(n42391) );
  NAND U43176 ( .A(n42377), .B(n42376), .Z(n42381) );
  ANDN U43177 ( .B(n42379), .A(n42378), .Z(n42380) );
  ANDN U43178 ( .B(n42381), .A(n42380), .Z(n42389) );
  AND U43179 ( .A(n42383), .B(n42382), .Z(n42387) );
  ANDN U43180 ( .B(n42385), .A(n42384), .Z(n42386) );
  OR U43181 ( .A(n42387), .B(n42386), .Z(n42388) );
  XNOR U43182 ( .A(n42389), .B(n42388), .Z(n42390) );
  XOR U43183 ( .A(n42391), .B(n42390), .Z(n42423) );
  NAND U43184 ( .A(n42393), .B(n42392), .Z(n42397) );
  NAND U43185 ( .A(n42395), .B(n42394), .Z(n42396) );
  AND U43186 ( .A(n42397), .B(n42396), .Z(n42405) );
  NAND U43187 ( .A(n42399), .B(n42398), .Z(n42403) );
  NAND U43188 ( .A(n42401), .B(n42400), .Z(n42402) );
  NAND U43189 ( .A(n42403), .B(n42402), .Z(n42404) );
  XNOR U43190 ( .A(n42405), .B(n42404), .Z(n42421) );
  NAND U43191 ( .A(n42407), .B(n42406), .Z(n42411) );
  NAND U43192 ( .A(n42409), .B(n42408), .Z(n42410) );
  AND U43193 ( .A(n42411), .B(n42410), .Z(n42419) );
  NAND U43194 ( .A(n42413), .B(n42412), .Z(n42417) );
  NAND U43195 ( .A(n42415), .B(n42414), .Z(n42416) );
  NAND U43196 ( .A(n42417), .B(n42416), .Z(n42418) );
  XNOR U43197 ( .A(n42419), .B(n42418), .Z(n42420) );
  XNOR U43198 ( .A(n42421), .B(n42420), .Z(n42422) );
  XNOR U43199 ( .A(n42423), .B(n42422), .Z(n42424) );
  XNOR U43200 ( .A(n42425), .B(n42424), .Z(n42426) );
  XNOR U43201 ( .A(n42427), .B(n42426), .Z(n42428) );
  NAND U43202 ( .A(n42431), .B(n42430), .Z(n42435) );
  NAND U43203 ( .A(n42433), .B(n42432), .Z(n42434) );
  NAND U43204 ( .A(n42437), .B(n42436), .Z(n42441) );
  NANDN U43205 ( .A(n42439), .B(n42438), .Z(n42440) );
  XNOR U43206 ( .A(n42451), .B(n42450), .Z(n42467) );
  NAND U43207 ( .A(n42453), .B(n42452), .Z(n42457) );
  NANDN U43208 ( .A(n42455), .B(n42454), .Z(n42456) );
  AND U43209 ( .A(n42457), .B(n42456), .Z(n42465) );
  NANDN U43210 ( .A(n42459), .B(n42458), .Z(n42463) );
  NANDN U43211 ( .A(n42461), .B(n42460), .Z(n42462) );
  NAND U43212 ( .A(n42463), .B(n42462), .Z(n42464) );
  XNOR U43213 ( .A(n42465), .B(n42464), .Z(n42466) );
  XNOR U43214 ( .A(n42467), .B(n42466), .Z(n42468) );
  XNOR U43215 ( .A(n42469), .B(n42468), .Z(n42485) );
  NANDN U43216 ( .A(n42471), .B(n42470), .Z(n42475) );
  NANDN U43217 ( .A(n42473), .B(n42472), .Z(n42474) );
  AND U43218 ( .A(n42475), .B(n42474), .Z(n42483) );
  NAND U43219 ( .A(n42477), .B(n42476), .Z(n42481) );
  NANDN U43220 ( .A(n42479), .B(n42478), .Z(n42480) );
  NAND U43221 ( .A(n42481), .B(n42480), .Z(n42482) );
  XNOR U43222 ( .A(n42483), .B(n42482), .Z(n42484) );
  XNOR U43223 ( .A(n42485), .B(n42484), .Z(n42486) );
  XNOR U43224 ( .A(n42487), .B(n42486), .Z(n42495) );
  ANDN U43225 ( .B(n42489), .A(n42488), .Z(n42493) );
  AND U43226 ( .A(n42491), .B(n42490), .Z(n42492) );
  NOR U43227 ( .A(n42493), .B(n42492), .Z(n42494) );
  XNOR U43228 ( .A(n42495), .B(n42494), .Z(N896) );
  AND U43229 ( .A(x[480]), .B(y[8128]), .Z(n43131) );
  XOR U43230 ( .A(n43131), .B(o[448]), .Z(N929) );
  AND U43231 ( .A(x[481]), .B(y[8128]), .Z(n42504) );
  AND U43232 ( .A(x[480]), .B(y[8129]), .Z(n42503) );
  XNOR U43233 ( .A(n42503), .B(o[449]), .Z(n42496) );
  XNOR U43234 ( .A(n42504), .B(n42496), .Z(n42498) );
  NAND U43235 ( .A(n43131), .B(o[448]), .Z(n42497) );
  XNOR U43236 ( .A(n42498), .B(n42497), .Z(N930) );
  NANDN U43237 ( .A(n42504), .B(n42496), .Z(n42500) );
  NAND U43238 ( .A(n42498), .B(n42497), .Z(n42499) );
  AND U43239 ( .A(n42500), .B(n42499), .Z(n42510) );
  AND U43240 ( .A(x[480]), .B(y[8130]), .Z(n42517) );
  XNOR U43241 ( .A(n42517), .B(o[450]), .Z(n42509) );
  XNOR U43242 ( .A(n42510), .B(n42509), .Z(n42512) );
  AND U43243 ( .A(y[8128]), .B(x[482]), .Z(n42502) );
  NAND U43244 ( .A(y[8129]), .B(x[481]), .Z(n42501) );
  XNOR U43245 ( .A(n42502), .B(n42501), .Z(n42506) );
  AND U43246 ( .A(n42503), .B(o[449]), .Z(n42505) );
  XNOR U43247 ( .A(n42506), .B(n42505), .Z(n42511) );
  XNOR U43248 ( .A(n42512), .B(n42511), .Z(N931) );
  AND U43249 ( .A(x[482]), .B(y[8129]), .Z(n42524) );
  NAND U43250 ( .A(n42524), .B(n42504), .Z(n42508) );
  NAND U43251 ( .A(n42506), .B(n42505), .Z(n42507) );
  AND U43252 ( .A(n42508), .B(n42507), .Z(n42527) );
  NANDN U43253 ( .A(n42510), .B(n42509), .Z(n42514) );
  NAND U43254 ( .A(n42512), .B(n42511), .Z(n42513) );
  AND U43255 ( .A(n42514), .B(n42513), .Z(n42526) );
  XNOR U43256 ( .A(n42527), .B(n42526), .Z(n42529) );
  AND U43257 ( .A(x[481]), .B(y[8130]), .Z(n42633) );
  XOR U43258 ( .A(n42524), .B(o[451]), .Z(n42532) );
  XOR U43259 ( .A(n42633), .B(n42532), .Z(n42534) );
  AND U43260 ( .A(y[8128]), .B(x[483]), .Z(n42516) );
  NAND U43261 ( .A(y[8131]), .B(x[480]), .Z(n42515) );
  XNOR U43262 ( .A(n42516), .B(n42515), .Z(n42519) );
  AND U43263 ( .A(n42517), .B(o[450]), .Z(n42518) );
  XOR U43264 ( .A(n42519), .B(n42518), .Z(n42533) );
  XOR U43265 ( .A(n42534), .B(n42533), .Z(n42528) );
  XOR U43266 ( .A(n42529), .B(n42528), .Z(N932) );
  AND U43267 ( .A(x[483]), .B(y[8131]), .Z(n42577) );
  NAND U43268 ( .A(n43131), .B(n42577), .Z(n42521) );
  NAND U43269 ( .A(n42519), .B(n42518), .Z(n42520) );
  NAND U43270 ( .A(n42521), .B(n42520), .Z(n42555) );
  AND U43271 ( .A(y[8132]), .B(x[480]), .Z(n42523) );
  NAND U43272 ( .A(y[8128]), .B(x[484]), .Z(n42522) );
  XNOR U43273 ( .A(n42523), .B(n42522), .Z(n42548) );
  AND U43274 ( .A(n42524), .B(o[451]), .Z(n42549) );
  XOR U43275 ( .A(n42548), .B(n42549), .Z(n42553) );
  AND U43276 ( .A(y[8130]), .B(x[482]), .Z(n42687) );
  NAND U43277 ( .A(y[8131]), .B(x[481]), .Z(n42525) );
  XNOR U43278 ( .A(n42687), .B(n42525), .Z(n42545) );
  AND U43279 ( .A(x[483]), .B(y[8129]), .Z(n42540) );
  XOR U43280 ( .A(o[452]), .B(n42540), .Z(n42544) );
  XOR U43281 ( .A(n42545), .B(n42544), .Z(n42552) );
  XOR U43282 ( .A(n42553), .B(n42552), .Z(n42554) );
  XOR U43283 ( .A(n42555), .B(n42554), .Z(n42559) );
  NANDN U43284 ( .A(n42527), .B(n42526), .Z(n42531) );
  NAND U43285 ( .A(n42529), .B(n42528), .Z(n42530) );
  NAND U43286 ( .A(n42531), .B(n42530), .Z(n42560) );
  NAND U43287 ( .A(n42633), .B(n42532), .Z(n42536) );
  NAND U43288 ( .A(n42534), .B(n42533), .Z(n42535) );
  NAND U43289 ( .A(n42536), .B(n42535), .Z(n42561) );
  IV U43290 ( .A(n42561), .Z(n42558) );
  XOR U43291 ( .A(n42560), .B(n42558), .Z(n42537) );
  XNOR U43292 ( .A(n42559), .B(n42537), .Z(N933) );
  AND U43293 ( .A(y[8128]), .B(x[485]), .Z(n42539) );
  NAND U43294 ( .A(y[8133]), .B(x[480]), .Z(n42538) );
  XNOR U43295 ( .A(n42539), .B(n42538), .Z(n42570) );
  AND U43296 ( .A(o[452]), .B(n42540), .Z(n42569) );
  XOR U43297 ( .A(n42570), .B(n42569), .Z(n42568) );
  NAND U43298 ( .A(x[482]), .B(y[8131]), .Z(n42640) );
  AND U43299 ( .A(y[8130]), .B(x[483]), .Z(n42542) );
  NAND U43300 ( .A(y[8132]), .B(x[481]), .Z(n42541) );
  XNOR U43301 ( .A(n42542), .B(n42541), .Z(n42564) );
  AND U43302 ( .A(x[484]), .B(y[8129]), .Z(n42575) );
  XOR U43303 ( .A(n42575), .B(o[453]), .Z(n42563) );
  XOR U43304 ( .A(n42564), .B(n42563), .Z(n42567) );
  XOR U43305 ( .A(n42640), .B(n42567), .Z(n42543) );
  XNOR U43306 ( .A(n42568), .B(n42543), .Z(n42585) );
  NANDN U43307 ( .A(n42640), .B(n42633), .Z(n42547) );
  NAND U43308 ( .A(n42545), .B(n42544), .Z(n42546) );
  NAND U43309 ( .A(n42547), .B(n42546), .Z(n42583) );
  AND U43310 ( .A(x[484]), .B(y[8132]), .Z(n43318) );
  NAND U43311 ( .A(n43318), .B(n43131), .Z(n42551) );
  NAND U43312 ( .A(n42549), .B(n42548), .Z(n42550) );
  NAND U43313 ( .A(n42551), .B(n42550), .Z(n42582) );
  XOR U43314 ( .A(n42583), .B(n42582), .Z(n42584) );
  XNOR U43315 ( .A(n42585), .B(n42584), .Z(n42581) );
  NAND U43316 ( .A(n42553), .B(n42552), .Z(n42557) );
  NAND U43317 ( .A(n42555), .B(n42554), .Z(n42556) );
  NAND U43318 ( .A(n42557), .B(n42556), .Z(n42580) );
  XOR U43319 ( .A(n42580), .B(n42579), .Z(n42562) );
  XNOR U43320 ( .A(n42581), .B(n42562), .Z(N934) );
  AND U43321 ( .A(x[483]), .B(y[8132]), .Z(n42641) );
  NAND U43322 ( .A(n42641), .B(n42633), .Z(n42566) );
  NAND U43323 ( .A(n42564), .B(n42563), .Z(n42565) );
  NAND U43324 ( .A(n42566), .B(n42565), .Z(n42614) );
  XOR U43325 ( .A(n42614), .B(n42613), .Z(n42616) );
  AND U43326 ( .A(x[485]), .B(y[8133]), .Z(n42811) );
  NAND U43327 ( .A(n43131), .B(n42811), .Z(n42572) );
  NAND U43328 ( .A(n42570), .B(n42569), .Z(n42571) );
  NAND U43329 ( .A(n42572), .B(n42571), .Z(n42590) );
  AND U43330 ( .A(y[8128]), .B(x[486]), .Z(n42574) );
  NAND U43331 ( .A(y[8134]), .B(x[480]), .Z(n42573) );
  XNOR U43332 ( .A(n42574), .B(n42573), .Z(n42596) );
  AND U43333 ( .A(n42575), .B(o[453]), .Z(n42597) );
  XOR U43334 ( .A(n42596), .B(n42597), .Z(n42589) );
  XOR U43335 ( .A(n42590), .B(n42589), .Z(n42592) );
  NAND U43336 ( .A(y[8132]), .B(x[482]), .Z(n42576) );
  XNOR U43337 ( .A(n42577), .B(n42576), .Z(n42601) );
  AND U43338 ( .A(y[8133]), .B(x[481]), .Z(n42852) );
  NAND U43339 ( .A(y[8130]), .B(x[484]), .Z(n42578) );
  XNOR U43340 ( .A(n42852), .B(n42578), .Z(n42605) );
  AND U43341 ( .A(x[485]), .B(y[8129]), .Z(n42612) );
  XOR U43342 ( .A(o[454]), .B(n42612), .Z(n42604) );
  XOR U43343 ( .A(n42605), .B(n42604), .Z(n42600) );
  XOR U43344 ( .A(n42601), .B(n42600), .Z(n42591) );
  XOR U43345 ( .A(n42592), .B(n42591), .Z(n42615) );
  XOR U43346 ( .A(n42616), .B(n42615), .Z(n42622) );
  NAND U43347 ( .A(n42583), .B(n42582), .Z(n42587) );
  NAND U43348 ( .A(n42585), .B(n42584), .Z(n42586) );
  AND U43349 ( .A(n42587), .B(n42586), .Z(n42621) );
  IV U43350 ( .A(n42621), .Z(n42619) );
  XOR U43351 ( .A(n42620), .B(n42619), .Z(n42588) );
  XNOR U43352 ( .A(n42622), .B(n42588), .Z(N935) );
  NAND U43353 ( .A(n42590), .B(n42589), .Z(n42594) );
  NAND U43354 ( .A(n42592), .B(n42591), .Z(n42593) );
  AND U43355 ( .A(n42594), .B(n42593), .Z(n42663) );
  AND U43356 ( .A(y[8130]), .B(x[485]), .Z(n42723) );
  NAND U43357 ( .A(y[8134]), .B(x[481]), .Z(n42595) );
  XNOR U43358 ( .A(n42723), .B(n42595), .Z(n42635) );
  AND U43359 ( .A(x[486]), .B(y[8129]), .Z(n42638) );
  XOR U43360 ( .A(o[455]), .B(n42638), .Z(n42634) );
  XOR U43361 ( .A(n42635), .B(n42634), .Z(n42652) );
  AND U43362 ( .A(x[486]), .B(y[8134]), .Z(n42870) );
  NAND U43363 ( .A(n43131), .B(n42870), .Z(n42599) );
  NAND U43364 ( .A(n42597), .B(n42596), .Z(n42598) );
  AND U43365 ( .A(n42599), .B(n42598), .Z(n42651) );
  NANDN U43366 ( .A(n42640), .B(n42641), .Z(n42603) );
  NAND U43367 ( .A(n42601), .B(n42600), .Z(n42602) );
  NAND U43368 ( .A(n42603), .B(n42602), .Z(n42654) );
  AND U43369 ( .A(x[484]), .B(y[8133]), .Z(n43136) );
  NAND U43370 ( .A(n43136), .B(n42633), .Z(n42607) );
  NAND U43371 ( .A(n42605), .B(n42604), .Z(n42606) );
  AND U43372 ( .A(n42607), .B(n42606), .Z(n42630) );
  AND U43373 ( .A(y[8133]), .B(x[482]), .Z(n42609) );
  NAND U43374 ( .A(y[8131]), .B(x[484]), .Z(n42608) );
  XNOR U43375 ( .A(n42609), .B(n42608), .Z(n42642) );
  XNOR U43376 ( .A(n42642), .B(n42641), .Z(n42628) );
  AND U43377 ( .A(y[8128]), .B(x[487]), .Z(n42611) );
  NAND U43378 ( .A(y[8135]), .B(x[480]), .Z(n42610) );
  XNOR U43379 ( .A(n42611), .B(n42610), .Z(n42646) );
  AND U43380 ( .A(o[454]), .B(n42612), .Z(n42645) );
  XNOR U43381 ( .A(n42646), .B(n42645), .Z(n42627) );
  XOR U43382 ( .A(n42628), .B(n42627), .Z(n42629) );
  XOR U43383 ( .A(n42630), .B(n42629), .Z(n42660) );
  XOR U43384 ( .A(n42661), .B(n42660), .Z(n42662) );
  XOR U43385 ( .A(n42663), .B(n42662), .Z(n42659) );
  NAND U43386 ( .A(n42614), .B(n42613), .Z(n42618) );
  NAND U43387 ( .A(n42616), .B(n42615), .Z(n42617) );
  NAND U43388 ( .A(n42618), .B(n42617), .Z(n42658) );
  NANDN U43389 ( .A(n42619), .B(n42620), .Z(n42625) );
  NOR U43390 ( .A(n42621), .B(n42620), .Z(n42623) );
  OR U43391 ( .A(n42623), .B(n42622), .Z(n42624) );
  AND U43392 ( .A(n42625), .B(n42624), .Z(n42657) );
  XOR U43393 ( .A(n42658), .B(n42657), .Z(n42626) );
  XNOR U43394 ( .A(n42659), .B(n42626), .Z(N936) );
  NAND U43395 ( .A(n42628), .B(n42627), .Z(n42632) );
  NAND U43396 ( .A(n42630), .B(n42629), .Z(n42631) );
  AND U43397 ( .A(n42632), .B(n42631), .Z(n42700) );
  AND U43398 ( .A(x[485]), .B(y[8134]), .Z(n42803) );
  NAND U43399 ( .A(n42803), .B(n42633), .Z(n42637) );
  NAND U43400 ( .A(n42635), .B(n42634), .Z(n42636) );
  NAND U43401 ( .A(n42637), .B(n42636), .Z(n42698) );
  AND U43402 ( .A(n42638), .B(o[455]), .Z(n42679) );
  AND U43403 ( .A(y[8131]), .B(x[485]), .Z(n43231) );
  AND U43404 ( .A(y[8135]), .B(x[481]), .Z(n43126) );
  XOR U43405 ( .A(n43231), .B(n43126), .Z(n42678) );
  XNOR U43406 ( .A(n42679), .B(n42678), .Z(n42683) );
  AND U43407 ( .A(x[483]), .B(y[8133]), .Z(n43463) );
  AND U43408 ( .A(x[486]), .B(y[8130]), .Z(n42639) );
  AND U43409 ( .A(y[8134]), .B(x[482]), .Z(n43541) );
  XOR U43410 ( .A(n42639), .B(n43541), .Z(n42688) );
  XNOR U43411 ( .A(n43318), .B(n42688), .Z(n42682) );
  XOR U43412 ( .A(n43463), .B(n42682), .Z(n42684) );
  XOR U43413 ( .A(n42683), .B(n42684), .Z(n42697) );
  XOR U43414 ( .A(n42698), .B(n42697), .Z(n42699) );
  XOR U43415 ( .A(n42700), .B(n42699), .Z(n42706) );
  NANDN U43416 ( .A(n42640), .B(n43136), .Z(n42644) );
  NAND U43417 ( .A(n42642), .B(n42641), .Z(n42643) );
  NAND U43418 ( .A(n42644), .B(n42643), .Z(n42694) );
  AND U43419 ( .A(x[487]), .B(y[8135]), .Z(n43018) );
  NAND U43420 ( .A(n43131), .B(n43018), .Z(n42648) );
  NAND U43421 ( .A(n42646), .B(n42645), .Z(n42647) );
  NAND U43422 ( .A(n42648), .B(n42647), .Z(n42692) );
  AND U43423 ( .A(y[8128]), .B(x[488]), .Z(n42650) );
  NAND U43424 ( .A(y[8136]), .B(x[480]), .Z(n42649) );
  XNOR U43425 ( .A(n42650), .B(n42649), .Z(n42669) );
  AND U43426 ( .A(x[487]), .B(y[8129]), .Z(n42674) );
  XOR U43427 ( .A(n42674), .B(o[456]), .Z(n42668) );
  XOR U43428 ( .A(n42669), .B(n42668), .Z(n42691) );
  XOR U43429 ( .A(n42692), .B(n42691), .Z(n42693) );
  XNOR U43430 ( .A(n42694), .B(n42693), .Z(n42704) );
  NANDN U43431 ( .A(n42652), .B(n42651), .Z(n42656) );
  NANDN U43432 ( .A(n42654), .B(n42653), .Z(n42655) );
  NAND U43433 ( .A(n42656), .B(n42655), .Z(n42703) );
  XOR U43434 ( .A(n42704), .B(n42703), .Z(n42705) );
  XOR U43435 ( .A(n42706), .B(n42705), .Z(n42712) );
  NAND U43436 ( .A(n42661), .B(n42660), .Z(n42665) );
  NAND U43437 ( .A(n42663), .B(n42662), .Z(n42664) );
  NAND U43438 ( .A(n42665), .B(n42664), .Z(n42711) );
  IV U43439 ( .A(n42711), .Z(n42709) );
  XOR U43440 ( .A(n42710), .B(n42709), .Z(n42666) );
  XNOR U43441 ( .A(n42712), .B(n42666), .Z(N937) );
  AND U43442 ( .A(x[488]), .B(y[8136]), .Z(n42667) );
  NAND U43443 ( .A(n42667), .B(n43131), .Z(n42671) );
  NAND U43444 ( .A(n42669), .B(n42668), .Z(n42670) );
  AND U43445 ( .A(n42671), .B(n42670), .Z(n42751) );
  AND U43446 ( .A(y[8132]), .B(x[485]), .Z(n42673) );
  NAND U43447 ( .A(y[8130]), .B(x[487]), .Z(n42672) );
  XNOR U43448 ( .A(n42673), .B(n42672), .Z(n42724) );
  NAND U43449 ( .A(n42674), .B(o[456]), .Z(n42725) );
  XOR U43450 ( .A(n42724), .B(n42725), .Z(n42749) );
  AND U43451 ( .A(y[8128]), .B(x[489]), .Z(n42676) );
  NAND U43452 ( .A(y[8137]), .B(x[480]), .Z(n42675) );
  XNOR U43453 ( .A(n42676), .B(n42675), .Z(n42732) );
  AND U43454 ( .A(x[488]), .B(y[8129]), .Z(n42741) );
  XOR U43455 ( .A(n42741), .B(o[457]), .Z(n42731) );
  XNOR U43456 ( .A(n42732), .B(n42731), .Z(n42750) );
  XNOR U43457 ( .A(n42749), .B(n42750), .Z(n42752) );
  XOR U43458 ( .A(n42751), .B(n42752), .Z(n42746) );
  AND U43459 ( .A(y[8131]), .B(x[486]), .Z(n43081) );
  NAND U43460 ( .A(y[8136]), .B(x[481]), .Z(n42677) );
  XOR U43461 ( .A(n43081), .B(n42677), .Z(n42736) );
  XOR U43462 ( .A(n43136), .B(n42736), .Z(n42755) );
  NAND U43463 ( .A(x[482]), .B(y[8135]), .Z(n43283) );
  NAND U43464 ( .A(x[483]), .B(y[8134]), .Z(n43089) );
  XOR U43465 ( .A(n43283), .B(n43089), .Z(n42756) );
  XNOR U43466 ( .A(n42755), .B(n42756), .Z(n42744) );
  NAND U43467 ( .A(x[485]), .B(y[8135]), .Z(n42931) );
  AND U43468 ( .A(x[481]), .B(y[8131]), .Z(n42735) );
  NANDN U43469 ( .A(n42931), .B(n42735), .Z(n42681) );
  NAND U43470 ( .A(n42679), .B(n42678), .Z(n42680) );
  NAND U43471 ( .A(n42681), .B(n42680), .Z(n42743) );
  XOR U43472 ( .A(n42744), .B(n42743), .Z(n42745) );
  XNOR U43473 ( .A(n42746), .B(n42745), .Z(n42719) );
  NANDN U43474 ( .A(n43463), .B(n42682), .Z(n42686) );
  NANDN U43475 ( .A(n42684), .B(n42683), .Z(n42685) );
  NAND U43476 ( .A(n42686), .B(n42685), .Z(n42717) );
  NAND U43477 ( .A(n42870), .B(n42687), .Z(n42690) );
  NAND U43478 ( .A(n43318), .B(n42688), .Z(n42689) );
  AND U43479 ( .A(n42690), .B(n42689), .Z(n42718) );
  XNOR U43480 ( .A(n42717), .B(n42718), .Z(n42720) );
  NAND U43481 ( .A(n42692), .B(n42691), .Z(n42696) );
  NAND U43482 ( .A(n42694), .B(n42693), .Z(n42695) );
  NAND U43483 ( .A(n42696), .B(n42695), .Z(n42760) );
  NAND U43484 ( .A(n42698), .B(n42697), .Z(n42702) );
  NAND U43485 ( .A(n42700), .B(n42699), .Z(n42701) );
  NAND U43486 ( .A(n42702), .B(n42701), .Z(n42759) );
  XOR U43487 ( .A(n42760), .B(n42759), .Z(n42762) );
  XOR U43488 ( .A(n42761), .B(n42762), .Z(n42767) );
  NAND U43489 ( .A(n42704), .B(n42703), .Z(n42708) );
  NANDN U43490 ( .A(n42706), .B(n42705), .Z(n42707) );
  NAND U43491 ( .A(n42708), .B(n42707), .Z(n42765) );
  NANDN U43492 ( .A(n42709), .B(n42710), .Z(n42715) );
  NOR U43493 ( .A(n42711), .B(n42710), .Z(n42713) );
  OR U43494 ( .A(n42713), .B(n42712), .Z(n42714) );
  AND U43495 ( .A(n42715), .B(n42714), .Z(n42766) );
  XOR U43496 ( .A(n42765), .B(n42766), .Z(n42716) );
  XNOR U43497 ( .A(n42767), .B(n42716), .Z(N938) );
  NAND U43498 ( .A(n42718), .B(n42717), .Z(n42722) );
  NANDN U43499 ( .A(n42720), .B(n42719), .Z(n42721) );
  NAND U43500 ( .A(n42722), .B(n42721), .Z(n42824) );
  AND U43501 ( .A(x[487]), .B(y[8132]), .Z(n42805) );
  NAND U43502 ( .A(n42805), .B(n42723), .Z(n42727) );
  NANDN U43503 ( .A(n42725), .B(n42724), .Z(n42726) );
  AND U43504 ( .A(n42727), .B(n42726), .Z(n42815) );
  AND U43505 ( .A(y[8131]), .B(x[487]), .Z(n42729) );
  NAND U43506 ( .A(y[8134]), .B(x[484]), .Z(n42728) );
  XNOR U43507 ( .A(n42729), .B(n42728), .Z(n42789) );
  AND U43508 ( .A(x[486]), .B(y[8132]), .Z(n42788) );
  XOR U43509 ( .A(n42789), .B(n42788), .Z(n42814) );
  AND U43510 ( .A(x[488]), .B(y[8130]), .Z(n42991) );
  AND U43511 ( .A(x[489]), .B(y[8129]), .Z(n42799) );
  XOR U43512 ( .A(o[458]), .B(n42799), .Z(n42810) );
  XOR U43513 ( .A(n42991), .B(n42810), .Z(n42812) );
  XNOR U43514 ( .A(n42812), .B(n42811), .Z(n42813) );
  XOR U43515 ( .A(n42814), .B(n42813), .Z(n42816) );
  XOR U43516 ( .A(n42815), .B(n42816), .Z(n42777) );
  AND U43517 ( .A(x[489]), .B(y[8137]), .Z(n42730) );
  NAND U43518 ( .A(n42730), .B(n43131), .Z(n42734) );
  NAND U43519 ( .A(n42732), .B(n42731), .Z(n42733) );
  NAND U43520 ( .A(n42734), .B(n42733), .Z(n42775) );
  AND U43521 ( .A(x[486]), .B(y[8136]), .Z(n43028) );
  NAND U43522 ( .A(n43028), .B(n42735), .Z(n42738) );
  NANDN U43523 ( .A(n42736), .B(n43136), .Z(n42737) );
  AND U43524 ( .A(n42738), .B(n42737), .Z(n42784) );
  AND U43525 ( .A(y[8128]), .B(x[490]), .Z(n42740) );
  NAND U43526 ( .A(y[8138]), .B(x[480]), .Z(n42739) );
  XNOR U43527 ( .A(n42740), .B(n42739), .Z(n42794) );
  AND U43528 ( .A(n42741), .B(o[457]), .Z(n42793) );
  XOR U43529 ( .A(n42794), .B(n42793), .Z(n42781) );
  AND U43530 ( .A(y[8135]), .B(x[483]), .Z(n43687) );
  NAND U43531 ( .A(y[8137]), .B(x[481]), .Z(n42742) );
  XNOR U43532 ( .A(n43687), .B(n42742), .Z(n42806) );
  NAND U43533 ( .A(x[482]), .B(y[8136]), .Z(n42807) );
  XOR U43534 ( .A(n42806), .B(n42807), .Z(n42782) );
  XNOR U43535 ( .A(n42781), .B(n42782), .Z(n42783) );
  XNOR U43536 ( .A(n42784), .B(n42783), .Z(n42776) );
  XOR U43537 ( .A(n42775), .B(n42776), .Z(n42778) );
  XOR U43538 ( .A(n42777), .B(n42778), .Z(n42823) );
  NAND U43539 ( .A(n42744), .B(n42743), .Z(n42748) );
  NAND U43540 ( .A(n42746), .B(n42745), .Z(n42747) );
  NAND U43541 ( .A(n42748), .B(n42747), .Z(n42771) );
  NAND U43542 ( .A(n42750), .B(n42749), .Z(n42754) );
  NANDN U43543 ( .A(n42752), .B(n42751), .Z(n42753) );
  AND U43544 ( .A(n42754), .B(n42753), .Z(n42770) );
  NAND U43545 ( .A(n42756), .B(n42755), .Z(n42758) );
  IV U43546 ( .A(n43283), .Z(n43365) );
  ANDN U43547 ( .B(n43089), .A(n43365), .Z(n42757) );
  ANDN U43548 ( .B(n42758), .A(n42757), .Z(n42769) );
  XOR U43549 ( .A(n42770), .B(n42769), .Z(n42772) );
  XNOR U43550 ( .A(n42771), .B(n42772), .Z(n42822) );
  XOR U43551 ( .A(n42824), .B(n42825), .Z(n42821) );
  NAND U43552 ( .A(n42760), .B(n42759), .Z(n42764) );
  NAND U43553 ( .A(n42762), .B(n42761), .Z(n42763) );
  NAND U43554 ( .A(n42764), .B(n42763), .Z(n42820) );
  XOR U43555 ( .A(n42820), .B(n42819), .Z(n42768) );
  XNOR U43556 ( .A(n42821), .B(n42768), .Z(N939) );
  NAND U43557 ( .A(n42770), .B(n42769), .Z(n42774) );
  NAND U43558 ( .A(n42772), .B(n42771), .Z(n42773) );
  NAND U43559 ( .A(n42774), .B(n42773), .Z(n42831) );
  NAND U43560 ( .A(n42776), .B(n42775), .Z(n42780) );
  NAND U43561 ( .A(n42778), .B(n42777), .Z(n42779) );
  NAND U43562 ( .A(n42780), .B(n42779), .Z(n42829) );
  NANDN U43563 ( .A(n42782), .B(n42781), .Z(n42786) );
  NANDN U43564 ( .A(n42784), .B(n42783), .Z(n42785) );
  NAND U43565 ( .A(n42786), .B(n42785), .Z(n42891) );
  AND U43566 ( .A(x[487]), .B(y[8134]), .Z(n42926) );
  AND U43567 ( .A(x[484]), .B(y[8131]), .Z(n42787) );
  NAND U43568 ( .A(n42926), .B(n42787), .Z(n42791) );
  NAND U43569 ( .A(n42789), .B(n42788), .Z(n42790) );
  NAND U43570 ( .A(n42791), .B(n42790), .Z(n42889) );
  AND U43571 ( .A(x[490]), .B(y[8138]), .Z(n42792) );
  NAND U43572 ( .A(n42792), .B(n43131), .Z(n42796) );
  NAND U43573 ( .A(n42794), .B(n42793), .Z(n42795) );
  NAND U43574 ( .A(n42796), .B(n42795), .Z(n42885) );
  AND U43575 ( .A(y[8128]), .B(x[491]), .Z(n42798) );
  NAND U43576 ( .A(y[8139]), .B(x[480]), .Z(n42797) );
  XNOR U43577 ( .A(n42798), .B(n42797), .Z(n42860) );
  AND U43578 ( .A(o[458]), .B(n42799), .Z(n42861) );
  XOR U43579 ( .A(n42860), .B(n42861), .Z(n42884) );
  AND U43580 ( .A(y[8133]), .B(x[486]), .Z(n42801) );
  NAND U43581 ( .A(y[8138]), .B(x[481]), .Z(n42800) );
  XNOR U43582 ( .A(n42801), .B(n42800), .Z(n42854) );
  AND U43583 ( .A(x[490]), .B(y[8129]), .Z(n42871) );
  XOR U43584 ( .A(o[459]), .B(n42871), .Z(n42853) );
  XOR U43585 ( .A(n42854), .B(n42853), .Z(n42883) );
  XOR U43586 ( .A(n42884), .B(n42883), .Z(n42886) );
  XNOR U43587 ( .A(n42885), .B(n42886), .Z(n42890) );
  XOR U43588 ( .A(n42891), .B(n42892), .Z(n42875) );
  NAND U43589 ( .A(x[483]), .B(y[8136]), .Z(n43816) );
  NAND U43590 ( .A(y[8137]), .B(x[482]), .Z(n42802) );
  XNOR U43591 ( .A(n42803), .B(n42802), .Z(n42849) );
  AND U43592 ( .A(x[484]), .B(y[8135]), .Z(n42848) );
  XNOR U43593 ( .A(n42849), .B(n42848), .Z(n42878) );
  XOR U43594 ( .A(n43816), .B(n42878), .Z(n42880) );
  NAND U43595 ( .A(y[8130]), .B(x[489]), .Z(n42804) );
  XNOR U43596 ( .A(n42805), .B(n42804), .Z(n42866) );
  AND U43597 ( .A(x[488]), .B(y[8131]), .Z(n42865) );
  XNOR U43598 ( .A(n42866), .B(n42865), .Z(n42879) );
  XOR U43599 ( .A(n42880), .B(n42879), .Z(n42844) );
  NAND U43600 ( .A(x[483]), .B(y[8137]), .Z(n42922) );
  NANDN U43601 ( .A(n42922), .B(n43126), .Z(n42809) );
  NANDN U43602 ( .A(n42807), .B(n42806), .Z(n42808) );
  AND U43603 ( .A(n42809), .B(n42808), .Z(n42843) );
  XOR U43604 ( .A(n42843), .B(n42842), .Z(n42845) );
  XOR U43605 ( .A(n42844), .B(n42845), .Z(n42873) );
  NANDN U43606 ( .A(n42814), .B(n42813), .Z(n42818) );
  NANDN U43607 ( .A(n42816), .B(n42815), .Z(n42817) );
  NAND U43608 ( .A(n42818), .B(n42817), .Z(n42872) );
  XNOR U43609 ( .A(n42873), .B(n42872), .Z(n42874) );
  XNOR U43610 ( .A(n42875), .B(n42874), .Z(n42830) );
  XNOR U43611 ( .A(n42829), .B(n42830), .Z(n42832) );
  XOR U43612 ( .A(n42831), .B(n42832), .Z(n42838) );
  NANDN U43613 ( .A(n42823), .B(n42822), .Z(n42827) );
  NAND U43614 ( .A(n42825), .B(n42824), .Z(n42826) );
  AND U43615 ( .A(n42827), .B(n42826), .Z(n42836) );
  IV U43616 ( .A(n42836), .Z(n42835) );
  XOR U43617 ( .A(n42837), .B(n42835), .Z(n42828) );
  XNOR U43618 ( .A(n42838), .B(n42828), .Z(N940) );
  NAND U43619 ( .A(n42830), .B(n42829), .Z(n42834) );
  NANDN U43620 ( .A(n42832), .B(n42831), .Z(n42833) );
  NAND U43621 ( .A(n42834), .B(n42833), .Z(n42896) );
  OR U43622 ( .A(n42837), .B(n42835), .Z(n42841) );
  ANDN U43623 ( .B(n42837), .A(n42836), .Z(n42839) );
  OR U43624 ( .A(n42839), .B(n42838), .Z(n42840) );
  AND U43625 ( .A(n42841), .B(n42840), .Z(n42897) );
  NANDN U43626 ( .A(n42843), .B(n42842), .Z(n42847) );
  OR U43627 ( .A(n42845), .B(n42844), .Z(n42846) );
  NAND U43628 ( .A(n42847), .B(n42846), .Z(n42962) );
  AND U43629 ( .A(x[485]), .B(y[8137]), .Z(n43356) );
  NAND U43630 ( .A(n43541), .B(n43356), .Z(n42851) );
  NAND U43631 ( .A(n42849), .B(n42848), .Z(n42850) );
  NAND U43632 ( .A(n42851), .B(n42850), .Z(n42910) );
  AND U43633 ( .A(x[486]), .B(y[8138]), .Z(n43143) );
  XOR U43634 ( .A(n42910), .B(n42909), .Z(n42912) );
  AND U43635 ( .A(x[489]), .B(y[8131]), .Z(n43536) );
  AND U43636 ( .A(y[8130]), .B(x[490]), .Z(n43591) );
  NAND U43637 ( .A(y[8136]), .B(x[484]), .Z(n42855) );
  XNOR U43638 ( .A(n43591), .B(n42855), .Z(n42953) );
  XOR U43639 ( .A(n43536), .B(n42953), .Z(n42932) );
  NAND U43640 ( .A(x[487]), .B(y[8133]), .Z(n42930) );
  XOR U43641 ( .A(n42931), .B(n42930), .Z(n42933) );
  AND U43642 ( .A(y[8128]), .B(x[492]), .Z(n42857) );
  NAND U43643 ( .A(y[8140]), .B(x[480]), .Z(n42856) );
  XNOR U43644 ( .A(n42857), .B(n42856), .Z(n42947) );
  AND U43645 ( .A(x[491]), .B(y[8129]), .Z(n42927) );
  XOR U43646 ( .A(o[460]), .B(n42927), .Z(n42946) );
  XOR U43647 ( .A(n42947), .B(n42946), .Z(n42916) );
  AND U43648 ( .A(y[8138]), .B(x[482]), .Z(n42859) );
  NAND U43649 ( .A(y[8132]), .B(x[488]), .Z(n42858) );
  XNOR U43650 ( .A(n42859), .B(n42858), .Z(n42921) );
  XOR U43651 ( .A(n42916), .B(n42915), .Z(n42918) );
  XOR U43652 ( .A(n42917), .B(n42918), .Z(n42911) );
  XOR U43653 ( .A(n42912), .B(n42911), .Z(n42961) );
  AND U43654 ( .A(x[491]), .B(y[8139]), .Z(n43939) );
  NAND U43655 ( .A(n43939), .B(n43131), .Z(n42863) );
  NAND U43656 ( .A(n42861), .B(n42860), .Z(n42862) );
  NAND U43657 ( .A(n42863), .B(n42862), .Z(n42939) );
  AND U43658 ( .A(x[487]), .B(y[8130]), .Z(n43069) );
  AND U43659 ( .A(x[489]), .B(y[8132]), .Z(n42864) );
  NAND U43660 ( .A(n43069), .B(n42864), .Z(n42868) );
  NAND U43661 ( .A(n42866), .B(n42865), .Z(n42867) );
  NAND U43662 ( .A(n42868), .B(n42867), .Z(n42937) );
  NAND U43663 ( .A(y[8139]), .B(x[481]), .Z(n42869) );
  XNOR U43664 ( .A(n42870), .B(n42869), .Z(n42943) );
  AND U43665 ( .A(o[459]), .B(n42871), .Z(n42942) );
  XOR U43666 ( .A(n42943), .B(n42942), .Z(n42936) );
  XOR U43667 ( .A(n42937), .B(n42936), .Z(n42938) );
  XOR U43668 ( .A(n42939), .B(n42938), .Z(n42960) );
  XOR U43669 ( .A(n42961), .B(n42960), .Z(n42963) );
  XNOR U43670 ( .A(n42962), .B(n42963), .Z(n42899) );
  NANDN U43671 ( .A(n42873), .B(n42872), .Z(n42877) );
  NAND U43672 ( .A(n42875), .B(n42874), .Z(n42876) );
  NAND U43673 ( .A(n42877), .B(n42876), .Z(n42900) );
  XOR U43674 ( .A(n42899), .B(n42900), .Z(n42902) );
  IV U43675 ( .A(n43816), .Z(n43550) );
  NANDN U43676 ( .A(n43550), .B(n42878), .Z(n42882) );
  NAND U43677 ( .A(n42880), .B(n42879), .Z(n42881) );
  NAND U43678 ( .A(n42882), .B(n42881), .Z(n42903) );
  NAND U43679 ( .A(n42884), .B(n42883), .Z(n42888) );
  NAND U43680 ( .A(n42886), .B(n42885), .Z(n42887) );
  AND U43681 ( .A(n42888), .B(n42887), .Z(n42904) );
  XOR U43682 ( .A(n42903), .B(n42904), .Z(n42906) );
  NANDN U43683 ( .A(n42890), .B(n42889), .Z(n42894) );
  NANDN U43684 ( .A(n42892), .B(n42891), .Z(n42893) );
  AND U43685 ( .A(n42894), .B(n42893), .Z(n42905) );
  XOR U43686 ( .A(n42906), .B(n42905), .Z(n42901) );
  XOR U43687 ( .A(n42902), .B(n42901), .Z(n42898) );
  XNOR U43688 ( .A(n42897), .B(n42898), .Z(n42895) );
  XNOR U43689 ( .A(n42896), .B(n42895), .Z(N941) );
  NAND U43690 ( .A(n42904), .B(n42903), .Z(n42908) );
  NAND U43691 ( .A(n42906), .B(n42905), .Z(n42907) );
  NAND U43692 ( .A(n42908), .B(n42907), .Z(n43040) );
  NAND U43693 ( .A(n42910), .B(n42909), .Z(n42914) );
  NAND U43694 ( .A(n42912), .B(n42911), .Z(n42913) );
  NAND U43695 ( .A(n42914), .B(n42913), .Z(n42968) );
  NAND U43696 ( .A(n42916), .B(n42915), .Z(n42920) );
  NAND U43697 ( .A(n42918), .B(n42917), .Z(n42919) );
  NAND U43698 ( .A(n42920), .B(n42919), .Z(n42975) );
  AND U43699 ( .A(y[8138]), .B(x[488]), .Z(n44190) );
  AND U43700 ( .A(x[482]), .B(y[8132]), .Z(n43077) );
  NAND U43701 ( .A(n44190), .B(n43077), .Z(n42924) );
  NANDN U43702 ( .A(n42922), .B(n42921), .Z(n42923) );
  NAND U43703 ( .A(n42924), .B(n42923), .Z(n43007) );
  NAND U43704 ( .A(y[8140]), .B(x[481]), .Z(n42925) );
  XNOR U43705 ( .A(n42926), .B(n42925), .Z(n42997) );
  AND U43706 ( .A(o[460]), .B(n42927), .Z(n42996) );
  XOR U43707 ( .A(n42997), .B(n42996), .Z(n43005) );
  AND U43708 ( .A(x[486]), .B(y[8135]), .Z(n43979) );
  AND U43709 ( .A(y[8139]), .B(x[482]), .Z(n42929) );
  NAND U43710 ( .A(y[8132]), .B(x[489]), .Z(n42928) );
  XNOR U43711 ( .A(n42929), .B(n42928), .Z(n43011) );
  XOR U43712 ( .A(n43979), .B(n43011), .Z(n43004) );
  XOR U43713 ( .A(n43005), .B(n43004), .Z(n43006) );
  XOR U43714 ( .A(n43007), .B(n43006), .Z(n42974) );
  NAND U43715 ( .A(n42931), .B(n42930), .Z(n42935) );
  ANDN U43716 ( .B(n42933), .A(n42932), .Z(n42934) );
  ANDN U43717 ( .B(n42935), .A(n42934), .Z(n42973) );
  XOR U43718 ( .A(n42974), .B(n42973), .Z(n42976) );
  XOR U43719 ( .A(n42975), .B(n42976), .Z(n42967) );
  XOR U43720 ( .A(n42968), .B(n42967), .Z(n42970) );
  NAND U43721 ( .A(n42937), .B(n42936), .Z(n42941) );
  NAND U43722 ( .A(n42939), .B(n42938), .Z(n42940) );
  NAND U43723 ( .A(n42941), .B(n42940), .Z(n42982) );
  AND U43724 ( .A(x[486]), .B(y[8139]), .Z(n43289) );
  IV U43725 ( .A(n43289), .Z(n43358) );
  AND U43726 ( .A(x[481]), .B(y[8134]), .Z(n42995) );
  NANDN U43727 ( .A(n43358), .B(n42995), .Z(n42945) );
  NAND U43728 ( .A(n42943), .B(n42942), .Z(n42944) );
  NAND U43729 ( .A(n42945), .B(n42944), .Z(n42988) );
  AND U43730 ( .A(x[492]), .B(y[8140]), .Z(n44196) );
  NAND U43731 ( .A(n44196), .B(n43131), .Z(n42949) );
  NAND U43732 ( .A(n42947), .B(n42946), .Z(n42948) );
  NAND U43733 ( .A(n42949), .B(n42948), .Z(n42986) );
  AND U43734 ( .A(x[490]), .B(y[8131]), .Z(n43828) );
  AND U43735 ( .A(y[8130]), .B(x[491]), .Z(n43789) );
  NAND U43736 ( .A(y[8133]), .B(x[488]), .Z(n42950) );
  XNOR U43737 ( .A(n43789), .B(n42950), .Z(n42992) );
  XOR U43738 ( .A(n43828), .B(n42992), .Z(n42985) );
  XOR U43739 ( .A(n42986), .B(n42985), .Z(n42987) );
  XOR U43740 ( .A(n42988), .B(n42987), .Z(n42980) );
  AND U43741 ( .A(x[490]), .B(y[8136]), .Z(n42952) );
  AND U43742 ( .A(x[484]), .B(y[8130]), .Z(n42951) );
  NAND U43743 ( .A(n42952), .B(n42951), .Z(n42955) );
  NAND U43744 ( .A(n42953), .B(n43536), .Z(n42954) );
  NAND U43745 ( .A(n42955), .B(n42954), .Z(n43032) );
  AND U43746 ( .A(y[8128]), .B(x[493]), .Z(n42957) );
  NAND U43747 ( .A(y[8141]), .B(x[480]), .Z(n42956) );
  XNOR U43748 ( .A(n42957), .B(n42956), .Z(n43023) );
  NAND U43749 ( .A(x[492]), .B(y[8129]), .Z(n43016) );
  XNOR U43750 ( .A(o[461]), .B(n43016), .Z(n43024) );
  XOR U43751 ( .A(n43023), .B(n43024), .Z(n43030) );
  AND U43752 ( .A(y[8136]), .B(x[485]), .Z(n42959) );
  NAND U43753 ( .A(y[8138]), .B(x[483]), .Z(n42958) );
  XNOR U43754 ( .A(n42959), .B(n42958), .Z(n43019) );
  AND U43755 ( .A(x[484]), .B(y[8137]), .Z(n43020) );
  XOR U43756 ( .A(n43019), .B(n43020), .Z(n43029) );
  XOR U43757 ( .A(n43030), .B(n43029), .Z(n43031) );
  XOR U43758 ( .A(n43032), .B(n43031), .Z(n42979) );
  XOR U43759 ( .A(n42980), .B(n42979), .Z(n42981) );
  XOR U43760 ( .A(n42982), .B(n42981), .Z(n42969) );
  XOR U43761 ( .A(n42970), .B(n42969), .Z(n43039) );
  NAND U43762 ( .A(n42961), .B(n42960), .Z(n42965) );
  NAND U43763 ( .A(n42963), .B(n42962), .Z(n42964) );
  AND U43764 ( .A(n42965), .B(n42964), .Z(n43038) );
  XOR U43765 ( .A(n43040), .B(n43041), .Z(n43037) );
  XNOR U43766 ( .A(n43036), .B(n43037), .Z(n42966) );
  XOR U43767 ( .A(n43035), .B(n42966), .Z(N942) );
  NAND U43768 ( .A(n42968), .B(n42967), .Z(n42972) );
  NAND U43769 ( .A(n42970), .B(n42969), .Z(n42971) );
  NAND U43770 ( .A(n42972), .B(n42971), .Z(n43120) );
  NAND U43771 ( .A(n42974), .B(n42973), .Z(n42978) );
  NAND U43772 ( .A(n42976), .B(n42975), .Z(n42977) );
  NAND U43773 ( .A(n42978), .B(n42977), .Z(n43119) );
  XOR U43774 ( .A(n43120), .B(n43119), .Z(n43122) );
  NAND U43775 ( .A(n42980), .B(n42979), .Z(n42984) );
  NAND U43776 ( .A(n42982), .B(n42981), .Z(n42983) );
  NAND U43777 ( .A(n42984), .B(n42983), .Z(n43048) );
  NAND U43778 ( .A(n42986), .B(n42985), .Z(n42990) );
  NAND U43779 ( .A(n42988), .B(n42987), .Z(n42989) );
  AND U43780 ( .A(n42990), .B(n42989), .Z(n43054) );
  AND U43781 ( .A(x[491]), .B(y[8133]), .Z(n43154) );
  NAND U43782 ( .A(n43154), .B(n42991), .Z(n42994) );
  NAND U43783 ( .A(n42992), .B(n43828), .Z(n42993) );
  NAND U43784 ( .A(n42994), .B(n42993), .Z(n43105) );
  NAND U43785 ( .A(x[487]), .B(y[8140]), .Z(n43552) );
  NANDN U43786 ( .A(n43552), .B(n42995), .Z(n42999) );
  NAND U43787 ( .A(n42997), .B(n42996), .Z(n42998) );
  NAND U43788 ( .A(n42999), .B(n42998), .Z(n43104) );
  XOR U43789 ( .A(n43105), .B(n43104), .Z(n43107) );
  AND U43790 ( .A(x[484]), .B(y[8138]), .Z(n43473) );
  AND U43791 ( .A(y[8139]), .B(x[483]), .Z(n43001) );
  NAND U43792 ( .A(y[8134]), .B(x[488]), .Z(n43000) );
  XNOR U43793 ( .A(n43001), .B(n43000), .Z(n43090) );
  XOR U43794 ( .A(n43356), .B(n43090), .Z(n43099) );
  XOR U43795 ( .A(n43473), .B(n43099), .Z(n43101) );
  AND U43796 ( .A(x[489]), .B(y[8133]), .Z(n43658) );
  AND U43797 ( .A(y[8140]), .B(x[482]), .Z(n43003) );
  NAND U43798 ( .A(y[8132]), .B(x[490]), .Z(n43002) );
  XNOR U43799 ( .A(n43003), .B(n43002), .Z(n43078) );
  XOR U43800 ( .A(n43658), .B(n43078), .Z(n43100) );
  XOR U43801 ( .A(n43101), .B(n43100), .Z(n43106) );
  XNOR U43802 ( .A(n43107), .B(n43106), .Z(n43052) );
  NAND U43803 ( .A(n43005), .B(n43004), .Z(n43009) );
  NAND U43804 ( .A(n43007), .B(n43006), .Z(n43008) );
  AND U43805 ( .A(n43009), .B(n43008), .Z(n43051) );
  XOR U43806 ( .A(n43052), .B(n43051), .Z(n43053) );
  XNOR U43807 ( .A(n43054), .B(n43053), .Z(n43046) );
  AND U43808 ( .A(x[489]), .B(y[8139]), .Z(n43010) );
  NAND U43809 ( .A(n43010), .B(n43077), .Z(n43013) );
  NAND U43810 ( .A(n43011), .B(n43979), .Z(n43012) );
  NAND U43811 ( .A(n43013), .B(n43012), .Z(n43065) );
  AND U43812 ( .A(y[8128]), .B(x[494]), .Z(n43015) );
  NAND U43813 ( .A(y[8142]), .B(x[480]), .Z(n43014) );
  XNOR U43814 ( .A(n43015), .B(n43014), .Z(n43087) );
  ANDN U43815 ( .B(o[461]), .A(n43016), .Z(n43086) );
  XOR U43816 ( .A(n43087), .B(n43086), .Z(n43064) );
  NAND U43817 ( .A(y[8130]), .B(x[492]), .Z(n43017) );
  XNOR U43818 ( .A(n43018), .B(n43017), .Z(n43071) );
  AND U43819 ( .A(x[493]), .B(y[8129]), .Z(n43076) );
  XOR U43820 ( .A(n43076), .B(o[462]), .Z(n43070) );
  XOR U43821 ( .A(n43071), .B(n43070), .Z(n43063) );
  XOR U43822 ( .A(n43064), .B(n43063), .Z(n43066) );
  XNOR U43823 ( .A(n43065), .B(n43066), .Z(n43111) );
  NAND U43824 ( .A(x[485]), .B(y[8138]), .Z(n43145) );
  NANDN U43825 ( .A(n43145), .B(n43550), .Z(n43022) );
  NAND U43826 ( .A(n43020), .B(n43019), .Z(n43021) );
  NAND U43827 ( .A(n43022), .B(n43021), .Z(n43059) );
  AND U43828 ( .A(x[493]), .B(y[8141]), .Z(n44573) );
  NAND U43829 ( .A(n44573), .B(n43131), .Z(n43026) );
  NAND U43830 ( .A(n43024), .B(n43023), .Z(n43025) );
  NAND U43831 ( .A(n43026), .B(n43025), .Z(n43057) );
  NAND U43832 ( .A(y[8131]), .B(x[491]), .Z(n43027) );
  XNOR U43833 ( .A(n43028), .B(n43027), .Z(n43083) );
  AND U43834 ( .A(x[481]), .B(y[8141]), .Z(n43082) );
  XOR U43835 ( .A(n43083), .B(n43082), .Z(n43058) );
  XNOR U43836 ( .A(n43057), .B(n43058), .Z(n43060) );
  XOR U43837 ( .A(n43059), .B(n43060), .Z(n43110) );
  XOR U43838 ( .A(n43111), .B(n43110), .Z(n43113) );
  NAND U43839 ( .A(n43030), .B(n43029), .Z(n43034) );
  NAND U43840 ( .A(n43032), .B(n43031), .Z(n43033) );
  AND U43841 ( .A(n43034), .B(n43033), .Z(n43112) );
  XNOR U43842 ( .A(n43113), .B(n43112), .Z(n43045) );
  XOR U43843 ( .A(n43046), .B(n43045), .Z(n43047) );
  XOR U43844 ( .A(n43048), .B(n43047), .Z(n43121) );
  XNOR U43845 ( .A(n43122), .B(n43121), .Z(n43118) );
  NANDN U43846 ( .A(n43039), .B(n43038), .Z(n43043) );
  NAND U43847 ( .A(n43041), .B(n43040), .Z(n43042) );
  AND U43848 ( .A(n43043), .B(n43042), .Z(n43117) );
  XOR U43849 ( .A(n43116), .B(n43117), .Z(n43044) );
  XNOR U43850 ( .A(n43118), .B(n43044), .Z(N943) );
  NAND U43851 ( .A(n43046), .B(n43045), .Z(n43050) );
  NAND U43852 ( .A(n43048), .B(n43047), .Z(n43049) );
  NAND U43853 ( .A(n43050), .B(n43049), .Z(n43204) );
  NAND U43854 ( .A(n43052), .B(n43051), .Z(n43056) );
  NAND U43855 ( .A(n43054), .B(n43053), .Z(n43055) );
  NAND U43856 ( .A(n43056), .B(n43055), .Z(n43179) );
  NAND U43857 ( .A(n43058), .B(n43057), .Z(n43062) );
  NANDN U43858 ( .A(n43060), .B(n43059), .Z(n43061) );
  NAND U43859 ( .A(n43062), .B(n43061), .Z(n43185) );
  NAND U43860 ( .A(n43064), .B(n43063), .Z(n43068) );
  NAND U43861 ( .A(n43066), .B(n43065), .Z(n43067) );
  NAND U43862 ( .A(n43068), .B(n43067), .Z(n43183) );
  NAND U43863 ( .A(x[492]), .B(y[8135]), .Z(n43543) );
  AND U43864 ( .A(y[8132]), .B(x[491]), .Z(n43073) );
  NAND U43865 ( .A(y[8130]), .B(x[493]), .Z(n43072) );
  XNOR U43866 ( .A(n43073), .B(n43072), .Z(n43163) );
  NAND U43867 ( .A(x[492]), .B(y[8131]), .Z(n43164) );
  XOR U43868 ( .A(n43163), .B(n43164), .Z(n43159) );
  AND U43869 ( .A(y[8128]), .B(x[495]), .Z(n43075) );
  NAND U43870 ( .A(y[8143]), .B(x[480]), .Z(n43074) );
  XNOR U43871 ( .A(n43075), .B(n43074), .Z(n43132) );
  NAND U43872 ( .A(n43076), .B(o[462]), .Z(n43133) );
  XOR U43873 ( .A(n43132), .B(n43133), .Z(n43160) );
  XNOR U43874 ( .A(n43159), .B(n43160), .Z(n43162) );
  XOR U43875 ( .A(n43161), .B(n43162), .Z(n43191) );
  AND U43876 ( .A(x[490]), .B(y[8140]), .Z(n43980) );
  NAND U43877 ( .A(n43077), .B(n43980), .Z(n43080) );
  NAND U43878 ( .A(n43658), .B(n43078), .Z(n43079) );
  NAND U43879 ( .A(n43080), .B(n43079), .Z(n43190) );
  AND U43880 ( .A(x[491]), .B(y[8136]), .Z(n43471) );
  NAND U43881 ( .A(n43471), .B(n43081), .Z(n43085) );
  NAND U43882 ( .A(n43083), .B(n43082), .Z(n43084) );
  NAND U43883 ( .A(n43085), .B(n43084), .Z(n43189) );
  XOR U43884 ( .A(n43190), .B(n43189), .Z(n43192) );
  XOR U43885 ( .A(n43191), .B(n43192), .Z(n43184) );
  XOR U43886 ( .A(n43183), .B(n43184), .Z(n43186) );
  XOR U43887 ( .A(n43185), .B(n43186), .Z(n43178) );
  AND U43888 ( .A(x[494]), .B(y[8142]), .Z(n44849) );
  AND U43889 ( .A(x[488]), .B(y[8139]), .Z(n43088) );
  NANDN U43890 ( .A(n43089), .B(n43088), .Z(n43092) );
  NAND U43891 ( .A(n43356), .B(n43090), .Z(n43091) );
  NAND U43892 ( .A(n43092), .B(n43091), .Z(n43156) );
  XOR U43893 ( .A(n43155), .B(n43156), .Z(n43157) );
  AND U43894 ( .A(y[8133]), .B(x[490]), .Z(n43094) );
  NAND U43895 ( .A(y[8139]), .B(x[484]), .Z(n43093) );
  XNOR U43896 ( .A(n43094), .B(n43093), .Z(n43138) );
  NAND U43897 ( .A(x[487]), .B(y[8136]), .Z(n43139) );
  XOR U43898 ( .A(n43138), .B(n43139), .Z(n43146) );
  NAND U43899 ( .A(x[486]), .B(y[8137]), .Z(n43144) );
  XOR U43900 ( .A(n43144), .B(n43145), .Z(n43147) );
  XOR U43901 ( .A(n43146), .B(n43147), .Z(n43174) );
  AND U43902 ( .A(y[8141]), .B(x[482]), .Z(n43096) );
  NAND U43903 ( .A(y[8134]), .B(x[489]), .Z(n43095) );
  XNOR U43904 ( .A(n43096), .B(n43095), .Z(n43149) );
  AND U43905 ( .A(x[483]), .B(y[8140]), .Z(n43148) );
  XOR U43906 ( .A(n43149), .B(n43148), .Z(n43172) );
  AND U43907 ( .A(y[8142]), .B(x[481]), .Z(n43098) );
  NAND U43908 ( .A(y[8135]), .B(x[488]), .Z(n43097) );
  XNOR U43909 ( .A(n43098), .B(n43097), .Z(n43127) );
  NAND U43910 ( .A(x[494]), .B(y[8129]), .Z(n43152) );
  XOR U43911 ( .A(o[463]), .B(n43152), .Z(n43128) );
  XNOR U43912 ( .A(n43127), .B(n43128), .Z(n43171) );
  XOR U43913 ( .A(n43172), .B(n43171), .Z(n43173) );
  XOR U43914 ( .A(n43174), .B(n43173), .Z(n43158) );
  XOR U43915 ( .A(n43157), .B(n43158), .Z(n43195) );
  NAND U43916 ( .A(n43473), .B(n43099), .Z(n43103) );
  NAND U43917 ( .A(n43101), .B(n43100), .Z(n43102) );
  AND U43918 ( .A(n43103), .B(n43102), .Z(n43196) );
  XOR U43919 ( .A(n43195), .B(n43196), .Z(n43198) );
  NAND U43920 ( .A(n43105), .B(n43104), .Z(n43109) );
  NAND U43921 ( .A(n43107), .B(n43106), .Z(n43108) );
  AND U43922 ( .A(n43109), .B(n43108), .Z(n43197) );
  XOR U43923 ( .A(n43198), .B(n43197), .Z(n43177) );
  XOR U43924 ( .A(n43179), .B(n43180), .Z(n43201) );
  NAND U43925 ( .A(n43111), .B(n43110), .Z(n43115) );
  NAND U43926 ( .A(n43113), .B(n43112), .Z(n43114) );
  AND U43927 ( .A(n43115), .B(n43114), .Z(n43202) );
  XOR U43928 ( .A(n43201), .B(n43202), .Z(n43203) );
  XOR U43929 ( .A(n43204), .B(n43203), .Z(n43210) );
  NAND U43930 ( .A(n43120), .B(n43119), .Z(n43124) );
  NAND U43931 ( .A(n43122), .B(n43121), .Z(n43123) );
  AND U43932 ( .A(n43124), .B(n43123), .Z(n43209) );
  IV U43933 ( .A(n43209), .Z(n43207) );
  XOR U43934 ( .A(n43208), .B(n43207), .Z(n43125) );
  XNOR U43935 ( .A(n43210), .B(n43125), .Z(N944) );
  AND U43936 ( .A(x[488]), .B(y[8142]), .Z(n43472) );
  NAND U43937 ( .A(n43472), .B(n43126), .Z(n43130) );
  NANDN U43938 ( .A(n43128), .B(n43127), .Z(n43129) );
  NAND U43939 ( .A(n43130), .B(n43129), .Z(n43268) );
  AND U43940 ( .A(x[495]), .B(y[8143]), .Z(n45162) );
  NAND U43941 ( .A(n45162), .B(n43131), .Z(n43135) );
  NANDN U43942 ( .A(n43133), .B(n43132), .Z(n43134) );
  NAND U43943 ( .A(n43135), .B(n43134), .Z(n43267) );
  XOR U43944 ( .A(n43268), .B(n43267), .Z(n43270) );
  AND U43945 ( .A(x[490]), .B(y[8139]), .Z(n43137) );
  NAND U43946 ( .A(n43137), .B(n43136), .Z(n43141) );
  NANDN U43947 ( .A(n43139), .B(n43138), .Z(n43140) );
  AND U43948 ( .A(n43141), .B(n43140), .Z(n43228) );
  AND U43949 ( .A(x[480]), .B(y[8144]), .Z(n43249) );
  AND U43950 ( .A(x[496]), .B(y[8128]), .Z(n43250) );
  XOR U43951 ( .A(n43249), .B(n43250), .Z(n43252) );
  AND U43952 ( .A(x[495]), .B(y[8129]), .Z(n43237) );
  XOR U43953 ( .A(o[464]), .B(n43237), .Z(n43251) );
  XOR U43954 ( .A(n43252), .B(n43251), .Z(n43225) );
  NAND U43955 ( .A(y[8137]), .B(x[487]), .Z(n43142) );
  XNOR U43956 ( .A(n43143), .B(n43142), .Z(n43242) );
  AND U43957 ( .A(x[490]), .B(y[8134]), .Z(n43241) );
  XNOR U43958 ( .A(n43242), .B(n43241), .Z(n43226) );
  XNOR U43959 ( .A(n43225), .B(n43226), .Z(n43227) );
  XNOR U43960 ( .A(n43228), .B(n43227), .Z(n43269) );
  XOR U43961 ( .A(n43270), .B(n43269), .Z(n43224) );
  IV U43962 ( .A(n43144), .Z(n43240) );
  AND U43963 ( .A(x[489]), .B(y[8141]), .Z(n43961) );
  AND U43964 ( .A(y[8143]), .B(x[481]), .Z(n43151) );
  NAND U43965 ( .A(y[8136]), .B(x[488]), .Z(n43150) );
  XNOR U43966 ( .A(n43151), .B(n43150), .Z(n43246) );
  ANDN U43967 ( .B(o[463]), .A(n43152), .Z(n43245) );
  XOR U43968 ( .A(n43246), .B(n43245), .Z(n43258) );
  NAND U43969 ( .A(y[8130]), .B(x[494]), .Z(n43153) );
  XNOR U43970 ( .A(n43154), .B(n43153), .Z(n43279) );
  AND U43971 ( .A(x[484]), .B(y[8140]), .Z(n43280) );
  XOR U43972 ( .A(n43279), .B(n43280), .Z(n43257) );
  XNOR U43973 ( .A(n43258), .B(n43257), .Z(n43260) );
  XOR U43974 ( .A(n43259), .B(n43260), .Z(n43222) );
  XOR U43975 ( .A(n43221), .B(n43222), .Z(n43223) );
  XNOR U43976 ( .A(n43224), .B(n43223), .Z(n43264) );
  XOR U43977 ( .A(n43264), .B(n43263), .Z(n43265) );
  AND U43978 ( .A(x[493]), .B(y[8132]), .Z(n43291) );
  NAND U43979 ( .A(n43291), .B(n43789), .Z(n43166) );
  NANDN U43980 ( .A(n43164), .B(n43163), .Z(n43165) );
  AND U43981 ( .A(n43166), .B(n43165), .Z(n43276) );
  AND U43982 ( .A(y[8142]), .B(x[482]), .Z(n43168) );
  NAND U43983 ( .A(y[8135]), .B(x[489]), .Z(n43167) );
  XNOR U43984 ( .A(n43168), .B(n43167), .Z(n43284) );
  NAND U43985 ( .A(x[483]), .B(y[8141]), .Z(n43285) );
  XNOR U43986 ( .A(n43284), .B(n43285), .Z(n43273) );
  AND U43987 ( .A(x[492]), .B(y[8132]), .Z(n43950) );
  AND U43988 ( .A(y[8139]), .B(x[485]), .Z(n43170) );
  NAND U43989 ( .A(y[8131]), .B(x[493]), .Z(n43169) );
  XOR U43990 ( .A(n43170), .B(n43169), .Z(n43232) );
  XOR U43991 ( .A(n43950), .B(n43232), .Z(n43274) );
  XNOR U43992 ( .A(n43273), .B(n43274), .Z(n43275) );
  XOR U43993 ( .A(n43276), .B(n43275), .Z(n43293) );
  NAND U43994 ( .A(n43172), .B(n43171), .Z(n43176) );
  NANDN U43995 ( .A(n43174), .B(n43173), .Z(n43175) );
  AND U43996 ( .A(n43176), .B(n43175), .Z(n43292) );
  XNOR U43997 ( .A(n43293), .B(n43292), .Z(n43295) );
  XOR U43998 ( .A(n43294), .B(n43295), .Z(n43266) );
  XOR U43999 ( .A(n43265), .B(n43266), .Z(n43296) );
  NANDN U44000 ( .A(n43178), .B(n43177), .Z(n43182) );
  NANDN U44001 ( .A(n43180), .B(n43179), .Z(n43181) );
  AND U44002 ( .A(n43182), .B(n43181), .Z(n43297) );
  XOR U44003 ( .A(n43296), .B(n43297), .Z(n43299) );
  NAND U44004 ( .A(n43184), .B(n43183), .Z(n43188) );
  NAND U44005 ( .A(n43186), .B(n43185), .Z(n43187) );
  NAND U44006 ( .A(n43188), .B(n43187), .Z(n43217) );
  NAND U44007 ( .A(n43190), .B(n43189), .Z(n43194) );
  NAND U44008 ( .A(n43192), .B(n43191), .Z(n43193) );
  NAND U44009 ( .A(n43194), .B(n43193), .Z(n43215) );
  NAND U44010 ( .A(n43196), .B(n43195), .Z(n43200) );
  NAND U44011 ( .A(n43198), .B(n43197), .Z(n43199) );
  AND U44012 ( .A(n43200), .B(n43199), .Z(n43216) );
  XOR U44013 ( .A(n43215), .B(n43216), .Z(n43218) );
  XOR U44014 ( .A(n43217), .B(n43218), .Z(n43298) );
  XNOR U44015 ( .A(n43299), .B(n43298), .Z(n43304) );
  NAND U44016 ( .A(n43202), .B(n43201), .Z(n43206) );
  NAND U44017 ( .A(n43204), .B(n43203), .Z(n43205) );
  NAND U44018 ( .A(n43206), .B(n43205), .Z(n43303) );
  NANDN U44019 ( .A(n43207), .B(n43208), .Z(n43213) );
  NOR U44020 ( .A(n43209), .B(n43208), .Z(n43211) );
  OR U44021 ( .A(n43211), .B(n43210), .Z(n43212) );
  AND U44022 ( .A(n43213), .B(n43212), .Z(n43302) );
  XOR U44023 ( .A(n43303), .B(n43302), .Z(n43214) );
  XNOR U44024 ( .A(n43304), .B(n43214), .Z(N945) );
  NAND U44025 ( .A(n43216), .B(n43215), .Z(n43220) );
  NAND U44026 ( .A(n43218), .B(n43217), .Z(n43219) );
  NAND U44027 ( .A(n43220), .B(n43219), .Z(n43401) );
  NANDN U44028 ( .A(n43226), .B(n43225), .Z(n43230) );
  NANDN U44029 ( .A(n43228), .B(n43227), .Z(n43229) );
  NAND U44030 ( .A(n43230), .B(n43229), .Z(n43393) );
  AND U44031 ( .A(x[493]), .B(y[8139]), .Z(n44204) );
  NAND U44032 ( .A(n44204), .B(n43231), .Z(n43234) );
  NANDN U44033 ( .A(n43232), .B(n43950), .Z(n43233) );
  NAND U44034 ( .A(n43234), .B(n43233), .Z(n43341) );
  AND U44035 ( .A(y[8144]), .B(x[481]), .Z(n43236) );
  NAND U44036 ( .A(y[8136]), .B(x[489]), .Z(n43235) );
  XNOR U44037 ( .A(n43236), .B(n43235), .Z(n43362) );
  AND U44038 ( .A(o[464]), .B(n43237), .Z(n43361) );
  XOR U44039 ( .A(n43362), .B(n43361), .Z(n43339) );
  AND U44040 ( .A(y[8130]), .B(x[495]), .Z(n43239) );
  NAND U44041 ( .A(y[8133]), .B(x[492]), .Z(n43238) );
  XNOR U44042 ( .A(n43239), .B(n43238), .Z(n43315) );
  AND U44043 ( .A(x[494]), .B(y[8131]), .Z(n43314) );
  XOR U44044 ( .A(n43315), .B(n43314), .Z(n43338) );
  XOR U44045 ( .A(n43339), .B(n43338), .Z(n43340) );
  XOR U44046 ( .A(n43341), .B(n43340), .Z(n43391) );
  NAND U44047 ( .A(x[487]), .B(y[8138]), .Z(n43373) );
  NANDN U44048 ( .A(n43373), .B(n43240), .Z(n43244) );
  NAND U44049 ( .A(n43242), .B(n43241), .Z(n43243) );
  NAND U44050 ( .A(n43244), .B(n43243), .Z(n43351) );
  NAND U44051 ( .A(x[488]), .B(y[8143]), .Z(n44044) );
  AND U44052 ( .A(x[481]), .B(y[8136]), .Z(n43451) );
  NANDN U44053 ( .A(n44044), .B(n43451), .Z(n43248) );
  NAND U44054 ( .A(n43246), .B(n43245), .Z(n43247) );
  NAND U44055 ( .A(n43248), .B(n43247), .Z(n43350) );
  XOR U44056 ( .A(n43351), .B(n43350), .Z(n43353) );
  NAND U44057 ( .A(n43250), .B(n43249), .Z(n43254) );
  NAND U44058 ( .A(n43252), .B(n43251), .Z(n43253) );
  NAND U44059 ( .A(n43254), .B(n43253), .Z(n43347) );
  AND U44060 ( .A(x[480]), .B(y[8145]), .Z(n43329) );
  AND U44061 ( .A(x[497]), .B(y[8128]), .Z(n43328) );
  XOR U44062 ( .A(n43329), .B(n43328), .Z(n43331) );
  AND U44063 ( .A(x[496]), .B(y[8129]), .Z(n43325) );
  XOR U44064 ( .A(n43325), .B(o[465]), .Z(n43330) );
  XOR U44065 ( .A(n43331), .B(n43330), .Z(n43345) );
  AND U44066 ( .A(y[8143]), .B(x[482]), .Z(n43256) );
  NAND U44067 ( .A(y[8135]), .B(x[490]), .Z(n43255) );
  XNOR U44068 ( .A(n43256), .B(n43255), .Z(n43366) );
  NAND U44069 ( .A(x[483]), .B(y[8142]), .Z(n43367) );
  XOR U44070 ( .A(n43345), .B(n43344), .Z(n43346) );
  XOR U44071 ( .A(n43347), .B(n43346), .Z(n43352) );
  XOR U44072 ( .A(n43353), .B(n43352), .Z(n43390) );
  XOR U44073 ( .A(n43391), .B(n43390), .Z(n43392) );
  XOR U44074 ( .A(n43393), .B(n43392), .Z(n43311) );
  NAND U44075 ( .A(n43258), .B(n43257), .Z(n43262) );
  NANDN U44076 ( .A(n43260), .B(n43259), .Z(n43261) );
  AND U44077 ( .A(n43262), .B(n43261), .Z(n43310) );
  XNOR U44078 ( .A(n43311), .B(n43310), .Z(n43313) );
  XNOR U44079 ( .A(n43312), .B(n43313), .Z(n43400) );
  NAND U44080 ( .A(n43268), .B(n43267), .Z(n43272) );
  NAND U44081 ( .A(n43270), .B(n43269), .Z(n43271) );
  AND U44082 ( .A(n43272), .B(n43271), .Z(n43387) );
  NANDN U44083 ( .A(n43274), .B(n43273), .Z(n43278) );
  NANDN U44084 ( .A(n43276), .B(n43275), .Z(n43277) );
  AND U44085 ( .A(n43278), .B(n43277), .Z(n43385) );
  NAND U44086 ( .A(x[494]), .B(y[8133]), .Z(n43588) );
  NANDN U44087 ( .A(n43588), .B(n43789), .Z(n43282) );
  NAND U44088 ( .A(n43280), .B(n43279), .Z(n43281) );
  AND U44089 ( .A(n43282), .B(n43281), .Z(n43379) );
  AND U44090 ( .A(x[489]), .B(y[8142]), .Z(n44185) );
  NANDN U44091 ( .A(n43283), .B(n44185), .Z(n43287) );
  NANDN U44092 ( .A(n43285), .B(n43284), .Z(n43286) );
  NAND U44093 ( .A(n43287), .B(n43286), .Z(n43378) );
  XNOR U44094 ( .A(n43379), .B(n43378), .Z(n43380) );
  AND U44095 ( .A(x[485]), .B(y[8140]), .Z(n43433) );
  NAND U44096 ( .A(y[8137]), .B(x[488]), .Z(n43288) );
  XNOR U44097 ( .A(n43433), .B(n43288), .Z(n43357) );
  XOR U44098 ( .A(n43357), .B(n43289), .Z(n43372) );
  XNOR U44099 ( .A(n43372), .B(n43373), .Z(n43374) );
  NAND U44100 ( .A(y[8141]), .B(x[484]), .Z(n43290) );
  XNOR U44101 ( .A(n43291), .B(n43290), .Z(n43319) );
  NAND U44102 ( .A(x[491]), .B(y[8134]), .Z(n43320) );
  XOR U44103 ( .A(n43319), .B(n43320), .Z(n43375) );
  XOR U44104 ( .A(n43374), .B(n43375), .Z(n43381) );
  XNOR U44105 ( .A(n43380), .B(n43381), .Z(n43384) );
  XNOR U44106 ( .A(n43385), .B(n43384), .Z(n43386) );
  XOR U44107 ( .A(n43387), .B(n43386), .Z(n43306) );
  XNOR U44108 ( .A(n43306), .B(n43307), .Z(n43309) );
  XOR U44109 ( .A(n43308), .B(n43309), .Z(n43399) );
  XOR U44110 ( .A(n43400), .B(n43399), .Z(n43402) );
  XOR U44111 ( .A(n43401), .B(n43402), .Z(n43398) );
  NAND U44112 ( .A(n43297), .B(n43296), .Z(n43301) );
  NAND U44113 ( .A(n43299), .B(n43298), .Z(n43300) );
  AND U44114 ( .A(n43301), .B(n43300), .Z(n43397) );
  XNOR U44115 ( .A(n43397), .B(n43396), .Z(n43305) );
  XNOR U44116 ( .A(n43398), .B(n43305), .Z(N946) );
  AND U44117 ( .A(x[495]), .B(y[8133]), .Z(n43549) );
  AND U44118 ( .A(x[492]), .B(y[8130]), .Z(n43648) );
  NAND U44119 ( .A(n43549), .B(n43648), .Z(n43317) );
  NAND U44120 ( .A(n43315), .B(n43314), .Z(n43316) );
  NAND U44121 ( .A(n43317), .B(n43316), .Z(n43499) );
  NAND U44122 ( .A(n44573), .B(n43318), .Z(n43322) );
  NANDN U44123 ( .A(n43320), .B(n43319), .Z(n43321) );
  AND U44124 ( .A(n43322), .B(n43321), .Z(n43490) );
  AND U44125 ( .A(y[8145]), .B(x[481]), .Z(n43324) );
  NAND U44126 ( .A(y[8136]), .B(x[490]), .Z(n43323) );
  XNOR U44127 ( .A(n43324), .B(n43323), .Z(n43452) );
  AND U44128 ( .A(n43325), .B(o[465]), .Z(n43453) );
  XOR U44129 ( .A(n43452), .B(n43453), .Z(n43488) );
  AND U44130 ( .A(y[8131]), .B(x[495]), .Z(n43327) );
  NAND U44131 ( .A(y[8137]), .B(x[489]), .Z(n43326) );
  XNOR U44132 ( .A(n43327), .B(n43326), .Z(n43443) );
  AND U44133 ( .A(x[494]), .B(y[8132]), .Z(n43444) );
  XOR U44134 ( .A(n43443), .B(n43444), .Z(n43487) );
  XOR U44135 ( .A(n43488), .B(n43487), .Z(n43489) );
  XOR U44136 ( .A(n43499), .B(n43500), .Z(n43502) );
  NAND U44137 ( .A(n43329), .B(n43328), .Z(n43333) );
  NAND U44138 ( .A(n43331), .B(n43330), .Z(n43332) );
  NAND U44139 ( .A(n43333), .B(n43332), .Z(n43511) );
  AND U44140 ( .A(y[8130]), .B(x[496]), .Z(n43335) );
  NAND U44141 ( .A(y[8135]), .B(x[491]), .Z(n43334) );
  XNOR U44142 ( .A(n43335), .B(n43334), .Z(n43439) );
  NAND U44143 ( .A(x[482]), .B(y[8144]), .Z(n43440) );
  XOR U44144 ( .A(n43511), .B(n43512), .Z(n43514) );
  AND U44145 ( .A(y[8141]), .B(x[485]), .Z(n43570) );
  NAND U44146 ( .A(y[8140]), .B(x[486]), .Z(n43336) );
  XNOR U44147 ( .A(n43570), .B(n43336), .Z(n43436) );
  NAND U44148 ( .A(y[8142]), .B(x[484]), .Z(n43337) );
  XNOR U44149 ( .A(n44190), .B(n43337), .Z(n43474) );
  AND U44150 ( .A(x[487]), .B(y[8139]), .Z(n43475) );
  XOR U44151 ( .A(n43474), .B(n43475), .Z(n43435) );
  XOR U44152 ( .A(n43436), .B(n43435), .Z(n43513) );
  XOR U44153 ( .A(n43514), .B(n43513), .Z(n43501) );
  XNOR U44154 ( .A(n43502), .B(n43501), .Z(n43422) );
  NAND U44155 ( .A(n43339), .B(n43338), .Z(n43343) );
  NAND U44156 ( .A(n43341), .B(n43340), .Z(n43342) );
  AND U44157 ( .A(n43343), .B(n43342), .Z(n43494) );
  NAND U44158 ( .A(n43345), .B(n43344), .Z(n43349) );
  NAND U44159 ( .A(n43347), .B(n43346), .Z(n43348) );
  AND U44160 ( .A(n43349), .B(n43348), .Z(n43493) );
  XOR U44161 ( .A(n43494), .B(n43493), .Z(n43496) );
  NAND U44162 ( .A(n43351), .B(n43350), .Z(n43355) );
  NAND U44163 ( .A(n43353), .B(n43352), .Z(n43354) );
  AND U44164 ( .A(n43355), .B(n43354), .Z(n43495) );
  XOR U44165 ( .A(n43496), .B(n43495), .Z(n43421) );
  XOR U44166 ( .A(n43422), .B(n43421), .Z(n43424) );
  AND U44167 ( .A(x[488]), .B(y[8140]), .Z(n43688) );
  NAND U44168 ( .A(n43688), .B(n43356), .Z(n43360) );
  NANDN U44169 ( .A(n43358), .B(n43357), .Z(n43359) );
  NAND U44170 ( .A(n43360), .B(n43359), .Z(n43506) );
  NAND U44171 ( .A(x[489]), .B(y[8144]), .Z(n44332) );
  NANDN U44172 ( .A(n44332), .B(n43451), .Z(n43364) );
  NAND U44173 ( .A(n43362), .B(n43361), .Z(n43363) );
  NAND U44174 ( .A(n43364), .B(n43363), .Z(n43505) );
  XOR U44175 ( .A(n43506), .B(n43505), .Z(n43508) );
  NAND U44176 ( .A(x[490]), .B(y[8143]), .Z(n44331) );
  NANDN U44177 ( .A(n44331), .B(n43365), .Z(n43369) );
  NANDN U44178 ( .A(n43367), .B(n43366), .Z(n43368) );
  AND U44179 ( .A(n43369), .B(n43368), .Z(n43484) );
  AND U44180 ( .A(x[480]), .B(y[8146]), .Z(n43456) );
  AND U44181 ( .A(x[498]), .B(y[8128]), .Z(n43457) );
  XOR U44182 ( .A(n43456), .B(n43457), .Z(n43459) );
  AND U44183 ( .A(x[497]), .B(y[8129]), .Z(n43478) );
  XOR U44184 ( .A(o[466]), .B(n43478), .Z(n43458) );
  XOR U44185 ( .A(n43459), .B(n43458), .Z(n43482) );
  AND U44186 ( .A(y[8133]), .B(x[493]), .Z(n43371) );
  NAND U44187 ( .A(y[8143]), .B(x[483]), .Z(n43370) );
  XNOR U44188 ( .A(n43371), .B(n43370), .Z(n43464) );
  AND U44189 ( .A(x[492]), .B(y[8134]), .Z(n43465) );
  XOR U44190 ( .A(n43464), .B(n43465), .Z(n43481) );
  XOR U44191 ( .A(n43482), .B(n43481), .Z(n43483) );
  XOR U44192 ( .A(n43508), .B(n43507), .Z(n43428) );
  NANDN U44193 ( .A(n43373), .B(n43372), .Z(n43377) );
  NANDN U44194 ( .A(n43375), .B(n43374), .Z(n43376) );
  AND U44195 ( .A(n43377), .B(n43376), .Z(n43427) );
  NANDN U44196 ( .A(n43379), .B(n43378), .Z(n43383) );
  NANDN U44197 ( .A(n43381), .B(n43380), .Z(n43382) );
  NAND U44198 ( .A(n43383), .B(n43382), .Z(n43430) );
  XNOR U44199 ( .A(n43424), .B(n43423), .Z(n43418) );
  NANDN U44200 ( .A(n43385), .B(n43384), .Z(n43389) );
  NANDN U44201 ( .A(n43387), .B(n43386), .Z(n43388) );
  NAND U44202 ( .A(n43389), .B(n43388), .Z(n43416) );
  NAND U44203 ( .A(n43391), .B(n43390), .Z(n43395) );
  NAND U44204 ( .A(n43393), .B(n43392), .Z(n43394) );
  NAND U44205 ( .A(n43395), .B(n43394), .Z(n43415) );
  XOR U44206 ( .A(n43416), .B(n43415), .Z(n43417) );
  XNOR U44207 ( .A(n43418), .B(n43417), .Z(n43407) );
  XNOR U44208 ( .A(n43406), .B(n43407), .Z(n43408) );
  XNOR U44209 ( .A(n43409), .B(n43408), .Z(n43414) );
  NAND U44210 ( .A(n43400), .B(n43399), .Z(n43404) );
  NAND U44211 ( .A(n43402), .B(n43401), .Z(n43403) );
  NAND U44212 ( .A(n43404), .B(n43403), .Z(n43413) );
  XOR U44213 ( .A(n43412), .B(n43413), .Z(n43405) );
  XNOR U44214 ( .A(n43414), .B(n43405), .Z(N947) );
  NANDN U44215 ( .A(n43407), .B(n43406), .Z(n43411) );
  NAND U44216 ( .A(n43409), .B(n43408), .Z(n43410) );
  AND U44217 ( .A(n43411), .B(n43410), .Z(n43633) );
  NAND U44218 ( .A(n43416), .B(n43415), .Z(n43420) );
  NAND U44219 ( .A(n43418), .B(n43417), .Z(n43419) );
  NAND U44220 ( .A(n43420), .B(n43419), .Z(n43629) );
  NAND U44221 ( .A(n43422), .B(n43421), .Z(n43426) );
  NAND U44222 ( .A(n43424), .B(n43423), .Z(n43425) );
  AND U44223 ( .A(n43426), .B(n43425), .Z(n43627) );
  NANDN U44224 ( .A(n43428), .B(n43427), .Z(n43432) );
  NANDN U44225 ( .A(n43430), .B(n43429), .Z(n43431) );
  AND U44226 ( .A(n43432), .B(n43431), .Z(n43521) );
  AND U44227 ( .A(x[486]), .B(y[8141]), .Z(n43434) );
  NAND U44228 ( .A(n43434), .B(n43433), .Z(n43438) );
  NAND U44229 ( .A(n43436), .B(n43435), .Z(n43437) );
  AND U44230 ( .A(n43438), .B(n43437), .Z(n43611) );
  AND U44231 ( .A(x[496]), .B(y[8135]), .Z(n43966) );
  NAND U44232 ( .A(n43966), .B(n43789), .Z(n43442) );
  NANDN U44233 ( .A(n43440), .B(n43439), .Z(n43441) );
  AND U44234 ( .A(n43442), .B(n43441), .Z(n43609) );
  AND U44235 ( .A(x[495]), .B(y[8137]), .Z(n44217) );
  NAND U44236 ( .A(n44217), .B(n43536), .Z(n43446) );
  NAND U44237 ( .A(n43444), .B(n43443), .Z(n43445) );
  NAND U44238 ( .A(n43446), .B(n43445), .Z(n43533) );
  AND U44239 ( .A(y[8146]), .B(x[481]), .Z(n43448) );
  NAND U44240 ( .A(y[8139]), .B(x[488]), .Z(n43447) );
  XNOR U44241 ( .A(n43448), .B(n43447), .Z(n43587) );
  AND U44242 ( .A(y[8134]), .B(x[493]), .Z(n43450) );
  NAND U44243 ( .A(y[8145]), .B(x[482]), .Z(n43449) );
  XNOR U44244 ( .A(n43450), .B(n43449), .Z(n43542) );
  XOR U44245 ( .A(n43531), .B(n43530), .Z(n43532) );
  XOR U44246 ( .A(n43533), .B(n43532), .Z(n43608) );
  NAND U44247 ( .A(x[490]), .B(y[8145]), .Z(n44710) );
  NANDN U44248 ( .A(n44710), .B(n43451), .Z(n43455) );
  NAND U44249 ( .A(n43453), .B(n43452), .Z(n43454) );
  NAND U44250 ( .A(n43455), .B(n43454), .Z(n43567) );
  NAND U44251 ( .A(n43457), .B(n43456), .Z(n43461) );
  NAND U44252 ( .A(n43459), .B(n43458), .Z(n43460) );
  NAND U44253 ( .A(n43461), .B(n43460), .Z(n43565) );
  AND U44254 ( .A(y[8131]), .B(x[496]), .Z(n44268) );
  NAND U44255 ( .A(y[8138]), .B(x[489]), .Z(n43462) );
  XNOR U44256 ( .A(n44268), .B(n43462), .Z(n43537) );
  AND U44257 ( .A(x[495]), .B(y[8132]), .Z(n43538) );
  XOR U44258 ( .A(n43537), .B(n43538), .Z(n43564) );
  XOR U44259 ( .A(n43565), .B(n43564), .Z(n43566) );
  XNOR U44260 ( .A(n43567), .B(n43566), .Z(n43604) );
  AND U44261 ( .A(x[493]), .B(y[8143]), .Z(n44864) );
  NAND U44262 ( .A(n43463), .B(n44864), .Z(n43467) );
  NAND U44263 ( .A(n43465), .B(n43464), .Z(n43466) );
  NAND U44264 ( .A(n43467), .B(n43466), .Z(n43561) );
  AND U44265 ( .A(y[8137]), .B(x[490]), .Z(n43469) );
  NAND U44266 ( .A(y[8130]), .B(x[497]), .Z(n43468) );
  XNOR U44267 ( .A(n43469), .B(n43468), .Z(n43593) );
  AND U44268 ( .A(x[498]), .B(y[8129]), .Z(n43557) );
  XOR U44269 ( .A(o[467]), .B(n43557), .Z(n43592) );
  XOR U44270 ( .A(n43593), .B(n43592), .Z(n43559) );
  NAND U44271 ( .A(y[8144]), .B(x[483]), .Z(n43470) );
  XNOR U44272 ( .A(n43471), .B(n43470), .Z(n43551) );
  XOR U44273 ( .A(n43559), .B(n43558), .Z(n43560) );
  XNOR U44274 ( .A(n43561), .B(n43560), .Z(n43603) );
  NAND U44275 ( .A(n43473), .B(n43472), .Z(n43477) );
  NAND U44276 ( .A(n43475), .B(n43474), .Z(n43476) );
  AND U44277 ( .A(n43477), .B(n43476), .Z(n43527) );
  AND U44278 ( .A(x[480]), .B(y[8147]), .Z(n43574) );
  AND U44279 ( .A(x[499]), .B(y[8128]), .Z(n43575) );
  XOR U44280 ( .A(n43574), .B(n43575), .Z(n43577) );
  AND U44281 ( .A(o[466]), .B(n43478), .Z(n43576) );
  XOR U44282 ( .A(n43577), .B(n43576), .Z(n43525) );
  AND U44283 ( .A(x[484]), .B(y[8143]), .Z(n43702) );
  AND U44284 ( .A(y[8142]), .B(x[485]), .Z(n43480) );
  NAND U44285 ( .A(y[8141]), .B(x[486]), .Z(n43479) );
  XNOR U44286 ( .A(n43480), .B(n43479), .Z(n43571) );
  XOR U44287 ( .A(n43702), .B(n43571), .Z(n43524) );
  XOR U44288 ( .A(n43525), .B(n43524), .Z(n43526) );
  XOR U44289 ( .A(n43527), .B(n43526), .Z(n43602) );
  XOR U44290 ( .A(n43603), .B(n43602), .Z(n43605) );
  XNOR U44291 ( .A(n43604), .B(n43605), .Z(n43598) );
  NAND U44292 ( .A(n43482), .B(n43481), .Z(n43486) );
  NANDN U44293 ( .A(n43484), .B(n43483), .Z(n43485) );
  AND U44294 ( .A(n43486), .B(n43485), .Z(n43597) );
  NAND U44295 ( .A(n43488), .B(n43487), .Z(n43492) );
  NANDN U44296 ( .A(n43490), .B(n43489), .Z(n43491) );
  NAND U44297 ( .A(n43492), .B(n43491), .Z(n43596) );
  XNOR U44298 ( .A(n43598), .B(n43599), .Z(n43518) );
  XOR U44299 ( .A(n43519), .B(n43518), .Z(n43520) );
  NAND U44300 ( .A(n43494), .B(n43493), .Z(n43498) );
  NAND U44301 ( .A(n43496), .B(n43495), .Z(n43497) );
  AND U44302 ( .A(n43498), .B(n43497), .Z(n43620) );
  NAND U44303 ( .A(n43500), .B(n43499), .Z(n43504) );
  NAND U44304 ( .A(n43502), .B(n43501), .Z(n43503) );
  NAND U44305 ( .A(n43504), .B(n43503), .Z(n43616) );
  NAND U44306 ( .A(n43506), .B(n43505), .Z(n43510) );
  NAND U44307 ( .A(n43508), .B(n43507), .Z(n43509) );
  NAND U44308 ( .A(n43510), .B(n43509), .Z(n43615) );
  NAND U44309 ( .A(n43512), .B(n43511), .Z(n43516) );
  NAND U44310 ( .A(n43514), .B(n43513), .Z(n43515) );
  NAND U44311 ( .A(n43516), .B(n43515), .Z(n43614) );
  XNOR U44312 ( .A(n43615), .B(n43614), .Z(n43617) );
  XNOR U44313 ( .A(n43620), .B(n43621), .Z(n43622) );
  XOR U44314 ( .A(n43627), .B(n43626), .Z(n43628) );
  XOR U44315 ( .A(n43629), .B(n43628), .Z(n43634) );
  XOR U44316 ( .A(n43632), .B(n43634), .Z(n43517) );
  XOR U44317 ( .A(n43633), .B(n43517), .Z(N948) );
  NAND U44318 ( .A(n43519), .B(n43518), .Z(n43523) );
  NANDN U44319 ( .A(n43521), .B(n43520), .Z(n43522) );
  AND U44320 ( .A(n43523), .B(n43522), .Z(n43740) );
  NAND U44321 ( .A(n43525), .B(n43524), .Z(n43529) );
  NANDN U44322 ( .A(n43527), .B(n43526), .Z(n43528) );
  NAND U44323 ( .A(n43529), .B(n43528), .Z(n43637) );
  NAND U44324 ( .A(n43531), .B(n43530), .Z(n43535) );
  NAND U44325 ( .A(n43533), .B(n43532), .Z(n43534) );
  NAND U44326 ( .A(n43535), .B(n43534), .Z(n43636) );
  XOR U44327 ( .A(n43637), .B(n43636), .Z(n43639) );
  AND U44328 ( .A(x[496]), .B(y[8138]), .Z(n44493) );
  NAND U44329 ( .A(n44493), .B(n43536), .Z(n43540) );
  NAND U44330 ( .A(n43538), .B(n43537), .Z(n43539) );
  NAND U44331 ( .A(n43540), .B(n43539), .Z(n43677) );
  AND U44332 ( .A(x[493]), .B(y[8145]), .Z(n45099) );
  NAND U44333 ( .A(n45099), .B(n43541), .Z(n43545) );
  NANDN U44334 ( .A(n43543), .B(n43542), .Z(n43544) );
  NAND U44335 ( .A(n43545), .B(n43544), .Z(n43722) );
  AND U44336 ( .A(y[8132]), .B(x[496]), .Z(n43547) );
  NAND U44337 ( .A(y[8138]), .B(x[490]), .Z(n43546) );
  XNOR U44338 ( .A(n43547), .B(n43546), .Z(n43683) );
  AND U44339 ( .A(x[482]), .B(y[8146]), .Z(n43684) );
  XOR U44340 ( .A(n43683), .B(n43684), .Z(n43720) );
  NAND U44341 ( .A(y[8139]), .B(x[489]), .Z(n43548) );
  XNOR U44342 ( .A(n43549), .B(n43548), .Z(n43659) );
  AND U44343 ( .A(x[494]), .B(y[8134]), .Z(n43660) );
  XOR U44344 ( .A(n43659), .B(n43660), .Z(n43719) );
  XOR U44345 ( .A(n43720), .B(n43719), .Z(n43721) );
  XOR U44346 ( .A(n43722), .B(n43721), .Z(n43676) );
  XOR U44347 ( .A(n43677), .B(n43676), .Z(n43679) );
  NAND U44348 ( .A(x[491]), .B(y[8144]), .Z(n44712) );
  NANDN U44349 ( .A(n44712), .B(n43550), .Z(n43554) );
  NANDN U44350 ( .A(n43552), .B(n43551), .Z(n43553) );
  NAND U44351 ( .A(n43554), .B(n43553), .Z(n43728) );
  AND U44352 ( .A(y[8137]), .B(x[491]), .Z(n43556) );
  NAND U44353 ( .A(y[8147]), .B(x[481]), .Z(n43555) );
  XNOR U44354 ( .A(n43556), .B(n43555), .Z(n43655) );
  AND U44355 ( .A(x[499]), .B(y[8129]), .Z(n43663) );
  XOR U44356 ( .A(o[468]), .B(n43663), .Z(n43654) );
  XOR U44357 ( .A(n43655), .B(n43654), .Z(n43726) );
  AND U44358 ( .A(x[480]), .B(y[8148]), .Z(n43707) );
  AND U44359 ( .A(x[500]), .B(y[8128]), .Z(n43708) );
  XOR U44360 ( .A(n43707), .B(n43708), .Z(n43710) );
  AND U44361 ( .A(o[467]), .B(n43557), .Z(n43709) );
  XOR U44362 ( .A(n43710), .B(n43709), .Z(n43725) );
  XOR U44363 ( .A(n43726), .B(n43725), .Z(n43727) );
  XOR U44364 ( .A(n43728), .B(n43727), .Z(n43678) );
  XOR U44365 ( .A(n43679), .B(n43678), .Z(n43638) );
  XNOR U44366 ( .A(n43639), .B(n43638), .Z(n43734) );
  NAND U44367 ( .A(n43559), .B(n43558), .Z(n43563) );
  NAND U44368 ( .A(n43561), .B(n43560), .Z(n43562) );
  AND U44369 ( .A(n43563), .B(n43562), .Z(n43732) );
  NAND U44370 ( .A(n43565), .B(n43564), .Z(n43569) );
  NAND U44371 ( .A(n43567), .B(n43566), .Z(n43568) );
  AND U44372 ( .A(n43569), .B(n43568), .Z(n43673) );
  NAND U44373 ( .A(x[486]), .B(y[8142]), .Z(n43643) );
  NANDN U44374 ( .A(n43643), .B(n43570), .Z(n43573) );
  NAND U44375 ( .A(n43571), .B(n43702), .Z(n43572) );
  NAND U44376 ( .A(n43573), .B(n43572), .Z(n43667) );
  NAND U44377 ( .A(n43575), .B(n43574), .Z(n43579) );
  NAND U44378 ( .A(n43577), .B(n43576), .Z(n43578) );
  NAND U44379 ( .A(n43579), .B(n43578), .Z(n43665) );
  AND U44380 ( .A(y[8130]), .B(x[498]), .Z(n43581) );
  NAND U44381 ( .A(y[8136]), .B(x[492]), .Z(n43580) );
  XNOR U44382 ( .A(n43581), .B(n43580), .Z(n43649) );
  AND U44383 ( .A(x[497]), .B(y[8131]), .Z(n43650) );
  XOR U44384 ( .A(n43649), .B(n43650), .Z(n43664) );
  XOR U44385 ( .A(n43665), .B(n43664), .Z(n43666) );
  XNOR U44386 ( .A(n43667), .B(n43666), .Z(n43671) );
  AND U44387 ( .A(y[8135]), .B(x[493]), .Z(n43583) );
  NAND U44388 ( .A(y[8145]), .B(x[483]), .Z(n43582) );
  XNOR U44389 ( .A(n43583), .B(n43582), .Z(n43689) );
  XNOR U44390 ( .A(n43689), .B(n43688), .Z(n43645) );
  AND U44391 ( .A(y[8143]), .B(x[485]), .Z(n43585) );
  NAND U44392 ( .A(y[8144]), .B(x[484]), .Z(n43584) );
  XNOR U44393 ( .A(n43585), .B(n43584), .Z(n43704) );
  AND U44394 ( .A(x[487]), .B(y[8141]), .Z(n43703) );
  XNOR U44395 ( .A(n43704), .B(n43703), .Z(n43642) );
  XOR U44396 ( .A(n43643), .B(n43642), .Z(n43644) );
  XNOR U44397 ( .A(n43645), .B(n43644), .Z(n43715) );
  AND U44398 ( .A(x[488]), .B(y[8146]), .Z(n44817) );
  AND U44399 ( .A(x[481]), .B(y[8139]), .Z(n43586) );
  NAND U44400 ( .A(n44817), .B(n43586), .Z(n43590) );
  NANDN U44401 ( .A(n43588), .B(n43587), .Z(n43589) );
  NAND U44402 ( .A(n43590), .B(n43589), .Z(n43714) );
  AND U44403 ( .A(x[497]), .B(y[8137]), .Z(n44501) );
  NAND U44404 ( .A(n44501), .B(n43591), .Z(n43595) );
  NAND U44405 ( .A(n43593), .B(n43592), .Z(n43594) );
  NAND U44406 ( .A(n43595), .B(n43594), .Z(n43713) );
  XOR U44407 ( .A(n43714), .B(n43713), .Z(n43716) );
  XNOR U44408 ( .A(n43715), .B(n43716), .Z(n43670) );
  XOR U44409 ( .A(n43671), .B(n43670), .Z(n43672) );
  XOR U44410 ( .A(n43673), .B(n43672), .Z(n43731) );
  XOR U44411 ( .A(n43732), .B(n43731), .Z(n43733) );
  XNOR U44412 ( .A(n43734), .B(n43733), .Z(n43738) );
  NANDN U44413 ( .A(n43597), .B(n43596), .Z(n43601) );
  NAND U44414 ( .A(n43599), .B(n43598), .Z(n43600) );
  AND U44415 ( .A(n43601), .B(n43600), .Z(n43746) );
  NAND U44416 ( .A(n43603), .B(n43602), .Z(n43607) );
  NAND U44417 ( .A(n43605), .B(n43604), .Z(n43606) );
  AND U44418 ( .A(n43607), .B(n43606), .Z(n43744) );
  NANDN U44419 ( .A(n43609), .B(n43608), .Z(n43613) );
  NANDN U44420 ( .A(n43611), .B(n43610), .Z(n43612) );
  AND U44421 ( .A(n43613), .B(n43612), .Z(n43743) );
  XNOR U44422 ( .A(n43746), .B(n43745), .Z(n43737) );
  XOR U44423 ( .A(n43738), .B(n43737), .Z(n43739) );
  XOR U44424 ( .A(n43740), .B(n43739), .Z(n43755) );
  NAND U44425 ( .A(n43615), .B(n43614), .Z(n43619) );
  NANDN U44426 ( .A(n43617), .B(n43616), .Z(n43618) );
  AND U44427 ( .A(n43619), .B(n43618), .Z(n43753) );
  NANDN U44428 ( .A(n43621), .B(n43620), .Z(n43625) );
  NANDN U44429 ( .A(n43623), .B(n43622), .Z(n43624) );
  AND U44430 ( .A(n43625), .B(n43624), .Z(n43752) );
  XOR U44431 ( .A(n43753), .B(n43752), .Z(n43754) );
  NAND U44432 ( .A(n43627), .B(n43626), .Z(n43631) );
  NAND U44433 ( .A(n43629), .B(n43628), .Z(n43630) );
  NAND U44434 ( .A(n43631), .B(n43630), .Z(n43750) );
  XOR U44435 ( .A(n43750), .B(n43749), .Z(n43635) );
  XNOR U44436 ( .A(n43751), .B(n43635), .Z(N949) );
  NAND U44437 ( .A(n43637), .B(n43636), .Z(n43641) );
  NAND U44438 ( .A(n43639), .B(n43638), .Z(n43640) );
  NAND U44439 ( .A(n43641), .B(n43640), .Z(n43768) );
  NAND U44440 ( .A(n43643), .B(n43642), .Z(n43647) );
  NAND U44441 ( .A(n43645), .B(n43644), .Z(n43646) );
  NAND U44442 ( .A(n43647), .B(n43646), .Z(n43839) );
  AND U44443 ( .A(x[498]), .B(y[8136]), .Z(n44500) );
  NAND U44444 ( .A(n44500), .B(n43648), .Z(n43652) );
  NAND U44445 ( .A(n43650), .B(n43649), .Z(n43651) );
  NAND U44446 ( .A(n43652), .B(n43651), .Z(n43845) );
  AND U44447 ( .A(x[491]), .B(y[8147]), .Z(n45278) );
  AND U44448 ( .A(x[481]), .B(y[8137]), .Z(n43653) );
  NAND U44449 ( .A(n45278), .B(n43653), .Z(n43657) );
  NAND U44450 ( .A(n43655), .B(n43654), .Z(n43656) );
  NAND U44451 ( .A(n43657), .B(n43656), .Z(n43844) );
  XOR U44452 ( .A(n43845), .B(n43844), .Z(n43847) );
  AND U44453 ( .A(x[495]), .B(y[8139]), .Z(n44488) );
  NAND U44454 ( .A(n44488), .B(n43658), .Z(n43662) );
  NAND U44455 ( .A(n43660), .B(n43659), .Z(n43661) );
  NAND U44456 ( .A(n43662), .B(n43661), .Z(n43803) );
  AND U44457 ( .A(o[468]), .B(n43663), .Z(n43825) );
  AND U44458 ( .A(x[480]), .B(y[8149]), .Z(n43822) );
  AND U44459 ( .A(x[501]), .B(y[8128]), .Z(n43823) );
  XOR U44460 ( .A(n43822), .B(n43823), .Z(n43824) );
  XOR U44461 ( .A(n43825), .B(n43824), .Z(n43801) );
  AND U44462 ( .A(x[485]), .B(y[8144]), .Z(n43809) );
  AND U44463 ( .A(x[496]), .B(y[8133]), .Z(n43808) );
  XOR U44464 ( .A(n43809), .B(n43808), .Z(n43807) );
  AND U44465 ( .A(x[495]), .B(y[8134]), .Z(n43806) );
  XOR U44466 ( .A(n43807), .B(n43806), .Z(n43800) );
  XOR U44467 ( .A(n43801), .B(n43800), .Z(n43802) );
  XOR U44468 ( .A(n43803), .B(n43802), .Z(n43846) );
  XNOR U44469 ( .A(n43847), .B(n43846), .Z(n43838) );
  XOR U44470 ( .A(n43839), .B(n43838), .Z(n43841) );
  NAND U44471 ( .A(n43665), .B(n43664), .Z(n43669) );
  NAND U44472 ( .A(n43667), .B(n43666), .Z(n43668) );
  AND U44473 ( .A(n43669), .B(n43668), .Z(n43840) );
  XNOR U44474 ( .A(n43841), .B(n43840), .Z(n43766) );
  NAND U44475 ( .A(n43671), .B(n43670), .Z(n43675) );
  NAND U44476 ( .A(n43673), .B(n43672), .Z(n43674) );
  AND U44477 ( .A(n43675), .B(n43674), .Z(n43765) );
  XOR U44478 ( .A(n43766), .B(n43765), .Z(n43767) );
  XNOR U44479 ( .A(n43768), .B(n43767), .Z(n43761) );
  NAND U44480 ( .A(n43677), .B(n43676), .Z(n43681) );
  NAND U44481 ( .A(n43679), .B(n43678), .Z(n43680) );
  NAND U44482 ( .A(n43681), .B(n43680), .Z(n43865) );
  AND U44483 ( .A(x[490]), .B(y[8132]), .Z(n43682) );
  NAND U44484 ( .A(n44493), .B(n43682), .Z(n43686) );
  NAND U44485 ( .A(n43684), .B(n43683), .Z(n43685) );
  NAND U44486 ( .A(n43686), .B(n43685), .Z(n43772) );
  NAND U44487 ( .A(n45099), .B(n43687), .Z(n43691) );
  NAND U44488 ( .A(n43689), .B(n43688), .Z(n43690) );
  NAND U44489 ( .A(n43691), .B(n43690), .Z(n43859) );
  AND U44490 ( .A(y[8130]), .B(x[499]), .Z(n43693) );
  NAND U44491 ( .A(y[8138]), .B(x[491]), .Z(n43692) );
  XNOR U44492 ( .A(n43693), .B(n43692), .Z(n43791) );
  AND U44493 ( .A(x[500]), .B(y[8129]), .Z(n43821) );
  XOR U44494 ( .A(o[469]), .B(n43821), .Z(n43790) );
  XOR U44495 ( .A(n43791), .B(n43790), .Z(n43857) );
  AND U44496 ( .A(y[8131]), .B(x[498]), .Z(n43695) );
  NAND U44497 ( .A(y[8139]), .B(x[490]), .Z(n43694) );
  XNOR U44498 ( .A(n43695), .B(n43694), .Z(n43829) );
  AND U44499 ( .A(x[481]), .B(y[8148]), .Z(n43830) );
  XOR U44500 ( .A(n43829), .B(n43830), .Z(n43856) );
  XOR U44501 ( .A(n43857), .B(n43856), .Z(n43858) );
  XOR U44502 ( .A(n43859), .B(n43858), .Z(n43771) );
  XOR U44503 ( .A(n43772), .B(n43771), .Z(n43774) );
  AND U44504 ( .A(x[487]), .B(y[8142]), .Z(n44042) );
  AND U44505 ( .A(y[8143]), .B(x[486]), .Z(n43697) );
  NAND U44506 ( .A(y[8135]), .B(x[494]), .Z(n43696) );
  XNOR U44507 ( .A(n43697), .B(n43696), .Z(n43833) );
  XNOR U44508 ( .A(n44042), .B(n43833), .Z(n43780) );
  NAND U44509 ( .A(x[489]), .B(y[8140]), .Z(n43778) );
  NAND U44510 ( .A(x[488]), .B(y[8141]), .Z(n43777) );
  XOR U44511 ( .A(n43778), .B(n43777), .Z(n43779) );
  XNOR U44512 ( .A(n43780), .B(n43779), .Z(n43796) );
  AND U44513 ( .A(y[8137]), .B(x[492]), .Z(n43699) );
  NAND U44514 ( .A(y[8132]), .B(x[497]), .Z(n43698) );
  XNOR U44515 ( .A(n43699), .B(n43698), .Z(n43783) );
  AND U44516 ( .A(x[482]), .B(y[8147]), .Z(n43784) );
  XOR U44517 ( .A(n43783), .B(n43784), .Z(n43795) );
  AND U44518 ( .A(y[8136]), .B(x[493]), .Z(n43701) );
  NAND U44519 ( .A(y[8146]), .B(x[483]), .Z(n43700) );
  XNOR U44520 ( .A(n43701), .B(n43700), .Z(n43817) );
  AND U44521 ( .A(x[484]), .B(y[8145]), .Z(n43818) );
  XOR U44522 ( .A(n43817), .B(n43818), .Z(n43794) );
  XOR U44523 ( .A(n43795), .B(n43794), .Z(n43797) );
  XOR U44524 ( .A(n43796), .B(n43797), .Z(n43853) );
  NAND U44525 ( .A(n43702), .B(n43809), .Z(n43706) );
  NAND U44526 ( .A(n43704), .B(n43703), .Z(n43705) );
  NAND U44527 ( .A(n43706), .B(n43705), .Z(n43851) );
  NAND U44528 ( .A(n43708), .B(n43707), .Z(n43712) );
  NAND U44529 ( .A(n43710), .B(n43709), .Z(n43711) );
  NAND U44530 ( .A(n43712), .B(n43711), .Z(n43850) );
  XOR U44531 ( .A(n43851), .B(n43850), .Z(n43852) );
  XOR U44532 ( .A(n43853), .B(n43852), .Z(n43773) );
  XOR U44533 ( .A(n43774), .B(n43773), .Z(n43863) );
  NAND U44534 ( .A(n43714), .B(n43713), .Z(n43718) );
  NAND U44535 ( .A(n43716), .B(n43715), .Z(n43717) );
  NAND U44536 ( .A(n43718), .B(n43717), .Z(n43870) );
  NAND U44537 ( .A(n43720), .B(n43719), .Z(n43724) );
  NAND U44538 ( .A(n43722), .B(n43721), .Z(n43723) );
  NAND U44539 ( .A(n43724), .B(n43723), .Z(n43869) );
  NAND U44540 ( .A(n43726), .B(n43725), .Z(n43730) );
  NAND U44541 ( .A(n43728), .B(n43727), .Z(n43729) );
  NAND U44542 ( .A(n43730), .B(n43729), .Z(n43868) );
  XOR U44543 ( .A(n43869), .B(n43868), .Z(n43871) );
  XOR U44544 ( .A(n43870), .B(n43871), .Z(n43862) );
  XOR U44545 ( .A(n43863), .B(n43862), .Z(n43864) );
  XNOR U44546 ( .A(n43865), .B(n43864), .Z(n43760) );
  NAND U44547 ( .A(n43732), .B(n43731), .Z(n43736) );
  NAND U44548 ( .A(n43734), .B(n43733), .Z(n43735) );
  NAND U44549 ( .A(n43736), .B(n43735), .Z(n43759) );
  XOR U44550 ( .A(n43760), .B(n43759), .Z(n43762) );
  XNOR U44551 ( .A(n43761), .B(n43762), .Z(n43883) );
  NAND U44552 ( .A(n43738), .B(n43737), .Z(n43742) );
  NAND U44553 ( .A(n43740), .B(n43739), .Z(n43741) );
  AND U44554 ( .A(n43742), .B(n43741), .Z(n43882) );
  NANDN U44555 ( .A(n43744), .B(n43743), .Z(n43748) );
  NAND U44556 ( .A(n43746), .B(n43745), .Z(n43747) );
  AND U44557 ( .A(n43748), .B(n43747), .Z(n43881) );
  XNOR U44558 ( .A(n43883), .B(n43884), .Z(n43877) );
  NAND U44559 ( .A(n43753), .B(n43752), .Z(n43757) );
  NANDN U44560 ( .A(n43755), .B(n43754), .Z(n43756) );
  AND U44561 ( .A(n43757), .B(n43756), .Z(n43875) );
  IV U44562 ( .A(n43875), .Z(n43874) );
  XOR U44563 ( .A(n43876), .B(n43874), .Z(n43758) );
  XNOR U44564 ( .A(n43877), .B(n43758), .Z(N950) );
  NAND U44565 ( .A(n43760), .B(n43759), .Z(n43764) );
  NAND U44566 ( .A(n43762), .B(n43761), .Z(n43763) );
  AND U44567 ( .A(n43764), .B(n43763), .Z(n44018) );
  NAND U44568 ( .A(n43766), .B(n43765), .Z(n43770) );
  NAND U44569 ( .A(n43768), .B(n43767), .Z(n43769) );
  NAND U44570 ( .A(n43770), .B(n43769), .Z(n44016) );
  NAND U44571 ( .A(n43772), .B(n43771), .Z(n43776) );
  NAND U44572 ( .A(n43774), .B(n43773), .Z(n43775) );
  NAND U44573 ( .A(n43776), .B(n43775), .Z(n44004) );
  NAND U44574 ( .A(n43778), .B(n43777), .Z(n43782) );
  NAND U44575 ( .A(n43780), .B(n43779), .Z(n43781) );
  NAND U44576 ( .A(n43782), .B(n43781), .Z(n43999) );
  NAND U44577 ( .A(n44501), .B(n43950), .Z(n43786) );
  NAND U44578 ( .A(n43784), .B(n43783), .Z(n43785) );
  NAND U44579 ( .A(n43786), .B(n43785), .Z(n43926) );
  AND U44580 ( .A(x[485]), .B(y[8145]), .Z(n43972) );
  AND U44581 ( .A(x[497]), .B(y[8133]), .Z(n43973) );
  XOR U44582 ( .A(n43972), .B(n43973), .Z(n43974) );
  AND U44583 ( .A(x[496]), .B(y[8134]), .Z(n43975) );
  XOR U44584 ( .A(n43974), .B(n43975), .Z(n43925) );
  AND U44585 ( .A(y[8132]), .B(x[498]), .Z(n43788) );
  NAND U44586 ( .A(y[8138]), .B(x[492]), .Z(n43787) );
  XNOR U44587 ( .A(n43788), .B(n43787), .Z(n43951) );
  AND U44588 ( .A(x[484]), .B(y[8146]), .Z(n43952) );
  XOR U44589 ( .A(n43951), .B(n43952), .Z(n43924) );
  XOR U44590 ( .A(n43925), .B(n43924), .Z(n43927) );
  XNOR U44591 ( .A(n43926), .B(n43927), .Z(n43996) );
  AND U44592 ( .A(x[499]), .B(y[8138]), .Z(n44990) );
  NAND U44593 ( .A(n44990), .B(n43789), .Z(n43793) );
  NAND U44594 ( .A(n43791), .B(n43790), .Z(n43792) );
  AND U44595 ( .A(n43793), .B(n43792), .Z(n43997) );
  XOR U44596 ( .A(n43996), .B(n43997), .Z(n43998) );
  XNOR U44597 ( .A(n43999), .B(n43998), .Z(n44003) );
  NAND U44598 ( .A(n43795), .B(n43794), .Z(n43799) );
  NAND U44599 ( .A(n43797), .B(n43796), .Z(n43798) );
  NAND U44600 ( .A(n43799), .B(n43798), .Z(n43985) );
  NAND U44601 ( .A(n43801), .B(n43800), .Z(n43805) );
  NAND U44602 ( .A(n43803), .B(n43802), .Z(n43804) );
  NAND U44603 ( .A(n43805), .B(n43804), .Z(n43984) );
  XOR U44604 ( .A(n43985), .B(n43984), .Z(n43987) );
  AND U44605 ( .A(n43807), .B(n43806), .Z(n43811) );
  NAND U44606 ( .A(n43809), .B(n43808), .Z(n43810) );
  NANDN U44607 ( .A(n43811), .B(n43810), .Z(n43947) );
  AND U44608 ( .A(y[8137]), .B(x[493]), .Z(n43813) );
  NAND U44609 ( .A(y[8130]), .B(x[500]), .Z(n43812) );
  XNOR U44610 ( .A(n43813), .B(n43812), .Z(n43968) );
  AND U44611 ( .A(x[482]), .B(y[8148]), .Z(n43969) );
  XOR U44612 ( .A(n43968), .B(n43969), .Z(n43945) );
  AND U44613 ( .A(y[8144]), .B(x[486]), .Z(n43815) );
  NAND U44614 ( .A(y[8135]), .B(x[495]), .Z(n43814) );
  XNOR U44615 ( .A(n43815), .B(n43814), .Z(n43981) );
  XOR U44616 ( .A(n43980), .B(n43981), .Z(n43944) );
  XOR U44617 ( .A(n43945), .B(n43944), .Z(n43946) );
  XOR U44618 ( .A(n43947), .B(n43946), .Z(n43991) );
  AND U44619 ( .A(x[493]), .B(y[8146]), .Z(n45279) );
  NANDN U44620 ( .A(n43816), .B(n45279), .Z(n43820) );
  NAND U44621 ( .A(n43818), .B(n43817), .Z(n43819) );
  NAND U44622 ( .A(n43820), .B(n43819), .Z(n43915) );
  AND U44623 ( .A(x[481]), .B(y[8149]), .Z(n43938) );
  XOR U44624 ( .A(n43939), .B(n43938), .Z(n43937) );
  AND U44625 ( .A(o[469]), .B(n43821), .Z(n43936) );
  XOR U44626 ( .A(n43937), .B(n43936), .Z(n43913) );
  AND U44627 ( .A(x[494]), .B(y[8136]), .Z(n43930) );
  AND U44628 ( .A(x[483]), .B(y[8147]), .Z(n43931) );
  XOR U44629 ( .A(n43930), .B(n43931), .Z(n43932) );
  AND U44630 ( .A(x[499]), .B(y[8131]), .Z(n43933) );
  XOR U44631 ( .A(n43932), .B(n43933), .Z(n43912) );
  XOR U44632 ( .A(n43913), .B(n43912), .Z(n43914) );
  XOR U44633 ( .A(n43915), .B(n43914), .Z(n43990) );
  XOR U44634 ( .A(n43991), .B(n43990), .Z(n43993) );
  NAND U44635 ( .A(n43823), .B(n43822), .Z(n43827) );
  NAND U44636 ( .A(n43825), .B(n43824), .Z(n43826) );
  NAND U44637 ( .A(n43827), .B(n43826), .Z(n43907) );
  AND U44638 ( .A(x[498]), .B(y[8139]), .Z(n44993) );
  NAND U44639 ( .A(n44993), .B(n43828), .Z(n43832) );
  NAND U44640 ( .A(n43830), .B(n43829), .Z(n43831) );
  NAND U44641 ( .A(n43832), .B(n43831), .Z(n43906) );
  XOR U44642 ( .A(n43907), .B(n43906), .Z(n43909) );
  AND U44643 ( .A(x[494]), .B(y[8143]), .Z(n45003) );
  NAND U44644 ( .A(n45003), .B(n43979), .Z(n43835) );
  NAND U44645 ( .A(n44042), .B(n43833), .Z(n43834) );
  NAND U44646 ( .A(n43835), .B(n43834), .Z(n43921) );
  AND U44647 ( .A(x[480]), .B(y[8150]), .Z(n43955) );
  AND U44648 ( .A(x[502]), .B(y[8128]), .Z(n43956) );
  XOR U44649 ( .A(n43955), .B(n43956), .Z(n43958) );
  AND U44650 ( .A(x[501]), .B(y[8129]), .Z(n43978) );
  XOR U44651 ( .A(o[470]), .B(n43978), .Z(n43957) );
  XOR U44652 ( .A(n43958), .B(n43957), .Z(n43919) );
  AND U44653 ( .A(y[8143]), .B(x[487]), .Z(n43837) );
  NAND U44654 ( .A(y[8142]), .B(x[488]), .Z(n43836) );
  XNOR U44655 ( .A(n43837), .B(n43836), .Z(n43962) );
  XOR U44656 ( .A(n43961), .B(n43962), .Z(n43918) );
  XOR U44657 ( .A(n43919), .B(n43918), .Z(n43920) );
  XOR U44658 ( .A(n43921), .B(n43920), .Z(n43908) );
  XOR U44659 ( .A(n43909), .B(n43908), .Z(n43992) );
  XOR U44660 ( .A(n43993), .B(n43992), .Z(n43986) );
  XOR U44661 ( .A(n43987), .B(n43986), .Z(n44002) );
  XOR U44662 ( .A(n44003), .B(n44002), .Z(n44005) );
  XNOR U44663 ( .A(n44004), .B(n44005), .Z(n43897) );
  NAND U44664 ( .A(n43839), .B(n43838), .Z(n43843) );
  NAND U44665 ( .A(n43841), .B(n43840), .Z(n43842) );
  NAND U44666 ( .A(n43843), .B(n43842), .Z(n43895) );
  NAND U44667 ( .A(n43845), .B(n43844), .Z(n43849) );
  NAND U44668 ( .A(n43847), .B(n43846), .Z(n43848) );
  AND U44669 ( .A(n43849), .B(n43848), .Z(n43903) );
  NAND U44670 ( .A(n43851), .B(n43850), .Z(n43855) );
  NAND U44671 ( .A(n43853), .B(n43852), .Z(n43854) );
  NAND U44672 ( .A(n43855), .B(n43854), .Z(n43901) );
  NAND U44673 ( .A(n43857), .B(n43856), .Z(n43861) );
  NAND U44674 ( .A(n43859), .B(n43858), .Z(n43860) );
  NAND U44675 ( .A(n43861), .B(n43860), .Z(n43900) );
  XOR U44676 ( .A(n43901), .B(n43900), .Z(n43902) );
  XOR U44677 ( .A(n43903), .B(n43902), .Z(n43894) );
  XOR U44678 ( .A(n43895), .B(n43894), .Z(n43896) );
  XNOR U44679 ( .A(n43897), .B(n43896), .Z(n43891) );
  NAND U44680 ( .A(n43863), .B(n43862), .Z(n43867) );
  NAND U44681 ( .A(n43865), .B(n43864), .Z(n43866) );
  NAND U44682 ( .A(n43867), .B(n43866), .Z(n43889) );
  NAND U44683 ( .A(n43869), .B(n43868), .Z(n43873) );
  NAND U44684 ( .A(n43871), .B(n43870), .Z(n43872) );
  NAND U44685 ( .A(n43873), .B(n43872), .Z(n43888) );
  XOR U44686 ( .A(n43889), .B(n43888), .Z(n43890) );
  XOR U44687 ( .A(n43891), .B(n43890), .Z(n44015) );
  XOR U44688 ( .A(n44016), .B(n44015), .Z(n44017) );
  XNOR U44689 ( .A(n44018), .B(n44017), .Z(n44011) );
  OR U44690 ( .A(n43876), .B(n43874), .Z(n43880) );
  ANDN U44691 ( .B(n43876), .A(n43875), .Z(n43878) );
  OR U44692 ( .A(n43878), .B(n43877), .Z(n43879) );
  AND U44693 ( .A(n43880), .B(n43879), .Z(n44010) );
  NANDN U44694 ( .A(n43882), .B(n43881), .Z(n43886) );
  NAND U44695 ( .A(n43884), .B(n43883), .Z(n43885) );
  NAND U44696 ( .A(n43886), .B(n43885), .Z(n44009) );
  IV U44697 ( .A(n44009), .Z(n44008) );
  XOR U44698 ( .A(n44010), .B(n44008), .Z(n43887) );
  XNOR U44699 ( .A(n44011), .B(n43887), .Z(N951) );
  NAND U44700 ( .A(n43889), .B(n43888), .Z(n43893) );
  NAND U44701 ( .A(n43891), .B(n43890), .Z(n43892) );
  AND U44702 ( .A(n43893), .B(n43892), .Z(n44163) );
  NAND U44703 ( .A(n43895), .B(n43894), .Z(n43899) );
  NAND U44704 ( .A(n43897), .B(n43896), .Z(n43898) );
  NAND U44705 ( .A(n43899), .B(n43898), .Z(n44160) );
  NAND U44706 ( .A(n43901), .B(n43900), .Z(n43905) );
  NANDN U44707 ( .A(n43903), .B(n43902), .Z(n43904) );
  NAND U44708 ( .A(n43905), .B(n43904), .Z(n44138) );
  NAND U44709 ( .A(n43907), .B(n43906), .Z(n43911) );
  NAND U44710 ( .A(n43909), .B(n43908), .Z(n43910) );
  NAND U44711 ( .A(n43911), .B(n43910), .Z(n44132) );
  NAND U44712 ( .A(n43913), .B(n43912), .Z(n43917) );
  NAND U44713 ( .A(n43915), .B(n43914), .Z(n43916) );
  NAND U44714 ( .A(n43917), .B(n43916), .Z(n44130) );
  NAND U44715 ( .A(n43919), .B(n43918), .Z(n43923) );
  NAND U44716 ( .A(n43921), .B(n43920), .Z(n43922) );
  NAND U44717 ( .A(n43923), .B(n43922), .Z(n44129) );
  XOR U44718 ( .A(n44130), .B(n44129), .Z(n44131) );
  XOR U44719 ( .A(n44132), .B(n44131), .Z(n44150) );
  NAND U44720 ( .A(n43925), .B(n43924), .Z(n43929) );
  NAND U44721 ( .A(n43927), .B(n43926), .Z(n43928) );
  NAND U44722 ( .A(n43929), .B(n43928), .Z(n44148) );
  NAND U44723 ( .A(n43931), .B(n43930), .Z(n43935) );
  NAND U44724 ( .A(n43933), .B(n43932), .Z(n43934) );
  NAND U44725 ( .A(n43935), .B(n43934), .Z(n44076) );
  AND U44726 ( .A(n43937), .B(n43936), .Z(n43941) );
  NAND U44727 ( .A(n43939), .B(n43938), .Z(n43940) );
  NANDN U44728 ( .A(n43941), .B(n43940), .Z(n44075) );
  XOR U44729 ( .A(n44076), .B(n44075), .Z(n44078) );
  AND U44730 ( .A(y[8144]), .B(x[487]), .Z(n43943) );
  NAND U44731 ( .A(y[8142]), .B(x[489]), .Z(n43942) );
  XNOR U44732 ( .A(n43943), .B(n43942), .Z(n44043) );
  NAND U44733 ( .A(x[490]), .B(y[8141]), .Z(n44082) );
  AND U44734 ( .A(x[486]), .B(y[8145]), .Z(n44034) );
  AND U44735 ( .A(x[495]), .B(y[8136]), .Z(n44035) );
  XOR U44736 ( .A(n44034), .B(n44035), .Z(n44036) );
  AND U44737 ( .A(x[491]), .B(y[8140]), .Z(n44037) );
  XOR U44738 ( .A(n44036), .B(n44037), .Z(n44083) );
  XOR U44739 ( .A(n44084), .B(n44083), .Z(n44077) );
  XOR U44740 ( .A(n44078), .B(n44077), .Z(n44147) );
  XOR U44741 ( .A(n44148), .B(n44147), .Z(n44149) );
  XOR U44742 ( .A(n44150), .B(n44149), .Z(n44136) );
  NAND U44743 ( .A(n43945), .B(n43944), .Z(n43949) );
  NAND U44744 ( .A(n43947), .B(n43946), .Z(n43948) );
  NAND U44745 ( .A(n43949), .B(n43948), .Z(n44070) );
  NAND U44746 ( .A(x[498]), .B(y[8138]), .Z(n44830) );
  NANDN U44747 ( .A(n44830), .B(n43950), .Z(n43954) );
  NAND U44748 ( .A(n43952), .B(n43951), .Z(n43953) );
  NAND U44749 ( .A(n43954), .B(n43953), .Z(n44106) );
  NAND U44750 ( .A(n43956), .B(n43955), .Z(n43960) );
  NAND U44751 ( .A(n43958), .B(n43957), .Z(n43959) );
  NAND U44752 ( .A(n43960), .B(n43959), .Z(n44105) );
  XOR U44753 ( .A(n44106), .B(n44105), .Z(n44107) );
  NANDN U44754 ( .A(n44044), .B(n44042), .Z(n43964) );
  NAND U44755 ( .A(n43962), .B(n43961), .Z(n43963) );
  NAND U44756 ( .A(n43964), .B(n43963), .Z(n44119) );
  AND U44757 ( .A(x[480]), .B(y[8151]), .Z(n44053) );
  NAND U44758 ( .A(x[503]), .B(y[8128]), .Z(n44054) );
  AND U44759 ( .A(x[502]), .B(y[8129]), .Z(n44033) );
  XOR U44760 ( .A(o[471]), .B(n44033), .Z(n44055) );
  XOR U44761 ( .A(n44056), .B(n44055), .Z(n44118) );
  NAND U44762 ( .A(y[8131]), .B(x[500]), .Z(n43965) );
  XNOR U44763 ( .A(n43966), .B(n43965), .Z(n44029) );
  AND U44764 ( .A(x[499]), .B(y[8132]), .Z(n44030) );
  XOR U44765 ( .A(n44029), .B(n44030), .Z(n44117) );
  XOR U44766 ( .A(n44118), .B(n44117), .Z(n44120) );
  XOR U44767 ( .A(n44119), .B(n44120), .Z(n44108) );
  XOR U44768 ( .A(n44107), .B(n44108), .Z(n44069) );
  XOR U44769 ( .A(n44070), .B(n44069), .Z(n44072) );
  AND U44770 ( .A(x[500]), .B(y[8137]), .Z(n45014) );
  AND U44771 ( .A(x[493]), .B(y[8130]), .Z(n43967) );
  NAND U44772 ( .A(n45014), .B(n43967), .Z(n43971) );
  NAND U44773 ( .A(n43969), .B(n43968), .Z(n43970) );
  NAND U44774 ( .A(n43971), .B(n43970), .Z(n44064) );
  NAND U44775 ( .A(n43973), .B(n43972), .Z(n43977) );
  NAND U44776 ( .A(n43975), .B(n43974), .Z(n43976) );
  NAND U44777 ( .A(n43977), .B(n43976), .Z(n44125) );
  AND U44778 ( .A(x[493]), .B(y[8138]), .Z(n44099) );
  AND U44779 ( .A(x[482]), .B(y[8149]), .Z(n44100) );
  XOR U44780 ( .A(n44099), .B(n44100), .Z(n44101) );
  AND U44781 ( .A(x[501]), .B(y[8130]), .Z(n44102) );
  XOR U44782 ( .A(n44101), .B(n44102), .Z(n44124) );
  AND U44783 ( .A(x[492]), .B(y[8139]), .Z(n44047) );
  AND U44784 ( .A(x[481]), .B(y[8150]), .Z(n44048) );
  XOR U44785 ( .A(n44047), .B(n44048), .Z(n44050) );
  AND U44786 ( .A(o[470]), .B(n43978), .Z(n44049) );
  XOR U44787 ( .A(n44050), .B(n44049), .Z(n44123) );
  XOR U44788 ( .A(n44124), .B(n44123), .Z(n44126) );
  XOR U44789 ( .A(n44125), .B(n44126), .Z(n44063) );
  XOR U44790 ( .A(n44064), .B(n44063), .Z(n44066) );
  AND U44791 ( .A(x[495]), .B(y[8144]), .Z(n45189) );
  NAND U44792 ( .A(n43979), .B(n45189), .Z(n43983) );
  NAND U44793 ( .A(n43981), .B(n43980), .Z(n43982) );
  NAND U44794 ( .A(n43983), .B(n43982), .Z(n44113) );
  AND U44795 ( .A(x[494]), .B(y[8137]), .Z(n44093) );
  AND U44796 ( .A(x[483]), .B(y[8148]), .Z(n44094) );
  XOR U44797 ( .A(n44093), .B(n44094), .Z(n44095) );
  AND U44798 ( .A(x[484]), .B(y[8147]), .Z(n44096) );
  XOR U44799 ( .A(n44095), .B(n44096), .Z(n44112) );
  AND U44800 ( .A(x[485]), .B(y[8146]), .Z(n44087) );
  AND U44801 ( .A(x[498]), .B(y[8133]), .Z(n44088) );
  XOR U44802 ( .A(n44087), .B(n44088), .Z(n44090) );
  AND U44803 ( .A(x[497]), .B(y[8134]), .Z(n44089) );
  XOR U44804 ( .A(n44090), .B(n44089), .Z(n44111) );
  XOR U44805 ( .A(n44112), .B(n44111), .Z(n44114) );
  XOR U44806 ( .A(n44113), .B(n44114), .Z(n44065) );
  XOR U44807 ( .A(n44066), .B(n44065), .Z(n44071) );
  XOR U44808 ( .A(n44072), .B(n44071), .Z(n44135) );
  XOR U44809 ( .A(n44136), .B(n44135), .Z(n44137) );
  XOR U44810 ( .A(n44138), .B(n44137), .Z(n44025) );
  NAND U44811 ( .A(n43985), .B(n43984), .Z(n43989) );
  NAND U44812 ( .A(n43987), .B(n43986), .Z(n43988) );
  NAND U44813 ( .A(n43989), .B(n43988), .Z(n44144) );
  NAND U44814 ( .A(n43991), .B(n43990), .Z(n43995) );
  NAND U44815 ( .A(n43993), .B(n43992), .Z(n43994) );
  NAND U44816 ( .A(n43995), .B(n43994), .Z(n44142) );
  NAND U44817 ( .A(n43997), .B(n43996), .Z(n44001) );
  NAND U44818 ( .A(n43999), .B(n43998), .Z(n44000) );
  AND U44819 ( .A(n44001), .B(n44000), .Z(n44141) );
  XOR U44820 ( .A(n44142), .B(n44141), .Z(n44143) );
  XOR U44821 ( .A(n44144), .B(n44143), .Z(n44023) );
  NAND U44822 ( .A(n44003), .B(n44002), .Z(n44007) );
  NAND U44823 ( .A(n44005), .B(n44004), .Z(n44006) );
  AND U44824 ( .A(n44007), .B(n44006), .Z(n44022) );
  XOR U44825 ( .A(n44160), .B(n44161), .Z(n44162) );
  XNOR U44826 ( .A(n44163), .B(n44162), .Z(n44156) );
  OR U44827 ( .A(n44010), .B(n44008), .Z(n44014) );
  ANDN U44828 ( .B(n44010), .A(n44009), .Z(n44012) );
  OR U44829 ( .A(n44012), .B(n44011), .Z(n44013) );
  AND U44830 ( .A(n44014), .B(n44013), .Z(n44154) );
  NAND U44831 ( .A(n44016), .B(n44015), .Z(n44020) );
  NAND U44832 ( .A(n44018), .B(n44017), .Z(n44019) );
  AND U44833 ( .A(n44020), .B(n44019), .Z(n44155) );
  IV U44834 ( .A(n44155), .Z(n44153) );
  XOR U44835 ( .A(n44154), .B(n44153), .Z(n44021) );
  XNOR U44836 ( .A(n44156), .B(n44021), .Z(N952) );
  NANDN U44837 ( .A(n44023), .B(n44022), .Z(n44027) );
  NANDN U44838 ( .A(n44025), .B(n44024), .Z(n44026) );
  AND U44839 ( .A(n44027), .B(n44026), .Z(n44302) );
  AND U44840 ( .A(x[500]), .B(y[8135]), .Z(n44028) );
  NAND U44841 ( .A(n44028), .B(n44268), .Z(n44032) );
  NAND U44842 ( .A(n44030), .B(n44029), .Z(n44031) );
  NAND U44843 ( .A(n44032), .B(n44031), .Z(n44288) );
  AND U44844 ( .A(x[502]), .B(y[8130]), .Z(n44195) );
  XOR U44845 ( .A(n44196), .B(n44195), .Z(n44198) );
  NAND U44846 ( .A(x[482]), .B(y[8150]), .Z(n44197) );
  AND U44847 ( .A(x[481]), .B(y[8151]), .Z(n44203) );
  XOR U44848 ( .A(n44204), .B(n44203), .Z(n44202) );
  AND U44849 ( .A(o[471]), .B(n44033), .Z(n44201) );
  XOR U44850 ( .A(n44202), .B(n44201), .Z(n44285) );
  XOR U44851 ( .A(n44286), .B(n44285), .Z(n44287) );
  XOR U44852 ( .A(n44288), .B(n44287), .Z(n44233) );
  NAND U44853 ( .A(n44035), .B(n44034), .Z(n44039) );
  NAND U44854 ( .A(n44037), .B(n44036), .Z(n44038) );
  NAND U44855 ( .A(n44039), .B(n44038), .Z(n44282) );
  AND U44856 ( .A(y[8136]), .B(x[496]), .Z(n44041) );
  NAND U44857 ( .A(y[8131]), .B(x[501]), .Z(n44040) );
  XNOR U44858 ( .A(n44041), .B(n44040), .Z(n44269) );
  AND U44859 ( .A(x[485]), .B(y[8147]), .Z(n44270) );
  XOR U44860 ( .A(n44269), .B(n44270), .Z(n44280) );
  AND U44861 ( .A(x[486]), .B(y[8146]), .Z(n44584) );
  AND U44862 ( .A(x[500]), .B(y[8132]), .Z(n44406) );
  XOR U44863 ( .A(n44584), .B(n44406), .Z(n44275) );
  AND U44864 ( .A(x[499]), .B(y[8133]), .Z(n44276) );
  XOR U44865 ( .A(n44275), .B(n44276), .Z(n44279) );
  XOR U44866 ( .A(n44280), .B(n44279), .Z(n44281) );
  XOR U44867 ( .A(n44282), .B(n44281), .Z(n44259) );
  NANDN U44868 ( .A(n44332), .B(n44042), .Z(n44046) );
  NANDN U44869 ( .A(n44044), .B(n44043), .Z(n44045) );
  NAND U44870 ( .A(n44046), .B(n44045), .Z(n44257) );
  NAND U44871 ( .A(n44048), .B(n44047), .Z(n44052) );
  NAND U44872 ( .A(n44050), .B(n44049), .Z(n44051) );
  NAND U44873 ( .A(n44052), .B(n44051), .Z(n44256) );
  XOR U44874 ( .A(n44257), .B(n44256), .Z(n44258) );
  XOR U44875 ( .A(n44259), .B(n44258), .Z(n44232) );
  XOR U44876 ( .A(n44233), .B(n44232), .Z(n44235) );
  NANDN U44877 ( .A(n44054), .B(n44053), .Z(n44058) );
  NAND U44878 ( .A(n44056), .B(n44055), .Z(n44057) );
  AND U44879 ( .A(n44058), .B(n44057), .Z(n44227) );
  AND U44880 ( .A(x[483]), .B(y[8149]), .Z(n44216) );
  XOR U44881 ( .A(n44217), .B(n44216), .Z(n44215) );
  AND U44882 ( .A(x[484]), .B(y[8148]), .Z(n44214) );
  XOR U44883 ( .A(n44215), .B(n44214), .Z(n44226) );
  AND U44884 ( .A(y[8143]), .B(x[489]), .Z(n44060) );
  NAND U44885 ( .A(y[8142]), .B(x[490]), .Z(n44059) );
  XNOR U44886 ( .A(n44060), .B(n44059), .Z(n44187) );
  AND U44887 ( .A(y[8138]), .B(x[494]), .Z(n44062) );
  NAND U44888 ( .A(y[8144]), .B(x[488]), .Z(n44061) );
  XNOR U44889 ( .A(n44062), .B(n44061), .Z(n44191) );
  AND U44890 ( .A(x[491]), .B(y[8141]), .Z(n44192) );
  XOR U44891 ( .A(n44191), .B(n44192), .Z(n44186) );
  XOR U44892 ( .A(n44187), .B(n44186), .Z(n44228) );
  XOR U44893 ( .A(n44229), .B(n44228), .Z(n44234) );
  XNOR U44894 ( .A(n44235), .B(n44234), .Z(n44180) );
  NAND U44895 ( .A(n44064), .B(n44063), .Z(n44068) );
  NAND U44896 ( .A(n44066), .B(n44065), .Z(n44067) );
  AND U44897 ( .A(n44068), .B(n44067), .Z(n44179) );
  XOR U44898 ( .A(n44180), .B(n44179), .Z(n44181) );
  NAND U44899 ( .A(n44070), .B(n44069), .Z(n44074) );
  NAND U44900 ( .A(n44072), .B(n44071), .Z(n44073) );
  AND U44901 ( .A(n44074), .B(n44073), .Z(n44182) );
  XOR U44902 ( .A(n44181), .B(n44182), .Z(n44176) );
  NAND U44903 ( .A(n44076), .B(n44075), .Z(n44080) );
  NAND U44904 ( .A(n44078), .B(n44077), .Z(n44079) );
  AND U44905 ( .A(n44080), .B(n44079), .Z(n44241) );
  NANDN U44906 ( .A(n44082), .B(n44081), .Z(n44086) );
  NAND U44907 ( .A(n44084), .B(n44083), .Z(n44085) );
  AND U44908 ( .A(n44086), .B(n44085), .Z(n44239) );
  NAND U44909 ( .A(n44088), .B(n44087), .Z(n44092) );
  NAND U44910 ( .A(n44090), .B(n44089), .Z(n44091) );
  NAND U44911 ( .A(n44092), .B(n44091), .Z(n44265) );
  AND U44912 ( .A(x[480]), .B(y[8152]), .Z(n44220) );
  AND U44913 ( .A(x[504]), .B(y[8128]), .Z(n44221) );
  XOR U44914 ( .A(n44220), .B(n44221), .Z(n44223) );
  AND U44915 ( .A(x[503]), .B(y[8129]), .Z(n44213) );
  XOR U44916 ( .A(o[472]), .B(n44213), .Z(n44222) );
  XOR U44917 ( .A(n44223), .B(n44222), .Z(n44263) );
  AND U44918 ( .A(x[487]), .B(y[8145]), .Z(n44207) );
  NAND U44919 ( .A(x[498]), .B(y[8134]), .Z(n44208) );
  NAND U44920 ( .A(x[497]), .B(y[8135]), .Z(n44210) );
  XOR U44921 ( .A(n44263), .B(n44262), .Z(n44264) );
  XOR U44922 ( .A(n44265), .B(n44264), .Z(n44253) );
  NAND U44923 ( .A(n44094), .B(n44093), .Z(n44098) );
  NAND U44924 ( .A(n44096), .B(n44095), .Z(n44097) );
  NAND U44925 ( .A(n44098), .B(n44097), .Z(n44251) );
  NAND U44926 ( .A(n44100), .B(n44099), .Z(n44104) );
  NAND U44927 ( .A(n44102), .B(n44101), .Z(n44103) );
  NAND U44928 ( .A(n44104), .B(n44103), .Z(n44250) );
  XOR U44929 ( .A(n44251), .B(n44250), .Z(n44252) );
  XOR U44930 ( .A(n44253), .B(n44252), .Z(n44238) );
  NAND U44931 ( .A(n44106), .B(n44105), .Z(n44110) );
  NAND U44932 ( .A(n44108), .B(n44107), .Z(n44109) );
  AND U44933 ( .A(n44110), .B(n44109), .Z(n44294) );
  NAND U44934 ( .A(n44112), .B(n44111), .Z(n44116) );
  NAND U44935 ( .A(n44114), .B(n44113), .Z(n44115) );
  AND U44936 ( .A(n44116), .B(n44115), .Z(n44292) );
  NAND U44937 ( .A(n44118), .B(n44117), .Z(n44122) );
  NAND U44938 ( .A(n44120), .B(n44119), .Z(n44121) );
  AND U44939 ( .A(n44122), .B(n44121), .Z(n44291) );
  XOR U44940 ( .A(n44292), .B(n44291), .Z(n44293) );
  XOR U44941 ( .A(n44294), .B(n44293), .Z(n44244) );
  NAND U44942 ( .A(n44124), .B(n44123), .Z(n44128) );
  NAND U44943 ( .A(n44126), .B(n44125), .Z(n44127) );
  AND U44944 ( .A(n44128), .B(n44127), .Z(n44245) );
  XOR U44945 ( .A(n44244), .B(n44245), .Z(n44247) );
  XOR U44946 ( .A(n44246), .B(n44247), .Z(n44173) );
  NAND U44947 ( .A(n44130), .B(n44129), .Z(n44134) );
  NAND U44948 ( .A(n44132), .B(n44131), .Z(n44133) );
  AND U44949 ( .A(n44134), .B(n44133), .Z(n44174) );
  XOR U44950 ( .A(n44173), .B(n44174), .Z(n44175) );
  XNOR U44951 ( .A(n44176), .B(n44175), .Z(n44300) );
  NAND U44952 ( .A(n44136), .B(n44135), .Z(n44140) );
  NAND U44953 ( .A(n44138), .B(n44137), .Z(n44139) );
  NAND U44954 ( .A(n44140), .B(n44139), .Z(n44170) );
  NAND U44955 ( .A(n44142), .B(n44141), .Z(n44146) );
  NAND U44956 ( .A(n44144), .B(n44143), .Z(n44145) );
  NAND U44957 ( .A(n44146), .B(n44145), .Z(n44168) );
  NAND U44958 ( .A(n44148), .B(n44147), .Z(n44152) );
  NAND U44959 ( .A(n44150), .B(n44149), .Z(n44151) );
  NAND U44960 ( .A(n44152), .B(n44151), .Z(n44167) );
  XOR U44961 ( .A(n44168), .B(n44167), .Z(n44169) );
  XNOR U44962 ( .A(n44170), .B(n44169), .Z(n44301) );
  XOR U44963 ( .A(n44300), .B(n44301), .Z(n44303) );
  XNOR U44964 ( .A(n44302), .B(n44303), .Z(n44299) );
  NANDN U44965 ( .A(n44153), .B(n44154), .Z(n44159) );
  NOR U44966 ( .A(n44155), .B(n44154), .Z(n44157) );
  OR U44967 ( .A(n44157), .B(n44156), .Z(n44158) );
  AND U44968 ( .A(n44159), .B(n44158), .Z(n44298) );
  NAND U44969 ( .A(n44161), .B(n44160), .Z(n44165) );
  NAND U44970 ( .A(n44163), .B(n44162), .Z(n44164) );
  NAND U44971 ( .A(n44165), .B(n44164), .Z(n44297) );
  XOR U44972 ( .A(n44298), .B(n44297), .Z(n44166) );
  XNOR U44973 ( .A(n44299), .B(n44166), .Z(N953) );
  NAND U44974 ( .A(n44168), .B(n44167), .Z(n44172) );
  NAND U44975 ( .A(n44170), .B(n44169), .Z(n44171) );
  AND U44976 ( .A(n44172), .B(n44171), .Z(n44453) );
  NAND U44977 ( .A(n44174), .B(n44173), .Z(n44178) );
  NAND U44978 ( .A(n44176), .B(n44175), .Z(n44177) );
  NAND U44979 ( .A(n44178), .B(n44177), .Z(n44451) );
  NAND U44980 ( .A(n44180), .B(n44179), .Z(n44184) );
  NAND U44981 ( .A(n44182), .B(n44181), .Z(n44183) );
  NAND U44982 ( .A(n44184), .B(n44183), .Z(n44308) );
  NANDN U44983 ( .A(n44331), .B(n44185), .Z(n44189) );
  NAND U44984 ( .A(n44187), .B(n44186), .Z(n44188) );
  NAND U44985 ( .A(n44189), .B(n44188), .Z(n44356) );
  AND U44986 ( .A(x[494]), .B(y[8144]), .Z(n45286) );
  NAND U44987 ( .A(n45286), .B(n44190), .Z(n44194) );
  NAND U44988 ( .A(n44192), .B(n44191), .Z(n44193) );
  NAND U44989 ( .A(n44194), .B(n44193), .Z(n44383) );
  NAND U44990 ( .A(x[491]), .B(y[8142]), .Z(n44402) );
  NAND U44991 ( .A(x[492]), .B(y[8141]), .Z(n44401) );
  NAND U44992 ( .A(x[487]), .B(y[8146]), .Z(n44400) );
  XOR U44993 ( .A(n44401), .B(n44400), .Z(n44403) );
  XNOR U44994 ( .A(n44402), .B(n44403), .Z(n44382) );
  NAND U44995 ( .A(x[504]), .B(y[8129]), .Z(n44399) );
  XNOR U44996 ( .A(o[473]), .B(n44399), .Z(n44370) );
  AND U44997 ( .A(x[481]), .B(y[8152]), .Z(n44369) );
  XOR U44998 ( .A(n44370), .B(n44369), .Z(n44372) );
  AND U44999 ( .A(x[493]), .B(y[8140]), .Z(n44371) );
  XOR U45000 ( .A(n44372), .B(n44371), .Z(n44381) );
  XOR U45001 ( .A(n44382), .B(n44381), .Z(n44384) );
  XOR U45002 ( .A(n44383), .B(n44384), .Z(n44355) );
  XOR U45003 ( .A(n44356), .B(n44355), .Z(n44358) );
  NAND U45004 ( .A(n44196), .B(n44195), .Z(n44200) );
  ANDN U45005 ( .B(n44198), .A(n44197), .Z(n44199) );
  ANDN U45006 ( .B(n44200), .A(n44199), .Z(n44344) );
  AND U45007 ( .A(n44202), .B(n44201), .Z(n44206) );
  NAND U45008 ( .A(n44204), .B(n44203), .Z(n44205) );
  NANDN U45009 ( .A(n44206), .B(n44205), .Z(n44343) );
  NANDN U45010 ( .A(n44208), .B(n44207), .Z(n44212) );
  NANDN U45011 ( .A(n44210), .B(n44209), .Z(n44211) );
  AND U45012 ( .A(n44212), .B(n44211), .Z(n44340) );
  NAND U45013 ( .A(x[488]), .B(y[8145]), .Z(n44333) );
  XOR U45014 ( .A(n44332), .B(n44331), .Z(n44334) );
  XNOR U45015 ( .A(n44333), .B(n44334), .Z(n44338) );
  NAND U45016 ( .A(n44213), .B(o[472]), .Z(n44327) );
  NAND U45017 ( .A(x[505]), .B(y[8128]), .Z(n44326) );
  NAND U45018 ( .A(x[480]), .B(y[8153]), .Z(n44325) );
  XNOR U45019 ( .A(n44326), .B(n44325), .Z(n44328) );
  XOR U45020 ( .A(n44327), .B(n44328), .Z(n44337) );
  XOR U45021 ( .A(n44338), .B(n44337), .Z(n44339) );
  XOR U45022 ( .A(n44346), .B(n44345), .Z(n44357) );
  XOR U45023 ( .A(n44358), .B(n44357), .Z(n44444) );
  AND U45024 ( .A(n44215), .B(n44214), .Z(n44219) );
  NAND U45025 ( .A(n44217), .B(n44216), .Z(n44218) );
  NANDN U45026 ( .A(n44219), .B(n44218), .Z(n44420) );
  NAND U45027 ( .A(n44221), .B(n44220), .Z(n44225) );
  NAND U45028 ( .A(n44223), .B(n44222), .Z(n44224) );
  NAND U45029 ( .A(n44225), .B(n44224), .Z(n44418) );
  AND U45030 ( .A(x[494]), .B(y[8139]), .Z(n44376) );
  AND U45031 ( .A(x[482]), .B(y[8151]), .Z(n44375) );
  XOR U45032 ( .A(n44376), .B(n44375), .Z(n44378) );
  AND U45033 ( .A(x[483]), .B(y[8150]), .Z(n44377) );
  XOR U45034 ( .A(n44378), .B(n44377), .Z(n44417) );
  XOR U45035 ( .A(n44418), .B(n44417), .Z(n44419) );
  XOR U45036 ( .A(n44420), .B(n44419), .Z(n44442) );
  NANDN U45037 ( .A(n44227), .B(n44226), .Z(n44231) );
  NAND U45038 ( .A(n44229), .B(n44228), .Z(n44230) );
  AND U45039 ( .A(n44231), .B(n44230), .Z(n44441) );
  NAND U45040 ( .A(n44233), .B(n44232), .Z(n44237) );
  NAND U45041 ( .A(n44235), .B(n44234), .Z(n44236) );
  NAND U45042 ( .A(n44237), .B(n44236), .Z(n44436) );
  NANDN U45043 ( .A(n44239), .B(n44238), .Z(n44243) );
  NANDN U45044 ( .A(n44241), .B(n44240), .Z(n44242) );
  NAND U45045 ( .A(n44243), .B(n44242), .Z(n44438) );
  XOR U45046 ( .A(n44308), .B(n44307), .Z(n44310) );
  NAND U45047 ( .A(n44245), .B(n44244), .Z(n44249) );
  NAND U45048 ( .A(n44247), .B(n44246), .Z(n44248) );
  NAND U45049 ( .A(n44249), .B(n44248), .Z(n44315) );
  NAND U45050 ( .A(n44251), .B(n44250), .Z(n44255) );
  NAND U45051 ( .A(n44253), .B(n44252), .Z(n44254) );
  AND U45052 ( .A(n44255), .B(n44254), .Z(n44320) );
  NAND U45053 ( .A(n44257), .B(n44256), .Z(n44261) );
  NAND U45054 ( .A(n44259), .B(n44258), .Z(n44260) );
  NAND U45055 ( .A(n44261), .B(n44260), .Z(n44319) );
  NAND U45056 ( .A(n44263), .B(n44262), .Z(n44267) );
  NAND U45057 ( .A(n44265), .B(n44264), .Z(n44266) );
  AND U45058 ( .A(n44267), .B(n44266), .Z(n44352) );
  AND U45059 ( .A(x[501]), .B(y[8136]), .Z(n45169) );
  NAND U45060 ( .A(n45169), .B(n44268), .Z(n44272) );
  NAND U45061 ( .A(n44270), .B(n44269), .Z(n44271) );
  NAND U45062 ( .A(n44272), .B(n44271), .Z(n44426) );
  NAND U45063 ( .A(x[502]), .B(y[8131]), .Z(n44395) );
  NAND U45064 ( .A(x[485]), .B(y[8148]), .Z(n44394) );
  NAND U45065 ( .A(x[497]), .B(y[8136]), .Z(n44393) );
  XOR U45066 ( .A(n44394), .B(n44393), .Z(n44396) );
  XNOR U45067 ( .A(n44395), .B(n44396), .Z(n44423) );
  AND U45068 ( .A(y[8133]), .B(x[500]), .Z(n44274) );
  NAND U45069 ( .A(y[8132]), .B(x[501]), .Z(n44273) );
  XNOR U45070 ( .A(n44274), .B(n44273), .Z(n44408) );
  AND U45071 ( .A(x[499]), .B(y[8134]), .Z(n44407) );
  XOR U45072 ( .A(n44408), .B(n44407), .Z(n44424) );
  XOR U45073 ( .A(n44423), .B(n44424), .Z(n44425) );
  XNOR U45074 ( .A(n44426), .B(n44425), .Z(n44350) );
  NAND U45075 ( .A(n44406), .B(n44584), .Z(n44278) );
  NAND U45076 ( .A(n44276), .B(n44275), .Z(n44277) );
  AND U45077 ( .A(n44278), .B(n44277), .Z(n44432) );
  NAND U45078 ( .A(x[495]), .B(y[8138]), .Z(n44413) );
  NAND U45079 ( .A(x[498]), .B(y[8135]), .Z(n44412) );
  NAND U45080 ( .A(x[486]), .B(y[8147]), .Z(n44411) );
  XOR U45081 ( .A(n44412), .B(n44411), .Z(n44414) );
  XNOR U45082 ( .A(n44413), .B(n44414), .Z(n44430) );
  NAND U45083 ( .A(x[503]), .B(y[8130]), .Z(n44389) );
  NAND U45084 ( .A(x[484]), .B(y[8149]), .Z(n44388) );
  NAND U45085 ( .A(x[496]), .B(y[8137]), .Z(n44387) );
  XNOR U45086 ( .A(n44388), .B(n44387), .Z(n44390) );
  XOR U45087 ( .A(n44389), .B(n44390), .Z(n44429) );
  XOR U45088 ( .A(n44430), .B(n44429), .Z(n44431) );
  XOR U45089 ( .A(n44432), .B(n44431), .Z(n44349) );
  XOR U45090 ( .A(n44350), .B(n44349), .Z(n44351) );
  XNOR U45091 ( .A(n44352), .B(n44351), .Z(n44364) );
  NAND U45092 ( .A(n44280), .B(n44279), .Z(n44284) );
  NAND U45093 ( .A(n44282), .B(n44281), .Z(n44283) );
  NAND U45094 ( .A(n44284), .B(n44283), .Z(n44362) );
  NAND U45095 ( .A(n44286), .B(n44285), .Z(n44290) );
  NAND U45096 ( .A(n44288), .B(n44287), .Z(n44289) );
  NAND U45097 ( .A(n44290), .B(n44289), .Z(n44361) );
  XOR U45098 ( .A(n44362), .B(n44361), .Z(n44363) );
  XOR U45099 ( .A(n44364), .B(n44363), .Z(n44321) );
  XNOR U45100 ( .A(n44322), .B(n44321), .Z(n44314) );
  NAND U45101 ( .A(n44292), .B(n44291), .Z(n44296) );
  NAND U45102 ( .A(n44294), .B(n44293), .Z(n44295) );
  NAND U45103 ( .A(n44296), .B(n44295), .Z(n44313) );
  XOR U45104 ( .A(n44314), .B(n44313), .Z(n44316) );
  XOR U45105 ( .A(n44315), .B(n44316), .Z(n44309) );
  XOR U45106 ( .A(n44310), .B(n44309), .Z(n44450) );
  XOR U45107 ( .A(n44451), .B(n44450), .Z(n44452) );
  XNOR U45108 ( .A(n44453), .B(n44452), .Z(n44449) );
  NANDN U45109 ( .A(n44301), .B(n44300), .Z(n44305) );
  NANDN U45110 ( .A(n44303), .B(n44302), .Z(n44304) );
  AND U45111 ( .A(n44305), .B(n44304), .Z(n44447) );
  XOR U45112 ( .A(n44448), .B(n44447), .Z(n44306) );
  XNOR U45113 ( .A(n44449), .B(n44306), .Z(N954) );
  NAND U45114 ( .A(n44308), .B(n44307), .Z(n44312) );
  NAND U45115 ( .A(n44310), .B(n44309), .Z(n44311) );
  AND U45116 ( .A(n44312), .B(n44311), .Z(n44607) );
  NAND U45117 ( .A(n44314), .B(n44313), .Z(n44318) );
  NAND U45118 ( .A(n44316), .B(n44315), .Z(n44317) );
  AND U45119 ( .A(n44318), .B(n44317), .Z(n44608) );
  XOR U45120 ( .A(n44607), .B(n44608), .Z(n44610) );
  NANDN U45121 ( .A(n44320), .B(n44319), .Z(n44324) );
  NAND U45122 ( .A(n44322), .B(n44321), .Z(n44323) );
  AND U45123 ( .A(n44324), .B(n44323), .Z(n44466) );
  AND U45124 ( .A(x[482]), .B(y[8152]), .Z(n44487) );
  XOR U45125 ( .A(n44488), .B(n44487), .Z(n44490) );
  NAND U45126 ( .A(x[504]), .B(y[8130]), .Z(n44489) );
  XNOR U45127 ( .A(n44490), .B(n44489), .Z(n44530) );
  NAND U45128 ( .A(n44326), .B(n44325), .Z(n44330) );
  NANDN U45129 ( .A(n44328), .B(n44327), .Z(n44329) );
  AND U45130 ( .A(n44330), .B(n44329), .Z(n44529) );
  XOR U45131 ( .A(n44530), .B(n44529), .Z(n44532) );
  NAND U45132 ( .A(n44332), .B(n44331), .Z(n44336) );
  NAND U45133 ( .A(n44334), .B(n44333), .Z(n44335) );
  AND U45134 ( .A(n44336), .B(n44335), .Z(n44531) );
  XOR U45135 ( .A(n44532), .B(n44531), .Z(n44561) );
  NAND U45136 ( .A(n44338), .B(n44337), .Z(n44342) );
  NANDN U45137 ( .A(n44340), .B(n44339), .Z(n44341) );
  AND U45138 ( .A(n44342), .B(n44341), .Z(n44560) );
  NANDN U45139 ( .A(n44344), .B(n44343), .Z(n44348) );
  NAND U45140 ( .A(n44346), .B(n44345), .Z(n44347) );
  NAND U45141 ( .A(n44348), .B(n44347), .Z(n44563) );
  NAND U45142 ( .A(n44350), .B(n44349), .Z(n44354) );
  NAND U45143 ( .A(n44352), .B(n44351), .Z(n44353) );
  NAND U45144 ( .A(n44354), .B(n44353), .Z(n44555) );
  NAND U45145 ( .A(n44356), .B(n44355), .Z(n44360) );
  NAND U45146 ( .A(n44358), .B(n44357), .Z(n44359) );
  AND U45147 ( .A(n44360), .B(n44359), .Z(n44554) );
  XOR U45148 ( .A(n44555), .B(n44554), .Z(n44556) );
  XOR U45149 ( .A(n44557), .B(n44556), .Z(n44464) );
  NAND U45150 ( .A(n44362), .B(n44361), .Z(n44366) );
  NAND U45151 ( .A(n44364), .B(n44363), .Z(n44365) );
  NAND U45152 ( .A(n44366), .B(n44365), .Z(n44472) );
  AND U45153 ( .A(x[492]), .B(y[8142]), .Z(n44720) );
  AND U45154 ( .A(x[485]), .B(y[8149]), .Z(n44543) );
  XOR U45155 ( .A(n44720), .B(n44543), .Z(n44545) );
  NAND U45156 ( .A(x[490]), .B(y[8144]), .Z(n44544) );
  XNOR U45157 ( .A(n44545), .B(n44544), .Z(n44569) );
  AND U45158 ( .A(x[487]), .B(y[8147]), .Z(n44566) );
  AND U45159 ( .A(y[8148]), .B(x[486]), .Z(n44368) );
  NAND U45160 ( .A(y[8146]), .B(x[488]), .Z(n44367) );
  XNOR U45161 ( .A(n44368), .B(n44367), .Z(n44585) );
  NAND U45162 ( .A(x[489]), .B(y[8145]), .Z(n44586) );
  XOR U45163 ( .A(n44585), .B(n44586), .Z(n44567) );
  XOR U45164 ( .A(n44569), .B(n44568), .Z(n44513) );
  NAND U45165 ( .A(n44370), .B(n44369), .Z(n44374) );
  NAND U45166 ( .A(n44372), .B(n44371), .Z(n44373) );
  NAND U45167 ( .A(n44374), .B(n44373), .Z(n44512) );
  NAND U45168 ( .A(n44376), .B(n44375), .Z(n44380) );
  NAND U45169 ( .A(n44378), .B(n44377), .Z(n44379) );
  NAND U45170 ( .A(n44380), .B(n44379), .Z(n44511) );
  XOR U45171 ( .A(n44512), .B(n44511), .Z(n44514) );
  XNOR U45172 ( .A(n44513), .B(n44514), .Z(n44518) );
  NAND U45173 ( .A(n44382), .B(n44381), .Z(n44386) );
  NAND U45174 ( .A(n44384), .B(n44383), .Z(n44385) );
  AND U45175 ( .A(n44386), .B(n44385), .Z(n44517) );
  XOR U45176 ( .A(n44518), .B(n44517), .Z(n44520) );
  NAND U45177 ( .A(n44388), .B(n44387), .Z(n44392) );
  NANDN U45178 ( .A(n44390), .B(n44389), .Z(n44391) );
  AND U45179 ( .A(n44392), .B(n44391), .Z(n44476) );
  NAND U45180 ( .A(n44394), .B(n44393), .Z(n44398) );
  NAND U45181 ( .A(n44396), .B(n44395), .Z(n44397) );
  AND U45182 ( .A(n44398), .B(n44397), .Z(n44475) );
  XOR U45183 ( .A(n44476), .B(n44475), .Z(n44478) );
  ANDN U45184 ( .B(o[473]), .A(n44399), .Z(n44578) );
  NAND U45185 ( .A(x[494]), .B(y[8140]), .Z(n44579) );
  XNOR U45186 ( .A(n44578), .B(n44579), .Z(n44580) );
  NAND U45187 ( .A(x[481]), .B(y[8153]), .Z(n44581) );
  XNOR U45188 ( .A(n44580), .B(n44581), .Z(n44536) );
  NAND U45189 ( .A(x[505]), .B(y[8129]), .Z(n44589) );
  XNOR U45190 ( .A(o[474]), .B(n44589), .Z(n44548) );
  NAND U45191 ( .A(x[506]), .B(y[8128]), .Z(n44549) );
  XNOR U45192 ( .A(n44548), .B(n44549), .Z(n44551) );
  AND U45193 ( .A(x[480]), .B(y[8154]), .Z(n44550) );
  XOR U45194 ( .A(n44551), .B(n44550), .Z(n44535) );
  XOR U45195 ( .A(n44536), .B(n44535), .Z(n44538) );
  NAND U45196 ( .A(n44401), .B(n44400), .Z(n44405) );
  NAND U45197 ( .A(n44403), .B(n44402), .Z(n44404) );
  AND U45198 ( .A(n44405), .B(n44404), .Z(n44537) );
  XOR U45199 ( .A(n44538), .B(n44537), .Z(n44477) );
  XOR U45200 ( .A(n44478), .B(n44477), .Z(n44526) );
  AND U45201 ( .A(x[501]), .B(y[8133]), .Z(n44572) );
  NAND U45202 ( .A(n44406), .B(n44572), .Z(n44410) );
  NAND U45203 ( .A(n44408), .B(n44407), .Z(n44409) );
  NAND U45204 ( .A(n44410), .B(n44409), .Z(n44507) );
  XOR U45205 ( .A(n44573), .B(n44572), .Z(n44575) );
  NAND U45206 ( .A(x[500]), .B(y[8134]), .Z(n44574) );
  XNOR U45207 ( .A(n44575), .B(n44574), .Z(n44506) );
  NAND U45208 ( .A(x[503]), .B(y[8131]), .Z(n44494) );
  XNOR U45209 ( .A(n44493), .B(n44494), .Z(n44496) );
  AND U45210 ( .A(x[502]), .B(y[8132]), .Z(n44495) );
  XOR U45211 ( .A(n44496), .B(n44495), .Z(n44505) );
  XOR U45212 ( .A(n44506), .B(n44505), .Z(n44508) );
  XOR U45213 ( .A(n44507), .B(n44508), .Z(n44524) );
  AND U45214 ( .A(x[499]), .B(y[8135]), .Z(n44590) );
  NAND U45215 ( .A(x[491]), .B(y[8143]), .Z(n44591) );
  XNOR U45216 ( .A(n44590), .B(n44591), .Z(n44592) );
  NAND U45217 ( .A(x[483]), .B(y[8151]), .Z(n44593) );
  XNOR U45218 ( .A(n44592), .B(n44593), .Z(n44482) );
  AND U45219 ( .A(x[484]), .B(y[8150]), .Z(n44499) );
  XOR U45220 ( .A(n44500), .B(n44499), .Z(n44502) );
  XOR U45221 ( .A(n44502), .B(n44501), .Z(n44481) );
  XOR U45222 ( .A(n44482), .B(n44481), .Z(n44484) );
  NAND U45223 ( .A(n44412), .B(n44411), .Z(n44416) );
  NAND U45224 ( .A(n44414), .B(n44413), .Z(n44415) );
  AND U45225 ( .A(n44416), .B(n44415), .Z(n44483) );
  XNOR U45226 ( .A(n44484), .B(n44483), .Z(n44523) );
  XNOR U45227 ( .A(n44520), .B(n44519), .Z(n44470) );
  NAND U45228 ( .A(n44418), .B(n44417), .Z(n44422) );
  NAND U45229 ( .A(n44420), .B(n44419), .Z(n44421) );
  AND U45230 ( .A(n44422), .B(n44421), .Z(n44601) );
  NAND U45231 ( .A(n44424), .B(n44423), .Z(n44428) );
  NAND U45232 ( .A(n44426), .B(n44425), .Z(n44427) );
  AND U45233 ( .A(n44428), .B(n44427), .Z(n44599) );
  NAND U45234 ( .A(n44430), .B(n44429), .Z(n44434) );
  NANDN U45235 ( .A(n44432), .B(n44431), .Z(n44433) );
  NAND U45236 ( .A(n44434), .B(n44433), .Z(n44598) );
  XOR U45237 ( .A(n44470), .B(n44469), .Z(n44471) );
  XOR U45238 ( .A(n44472), .B(n44471), .Z(n44463) );
  NANDN U45239 ( .A(n44436), .B(n44435), .Z(n44440) );
  NANDN U45240 ( .A(n44438), .B(n44437), .Z(n44439) );
  AND U45241 ( .A(n44440), .B(n44439), .Z(n44457) );
  NANDN U45242 ( .A(n44442), .B(n44441), .Z(n44446) );
  NANDN U45243 ( .A(n44444), .B(n44443), .Z(n44445) );
  NAND U45244 ( .A(n44446), .B(n44445), .Z(n44458) );
  XOR U45245 ( .A(n44460), .B(n44459), .Z(n44609) );
  XNOR U45246 ( .A(n44610), .B(n44609), .Z(n44606) );
  NAND U45247 ( .A(n44451), .B(n44450), .Z(n44455) );
  NAND U45248 ( .A(n44453), .B(n44452), .Z(n44454) );
  AND U45249 ( .A(n44455), .B(n44454), .Z(n44605) );
  XOR U45250 ( .A(n44604), .B(n44605), .Z(n44456) );
  XNOR U45251 ( .A(n44606), .B(n44456), .Z(N955) );
  NANDN U45252 ( .A(n44458), .B(n44457), .Z(n44462) );
  NAND U45253 ( .A(n44460), .B(n44459), .Z(n44461) );
  AND U45254 ( .A(n44462), .B(n44461), .Z(n44758) );
  NANDN U45255 ( .A(n44464), .B(n44463), .Z(n44468) );
  NANDN U45256 ( .A(n44466), .B(n44465), .Z(n44467) );
  AND U45257 ( .A(n44468), .B(n44467), .Z(n44756) );
  NAND U45258 ( .A(n44470), .B(n44469), .Z(n44474) );
  NAND U45259 ( .A(n44472), .B(n44471), .Z(n44473) );
  NAND U45260 ( .A(n44474), .B(n44473), .Z(n44616) );
  NAND U45261 ( .A(n44476), .B(n44475), .Z(n44480) );
  NAND U45262 ( .A(n44478), .B(n44477), .Z(n44479) );
  NAND U45263 ( .A(n44480), .B(n44479), .Z(n44640) );
  NAND U45264 ( .A(n44482), .B(n44481), .Z(n44486) );
  NAND U45265 ( .A(n44484), .B(n44483), .Z(n44485) );
  NAND U45266 ( .A(n44486), .B(n44485), .Z(n44638) );
  NAND U45267 ( .A(n44488), .B(n44487), .Z(n44492) );
  ANDN U45268 ( .B(n44490), .A(n44489), .Z(n44491) );
  ANDN U45269 ( .B(n44492), .A(n44491), .Z(n44693) );
  NANDN U45270 ( .A(n44494), .B(n44493), .Z(n44498) );
  NAND U45271 ( .A(n44496), .B(n44495), .Z(n44497) );
  NAND U45272 ( .A(n44498), .B(n44497), .Z(n44692) );
  XNOR U45273 ( .A(n44693), .B(n44692), .Z(n44694) );
  NAND U45274 ( .A(n44500), .B(n44499), .Z(n44504) );
  AND U45275 ( .A(n44502), .B(n44501), .Z(n44503) );
  ANDN U45276 ( .B(n44504), .A(n44503), .Z(n44707) );
  AND U45277 ( .A(x[480]), .B(y[8155]), .Z(n44661) );
  NAND U45278 ( .A(x[507]), .B(y[8128]), .Z(n44662) );
  XNOR U45279 ( .A(n44661), .B(n44662), .Z(n44664) );
  NAND U45280 ( .A(x[506]), .B(y[8129]), .Z(n44671) );
  XOR U45281 ( .A(n44664), .B(n44663), .Z(n44704) );
  AND U45282 ( .A(x[489]), .B(y[8146]), .Z(n44665) );
  NAND U45283 ( .A(x[501]), .B(y[8134]), .Z(n44666) );
  XNOR U45284 ( .A(n44665), .B(n44666), .Z(n44667) );
  NAND U45285 ( .A(x[498]), .B(y[8137]), .Z(n44668) );
  XOR U45286 ( .A(n44667), .B(n44668), .Z(n44705) );
  XNOR U45287 ( .A(n44704), .B(n44705), .Z(n44706) );
  XOR U45288 ( .A(n44707), .B(n44706), .Z(n44695) );
  XNOR U45289 ( .A(n44694), .B(n44695), .Z(n44639) );
  XOR U45290 ( .A(n44638), .B(n44639), .Z(n44641) );
  XOR U45291 ( .A(n44640), .B(n44641), .Z(n44752) );
  NAND U45292 ( .A(n44506), .B(n44505), .Z(n44510) );
  NAND U45293 ( .A(n44508), .B(n44507), .Z(n44509) );
  AND U45294 ( .A(n44510), .B(n44509), .Z(n44750) );
  NAND U45295 ( .A(n44512), .B(n44511), .Z(n44516) );
  NAND U45296 ( .A(n44514), .B(n44513), .Z(n44515) );
  AND U45297 ( .A(n44516), .B(n44515), .Z(n44749) );
  XOR U45298 ( .A(n44750), .B(n44749), .Z(n44751) );
  NAND U45299 ( .A(n44518), .B(n44517), .Z(n44522) );
  NAND U45300 ( .A(n44520), .B(n44519), .Z(n44521) );
  AND U45301 ( .A(n44522), .B(n44521), .Z(n44740) );
  NANDN U45302 ( .A(n44524), .B(n44523), .Z(n44528) );
  NANDN U45303 ( .A(n44526), .B(n44525), .Z(n44527) );
  AND U45304 ( .A(n44528), .B(n44527), .Z(n44737) );
  NAND U45305 ( .A(n44530), .B(n44529), .Z(n44534) );
  NAND U45306 ( .A(n44532), .B(n44531), .Z(n44533) );
  NAND U45307 ( .A(n44534), .B(n44533), .Z(n44634) );
  NAND U45308 ( .A(n44536), .B(n44535), .Z(n44540) );
  NAND U45309 ( .A(n44538), .B(n44537), .Z(n44539) );
  NAND U45310 ( .A(n44540), .B(n44539), .Z(n44632) );
  AND U45311 ( .A(x[499]), .B(y[8136]), .Z(n44649) );
  NAND U45312 ( .A(x[505]), .B(y[8130]), .Z(n44650) );
  XNOR U45313 ( .A(n44649), .B(n44650), .Z(n44651) );
  NAND U45314 ( .A(x[486]), .B(y[8149]), .Z(n44652) );
  XNOR U45315 ( .A(n44651), .B(n44652), .Z(n44683) );
  AND U45316 ( .A(x[495]), .B(y[8140]), .Z(n44725) );
  NAND U45317 ( .A(x[482]), .B(y[8153]), .Z(n44726) );
  NAND U45318 ( .A(x[483]), .B(y[8152]), .Z(n44728) );
  XOR U45319 ( .A(n44683), .B(n44682), .Z(n44685) );
  NAND U45320 ( .A(x[496]), .B(y[8139]), .Z(n44711) );
  XNOR U45321 ( .A(n44711), .B(n44710), .Z(n44713) );
  XOR U45322 ( .A(n44712), .B(n44713), .Z(n44721) );
  AND U45323 ( .A(y[8142]), .B(x[493]), .Z(n44542) );
  NAND U45324 ( .A(y[8143]), .B(x[492]), .Z(n44541) );
  XNOR U45325 ( .A(n44542), .B(n44541), .Z(n44722) );
  XOR U45326 ( .A(n44721), .B(n44722), .Z(n44684) );
  XOR U45327 ( .A(n44685), .B(n44684), .Z(n44689) );
  NAND U45328 ( .A(n44720), .B(n44543), .Z(n44547) );
  ANDN U45329 ( .B(n44545), .A(n44544), .Z(n44546) );
  ANDN U45330 ( .B(n44547), .A(n44546), .Z(n44687) );
  NANDN U45331 ( .A(n44549), .B(n44548), .Z(n44553) );
  NAND U45332 ( .A(n44551), .B(n44550), .Z(n44552) );
  NAND U45333 ( .A(n44553), .B(n44552), .Z(n44686) );
  XNOR U45334 ( .A(n44687), .B(n44686), .Z(n44688) );
  XOR U45335 ( .A(n44689), .B(n44688), .Z(n44633) );
  XNOR U45336 ( .A(n44632), .B(n44633), .Z(n44635) );
  XNOR U45337 ( .A(n44737), .B(n44738), .Z(n44739) );
  XOR U45338 ( .A(n44740), .B(n44739), .Z(n44614) );
  XNOR U45339 ( .A(n44615), .B(n44614), .Z(n44617) );
  XOR U45340 ( .A(n44616), .B(n44617), .Z(n44622) );
  NAND U45341 ( .A(n44555), .B(n44554), .Z(n44559) );
  NAND U45342 ( .A(n44557), .B(n44556), .Z(n44558) );
  NAND U45343 ( .A(n44559), .B(n44558), .Z(n44621) );
  NANDN U45344 ( .A(n44561), .B(n44560), .Z(n44565) );
  NANDN U45345 ( .A(n44563), .B(n44562), .Z(n44564) );
  NAND U45346 ( .A(n44565), .B(n44564), .Z(n44627) );
  NANDN U45347 ( .A(n44567), .B(n44566), .Z(n44571) );
  NAND U45348 ( .A(n44569), .B(n44568), .Z(n44570) );
  NAND U45349 ( .A(n44571), .B(n44570), .Z(n44745) );
  NAND U45350 ( .A(n44573), .B(n44572), .Z(n44577) );
  ANDN U45351 ( .B(n44575), .A(n44574), .Z(n44576) );
  ANDN U45352 ( .B(n44577), .A(n44576), .Z(n44675) );
  NANDN U45353 ( .A(n44579), .B(n44578), .Z(n44583) );
  NANDN U45354 ( .A(n44581), .B(n44580), .Z(n44582) );
  NAND U45355 ( .A(n44583), .B(n44582), .Z(n44674) );
  XNOR U45356 ( .A(n44675), .B(n44674), .Z(n44677) );
  AND U45357 ( .A(y[8148]), .B(x[488]), .Z(n44673) );
  NAND U45358 ( .A(n44584), .B(n44673), .Z(n44588) );
  NANDN U45359 ( .A(n44586), .B(n44585), .Z(n44587) );
  NAND U45360 ( .A(n44588), .B(n44587), .Z(n44700) );
  AND U45361 ( .A(x[494]), .B(y[8141]), .Z(n44731) );
  NAND U45362 ( .A(x[481]), .B(y[8154]), .Z(n44732) );
  ANDN U45363 ( .B(o[474]), .A(n44589), .Z(n44733) );
  XOR U45364 ( .A(n44734), .B(n44733), .Z(n44699) );
  AND U45365 ( .A(x[497]), .B(y[8138]), .Z(n44655) );
  NAND U45366 ( .A(x[484]), .B(y[8151]), .Z(n44656) );
  XNOR U45367 ( .A(n44655), .B(n44656), .Z(n44658) );
  AND U45368 ( .A(x[485]), .B(y[8150]), .Z(n44657) );
  XOR U45369 ( .A(n44658), .B(n44657), .Z(n44698) );
  XOR U45370 ( .A(n44699), .B(n44698), .Z(n44701) );
  XOR U45371 ( .A(n44700), .B(n44701), .Z(n44676) );
  XOR U45372 ( .A(n44677), .B(n44676), .Z(n44744) );
  NANDN U45373 ( .A(n44591), .B(n44590), .Z(n44595) );
  NANDN U45374 ( .A(n44593), .B(n44592), .Z(n44594) );
  AND U45375 ( .A(n44595), .B(n44594), .Z(n44681) );
  AND U45376 ( .A(y[8131]), .B(x[504]), .Z(n44597) );
  NAND U45377 ( .A(y[8135]), .B(x[500]), .Z(n44596) );
  XNOR U45378 ( .A(n44597), .B(n44596), .Z(n44645) );
  NAND U45379 ( .A(x[487]), .B(y[8148]), .Z(n44646) );
  XNOR U45380 ( .A(n44645), .B(n44646), .Z(n44679) );
  AND U45381 ( .A(x[488]), .B(y[8147]), .Z(n44714) );
  NAND U45382 ( .A(x[503]), .B(y[8132]), .Z(n44715) );
  NAND U45383 ( .A(x[502]), .B(y[8133]), .Z(n44717) );
  XOR U45384 ( .A(n44679), .B(n44678), .Z(n44680) );
  XNOR U45385 ( .A(n44681), .B(n44680), .Z(n44743) );
  XOR U45386 ( .A(n44744), .B(n44743), .Z(n44746) );
  XNOR U45387 ( .A(n44745), .B(n44746), .Z(n44626) );
  XOR U45388 ( .A(n44627), .B(n44626), .Z(n44629) );
  NANDN U45389 ( .A(n44599), .B(n44598), .Z(n44603) );
  NANDN U45390 ( .A(n44601), .B(n44600), .Z(n44602) );
  AND U45391 ( .A(n44603), .B(n44602), .Z(n44628) );
  XOR U45392 ( .A(n44629), .B(n44628), .Z(n44620) );
  XOR U45393 ( .A(n44621), .B(n44620), .Z(n44623) );
  XOR U45394 ( .A(n44622), .B(n44623), .Z(n44755) );
  XOR U45395 ( .A(n44756), .B(n44755), .Z(n44757) );
  XNOR U45396 ( .A(n44758), .B(n44757), .Z(n44764) );
  NAND U45397 ( .A(n44608), .B(n44607), .Z(n44612) );
  NAND U45398 ( .A(n44610), .B(n44609), .Z(n44611) );
  AND U45399 ( .A(n44612), .B(n44611), .Z(n44763) );
  IV U45400 ( .A(n44763), .Z(n44761) );
  XOR U45401 ( .A(n44762), .B(n44761), .Z(n44613) );
  XNOR U45402 ( .A(n44764), .B(n44613), .Z(N956) );
  NAND U45403 ( .A(n44615), .B(n44614), .Z(n44619) );
  NANDN U45404 ( .A(n44617), .B(n44616), .Z(n44618) );
  NAND U45405 ( .A(n44619), .B(n44618), .Z(n44925) );
  NAND U45406 ( .A(n44621), .B(n44620), .Z(n44625) );
  NAND U45407 ( .A(n44623), .B(n44622), .Z(n44624) );
  AND U45408 ( .A(n44625), .B(n44624), .Z(n44924) );
  XOR U45409 ( .A(n44925), .B(n44924), .Z(n44927) );
  NAND U45410 ( .A(n44627), .B(n44626), .Z(n44631) );
  NAND U45411 ( .A(n44629), .B(n44628), .Z(n44630) );
  AND U45412 ( .A(n44631), .B(n44630), .Z(n44770) );
  NAND U45413 ( .A(n44633), .B(n44632), .Z(n44637) );
  NANDN U45414 ( .A(n44635), .B(n44634), .Z(n44636) );
  NAND U45415 ( .A(n44637), .B(n44636), .Z(n44782) );
  NAND U45416 ( .A(n44639), .B(n44638), .Z(n44643) );
  NAND U45417 ( .A(n44641), .B(n44640), .Z(n44642) );
  NAND U45418 ( .A(n44643), .B(n44642), .Z(n44781) );
  XOR U45419 ( .A(n44782), .B(n44781), .Z(n44784) );
  AND U45420 ( .A(x[504]), .B(y[8135]), .Z(n45179) );
  AND U45421 ( .A(x[500]), .B(y[8131]), .Z(n44644) );
  NAND U45422 ( .A(n45179), .B(n44644), .Z(n44648) );
  NANDN U45423 ( .A(n44646), .B(n44645), .Z(n44647) );
  AND U45424 ( .A(n44648), .B(n44647), .Z(n44921) );
  AND U45425 ( .A(x[505]), .B(y[8131]), .Z(n44848) );
  XOR U45426 ( .A(n44849), .B(n44848), .Z(n44847) );
  NAND U45427 ( .A(x[481]), .B(y[8155]), .Z(n44846) );
  AND U45428 ( .A(x[496]), .B(y[8140]), .Z(n44840) );
  NAND U45429 ( .A(x[504]), .B(y[8132]), .Z(n44841) );
  NAND U45430 ( .A(x[482]), .B(y[8154]), .Z(n44843) );
  XOR U45431 ( .A(n44919), .B(n44918), .Z(n44920) );
  NANDN U45432 ( .A(n44650), .B(n44649), .Z(n44654) );
  NANDN U45433 ( .A(n44652), .B(n44651), .Z(n44653) );
  AND U45434 ( .A(n44654), .B(n44653), .Z(n44915) );
  NAND U45435 ( .A(x[483]), .B(y[8153]), .Z(n44865) );
  NAND U45436 ( .A(x[503]), .B(y[8133]), .Z(n44867) );
  AND U45437 ( .A(x[485]), .B(y[8151]), .Z(n44833) );
  NAND U45438 ( .A(x[501]), .B(y[8135]), .Z(n44834) );
  NAND U45439 ( .A(x[500]), .B(y[8136]), .Z(n44836) );
  XOR U45440 ( .A(n44913), .B(n44912), .Z(n44914) );
  NANDN U45441 ( .A(n44656), .B(n44655), .Z(n44660) );
  NAND U45442 ( .A(n44658), .B(n44657), .Z(n44659) );
  AND U45443 ( .A(n44660), .B(n44659), .Z(n44907) );
  NANDN U45444 ( .A(n44666), .B(n44665), .Z(n44670) );
  NANDN U45445 ( .A(n44668), .B(n44667), .Z(n44669) );
  AND U45446 ( .A(n44670), .B(n44669), .Z(n44802) );
  ANDN U45447 ( .B(o[475]), .A(n44671), .Z(n44814) );
  AND U45448 ( .A(x[480]), .B(y[8156]), .Z(n44812) );
  AND U45449 ( .A(x[508]), .B(y[8128]), .Z(n44811) );
  XOR U45450 ( .A(n44812), .B(n44811), .Z(n44813) );
  XOR U45451 ( .A(n44814), .B(n44813), .Z(n44800) );
  NAND U45452 ( .A(y[8146]), .B(x[490]), .Z(n44672) );
  XNOR U45453 ( .A(n44673), .B(n44672), .Z(n44819) );
  AND U45454 ( .A(x[489]), .B(y[8147]), .Z(n44818) );
  XOR U45455 ( .A(n44819), .B(n44818), .Z(n44799) );
  XOR U45456 ( .A(n44800), .B(n44799), .Z(n44801) );
  XNOR U45457 ( .A(n44909), .B(n44908), .Z(n44890) );
  XOR U45458 ( .A(n44891), .B(n44890), .Z(n44892) );
  XOR U45459 ( .A(n44893), .B(n44892), .Z(n44788) );
  XNOR U45460 ( .A(n44885), .B(n44884), .Z(n44886) );
  XNOR U45461 ( .A(n44887), .B(n44886), .Z(n44787) );
  NANDN U45462 ( .A(n44687), .B(n44686), .Z(n44691) );
  NAND U45463 ( .A(n44689), .B(n44688), .Z(n44690) );
  AND U45464 ( .A(n44691), .B(n44690), .Z(n44794) );
  NANDN U45465 ( .A(n44693), .B(n44692), .Z(n44697) );
  NANDN U45466 ( .A(n44695), .B(n44694), .Z(n44696) );
  AND U45467 ( .A(n44697), .B(n44696), .Z(n44899) );
  NAND U45468 ( .A(n44699), .B(n44698), .Z(n44703) );
  NAND U45469 ( .A(n44701), .B(n44700), .Z(n44702) );
  AND U45470 ( .A(n44703), .B(n44702), .Z(n44897) );
  NANDN U45471 ( .A(n44705), .B(n44704), .Z(n44709) );
  NANDN U45472 ( .A(n44707), .B(n44706), .Z(n44708) );
  NAND U45473 ( .A(n44709), .B(n44708), .Z(n44896) );
  XNOR U45474 ( .A(n44897), .B(n44896), .Z(n44898) );
  XNOR U45475 ( .A(n44899), .B(n44898), .Z(n44793) );
  XNOR U45476 ( .A(n44794), .B(n44793), .Z(n44796) );
  AND U45477 ( .A(x[495]), .B(y[8141]), .Z(n44873) );
  NAND U45478 ( .A(x[507]), .B(y[8129]), .Z(n44839) );
  AND U45479 ( .A(x[506]), .B(y[8130]), .Z(n44870) );
  XOR U45480 ( .A(n44871), .B(n44870), .Z(n44872) );
  XOR U45481 ( .A(n44873), .B(n44872), .Z(n44859) );
  AND U45482 ( .A(x[487]), .B(y[8149]), .Z(n44852) );
  NAND U45483 ( .A(x[492]), .B(y[8144]), .Z(n44853) );
  AND U45484 ( .A(x[491]), .B(y[8145]), .Z(n44854) );
  XNOR U45485 ( .A(n44855), .B(n44854), .Z(n44858) );
  AND U45486 ( .A(x[497]), .B(y[8139]), .Z(n44805) );
  NAND U45487 ( .A(x[502]), .B(y[8134]), .Z(n44806) );
  NAND U45488 ( .A(x[484]), .B(y[8152]), .Z(n44808) );
  AND U45489 ( .A(x[486]), .B(y[8150]), .Z(n45032) );
  NAND U45490 ( .A(x[499]), .B(y[8137]), .Z(n44828) );
  XOR U45491 ( .A(n44879), .B(n44878), .Z(n44880) );
  NANDN U45492 ( .A(n44715), .B(n44714), .Z(n44719) );
  NANDN U45493 ( .A(n44717), .B(n44716), .Z(n44718) );
  AND U45494 ( .A(n44719), .B(n44718), .Z(n44881) );
  XOR U45495 ( .A(n44903), .B(n44902), .Z(n44905) );
  NAND U45496 ( .A(n44864), .B(n44720), .Z(n44724) );
  NAND U45497 ( .A(n44722), .B(n44721), .Z(n44723) );
  AND U45498 ( .A(n44724), .B(n44723), .Z(n44825) );
  NANDN U45499 ( .A(n44726), .B(n44725), .Z(n44730) );
  NANDN U45500 ( .A(n44728), .B(n44727), .Z(n44729) );
  AND U45501 ( .A(n44730), .B(n44729), .Z(n44823) );
  NANDN U45502 ( .A(n44732), .B(n44731), .Z(n44736) );
  NAND U45503 ( .A(n44734), .B(n44733), .Z(n44735) );
  NAND U45504 ( .A(n44736), .B(n44735), .Z(n44822) );
  XOR U45505 ( .A(n44905), .B(n44904), .Z(n44795) );
  XOR U45506 ( .A(n44796), .B(n44795), .Z(n44789) );
  XOR U45507 ( .A(n44790), .B(n44789), .Z(n44783) );
  XOR U45508 ( .A(n44784), .B(n44783), .Z(n44769) );
  XOR U45509 ( .A(n44770), .B(n44769), .Z(n44771) );
  NANDN U45510 ( .A(n44738), .B(n44737), .Z(n44742) );
  NAND U45511 ( .A(n44740), .B(n44739), .Z(n44741) );
  NAND U45512 ( .A(n44742), .B(n44741), .Z(n44777) );
  NAND U45513 ( .A(n44744), .B(n44743), .Z(n44748) );
  NAND U45514 ( .A(n44746), .B(n44745), .Z(n44747) );
  NAND U45515 ( .A(n44748), .B(n44747), .Z(n44775) );
  NAND U45516 ( .A(n44750), .B(n44749), .Z(n44754) );
  NANDN U45517 ( .A(n44752), .B(n44751), .Z(n44753) );
  AND U45518 ( .A(n44754), .B(n44753), .Z(n44776) );
  XNOR U45519 ( .A(n44775), .B(n44776), .Z(n44778) );
  XNOR U45520 ( .A(n44771), .B(n44772), .Z(n44926) );
  XOR U45521 ( .A(n44927), .B(n44926), .Z(n44932) );
  NAND U45522 ( .A(n44756), .B(n44755), .Z(n44760) );
  NAND U45523 ( .A(n44758), .B(n44757), .Z(n44759) );
  NAND U45524 ( .A(n44760), .B(n44759), .Z(n44930) );
  NANDN U45525 ( .A(n44761), .B(n44762), .Z(n44767) );
  NOR U45526 ( .A(n44763), .B(n44762), .Z(n44765) );
  OR U45527 ( .A(n44765), .B(n44764), .Z(n44766) );
  AND U45528 ( .A(n44767), .B(n44766), .Z(n44931) );
  XOR U45529 ( .A(n44930), .B(n44931), .Z(n44768) );
  XNOR U45530 ( .A(n44932), .B(n44768), .Z(N957) );
  NAND U45531 ( .A(n44770), .B(n44769), .Z(n44774) );
  NANDN U45532 ( .A(n44772), .B(n44771), .Z(n44773) );
  NAND U45533 ( .A(n44774), .B(n44773), .Z(n44939) );
  NAND U45534 ( .A(n44776), .B(n44775), .Z(n44780) );
  NANDN U45535 ( .A(n44778), .B(n44777), .Z(n44779) );
  NAND U45536 ( .A(n44780), .B(n44779), .Z(n44937) );
  NAND U45537 ( .A(n44782), .B(n44781), .Z(n44786) );
  NAND U45538 ( .A(n44784), .B(n44783), .Z(n44785) );
  NAND U45539 ( .A(n44786), .B(n44785), .Z(n44944) );
  NANDN U45540 ( .A(n44788), .B(n44787), .Z(n44792) );
  NAND U45541 ( .A(n44790), .B(n44789), .Z(n44791) );
  NAND U45542 ( .A(n44792), .B(n44791), .Z(n44943) );
  XOR U45543 ( .A(n44944), .B(n44943), .Z(n44946) );
  NANDN U45544 ( .A(n44794), .B(n44793), .Z(n44798) );
  NAND U45545 ( .A(n44796), .B(n44795), .Z(n44797) );
  AND U45546 ( .A(n44798), .B(n44797), .Z(n44954) );
  NAND U45547 ( .A(n44800), .B(n44799), .Z(n44804) );
  NANDN U45548 ( .A(n44802), .B(n44801), .Z(n44803) );
  AND U45549 ( .A(n44804), .B(n44803), .Z(n45063) );
  NANDN U45550 ( .A(n44806), .B(n44805), .Z(n44810) );
  NANDN U45551 ( .A(n44808), .B(n44807), .Z(n44809) );
  NAND U45552 ( .A(n44810), .B(n44809), .Z(n45103) );
  NAND U45553 ( .A(n44812), .B(n44811), .Z(n44816) );
  NAND U45554 ( .A(n44814), .B(n44813), .Z(n44815) );
  NAND U45555 ( .A(n44816), .B(n44815), .Z(n45102) );
  XOR U45556 ( .A(n45103), .B(n45102), .Z(n45105) );
  AND U45557 ( .A(y[8148]), .B(x[490]), .Z(n45100) );
  NAND U45558 ( .A(n44817), .B(n45100), .Z(n44821) );
  NAND U45559 ( .A(n44819), .B(n44818), .Z(n44820) );
  NAND U45560 ( .A(n44821), .B(n44820), .Z(n45071) );
  AND U45561 ( .A(x[502]), .B(y[8135]), .Z(n45010) );
  AND U45562 ( .A(x[492]), .B(y[8145]), .Z(n45280) );
  AND U45563 ( .A(x[481]), .B(y[8156]), .Z(n45008) );
  XOR U45564 ( .A(n45280), .B(n45008), .Z(n45009) );
  XOR U45565 ( .A(n45010), .B(n45009), .Z(n45070) );
  AND U45566 ( .A(x[495]), .B(y[8142]), .Z(n45013) );
  XOR U45567 ( .A(n45013), .B(n45169), .Z(n45015) );
  XOR U45568 ( .A(n45015), .B(n45014), .Z(n45069) );
  XOR U45569 ( .A(n45070), .B(n45069), .Z(n45072) );
  XOR U45570 ( .A(n45071), .B(n45072), .Z(n45104) );
  XOR U45571 ( .A(n45105), .B(n45104), .Z(n45064) );
  NANDN U45572 ( .A(n44823), .B(n44822), .Z(n44827) );
  NANDN U45573 ( .A(n44825), .B(n44824), .Z(n44826) );
  AND U45574 ( .A(n44827), .B(n44826), .Z(n45065) );
  XOR U45575 ( .A(n45066), .B(n45065), .Z(n45060) );
  NANDN U45576 ( .A(n44828), .B(n45032), .Z(n44832) );
  NANDN U45577 ( .A(n44830), .B(n44829), .Z(n44831) );
  AND U45578 ( .A(n44832), .B(n44831), .Z(n45084) );
  AND U45579 ( .A(x[505]), .B(y[8132]), .Z(n45005) );
  AND U45580 ( .A(x[506]), .B(y[8131]), .Z(n45002) );
  XOR U45581 ( .A(n45003), .B(n45002), .Z(n45004) );
  XOR U45582 ( .A(n45005), .B(n45004), .Z(n45082) );
  AND U45583 ( .A(x[508]), .B(y[8129]), .Z(n45020) );
  XOR U45584 ( .A(o[477]), .B(n45020), .Z(n45095) );
  AND U45585 ( .A(x[480]), .B(y[8157]), .Z(n45093) );
  AND U45586 ( .A(x[509]), .B(y[8128]), .Z(n45092) );
  XOR U45587 ( .A(n45093), .B(n45092), .Z(n45094) );
  XNOR U45588 ( .A(n45095), .B(n45094), .Z(n45081) );
  XOR U45589 ( .A(n45084), .B(n45083), .Z(n45051) );
  NANDN U45590 ( .A(n44834), .B(n44833), .Z(n44838) );
  NANDN U45591 ( .A(n44836), .B(n44835), .Z(n44837) );
  NAND U45592 ( .A(n44838), .B(n44837), .Z(n45041) );
  ANDN U45593 ( .B(o[476]), .A(n44839), .Z(n44981) );
  AND U45594 ( .A(x[496]), .B(y[8141]), .Z(n44979) );
  AND U45595 ( .A(x[507]), .B(y[8130]), .Z(n44978) );
  XOR U45596 ( .A(n44979), .B(n44978), .Z(n44980) );
  XOR U45597 ( .A(n44981), .B(n44980), .Z(n45040) );
  AND U45598 ( .A(x[482]), .B(y[8155]), .Z(n44991) );
  XOR U45599 ( .A(n44991), .B(n44990), .Z(n44992) );
  XOR U45600 ( .A(n44993), .B(n44992), .Z(n45039) );
  XOR U45601 ( .A(n45040), .B(n45039), .Z(n45042) );
  XOR U45602 ( .A(n45041), .B(n45042), .Z(n45052) );
  NANDN U45603 ( .A(n44841), .B(n44840), .Z(n44845) );
  NANDN U45604 ( .A(n44843), .B(n44842), .Z(n44844) );
  AND U45605 ( .A(n44845), .B(n44844), .Z(n45076) );
  ANDN U45606 ( .B(n44847), .A(n44846), .Z(n44851) );
  NAND U45607 ( .A(n44849), .B(n44848), .Z(n44850) );
  NANDN U45608 ( .A(n44851), .B(n44850), .Z(n45075) );
  NANDN U45609 ( .A(n44853), .B(n44852), .Z(n44857) );
  NAND U45610 ( .A(n44855), .B(n44854), .Z(n44856) );
  NAND U45611 ( .A(n44857), .B(n44856), .Z(n44974) );
  AND U45612 ( .A(x[491]), .B(y[8146]), .Z(n45029) );
  AND U45613 ( .A(x[483]), .B(y[8154]), .Z(n45027) );
  AND U45614 ( .A(x[497]), .B(y[8140]), .Z(n45026) );
  XOR U45615 ( .A(n45027), .B(n45026), .Z(n45028) );
  XOR U45616 ( .A(n45029), .B(n45028), .Z(n44973) );
  AND U45617 ( .A(x[503]), .B(y[8134]), .Z(n45023) );
  AND U45618 ( .A(x[493]), .B(y[8144]), .Z(n45021) );
  AND U45619 ( .A(x[504]), .B(y[8133]), .Z(n45236) );
  XOR U45620 ( .A(n45021), .B(n45236), .Z(n45022) );
  XOR U45621 ( .A(n45023), .B(n45022), .Z(n44972) );
  XOR U45622 ( .A(n44973), .B(n44972), .Z(n44975) );
  XOR U45623 ( .A(n44974), .B(n44975), .Z(n45077) );
  XOR U45624 ( .A(n45078), .B(n45077), .Z(n45054) );
  NANDN U45625 ( .A(n44859), .B(n44858), .Z(n44863) );
  NANDN U45626 ( .A(n44861), .B(n44860), .Z(n44862) );
  NAND U45627 ( .A(n44863), .B(n44862), .Z(n44967) );
  NANDN U45628 ( .A(n44865), .B(n44864), .Z(n44869) );
  NANDN U45629 ( .A(n44867), .B(n44866), .Z(n44868) );
  NAND U45630 ( .A(n44869), .B(n44868), .Z(n44997) );
  NAND U45631 ( .A(n44871), .B(n44870), .Z(n44875) );
  NAND U45632 ( .A(n44873), .B(n44872), .Z(n44874) );
  NAND U45633 ( .A(n44875), .B(n44874), .Z(n44996) );
  XOR U45634 ( .A(n44997), .B(n44996), .Z(n44999) );
  AND U45635 ( .A(x[488]), .B(y[8149]), .Z(n45034) );
  AND U45636 ( .A(x[486]), .B(y[8151]), .Z(n44877) );
  AND U45637 ( .A(y[8150]), .B(x[487]), .Z(n44876) );
  XOR U45638 ( .A(n44877), .B(n44876), .Z(n45033) );
  XOR U45639 ( .A(n45034), .B(n45033), .Z(n45087) );
  NAND U45640 ( .A(x[489]), .B(y[8148]), .Z(n45176) );
  AND U45641 ( .A(x[485]), .B(y[8152]), .Z(n44987) );
  AND U45642 ( .A(x[484]), .B(y[8153]), .Z(n44985) );
  AND U45643 ( .A(x[490]), .B(y[8147]), .Z(n44984) );
  XOR U45644 ( .A(n44985), .B(n44984), .Z(n44986) );
  XOR U45645 ( .A(n44987), .B(n44986), .Z(n45088) );
  XOR U45646 ( .A(n45089), .B(n45088), .Z(n44998) );
  XNOR U45647 ( .A(n44999), .B(n44998), .Z(n44966) );
  XOR U45648 ( .A(n44967), .B(n44966), .Z(n44968) );
  XOR U45649 ( .A(n44969), .B(n44968), .Z(n45058) );
  NAND U45650 ( .A(n44879), .B(n44878), .Z(n44883) );
  NANDN U45651 ( .A(n44881), .B(n44880), .Z(n44882) );
  NAND U45652 ( .A(n44883), .B(n44882), .Z(n45057) );
  XNOR U45653 ( .A(n44954), .B(n44953), .Z(n44956) );
  NANDN U45654 ( .A(n44885), .B(n44884), .Z(n44889) );
  NANDN U45655 ( .A(n44887), .B(n44886), .Z(n44888) );
  AND U45656 ( .A(n44889), .B(n44888), .Z(n44950) );
  NAND U45657 ( .A(n44891), .B(n44890), .Z(n44895) );
  NAND U45658 ( .A(n44893), .B(n44892), .Z(n44894) );
  AND U45659 ( .A(n44895), .B(n44894), .Z(n44949) );
  XNOR U45660 ( .A(n44950), .B(n44949), .Z(n44952) );
  NANDN U45661 ( .A(n44897), .B(n44896), .Z(n44901) );
  NANDN U45662 ( .A(n44899), .B(n44898), .Z(n44900) );
  NAND U45663 ( .A(n44901), .B(n44900), .Z(n44962) );
  NANDN U45664 ( .A(n44907), .B(n44906), .Z(n44911) );
  NAND U45665 ( .A(n44909), .B(n44908), .Z(n44910) );
  AND U45666 ( .A(n44911), .B(n44910), .Z(n45048) );
  NAND U45667 ( .A(n44913), .B(n44912), .Z(n44917) );
  NANDN U45668 ( .A(n44915), .B(n44914), .Z(n44916) );
  AND U45669 ( .A(n44917), .B(n44916), .Z(n45046) );
  NAND U45670 ( .A(n44919), .B(n44918), .Z(n44923) );
  NANDN U45671 ( .A(n44921), .B(n44920), .Z(n44922) );
  NAND U45672 ( .A(n44923), .B(n44922), .Z(n45045) );
  XOR U45673 ( .A(n44960), .B(n44961), .Z(n44963) );
  XOR U45674 ( .A(n44962), .B(n44963), .Z(n44951) );
  XOR U45675 ( .A(n44952), .B(n44951), .Z(n44955) );
  XOR U45676 ( .A(n44956), .B(n44955), .Z(n44945) );
  XOR U45677 ( .A(n44946), .B(n44945), .Z(n44938) );
  XNOR U45678 ( .A(n44937), .B(n44938), .Z(n44940) );
  XOR U45679 ( .A(n44939), .B(n44940), .Z(n44936) );
  NAND U45680 ( .A(n44925), .B(n44924), .Z(n44929) );
  NAND U45681 ( .A(n44927), .B(n44926), .Z(n44928) );
  NAND U45682 ( .A(n44929), .B(n44928), .Z(n44935) );
  XOR U45683 ( .A(n44935), .B(n44934), .Z(n44933) );
  XNOR U45684 ( .A(n44936), .B(n44933), .Z(N958) );
  NAND U45685 ( .A(n44938), .B(n44937), .Z(n44942) );
  NANDN U45686 ( .A(n44940), .B(n44939), .Z(n44941) );
  NAND U45687 ( .A(n44942), .B(n44941), .Z(n45366) );
  NAND U45688 ( .A(n44944), .B(n44943), .Z(n44948) );
  NAND U45689 ( .A(n44946), .B(n44945), .Z(n44947) );
  NAND U45690 ( .A(n44948), .B(n44947), .Z(n45369) );
  NANDN U45691 ( .A(n44954), .B(n44953), .Z(n44959) );
  IV U45692 ( .A(n44955), .Z(n44957) );
  NANDN U45693 ( .A(n44957), .B(n44956), .Z(n44958) );
  NAND U45694 ( .A(n44959), .B(n44958), .Z(n45111) );
  NAND U45695 ( .A(n44961), .B(n44960), .Z(n44965) );
  NAND U45696 ( .A(n44963), .B(n44962), .Z(n44964) );
  AND U45697 ( .A(n44965), .B(n44964), .Z(n45108) );
  XOR U45698 ( .A(n45109), .B(n45108), .Z(n45372) );
  NAND U45699 ( .A(n44967), .B(n44966), .Z(n44971) );
  NAND U45700 ( .A(n44969), .B(n44968), .Z(n44970) );
  AND U45701 ( .A(n44971), .B(n44970), .Z(n45351) );
  NAND U45702 ( .A(n44973), .B(n44972), .Z(n44977) );
  NAND U45703 ( .A(n44975), .B(n44974), .Z(n44976) );
  AND U45704 ( .A(n44977), .B(n44976), .Z(n45117) );
  NAND U45705 ( .A(n44979), .B(n44978), .Z(n44983) );
  NAND U45706 ( .A(n44981), .B(n44980), .Z(n44982) );
  NAND U45707 ( .A(n44983), .B(n44982), .Z(n45127) );
  NAND U45708 ( .A(n44985), .B(n44984), .Z(n44989) );
  NAND U45709 ( .A(n44987), .B(n44986), .Z(n44988) );
  NAND U45710 ( .A(n44989), .B(n44988), .Z(n45130) );
  AND U45711 ( .A(x[486]), .B(y[8152]), .Z(n45240) );
  AND U45712 ( .A(x[485]), .B(y[8153]), .Z(n45242) );
  AND U45713 ( .A(x[499]), .B(y[8139]), .Z(n45241) );
  XOR U45714 ( .A(n45242), .B(n45241), .Z(n45239) );
  XNOR U45715 ( .A(n45240), .B(n45239), .Z(n45272) );
  AND U45716 ( .A(x[484]), .B(y[8154]), .Z(n45298) );
  AND U45717 ( .A(x[483]), .B(y[8155]), .Z(n45300) );
  AND U45718 ( .A(x[498]), .B(y[8140]), .Z(n45299) );
  XOR U45719 ( .A(n45300), .B(n45299), .Z(n45297) );
  XOR U45720 ( .A(n45298), .B(n45297), .Z(n45269) );
  NAND U45721 ( .A(n44991), .B(n44990), .Z(n44995) );
  NAND U45722 ( .A(n44993), .B(n44992), .Z(n44994) );
  AND U45723 ( .A(n44995), .B(n44994), .Z(n45270) );
  XOR U45724 ( .A(n45272), .B(n45271), .Z(n45129) );
  XOR U45725 ( .A(n45130), .B(n45129), .Z(n45128) );
  XOR U45726 ( .A(n45127), .B(n45128), .Z(n45118) );
  NAND U45727 ( .A(n44997), .B(n44996), .Z(n45001) );
  NAND U45728 ( .A(n44999), .B(n44998), .Z(n45000) );
  AND U45729 ( .A(n45001), .B(n45000), .Z(n45114) );
  XOR U45730 ( .A(n45115), .B(n45114), .Z(n45354) );
  AND U45731 ( .A(n45003), .B(n45002), .Z(n45007) );
  NAND U45732 ( .A(n45005), .B(n45004), .Z(n45006) );
  NANDN U45733 ( .A(n45007), .B(n45006), .Z(n45153) );
  AND U45734 ( .A(n45280), .B(n45008), .Z(n45012) );
  NAND U45735 ( .A(n45010), .B(n45009), .Z(n45011) );
  NANDN U45736 ( .A(n45012), .B(n45011), .Z(n45156) );
  NAND U45737 ( .A(n45013), .B(n45169), .Z(n45017) );
  NAND U45738 ( .A(n45015), .B(n45014), .Z(n45016) );
  AND U45739 ( .A(n45017), .B(n45016), .Z(n45134) );
  AND U45740 ( .A(x[503]), .B(y[8135]), .Z(n45234) );
  AND U45741 ( .A(y[8134]), .B(x[504]), .Z(n45019) );
  AND U45742 ( .A(y[8133]), .B(x[505]), .Z(n45018) );
  XOR U45743 ( .A(n45019), .B(n45018), .Z(n45233) );
  XOR U45744 ( .A(n45234), .B(n45233), .Z(n45136) );
  AND U45745 ( .A(n45020), .B(o[477]), .Z(n45228) );
  AND U45746 ( .A(x[508]), .B(y[8130]), .Z(n45230) );
  AND U45747 ( .A(x[496]), .B(y[8142]), .Z(n45229) );
  XOR U45748 ( .A(n45230), .B(n45229), .Z(n45227) );
  XNOR U45749 ( .A(n45228), .B(n45227), .Z(n45135) );
  XNOR U45750 ( .A(n45134), .B(n45133), .Z(n45155) );
  XOR U45751 ( .A(n45156), .B(n45155), .Z(n45154) );
  XOR U45752 ( .A(n45153), .B(n45154), .Z(n45334) );
  NAND U45753 ( .A(n45021), .B(n45236), .Z(n45025) );
  NAND U45754 ( .A(n45023), .B(n45022), .Z(n45024) );
  NAND U45755 ( .A(n45025), .B(n45024), .Z(n45124) );
  NAND U45756 ( .A(n45027), .B(n45026), .Z(n45031) );
  NAND U45757 ( .A(n45029), .B(n45028), .Z(n45030) );
  AND U45758 ( .A(n45031), .B(n45030), .Z(n45146) );
  AND U45759 ( .A(x[480]), .B(y[8158]), .Z(n45158) );
  AND U45760 ( .A(x[509]), .B(y[8129]), .Z(n45177) );
  XOR U45761 ( .A(o[478]), .B(n45177), .Z(n45160) );
  AND U45762 ( .A(x[510]), .B(y[8128]), .Z(n45159) );
  XOR U45763 ( .A(n45160), .B(n45159), .Z(n45157) );
  XOR U45764 ( .A(n45158), .B(n45157), .Z(n45148) );
  AND U45765 ( .A(x[500]), .B(y[8138]), .Z(n45285) );
  XOR U45766 ( .A(n45286), .B(n45285), .Z(n45284) );
  AND U45767 ( .A(x[488]), .B(y[8150]), .Z(n45283) );
  XNOR U45768 ( .A(n45284), .B(n45283), .Z(n45147) );
  XNOR U45769 ( .A(n45146), .B(n45145), .Z(n45123) );
  XOR U45770 ( .A(n45124), .B(n45123), .Z(n45121) );
  AND U45771 ( .A(x[487]), .B(y[8151]), .Z(n45168) );
  NAND U45772 ( .A(n45032), .B(n45168), .Z(n45036) );
  NAND U45773 ( .A(n45034), .B(n45033), .Z(n45035) );
  AND U45774 ( .A(n45036), .B(n45035), .Z(n45139) );
  AND U45775 ( .A(y[8137]), .B(x[501]), .Z(n45038) );
  AND U45776 ( .A(y[8136]), .B(x[502]), .Z(n45037) );
  XOR U45777 ( .A(n45038), .B(n45037), .Z(n45167) );
  XOR U45778 ( .A(n45168), .B(n45167), .Z(n45142) );
  AND U45779 ( .A(x[497]), .B(y[8141]), .Z(n45292) );
  AND U45780 ( .A(x[482]), .B(y[8156]), .Z(n45294) );
  AND U45781 ( .A(x[506]), .B(y[8132]), .Z(n45293) );
  XOR U45782 ( .A(n45294), .B(n45293), .Z(n45291) );
  XNOR U45783 ( .A(n45292), .B(n45291), .Z(n45141) );
  XNOR U45784 ( .A(n45139), .B(n45140), .Z(n45122) );
  XNOR U45785 ( .A(n45121), .B(n45122), .Z(n45336) );
  NAND U45786 ( .A(n45040), .B(n45039), .Z(n45044) );
  NAND U45787 ( .A(n45042), .B(n45041), .Z(n45043) );
  NAND U45788 ( .A(n45044), .B(n45043), .Z(n45335) );
  XOR U45789 ( .A(n45336), .B(n45335), .Z(n45333) );
  XOR U45790 ( .A(n45334), .B(n45333), .Z(n45353) );
  XNOR U45791 ( .A(n45351), .B(n45352), .Z(n45346) );
  NANDN U45792 ( .A(n45046), .B(n45045), .Z(n45050) );
  NANDN U45793 ( .A(n45048), .B(n45047), .Z(n45049) );
  AND U45794 ( .A(n45050), .B(n45049), .Z(n45348) );
  NANDN U45795 ( .A(n45052), .B(n45051), .Z(n45056) );
  NANDN U45796 ( .A(n45054), .B(n45053), .Z(n45055) );
  NAND U45797 ( .A(n45056), .B(n45055), .Z(n45347) );
  XOR U45798 ( .A(n45348), .B(n45347), .Z(n45345) );
  XOR U45799 ( .A(n45346), .B(n45345), .Z(n45381) );
  NANDN U45800 ( .A(n45058), .B(n45057), .Z(n45062) );
  NANDN U45801 ( .A(n45060), .B(n45059), .Z(n45061) );
  AND U45802 ( .A(n45062), .B(n45061), .Z(n45384) );
  NANDN U45803 ( .A(n45064), .B(n45063), .Z(n45068) );
  NAND U45804 ( .A(n45066), .B(n45065), .Z(n45067) );
  AND U45805 ( .A(n45068), .B(n45067), .Z(n45327) );
  NAND U45806 ( .A(n45070), .B(n45069), .Z(n45074) );
  NAND U45807 ( .A(n45072), .B(n45071), .Z(n45073) );
  AND U45808 ( .A(n45074), .B(n45073), .Z(n45318) );
  NANDN U45809 ( .A(n45076), .B(n45075), .Z(n45080) );
  NAND U45810 ( .A(n45078), .B(n45077), .Z(n45079) );
  AND U45811 ( .A(n45080), .B(n45079), .Z(n45317) );
  XOR U45812 ( .A(n45318), .B(n45317), .Z(n45316) );
  NANDN U45813 ( .A(n45082), .B(n45081), .Z(n45086) );
  NAND U45814 ( .A(n45084), .B(n45083), .Z(n45085) );
  NAND U45815 ( .A(n45086), .B(n45085), .Z(n45315) );
  XOR U45816 ( .A(n45316), .B(n45315), .Z(n45330) );
  NANDN U45817 ( .A(n45176), .B(n45087), .Z(n45091) );
  NAND U45818 ( .A(n45089), .B(n45088), .Z(n45090) );
  AND U45819 ( .A(n45091), .B(n45090), .Z(n45311) );
  NAND U45820 ( .A(n45093), .B(n45092), .Z(n45097) );
  NAND U45821 ( .A(n45095), .B(n45094), .Z(n45096) );
  NAND U45822 ( .A(n45097), .B(n45096), .Z(n45265) );
  AND U45823 ( .A(y[8146]), .B(x[492]), .Z(n45098) );
  XOR U45824 ( .A(n45099), .B(n45098), .Z(n45277) );
  XOR U45825 ( .A(n45278), .B(n45277), .Z(n45175) );
  AND U45826 ( .A(y[8149]), .B(x[489]), .Z(n45101) );
  XOR U45827 ( .A(n45101), .B(n45100), .Z(n45174) );
  XOR U45828 ( .A(n45175), .B(n45174), .Z(n45268) );
  AND U45829 ( .A(x[507]), .B(y[8131]), .Z(n45164) );
  AND U45830 ( .A(x[481]), .B(y[8157]), .Z(n45163) );
  XOR U45831 ( .A(n45164), .B(n45163), .Z(n45161) );
  XOR U45832 ( .A(n45162), .B(n45161), .Z(n45267) );
  XOR U45833 ( .A(n45268), .B(n45267), .Z(n45266) );
  XOR U45834 ( .A(n45265), .B(n45266), .Z(n45312) );
  NAND U45835 ( .A(n45103), .B(n45102), .Z(n45107) );
  NAND U45836 ( .A(n45105), .B(n45104), .Z(n45106) );
  AND U45837 ( .A(n45107), .B(n45106), .Z(n45310) );
  XNOR U45838 ( .A(n45309), .B(n45310), .Z(n45329) );
  XNOR U45839 ( .A(n45327), .B(n45328), .Z(n45383) );
  XOR U45840 ( .A(n45381), .B(n45382), .Z(n45371) );
  XOR U45841 ( .A(n45369), .B(n45370), .Z(n45363) );
  XNOR U45842 ( .A(n45364), .B(n45363), .Z(N959) );
  NAND U45843 ( .A(n45109), .B(n45108), .Z(n45113) );
  NANDN U45844 ( .A(n45111), .B(n45110), .Z(n45112) );
  AND U45845 ( .A(n45113), .B(n45112), .Z(n45380) );
  IV U45846 ( .A(n45114), .Z(n45116) );
  NANDN U45847 ( .A(n45116), .B(n45115), .Z(n45120) );
  NANDN U45848 ( .A(n45118), .B(n45117), .Z(n45119) );
  AND U45849 ( .A(n45120), .B(n45119), .Z(n45362) );
  NANDN U45850 ( .A(n45122), .B(n45121), .Z(n45126) );
  NAND U45851 ( .A(n45124), .B(n45123), .Z(n45125) );
  AND U45852 ( .A(n45126), .B(n45125), .Z(n45344) );
  NAND U45853 ( .A(n45128), .B(n45127), .Z(n45132) );
  NAND U45854 ( .A(n45130), .B(n45129), .Z(n45131) );
  AND U45855 ( .A(n45132), .B(n45131), .Z(n45326) );
  NAND U45856 ( .A(n45134), .B(n45133), .Z(n45138) );
  NANDN U45857 ( .A(n45136), .B(n45135), .Z(n45137) );
  AND U45858 ( .A(n45138), .B(n45137), .Z(n45308) );
  NANDN U45859 ( .A(n45140), .B(n45139), .Z(n45144) );
  NANDN U45860 ( .A(n45142), .B(n45141), .Z(n45143) );
  AND U45861 ( .A(n45144), .B(n45143), .Z(n45152) );
  NAND U45862 ( .A(n45146), .B(n45145), .Z(n45150) );
  NANDN U45863 ( .A(n45148), .B(n45147), .Z(n45149) );
  NAND U45864 ( .A(n45150), .B(n45149), .Z(n45151) );
  XNOR U45865 ( .A(n45152), .B(n45151), .Z(n45306) );
  NAND U45866 ( .A(n45162), .B(n45161), .Z(n45166) );
  NAND U45867 ( .A(n45164), .B(n45163), .Z(n45165) );
  AND U45868 ( .A(n45166), .B(n45165), .Z(n45173) );
  NAND U45869 ( .A(n45168), .B(n45167), .Z(n45171) );
  AND U45870 ( .A(x[502]), .B(y[8137]), .Z(n45178) );
  NAND U45871 ( .A(n45169), .B(n45178), .Z(n45170) );
  NAND U45872 ( .A(n45171), .B(n45170), .Z(n45172) );
  AND U45873 ( .A(x[490]), .B(y[8149]), .Z(n45200) );
  AND U45874 ( .A(y[8154]), .B(x[485]), .Z(n45185) );
  AND U45875 ( .A(n45177), .B(o[478]), .Z(n45183) );
  XOR U45876 ( .A(n45178), .B(o[479]), .Z(n45181) );
  AND U45877 ( .A(x[505]), .B(y[8134]), .Z(n45235) );
  XNOR U45878 ( .A(n45179), .B(n45235), .Z(n45180) );
  XNOR U45879 ( .A(n45181), .B(n45180), .Z(n45182) );
  XNOR U45880 ( .A(n45183), .B(n45182), .Z(n45184) );
  XNOR U45881 ( .A(n45185), .B(n45184), .Z(n45224) );
  AND U45882 ( .A(y[8143]), .B(x[496]), .Z(n45191) );
  AND U45883 ( .A(y[8148]), .B(x[491]), .Z(n45187) );
  NAND U45884 ( .A(y[8147]), .B(x[492]), .Z(n45186) );
  XNOR U45885 ( .A(n45187), .B(n45186), .Z(n45188) );
  XNOR U45886 ( .A(n45189), .B(n45188), .Z(n45190) );
  XNOR U45887 ( .A(n45191), .B(n45190), .Z(n45214) );
  AND U45888 ( .A(y[8138]), .B(x[501]), .Z(n45193) );
  NAND U45889 ( .A(y[8151]), .B(x[488]), .Z(n45192) );
  XNOR U45890 ( .A(n45193), .B(n45192), .Z(n45204) );
  AND U45891 ( .A(y[8140]), .B(x[499]), .Z(n45195) );
  NAND U45892 ( .A(y[8157]), .B(x[482]), .Z(n45194) );
  XNOR U45893 ( .A(n45195), .B(n45194), .Z(n45199) );
  AND U45894 ( .A(y[8136]), .B(x[503]), .Z(n45197) );
  NAND U45895 ( .A(y[8142]), .B(x[497]), .Z(n45196) );
  XNOR U45896 ( .A(n45197), .B(n45196), .Z(n45198) );
  XOR U45897 ( .A(n45199), .B(n45198), .Z(n45202) );
  XNOR U45898 ( .A(n45279), .B(n45200), .Z(n45201) );
  XNOR U45899 ( .A(n45202), .B(n45201), .Z(n45203) );
  XOR U45900 ( .A(n45204), .B(n45203), .Z(n45212) );
  AND U45901 ( .A(y[8153]), .B(x[486]), .Z(n45206) );
  NAND U45902 ( .A(y[8152]), .B(x[487]), .Z(n45205) );
  XNOR U45903 ( .A(n45206), .B(n45205), .Z(n45210) );
  AND U45904 ( .A(y[8128]), .B(x[511]), .Z(n45208) );
  NAND U45905 ( .A(y[8155]), .B(x[484]), .Z(n45207) );
  XNOR U45906 ( .A(n45208), .B(n45207), .Z(n45209) );
  XNOR U45907 ( .A(n45210), .B(n45209), .Z(n45211) );
  XNOR U45908 ( .A(n45212), .B(n45211), .Z(n45213) );
  XOR U45909 ( .A(n45214), .B(n45213), .Z(n45222) );
  AND U45910 ( .A(y[8132]), .B(x[507]), .Z(n45216) );
  NAND U45911 ( .A(y[8150]), .B(x[489]), .Z(n45215) );
  XNOR U45912 ( .A(n45216), .B(n45215), .Z(n45220) );
  AND U45913 ( .A(y[8145]), .B(x[494]), .Z(n45218) );
  NAND U45914 ( .A(y[8133]), .B(x[506]), .Z(n45217) );
  XNOR U45915 ( .A(n45218), .B(n45217), .Z(n45219) );
  XNOR U45916 ( .A(n45220), .B(n45219), .Z(n45221) );
  XNOR U45917 ( .A(n45222), .B(n45221), .Z(n45223) );
  XNOR U45918 ( .A(n45224), .B(n45223), .Z(n45225) );
  NAND U45919 ( .A(n45228), .B(n45227), .Z(n45232) );
  NAND U45920 ( .A(n45230), .B(n45229), .Z(n45231) );
  AND U45921 ( .A(n45232), .B(n45231), .Z(n45264) );
  NAND U45922 ( .A(n45234), .B(n45233), .Z(n45238) );
  NAND U45923 ( .A(n45236), .B(n45235), .Z(n45237) );
  AND U45924 ( .A(n45238), .B(n45237), .Z(n45246) );
  NAND U45925 ( .A(n45240), .B(n45239), .Z(n45244) );
  NAND U45926 ( .A(n45242), .B(n45241), .Z(n45243) );
  NAND U45927 ( .A(n45244), .B(n45243), .Z(n45245) );
  XNOR U45928 ( .A(n45246), .B(n45245), .Z(n45262) );
  AND U45929 ( .A(y[8129]), .B(x[510]), .Z(n45248) );
  NAND U45930 ( .A(y[8131]), .B(x[508]), .Z(n45247) );
  XNOR U45931 ( .A(n45248), .B(n45247), .Z(n45252) );
  AND U45932 ( .A(y[8130]), .B(x[509]), .Z(n45250) );
  NAND U45933 ( .A(y[8139]), .B(x[500]), .Z(n45249) );
  XNOR U45934 ( .A(n45250), .B(n45249), .Z(n45251) );
  XOR U45935 ( .A(n45252), .B(n45251), .Z(n45260) );
  AND U45936 ( .A(y[8158]), .B(x[481]), .Z(n45254) );
  NAND U45937 ( .A(y[8159]), .B(x[480]), .Z(n45253) );
  XNOR U45938 ( .A(n45254), .B(n45253), .Z(n45258) );
  AND U45939 ( .A(y[8156]), .B(x[483]), .Z(n45256) );
  NAND U45940 ( .A(y[8141]), .B(x[498]), .Z(n45255) );
  XNOR U45941 ( .A(n45256), .B(n45255), .Z(n45257) );
  XNOR U45942 ( .A(n45258), .B(n45257), .Z(n45259) );
  XNOR U45943 ( .A(n45260), .B(n45259), .Z(n45261) );
  XNOR U45944 ( .A(n45262), .B(n45261), .Z(n45263) );
  ANDN U45945 ( .B(n45270), .A(n45269), .Z(n45274) );
  ANDN U45946 ( .B(n45272), .A(n45271), .Z(n45273) );
  OR U45947 ( .A(n45274), .B(n45273), .Z(n45275) );
  NAND U45948 ( .A(n45278), .B(n45277), .Z(n45282) );
  NAND U45949 ( .A(n45280), .B(n45279), .Z(n45281) );
  AND U45950 ( .A(n45282), .B(n45281), .Z(n45290) );
  NAND U45951 ( .A(n45284), .B(n45283), .Z(n45288) );
  NAND U45952 ( .A(n45286), .B(n45285), .Z(n45287) );
  NAND U45953 ( .A(n45288), .B(n45287), .Z(n45289) );
  NAND U45954 ( .A(n45292), .B(n45291), .Z(n45296) );
  NAND U45955 ( .A(n45294), .B(n45293), .Z(n45295) );
  AND U45956 ( .A(n45296), .B(n45295), .Z(n45304) );
  NAND U45957 ( .A(n45298), .B(n45297), .Z(n45302) );
  NAND U45958 ( .A(n45300), .B(n45299), .Z(n45301) );
  NAND U45959 ( .A(n45302), .B(n45301), .Z(n45303) );
  XNOR U45960 ( .A(n45306), .B(n45305), .Z(n45307) );
  XNOR U45961 ( .A(n45308), .B(n45307), .Z(n45324) );
  NAND U45962 ( .A(n45310), .B(n45309), .Z(n45314) );
  NANDN U45963 ( .A(n45312), .B(n45311), .Z(n45313) );
  AND U45964 ( .A(n45314), .B(n45313), .Z(n45322) );
  NAND U45965 ( .A(n45318), .B(n45317), .Z(n45319) );
  NAND U45966 ( .A(n45320), .B(n45319), .Z(n45321) );
  XNOR U45967 ( .A(n45322), .B(n45321), .Z(n45323) );
  XNOR U45968 ( .A(n45324), .B(n45323), .Z(n45325) );
  XNOR U45969 ( .A(n45326), .B(n45325), .Z(n45342) );
  NANDN U45970 ( .A(n45328), .B(n45327), .Z(n45332) );
  NANDN U45971 ( .A(n45330), .B(n45329), .Z(n45331) );
  AND U45972 ( .A(n45332), .B(n45331), .Z(n45340) );
  NAND U45973 ( .A(n45334), .B(n45333), .Z(n45338) );
  NAND U45974 ( .A(n45336), .B(n45335), .Z(n45337) );
  NAND U45975 ( .A(n45338), .B(n45337), .Z(n45339) );
  XNOR U45976 ( .A(n45340), .B(n45339), .Z(n45341) );
  XNOR U45977 ( .A(n45342), .B(n45341), .Z(n45343) );
  XNOR U45978 ( .A(n45344), .B(n45343), .Z(n45360) );
  NANDN U45979 ( .A(n45346), .B(n45345), .Z(n45350) );
  NAND U45980 ( .A(n45348), .B(n45347), .Z(n45349) );
  AND U45981 ( .A(n45350), .B(n45349), .Z(n45358) );
  NANDN U45982 ( .A(n45352), .B(n45351), .Z(n45356) );
  NANDN U45983 ( .A(n45354), .B(n45353), .Z(n45355) );
  NAND U45984 ( .A(n45356), .B(n45355), .Z(n45357) );
  XNOR U45985 ( .A(n45358), .B(n45357), .Z(n45359) );
  XNOR U45986 ( .A(n45360), .B(n45359), .Z(n45361) );
  XNOR U45987 ( .A(n45362), .B(n45361), .Z(n45378) );
  NAND U45988 ( .A(n45364), .B(n45363), .Z(n45368) );
  NANDN U45989 ( .A(n45366), .B(n45365), .Z(n45367) );
  AND U45990 ( .A(n45368), .B(n45367), .Z(n45376) );
  NANDN U45991 ( .A(n45370), .B(n45369), .Z(n45374) );
  NANDN U45992 ( .A(n45372), .B(n45371), .Z(n45373) );
  NAND U45993 ( .A(n45374), .B(n45373), .Z(n45375) );
  XNOR U45994 ( .A(n45376), .B(n45375), .Z(n45377) );
  XNOR U45995 ( .A(n45378), .B(n45377), .Z(n45379) );
  XNOR U45996 ( .A(n45380), .B(n45379), .Z(n45388) );
  NAND U45997 ( .A(n45382), .B(n45381), .Z(n45386) );
  NANDN U45998 ( .A(n45384), .B(n45383), .Z(n45385) );
  NAND U45999 ( .A(n45386), .B(n45385), .Z(n45387) );
  XNOR U46000 ( .A(n45388), .B(n45387), .Z(N960) );
  AND U46001 ( .A(x[480]), .B(y[8160]), .Z(n46060) );
  XOR U46002 ( .A(n46060), .B(o[480]), .Z(N993) );
  AND U46003 ( .A(x[481]), .B(y[8160]), .Z(n45397) );
  AND U46004 ( .A(x[480]), .B(y[8161]), .Z(n45396) );
  XNOR U46005 ( .A(n45396), .B(o[481]), .Z(n45389) );
  XNOR U46006 ( .A(n45397), .B(n45389), .Z(n45391) );
  NAND U46007 ( .A(n46060), .B(o[480]), .Z(n45390) );
  XNOR U46008 ( .A(n45391), .B(n45390), .Z(N994) );
  NANDN U46009 ( .A(n45397), .B(n45389), .Z(n45393) );
  NAND U46010 ( .A(n45391), .B(n45390), .Z(n45392) );
  AND U46011 ( .A(n45393), .B(n45392), .Z(n45403) );
  AND U46012 ( .A(x[480]), .B(y[8162]), .Z(n45410) );
  XNOR U46013 ( .A(n45410), .B(o[482]), .Z(n45402) );
  XNOR U46014 ( .A(n45403), .B(n45402), .Z(n45405) );
  AND U46015 ( .A(y[8160]), .B(x[482]), .Z(n45395) );
  NAND U46016 ( .A(y[8161]), .B(x[481]), .Z(n45394) );
  XNOR U46017 ( .A(n45395), .B(n45394), .Z(n45399) );
  AND U46018 ( .A(n45396), .B(o[481]), .Z(n45398) );
  XNOR U46019 ( .A(n45399), .B(n45398), .Z(n45404) );
  XNOR U46020 ( .A(n45405), .B(n45404), .Z(N995) );
  AND U46021 ( .A(x[482]), .B(y[8161]), .Z(n45417) );
  NAND U46022 ( .A(n45417), .B(n45397), .Z(n45401) );
  NAND U46023 ( .A(n45399), .B(n45398), .Z(n45400) );
  AND U46024 ( .A(n45401), .B(n45400), .Z(n45420) );
  NANDN U46025 ( .A(n45403), .B(n45402), .Z(n45407) );
  NAND U46026 ( .A(n45405), .B(n45404), .Z(n45406) );
  AND U46027 ( .A(n45407), .B(n45406), .Z(n45419) );
  XNOR U46028 ( .A(n45420), .B(n45419), .Z(n45422) );
  AND U46029 ( .A(x[481]), .B(y[8162]), .Z(n45522) );
  XOR U46030 ( .A(n45417), .B(o[483]), .Z(n45425) );
  XOR U46031 ( .A(n45522), .B(n45425), .Z(n45427) );
  AND U46032 ( .A(y[8160]), .B(x[483]), .Z(n45409) );
  NAND U46033 ( .A(y[8163]), .B(x[480]), .Z(n45408) );
  XNOR U46034 ( .A(n45409), .B(n45408), .Z(n45412) );
  AND U46035 ( .A(n45410), .B(o[482]), .Z(n45411) );
  XOR U46036 ( .A(n45412), .B(n45411), .Z(n45426) );
  XOR U46037 ( .A(n45427), .B(n45426), .Z(n45421) );
  XOR U46038 ( .A(n45422), .B(n45421), .Z(N996) );
  AND U46039 ( .A(x[483]), .B(y[8163]), .Z(n45470) );
  NAND U46040 ( .A(n46060), .B(n45470), .Z(n45414) );
  NAND U46041 ( .A(n45412), .B(n45411), .Z(n45413) );
  NAND U46042 ( .A(n45414), .B(n45413), .Z(n45433) );
  AND U46043 ( .A(y[8164]), .B(x[480]), .Z(n45416) );
  NAND U46044 ( .A(y[8160]), .B(x[484]), .Z(n45415) );
  XNOR U46045 ( .A(n45416), .B(n45415), .Z(n45451) );
  NAND U46046 ( .A(n45417), .B(o[483]), .Z(n45452) );
  XNOR U46047 ( .A(n45451), .B(n45452), .Z(n45432) );
  AND U46048 ( .A(y[8162]), .B(x[482]), .Z(n45581) );
  NAND U46049 ( .A(y[8163]), .B(x[481]), .Z(n45418) );
  XNOR U46050 ( .A(n45581), .B(n45418), .Z(n45448) );
  AND U46051 ( .A(x[483]), .B(y[8161]), .Z(n45443) );
  XOR U46052 ( .A(o[484]), .B(n45443), .Z(n45447) );
  XOR U46053 ( .A(n45448), .B(n45447), .Z(n45431) );
  XOR U46054 ( .A(n45432), .B(n45431), .Z(n45434) );
  XOR U46055 ( .A(n45433), .B(n45434), .Z(n45438) );
  NANDN U46056 ( .A(n45420), .B(n45419), .Z(n45424) );
  NAND U46057 ( .A(n45422), .B(n45421), .Z(n45423) );
  NAND U46058 ( .A(n45424), .B(n45423), .Z(n45439) );
  NAND U46059 ( .A(n45522), .B(n45425), .Z(n45429) );
  NAND U46060 ( .A(n45427), .B(n45426), .Z(n45428) );
  NAND U46061 ( .A(n45429), .B(n45428), .Z(n45440) );
  IV U46062 ( .A(n45440), .Z(n45437) );
  XOR U46063 ( .A(n45439), .B(n45437), .Z(n45430) );
  XNOR U46064 ( .A(n45438), .B(n45430), .Z(N997) );
  NAND U46065 ( .A(n45432), .B(n45431), .Z(n45436) );
  NAND U46066 ( .A(n45434), .B(n45433), .Z(n45435) );
  AND U46067 ( .A(n45436), .B(n45435), .Z(n45478) );
  AND U46068 ( .A(y[8160]), .B(x[485]), .Z(n45442) );
  NAND U46069 ( .A(y[8165]), .B(x[480]), .Z(n45441) );
  XNOR U46070 ( .A(n45442), .B(n45441), .Z(n45463) );
  AND U46071 ( .A(o[484]), .B(n45443), .Z(n45462) );
  XOR U46072 ( .A(n45463), .B(n45462), .Z(n45461) );
  NAND U46073 ( .A(x[482]), .B(y[8163]), .Z(n45530) );
  AND U46074 ( .A(y[8162]), .B(x[483]), .Z(n45445) );
  NAND U46075 ( .A(y[8164]), .B(x[481]), .Z(n45444) );
  XNOR U46076 ( .A(n45445), .B(n45444), .Z(n45457) );
  AND U46077 ( .A(x[484]), .B(y[8161]), .Z(n45468) );
  XOR U46078 ( .A(n45468), .B(o[485]), .Z(n45456) );
  XOR U46079 ( .A(n45457), .B(n45456), .Z(n45460) );
  XOR U46080 ( .A(n45530), .B(n45460), .Z(n45446) );
  XNOR U46081 ( .A(n45461), .B(n45446), .Z(n45474) );
  NANDN U46082 ( .A(n45530), .B(n45522), .Z(n45450) );
  NAND U46083 ( .A(n45448), .B(n45447), .Z(n45449) );
  AND U46084 ( .A(n45450), .B(n45449), .Z(n45473) );
  AND U46085 ( .A(x[484]), .B(y[8164]), .Z(n46274) );
  NAND U46086 ( .A(n46274), .B(n46060), .Z(n45454) );
  NANDN U46087 ( .A(n45452), .B(n45451), .Z(n45453) );
  NAND U46088 ( .A(n45454), .B(n45453), .Z(n45472) );
  XOR U46089 ( .A(n45473), .B(n45472), .Z(n45475) );
  XNOR U46090 ( .A(n45474), .B(n45475), .Z(n45480) );
  XNOR U46091 ( .A(n45479), .B(n45480), .Z(n45455) );
  XOR U46092 ( .A(n45478), .B(n45455), .Z(N998) );
  AND U46093 ( .A(x[483]), .B(y[8164]), .Z(n45531) );
  NAND U46094 ( .A(n45531), .B(n45522), .Z(n45459) );
  NAND U46095 ( .A(n45457), .B(n45456), .Z(n45458) );
  AND U46096 ( .A(n45459), .B(n45458), .Z(n45483) );
  AND U46097 ( .A(x[485]), .B(y[8165]), .Z(n45704) );
  NAND U46098 ( .A(n46060), .B(n45704), .Z(n45465) );
  NAND U46099 ( .A(n45463), .B(n45462), .Z(n45464) );
  NAND U46100 ( .A(n45465), .B(n45464), .Z(n45492) );
  AND U46101 ( .A(y[8160]), .B(x[486]), .Z(n45467) );
  NAND U46102 ( .A(y[8166]), .B(x[480]), .Z(n45466) );
  XNOR U46103 ( .A(n45467), .B(n45466), .Z(n45498) );
  AND U46104 ( .A(n45468), .B(o[485]), .Z(n45499) );
  XOR U46105 ( .A(n45498), .B(n45499), .Z(n45491) );
  XOR U46106 ( .A(n45492), .B(n45491), .Z(n45494) );
  NAND U46107 ( .A(y[8164]), .B(x[482]), .Z(n45469) );
  XNOR U46108 ( .A(n45470), .B(n45469), .Z(n45503) );
  AND U46109 ( .A(y[8165]), .B(x[481]), .Z(n45733) );
  NAND U46110 ( .A(y[8162]), .B(x[484]), .Z(n45471) );
  XNOR U46111 ( .A(n45733), .B(n45471), .Z(n45507) );
  AND U46112 ( .A(x[485]), .B(y[8161]), .Z(n45514) );
  XOR U46113 ( .A(o[486]), .B(n45514), .Z(n45506) );
  XOR U46114 ( .A(n45507), .B(n45506), .Z(n45502) );
  XOR U46115 ( .A(n45503), .B(n45502), .Z(n45493) );
  XOR U46116 ( .A(n45494), .B(n45493), .Z(n45484) );
  XNOR U46117 ( .A(n45485), .B(n45484), .Z(n45490) );
  NANDN U46118 ( .A(n45473), .B(n45472), .Z(n45477) );
  NANDN U46119 ( .A(n45475), .B(n45474), .Z(n45476) );
  NAND U46120 ( .A(n45477), .B(n45476), .Z(n45488) );
  XOR U46121 ( .A(n45488), .B(n45489), .Z(n45481) );
  XNOR U46122 ( .A(n45490), .B(n45481), .Z(N999) );
  NANDN U46123 ( .A(n45483), .B(n45482), .Z(n45487) );
  NAND U46124 ( .A(n45485), .B(n45484), .Z(n45486) );
  NAND U46125 ( .A(n45487), .B(n45486), .Z(n45548) );
  IV U46126 ( .A(n45548), .Z(n45547) );
  NAND U46127 ( .A(n45492), .B(n45491), .Z(n45496) );
  NAND U46128 ( .A(n45494), .B(n45493), .Z(n45495) );
  AND U46129 ( .A(n45496), .B(n45495), .Z(n45557) );
  AND U46130 ( .A(y[8162]), .B(x[485]), .Z(n45617) );
  NAND U46131 ( .A(y[8166]), .B(x[481]), .Z(n45497) );
  XNOR U46132 ( .A(n45617), .B(n45497), .Z(n45524) );
  AND U46133 ( .A(x[486]), .B(y[8161]), .Z(n45527) );
  XOR U46134 ( .A(o[487]), .B(n45527), .Z(n45523) );
  XOR U46135 ( .A(n45524), .B(n45523), .Z(n45542) );
  AND U46136 ( .A(x[486]), .B(y[8166]), .Z(n45753) );
  NAND U46137 ( .A(n46060), .B(n45753), .Z(n45501) );
  NAND U46138 ( .A(n45499), .B(n45498), .Z(n45500) );
  AND U46139 ( .A(n45501), .B(n45500), .Z(n45541) );
  NANDN U46140 ( .A(n45530), .B(n45531), .Z(n45505) );
  NAND U46141 ( .A(n45503), .B(n45502), .Z(n45504) );
  NAND U46142 ( .A(n45505), .B(n45504), .Z(n45544) );
  AND U46143 ( .A(x[484]), .B(y[8165]), .Z(n46065) );
  NAND U46144 ( .A(n46065), .B(n45522), .Z(n45509) );
  NAND U46145 ( .A(n45507), .B(n45506), .Z(n45508) );
  AND U46146 ( .A(n45509), .B(n45508), .Z(n45519) );
  AND U46147 ( .A(y[8165]), .B(x[482]), .Z(n45511) );
  NAND U46148 ( .A(y[8163]), .B(x[484]), .Z(n45510) );
  XNOR U46149 ( .A(n45511), .B(n45510), .Z(n45532) );
  XNOR U46150 ( .A(n45532), .B(n45531), .Z(n45517) );
  AND U46151 ( .A(y[8160]), .B(x[487]), .Z(n45513) );
  NAND U46152 ( .A(y[8167]), .B(x[480]), .Z(n45512) );
  XNOR U46153 ( .A(n45513), .B(n45512), .Z(n45536) );
  AND U46154 ( .A(o[486]), .B(n45514), .Z(n45535) );
  XNOR U46155 ( .A(n45536), .B(n45535), .Z(n45516) );
  XOR U46156 ( .A(n45517), .B(n45516), .Z(n45518) );
  XOR U46157 ( .A(n45519), .B(n45518), .Z(n45554) );
  XOR U46158 ( .A(n45555), .B(n45554), .Z(n45556) );
  XOR U46159 ( .A(n45557), .B(n45556), .Z(n45550) );
  XNOR U46160 ( .A(n45549), .B(n45550), .Z(n45515) );
  XOR U46161 ( .A(n45547), .B(n45515), .Z(N1000) );
  NAND U46162 ( .A(n45517), .B(n45516), .Z(n45521) );
  NAND U46163 ( .A(n45519), .B(n45518), .Z(n45520) );
  AND U46164 ( .A(n45521), .B(n45520), .Z(n45594) );
  AND U46165 ( .A(x[485]), .B(y[8166]), .Z(n45695) );
  NAND U46166 ( .A(n45695), .B(n45522), .Z(n45526) );
  NAND U46167 ( .A(n45524), .B(n45523), .Z(n45525) );
  NAND U46168 ( .A(n45526), .B(n45525), .Z(n45592) );
  AND U46169 ( .A(o[487]), .B(n45527), .Z(n45572) );
  AND U46170 ( .A(y[8163]), .B(x[485]), .Z(n46149) );
  NAND U46171 ( .A(y[8167]), .B(x[481]), .Z(n45528) );
  XNOR U46172 ( .A(n46149), .B(n45528), .Z(n45573) );
  XNOR U46173 ( .A(n45572), .B(n45573), .Z(n45577) );
  NAND U46174 ( .A(x[483]), .B(y[8165]), .Z(n46382) );
  AND U46175 ( .A(x[486]), .B(y[8162]), .Z(n45529) );
  AND U46176 ( .A(y[8166]), .B(x[482]), .Z(n46502) );
  XOR U46177 ( .A(n45529), .B(n46502), .Z(n45582) );
  XOR U46178 ( .A(n46274), .B(n45582), .Z(n45576) );
  XOR U46179 ( .A(n45577), .B(n45578), .Z(n45591) );
  XOR U46180 ( .A(n45592), .B(n45591), .Z(n45593) );
  XOR U46181 ( .A(n45594), .B(n45593), .Z(n45600) );
  NANDN U46182 ( .A(n45530), .B(n46065), .Z(n45534) );
  NAND U46183 ( .A(n45532), .B(n45531), .Z(n45533) );
  NAND U46184 ( .A(n45534), .B(n45533), .Z(n45588) );
  AND U46185 ( .A(x[487]), .B(y[8167]), .Z(n45919) );
  NAND U46186 ( .A(n46060), .B(n45919), .Z(n45538) );
  NAND U46187 ( .A(n45536), .B(n45535), .Z(n45537) );
  NAND U46188 ( .A(n45538), .B(n45537), .Z(n45586) );
  AND U46189 ( .A(y[8160]), .B(x[488]), .Z(n45540) );
  NAND U46190 ( .A(y[8168]), .B(x[480]), .Z(n45539) );
  XNOR U46191 ( .A(n45540), .B(n45539), .Z(n45563) );
  AND U46192 ( .A(x[487]), .B(y[8161]), .Z(n45566) );
  XOR U46193 ( .A(o[488]), .B(n45566), .Z(n45562) );
  XOR U46194 ( .A(n45563), .B(n45562), .Z(n45585) );
  XOR U46195 ( .A(n45586), .B(n45585), .Z(n45587) );
  XNOR U46196 ( .A(n45588), .B(n45587), .Z(n45598) );
  NANDN U46197 ( .A(n45542), .B(n45541), .Z(n45546) );
  NANDN U46198 ( .A(n45544), .B(n45543), .Z(n45545) );
  NAND U46199 ( .A(n45546), .B(n45545), .Z(n45597) );
  XOR U46200 ( .A(n45598), .B(n45597), .Z(n45599) );
  XOR U46201 ( .A(n45600), .B(n45599), .Z(n45606) );
  OR U46202 ( .A(n45549), .B(n45547), .Z(n45553) );
  ANDN U46203 ( .B(n45549), .A(n45548), .Z(n45551) );
  OR U46204 ( .A(n45551), .B(n45550), .Z(n45552) );
  AND U46205 ( .A(n45553), .B(n45552), .Z(n45604) );
  NAND U46206 ( .A(n45555), .B(n45554), .Z(n45559) );
  NAND U46207 ( .A(n45557), .B(n45556), .Z(n45558) );
  NAND U46208 ( .A(n45559), .B(n45558), .Z(n45605) );
  IV U46209 ( .A(n45605), .Z(n45603) );
  XOR U46210 ( .A(n45604), .B(n45603), .Z(n45560) );
  XNOR U46211 ( .A(n45606), .B(n45560), .Z(N1001) );
  AND U46212 ( .A(x[488]), .B(y[8168]), .Z(n45561) );
  NAND U46213 ( .A(n45561), .B(n46060), .Z(n45565) );
  NAND U46214 ( .A(n45563), .B(n45562), .Z(n45564) );
  AND U46215 ( .A(n45565), .B(n45564), .Z(n45646) );
  AND U46216 ( .A(o[488]), .B(n45566), .Z(n45619) );
  AND U46217 ( .A(y[8164]), .B(x[485]), .Z(n45568) );
  NAND U46218 ( .A(y[8162]), .B(x[487]), .Z(n45567) );
  XNOR U46219 ( .A(n45568), .B(n45567), .Z(n45618) );
  XNOR U46220 ( .A(n45619), .B(n45618), .Z(n45644) );
  AND U46221 ( .A(y[8160]), .B(x[489]), .Z(n45570) );
  NAND U46222 ( .A(y[8169]), .B(x[480]), .Z(n45569) );
  XNOR U46223 ( .A(n45570), .B(n45569), .Z(n45626) );
  AND U46224 ( .A(x[488]), .B(y[8161]), .Z(n45633) );
  XOR U46225 ( .A(o[489]), .B(n45633), .Z(n45625) );
  XNOR U46226 ( .A(n45626), .B(n45625), .Z(n45643) );
  XOR U46227 ( .A(n45644), .B(n45643), .Z(n45645) );
  XNOR U46228 ( .A(n45646), .B(n45645), .Z(n45640) );
  AND U46229 ( .A(y[8163]), .B(x[486]), .Z(n45984) );
  NAND U46230 ( .A(y[8168]), .B(x[481]), .Z(n45571) );
  XNOR U46231 ( .A(n45984), .B(n45571), .Z(n45630) );
  XNOR U46232 ( .A(n46065), .B(n45630), .Z(n45650) );
  AND U46233 ( .A(x[482]), .B(y[8167]), .Z(n46251) );
  NAND U46234 ( .A(x[483]), .B(y[8166]), .Z(n45994) );
  XNOR U46235 ( .A(n46251), .B(n45994), .Z(n45649) );
  XNOR U46236 ( .A(n45650), .B(n45649), .Z(n45638) );
  NAND U46237 ( .A(x[485]), .B(y[8167]), .Z(n45833) );
  AND U46238 ( .A(x[481]), .B(y[8163]), .Z(n45629) );
  NANDN U46239 ( .A(n45833), .B(n45629), .Z(n45575) );
  NAND U46240 ( .A(n45573), .B(n45572), .Z(n45574) );
  NAND U46241 ( .A(n45575), .B(n45574), .Z(n45637) );
  XOR U46242 ( .A(n45638), .B(n45637), .Z(n45639) );
  XNOR U46243 ( .A(n45640), .B(n45639), .Z(n45613) );
  NANDN U46244 ( .A(n45576), .B(n46382), .Z(n45580) );
  NANDN U46245 ( .A(n45578), .B(n45577), .Z(n45579) );
  NAND U46246 ( .A(n45580), .B(n45579), .Z(n45611) );
  NAND U46247 ( .A(n45753), .B(n45581), .Z(n45584) );
  NAND U46248 ( .A(n46274), .B(n45582), .Z(n45583) );
  AND U46249 ( .A(n45584), .B(n45583), .Z(n45612) );
  XNOR U46250 ( .A(n45611), .B(n45612), .Z(n45614) );
  NAND U46251 ( .A(n45586), .B(n45585), .Z(n45590) );
  NAND U46252 ( .A(n45588), .B(n45587), .Z(n45589) );
  NAND U46253 ( .A(n45590), .B(n45589), .Z(n45652) );
  NAND U46254 ( .A(n45592), .B(n45591), .Z(n45596) );
  NAND U46255 ( .A(n45594), .B(n45593), .Z(n45595) );
  NAND U46256 ( .A(n45596), .B(n45595), .Z(n45651) );
  XOR U46257 ( .A(n45652), .B(n45651), .Z(n45654) );
  XOR U46258 ( .A(n45653), .B(n45654), .Z(n45659) );
  NAND U46259 ( .A(n45598), .B(n45597), .Z(n45602) );
  NANDN U46260 ( .A(n45600), .B(n45599), .Z(n45601) );
  NAND U46261 ( .A(n45602), .B(n45601), .Z(n45657) );
  NANDN U46262 ( .A(n45603), .B(n45604), .Z(n45609) );
  NOR U46263 ( .A(n45605), .B(n45604), .Z(n45607) );
  OR U46264 ( .A(n45607), .B(n45606), .Z(n45608) );
  AND U46265 ( .A(n45609), .B(n45608), .Z(n45658) );
  XOR U46266 ( .A(n45657), .B(n45658), .Z(n45610) );
  XNOR U46267 ( .A(n45659), .B(n45610), .Z(N1002) );
  NAND U46268 ( .A(n45612), .B(n45611), .Z(n45616) );
  NANDN U46269 ( .A(n45614), .B(n45613), .Z(n45615) );
  NAND U46270 ( .A(n45616), .B(n45615), .Z(n45718) );
  AND U46271 ( .A(x[487]), .B(y[8164]), .Z(n45697) );
  NAND U46272 ( .A(n45697), .B(n45617), .Z(n45621) );
  NAND U46273 ( .A(n45619), .B(n45618), .Z(n45620) );
  AND U46274 ( .A(n45621), .B(n45620), .Z(n45710) );
  AND U46275 ( .A(y[8163]), .B(x[487]), .Z(n45623) );
  NAND U46276 ( .A(y[8166]), .B(x[484]), .Z(n45622) );
  XNOR U46277 ( .A(n45623), .B(n45622), .Z(n45681) );
  AND U46278 ( .A(x[486]), .B(y[8164]), .Z(n45680) );
  XNOR U46279 ( .A(n45681), .B(n45680), .Z(n45708) );
  AND U46280 ( .A(x[488]), .B(y[8162]), .Z(n45893) );
  AND U46281 ( .A(x[489]), .B(y[8161]), .Z(n45691) );
  XOR U46282 ( .A(o[490]), .B(n45691), .Z(n45702) );
  XOR U46283 ( .A(n45893), .B(n45702), .Z(n45703) );
  XNOR U46284 ( .A(n45704), .B(n45703), .Z(n45707) );
  XOR U46285 ( .A(n45708), .B(n45707), .Z(n45709) );
  XNOR U46286 ( .A(n45710), .B(n45709), .Z(n45670) );
  AND U46287 ( .A(x[489]), .B(y[8169]), .Z(n45624) );
  NAND U46288 ( .A(n45624), .B(n46060), .Z(n45628) );
  NAND U46289 ( .A(n45626), .B(n45625), .Z(n45627) );
  NAND U46290 ( .A(n45628), .B(n45627), .Z(n45668) );
  AND U46291 ( .A(x[486]), .B(y[8168]), .Z(n45929) );
  NAND U46292 ( .A(n45929), .B(n45629), .Z(n45632) );
  NAND U46293 ( .A(n46065), .B(n45630), .Z(n45631) );
  NAND U46294 ( .A(n45632), .B(n45631), .Z(n45676) );
  AND U46295 ( .A(o[489]), .B(n45633), .Z(n45686) );
  AND U46296 ( .A(y[8160]), .B(x[490]), .Z(n45635) );
  AND U46297 ( .A(y[8170]), .B(x[480]), .Z(n45634) );
  XOR U46298 ( .A(n45635), .B(n45634), .Z(n45685) );
  XOR U46299 ( .A(n45686), .B(n45685), .Z(n45674) );
  AND U46300 ( .A(y[8167]), .B(x[483]), .Z(n46618) );
  NAND U46301 ( .A(y[8169]), .B(x[481]), .Z(n45636) );
  XNOR U46302 ( .A(n46618), .B(n45636), .Z(n45698) );
  AND U46303 ( .A(x[482]), .B(y[8168]), .Z(n45699) );
  XOR U46304 ( .A(n45698), .B(n45699), .Z(n45673) );
  XOR U46305 ( .A(n45674), .B(n45673), .Z(n45675) );
  XOR U46306 ( .A(n45676), .B(n45675), .Z(n45667) );
  XOR U46307 ( .A(n45668), .B(n45667), .Z(n45669) );
  XOR U46308 ( .A(n45670), .B(n45669), .Z(n45717) );
  NAND U46309 ( .A(n45638), .B(n45637), .Z(n45642) );
  NAND U46310 ( .A(n45640), .B(n45639), .Z(n45641) );
  AND U46311 ( .A(n45642), .B(n45641), .Z(n45664) );
  NAND U46312 ( .A(n45644), .B(n45643), .Z(n45648) );
  NAND U46313 ( .A(n45646), .B(n45645), .Z(n45647) );
  AND U46314 ( .A(n45648), .B(n45647), .Z(n45661) );
  XOR U46315 ( .A(n45661), .B(n45662), .Z(n45663) );
  XOR U46316 ( .A(n45664), .B(n45663), .Z(n45716) );
  XOR U46317 ( .A(n45718), .B(n45719), .Z(n45715) );
  NAND U46318 ( .A(n45652), .B(n45651), .Z(n45656) );
  NAND U46319 ( .A(n45654), .B(n45653), .Z(n45655) );
  NAND U46320 ( .A(n45656), .B(n45655), .Z(n45714) );
  XOR U46321 ( .A(n45714), .B(n45713), .Z(n45660) );
  XNOR U46322 ( .A(n45715), .B(n45660), .Z(N1003) );
  NAND U46323 ( .A(n45662), .B(n45661), .Z(n45666) );
  NANDN U46324 ( .A(n45664), .B(n45663), .Z(n45665) );
  AND U46325 ( .A(n45666), .B(n45665), .Z(n45788) );
  NAND U46326 ( .A(n45668), .B(n45667), .Z(n45672) );
  NAND U46327 ( .A(n45670), .B(n45669), .Z(n45671) );
  NAND U46328 ( .A(n45672), .B(n45671), .Z(n45786) );
  NAND U46329 ( .A(n45674), .B(n45673), .Z(n45678) );
  NAND U46330 ( .A(n45676), .B(n45675), .Z(n45677) );
  NAND U46331 ( .A(n45678), .B(n45677), .Z(n45774) );
  AND U46332 ( .A(x[487]), .B(y[8166]), .Z(n45828) );
  AND U46333 ( .A(x[484]), .B(y[8163]), .Z(n45679) );
  NAND U46334 ( .A(n45828), .B(n45679), .Z(n45683) );
  NAND U46335 ( .A(n45681), .B(n45680), .Z(n45682) );
  NAND U46336 ( .A(n45683), .B(n45682), .Z(n45772) );
  AND U46337 ( .A(x[490]), .B(y[8170]), .Z(n45684) );
  NAND U46338 ( .A(n45684), .B(n46060), .Z(n45688) );
  NAND U46339 ( .A(n45686), .B(n45685), .Z(n45687) );
  NAND U46340 ( .A(n45688), .B(n45687), .Z(n45768) );
  AND U46341 ( .A(y[8160]), .B(x[491]), .Z(n45690) );
  NAND U46342 ( .A(y[8171]), .B(x[480]), .Z(n45689) );
  XNOR U46343 ( .A(n45690), .B(n45689), .Z(n45744) );
  AND U46344 ( .A(o[490]), .B(n45691), .Z(n45743) );
  XOR U46345 ( .A(n45744), .B(n45743), .Z(n45767) );
  AND U46346 ( .A(y[8165]), .B(x[486]), .Z(n45693) );
  NAND U46347 ( .A(y[8170]), .B(x[481]), .Z(n45692) );
  XNOR U46348 ( .A(n45693), .B(n45692), .Z(n45735) );
  AND U46349 ( .A(x[490]), .B(y[8161]), .Z(n45754) );
  XOR U46350 ( .A(o[491]), .B(n45754), .Z(n45734) );
  XOR U46351 ( .A(n45735), .B(n45734), .Z(n45766) );
  XOR U46352 ( .A(n45767), .B(n45766), .Z(n45769) );
  XNOR U46353 ( .A(n45768), .B(n45769), .Z(n45773) );
  XOR U46354 ( .A(n45774), .B(n45775), .Z(n45757) );
  AND U46355 ( .A(x[483]), .B(y[8168]), .Z(n46751) );
  NAND U46356 ( .A(y[8169]), .B(x[482]), .Z(n45694) );
  XNOR U46357 ( .A(n45695), .B(n45694), .Z(n45730) );
  AND U46358 ( .A(x[484]), .B(y[8167]), .Z(n45729) );
  XNOR U46359 ( .A(n45730), .B(n45729), .Z(n45761) );
  XNOR U46360 ( .A(n46751), .B(n45761), .Z(n45763) );
  NAND U46361 ( .A(y[8162]), .B(x[489]), .Z(n45696) );
  XNOR U46362 ( .A(n45697), .B(n45696), .Z(n45749) );
  AND U46363 ( .A(x[488]), .B(y[8163]), .Z(n45748) );
  XNOR U46364 ( .A(n45749), .B(n45748), .Z(n45762) );
  XNOR U46365 ( .A(n45763), .B(n45762), .Z(n45726) );
  AND U46366 ( .A(x[483]), .B(y[8169]), .Z(n45824) );
  AND U46367 ( .A(x[481]), .B(y[8167]), .Z(n46055) );
  NAND U46368 ( .A(n45824), .B(n46055), .Z(n45701) );
  NAND U46369 ( .A(n45699), .B(n45698), .Z(n45700) );
  NAND U46370 ( .A(n45701), .B(n45700), .Z(n45724) );
  NAND U46371 ( .A(n45893), .B(n45702), .Z(n45706) );
  NAND U46372 ( .A(n45704), .B(n45703), .Z(n45705) );
  NAND U46373 ( .A(n45706), .B(n45705), .Z(n45723) );
  XOR U46374 ( .A(n45724), .B(n45723), .Z(n45725) );
  XNOR U46375 ( .A(n45726), .B(n45725), .Z(n45756) );
  NAND U46376 ( .A(n45708), .B(n45707), .Z(n45712) );
  NAND U46377 ( .A(n45710), .B(n45709), .Z(n45711) );
  NAND U46378 ( .A(n45712), .B(n45711), .Z(n45755) );
  XOR U46379 ( .A(n45756), .B(n45755), .Z(n45758) );
  XNOR U46380 ( .A(n45757), .B(n45758), .Z(n45785) );
  XOR U46381 ( .A(n45786), .B(n45785), .Z(n45787) );
  XOR U46382 ( .A(n45788), .B(n45787), .Z(n45781) );
  NANDN U46383 ( .A(n45717), .B(n45716), .Z(n45721) );
  NAND U46384 ( .A(n45719), .B(n45718), .Z(n45720) );
  AND U46385 ( .A(n45721), .B(n45720), .Z(n45779) );
  IV U46386 ( .A(n45779), .Z(n45778) );
  XOR U46387 ( .A(n45780), .B(n45778), .Z(n45722) );
  XNOR U46388 ( .A(n45781), .B(n45722), .Z(N1004) );
  NAND U46389 ( .A(n45724), .B(n45723), .Z(n45728) );
  NAND U46390 ( .A(n45726), .B(n45725), .Z(n45727) );
  NAND U46391 ( .A(n45728), .B(n45727), .Z(n45864) );
  AND U46392 ( .A(x[485]), .B(y[8169]), .Z(n46242) );
  NAND U46393 ( .A(n46502), .B(n46242), .Z(n45732) );
  NAND U46394 ( .A(n45730), .B(n45729), .Z(n45731) );
  AND U46395 ( .A(n45732), .B(n45731), .Z(n45812) );
  AND U46396 ( .A(x[486]), .B(y[8170]), .Z(n46072) );
  NAND U46397 ( .A(n46072), .B(n45733), .Z(n45737) );
  NAND U46398 ( .A(n45735), .B(n45734), .Z(n45736) );
  NAND U46399 ( .A(n45737), .B(n45736), .Z(n45811) );
  AND U46400 ( .A(x[489]), .B(y[8163]), .Z(n46497) );
  AND U46401 ( .A(y[8162]), .B(x[490]), .Z(n46492) );
  NAND U46402 ( .A(y[8168]), .B(x[484]), .Z(n45738) );
  XNOR U46403 ( .A(n46492), .B(n45738), .Z(n45855) );
  XOR U46404 ( .A(n46497), .B(n45855), .Z(n45834) );
  NAND U46405 ( .A(x[487]), .B(y[8165]), .Z(n45832) );
  XOR U46406 ( .A(n45833), .B(n45832), .Z(n45835) );
  AND U46407 ( .A(y[8160]), .B(x[492]), .Z(n45740) );
  NAND U46408 ( .A(y[8172]), .B(x[480]), .Z(n45739) );
  XNOR U46409 ( .A(n45740), .B(n45739), .Z(n45849) );
  AND U46410 ( .A(x[491]), .B(y[8161]), .Z(n45829) );
  XOR U46411 ( .A(o[492]), .B(n45829), .Z(n45848) );
  XOR U46412 ( .A(n45849), .B(n45848), .Z(n45818) );
  AND U46413 ( .A(y[8170]), .B(x[482]), .Z(n45742) );
  NAND U46414 ( .A(y[8164]), .B(x[488]), .Z(n45741) );
  XNOR U46415 ( .A(n45742), .B(n45741), .Z(n45823) );
  XOR U46416 ( .A(n45823), .B(n45824), .Z(n45817) );
  XOR U46417 ( .A(n45818), .B(n45817), .Z(n45820) );
  XOR U46418 ( .A(n45819), .B(n45820), .Z(n45813) );
  XOR U46419 ( .A(n45814), .B(n45813), .Z(n45863) );
  AND U46420 ( .A(x[491]), .B(y[8171]), .Z(n46874) );
  NAND U46421 ( .A(n46874), .B(n46060), .Z(n45746) );
  NAND U46422 ( .A(n45744), .B(n45743), .Z(n45745) );
  NAND U46423 ( .A(n45746), .B(n45745), .Z(n45841) );
  AND U46424 ( .A(x[487]), .B(y[8162]), .Z(n45970) );
  AND U46425 ( .A(x[489]), .B(y[8164]), .Z(n45747) );
  NAND U46426 ( .A(n45970), .B(n45747), .Z(n45751) );
  NAND U46427 ( .A(n45749), .B(n45748), .Z(n45750) );
  NAND U46428 ( .A(n45751), .B(n45750), .Z(n45839) );
  NAND U46429 ( .A(y[8171]), .B(x[481]), .Z(n45752) );
  XNOR U46430 ( .A(n45753), .B(n45752), .Z(n45845) );
  AND U46431 ( .A(o[491]), .B(n45754), .Z(n45844) );
  XOR U46432 ( .A(n45845), .B(n45844), .Z(n45838) );
  XOR U46433 ( .A(n45839), .B(n45838), .Z(n45840) );
  XOR U46434 ( .A(n45841), .B(n45840), .Z(n45862) );
  XOR U46435 ( .A(n45863), .B(n45862), .Z(n45865) );
  XNOR U46436 ( .A(n45864), .B(n45865), .Z(n45793) );
  NAND U46437 ( .A(n45756), .B(n45755), .Z(n45760) );
  NAND U46438 ( .A(n45758), .B(n45757), .Z(n45759) );
  NAND U46439 ( .A(n45760), .B(n45759), .Z(n45792) );
  XOR U46440 ( .A(n45793), .B(n45792), .Z(n45795) );
  NANDN U46441 ( .A(n46751), .B(n45761), .Z(n45765) );
  NAND U46442 ( .A(n45763), .B(n45762), .Z(n45764) );
  NAND U46443 ( .A(n45765), .B(n45764), .Z(n45805) );
  NAND U46444 ( .A(n45767), .B(n45766), .Z(n45771) );
  NAND U46445 ( .A(n45769), .B(n45768), .Z(n45770) );
  AND U46446 ( .A(n45771), .B(n45770), .Z(n45806) );
  XOR U46447 ( .A(n45805), .B(n45806), .Z(n45808) );
  NANDN U46448 ( .A(n45773), .B(n45772), .Z(n45777) );
  NANDN U46449 ( .A(n45775), .B(n45774), .Z(n45776) );
  AND U46450 ( .A(n45777), .B(n45776), .Z(n45807) );
  XOR U46451 ( .A(n45808), .B(n45807), .Z(n45794) );
  XNOR U46452 ( .A(n45795), .B(n45794), .Z(n45802) );
  OR U46453 ( .A(n45780), .B(n45778), .Z(n45784) );
  ANDN U46454 ( .B(n45780), .A(n45779), .Z(n45782) );
  OR U46455 ( .A(n45782), .B(n45781), .Z(n45783) );
  AND U46456 ( .A(n45784), .B(n45783), .Z(n45799) );
  NAND U46457 ( .A(n45786), .B(n45785), .Z(n45790) );
  NANDN U46458 ( .A(n45788), .B(n45787), .Z(n45789) );
  AND U46459 ( .A(n45790), .B(n45789), .Z(n45800) );
  IV U46460 ( .A(n45800), .Z(n45798) );
  XOR U46461 ( .A(n45799), .B(n45798), .Z(n45791) );
  XNOR U46462 ( .A(n45802), .B(n45791), .Z(N1005) );
  NAND U46463 ( .A(n45793), .B(n45792), .Z(n45797) );
  NAND U46464 ( .A(n45795), .B(n45794), .Z(n45796) );
  AND U46465 ( .A(n45797), .B(n45796), .Z(n45937) );
  NANDN U46466 ( .A(n45798), .B(n45799), .Z(n45804) );
  NOR U46467 ( .A(n45800), .B(n45799), .Z(n45801) );
  OR U46468 ( .A(n45802), .B(n45801), .Z(n45803) );
  AND U46469 ( .A(n45804), .B(n45803), .Z(n45936) );
  NAND U46470 ( .A(n45806), .B(n45805), .Z(n45810) );
  NAND U46471 ( .A(n45808), .B(n45807), .Z(n45809) );
  NAND U46472 ( .A(n45810), .B(n45809), .Z(n45941) );
  NANDN U46473 ( .A(n45812), .B(n45811), .Z(n45816) );
  NAND U46474 ( .A(n45814), .B(n45813), .Z(n45815) );
  AND U46475 ( .A(n45816), .B(n45815), .Z(n45870) );
  NAND U46476 ( .A(n45818), .B(n45817), .Z(n45822) );
  NAND U46477 ( .A(n45820), .B(n45819), .Z(n45821) );
  NAND U46478 ( .A(n45822), .B(n45821), .Z(n45877) );
  AND U46479 ( .A(y[8170]), .B(x[488]), .Z(n47161) );
  AND U46480 ( .A(x[482]), .B(y[8164]), .Z(n45980) );
  NAND U46481 ( .A(n47161), .B(n45980), .Z(n45826) );
  NAND U46482 ( .A(n45824), .B(n45823), .Z(n45825) );
  NAND U46483 ( .A(n45826), .B(n45825), .Z(n45908) );
  NAND U46484 ( .A(y[8172]), .B(x[481]), .Z(n45827) );
  XNOR U46485 ( .A(n45828), .B(n45827), .Z(n45899) );
  AND U46486 ( .A(o[492]), .B(n45829), .Z(n45898) );
  XOR U46487 ( .A(n45899), .B(n45898), .Z(n45906) );
  AND U46488 ( .A(x[486]), .B(y[8167]), .Z(n46914) );
  AND U46489 ( .A(y[8171]), .B(x[482]), .Z(n45831) );
  NAND U46490 ( .A(y[8164]), .B(x[489]), .Z(n45830) );
  XNOR U46491 ( .A(n45831), .B(n45830), .Z(n45912) );
  XOR U46492 ( .A(n46914), .B(n45912), .Z(n45905) );
  XOR U46493 ( .A(n45906), .B(n45905), .Z(n45907) );
  XOR U46494 ( .A(n45908), .B(n45907), .Z(n45876) );
  NAND U46495 ( .A(n45833), .B(n45832), .Z(n45837) );
  ANDN U46496 ( .B(n45835), .A(n45834), .Z(n45836) );
  ANDN U46497 ( .B(n45837), .A(n45836), .Z(n45875) );
  XOR U46498 ( .A(n45876), .B(n45875), .Z(n45878) );
  XOR U46499 ( .A(n45877), .B(n45878), .Z(n45869) );
  NAND U46500 ( .A(n45839), .B(n45838), .Z(n45843) );
  NAND U46501 ( .A(n45841), .B(n45840), .Z(n45842) );
  NAND U46502 ( .A(n45843), .B(n45842), .Z(n45884) );
  AND U46503 ( .A(x[486]), .B(y[8171]), .Z(n46243) );
  AND U46504 ( .A(x[481]), .B(y[8166]), .Z(n45897) );
  NAND U46505 ( .A(n46243), .B(n45897), .Z(n45847) );
  NAND U46506 ( .A(n45845), .B(n45844), .Z(n45846) );
  NAND U46507 ( .A(n45847), .B(n45846), .Z(n45890) );
  AND U46508 ( .A(x[492]), .B(y[8172]), .Z(n47167) );
  NAND U46509 ( .A(n47167), .B(n46060), .Z(n45851) );
  NAND U46510 ( .A(n45849), .B(n45848), .Z(n45850) );
  NAND U46511 ( .A(n45851), .B(n45850), .Z(n45888) );
  AND U46512 ( .A(x[490]), .B(y[8163]), .Z(n46763) );
  AND U46513 ( .A(y[8162]), .B(x[491]), .Z(n46724) );
  NAND U46514 ( .A(y[8165]), .B(x[488]), .Z(n45852) );
  XNOR U46515 ( .A(n46724), .B(n45852), .Z(n45894) );
  XOR U46516 ( .A(n46763), .B(n45894), .Z(n45887) );
  XOR U46517 ( .A(n45888), .B(n45887), .Z(n45889) );
  XOR U46518 ( .A(n45890), .B(n45889), .Z(n45882) );
  AND U46519 ( .A(x[490]), .B(y[8168]), .Z(n45854) );
  AND U46520 ( .A(x[484]), .B(y[8162]), .Z(n45853) );
  NAND U46521 ( .A(n45854), .B(n45853), .Z(n45857) );
  NAND U46522 ( .A(n45855), .B(n46497), .Z(n45856) );
  NAND U46523 ( .A(n45857), .B(n45856), .Z(n45933) );
  AND U46524 ( .A(y[8160]), .B(x[493]), .Z(n45859) );
  NAND U46525 ( .A(y[8173]), .B(x[480]), .Z(n45858) );
  XNOR U46526 ( .A(n45859), .B(n45858), .Z(n45925) );
  AND U46527 ( .A(x[492]), .B(y[8161]), .Z(n45917) );
  XOR U46528 ( .A(o[493]), .B(n45917), .Z(n45924) );
  XOR U46529 ( .A(n45925), .B(n45924), .Z(n45931) );
  AND U46530 ( .A(y[8168]), .B(x[485]), .Z(n45861) );
  NAND U46531 ( .A(y[8170]), .B(x[483]), .Z(n45860) );
  XNOR U46532 ( .A(n45861), .B(n45860), .Z(n45920) );
  AND U46533 ( .A(x[484]), .B(y[8169]), .Z(n45921) );
  XOR U46534 ( .A(n45920), .B(n45921), .Z(n45930) );
  XOR U46535 ( .A(n45931), .B(n45930), .Z(n45932) );
  XOR U46536 ( .A(n45933), .B(n45932), .Z(n45881) );
  XOR U46537 ( .A(n45882), .B(n45881), .Z(n45883) );
  XOR U46538 ( .A(n45884), .B(n45883), .Z(n45871) );
  XOR U46539 ( .A(n45872), .B(n45871), .Z(n45940) );
  NAND U46540 ( .A(n45863), .B(n45862), .Z(n45867) );
  NAND U46541 ( .A(n45865), .B(n45864), .Z(n45866) );
  AND U46542 ( .A(n45867), .B(n45866), .Z(n45939) );
  XOR U46543 ( .A(n45941), .B(n45942), .Z(n45938) );
  XNOR U46544 ( .A(n45936), .B(n45938), .Z(n45868) );
  XOR U46545 ( .A(n45937), .B(n45868), .Z(N1006) );
  NANDN U46546 ( .A(n45870), .B(n45869), .Z(n45874) );
  NAND U46547 ( .A(n45872), .B(n45871), .Z(n45873) );
  AND U46548 ( .A(n45874), .B(n45873), .Z(n46029) );
  NAND U46549 ( .A(n45876), .B(n45875), .Z(n45880) );
  NAND U46550 ( .A(n45878), .B(n45877), .Z(n45879) );
  NAND U46551 ( .A(n45880), .B(n45879), .Z(n46028) );
  NAND U46552 ( .A(n45882), .B(n45881), .Z(n45886) );
  NAND U46553 ( .A(n45884), .B(n45883), .Z(n45885) );
  NAND U46554 ( .A(n45886), .B(n45885), .Z(n45949) );
  NAND U46555 ( .A(n45888), .B(n45887), .Z(n45892) );
  NAND U46556 ( .A(n45890), .B(n45889), .Z(n45891) );
  AND U46557 ( .A(n45892), .B(n45891), .Z(n45955) );
  AND U46558 ( .A(x[491]), .B(y[8165]), .Z(n46086) );
  NAND U46559 ( .A(n46086), .B(n45893), .Z(n45896) );
  NAND U46560 ( .A(n45894), .B(n46763), .Z(n45895) );
  NAND U46561 ( .A(n45896), .B(n45895), .Z(n46010) );
  NAND U46562 ( .A(x[487]), .B(y[8172]), .Z(n46512) );
  NANDN U46563 ( .A(n46512), .B(n45897), .Z(n45901) );
  NAND U46564 ( .A(n45899), .B(n45898), .Z(n45900) );
  NAND U46565 ( .A(n45901), .B(n45900), .Z(n46009) );
  XOR U46566 ( .A(n46010), .B(n46009), .Z(n46012) );
  AND U46567 ( .A(x[484]), .B(y[8170]), .Z(n46391) );
  AND U46568 ( .A(y[8171]), .B(x[483]), .Z(n45903) );
  NAND U46569 ( .A(y[8166]), .B(x[488]), .Z(n45902) );
  XNOR U46570 ( .A(n45903), .B(n45902), .Z(n45995) );
  XOR U46571 ( .A(n46242), .B(n45995), .Z(n46004) );
  XOR U46572 ( .A(n46391), .B(n46004), .Z(n46006) );
  AND U46573 ( .A(x[489]), .B(y[8165]), .Z(n46573) );
  AND U46574 ( .A(y[8172]), .B(x[482]), .Z(n45904) );
  AND U46575 ( .A(y[8164]), .B(x[490]), .Z(n46613) );
  XOR U46576 ( .A(n45904), .B(n46613), .Z(n45981) );
  XOR U46577 ( .A(n46573), .B(n45981), .Z(n46005) );
  XOR U46578 ( .A(n46006), .B(n46005), .Z(n46011) );
  XNOR U46579 ( .A(n46012), .B(n46011), .Z(n45953) );
  NAND U46580 ( .A(n45906), .B(n45905), .Z(n45910) );
  NAND U46581 ( .A(n45908), .B(n45907), .Z(n45909) );
  AND U46582 ( .A(n45910), .B(n45909), .Z(n45952) );
  XOR U46583 ( .A(n45953), .B(n45952), .Z(n45954) );
  XNOR U46584 ( .A(n45955), .B(n45954), .Z(n45947) );
  AND U46585 ( .A(x[489]), .B(y[8171]), .Z(n45911) );
  NAND U46586 ( .A(n45911), .B(n45980), .Z(n45914) );
  NAND U46587 ( .A(n45912), .B(n46914), .Z(n45913) );
  NAND U46588 ( .A(n45914), .B(n45913), .Z(n45967) );
  AND U46589 ( .A(y[8160]), .B(x[494]), .Z(n45916) );
  NAND U46590 ( .A(y[8174]), .B(x[480]), .Z(n45915) );
  XNOR U46591 ( .A(n45916), .B(n45915), .Z(n45990) );
  AND U46592 ( .A(o[493]), .B(n45917), .Z(n45989) );
  XOR U46593 ( .A(n45990), .B(n45989), .Z(n45965) );
  NAND U46594 ( .A(y[8162]), .B(x[492]), .Z(n45918) );
  XNOR U46595 ( .A(n45919), .B(n45918), .Z(n45972) );
  AND U46596 ( .A(x[493]), .B(y[8161]), .Z(n45979) );
  XOR U46597 ( .A(o[494]), .B(n45979), .Z(n45971) );
  XOR U46598 ( .A(n45972), .B(n45971), .Z(n45964) );
  XOR U46599 ( .A(n45965), .B(n45964), .Z(n45966) );
  XNOR U46600 ( .A(n45967), .B(n45966), .Z(n46016) );
  AND U46601 ( .A(x[485]), .B(y[8170]), .Z(n46073) );
  NAND U46602 ( .A(n46751), .B(n46073), .Z(n45923) );
  NAND U46603 ( .A(n45921), .B(n45920), .Z(n45922) );
  AND U46604 ( .A(n45923), .B(n45922), .Z(n45961) );
  AND U46605 ( .A(x[493]), .B(y[8173]), .Z(n47486) );
  NAND U46606 ( .A(n47486), .B(n46060), .Z(n45927) );
  NAND U46607 ( .A(n45925), .B(n45924), .Z(n45926) );
  NAND U46608 ( .A(n45927), .B(n45926), .Z(n45959) );
  NAND U46609 ( .A(y[8163]), .B(x[491]), .Z(n45928) );
  XNOR U46610 ( .A(n45929), .B(n45928), .Z(n45985) );
  AND U46611 ( .A(x[481]), .B(y[8173]), .Z(n45986) );
  XOR U46612 ( .A(n45985), .B(n45986), .Z(n45958) );
  XOR U46613 ( .A(n45959), .B(n45958), .Z(n45960) );
  XOR U46614 ( .A(n45961), .B(n45960), .Z(n46015) );
  XOR U46615 ( .A(n46016), .B(n46015), .Z(n46018) );
  NAND U46616 ( .A(n45931), .B(n45930), .Z(n45935) );
  NAND U46617 ( .A(n45933), .B(n45932), .Z(n45934) );
  AND U46618 ( .A(n45935), .B(n45934), .Z(n46017) );
  XNOR U46619 ( .A(n46018), .B(n46017), .Z(n45946) );
  XOR U46620 ( .A(n45947), .B(n45946), .Z(n45948) );
  XOR U46621 ( .A(n45949), .B(n45948), .Z(n46030) );
  XNOR U46622 ( .A(n46031), .B(n46030), .Z(n46024) );
  NANDN U46623 ( .A(n45940), .B(n45939), .Z(n45944) );
  NAND U46624 ( .A(n45942), .B(n45941), .Z(n45943) );
  AND U46625 ( .A(n45944), .B(n45943), .Z(n46022) );
  IV U46626 ( .A(n46022), .Z(n46021) );
  XOR U46627 ( .A(n46023), .B(n46021), .Z(n45945) );
  XNOR U46628 ( .A(n46024), .B(n45945), .Z(N1007) );
  NAND U46629 ( .A(n45947), .B(n45946), .Z(n45951) );
  NAND U46630 ( .A(n45949), .B(n45948), .Z(n45950) );
  AND U46631 ( .A(n45951), .B(n45950), .Z(n46127) );
  NAND U46632 ( .A(n45953), .B(n45952), .Z(n45957) );
  NAND U46633 ( .A(n45955), .B(n45954), .Z(n45956) );
  NAND U46634 ( .A(n45957), .B(n45956), .Z(n46096) );
  NAND U46635 ( .A(n45959), .B(n45958), .Z(n45963) );
  NANDN U46636 ( .A(n45961), .B(n45960), .Z(n45962) );
  NAND U46637 ( .A(n45963), .B(n45962), .Z(n46102) );
  NAND U46638 ( .A(n45965), .B(n45964), .Z(n45969) );
  NAND U46639 ( .A(n45967), .B(n45966), .Z(n45968) );
  NAND U46640 ( .A(n45969), .B(n45968), .Z(n46100) );
  NAND U46641 ( .A(x[492]), .B(y[8167]), .Z(n46504) );
  NANDN U46642 ( .A(n46504), .B(n45970), .Z(n45974) );
  NAND U46643 ( .A(n45972), .B(n45971), .Z(n45973) );
  AND U46644 ( .A(n45974), .B(n45973), .Z(n46038) );
  AND U46645 ( .A(y[8164]), .B(x[491]), .Z(n45976) );
  NAND U46646 ( .A(y[8162]), .B(x[493]), .Z(n45975) );
  XNOR U46647 ( .A(n45976), .B(n45975), .Z(n46042) );
  AND U46648 ( .A(x[492]), .B(y[8163]), .Z(n46041) );
  XNOR U46649 ( .A(n46042), .B(n46041), .Z(n46036) );
  AND U46650 ( .A(y[8160]), .B(x[495]), .Z(n45978) );
  NAND U46651 ( .A(y[8175]), .B(x[480]), .Z(n45977) );
  XNOR U46652 ( .A(n45978), .B(n45977), .Z(n46062) );
  AND U46653 ( .A(o[494]), .B(n45979), .Z(n46061) );
  XNOR U46654 ( .A(n46062), .B(n46061), .Z(n46035) );
  XOR U46655 ( .A(n46036), .B(n46035), .Z(n46037) );
  XNOR U46656 ( .A(n46038), .B(n46037), .Z(n46108) );
  NAND U46657 ( .A(x[490]), .B(y[8172]), .Z(n46916) );
  NANDN U46658 ( .A(n46916), .B(n45980), .Z(n45983) );
  NAND U46659 ( .A(n46573), .B(n45981), .Z(n45982) );
  NAND U46660 ( .A(n45983), .B(n45982), .Z(n46106) );
  AND U46661 ( .A(x[491]), .B(y[8168]), .Z(n46390) );
  NAND U46662 ( .A(n46390), .B(n45984), .Z(n45988) );
  NAND U46663 ( .A(n45986), .B(n45985), .Z(n45987) );
  NAND U46664 ( .A(n45988), .B(n45987), .Z(n46105) );
  XOR U46665 ( .A(n46106), .B(n46105), .Z(n46107) );
  XOR U46666 ( .A(n46108), .B(n46107), .Z(n46099) );
  XOR U46667 ( .A(n46100), .B(n46099), .Z(n46101) );
  XNOR U46668 ( .A(n46102), .B(n46101), .Z(n46093) );
  AND U46669 ( .A(x[494]), .B(y[8174]), .Z(n47739) );
  NAND U46670 ( .A(n47739), .B(n46060), .Z(n45992) );
  NAND U46671 ( .A(n45990), .B(n45989), .Z(n45991) );
  NAND U46672 ( .A(n45992), .B(n45991), .Z(n46088) );
  AND U46673 ( .A(x[488]), .B(y[8171]), .Z(n45993) );
  NANDN U46674 ( .A(n45994), .B(n45993), .Z(n45997) );
  NAND U46675 ( .A(n45995), .B(n46242), .Z(n45996) );
  NAND U46676 ( .A(n45997), .B(n45996), .Z(n46087) );
  XOR U46677 ( .A(n46088), .B(n46087), .Z(n46090) );
  AND U46678 ( .A(y[8165]), .B(x[490]), .Z(n45999) );
  NAND U46679 ( .A(y[8171]), .B(x[484]), .Z(n45998) );
  XNOR U46680 ( .A(n45999), .B(n45998), .Z(n46068) );
  AND U46681 ( .A(x[487]), .B(y[8168]), .Z(n46067) );
  XNOR U46682 ( .A(n46068), .B(n46067), .Z(n46075) );
  NAND U46683 ( .A(x[486]), .B(y[8169]), .Z(n46158) );
  XNOR U46684 ( .A(n46158), .B(n46073), .Z(n46074) );
  XNOR U46685 ( .A(n46075), .B(n46074), .Z(n46051) );
  AND U46686 ( .A(y[8173]), .B(x[482]), .Z(n46001) );
  NAND U46687 ( .A(y[8166]), .B(x[489]), .Z(n46000) );
  XNOR U46688 ( .A(n46001), .B(n46000), .Z(n46078) );
  AND U46689 ( .A(x[483]), .B(y[8172]), .Z(n46079) );
  XOR U46690 ( .A(n46078), .B(n46079), .Z(n46050) );
  AND U46691 ( .A(y[8174]), .B(x[481]), .Z(n46003) );
  NAND U46692 ( .A(y[8167]), .B(x[488]), .Z(n46002) );
  XNOR U46693 ( .A(n46003), .B(n46002), .Z(n46057) );
  AND U46694 ( .A(x[494]), .B(y[8161]), .Z(n46084) );
  XOR U46695 ( .A(o[495]), .B(n46084), .Z(n46056) );
  XOR U46696 ( .A(n46057), .B(n46056), .Z(n46049) );
  XOR U46697 ( .A(n46050), .B(n46049), .Z(n46052) );
  XOR U46698 ( .A(n46051), .B(n46052), .Z(n46089) );
  XNOR U46699 ( .A(n46090), .B(n46089), .Z(n46112) );
  NAND U46700 ( .A(n46391), .B(n46004), .Z(n46008) );
  NAND U46701 ( .A(n46006), .B(n46005), .Z(n46007) );
  AND U46702 ( .A(n46008), .B(n46007), .Z(n46111) );
  XOR U46703 ( .A(n46112), .B(n46111), .Z(n46113) );
  NAND U46704 ( .A(n46010), .B(n46009), .Z(n46014) );
  NAND U46705 ( .A(n46012), .B(n46011), .Z(n46013) );
  AND U46706 ( .A(n46014), .B(n46013), .Z(n46114) );
  XOR U46707 ( .A(n46113), .B(n46114), .Z(n46094) );
  XOR U46708 ( .A(n46093), .B(n46094), .Z(n46095) );
  XNOR U46709 ( .A(n46096), .B(n46095), .Z(n46124) );
  NAND U46710 ( .A(n46016), .B(n46015), .Z(n46020) );
  NAND U46711 ( .A(n46018), .B(n46017), .Z(n46019) );
  AND U46712 ( .A(n46020), .B(n46019), .Z(n46125) );
  XOR U46713 ( .A(n46124), .B(n46125), .Z(n46126) );
  XOR U46714 ( .A(n46127), .B(n46126), .Z(n46120) );
  OR U46715 ( .A(n46023), .B(n46021), .Z(n46027) );
  ANDN U46716 ( .B(n46023), .A(n46022), .Z(n46025) );
  OR U46717 ( .A(n46025), .B(n46024), .Z(n46026) );
  AND U46718 ( .A(n46027), .B(n46026), .Z(n46119) );
  NANDN U46719 ( .A(n46029), .B(n46028), .Z(n46033) );
  NAND U46720 ( .A(n46031), .B(n46030), .Z(n46032) );
  NAND U46721 ( .A(n46033), .B(n46032), .Z(n46118) );
  IV U46722 ( .A(n46118), .Z(n46117) );
  XOR U46723 ( .A(n46119), .B(n46117), .Z(n46034) );
  XNOR U46724 ( .A(n46120), .B(n46034), .Z(N1008) );
  NAND U46725 ( .A(n46036), .B(n46035), .Z(n46040) );
  NAND U46726 ( .A(n46038), .B(n46037), .Z(n46039) );
  NAND U46727 ( .A(n46040), .B(n46039), .Z(n46213) );
  AND U46728 ( .A(x[493]), .B(y[8164]), .Z(n46209) );
  NAND U46729 ( .A(n46724), .B(n46209), .Z(n46044) );
  NAND U46730 ( .A(n46042), .B(n46041), .Z(n46043) );
  NAND U46731 ( .A(n46044), .B(n46043), .Z(n46196) );
  AND U46732 ( .A(y[8174]), .B(x[482]), .Z(n46046) );
  NAND U46733 ( .A(y[8167]), .B(x[489]), .Z(n46045) );
  XNOR U46734 ( .A(n46046), .B(n46045), .Z(n46203) );
  NAND U46735 ( .A(x[483]), .B(y[8173]), .Z(n46204) );
  XNOR U46736 ( .A(n46203), .B(n46204), .Z(n46194) );
  AND U46737 ( .A(x[492]), .B(y[8164]), .Z(n46885) );
  AND U46738 ( .A(y[8171]), .B(x[485]), .Z(n46048) );
  NAND U46739 ( .A(y[8163]), .B(x[493]), .Z(n46047) );
  XNOR U46740 ( .A(n46048), .B(n46047), .Z(n46150) );
  XOR U46741 ( .A(n46885), .B(n46150), .Z(n46193) );
  XOR U46742 ( .A(n46194), .B(n46193), .Z(n46195) );
  XNOR U46743 ( .A(n46196), .B(n46195), .Z(n46210) );
  NAND U46744 ( .A(n46050), .B(n46049), .Z(n46054) );
  NAND U46745 ( .A(n46052), .B(n46051), .Z(n46053) );
  AND U46746 ( .A(n46054), .B(n46053), .Z(n46211) );
  XOR U46747 ( .A(n46210), .B(n46211), .Z(n46212) );
  XOR U46748 ( .A(n46213), .B(n46212), .Z(n46184) );
  AND U46749 ( .A(x[488]), .B(y[8174]), .Z(n46392) );
  NAND U46750 ( .A(n46392), .B(n46055), .Z(n46059) );
  NAND U46751 ( .A(n46057), .B(n46056), .Z(n46058) );
  AND U46752 ( .A(n46059), .B(n46058), .Z(n46188) );
  AND U46753 ( .A(x[495]), .B(y[8175]), .Z(n48167) );
  NAND U46754 ( .A(n48167), .B(n46060), .Z(n46064) );
  NAND U46755 ( .A(n46062), .B(n46061), .Z(n46063) );
  NAND U46756 ( .A(n46064), .B(n46063), .Z(n46187) );
  AND U46757 ( .A(x[490]), .B(y[8171]), .Z(n46066) );
  NAND U46758 ( .A(n46066), .B(n46065), .Z(n46070) );
  NAND U46759 ( .A(n46068), .B(n46067), .Z(n46069) );
  NAND U46760 ( .A(n46070), .B(n46069), .Z(n46145) );
  AND U46761 ( .A(x[480]), .B(y[8176]), .Z(n46167) );
  NAND U46762 ( .A(x[496]), .B(y[8160]), .Z(n46168) );
  NAND U46763 ( .A(x[495]), .B(y[8161]), .Z(n46155) );
  XOR U46764 ( .A(o[496]), .B(n46155), .Z(n46170) );
  NAND U46765 ( .A(y[8169]), .B(x[487]), .Z(n46071) );
  XNOR U46766 ( .A(n46072), .B(n46071), .Z(n46160) );
  AND U46767 ( .A(x[490]), .B(y[8166]), .Z(n46159) );
  XOR U46768 ( .A(n46160), .B(n46159), .Z(n46143) );
  XOR U46769 ( .A(n46144), .B(n46143), .Z(n46146) );
  XOR U46770 ( .A(n46145), .B(n46146), .Z(n46189) );
  XNOR U46771 ( .A(n46190), .B(n46189), .Z(n46140) );
  NANDN U46772 ( .A(n46073), .B(n46158), .Z(n46077) );
  NAND U46773 ( .A(n46075), .B(n46074), .Z(n46076) );
  NAND U46774 ( .A(n46077), .B(n46076), .Z(n46138) );
  NAND U46775 ( .A(x[489]), .B(y[8173]), .Z(n46897) );
  NANDN U46776 ( .A(n46897), .B(n46502), .Z(n46081) );
  NAND U46777 ( .A(n46079), .B(n46078), .Z(n46080) );
  AND U46778 ( .A(n46081), .B(n46080), .Z(n46178) );
  AND U46779 ( .A(y[8175]), .B(x[481]), .Z(n46083) );
  NAND U46780 ( .A(y[8168]), .B(x[488]), .Z(n46082) );
  XNOR U46781 ( .A(n46083), .B(n46082), .Z(n46164) );
  AND U46782 ( .A(o[495]), .B(n46084), .Z(n46163) );
  XOR U46783 ( .A(n46164), .B(n46163), .Z(n46175) );
  NAND U46784 ( .A(y[8162]), .B(x[494]), .Z(n46085) );
  XNOR U46785 ( .A(n46086), .B(n46085), .Z(n46199) );
  NAND U46786 ( .A(x[484]), .B(y[8172]), .Z(n46200) );
  XNOR U46787 ( .A(n46199), .B(n46200), .Z(n46176) );
  XOR U46788 ( .A(n46175), .B(n46176), .Z(n46177) );
  XOR U46789 ( .A(n46178), .B(n46177), .Z(n46137) );
  XOR U46790 ( .A(n46138), .B(n46137), .Z(n46139) );
  XOR U46791 ( .A(n46140), .B(n46139), .Z(n46181) );
  NAND U46792 ( .A(n46088), .B(n46087), .Z(n46092) );
  NAND U46793 ( .A(n46090), .B(n46089), .Z(n46091) );
  AND U46794 ( .A(n46092), .B(n46091), .Z(n46182) );
  XOR U46795 ( .A(n46181), .B(n46182), .Z(n46183) );
  XNOR U46796 ( .A(n46184), .B(n46183), .Z(n46217) );
  NAND U46797 ( .A(n46094), .B(n46093), .Z(n46098) );
  NAND U46798 ( .A(n46096), .B(n46095), .Z(n46097) );
  AND U46799 ( .A(n46098), .B(n46097), .Z(n46216) );
  XOR U46800 ( .A(n46217), .B(n46216), .Z(n46219) );
  NAND U46801 ( .A(n46100), .B(n46099), .Z(n46104) );
  NAND U46802 ( .A(n46102), .B(n46101), .Z(n46103) );
  NAND U46803 ( .A(n46104), .B(n46103), .Z(n46134) );
  NAND U46804 ( .A(n46106), .B(n46105), .Z(n46110) );
  NAND U46805 ( .A(n46108), .B(n46107), .Z(n46109) );
  NAND U46806 ( .A(n46110), .B(n46109), .Z(n46132) );
  NAND U46807 ( .A(n46112), .B(n46111), .Z(n46116) );
  NAND U46808 ( .A(n46114), .B(n46113), .Z(n46115) );
  AND U46809 ( .A(n46116), .B(n46115), .Z(n46131) );
  XOR U46810 ( .A(n46132), .B(n46131), .Z(n46133) );
  XOR U46811 ( .A(n46134), .B(n46133), .Z(n46218) );
  XOR U46812 ( .A(n46219), .B(n46218), .Z(n46225) );
  OR U46813 ( .A(n46119), .B(n46117), .Z(n46123) );
  ANDN U46814 ( .B(n46119), .A(n46118), .Z(n46121) );
  OR U46815 ( .A(n46121), .B(n46120), .Z(n46122) );
  AND U46816 ( .A(n46123), .B(n46122), .Z(n46223) );
  NAND U46817 ( .A(n46125), .B(n46124), .Z(n46129) );
  NANDN U46818 ( .A(n46127), .B(n46126), .Z(n46128) );
  AND U46819 ( .A(n46129), .B(n46128), .Z(n46224) );
  IV U46820 ( .A(n46224), .Z(n46222) );
  XOR U46821 ( .A(n46223), .B(n46222), .Z(n46130) );
  XNOR U46822 ( .A(n46225), .B(n46130), .Z(N1009) );
  NAND U46823 ( .A(n46132), .B(n46131), .Z(n46136) );
  NAND U46824 ( .A(n46134), .B(n46133), .Z(n46135) );
  AND U46825 ( .A(n46136), .B(n46135), .Z(n46330) );
  NAND U46826 ( .A(n46138), .B(n46137), .Z(n46142) );
  NAND U46827 ( .A(n46140), .B(n46139), .Z(n46141) );
  NAND U46828 ( .A(n46142), .B(n46141), .Z(n46239) );
  NAND U46829 ( .A(n46144), .B(n46143), .Z(n46148) );
  NAND U46830 ( .A(n46146), .B(n46145), .Z(n46147) );
  AND U46831 ( .A(n46148), .B(n46147), .Z(n46321) );
  AND U46832 ( .A(x[493]), .B(y[8171]), .Z(n47175) );
  NAND U46833 ( .A(n47175), .B(n46149), .Z(n46152) );
  NAND U46834 ( .A(n46150), .B(n46885), .Z(n46151) );
  AND U46835 ( .A(n46152), .B(n46151), .Z(n46297) );
  AND U46836 ( .A(y[8176]), .B(x[481]), .Z(n46154) );
  NAND U46837 ( .A(y[8168]), .B(x[489]), .Z(n46153) );
  XNOR U46838 ( .A(n46154), .B(n46153), .Z(n46247) );
  NANDN U46839 ( .A(n46155), .B(o[496]), .Z(n46248) );
  XNOR U46840 ( .A(n46247), .B(n46248), .Z(n46295) );
  AND U46841 ( .A(y[8162]), .B(x[495]), .Z(n46157) );
  NAND U46842 ( .A(y[8165]), .B(x[492]), .Z(n46156) );
  XNOR U46843 ( .A(n46157), .B(n46156), .Z(n46271) );
  AND U46844 ( .A(x[494]), .B(y[8163]), .Z(n46270) );
  XOR U46845 ( .A(n46271), .B(n46270), .Z(n46294) );
  XOR U46846 ( .A(n46295), .B(n46294), .Z(n46296) );
  AND U46847 ( .A(x[487]), .B(y[8170]), .Z(n46259) );
  NANDN U46848 ( .A(n46158), .B(n46259), .Z(n46162) );
  NAND U46849 ( .A(n46160), .B(n46159), .Z(n46161) );
  AND U46850 ( .A(n46162), .B(n46161), .Z(n46307) );
  NAND U46851 ( .A(x[488]), .B(y[8175]), .Z(n46975) );
  AND U46852 ( .A(x[481]), .B(y[8168]), .Z(n46370) );
  NANDN U46853 ( .A(n46975), .B(n46370), .Z(n46166) );
  NAND U46854 ( .A(n46164), .B(n46163), .Z(n46165) );
  NAND U46855 ( .A(n46166), .B(n46165), .Z(n46306) );
  NANDN U46856 ( .A(n46168), .B(n46167), .Z(n46172) );
  NANDN U46857 ( .A(n46170), .B(n46169), .Z(n46171) );
  AND U46858 ( .A(n46172), .B(n46171), .Z(n46303) );
  AND U46859 ( .A(x[480]), .B(y[8177]), .Z(n46285) );
  AND U46860 ( .A(x[497]), .B(y[8160]), .Z(n46284) );
  XOR U46861 ( .A(n46285), .B(n46284), .Z(n46287) );
  AND U46862 ( .A(x[496]), .B(y[8161]), .Z(n46281) );
  XOR U46863 ( .A(n46281), .B(o[497]), .Z(n46286) );
  XOR U46864 ( .A(n46287), .B(n46286), .Z(n46300) );
  AND U46865 ( .A(y[8175]), .B(x[482]), .Z(n46174) );
  NAND U46866 ( .A(y[8167]), .B(x[490]), .Z(n46173) );
  XNOR U46867 ( .A(n46174), .B(n46173), .Z(n46252) );
  NAND U46868 ( .A(x[483]), .B(y[8174]), .Z(n46253) );
  XOR U46869 ( .A(n46252), .B(n46253), .Z(n46301) );
  XOR U46870 ( .A(n46309), .B(n46308), .Z(n46318) );
  XOR U46871 ( .A(n46319), .B(n46318), .Z(n46320) );
  NAND U46872 ( .A(n46176), .B(n46175), .Z(n46180) );
  NANDN U46873 ( .A(n46178), .B(n46177), .Z(n46179) );
  AND U46874 ( .A(n46180), .B(n46179), .Z(n46237) );
  XOR U46875 ( .A(n46236), .B(n46237), .Z(n46238) );
  XNOR U46876 ( .A(n46239), .B(n46238), .Z(n46328) );
  NAND U46877 ( .A(n46182), .B(n46181), .Z(n46186) );
  NAND U46878 ( .A(n46184), .B(n46183), .Z(n46185) );
  AND U46879 ( .A(n46186), .B(n46185), .Z(n46233) );
  NANDN U46880 ( .A(n46188), .B(n46187), .Z(n46192) );
  NAND U46881 ( .A(n46190), .B(n46189), .Z(n46191) );
  NAND U46882 ( .A(n46192), .B(n46191), .Z(n46315) );
  NAND U46883 ( .A(n46194), .B(n46193), .Z(n46198) );
  NAND U46884 ( .A(n46196), .B(n46195), .Z(n46197) );
  NAND U46885 ( .A(n46198), .B(n46197), .Z(n46313) );
  NAND U46886 ( .A(x[494]), .B(y[8165]), .Z(n46489) );
  NANDN U46887 ( .A(n46489), .B(n46724), .Z(n46202) );
  NANDN U46888 ( .A(n46200), .B(n46199), .Z(n46201) );
  AND U46889 ( .A(n46202), .B(n46201), .Z(n46265) );
  AND U46890 ( .A(x[489]), .B(y[8174]), .Z(n47156) );
  NAND U46891 ( .A(n46251), .B(n47156), .Z(n46206) );
  NANDN U46892 ( .A(n46204), .B(n46203), .Z(n46205) );
  NAND U46893 ( .A(n46206), .B(n46205), .Z(n46264) );
  XNOR U46894 ( .A(n46265), .B(n46264), .Z(n46266) );
  AND U46895 ( .A(x[485]), .B(y[8172]), .Z(n46352) );
  NAND U46896 ( .A(y[8169]), .B(x[488]), .Z(n46207) );
  XNOR U46897 ( .A(n46352), .B(n46207), .Z(n46244) );
  XOR U46898 ( .A(n46244), .B(n46243), .Z(n46258) );
  XOR U46899 ( .A(n46258), .B(n46259), .Z(n46260) );
  NAND U46900 ( .A(y[8173]), .B(x[484]), .Z(n46208) );
  XNOR U46901 ( .A(n46209), .B(n46208), .Z(n46275) );
  NAND U46902 ( .A(x[491]), .B(y[8166]), .Z(n46276) );
  XOR U46903 ( .A(n46275), .B(n46276), .Z(n46261) );
  XOR U46904 ( .A(n46260), .B(n46261), .Z(n46267) );
  XNOR U46905 ( .A(n46266), .B(n46267), .Z(n46312) );
  XOR U46906 ( .A(n46313), .B(n46312), .Z(n46314) );
  XNOR U46907 ( .A(n46315), .B(n46314), .Z(n46231) );
  NAND U46908 ( .A(n46211), .B(n46210), .Z(n46215) );
  NAND U46909 ( .A(n46213), .B(n46212), .Z(n46214) );
  NAND U46910 ( .A(n46215), .B(n46214), .Z(n46230) );
  XOR U46911 ( .A(n46231), .B(n46230), .Z(n46232) );
  XOR U46912 ( .A(n46233), .B(n46232), .Z(n46327) );
  XOR U46913 ( .A(n46328), .B(n46327), .Z(n46329) );
  XOR U46914 ( .A(n46330), .B(n46329), .Z(n46326) );
  NAND U46915 ( .A(n46217), .B(n46216), .Z(n46221) );
  NAND U46916 ( .A(n46219), .B(n46218), .Z(n46220) );
  NAND U46917 ( .A(n46221), .B(n46220), .Z(n46325) );
  NANDN U46918 ( .A(n46222), .B(n46223), .Z(n46228) );
  NOR U46919 ( .A(n46224), .B(n46223), .Z(n46226) );
  OR U46920 ( .A(n46226), .B(n46225), .Z(n46227) );
  AND U46921 ( .A(n46228), .B(n46227), .Z(n46324) );
  XOR U46922 ( .A(n46325), .B(n46324), .Z(n46229) );
  XNOR U46923 ( .A(n46326), .B(n46229), .Z(N1010) );
  NAND U46924 ( .A(n46231), .B(n46230), .Z(n46235) );
  NANDN U46925 ( .A(n46233), .B(n46232), .Z(n46234) );
  AND U46926 ( .A(n46235), .B(n46234), .Z(n46439) );
  NAND U46927 ( .A(n46237), .B(n46236), .Z(n46241) );
  NAND U46928 ( .A(n46239), .B(n46238), .Z(n46240) );
  AND U46929 ( .A(n46241), .B(n46240), .Z(n46437) );
  AND U46930 ( .A(x[488]), .B(y[8172]), .Z(n46619) );
  NAND U46931 ( .A(n46619), .B(n46242), .Z(n46246) );
  NAND U46932 ( .A(n46244), .B(n46243), .Z(n46245) );
  NAND U46933 ( .A(n46246), .B(n46245), .Z(n46425) );
  AND U46934 ( .A(x[489]), .B(y[8176]), .Z(n47252) );
  NAND U46935 ( .A(n47252), .B(n46370), .Z(n46250) );
  NANDN U46936 ( .A(n46248), .B(n46247), .Z(n46249) );
  NAND U46937 ( .A(n46250), .B(n46249), .Z(n46424) );
  XOR U46938 ( .A(n46425), .B(n46424), .Z(n46427) );
  NAND U46939 ( .A(x[490]), .B(y[8175]), .Z(n47251) );
  NANDN U46940 ( .A(n47251), .B(n46251), .Z(n46255) );
  NANDN U46941 ( .A(n46253), .B(n46252), .Z(n46254) );
  AND U46942 ( .A(n46255), .B(n46254), .Z(n46403) );
  AND U46943 ( .A(x[480]), .B(y[8178]), .Z(n46375) );
  NAND U46944 ( .A(x[498]), .B(y[8160]), .Z(n46376) );
  XNOR U46945 ( .A(n46375), .B(n46376), .Z(n46377) );
  NAND U46946 ( .A(x[497]), .B(y[8161]), .Z(n46397) );
  XOR U46947 ( .A(o[498]), .B(n46397), .Z(n46378) );
  XNOR U46948 ( .A(n46377), .B(n46378), .Z(n46400) );
  AND U46949 ( .A(y[8165]), .B(x[493]), .Z(n46257) );
  NAND U46950 ( .A(y[8175]), .B(x[483]), .Z(n46256) );
  XNOR U46951 ( .A(n46257), .B(n46256), .Z(n46383) );
  NAND U46952 ( .A(x[492]), .B(y[8166]), .Z(n46384) );
  XOR U46953 ( .A(n46383), .B(n46384), .Z(n46401) );
  XNOR U46954 ( .A(n46400), .B(n46401), .Z(n46402) );
  XNOR U46955 ( .A(n46403), .B(n46402), .Z(n46426) );
  XOR U46956 ( .A(n46427), .B(n46426), .Z(n46347) );
  NAND U46957 ( .A(n46259), .B(n46258), .Z(n46263) );
  NANDN U46958 ( .A(n46261), .B(n46260), .Z(n46262) );
  AND U46959 ( .A(n46263), .B(n46262), .Z(n46346) );
  XNOR U46960 ( .A(n46347), .B(n46346), .Z(n46348) );
  NANDN U46961 ( .A(n46265), .B(n46264), .Z(n46269) );
  NANDN U46962 ( .A(n46267), .B(n46266), .Z(n46268) );
  NAND U46963 ( .A(n46269), .B(n46268), .Z(n46349) );
  XNOR U46964 ( .A(n46348), .B(n46349), .Z(n46343) );
  AND U46965 ( .A(x[495]), .B(y[8165]), .Z(n46510) );
  AND U46966 ( .A(x[492]), .B(y[8162]), .Z(n46579) );
  NAND U46967 ( .A(n46510), .B(n46579), .Z(n46273) );
  NAND U46968 ( .A(n46271), .B(n46270), .Z(n46272) );
  NAND U46969 ( .A(n46273), .B(n46272), .Z(n46418) );
  NAND U46970 ( .A(n47486), .B(n46274), .Z(n46278) );
  NANDN U46971 ( .A(n46276), .B(n46275), .Z(n46277) );
  AND U46972 ( .A(n46278), .B(n46277), .Z(n46409) );
  AND U46973 ( .A(y[8177]), .B(x[481]), .Z(n46280) );
  NAND U46974 ( .A(y[8168]), .B(x[490]), .Z(n46279) );
  XNOR U46975 ( .A(n46280), .B(n46279), .Z(n46371) );
  NAND U46976 ( .A(n46281), .B(o[497]), .Z(n46372) );
  XNOR U46977 ( .A(n46371), .B(n46372), .Z(n46406) );
  AND U46978 ( .A(y[8163]), .B(x[495]), .Z(n46283) );
  NAND U46979 ( .A(y[8169]), .B(x[489]), .Z(n46282) );
  XNOR U46980 ( .A(n46283), .B(n46282), .Z(n46362) );
  NAND U46981 ( .A(x[494]), .B(y[8164]), .Z(n46363) );
  XOR U46982 ( .A(n46362), .B(n46363), .Z(n46407) );
  XNOR U46983 ( .A(n46406), .B(n46407), .Z(n46408) );
  XNOR U46984 ( .A(n46409), .B(n46408), .Z(n46419) );
  XOR U46985 ( .A(n46418), .B(n46419), .Z(n46421) );
  NAND U46986 ( .A(n46285), .B(n46284), .Z(n46289) );
  NAND U46987 ( .A(n46287), .B(n46286), .Z(n46288) );
  NAND U46988 ( .A(n46289), .B(n46288), .Z(n46430) );
  AND U46989 ( .A(y[8162]), .B(x[496]), .Z(n46291) );
  NAND U46990 ( .A(y[8167]), .B(x[491]), .Z(n46290) );
  XNOR U46991 ( .A(n46291), .B(n46290), .Z(n46358) );
  NAND U46992 ( .A(x[482]), .B(y[8176]), .Z(n46359) );
  XNOR U46993 ( .A(n46358), .B(n46359), .Z(n46431) );
  XOR U46994 ( .A(n46430), .B(n46431), .Z(n46433) );
  AND U46995 ( .A(y[8173]), .B(x[485]), .Z(n46471) );
  NAND U46996 ( .A(y[8172]), .B(x[486]), .Z(n46292) );
  XNOR U46997 ( .A(n46471), .B(n46292), .Z(n46355) );
  NAND U46998 ( .A(y[8174]), .B(x[484]), .Z(n46293) );
  XNOR U46999 ( .A(n47161), .B(n46293), .Z(n46393) );
  AND U47000 ( .A(x[487]), .B(y[8171]), .Z(n46394) );
  XOR U47001 ( .A(n46393), .B(n46394), .Z(n46354) );
  XOR U47002 ( .A(n46355), .B(n46354), .Z(n46432) );
  XOR U47003 ( .A(n46433), .B(n46432), .Z(n46420) );
  XOR U47004 ( .A(n46421), .B(n46420), .Z(n46341) );
  NAND U47005 ( .A(n46295), .B(n46294), .Z(n46299) );
  NANDN U47006 ( .A(n46297), .B(n46296), .Z(n46298) );
  AND U47007 ( .A(n46299), .B(n46298), .Z(n46413) );
  NANDN U47008 ( .A(n46301), .B(n46300), .Z(n46305) );
  NANDN U47009 ( .A(n46303), .B(n46302), .Z(n46304) );
  AND U47010 ( .A(n46305), .B(n46304), .Z(n46412) );
  XOR U47011 ( .A(n46413), .B(n46412), .Z(n46415) );
  NANDN U47012 ( .A(n46307), .B(n46306), .Z(n46311) );
  NAND U47013 ( .A(n46309), .B(n46308), .Z(n46310) );
  AND U47014 ( .A(n46311), .B(n46310), .Z(n46414) );
  XOR U47015 ( .A(n46415), .B(n46414), .Z(n46340) );
  XOR U47016 ( .A(n46343), .B(n46342), .Z(n46337) );
  NAND U47017 ( .A(n46313), .B(n46312), .Z(n46317) );
  NAND U47018 ( .A(n46315), .B(n46314), .Z(n46316) );
  AND U47019 ( .A(n46317), .B(n46316), .Z(n46335) );
  NAND U47020 ( .A(n46319), .B(n46318), .Z(n46323) );
  NANDN U47021 ( .A(n46321), .B(n46320), .Z(n46322) );
  NAND U47022 ( .A(n46323), .B(n46322), .Z(n46334) );
  XOR U47023 ( .A(n46437), .B(n46436), .Z(n46438) );
  XOR U47024 ( .A(n46439), .B(n46438), .Z(n46445) );
  NAND U47025 ( .A(n46328), .B(n46327), .Z(n46332) );
  NANDN U47026 ( .A(n46330), .B(n46329), .Z(n46331) );
  AND U47027 ( .A(n46332), .B(n46331), .Z(n46444) );
  IV U47028 ( .A(n46444), .Z(n46442) );
  XOR U47029 ( .A(n46443), .B(n46442), .Z(n46333) );
  XNOR U47030 ( .A(n46445), .B(n46333), .Z(N1011) );
  NANDN U47031 ( .A(n46335), .B(n46334), .Z(n46339) );
  NANDN U47032 ( .A(n46337), .B(n46336), .Z(n46338) );
  AND U47033 ( .A(n46339), .B(n46338), .Z(n46453) );
  NANDN U47034 ( .A(n46341), .B(n46340), .Z(n46345) );
  NAND U47035 ( .A(n46343), .B(n46342), .Z(n46344) );
  AND U47036 ( .A(n46345), .B(n46344), .Z(n46451) );
  NANDN U47037 ( .A(n46347), .B(n46346), .Z(n46351) );
  NANDN U47038 ( .A(n46349), .B(n46348), .Z(n46350) );
  AND U47039 ( .A(n46351), .B(n46350), .Z(n46551) );
  AND U47040 ( .A(x[486]), .B(y[8173]), .Z(n46353) );
  NAND U47041 ( .A(n46353), .B(n46352), .Z(n46357) );
  NAND U47042 ( .A(n46355), .B(n46354), .Z(n46356) );
  AND U47043 ( .A(n46357), .B(n46356), .Z(n46544) );
  AND U47044 ( .A(x[496]), .B(y[8167]), .Z(n46901) );
  NAND U47045 ( .A(n46901), .B(n46724), .Z(n46361) );
  NANDN U47046 ( .A(n46359), .B(n46358), .Z(n46360) );
  AND U47047 ( .A(n46361), .B(n46360), .Z(n46543) );
  AND U47048 ( .A(x[495]), .B(y[8169]), .Z(n47186) );
  NAND U47049 ( .A(n47186), .B(n46497), .Z(n46365) );
  NANDN U47050 ( .A(n46363), .B(n46362), .Z(n46364) );
  NAND U47051 ( .A(n46365), .B(n46364), .Z(n46527) );
  AND U47052 ( .A(y[8178]), .B(x[481]), .Z(n46367) );
  NAND U47053 ( .A(y[8171]), .B(x[488]), .Z(n46366) );
  XNOR U47054 ( .A(n46367), .B(n46366), .Z(n46488) );
  AND U47055 ( .A(y[8166]), .B(x[493]), .Z(n46369) );
  NAND U47056 ( .A(y[8177]), .B(x[482]), .Z(n46368) );
  XNOR U47057 ( .A(n46369), .B(n46368), .Z(n46503) );
  XOR U47058 ( .A(n46525), .B(n46524), .Z(n46526) );
  XOR U47059 ( .A(n46527), .B(n46526), .Z(n46542) );
  XOR U47060 ( .A(n46543), .B(n46542), .Z(n46545) );
  XOR U47061 ( .A(n46544), .B(n46545), .Z(n46549) );
  AND U47062 ( .A(x[490]), .B(y[8177]), .Z(n47406) );
  IV U47063 ( .A(n47406), .Z(n47541) );
  NANDN U47064 ( .A(n47541), .B(n46370), .Z(n46374) );
  NANDN U47065 ( .A(n46372), .B(n46371), .Z(n46373) );
  NAND U47066 ( .A(n46374), .B(n46373), .Z(n46468) );
  NANDN U47067 ( .A(n46376), .B(n46375), .Z(n46380) );
  NANDN U47068 ( .A(n46378), .B(n46377), .Z(n46379) );
  NAND U47069 ( .A(n46380), .B(n46379), .Z(n46466) );
  AND U47070 ( .A(y[8163]), .B(x[496]), .Z(n47132) );
  NAND U47071 ( .A(y[8170]), .B(x[489]), .Z(n46381) );
  XNOR U47072 ( .A(n47132), .B(n46381), .Z(n46498) );
  AND U47073 ( .A(x[495]), .B(y[8164]), .Z(n46499) );
  XOR U47074 ( .A(n46498), .B(n46499), .Z(n46465) );
  XOR U47075 ( .A(n46466), .B(n46465), .Z(n46467) );
  XNOR U47076 ( .A(n46468), .B(n46467), .Z(n46538) );
  AND U47077 ( .A(x[493]), .B(y[8175]), .Z(n47760) );
  NANDN U47078 ( .A(n46382), .B(n47760), .Z(n46386) );
  NANDN U47079 ( .A(n46384), .B(n46383), .Z(n46385) );
  NAND U47080 ( .A(n46386), .B(n46385), .Z(n46462) );
  AND U47081 ( .A(y[8169]), .B(x[490]), .Z(n46388) );
  NAND U47082 ( .A(y[8162]), .B(x[497]), .Z(n46387) );
  XNOR U47083 ( .A(n46388), .B(n46387), .Z(n46494) );
  AND U47084 ( .A(x[498]), .B(y[8161]), .Z(n46517) );
  XOR U47085 ( .A(o[499]), .B(n46517), .Z(n46493) );
  XOR U47086 ( .A(n46494), .B(n46493), .Z(n46460) );
  NAND U47087 ( .A(y[8176]), .B(x[483]), .Z(n46389) );
  XNOR U47088 ( .A(n46390), .B(n46389), .Z(n46511) );
  XOR U47089 ( .A(n46460), .B(n46459), .Z(n46461) );
  XNOR U47090 ( .A(n46462), .B(n46461), .Z(n46537) );
  NAND U47091 ( .A(n46392), .B(n46391), .Z(n46396) );
  NAND U47092 ( .A(n46394), .B(n46393), .Z(n46395) );
  AND U47093 ( .A(n46396), .B(n46395), .Z(n46521) );
  ANDN U47094 ( .B(o[498]), .A(n46397), .Z(n46478) );
  AND U47095 ( .A(x[480]), .B(y[8179]), .Z(n46475) );
  AND U47096 ( .A(x[499]), .B(y[8160]), .Z(n46476) );
  XOR U47097 ( .A(n46475), .B(n46476), .Z(n46477) );
  XOR U47098 ( .A(n46478), .B(n46477), .Z(n46519) );
  AND U47099 ( .A(x[484]), .B(y[8175]), .Z(n46633) );
  AND U47100 ( .A(y[8174]), .B(x[485]), .Z(n46399) );
  NAND U47101 ( .A(y[8173]), .B(x[486]), .Z(n46398) );
  XNOR U47102 ( .A(n46399), .B(n46398), .Z(n46472) );
  XOR U47103 ( .A(n46633), .B(n46472), .Z(n46518) );
  XOR U47104 ( .A(n46519), .B(n46518), .Z(n46520) );
  XOR U47105 ( .A(n46521), .B(n46520), .Z(n46536) );
  XNOR U47106 ( .A(n46537), .B(n46536), .Z(n46539) );
  XOR U47107 ( .A(n46538), .B(n46539), .Z(n46532) );
  NANDN U47108 ( .A(n46401), .B(n46400), .Z(n46405) );
  NANDN U47109 ( .A(n46403), .B(n46402), .Z(n46404) );
  AND U47110 ( .A(n46405), .B(n46404), .Z(n46531) );
  NANDN U47111 ( .A(n46407), .B(n46406), .Z(n46411) );
  NANDN U47112 ( .A(n46409), .B(n46408), .Z(n46410) );
  NAND U47113 ( .A(n46411), .B(n46410), .Z(n46530) );
  XOR U47114 ( .A(n46531), .B(n46530), .Z(n46533) );
  XOR U47115 ( .A(n46532), .B(n46533), .Z(n46548) );
  XNOR U47116 ( .A(n46549), .B(n46548), .Z(n46550) );
  XOR U47117 ( .A(n46551), .B(n46550), .Z(n46562) );
  NAND U47118 ( .A(n46413), .B(n46412), .Z(n46417) );
  NAND U47119 ( .A(n46415), .B(n46414), .Z(n46416) );
  AND U47120 ( .A(n46417), .B(n46416), .Z(n46560) );
  NAND U47121 ( .A(n46419), .B(n46418), .Z(n46423) );
  NAND U47122 ( .A(n46421), .B(n46420), .Z(n46422) );
  NAND U47123 ( .A(n46423), .B(n46422), .Z(n46556) );
  NAND U47124 ( .A(n46425), .B(n46424), .Z(n46429) );
  NAND U47125 ( .A(n46427), .B(n46426), .Z(n46428) );
  NAND U47126 ( .A(n46429), .B(n46428), .Z(n46555) );
  NAND U47127 ( .A(n46431), .B(n46430), .Z(n46435) );
  NAND U47128 ( .A(n46433), .B(n46432), .Z(n46434) );
  NAND U47129 ( .A(n46435), .B(n46434), .Z(n46554) );
  XNOR U47130 ( .A(n46555), .B(n46554), .Z(n46557) );
  XNOR U47131 ( .A(n46560), .B(n46561), .Z(n46563) );
  XOR U47132 ( .A(n46562), .B(n46563), .Z(n46450) );
  XOR U47133 ( .A(n46451), .B(n46450), .Z(n46452) );
  XOR U47134 ( .A(n46453), .B(n46452), .Z(n46458) );
  NAND U47135 ( .A(n46437), .B(n46436), .Z(n46441) );
  NAND U47136 ( .A(n46439), .B(n46438), .Z(n46440) );
  NAND U47137 ( .A(n46441), .B(n46440), .Z(n46457) );
  NANDN U47138 ( .A(n46442), .B(n46443), .Z(n46448) );
  NOR U47139 ( .A(n46444), .B(n46443), .Z(n46446) );
  OR U47140 ( .A(n46446), .B(n46445), .Z(n46447) );
  AND U47141 ( .A(n46448), .B(n46447), .Z(n46456) );
  XOR U47142 ( .A(n46457), .B(n46456), .Z(n46449) );
  XNOR U47143 ( .A(n46458), .B(n46449), .Z(N1012) );
  NAND U47144 ( .A(n46451), .B(n46450), .Z(n46455) );
  NANDN U47145 ( .A(n46453), .B(n46452), .Z(n46454) );
  NAND U47146 ( .A(n46455), .B(n46454), .Z(n46681) );
  IV U47147 ( .A(n46681), .Z(n46680) );
  NAND U47148 ( .A(n46460), .B(n46459), .Z(n46464) );
  NAND U47149 ( .A(n46462), .B(n46461), .Z(n46463) );
  AND U47150 ( .A(n46464), .B(n46463), .Z(n46663) );
  NAND U47151 ( .A(n46466), .B(n46465), .Z(n46470) );
  NAND U47152 ( .A(n46468), .B(n46467), .Z(n46469) );
  AND U47153 ( .A(n46470), .B(n46469), .Z(n46604) );
  NAND U47154 ( .A(x[486]), .B(y[8174]), .Z(n46590) );
  NANDN U47155 ( .A(n46590), .B(n46471), .Z(n46474) );
  NAND U47156 ( .A(n46472), .B(n46633), .Z(n46473) );
  NAND U47157 ( .A(n46474), .B(n46473), .Z(n46598) );
  NAND U47158 ( .A(n46476), .B(n46475), .Z(n46480) );
  NAND U47159 ( .A(n46478), .B(n46477), .Z(n46479) );
  NAND U47160 ( .A(n46480), .B(n46479), .Z(n46596) );
  AND U47161 ( .A(y[8162]), .B(x[498]), .Z(n46482) );
  NAND U47162 ( .A(y[8168]), .B(x[492]), .Z(n46481) );
  XNOR U47163 ( .A(n46482), .B(n46481), .Z(n46580) );
  AND U47164 ( .A(x[497]), .B(y[8163]), .Z(n46581) );
  XOR U47165 ( .A(n46580), .B(n46581), .Z(n46595) );
  XOR U47166 ( .A(n46596), .B(n46595), .Z(n46597) );
  XNOR U47167 ( .A(n46598), .B(n46597), .Z(n46602) );
  AND U47168 ( .A(y[8167]), .B(x[493]), .Z(n46484) );
  NAND U47169 ( .A(y[8177]), .B(x[483]), .Z(n46483) );
  XNOR U47170 ( .A(n46484), .B(n46483), .Z(n46620) );
  XNOR U47171 ( .A(n46620), .B(n46619), .Z(n46592) );
  AND U47172 ( .A(y[8175]), .B(x[485]), .Z(n46486) );
  NAND U47173 ( .A(y[8176]), .B(x[484]), .Z(n46485) );
  XNOR U47174 ( .A(n46486), .B(n46485), .Z(n46635) );
  AND U47175 ( .A(x[487]), .B(y[8173]), .Z(n46634) );
  XNOR U47176 ( .A(n46635), .B(n46634), .Z(n46589) );
  XOR U47177 ( .A(n46590), .B(n46589), .Z(n46591) );
  XNOR U47178 ( .A(n46592), .B(n46591), .Z(n46646) );
  AND U47179 ( .A(x[488]), .B(y[8178]), .Z(n47713) );
  AND U47180 ( .A(x[481]), .B(y[8171]), .Z(n46487) );
  NAND U47181 ( .A(n47713), .B(n46487), .Z(n46491) );
  NANDN U47182 ( .A(n46489), .B(n46488), .Z(n46490) );
  NAND U47183 ( .A(n46491), .B(n46490), .Z(n46645) );
  NAND U47184 ( .A(x[497]), .B(y[8169]), .Z(n47452) );
  NANDN U47185 ( .A(n47452), .B(n46492), .Z(n46496) );
  NAND U47186 ( .A(n46494), .B(n46493), .Z(n46495) );
  NAND U47187 ( .A(n46496), .B(n46495), .Z(n46644) );
  XOR U47188 ( .A(n46645), .B(n46644), .Z(n46647) );
  XNOR U47189 ( .A(n46646), .B(n46647), .Z(n46601) );
  XOR U47190 ( .A(n46602), .B(n46601), .Z(n46603) );
  XOR U47191 ( .A(n46604), .B(n46603), .Z(n46662) );
  XOR U47192 ( .A(n46663), .B(n46662), .Z(n46665) );
  AND U47193 ( .A(x[496]), .B(y[8170]), .Z(n47444) );
  NAND U47194 ( .A(n47444), .B(n46497), .Z(n46501) );
  NAND U47195 ( .A(n46499), .B(n46498), .Z(n46500) );
  NAND U47196 ( .A(n46501), .B(n46500), .Z(n46608) );
  AND U47197 ( .A(x[493]), .B(y[8177]), .Z(n47999) );
  NAND U47198 ( .A(n47999), .B(n46502), .Z(n46506) );
  NANDN U47199 ( .A(n46504), .B(n46503), .Z(n46505) );
  NAND U47200 ( .A(n46506), .B(n46505), .Z(n46653) );
  AND U47201 ( .A(y[8164]), .B(x[496]), .Z(n46508) );
  NAND U47202 ( .A(y[8170]), .B(x[490]), .Z(n46507) );
  XNOR U47203 ( .A(n46508), .B(n46507), .Z(n46614) );
  AND U47204 ( .A(x[482]), .B(y[8178]), .Z(n46615) );
  XOR U47205 ( .A(n46614), .B(n46615), .Z(n46651) );
  NAND U47206 ( .A(y[8171]), .B(x[489]), .Z(n46509) );
  XNOR U47207 ( .A(n46510), .B(n46509), .Z(n46574) );
  AND U47208 ( .A(x[494]), .B(y[8166]), .Z(n46575) );
  XOR U47209 ( .A(n46574), .B(n46575), .Z(n46650) );
  XOR U47210 ( .A(n46651), .B(n46650), .Z(n46652) );
  XOR U47211 ( .A(n46653), .B(n46652), .Z(n46607) );
  XOR U47212 ( .A(n46608), .B(n46607), .Z(n46610) );
  AND U47213 ( .A(x[491]), .B(y[8176]), .Z(n47544) );
  NAND U47214 ( .A(n46751), .B(n47544), .Z(n46514) );
  NANDN U47215 ( .A(n46512), .B(n46511), .Z(n46513) );
  NAND U47216 ( .A(n46514), .B(n46513), .Z(n46659) );
  AND U47217 ( .A(y[8169]), .B(x[491]), .Z(n46516) );
  NAND U47218 ( .A(y[8179]), .B(x[481]), .Z(n46515) );
  XNOR U47219 ( .A(n46516), .B(n46515), .Z(n46586) );
  AND U47220 ( .A(x[499]), .B(y[8161]), .Z(n46578) );
  XOR U47221 ( .A(o[500]), .B(n46578), .Z(n46585) );
  XOR U47222 ( .A(n46586), .B(n46585), .Z(n46657) );
  AND U47223 ( .A(x[480]), .B(y[8180]), .Z(n46638) );
  AND U47224 ( .A(x[500]), .B(y[8160]), .Z(n46639) );
  XOR U47225 ( .A(n46638), .B(n46639), .Z(n46641) );
  AND U47226 ( .A(o[499]), .B(n46517), .Z(n46640) );
  XOR U47227 ( .A(n46641), .B(n46640), .Z(n46656) );
  XOR U47228 ( .A(n46657), .B(n46656), .Z(n46658) );
  XOR U47229 ( .A(n46659), .B(n46658), .Z(n46609) );
  XNOR U47230 ( .A(n46610), .B(n46609), .Z(n46570) );
  NAND U47231 ( .A(n46519), .B(n46518), .Z(n46523) );
  NANDN U47232 ( .A(n46521), .B(n46520), .Z(n46522) );
  AND U47233 ( .A(n46523), .B(n46522), .Z(n46567) );
  NAND U47234 ( .A(n46525), .B(n46524), .Z(n46529) );
  NAND U47235 ( .A(n46527), .B(n46526), .Z(n46528) );
  AND U47236 ( .A(n46529), .B(n46528), .Z(n46568) );
  XOR U47237 ( .A(n46567), .B(n46568), .Z(n46569) );
  XOR U47238 ( .A(n46570), .B(n46569), .Z(n46664) );
  XOR U47239 ( .A(n46665), .B(n46664), .Z(n46669) );
  NANDN U47240 ( .A(n46531), .B(n46530), .Z(n46535) );
  NANDN U47241 ( .A(n46533), .B(n46532), .Z(n46534) );
  AND U47242 ( .A(n46535), .B(n46534), .Z(n46677) );
  NAND U47243 ( .A(n46537), .B(n46536), .Z(n46541) );
  NANDN U47244 ( .A(n46539), .B(n46538), .Z(n46540) );
  AND U47245 ( .A(n46541), .B(n46540), .Z(n46675) );
  NANDN U47246 ( .A(n46543), .B(n46542), .Z(n46547) );
  OR U47247 ( .A(n46545), .B(n46544), .Z(n46546) );
  AND U47248 ( .A(n46547), .B(n46546), .Z(n46674) );
  XNOR U47249 ( .A(n46675), .B(n46674), .Z(n46676) );
  XNOR U47250 ( .A(n46677), .B(n46676), .Z(n46668) );
  XNOR U47251 ( .A(n46669), .B(n46668), .Z(n46670) );
  NANDN U47252 ( .A(n46549), .B(n46548), .Z(n46553) );
  NANDN U47253 ( .A(n46551), .B(n46550), .Z(n46552) );
  NAND U47254 ( .A(n46553), .B(n46552), .Z(n46671) );
  XOR U47255 ( .A(n46670), .B(n46671), .Z(n46689) );
  NAND U47256 ( .A(n46555), .B(n46554), .Z(n46559) );
  NANDN U47257 ( .A(n46557), .B(n46556), .Z(n46558) );
  AND U47258 ( .A(n46559), .B(n46558), .Z(n46688) );
  NANDN U47259 ( .A(n46561), .B(n46560), .Z(n46565) );
  NAND U47260 ( .A(n46563), .B(n46562), .Z(n46564) );
  AND U47261 ( .A(n46565), .B(n46564), .Z(n46687) );
  XOR U47262 ( .A(n46688), .B(n46687), .Z(n46690) );
  XOR U47263 ( .A(n46689), .B(n46690), .Z(n46683) );
  XNOR U47264 ( .A(n46682), .B(n46683), .Z(n46566) );
  XOR U47265 ( .A(n46680), .B(n46566), .Z(N1013) );
  NAND U47266 ( .A(n46568), .B(n46567), .Z(n46572) );
  NAND U47267 ( .A(n46570), .B(n46569), .Z(n46571) );
  AND U47268 ( .A(n46572), .B(n46571), .Z(n46703) );
  AND U47269 ( .A(x[495]), .B(y[8171]), .Z(n47439) );
  NAND U47270 ( .A(n47439), .B(n46573), .Z(n46577) );
  NAND U47271 ( .A(n46575), .B(n46574), .Z(n46576) );
  AND U47272 ( .A(n46577), .B(n46576), .Z(n46738) );
  AND U47273 ( .A(x[480]), .B(y[8181]), .Z(n46757) );
  AND U47274 ( .A(x[501]), .B(y[8160]), .Z(n46758) );
  XOR U47275 ( .A(n46757), .B(n46758), .Z(n46760) );
  AND U47276 ( .A(o[500]), .B(n46578), .Z(n46759) );
  XOR U47277 ( .A(n46760), .B(n46759), .Z(n46736) );
  AND U47278 ( .A(x[485]), .B(y[8176]), .Z(n46744) );
  AND U47279 ( .A(x[496]), .B(y[8165]), .Z(n46743) );
  XOR U47280 ( .A(n46744), .B(n46743), .Z(n46742) );
  AND U47281 ( .A(x[495]), .B(y[8166]), .Z(n46741) );
  XOR U47282 ( .A(n46742), .B(n46741), .Z(n46735) );
  XOR U47283 ( .A(n46736), .B(n46735), .Z(n46737) );
  AND U47284 ( .A(x[498]), .B(y[8168]), .Z(n47451) );
  NAND U47285 ( .A(n47451), .B(n46579), .Z(n46583) );
  NAND U47286 ( .A(n46581), .B(n46580), .Z(n46582) );
  NAND U47287 ( .A(n46583), .B(n46582), .Z(n46780) );
  AND U47288 ( .A(x[491]), .B(y[8179]), .Z(n48161) );
  AND U47289 ( .A(x[481]), .B(y[8169]), .Z(n46584) );
  NAND U47290 ( .A(n48161), .B(n46584), .Z(n46588) );
  NAND U47291 ( .A(n46586), .B(n46585), .Z(n46587) );
  NAND U47292 ( .A(n46588), .B(n46587), .Z(n46779) );
  XOR U47293 ( .A(n46780), .B(n46779), .Z(n46781) );
  XNOR U47294 ( .A(n46782), .B(n46781), .Z(n46774) );
  NAND U47295 ( .A(n46590), .B(n46589), .Z(n46594) );
  NAND U47296 ( .A(n46592), .B(n46591), .Z(n46593) );
  NAND U47297 ( .A(n46594), .B(n46593), .Z(n46773) );
  XOR U47298 ( .A(n46774), .B(n46773), .Z(n46776) );
  NAND U47299 ( .A(n46596), .B(n46595), .Z(n46600) );
  NAND U47300 ( .A(n46598), .B(n46597), .Z(n46599) );
  AND U47301 ( .A(n46600), .B(n46599), .Z(n46775) );
  XNOR U47302 ( .A(n46776), .B(n46775), .Z(n46701) );
  NAND U47303 ( .A(n46602), .B(n46601), .Z(n46606) );
  NAND U47304 ( .A(n46604), .B(n46603), .Z(n46605) );
  AND U47305 ( .A(n46606), .B(n46605), .Z(n46700) );
  XOR U47306 ( .A(n46701), .B(n46700), .Z(n46702) );
  XNOR U47307 ( .A(n46703), .B(n46702), .Z(n46697) );
  NAND U47308 ( .A(n46608), .B(n46607), .Z(n46612) );
  NAND U47309 ( .A(n46610), .B(n46609), .Z(n46611) );
  NAND U47310 ( .A(n46612), .B(n46611), .Z(n46800) );
  NAND U47311 ( .A(n47444), .B(n46613), .Z(n46617) );
  NAND U47312 ( .A(n46615), .B(n46614), .Z(n46616) );
  NAND U47313 ( .A(n46617), .B(n46616), .Z(n46707) );
  NAND U47314 ( .A(n47999), .B(n46618), .Z(n46622) );
  NAND U47315 ( .A(n46620), .B(n46619), .Z(n46621) );
  NAND U47316 ( .A(n46622), .B(n46621), .Z(n46794) );
  AND U47317 ( .A(y[8162]), .B(x[499]), .Z(n46624) );
  NAND U47318 ( .A(y[8170]), .B(x[491]), .Z(n46623) );
  XNOR U47319 ( .A(n46624), .B(n46623), .Z(n46726) );
  AND U47320 ( .A(x[500]), .B(y[8161]), .Z(n46756) );
  XOR U47321 ( .A(o[501]), .B(n46756), .Z(n46725) );
  XOR U47322 ( .A(n46726), .B(n46725), .Z(n46792) );
  AND U47323 ( .A(y[8163]), .B(x[498]), .Z(n46626) );
  NAND U47324 ( .A(y[8171]), .B(x[490]), .Z(n46625) );
  XNOR U47325 ( .A(n46626), .B(n46625), .Z(n46764) );
  AND U47326 ( .A(x[481]), .B(y[8180]), .Z(n46765) );
  XOR U47327 ( .A(n46764), .B(n46765), .Z(n46791) );
  XOR U47328 ( .A(n46792), .B(n46791), .Z(n46793) );
  XOR U47329 ( .A(n46794), .B(n46793), .Z(n46706) );
  XOR U47330 ( .A(n46707), .B(n46706), .Z(n46709) );
  AND U47331 ( .A(x[487]), .B(y[8174]), .Z(n46973) );
  AND U47332 ( .A(y[8175]), .B(x[486]), .Z(n46628) );
  NAND U47333 ( .A(y[8167]), .B(x[494]), .Z(n46627) );
  XNOR U47334 ( .A(n46628), .B(n46627), .Z(n46768) );
  XOR U47335 ( .A(n46973), .B(n46768), .Z(n46715) );
  AND U47336 ( .A(x[489]), .B(y[8172]), .Z(n46713) );
  NAND U47337 ( .A(x[488]), .B(y[8173]), .Z(n46712) );
  AND U47338 ( .A(y[8169]), .B(x[492]), .Z(n46630) );
  NAND U47339 ( .A(y[8164]), .B(x[497]), .Z(n46629) );
  XNOR U47340 ( .A(n46630), .B(n46629), .Z(n46718) );
  AND U47341 ( .A(x[482]), .B(y[8179]), .Z(n46719) );
  XOR U47342 ( .A(n46718), .B(n46719), .Z(n46730) );
  AND U47343 ( .A(y[8168]), .B(x[493]), .Z(n46632) );
  NAND U47344 ( .A(y[8178]), .B(x[483]), .Z(n46631) );
  XNOR U47345 ( .A(n46632), .B(n46631), .Z(n46752) );
  AND U47346 ( .A(x[484]), .B(y[8177]), .Z(n46753) );
  XOR U47347 ( .A(n46752), .B(n46753), .Z(n46729) );
  XOR U47348 ( .A(n46730), .B(n46729), .Z(n46732) );
  XOR U47349 ( .A(n46731), .B(n46732), .Z(n46788) );
  NAND U47350 ( .A(n46744), .B(n46633), .Z(n46637) );
  NAND U47351 ( .A(n46635), .B(n46634), .Z(n46636) );
  NAND U47352 ( .A(n46637), .B(n46636), .Z(n46786) );
  NAND U47353 ( .A(n46639), .B(n46638), .Z(n46643) );
  NAND U47354 ( .A(n46641), .B(n46640), .Z(n46642) );
  NAND U47355 ( .A(n46643), .B(n46642), .Z(n46785) );
  XOR U47356 ( .A(n46786), .B(n46785), .Z(n46787) );
  XOR U47357 ( .A(n46788), .B(n46787), .Z(n46708) );
  XOR U47358 ( .A(n46709), .B(n46708), .Z(n46798) );
  NAND U47359 ( .A(n46645), .B(n46644), .Z(n46649) );
  NAND U47360 ( .A(n46647), .B(n46646), .Z(n46648) );
  NAND U47361 ( .A(n46649), .B(n46648), .Z(n46805) );
  NAND U47362 ( .A(n46651), .B(n46650), .Z(n46655) );
  NAND U47363 ( .A(n46653), .B(n46652), .Z(n46654) );
  NAND U47364 ( .A(n46655), .B(n46654), .Z(n46804) );
  NAND U47365 ( .A(n46657), .B(n46656), .Z(n46661) );
  NAND U47366 ( .A(n46659), .B(n46658), .Z(n46660) );
  NAND U47367 ( .A(n46661), .B(n46660), .Z(n46803) );
  XOR U47368 ( .A(n46804), .B(n46803), .Z(n46806) );
  XOR U47369 ( .A(n46805), .B(n46806), .Z(n46797) );
  XOR U47370 ( .A(n46798), .B(n46797), .Z(n46799) );
  XNOR U47371 ( .A(n46800), .B(n46799), .Z(n46695) );
  NAND U47372 ( .A(n46663), .B(n46662), .Z(n46667) );
  NAND U47373 ( .A(n46665), .B(n46664), .Z(n46666) );
  NAND U47374 ( .A(n46667), .B(n46666), .Z(n46694) );
  XOR U47375 ( .A(n46695), .B(n46694), .Z(n46696) );
  XNOR U47376 ( .A(n46697), .B(n46696), .Z(n46818) );
  NANDN U47377 ( .A(n46669), .B(n46668), .Z(n46673) );
  NANDN U47378 ( .A(n46671), .B(n46670), .Z(n46672) );
  AND U47379 ( .A(n46673), .B(n46672), .Z(n46817) );
  NANDN U47380 ( .A(n46675), .B(n46674), .Z(n46679) );
  NAND U47381 ( .A(n46677), .B(n46676), .Z(n46678) );
  AND U47382 ( .A(n46679), .B(n46678), .Z(n46816) );
  XOR U47383 ( .A(n46817), .B(n46816), .Z(n46819) );
  XOR U47384 ( .A(n46818), .B(n46819), .Z(n46812) );
  OR U47385 ( .A(n46682), .B(n46680), .Z(n46686) );
  ANDN U47386 ( .B(n46682), .A(n46681), .Z(n46684) );
  OR U47387 ( .A(n46684), .B(n46683), .Z(n46685) );
  AND U47388 ( .A(n46686), .B(n46685), .Z(n46811) );
  NAND U47389 ( .A(n46688), .B(n46687), .Z(n46692) );
  NAND U47390 ( .A(n46690), .B(n46689), .Z(n46691) );
  AND U47391 ( .A(n46692), .B(n46691), .Z(n46810) );
  IV U47392 ( .A(n46810), .Z(n46809) );
  XOR U47393 ( .A(n46811), .B(n46809), .Z(n46693) );
  XNOR U47394 ( .A(n46812), .B(n46693), .Z(N1014) );
  NAND U47395 ( .A(n46695), .B(n46694), .Z(n46699) );
  NAND U47396 ( .A(n46697), .B(n46696), .Z(n46698) );
  AND U47397 ( .A(n46699), .B(n46698), .Z(n46949) );
  NAND U47398 ( .A(n46701), .B(n46700), .Z(n46705) );
  NAND U47399 ( .A(n46703), .B(n46702), .Z(n46704) );
  NAND U47400 ( .A(n46705), .B(n46704), .Z(n46947) );
  NAND U47401 ( .A(n46707), .B(n46706), .Z(n46711) );
  NAND U47402 ( .A(n46709), .B(n46708), .Z(n46710) );
  NAND U47403 ( .A(n46711), .B(n46710), .Z(n46940) );
  NANDN U47404 ( .A(n46713), .B(n46712), .Z(n46717) );
  NANDN U47405 ( .A(n46715), .B(n46714), .Z(n46716) );
  NAND U47406 ( .A(n46717), .B(n46716), .Z(n46934) );
  NANDN U47407 ( .A(n47452), .B(n46885), .Z(n46721) );
  NAND U47408 ( .A(n46719), .B(n46718), .Z(n46720) );
  NAND U47409 ( .A(n46721), .B(n46720), .Z(n46861) );
  AND U47410 ( .A(x[485]), .B(y[8177]), .Z(n46907) );
  AND U47411 ( .A(x[497]), .B(y[8165]), .Z(n46908) );
  XOR U47412 ( .A(n46907), .B(n46908), .Z(n46909) );
  AND U47413 ( .A(x[496]), .B(y[8166]), .Z(n46910) );
  XOR U47414 ( .A(n46909), .B(n46910), .Z(n46860) );
  AND U47415 ( .A(y[8164]), .B(x[498]), .Z(n46723) );
  NAND U47416 ( .A(y[8170]), .B(x[492]), .Z(n46722) );
  XNOR U47417 ( .A(n46723), .B(n46722), .Z(n46886) );
  AND U47418 ( .A(x[484]), .B(y[8178]), .Z(n46887) );
  XOR U47419 ( .A(n46886), .B(n46887), .Z(n46859) );
  XOR U47420 ( .A(n46860), .B(n46859), .Z(n46862) );
  XNOR U47421 ( .A(n46861), .B(n46862), .Z(n46931) );
  AND U47422 ( .A(x[499]), .B(y[8170]), .Z(n47884) );
  NAND U47423 ( .A(n47884), .B(n46724), .Z(n46728) );
  NAND U47424 ( .A(n46726), .B(n46725), .Z(n46727) );
  AND U47425 ( .A(n46728), .B(n46727), .Z(n46932) );
  XOR U47426 ( .A(n46931), .B(n46932), .Z(n46933) );
  XNOR U47427 ( .A(n46934), .B(n46933), .Z(n46937) );
  NAND U47428 ( .A(n46730), .B(n46729), .Z(n46734) );
  NAND U47429 ( .A(n46732), .B(n46731), .Z(n46733) );
  NAND U47430 ( .A(n46734), .B(n46733), .Z(n46920) );
  NAND U47431 ( .A(n46736), .B(n46735), .Z(n46740) );
  NANDN U47432 ( .A(n46738), .B(n46737), .Z(n46739) );
  NAND U47433 ( .A(n46740), .B(n46739), .Z(n46919) );
  XOR U47434 ( .A(n46920), .B(n46919), .Z(n46922) );
  AND U47435 ( .A(n46742), .B(n46741), .Z(n46746) );
  NAND U47436 ( .A(n46744), .B(n46743), .Z(n46745) );
  NANDN U47437 ( .A(n46746), .B(n46745), .Z(n46882) );
  AND U47438 ( .A(y[8169]), .B(x[493]), .Z(n46748) );
  NAND U47439 ( .A(y[8162]), .B(x[500]), .Z(n46747) );
  XNOR U47440 ( .A(n46748), .B(n46747), .Z(n46903) );
  AND U47441 ( .A(x[482]), .B(y[8180]), .Z(n46904) );
  XOR U47442 ( .A(n46903), .B(n46904), .Z(n46880) );
  AND U47443 ( .A(y[8176]), .B(x[486]), .Z(n46750) );
  NAND U47444 ( .A(y[8167]), .B(x[495]), .Z(n46749) );
  XNOR U47445 ( .A(n46750), .B(n46749), .Z(n46915) );
  XOR U47446 ( .A(n46880), .B(n46879), .Z(n46881) );
  XOR U47447 ( .A(n46882), .B(n46881), .Z(n46926) );
  AND U47448 ( .A(x[493]), .B(y[8178]), .Z(n48158) );
  NAND U47449 ( .A(n46751), .B(n48158), .Z(n46755) );
  NAND U47450 ( .A(n46753), .B(n46752), .Z(n46754) );
  NAND U47451 ( .A(n46755), .B(n46754), .Z(n46850) );
  AND U47452 ( .A(x[481]), .B(y[8181]), .Z(n46873) );
  XOR U47453 ( .A(n46874), .B(n46873), .Z(n46872) );
  AND U47454 ( .A(o[501]), .B(n46756), .Z(n46871) );
  XOR U47455 ( .A(n46872), .B(n46871), .Z(n46848) );
  AND U47456 ( .A(x[494]), .B(y[8168]), .Z(n46865) );
  AND U47457 ( .A(x[483]), .B(y[8179]), .Z(n46866) );
  XOR U47458 ( .A(n46865), .B(n46866), .Z(n46867) );
  AND U47459 ( .A(x[499]), .B(y[8163]), .Z(n46868) );
  XOR U47460 ( .A(n46867), .B(n46868), .Z(n46847) );
  XOR U47461 ( .A(n46848), .B(n46847), .Z(n46849) );
  XOR U47462 ( .A(n46850), .B(n46849), .Z(n46925) );
  XOR U47463 ( .A(n46926), .B(n46925), .Z(n46928) );
  NAND U47464 ( .A(n46758), .B(n46757), .Z(n46762) );
  NAND U47465 ( .A(n46760), .B(n46759), .Z(n46761) );
  NAND U47466 ( .A(n46762), .B(n46761), .Z(n46842) );
  AND U47467 ( .A(x[498]), .B(y[8171]), .Z(n47887) );
  NAND U47468 ( .A(n47887), .B(n46763), .Z(n46767) );
  NAND U47469 ( .A(n46765), .B(n46764), .Z(n46766) );
  NAND U47470 ( .A(n46767), .B(n46766), .Z(n46841) );
  XOR U47471 ( .A(n46842), .B(n46841), .Z(n46844) );
  AND U47472 ( .A(x[494]), .B(y[8175]), .Z(n47927) );
  NAND U47473 ( .A(n47927), .B(n46914), .Z(n46770) );
  NAND U47474 ( .A(n46973), .B(n46768), .Z(n46769) );
  NAND U47475 ( .A(n46770), .B(n46769), .Z(n46856) );
  AND U47476 ( .A(x[480]), .B(y[8182]), .Z(n46890) );
  AND U47477 ( .A(x[502]), .B(y[8160]), .Z(n46891) );
  XOR U47478 ( .A(n46890), .B(n46891), .Z(n46893) );
  AND U47479 ( .A(x[501]), .B(y[8161]), .Z(n46913) );
  XOR U47480 ( .A(o[502]), .B(n46913), .Z(n46892) );
  XOR U47481 ( .A(n46893), .B(n46892), .Z(n46854) );
  AND U47482 ( .A(y[8175]), .B(x[487]), .Z(n46772) );
  NAND U47483 ( .A(y[8174]), .B(x[488]), .Z(n46771) );
  XNOR U47484 ( .A(n46772), .B(n46771), .Z(n46896) );
  XOR U47485 ( .A(n46854), .B(n46853), .Z(n46855) );
  XOR U47486 ( .A(n46856), .B(n46855), .Z(n46843) );
  XOR U47487 ( .A(n46844), .B(n46843), .Z(n46927) );
  XOR U47488 ( .A(n46928), .B(n46927), .Z(n46921) );
  XOR U47489 ( .A(n46922), .B(n46921), .Z(n46938) );
  XOR U47490 ( .A(n46937), .B(n46938), .Z(n46939) );
  XNOR U47491 ( .A(n46940), .B(n46939), .Z(n46831) );
  NAND U47492 ( .A(n46774), .B(n46773), .Z(n46778) );
  NAND U47493 ( .A(n46776), .B(n46775), .Z(n46777) );
  NAND U47494 ( .A(n46778), .B(n46777), .Z(n46830) );
  NAND U47495 ( .A(n46780), .B(n46779), .Z(n46784) );
  NAND U47496 ( .A(n46782), .B(n46781), .Z(n46783) );
  AND U47497 ( .A(n46784), .B(n46783), .Z(n46838) );
  NAND U47498 ( .A(n46786), .B(n46785), .Z(n46790) );
  NAND U47499 ( .A(n46788), .B(n46787), .Z(n46789) );
  NAND U47500 ( .A(n46790), .B(n46789), .Z(n46836) );
  NAND U47501 ( .A(n46792), .B(n46791), .Z(n46796) );
  NAND U47502 ( .A(n46794), .B(n46793), .Z(n46795) );
  NAND U47503 ( .A(n46796), .B(n46795), .Z(n46835) );
  XOR U47504 ( .A(n46836), .B(n46835), .Z(n46837) );
  XOR U47505 ( .A(n46838), .B(n46837), .Z(n46829) );
  XOR U47506 ( .A(n46830), .B(n46829), .Z(n46832) );
  XNOR U47507 ( .A(n46831), .B(n46832), .Z(n46825) );
  NAND U47508 ( .A(n46798), .B(n46797), .Z(n46802) );
  NAND U47509 ( .A(n46800), .B(n46799), .Z(n46801) );
  NAND U47510 ( .A(n46802), .B(n46801), .Z(n46824) );
  NAND U47511 ( .A(n46804), .B(n46803), .Z(n46808) );
  NAND U47512 ( .A(n46806), .B(n46805), .Z(n46807) );
  NAND U47513 ( .A(n46808), .B(n46807), .Z(n46823) );
  XOR U47514 ( .A(n46824), .B(n46823), .Z(n46826) );
  XOR U47515 ( .A(n46825), .B(n46826), .Z(n46946) );
  XOR U47516 ( .A(n46947), .B(n46946), .Z(n46948) );
  XNOR U47517 ( .A(n46949), .B(n46948), .Z(n46943) );
  OR U47518 ( .A(n46811), .B(n46809), .Z(n46815) );
  ANDN U47519 ( .B(n46811), .A(n46810), .Z(n46813) );
  OR U47520 ( .A(n46813), .B(n46812), .Z(n46814) );
  AND U47521 ( .A(n46815), .B(n46814), .Z(n46944) );
  NANDN U47522 ( .A(n46817), .B(n46816), .Z(n46821) );
  NANDN U47523 ( .A(n46819), .B(n46818), .Z(n46820) );
  AND U47524 ( .A(n46821), .B(n46820), .Z(n46945) );
  XOR U47525 ( .A(n46944), .B(n46945), .Z(n46822) );
  XNOR U47526 ( .A(n46943), .B(n46822), .Z(N1015) );
  NAND U47527 ( .A(n46824), .B(n46823), .Z(n46828) );
  NAND U47528 ( .A(n46826), .B(n46825), .Z(n46827) );
  AND U47529 ( .A(n46828), .B(n46827), .Z(n47094) );
  NAND U47530 ( .A(n46830), .B(n46829), .Z(n46834) );
  NAND U47531 ( .A(n46832), .B(n46831), .Z(n46833) );
  NAND U47532 ( .A(n46834), .B(n46833), .Z(n47092) );
  NAND U47533 ( .A(n46836), .B(n46835), .Z(n46840) );
  NANDN U47534 ( .A(n46838), .B(n46837), .Z(n46839) );
  NAND U47535 ( .A(n46840), .B(n46839), .Z(n47069) );
  NAND U47536 ( .A(n46842), .B(n46841), .Z(n46846) );
  NAND U47537 ( .A(n46844), .B(n46843), .Z(n46845) );
  NAND U47538 ( .A(n46846), .B(n46845), .Z(n47063) );
  NAND U47539 ( .A(n46848), .B(n46847), .Z(n46852) );
  NAND U47540 ( .A(n46850), .B(n46849), .Z(n46851) );
  NAND U47541 ( .A(n46852), .B(n46851), .Z(n47061) );
  NAND U47542 ( .A(n46854), .B(n46853), .Z(n46858) );
  NAND U47543 ( .A(n46856), .B(n46855), .Z(n46857) );
  NAND U47544 ( .A(n46858), .B(n46857), .Z(n47060) );
  XOR U47545 ( .A(n47061), .B(n47060), .Z(n47062) );
  XOR U47546 ( .A(n47063), .B(n47062), .Z(n47081) );
  NAND U47547 ( .A(n46860), .B(n46859), .Z(n46864) );
  NAND U47548 ( .A(n46862), .B(n46861), .Z(n46863) );
  AND U47549 ( .A(n46864), .B(n46863), .Z(n47079) );
  NAND U47550 ( .A(n46866), .B(n46865), .Z(n46870) );
  NAND U47551 ( .A(n46868), .B(n46867), .Z(n46869) );
  NAND U47552 ( .A(n46870), .B(n46869), .Z(n47007) );
  AND U47553 ( .A(n46872), .B(n46871), .Z(n46876) );
  NAND U47554 ( .A(n46874), .B(n46873), .Z(n46875) );
  NANDN U47555 ( .A(n46876), .B(n46875), .Z(n47006) );
  XOR U47556 ( .A(n47007), .B(n47006), .Z(n47009) );
  AND U47557 ( .A(y[8176]), .B(x[487]), .Z(n46878) );
  NAND U47558 ( .A(y[8174]), .B(x[489]), .Z(n46877) );
  XNOR U47559 ( .A(n46878), .B(n46877), .Z(n46974) );
  AND U47560 ( .A(x[490]), .B(y[8173]), .Z(n47012) );
  XOR U47561 ( .A(n47013), .B(n47012), .Z(n47015) );
  AND U47562 ( .A(x[486]), .B(y[8177]), .Z(n46965) );
  NAND U47563 ( .A(x[495]), .B(y[8168]), .Z(n46966) );
  XNOR U47564 ( .A(n46965), .B(n46966), .Z(n46968) );
  AND U47565 ( .A(x[491]), .B(y[8172]), .Z(n46967) );
  XOR U47566 ( .A(n46968), .B(n46967), .Z(n47014) );
  XOR U47567 ( .A(n47015), .B(n47014), .Z(n47008) );
  XOR U47568 ( .A(n47009), .B(n47008), .Z(n47078) );
  XOR U47569 ( .A(n47081), .B(n47080), .Z(n47067) );
  NAND U47570 ( .A(n46880), .B(n46879), .Z(n46884) );
  NAND U47571 ( .A(n46882), .B(n46881), .Z(n46883) );
  NAND U47572 ( .A(n46884), .B(n46883), .Z(n47001) );
  NAND U47573 ( .A(x[498]), .B(y[8170]), .Z(n47750) );
  NANDN U47574 ( .A(n47750), .B(n46885), .Z(n46889) );
  NAND U47575 ( .A(n46887), .B(n46886), .Z(n46888) );
  AND U47576 ( .A(n46889), .B(n46888), .Z(n47037) );
  NAND U47577 ( .A(n46891), .B(n46890), .Z(n46895) );
  NAND U47578 ( .A(n46893), .B(n46892), .Z(n46894) );
  NAND U47579 ( .A(n46895), .B(n46894), .Z(n47036) );
  NANDN U47580 ( .A(n46975), .B(n46973), .Z(n46899) );
  NANDN U47581 ( .A(n46897), .B(n46896), .Z(n46898) );
  AND U47582 ( .A(n46899), .B(n46898), .Z(n47051) );
  AND U47583 ( .A(x[480]), .B(y[8183]), .Z(n46985) );
  AND U47584 ( .A(x[503]), .B(y[8160]), .Z(n46984) );
  XOR U47585 ( .A(n46985), .B(n46984), .Z(n46987) );
  AND U47586 ( .A(x[502]), .B(y[8161]), .Z(n46964) );
  XOR U47587 ( .A(n46964), .B(o[503]), .Z(n46986) );
  XOR U47588 ( .A(n46987), .B(n46986), .Z(n47048) );
  NAND U47589 ( .A(y[8163]), .B(x[500]), .Z(n46900) );
  XNOR U47590 ( .A(n46901), .B(n46900), .Z(n46960) );
  NAND U47591 ( .A(x[499]), .B(y[8164]), .Z(n46961) );
  XOR U47592 ( .A(n46960), .B(n46961), .Z(n47049) );
  XOR U47593 ( .A(n47039), .B(n47038), .Z(n47000) );
  XOR U47594 ( .A(n47001), .B(n47000), .Z(n47003) );
  NAND U47595 ( .A(x[500]), .B(y[8169]), .Z(n47937) );
  AND U47596 ( .A(x[493]), .B(y[8162]), .Z(n46902) );
  NANDN U47597 ( .A(n47937), .B(n46902), .Z(n46906) );
  NAND U47598 ( .A(n46904), .B(n46903), .Z(n46905) );
  NAND U47599 ( .A(n46906), .B(n46905), .Z(n46995) );
  NAND U47600 ( .A(n46908), .B(n46907), .Z(n46912) );
  NAND U47601 ( .A(n46910), .B(n46909), .Z(n46911) );
  AND U47602 ( .A(n46912), .B(n46911), .Z(n47057) );
  AND U47603 ( .A(x[493]), .B(y[8170]), .Z(n47030) );
  AND U47604 ( .A(x[482]), .B(y[8181]), .Z(n47031) );
  XOR U47605 ( .A(n47030), .B(n47031), .Z(n47032) );
  AND U47606 ( .A(x[501]), .B(y[8162]), .Z(n47033) );
  XOR U47607 ( .A(n47032), .B(n47033), .Z(n47055) );
  AND U47608 ( .A(x[492]), .B(y[8171]), .Z(n46978) );
  AND U47609 ( .A(x[481]), .B(y[8182]), .Z(n46979) );
  XOR U47610 ( .A(n46978), .B(n46979), .Z(n46981) );
  AND U47611 ( .A(o[502]), .B(n46913), .Z(n46980) );
  XOR U47612 ( .A(n46981), .B(n46980), .Z(n47054) );
  XOR U47613 ( .A(n47055), .B(n47054), .Z(n47056) );
  XOR U47614 ( .A(n46995), .B(n46994), .Z(n46997) );
  AND U47615 ( .A(x[495]), .B(y[8176]), .Z(n48116) );
  NAND U47616 ( .A(n48116), .B(n46914), .Z(n46918) );
  NANDN U47617 ( .A(n46916), .B(n46915), .Z(n46917) );
  AND U47618 ( .A(n46918), .B(n46917), .Z(n47045) );
  AND U47619 ( .A(x[494]), .B(y[8169]), .Z(n47024) );
  AND U47620 ( .A(x[483]), .B(y[8180]), .Z(n47025) );
  XOR U47621 ( .A(n47024), .B(n47025), .Z(n47026) );
  AND U47622 ( .A(x[484]), .B(y[8179]), .Z(n47027) );
  XOR U47623 ( .A(n47026), .B(n47027), .Z(n47042) );
  AND U47624 ( .A(x[485]), .B(y[8178]), .Z(n47018) );
  NAND U47625 ( .A(x[498]), .B(y[8165]), .Z(n47019) );
  XNOR U47626 ( .A(n47018), .B(n47019), .Z(n47020) );
  NAND U47627 ( .A(x[497]), .B(y[8166]), .Z(n47021) );
  XOR U47628 ( .A(n47020), .B(n47021), .Z(n47043) );
  XOR U47629 ( .A(n46997), .B(n46996), .Z(n47002) );
  XOR U47630 ( .A(n47003), .B(n47002), .Z(n47066) );
  XOR U47631 ( .A(n47067), .B(n47066), .Z(n47068) );
  XNOR U47632 ( .A(n47069), .B(n47068), .Z(n46955) );
  NAND U47633 ( .A(n46920), .B(n46919), .Z(n46924) );
  NAND U47634 ( .A(n46922), .B(n46921), .Z(n46923) );
  NAND U47635 ( .A(n46924), .B(n46923), .Z(n47075) );
  NAND U47636 ( .A(n46926), .B(n46925), .Z(n46930) );
  NAND U47637 ( .A(n46928), .B(n46927), .Z(n46929) );
  NAND U47638 ( .A(n46930), .B(n46929), .Z(n47073) );
  NAND U47639 ( .A(n46932), .B(n46931), .Z(n46936) );
  NAND U47640 ( .A(n46934), .B(n46933), .Z(n46935) );
  AND U47641 ( .A(n46936), .B(n46935), .Z(n47072) );
  XOR U47642 ( .A(n47073), .B(n47072), .Z(n47074) );
  XNOR U47643 ( .A(n47075), .B(n47074), .Z(n46953) );
  NAND U47644 ( .A(n46938), .B(n46937), .Z(n46942) );
  NAND U47645 ( .A(n46940), .B(n46939), .Z(n46941) );
  AND U47646 ( .A(n46942), .B(n46941), .Z(n46954) );
  XOR U47647 ( .A(n46953), .B(n46954), .Z(n46956) );
  XOR U47648 ( .A(n46955), .B(n46956), .Z(n47091) );
  XOR U47649 ( .A(n47092), .B(n47091), .Z(n47093) );
  XNOR U47650 ( .A(n47094), .B(n47093), .Z(n47087) );
  NAND U47651 ( .A(n46947), .B(n46946), .Z(n46951) );
  NAND U47652 ( .A(n46949), .B(n46948), .Z(n46950) );
  AND U47653 ( .A(n46951), .B(n46950), .Z(n47086) );
  IV U47654 ( .A(n47086), .Z(n47084) );
  XOR U47655 ( .A(n47085), .B(n47084), .Z(n46952) );
  XNOR U47656 ( .A(n47087), .B(n46952), .Z(N1016) );
  NAND U47657 ( .A(n46954), .B(n46953), .Z(n46958) );
  NAND U47658 ( .A(n46956), .B(n46955), .Z(n46957) );
  AND U47659 ( .A(n46958), .B(n46957), .Z(n47223) );
  AND U47660 ( .A(x[500]), .B(y[8167]), .Z(n46959) );
  NAND U47661 ( .A(n46959), .B(n47132), .Z(n46963) );
  NANDN U47662 ( .A(n46961), .B(n46960), .Z(n46962) );
  AND U47663 ( .A(n46963), .B(n46962), .Z(n47149) );
  AND U47664 ( .A(x[502]), .B(y[8162]), .Z(n47166) );
  XOR U47665 ( .A(n47167), .B(n47166), .Z(n47169) );
  AND U47666 ( .A(x[482]), .B(y[8182]), .Z(n47168) );
  XOR U47667 ( .A(n47169), .B(n47168), .Z(n47147) );
  AND U47668 ( .A(x[481]), .B(y[8183]), .Z(n47174) );
  XOR U47669 ( .A(n47175), .B(n47174), .Z(n47173) );
  AND U47670 ( .A(n46964), .B(o[503]), .Z(n47172) );
  XOR U47671 ( .A(n47173), .B(n47172), .Z(n47146) );
  XOR U47672 ( .A(n47147), .B(n47146), .Z(n47148) );
  XNOR U47673 ( .A(n47149), .B(n47148), .Z(n47200) );
  NANDN U47674 ( .A(n46966), .B(n46965), .Z(n46970) );
  NAND U47675 ( .A(n46968), .B(n46967), .Z(n46969) );
  NAND U47676 ( .A(n46970), .B(n46969), .Z(n47144) );
  AND U47677 ( .A(y[8168]), .B(x[496]), .Z(n46972) );
  NAND U47678 ( .A(y[8163]), .B(x[501]), .Z(n46971) );
  XNOR U47679 ( .A(n46972), .B(n46971), .Z(n47134) );
  AND U47680 ( .A(x[485]), .B(y[8179]), .Z(n47133) );
  XOR U47681 ( .A(n47134), .B(n47133), .Z(n47143) );
  AND U47682 ( .A(x[486]), .B(y[8178]), .Z(n47497) );
  AND U47683 ( .A(x[500]), .B(y[8164]), .Z(n47137) );
  XOR U47684 ( .A(n47497), .B(n47137), .Z(n47139) );
  AND U47685 ( .A(x[499]), .B(y[8165]), .Z(n47138) );
  XOR U47686 ( .A(n47139), .B(n47138), .Z(n47142) );
  XOR U47687 ( .A(n47143), .B(n47142), .Z(n47145) );
  XOR U47688 ( .A(n47144), .B(n47145), .Z(n47125) );
  NAND U47689 ( .A(n47252), .B(n46973), .Z(n46977) );
  NANDN U47690 ( .A(n46975), .B(n46974), .Z(n46976) );
  NAND U47691 ( .A(n46977), .B(n46976), .Z(n47123) );
  NAND U47692 ( .A(n46979), .B(n46978), .Z(n46983) );
  NAND U47693 ( .A(n46981), .B(n46980), .Z(n46982) );
  NAND U47694 ( .A(n46983), .B(n46982), .Z(n47122) );
  XOR U47695 ( .A(n47123), .B(n47122), .Z(n47124) );
  XOR U47696 ( .A(n47125), .B(n47124), .Z(n47199) );
  XOR U47697 ( .A(n47200), .B(n47199), .Z(n47202) );
  NAND U47698 ( .A(n46985), .B(n46984), .Z(n46989) );
  NAND U47699 ( .A(n46987), .B(n46986), .Z(n46988) );
  NAND U47700 ( .A(n46989), .B(n46988), .Z(n47193) );
  AND U47701 ( .A(x[483]), .B(y[8181]), .Z(n47185) );
  XOR U47702 ( .A(n47186), .B(n47185), .Z(n47188) );
  AND U47703 ( .A(x[484]), .B(y[8180]), .Z(n47187) );
  XOR U47704 ( .A(n47188), .B(n47187), .Z(n47194) );
  XOR U47705 ( .A(n47193), .B(n47194), .Z(n47196) );
  AND U47706 ( .A(y[8175]), .B(x[489]), .Z(n46991) );
  NAND U47707 ( .A(y[8174]), .B(x[490]), .Z(n46990) );
  XNOR U47708 ( .A(n46991), .B(n46990), .Z(n47158) );
  AND U47709 ( .A(y[8170]), .B(x[494]), .Z(n46993) );
  NAND U47710 ( .A(y[8176]), .B(x[488]), .Z(n46992) );
  XNOR U47711 ( .A(n46993), .B(n46992), .Z(n47162) );
  NAND U47712 ( .A(x[491]), .B(y[8173]), .Z(n47163) );
  XNOR U47713 ( .A(n47162), .B(n47163), .Z(n47157) );
  XOR U47714 ( .A(n47158), .B(n47157), .Z(n47195) );
  XOR U47715 ( .A(n47196), .B(n47195), .Z(n47201) );
  XNOR U47716 ( .A(n47202), .B(n47201), .Z(n47212) );
  NAND U47717 ( .A(n46995), .B(n46994), .Z(n46999) );
  NAND U47718 ( .A(n46997), .B(n46996), .Z(n46998) );
  AND U47719 ( .A(n46999), .B(n46998), .Z(n47211) );
  XOR U47720 ( .A(n47212), .B(n47211), .Z(n47213) );
  NAND U47721 ( .A(n47001), .B(n47000), .Z(n47005) );
  NAND U47722 ( .A(n47003), .B(n47002), .Z(n47004) );
  AND U47723 ( .A(n47005), .B(n47004), .Z(n47214) );
  XOR U47724 ( .A(n47213), .B(n47214), .Z(n47107) );
  NAND U47725 ( .A(n47007), .B(n47006), .Z(n47011) );
  NAND U47726 ( .A(n47009), .B(n47008), .Z(n47010) );
  NAND U47727 ( .A(n47011), .B(n47010), .Z(n47207) );
  NAND U47728 ( .A(n47013), .B(n47012), .Z(n47017) );
  NAND U47729 ( .A(n47015), .B(n47014), .Z(n47016) );
  NAND U47730 ( .A(n47017), .B(n47016), .Z(n47205) );
  NANDN U47731 ( .A(n47019), .B(n47018), .Z(n47023) );
  NANDN U47732 ( .A(n47021), .B(n47020), .Z(n47022) );
  NAND U47733 ( .A(n47023), .B(n47022), .Z(n47130) );
  AND U47734 ( .A(x[480]), .B(y[8184]), .Z(n47190) );
  AND U47735 ( .A(x[504]), .B(y[8160]), .Z(n47189) );
  XOR U47736 ( .A(n47190), .B(n47189), .Z(n47192) );
  AND U47737 ( .A(x[503]), .B(y[8161]), .Z(n47184) );
  XOR U47738 ( .A(n47184), .B(o[504]), .Z(n47191) );
  XOR U47739 ( .A(n47192), .B(n47191), .Z(n47129) );
  AND U47740 ( .A(x[487]), .B(y[8177]), .Z(n47179) );
  AND U47741 ( .A(x[498]), .B(y[8166]), .Z(n47178) );
  XOR U47742 ( .A(n47179), .B(n47178), .Z(n47181) );
  AND U47743 ( .A(x[497]), .B(y[8167]), .Z(n47180) );
  XOR U47744 ( .A(n47181), .B(n47180), .Z(n47128) );
  XOR U47745 ( .A(n47129), .B(n47128), .Z(n47131) );
  XOR U47746 ( .A(n47130), .B(n47131), .Z(n47119) );
  NAND U47747 ( .A(n47025), .B(n47024), .Z(n47029) );
  NAND U47748 ( .A(n47027), .B(n47026), .Z(n47028) );
  NAND U47749 ( .A(n47029), .B(n47028), .Z(n47117) );
  NAND U47750 ( .A(n47031), .B(n47030), .Z(n47035) );
  NAND U47751 ( .A(n47033), .B(n47032), .Z(n47034) );
  NAND U47752 ( .A(n47035), .B(n47034), .Z(n47116) );
  XOR U47753 ( .A(n47117), .B(n47116), .Z(n47118) );
  XOR U47754 ( .A(n47119), .B(n47118), .Z(n47206) );
  XOR U47755 ( .A(n47205), .B(n47206), .Z(n47208) );
  XNOR U47756 ( .A(n47207), .B(n47208), .Z(n47112) );
  NANDN U47757 ( .A(n47037), .B(n47036), .Z(n47041) );
  NAND U47758 ( .A(n47039), .B(n47038), .Z(n47040) );
  AND U47759 ( .A(n47041), .B(n47040), .Z(n47153) );
  NANDN U47760 ( .A(n47043), .B(n47042), .Z(n47047) );
  NANDN U47761 ( .A(n47045), .B(n47044), .Z(n47046) );
  AND U47762 ( .A(n47047), .B(n47046), .Z(n47150) );
  NANDN U47763 ( .A(n47049), .B(n47048), .Z(n47053) );
  NANDN U47764 ( .A(n47051), .B(n47050), .Z(n47052) );
  NAND U47765 ( .A(n47053), .B(n47052), .Z(n47151) );
  XOR U47766 ( .A(n47153), .B(n47152), .Z(n47110) );
  NAND U47767 ( .A(n47055), .B(n47054), .Z(n47059) );
  NANDN U47768 ( .A(n47057), .B(n47056), .Z(n47058) );
  AND U47769 ( .A(n47059), .B(n47058), .Z(n47111) );
  XOR U47770 ( .A(n47110), .B(n47111), .Z(n47113) );
  XOR U47771 ( .A(n47112), .B(n47113), .Z(n47104) );
  NAND U47772 ( .A(n47061), .B(n47060), .Z(n47065) );
  NAND U47773 ( .A(n47063), .B(n47062), .Z(n47064) );
  NAND U47774 ( .A(n47065), .B(n47064), .Z(n47105) );
  XNOR U47775 ( .A(n47107), .B(n47106), .Z(n47221) );
  NAND U47776 ( .A(n47067), .B(n47066), .Z(n47071) );
  NAND U47777 ( .A(n47069), .B(n47068), .Z(n47070) );
  AND U47778 ( .A(n47071), .B(n47070), .Z(n47101) );
  NAND U47779 ( .A(n47073), .B(n47072), .Z(n47077) );
  NAND U47780 ( .A(n47075), .B(n47074), .Z(n47076) );
  AND U47781 ( .A(n47077), .B(n47076), .Z(n47099) );
  NANDN U47782 ( .A(n47079), .B(n47078), .Z(n47083) );
  NAND U47783 ( .A(n47081), .B(n47080), .Z(n47082) );
  NAND U47784 ( .A(n47083), .B(n47082), .Z(n47098) );
  XOR U47785 ( .A(n47221), .B(n47220), .Z(n47222) );
  XNOR U47786 ( .A(n47223), .B(n47222), .Z(n47219) );
  NANDN U47787 ( .A(n47084), .B(n47085), .Z(n47090) );
  NOR U47788 ( .A(n47086), .B(n47085), .Z(n47088) );
  OR U47789 ( .A(n47088), .B(n47087), .Z(n47089) );
  AND U47790 ( .A(n47090), .B(n47089), .Z(n47217) );
  NAND U47791 ( .A(n47092), .B(n47091), .Z(n47096) );
  NAND U47792 ( .A(n47094), .B(n47093), .Z(n47095) );
  AND U47793 ( .A(n47096), .B(n47095), .Z(n47218) );
  XOR U47794 ( .A(n47217), .B(n47218), .Z(n47097) );
  XNOR U47795 ( .A(n47219), .B(n47097), .Z(N1017) );
  NANDN U47796 ( .A(n47099), .B(n47098), .Z(n47103) );
  NANDN U47797 ( .A(n47101), .B(n47100), .Z(n47102) );
  AND U47798 ( .A(n47103), .B(n47102), .Z(n47361) );
  NANDN U47799 ( .A(n47105), .B(n47104), .Z(n47109) );
  NAND U47800 ( .A(n47107), .B(n47106), .Z(n47108) );
  AND U47801 ( .A(n47109), .B(n47108), .Z(n47359) );
  NAND U47802 ( .A(n47111), .B(n47110), .Z(n47115) );
  NAND U47803 ( .A(n47113), .B(n47112), .Z(n47114) );
  AND U47804 ( .A(n47115), .B(n47114), .Z(n47236) );
  NAND U47805 ( .A(n47117), .B(n47116), .Z(n47121) );
  NAND U47806 ( .A(n47119), .B(n47118), .Z(n47120) );
  NAND U47807 ( .A(n47121), .B(n47120), .Z(n47240) );
  NAND U47808 ( .A(n47123), .B(n47122), .Z(n47127) );
  NAND U47809 ( .A(n47125), .B(n47124), .Z(n47126) );
  NAND U47810 ( .A(n47127), .B(n47126), .Z(n47239) );
  XOR U47811 ( .A(n47240), .B(n47239), .Z(n47242) );
  AND U47812 ( .A(x[501]), .B(y[8168]), .Z(n48097) );
  AND U47813 ( .A(x[502]), .B(y[8163]), .Z(n47313) );
  AND U47814 ( .A(x[485]), .B(y[8180]), .Z(n47311) );
  NAND U47815 ( .A(x[497]), .B(y[8168]), .Z(n47310) );
  XNOR U47816 ( .A(n47311), .B(n47310), .Z(n47312) );
  XOR U47817 ( .A(n47313), .B(n47312), .Z(n47338) );
  AND U47818 ( .A(y[8165]), .B(x[500]), .Z(n47136) );
  NAND U47819 ( .A(y[8164]), .B(x[501]), .Z(n47135) );
  XNOR U47820 ( .A(n47136), .B(n47135), .Z(n47324) );
  NAND U47821 ( .A(x[499]), .B(y[8166]), .Z(n47325) );
  XNOR U47822 ( .A(n47324), .B(n47325), .Z(n47339) );
  XOR U47823 ( .A(n47338), .B(n47339), .Z(n47341) );
  XNOR U47824 ( .A(n47340), .B(n47341), .Z(n47270) );
  IV U47825 ( .A(n47137), .Z(n47323) );
  NANDN U47826 ( .A(n47323), .B(n47497), .Z(n47141) );
  NAND U47827 ( .A(n47139), .B(n47138), .Z(n47140) );
  NAND U47828 ( .A(n47141), .B(n47140), .Z(n47345) );
  AND U47829 ( .A(x[495]), .B(y[8170]), .Z(n47331) );
  AND U47830 ( .A(x[498]), .B(y[8167]), .Z(n47329) );
  NAND U47831 ( .A(x[486]), .B(y[8179]), .Z(n47328) );
  XNOR U47832 ( .A(n47329), .B(n47328), .Z(n47330) );
  XOR U47833 ( .A(n47331), .B(n47330), .Z(n47342) );
  AND U47834 ( .A(x[503]), .B(y[8162]), .Z(n47306) );
  AND U47835 ( .A(x[484]), .B(y[8181]), .Z(n47305) );
  NAND U47836 ( .A(x[496]), .B(y[8169]), .Z(n47304) );
  XOR U47837 ( .A(n47305), .B(n47304), .Z(n47307) );
  XNOR U47838 ( .A(n47306), .B(n47307), .Z(n47343) );
  XOR U47839 ( .A(n47342), .B(n47343), .Z(n47344) );
  XNOR U47840 ( .A(n47345), .B(n47344), .Z(n47269) );
  XNOR U47841 ( .A(n47270), .B(n47269), .Z(n47272) );
  XNOR U47842 ( .A(n47271), .B(n47272), .Z(n47282) );
  XOR U47843 ( .A(n47279), .B(n47280), .Z(n47281) );
  XNOR U47844 ( .A(n47282), .B(n47281), .Z(n47241) );
  XOR U47845 ( .A(n47242), .B(n47241), .Z(n47234) );
  NANDN U47846 ( .A(n47151), .B(n47150), .Z(n47155) );
  NAND U47847 ( .A(n47153), .B(n47152), .Z(n47154) );
  NAND U47848 ( .A(n47155), .B(n47154), .Z(n47233) );
  NANDN U47849 ( .A(n47251), .B(n47156), .Z(n47160) );
  NAND U47850 ( .A(n47158), .B(n47157), .Z(n47159) );
  NAND U47851 ( .A(n47160), .B(n47159), .Z(n47275) );
  AND U47852 ( .A(x[494]), .B(y[8176]), .Z(n48173) );
  NAND U47853 ( .A(n48173), .B(n47161), .Z(n47165) );
  NANDN U47854 ( .A(n47163), .B(n47162), .Z(n47164) );
  AND U47855 ( .A(n47165), .B(n47164), .Z(n47301) );
  AND U47856 ( .A(x[491]), .B(y[8174]), .Z(n47320) );
  AND U47857 ( .A(x[492]), .B(y[8173]), .Z(n47318) );
  NAND U47858 ( .A(x[487]), .B(y[8178]), .Z(n47317) );
  XNOR U47859 ( .A(n47318), .B(n47317), .Z(n47319) );
  XNOR U47860 ( .A(n47320), .B(n47319), .Z(n47299) );
  NAND U47861 ( .A(x[504]), .B(y[8161]), .Z(n47316) );
  XNOR U47862 ( .A(o[505]), .B(n47316), .Z(n47286) );
  NAND U47863 ( .A(x[481]), .B(y[8184]), .Z(n47287) );
  XNOR U47864 ( .A(n47286), .B(n47287), .Z(n47288) );
  NAND U47865 ( .A(x[493]), .B(y[8172]), .Z(n47289) );
  XNOR U47866 ( .A(n47288), .B(n47289), .Z(n47298) );
  XNOR U47867 ( .A(n47299), .B(n47298), .Z(n47300) );
  XNOR U47868 ( .A(n47301), .B(n47300), .Z(n47276) );
  XOR U47869 ( .A(n47275), .B(n47276), .Z(n47278) );
  AND U47870 ( .A(n47167), .B(n47166), .Z(n47171) );
  NAND U47871 ( .A(n47169), .B(n47168), .Z(n47170) );
  NANDN U47872 ( .A(n47171), .B(n47170), .Z(n47264) );
  AND U47873 ( .A(n47173), .B(n47172), .Z(n47177) );
  NAND U47874 ( .A(n47175), .B(n47174), .Z(n47176) );
  NANDN U47875 ( .A(n47177), .B(n47176), .Z(n47263) );
  XOR U47876 ( .A(n47264), .B(n47263), .Z(n47266) );
  NAND U47877 ( .A(n47179), .B(n47178), .Z(n47183) );
  NAND U47878 ( .A(n47181), .B(n47180), .Z(n47182) );
  NAND U47879 ( .A(n47183), .B(n47182), .Z(n47259) );
  AND U47880 ( .A(x[488]), .B(y[8177]), .Z(n47254) );
  XNOR U47881 ( .A(n47252), .B(n47251), .Z(n47253) );
  XOR U47882 ( .A(n47254), .B(n47253), .Z(n47258) );
  AND U47883 ( .A(n47184), .B(o[504]), .Z(n47247) );
  AND U47884 ( .A(x[505]), .B(y[8160]), .Z(n47246) );
  NAND U47885 ( .A(x[480]), .B(y[8185]), .Z(n47245) );
  XOR U47886 ( .A(n47246), .B(n47245), .Z(n47248) );
  XNOR U47887 ( .A(n47247), .B(n47248), .Z(n47257) );
  XOR U47888 ( .A(n47258), .B(n47257), .Z(n47260) );
  XOR U47889 ( .A(n47259), .B(n47260), .Z(n47265) );
  XOR U47890 ( .A(n47266), .B(n47265), .Z(n47277) );
  XOR U47891 ( .A(n47278), .B(n47277), .Z(n47355) );
  AND U47892 ( .A(x[494]), .B(y[8171]), .Z(n47292) );
  NAND U47893 ( .A(x[482]), .B(y[8183]), .Z(n47293) );
  XNOR U47894 ( .A(n47292), .B(n47293), .Z(n47294) );
  NAND U47895 ( .A(x[483]), .B(y[8182]), .Z(n47295) );
  XNOR U47896 ( .A(n47294), .B(n47295), .Z(n47335) );
  XOR U47897 ( .A(n47334), .B(n47335), .Z(n47337) );
  XOR U47898 ( .A(n47336), .B(n47337), .Z(n47353) );
  NAND U47899 ( .A(n47194), .B(n47193), .Z(n47198) );
  NAND U47900 ( .A(n47196), .B(n47195), .Z(n47197) );
  AND U47901 ( .A(n47198), .B(n47197), .Z(n47352) );
  NAND U47902 ( .A(n47200), .B(n47199), .Z(n47204) );
  NAND U47903 ( .A(n47202), .B(n47201), .Z(n47203) );
  AND U47904 ( .A(n47204), .B(n47203), .Z(n47346) );
  XOR U47905 ( .A(n47347), .B(n47346), .Z(n47349) );
  NAND U47906 ( .A(n47206), .B(n47205), .Z(n47210) );
  NAND U47907 ( .A(n47208), .B(n47207), .Z(n47209) );
  AND U47908 ( .A(n47210), .B(n47209), .Z(n47348) );
  XNOR U47909 ( .A(n47349), .B(n47348), .Z(n47228) );
  NAND U47910 ( .A(n47212), .B(n47211), .Z(n47216) );
  NAND U47911 ( .A(n47214), .B(n47213), .Z(n47215) );
  AND U47912 ( .A(n47216), .B(n47215), .Z(n47227) );
  XOR U47913 ( .A(n47228), .B(n47227), .Z(n47230) );
  XNOR U47914 ( .A(n47229), .B(n47230), .Z(n47358) );
  XNOR U47915 ( .A(n47361), .B(n47360), .Z(n47367) );
  NAND U47916 ( .A(n47221), .B(n47220), .Z(n47225) );
  NAND U47917 ( .A(n47223), .B(n47222), .Z(n47224) );
  AND U47918 ( .A(n47225), .B(n47224), .Z(n47366) );
  IV U47919 ( .A(n47366), .Z(n47364) );
  XOR U47920 ( .A(n47365), .B(n47364), .Z(n47226) );
  XNOR U47921 ( .A(n47367), .B(n47226), .Z(N1018) );
  NAND U47922 ( .A(n47228), .B(n47227), .Z(n47232) );
  NAND U47923 ( .A(n47230), .B(n47229), .Z(n47231) );
  NAND U47924 ( .A(n47232), .B(n47231), .Z(n47514) );
  NANDN U47925 ( .A(n47234), .B(n47233), .Z(n47238) );
  NANDN U47926 ( .A(n47236), .B(n47235), .Z(n47237) );
  AND U47927 ( .A(n47238), .B(n47237), .Z(n47513) );
  XOR U47928 ( .A(n47514), .B(n47513), .Z(n47516) );
  NAND U47929 ( .A(n47240), .B(n47239), .Z(n47244) );
  NAND U47930 ( .A(n47242), .B(n47241), .Z(n47243) );
  NAND U47931 ( .A(n47244), .B(n47243), .Z(n47380) );
  AND U47932 ( .A(x[482]), .B(y[8184]), .Z(n47438) );
  XOR U47933 ( .A(n47439), .B(n47438), .Z(n47441) );
  NAND U47934 ( .A(x[504]), .B(y[8162]), .Z(n47440) );
  XNOR U47935 ( .A(n47441), .B(n47440), .Z(n47394) );
  NANDN U47936 ( .A(n47246), .B(n47245), .Z(n47250) );
  OR U47937 ( .A(n47248), .B(n47247), .Z(n47249) );
  NAND U47938 ( .A(n47250), .B(n47249), .Z(n47395) );
  XNOR U47939 ( .A(n47394), .B(n47395), .Z(n47396) );
  NANDN U47940 ( .A(n47252), .B(n47251), .Z(n47256) );
  NANDN U47941 ( .A(n47254), .B(n47253), .Z(n47255) );
  NAND U47942 ( .A(n47256), .B(n47255), .Z(n47397) );
  XOR U47943 ( .A(n47396), .B(n47397), .Z(n47468) );
  NAND U47944 ( .A(n47258), .B(n47257), .Z(n47262) );
  NAND U47945 ( .A(n47260), .B(n47259), .Z(n47261) );
  AND U47946 ( .A(n47262), .B(n47261), .Z(n47469) );
  XOR U47947 ( .A(n47468), .B(n47469), .Z(n47471) );
  NAND U47948 ( .A(n47264), .B(n47263), .Z(n47268) );
  NAND U47949 ( .A(n47266), .B(n47265), .Z(n47267) );
  AND U47950 ( .A(n47268), .B(n47267), .Z(n47470) );
  XOR U47951 ( .A(n47471), .B(n47470), .Z(n47511) );
  NAND U47952 ( .A(n47270), .B(n47269), .Z(n47274) );
  NANDN U47953 ( .A(n47272), .B(n47271), .Z(n47273) );
  NAND U47954 ( .A(n47274), .B(n47273), .Z(n47510) );
  XNOR U47955 ( .A(n47510), .B(n47509), .Z(n47512) );
  XOR U47956 ( .A(n47511), .B(n47512), .Z(n47378) );
  AND U47957 ( .A(y[8180]), .B(x[486]), .Z(n47284) );
  NAND U47958 ( .A(y[8178]), .B(x[488]), .Z(n47283) );
  XNOR U47959 ( .A(n47284), .B(n47283), .Z(n47498) );
  NAND U47960 ( .A(x[489]), .B(y[8177]), .Z(n47499) );
  XOR U47961 ( .A(n47498), .B(n47499), .Z(n47474) );
  AND U47962 ( .A(x[492]), .B(y[8174]), .Z(n47553) );
  AND U47963 ( .A(x[485]), .B(y[8181]), .Z(n47409) );
  XOR U47964 ( .A(n47553), .B(n47409), .Z(n47411) );
  NAND U47965 ( .A(x[490]), .B(y[8176]), .Z(n47410) );
  XNOR U47966 ( .A(n47411), .B(n47410), .Z(n47476) );
  AND U47967 ( .A(x[487]), .B(y[8179]), .Z(n47475) );
  XNOR U47968 ( .A(n47476), .B(n47475), .Z(n47285) );
  XOR U47969 ( .A(n47474), .B(n47285), .Z(n47464) );
  NANDN U47970 ( .A(n47287), .B(n47286), .Z(n47291) );
  NANDN U47971 ( .A(n47289), .B(n47288), .Z(n47290) );
  AND U47972 ( .A(n47291), .B(n47290), .Z(n47463) );
  NANDN U47973 ( .A(n47293), .B(n47292), .Z(n47297) );
  NANDN U47974 ( .A(n47295), .B(n47294), .Z(n47296) );
  NAND U47975 ( .A(n47297), .B(n47296), .Z(n47462) );
  XOR U47976 ( .A(n47463), .B(n47462), .Z(n47465) );
  XNOR U47977 ( .A(n47464), .B(n47465), .Z(n47421) );
  NANDN U47978 ( .A(n47299), .B(n47298), .Z(n47303) );
  NANDN U47979 ( .A(n47301), .B(n47300), .Z(n47302) );
  AND U47980 ( .A(n47303), .B(n47302), .Z(n47420) );
  XNOR U47981 ( .A(n47421), .B(n47420), .Z(n47422) );
  NANDN U47982 ( .A(n47305), .B(n47304), .Z(n47309) );
  OR U47983 ( .A(n47307), .B(n47306), .Z(n47308) );
  AND U47984 ( .A(n47309), .B(n47308), .Z(n47426) );
  NANDN U47985 ( .A(n47311), .B(n47310), .Z(n47315) );
  NANDN U47986 ( .A(n47313), .B(n47312), .Z(n47314) );
  NAND U47987 ( .A(n47315), .B(n47314), .Z(n47427) );
  XNOR U47988 ( .A(n47426), .B(n47427), .Z(n47428) );
  ANDN U47989 ( .B(o[505]), .A(n47316), .Z(n47491) );
  NAND U47990 ( .A(x[494]), .B(y[8172]), .Z(n47492) );
  XNOR U47991 ( .A(n47491), .B(n47492), .Z(n47493) );
  NAND U47992 ( .A(x[481]), .B(y[8185]), .Z(n47494) );
  XNOR U47993 ( .A(n47493), .B(n47494), .Z(n47400) );
  NAND U47994 ( .A(x[505]), .B(y[8161]), .Z(n47502) );
  XNOR U47995 ( .A(o[506]), .B(n47502), .Z(n47414) );
  NAND U47996 ( .A(x[506]), .B(y[8160]), .Z(n47415) );
  XNOR U47997 ( .A(n47414), .B(n47415), .Z(n47416) );
  NAND U47998 ( .A(x[480]), .B(y[8186]), .Z(n47417) );
  XOR U47999 ( .A(n47416), .B(n47417), .Z(n47401) );
  NANDN U48000 ( .A(n47318), .B(n47317), .Z(n47322) );
  NANDN U48001 ( .A(n47320), .B(n47319), .Z(n47321) );
  NAND U48002 ( .A(n47322), .B(n47321), .Z(n47403) );
  XNOR U48003 ( .A(n47428), .B(n47429), .Z(n47390) );
  AND U48004 ( .A(x[501]), .B(y[8165]), .Z(n47485) );
  NANDN U48005 ( .A(n47323), .B(n47485), .Z(n47327) );
  NANDN U48006 ( .A(n47325), .B(n47324), .Z(n47326) );
  AND U48007 ( .A(n47327), .B(n47326), .Z(n47459) );
  XOR U48008 ( .A(n47486), .B(n47485), .Z(n47488) );
  NAND U48009 ( .A(x[500]), .B(y[8166]), .Z(n47487) );
  XNOR U48010 ( .A(n47488), .B(n47487), .Z(n47456) );
  NAND U48011 ( .A(x[503]), .B(y[8163]), .Z(n47445) );
  XNOR U48012 ( .A(n47444), .B(n47445), .Z(n47447) );
  AND U48013 ( .A(x[502]), .B(y[8164]), .Z(n47446) );
  XNOR U48014 ( .A(n47447), .B(n47446), .Z(n47457) );
  XNOR U48015 ( .A(n47456), .B(n47457), .Z(n47458) );
  XNOR U48016 ( .A(n47459), .B(n47458), .Z(n47389) );
  AND U48017 ( .A(x[484]), .B(y[8182]), .Z(n47450) );
  XOR U48018 ( .A(n47451), .B(n47450), .Z(n47453) );
  AND U48019 ( .A(x[491]), .B(y[8175]), .Z(n47477) );
  NAND U48020 ( .A(x[499]), .B(y[8167]), .Z(n47478) );
  XNOR U48021 ( .A(n47477), .B(n47478), .Z(n47479) );
  NAND U48022 ( .A(x[483]), .B(y[8183]), .Z(n47480) );
  XOR U48023 ( .A(n47479), .B(n47480), .Z(n47433) );
  XNOR U48024 ( .A(n47432), .B(n47433), .Z(n47434) );
  NANDN U48025 ( .A(n47329), .B(n47328), .Z(n47333) );
  NANDN U48026 ( .A(n47331), .B(n47330), .Z(n47332) );
  NAND U48027 ( .A(n47333), .B(n47332), .Z(n47435) );
  XOR U48028 ( .A(n47434), .B(n47435), .Z(n47388) );
  XOR U48029 ( .A(n47389), .B(n47388), .Z(n47391) );
  XNOR U48030 ( .A(n47390), .B(n47391), .Z(n47423) );
  XNOR U48031 ( .A(n47422), .B(n47423), .Z(n47385) );
  XOR U48032 ( .A(n47504), .B(n47503), .Z(n47506) );
  XOR U48033 ( .A(n47505), .B(n47506), .Z(n47384) );
  XNOR U48034 ( .A(n47385), .B(n47384), .Z(n47387) );
  XOR U48035 ( .A(n47386), .B(n47387), .Z(n47379) );
  XOR U48036 ( .A(n47378), .B(n47379), .Z(n47381) );
  XOR U48037 ( .A(n47380), .B(n47381), .Z(n47375) );
  NAND U48038 ( .A(n47347), .B(n47346), .Z(n47351) );
  NAND U48039 ( .A(n47349), .B(n47348), .Z(n47350) );
  AND U48040 ( .A(n47351), .B(n47350), .Z(n47373) );
  NANDN U48041 ( .A(n47353), .B(n47352), .Z(n47357) );
  NANDN U48042 ( .A(n47355), .B(n47354), .Z(n47356) );
  AND U48043 ( .A(n47357), .B(n47356), .Z(n47372) );
  XOR U48044 ( .A(n47373), .B(n47372), .Z(n47374) );
  XOR U48045 ( .A(n47375), .B(n47374), .Z(n47515) );
  XOR U48046 ( .A(n47516), .B(n47515), .Z(n47521) );
  NANDN U48047 ( .A(n47359), .B(n47358), .Z(n47363) );
  NAND U48048 ( .A(n47361), .B(n47360), .Z(n47362) );
  NAND U48049 ( .A(n47363), .B(n47362), .Z(n47519) );
  NANDN U48050 ( .A(n47364), .B(n47365), .Z(n47370) );
  NOR U48051 ( .A(n47366), .B(n47365), .Z(n47368) );
  OR U48052 ( .A(n47368), .B(n47367), .Z(n47369) );
  AND U48053 ( .A(n47370), .B(n47369), .Z(n47520) );
  XOR U48054 ( .A(n47519), .B(n47520), .Z(n47371) );
  XNOR U48055 ( .A(n47521), .B(n47371), .Z(N1019) );
  NAND U48056 ( .A(n47373), .B(n47372), .Z(n47377) );
  NAND U48057 ( .A(n47375), .B(n47374), .Z(n47376) );
  NAND U48058 ( .A(n47377), .B(n47376), .Z(n47671) );
  NAND U48059 ( .A(n47379), .B(n47378), .Z(n47383) );
  NAND U48060 ( .A(n47381), .B(n47380), .Z(n47382) );
  NAND U48061 ( .A(n47383), .B(n47382), .Z(n47669) );
  NANDN U48062 ( .A(n47389), .B(n47388), .Z(n47393) );
  OR U48063 ( .A(n47391), .B(n47390), .Z(n47392) );
  AND U48064 ( .A(n47393), .B(n47392), .Z(n47648) );
  NANDN U48065 ( .A(n47395), .B(n47394), .Z(n47399) );
  NANDN U48066 ( .A(n47397), .B(n47396), .Z(n47398) );
  AND U48067 ( .A(n47399), .B(n47398), .Z(n47639) );
  NANDN U48068 ( .A(n47401), .B(n47400), .Z(n47405) );
  NANDN U48069 ( .A(n47403), .B(n47402), .Z(n47404) );
  AND U48070 ( .A(n47405), .B(n47404), .Z(n47637) );
  AND U48071 ( .A(x[486]), .B(y[8181]), .Z(n47613) );
  AND U48072 ( .A(x[499]), .B(y[8168]), .Z(n47611) );
  NAND U48073 ( .A(x[505]), .B(y[8162]), .Z(n47612) );
  XOR U48074 ( .A(n47611), .B(n47612), .Z(n47614) );
  XNOR U48075 ( .A(n47613), .B(n47614), .Z(n47602) );
  AND U48076 ( .A(x[495]), .B(y[8172]), .Z(n47562) );
  NAND U48077 ( .A(x[482]), .B(y[8185]), .Z(n47563) );
  XNOR U48078 ( .A(n47562), .B(n47563), .Z(n47564) );
  NAND U48079 ( .A(x[483]), .B(y[8184]), .Z(n47565) );
  XOR U48080 ( .A(n47564), .B(n47565), .Z(n47603) );
  XNOR U48081 ( .A(n47602), .B(n47603), .Z(n47605) );
  AND U48082 ( .A(x[496]), .B(y[8171]), .Z(n47542) );
  XOR U48083 ( .A(n47542), .B(n47406), .Z(n47543) );
  XOR U48084 ( .A(n47544), .B(n47543), .Z(n47554) );
  AND U48085 ( .A(y[8174]), .B(x[493]), .Z(n47408) );
  NAND U48086 ( .A(y[8175]), .B(x[492]), .Z(n47407) );
  XNOR U48087 ( .A(n47408), .B(n47407), .Z(n47555) );
  XOR U48088 ( .A(n47554), .B(n47555), .Z(n47604) );
  XOR U48089 ( .A(n47605), .B(n47604), .Z(n47570) );
  NAND U48090 ( .A(n47553), .B(n47409), .Z(n47413) );
  ANDN U48091 ( .B(n47411), .A(n47410), .Z(n47412) );
  ANDN U48092 ( .B(n47413), .A(n47412), .Z(n47569) );
  NANDN U48093 ( .A(n47415), .B(n47414), .Z(n47419) );
  NANDN U48094 ( .A(n47417), .B(n47416), .Z(n47418) );
  NAND U48095 ( .A(n47419), .B(n47418), .Z(n47568) );
  XOR U48096 ( .A(n47569), .B(n47568), .Z(n47571) );
  XNOR U48097 ( .A(n47570), .B(n47571), .Z(n47636) );
  XNOR U48098 ( .A(n47648), .B(n47649), .Z(n47651) );
  NANDN U48099 ( .A(n47421), .B(n47420), .Z(n47425) );
  NANDN U48100 ( .A(n47423), .B(n47422), .Z(n47424) );
  AND U48101 ( .A(n47425), .B(n47424), .Z(n47650) );
  XOR U48102 ( .A(n47651), .B(n47650), .Z(n47529) );
  NANDN U48103 ( .A(n47427), .B(n47426), .Z(n47431) );
  NANDN U48104 ( .A(n47429), .B(n47428), .Z(n47430) );
  AND U48105 ( .A(n47431), .B(n47430), .Z(n47645) );
  NANDN U48106 ( .A(n47433), .B(n47432), .Z(n47437) );
  NANDN U48107 ( .A(n47435), .B(n47434), .Z(n47436) );
  AND U48108 ( .A(n47437), .B(n47436), .Z(n47643) );
  NAND U48109 ( .A(n47439), .B(n47438), .Z(n47443) );
  ANDN U48110 ( .B(n47441), .A(n47440), .Z(n47442) );
  ANDN U48111 ( .B(n47443), .A(n47442), .Z(n47575) );
  NANDN U48112 ( .A(n47445), .B(n47444), .Z(n47449) );
  NAND U48113 ( .A(n47447), .B(n47446), .Z(n47448) );
  NAND U48114 ( .A(n47449), .B(n47448), .Z(n47574) );
  XNOR U48115 ( .A(n47575), .B(n47574), .Z(n47576) );
  NAND U48116 ( .A(n47451), .B(n47450), .Z(n47455) );
  ANDN U48117 ( .B(n47453), .A(n47452), .Z(n47454) );
  ANDN U48118 ( .B(n47455), .A(n47454), .Z(n47589) );
  AND U48119 ( .A(x[480]), .B(y[8187]), .Z(n47632) );
  NAND U48120 ( .A(x[507]), .B(y[8160]), .Z(n47633) );
  XNOR U48121 ( .A(n47632), .B(n47633), .Z(n47635) );
  AND U48122 ( .A(x[506]), .B(y[8161]), .Z(n47623) );
  XOR U48123 ( .A(o[507]), .B(n47623), .Z(n47634) );
  XOR U48124 ( .A(n47635), .B(n47634), .Z(n47586) );
  AND U48125 ( .A(x[489]), .B(y[8178]), .Z(n47617) );
  NAND U48126 ( .A(x[501]), .B(y[8166]), .Z(n47618) );
  XNOR U48127 ( .A(n47617), .B(n47618), .Z(n47619) );
  NAND U48128 ( .A(x[498]), .B(y[8169]), .Z(n47620) );
  XOR U48129 ( .A(n47619), .B(n47620), .Z(n47587) );
  XNOR U48130 ( .A(n47586), .B(n47587), .Z(n47588) );
  XOR U48131 ( .A(n47589), .B(n47588), .Z(n47577) );
  XNOR U48132 ( .A(n47576), .B(n47577), .Z(n47642) );
  NANDN U48133 ( .A(n47457), .B(n47456), .Z(n47461) );
  NANDN U48134 ( .A(n47459), .B(n47458), .Z(n47460) );
  AND U48135 ( .A(n47461), .B(n47460), .Z(n47655) );
  NANDN U48136 ( .A(n47463), .B(n47462), .Z(n47467) );
  NANDN U48137 ( .A(n47465), .B(n47464), .Z(n47466) );
  AND U48138 ( .A(n47467), .B(n47466), .Z(n47654) );
  XOR U48139 ( .A(n47655), .B(n47654), .Z(n47656) );
  XNOR U48140 ( .A(n47529), .B(n47530), .Z(n47532) );
  XNOR U48141 ( .A(n47531), .B(n47532), .Z(n47525) );
  NAND U48142 ( .A(n47469), .B(n47468), .Z(n47473) );
  NAND U48143 ( .A(n47471), .B(n47470), .Z(n47472) );
  NAND U48144 ( .A(n47473), .B(n47472), .Z(n47535) );
  NANDN U48145 ( .A(n47478), .B(n47477), .Z(n47482) );
  NANDN U48146 ( .A(n47480), .B(n47479), .Z(n47481) );
  AND U48147 ( .A(n47482), .B(n47481), .Z(n47601) );
  AND U48148 ( .A(x[487]), .B(y[8180]), .Z(n47607) );
  AND U48149 ( .A(y[8163]), .B(x[504]), .Z(n47484) );
  NAND U48150 ( .A(y[8167]), .B(x[500]), .Z(n47483) );
  XOR U48151 ( .A(n47484), .B(n47483), .Z(n47608) );
  XNOR U48152 ( .A(n47607), .B(n47608), .Z(n47599) );
  AND U48153 ( .A(x[502]), .B(y[8165]), .Z(n47550) );
  AND U48154 ( .A(x[488]), .B(y[8179]), .Z(n47547) );
  NAND U48155 ( .A(x[503]), .B(y[8164]), .Z(n47548) );
  XOR U48156 ( .A(n47550), .B(n47549), .Z(n47598) );
  XOR U48157 ( .A(n47599), .B(n47598), .Z(n47600) );
  XOR U48158 ( .A(n47601), .B(n47600), .Z(n47661) );
  NAND U48159 ( .A(n47486), .B(n47485), .Z(n47490) );
  ANDN U48160 ( .B(n47488), .A(n47487), .Z(n47489) );
  ANDN U48161 ( .B(n47490), .A(n47489), .Z(n47593) );
  NANDN U48162 ( .A(n47492), .B(n47491), .Z(n47496) );
  NANDN U48163 ( .A(n47494), .B(n47493), .Z(n47495) );
  NAND U48164 ( .A(n47496), .B(n47495), .Z(n47592) );
  XNOR U48165 ( .A(n47593), .B(n47592), .Z(n47595) );
  AND U48166 ( .A(x[488]), .B(y[8180]), .Z(n47625) );
  NAND U48167 ( .A(n47497), .B(n47625), .Z(n47501) );
  NANDN U48168 ( .A(n47499), .B(n47498), .Z(n47500) );
  NAND U48169 ( .A(n47501), .B(n47500), .Z(n47582) );
  ANDN U48170 ( .B(o[506]), .A(n47502), .Z(n47558) );
  AND U48171 ( .A(x[481]), .B(y[8186]), .Z(n47556) );
  NAND U48172 ( .A(x[494]), .B(y[8173]), .Z(n47557) );
  XOR U48173 ( .A(n47556), .B(n47557), .Z(n47559) );
  XNOR U48174 ( .A(n47558), .B(n47559), .Z(n47581) );
  AND U48175 ( .A(x[497]), .B(y[8170]), .Z(n47626) );
  NAND U48176 ( .A(x[484]), .B(y[8183]), .Z(n47627) );
  XNOR U48177 ( .A(n47626), .B(n47627), .Z(n47629) );
  AND U48178 ( .A(x[485]), .B(y[8182]), .Z(n47628) );
  XOR U48179 ( .A(n47629), .B(n47628), .Z(n47580) );
  XOR U48180 ( .A(n47581), .B(n47580), .Z(n47583) );
  XOR U48181 ( .A(n47582), .B(n47583), .Z(n47594) );
  XNOR U48182 ( .A(n47595), .B(n47594), .Z(n47660) );
  XOR U48183 ( .A(n47661), .B(n47660), .Z(n47662) );
  XNOR U48184 ( .A(n47663), .B(n47662), .Z(n47536) );
  XOR U48185 ( .A(n47535), .B(n47536), .Z(n47538) );
  NAND U48186 ( .A(n47504), .B(n47503), .Z(n47508) );
  NAND U48187 ( .A(n47506), .B(n47505), .Z(n47507) );
  AND U48188 ( .A(n47508), .B(n47507), .Z(n47537) );
  XOR U48189 ( .A(n47538), .B(n47537), .Z(n47524) );
  XOR U48190 ( .A(n47524), .B(n47523), .Z(n47526) );
  XOR U48191 ( .A(n47525), .B(n47526), .Z(n47670) );
  XNOR U48192 ( .A(n47669), .B(n47670), .Z(n47672) );
  XOR U48193 ( .A(n47671), .B(n47672), .Z(n47668) );
  NAND U48194 ( .A(n47514), .B(n47513), .Z(n47518) );
  NAND U48195 ( .A(n47516), .B(n47515), .Z(n47517) );
  NAND U48196 ( .A(n47518), .B(n47517), .Z(n47667) );
  XOR U48197 ( .A(n47667), .B(n47666), .Z(n47522) );
  XNOR U48198 ( .A(n47668), .B(n47522), .Z(N1020) );
  NANDN U48199 ( .A(n47524), .B(n47523), .Z(n47528) );
  OR U48200 ( .A(n47526), .B(n47525), .Z(n47527) );
  NAND U48201 ( .A(n47528), .B(n47527), .Z(n47676) );
  OR U48202 ( .A(n47530), .B(n47529), .Z(n47534) );
  NANDN U48203 ( .A(n47532), .B(n47531), .Z(n47533) );
  AND U48204 ( .A(n47534), .B(n47533), .Z(n47677) );
  XOR U48205 ( .A(n47676), .B(n47677), .Z(n47679) );
  NAND U48206 ( .A(n47536), .B(n47535), .Z(n47540) );
  NAND U48207 ( .A(n47538), .B(n47537), .Z(n47539) );
  AND U48208 ( .A(n47540), .B(n47539), .Z(n47683) );
  NANDN U48209 ( .A(n47542), .B(n47541), .Z(n47546) );
  NANDN U48210 ( .A(n47544), .B(n47543), .Z(n47545) );
  AND U48211 ( .A(n47546), .B(n47545), .Z(n47776) );
  AND U48212 ( .A(x[487]), .B(y[8181]), .Z(n47743) );
  AND U48213 ( .A(x[492]), .B(y[8176]), .Z(n47742) );
  XOR U48214 ( .A(n47743), .B(n47742), .Z(n47745) );
  AND U48215 ( .A(x[491]), .B(y[8177]), .Z(n47744) );
  XOR U48216 ( .A(n47745), .B(n47744), .Z(n47775) );
  AND U48217 ( .A(x[495]), .B(y[8173]), .Z(n47769) );
  AND U48218 ( .A(x[507]), .B(y[8161]), .Z(n47759) );
  XOR U48219 ( .A(o[508]), .B(n47759), .Z(n47766) );
  NAND U48220 ( .A(x[506]), .B(y[8162]), .Z(n47767) );
  XNOR U48221 ( .A(n47766), .B(n47767), .Z(n47768) );
  XNOR U48222 ( .A(n47769), .B(n47768), .Z(n47774) );
  XOR U48223 ( .A(n47775), .B(n47774), .Z(n47777) );
  XOR U48224 ( .A(n47776), .B(n47777), .Z(n47817) );
  NANDN U48225 ( .A(n47548), .B(n47547), .Z(n47552) );
  NAND U48226 ( .A(n47550), .B(n47549), .Z(n47551) );
  AND U48227 ( .A(n47552), .B(n47551), .Z(n47727) );
  AND U48228 ( .A(x[497]), .B(y[8171]), .Z(n47706) );
  AND U48229 ( .A(x[502]), .B(y[8166]), .Z(n47705) );
  XOR U48230 ( .A(n47706), .B(n47705), .Z(n47708) );
  AND U48231 ( .A(x[484]), .B(y[8184]), .Z(n47707) );
  XOR U48232 ( .A(n47708), .B(n47707), .Z(n47725) );
  AND U48233 ( .A(x[486]), .B(y[8182]), .Z(n47902) );
  NAND U48234 ( .A(x[499]), .B(y[8169]), .Z(n47748) );
  XNOR U48235 ( .A(n47902), .B(n47748), .Z(n47749) );
  XOR U48236 ( .A(n47725), .B(n47724), .Z(n47726) );
  XNOR U48237 ( .A(n47817), .B(n47816), .Z(n47818) );
  NANDN U48238 ( .A(n47557), .B(n47556), .Z(n47561) );
  NANDN U48239 ( .A(n47559), .B(n47558), .Z(n47560) );
  AND U48240 ( .A(n47561), .B(n47560), .Z(n47719) );
  NANDN U48241 ( .A(n47563), .B(n47562), .Z(n47567) );
  NANDN U48242 ( .A(n47565), .B(n47564), .Z(n47566) );
  NAND U48243 ( .A(n47567), .B(n47566), .Z(n47718) );
  XNOR U48244 ( .A(n47719), .B(n47718), .Z(n47720) );
  XOR U48245 ( .A(n47721), .B(n47720), .Z(n47819) );
  XNOR U48246 ( .A(n47818), .B(n47819), .Z(n47697) );
  NANDN U48247 ( .A(n47569), .B(n47568), .Z(n47573) );
  NANDN U48248 ( .A(n47571), .B(n47570), .Z(n47572) );
  AND U48249 ( .A(n47573), .B(n47572), .Z(n47696) );
  NANDN U48250 ( .A(n47575), .B(n47574), .Z(n47579) );
  NANDN U48251 ( .A(n47577), .B(n47576), .Z(n47578) );
  AND U48252 ( .A(n47579), .B(n47578), .Z(n47795) );
  NAND U48253 ( .A(n47581), .B(n47580), .Z(n47585) );
  NAND U48254 ( .A(n47583), .B(n47582), .Z(n47584) );
  AND U48255 ( .A(n47585), .B(n47584), .Z(n47793) );
  NANDN U48256 ( .A(n47587), .B(n47586), .Z(n47591) );
  NANDN U48257 ( .A(n47589), .B(n47588), .Z(n47590) );
  NAND U48258 ( .A(n47591), .B(n47590), .Z(n47792) );
  XNOR U48259 ( .A(n47793), .B(n47792), .Z(n47794) );
  XNOR U48260 ( .A(n47795), .B(n47794), .Z(n47695) );
  XOR U48261 ( .A(n47696), .B(n47695), .Z(n47698) );
  XOR U48262 ( .A(n47697), .B(n47698), .Z(n47824) );
  NANDN U48263 ( .A(n47593), .B(n47592), .Z(n47597) );
  NAND U48264 ( .A(n47595), .B(n47594), .Z(n47596) );
  AND U48265 ( .A(n47597), .B(n47596), .Z(n47783) );
  XNOR U48266 ( .A(n47781), .B(n47780), .Z(n47782) );
  XOR U48267 ( .A(n47783), .B(n47782), .Z(n47822) );
  AND U48268 ( .A(x[504]), .B(y[8167]), .Z(n48108) );
  AND U48269 ( .A(x[500]), .B(y[8163]), .Z(n47606) );
  NAND U48270 ( .A(n48108), .B(n47606), .Z(n47610) );
  NANDN U48271 ( .A(n47608), .B(n47607), .Z(n47609) );
  AND U48272 ( .A(n47610), .B(n47609), .Z(n47806) );
  AND U48273 ( .A(x[505]), .B(y[8163]), .Z(n47738) );
  XOR U48274 ( .A(n47739), .B(n47738), .Z(n47737) );
  NAND U48275 ( .A(x[481]), .B(y[8187]), .Z(n47736) );
  XNOR U48276 ( .A(n47737), .B(n47736), .Z(n47804) );
  AND U48277 ( .A(x[496]), .B(y[8172]), .Z(n47730) );
  NAND U48278 ( .A(x[504]), .B(y[8164]), .Z(n47731) );
  XNOR U48279 ( .A(n47730), .B(n47731), .Z(n47732) );
  NAND U48280 ( .A(x[482]), .B(y[8186]), .Z(n47733) );
  XOR U48281 ( .A(n47732), .B(n47733), .Z(n47805) );
  XOR U48282 ( .A(n47804), .B(n47805), .Z(n47807) );
  XOR U48283 ( .A(n47806), .B(n47807), .Z(n47788) );
  NANDN U48284 ( .A(n47612), .B(n47611), .Z(n47616) );
  NANDN U48285 ( .A(n47614), .B(n47613), .Z(n47615) );
  AND U48286 ( .A(n47616), .B(n47615), .Z(n47812) );
  NAND U48287 ( .A(x[483]), .B(y[8185]), .Z(n47761) );
  XNOR U48288 ( .A(n47760), .B(n47761), .Z(n47762) );
  NAND U48289 ( .A(x[503]), .B(y[8165]), .Z(n47763) );
  XNOR U48290 ( .A(n47762), .B(n47763), .Z(n47810) );
  AND U48291 ( .A(x[485]), .B(y[8183]), .Z(n47753) );
  NAND U48292 ( .A(x[501]), .B(y[8167]), .Z(n47754) );
  XNOR U48293 ( .A(n47753), .B(n47754), .Z(n47755) );
  NAND U48294 ( .A(x[500]), .B(y[8168]), .Z(n47756) );
  XOR U48295 ( .A(n47755), .B(n47756), .Z(n47811) );
  XOR U48296 ( .A(n47810), .B(n47811), .Z(n47813) );
  XOR U48297 ( .A(n47812), .B(n47813), .Z(n47787) );
  NANDN U48298 ( .A(n47618), .B(n47617), .Z(n47622) );
  NANDN U48299 ( .A(n47620), .B(n47619), .Z(n47621) );
  NAND U48300 ( .A(n47622), .B(n47621), .Z(n47703) );
  AND U48301 ( .A(x[480]), .B(y[8188]), .Z(n47710) );
  AND U48302 ( .A(x[508]), .B(y[8160]), .Z(n47709) );
  XOR U48303 ( .A(n47710), .B(n47709), .Z(n47711) );
  XOR U48304 ( .A(n47711), .B(n47712), .Z(n47702) );
  NAND U48305 ( .A(y[8178]), .B(x[490]), .Z(n47624) );
  XNOR U48306 ( .A(n47625), .B(n47624), .Z(n47715) );
  AND U48307 ( .A(x[489]), .B(y[8179]), .Z(n47714) );
  XOR U48308 ( .A(n47715), .B(n47714), .Z(n47701) );
  XOR U48309 ( .A(n47702), .B(n47701), .Z(n47704) );
  XOR U48310 ( .A(n47703), .B(n47704), .Z(n47801) );
  NANDN U48311 ( .A(n47627), .B(n47626), .Z(n47631) );
  NAND U48312 ( .A(n47629), .B(n47628), .Z(n47630) );
  AND U48313 ( .A(n47631), .B(n47630), .Z(n47799) );
  XNOR U48314 ( .A(n47799), .B(n47798), .Z(n47800) );
  XNOR U48315 ( .A(n47801), .B(n47800), .Z(n47786) );
  XOR U48316 ( .A(n47787), .B(n47786), .Z(n47789) );
  XOR U48317 ( .A(n47788), .B(n47789), .Z(n47823) );
  XNOR U48318 ( .A(n47822), .B(n47823), .Z(n47825) );
  NANDN U48319 ( .A(n47637), .B(n47636), .Z(n47641) );
  NANDN U48320 ( .A(n47639), .B(n47638), .Z(n47640) );
  AND U48321 ( .A(n47641), .B(n47640), .Z(n47829) );
  NANDN U48322 ( .A(n47643), .B(n47642), .Z(n47647) );
  NANDN U48323 ( .A(n47645), .B(n47644), .Z(n47646) );
  NAND U48324 ( .A(n47647), .B(n47646), .Z(n47828) );
  XNOR U48325 ( .A(n47830), .B(n47831), .Z(n47684) );
  NANDN U48326 ( .A(n47649), .B(n47648), .Z(n47653) );
  NAND U48327 ( .A(n47651), .B(n47650), .Z(n47652) );
  NAND U48328 ( .A(n47653), .B(n47652), .Z(n47691) );
  NAND U48329 ( .A(n47655), .B(n47654), .Z(n47659) );
  NANDN U48330 ( .A(n47657), .B(n47656), .Z(n47658) );
  AND U48331 ( .A(n47659), .B(n47658), .Z(n47690) );
  NAND U48332 ( .A(n47661), .B(n47660), .Z(n47665) );
  NANDN U48333 ( .A(n47663), .B(n47662), .Z(n47664) );
  AND U48334 ( .A(n47665), .B(n47664), .Z(n47689) );
  XOR U48335 ( .A(n47690), .B(n47689), .Z(n47692) );
  XNOR U48336 ( .A(n47691), .B(n47692), .Z(n47686) );
  XNOR U48337 ( .A(n47679), .B(n47678), .Z(n47682) );
  NAND U48338 ( .A(n47670), .B(n47669), .Z(n47674) );
  NANDN U48339 ( .A(n47672), .B(n47671), .Z(n47673) );
  NAND U48340 ( .A(n47674), .B(n47673), .Z(n47680) );
  XNOR U48341 ( .A(n47681), .B(n47680), .Z(n47675) );
  XNOR U48342 ( .A(n47682), .B(n47675), .Z(N1021) );
  NANDN U48343 ( .A(n47684), .B(n47683), .Z(n47688) );
  NANDN U48344 ( .A(n47686), .B(n47685), .Z(n47687) );
  NAND U48345 ( .A(n47688), .B(n47687), .Z(n47840) );
  NAND U48346 ( .A(n47690), .B(n47689), .Z(n47694) );
  NAND U48347 ( .A(n47692), .B(n47691), .Z(n47693) );
  NAND U48348 ( .A(n47694), .B(n47693), .Z(n47839) );
  NANDN U48349 ( .A(n47696), .B(n47695), .Z(n47700) );
  NANDN U48350 ( .A(n47698), .B(n47697), .Z(n47699) );
  AND U48351 ( .A(n47700), .B(n47699), .Z(n47855) );
  XOR U48352 ( .A(n47983), .B(n47984), .Z(n47985) );
  AND U48353 ( .A(x[490]), .B(y[8180]), .Z(n48000) );
  NAND U48354 ( .A(n47713), .B(n48000), .Z(n47717) );
  NAND U48355 ( .A(n47715), .B(n47714), .Z(n47716) );
  NAND U48356 ( .A(n47717), .B(n47716), .Z(n47967) );
  AND U48357 ( .A(x[502]), .B(y[8167]), .Z(n47934) );
  AND U48358 ( .A(x[481]), .B(y[8188]), .Z(n47932) );
  NAND U48359 ( .A(x[492]), .B(y[8177]), .Z(n48159) );
  XOR U48360 ( .A(n47934), .B(n47933), .Z(n47966) );
  NAND U48361 ( .A(x[495]), .B(y[8174]), .Z(n47935) );
  XNOR U48362 ( .A(n48097), .B(n47935), .Z(n47936) );
  XOR U48363 ( .A(n47966), .B(n47965), .Z(n47968) );
  XNOR U48364 ( .A(n47967), .B(n47968), .Z(n47986) );
  XOR U48365 ( .A(n47985), .B(n47986), .Z(n47961) );
  XOR U48366 ( .A(n47962), .B(n47961), .Z(n47964) );
  NANDN U48367 ( .A(n47719), .B(n47718), .Z(n47723) );
  NANDN U48368 ( .A(n47721), .B(n47720), .Z(n47722) );
  AND U48369 ( .A(n47723), .B(n47722), .Z(n47963) );
  XOR U48370 ( .A(n47964), .B(n47963), .Z(n47958) );
  NAND U48371 ( .A(n47725), .B(n47724), .Z(n47729) );
  NANDN U48372 ( .A(n47727), .B(n47726), .Z(n47728) );
  AND U48373 ( .A(n47729), .B(n47728), .Z(n47956) );
  NANDN U48374 ( .A(n47731), .B(n47730), .Z(n47735) );
  NANDN U48375 ( .A(n47733), .B(n47732), .Z(n47734) );
  NAND U48376 ( .A(n47735), .B(n47734), .Z(n47972) );
  ANDN U48377 ( .B(n47737), .A(n47736), .Z(n47741) );
  NAND U48378 ( .A(n47739), .B(n47738), .Z(n47740) );
  NANDN U48379 ( .A(n47741), .B(n47740), .Z(n47971) );
  XOR U48380 ( .A(n47972), .B(n47971), .Z(n47973) );
  NAND U48381 ( .A(n47743), .B(n47742), .Z(n47747) );
  NAND U48382 ( .A(n47745), .B(n47744), .Z(n47746) );
  NAND U48383 ( .A(n47747), .B(n47746), .Z(n47874) );
  AND U48384 ( .A(x[491]), .B(y[8178]), .Z(n47917) );
  AND U48385 ( .A(x[483]), .B(y[8186]), .Z(n47915) );
  AND U48386 ( .A(x[497]), .B(y[8172]), .Z(n47914) );
  XOR U48387 ( .A(n47915), .B(n47914), .Z(n47916) );
  XOR U48388 ( .A(n47917), .B(n47916), .Z(n47873) );
  AND U48389 ( .A(x[503]), .B(y[8166]), .Z(n47911) );
  AND U48390 ( .A(x[493]), .B(y[8176]), .Z(n47909) );
  AND U48391 ( .A(x[504]), .B(y[8165]), .Z(n48054) );
  XOR U48392 ( .A(n47909), .B(n48054), .Z(n47910) );
  XOR U48393 ( .A(n47911), .B(n47910), .Z(n47872) );
  XOR U48394 ( .A(n47873), .B(n47872), .Z(n47875) );
  XNOR U48395 ( .A(n47874), .B(n47875), .Z(n47974) );
  NANDN U48396 ( .A(n47748), .B(n47902), .Z(n47752) );
  NANDN U48397 ( .A(n47750), .B(n47749), .Z(n47751) );
  NAND U48398 ( .A(n47752), .B(n47751), .Z(n47980) );
  AND U48399 ( .A(x[505]), .B(y[8164]), .Z(n47929) );
  AND U48400 ( .A(x[506]), .B(y[8163]), .Z(n47926) );
  XOR U48401 ( .A(n47927), .B(n47926), .Z(n47928) );
  XOR U48402 ( .A(n47929), .B(n47928), .Z(n47978) );
  AND U48403 ( .A(x[508]), .B(y[8161]), .Z(n47942) );
  XOR U48404 ( .A(o[509]), .B(n47942), .Z(n47995) );
  AND U48405 ( .A(x[480]), .B(y[8189]), .Z(n47993) );
  AND U48406 ( .A(x[509]), .B(y[8160]), .Z(n47992) );
  XOR U48407 ( .A(n47993), .B(n47992), .Z(n47994) );
  XNOR U48408 ( .A(n47995), .B(n47994), .Z(n47977) );
  XOR U48409 ( .A(n47980), .B(n47979), .Z(n47949) );
  NANDN U48410 ( .A(n47754), .B(n47753), .Z(n47758) );
  NANDN U48411 ( .A(n47756), .B(n47755), .Z(n47757) );
  NAND U48412 ( .A(n47758), .B(n47757), .Z(n47922) );
  AND U48413 ( .A(x[482]), .B(y[8187]), .Z(n47885) );
  XOR U48414 ( .A(n47885), .B(n47884), .Z(n47886) );
  XOR U48415 ( .A(n47887), .B(n47886), .Z(n47921) );
  AND U48416 ( .A(n47759), .B(o[508]), .Z(n47893) );
  AND U48417 ( .A(x[496]), .B(y[8173]), .Z(n47891) );
  AND U48418 ( .A(x[507]), .B(y[8162]), .Z(n47890) );
  XOR U48419 ( .A(n47891), .B(n47890), .Z(n47892) );
  XOR U48420 ( .A(n47893), .B(n47892), .Z(n47920) );
  XOR U48421 ( .A(n47921), .B(n47920), .Z(n47923) );
  XOR U48422 ( .A(n47922), .B(n47923), .Z(n47950) );
  NANDN U48423 ( .A(n47761), .B(n47760), .Z(n47765) );
  NANDN U48424 ( .A(n47763), .B(n47762), .Z(n47764) );
  NAND U48425 ( .A(n47765), .B(n47764), .Z(n47897) );
  NANDN U48426 ( .A(n47767), .B(n47766), .Z(n47771) );
  NAND U48427 ( .A(n47769), .B(n47768), .Z(n47770) );
  NAND U48428 ( .A(n47771), .B(n47770), .Z(n47896) );
  XOR U48429 ( .A(n47897), .B(n47896), .Z(n47899) );
  AND U48430 ( .A(x[488]), .B(y[8181]), .Z(n47904) );
  AND U48431 ( .A(x[486]), .B(y[8183]), .Z(n47773) );
  AND U48432 ( .A(y[8182]), .B(x[487]), .Z(n47772) );
  XOR U48433 ( .A(n47773), .B(n47772), .Z(n47903) );
  XOR U48434 ( .A(n47904), .B(n47903), .Z(n47987) );
  AND U48435 ( .A(x[489]), .B(y[8180]), .Z(n48104) );
  XOR U48436 ( .A(n47987), .B(n48104), .Z(n47989) );
  AND U48437 ( .A(x[485]), .B(y[8184]), .Z(n47881) );
  AND U48438 ( .A(x[484]), .B(y[8185]), .Z(n47879) );
  AND U48439 ( .A(x[490]), .B(y[8179]), .Z(n47878) );
  XOR U48440 ( .A(n47879), .B(n47878), .Z(n47880) );
  XOR U48441 ( .A(n47881), .B(n47880), .Z(n47988) );
  XOR U48442 ( .A(n47989), .B(n47988), .Z(n47898) );
  XOR U48443 ( .A(n47899), .B(n47898), .Z(n47867) );
  NANDN U48444 ( .A(n47775), .B(n47774), .Z(n47779) );
  OR U48445 ( .A(n47777), .B(n47776), .Z(n47778) );
  NAND U48446 ( .A(n47779), .B(n47778), .Z(n47866) );
  XNOR U48447 ( .A(n47867), .B(n47866), .Z(n47868) );
  XNOR U48448 ( .A(n47869), .B(n47868), .Z(n47955) );
  XNOR U48449 ( .A(n47855), .B(n47854), .Z(n47857) );
  NANDN U48450 ( .A(n47781), .B(n47780), .Z(n47785) );
  NANDN U48451 ( .A(n47783), .B(n47782), .Z(n47784) );
  AND U48452 ( .A(n47785), .B(n47784), .Z(n47851) );
  NANDN U48453 ( .A(n47787), .B(n47786), .Z(n47791) );
  OR U48454 ( .A(n47789), .B(n47788), .Z(n47790) );
  AND U48455 ( .A(n47791), .B(n47790), .Z(n47850) );
  XNOR U48456 ( .A(n47851), .B(n47850), .Z(n47853) );
  NANDN U48457 ( .A(n47793), .B(n47792), .Z(n47797) );
  NANDN U48458 ( .A(n47795), .B(n47794), .Z(n47796) );
  NAND U48459 ( .A(n47797), .B(n47796), .Z(n47862) );
  NANDN U48460 ( .A(n47799), .B(n47798), .Z(n47803) );
  NAND U48461 ( .A(n47801), .B(n47800), .Z(n47802) );
  AND U48462 ( .A(n47803), .B(n47802), .Z(n47946) );
  NANDN U48463 ( .A(n47805), .B(n47804), .Z(n47809) );
  OR U48464 ( .A(n47807), .B(n47806), .Z(n47808) );
  AND U48465 ( .A(n47809), .B(n47808), .Z(n47944) );
  NANDN U48466 ( .A(n47811), .B(n47810), .Z(n47815) );
  OR U48467 ( .A(n47813), .B(n47812), .Z(n47814) );
  NAND U48468 ( .A(n47815), .B(n47814), .Z(n47943) );
  XNOR U48469 ( .A(n47944), .B(n47943), .Z(n47945) );
  XNOR U48470 ( .A(n47946), .B(n47945), .Z(n47861) );
  NANDN U48471 ( .A(n47817), .B(n47816), .Z(n47821) );
  NANDN U48472 ( .A(n47819), .B(n47818), .Z(n47820) );
  NAND U48473 ( .A(n47821), .B(n47820), .Z(n47860) );
  XOR U48474 ( .A(n47861), .B(n47860), .Z(n47863) );
  XOR U48475 ( .A(n47862), .B(n47863), .Z(n47852) );
  XOR U48476 ( .A(n47853), .B(n47852), .Z(n47856) );
  XOR U48477 ( .A(n47857), .B(n47856), .Z(n47847) );
  NAND U48478 ( .A(n47823), .B(n47822), .Z(n47827) );
  NANDN U48479 ( .A(n47825), .B(n47824), .Z(n47826) );
  AND U48480 ( .A(n47827), .B(n47826), .Z(n47845) );
  NANDN U48481 ( .A(n47829), .B(n47828), .Z(n47833) );
  NAND U48482 ( .A(n47831), .B(n47830), .Z(n47832) );
  AND U48483 ( .A(n47833), .B(n47832), .Z(n47844) );
  XOR U48484 ( .A(n47847), .B(n47846), .Z(n47838) );
  XOR U48485 ( .A(n47839), .B(n47838), .Z(n47841) );
  XOR U48486 ( .A(n47840), .B(n47841), .Z(n47837) );
  XOR U48487 ( .A(n47835), .B(n47837), .Z(n47834) );
  XOR U48488 ( .A(n47836), .B(n47834), .Z(N1022) );
  NAND U48489 ( .A(n47839), .B(n47838), .Z(n47843) );
  NAND U48490 ( .A(n47841), .B(n47840), .Z(n47842) );
  AND U48491 ( .A(n47843), .B(n47842), .Z(n48258) );
  XNOR U48492 ( .A(n48259), .B(n48258), .Z(n48257) );
  NANDN U48493 ( .A(n47845), .B(n47844), .Z(n47849) );
  NANDN U48494 ( .A(n47847), .B(n47846), .Z(n47848) );
  AND U48495 ( .A(n47849), .B(n47848), .Z(n48275) );
  NANDN U48496 ( .A(n47855), .B(n47854), .Z(n47859) );
  NAND U48497 ( .A(n47857), .B(n47856), .Z(n47858) );
  AND U48498 ( .A(n47859), .B(n47858), .Z(n48246) );
  XOR U48499 ( .A(n48247), .B(n48246), .Z(n48245) );
  NAND U48500 ( .A(n47861), .B(n47860), .Z(n47865) );
  NAND U48501 ( .A(n47863), .B(n47862), .Z(n47864) );
  AND U48502 ( .A(n47865), .B(n47864), .Z(n48244) );
  XOR U48503 ( .A(n48245), .B(n48244), .Z(n48277) );
  NANDN U48504 ( .A(n47867), .B(n47866), .Z(n47871) );
  NAND U48505 ( .A(n47869), .B(n47868), .Z(n47870) );
  AND U48506 ( .A(n47871), .B(n47870), .Z(n48002) );
  NAND U48507 ( .A(n47873), .B(n47872), .Z(n47877) );
  NAND U48508 ( .A(n47875), .B(n47874), .Z(n47876) );
  AND U48509 ( .A(n47877), .B(n47876), .Z(n48010) );
  NAND U48510 ( .A(n47879), .B(n47878), .Z(n47883) );
  NAND U48511 ( .A(n47881), .B(n47880), .Z(n47882) );
  NAND U48512 ( .A(n47883), .B(n47882), .Z(n48023) );
  AND U48513 ( .A(x[486]), .B(y[8184]), .Z(n48153) );
  AND U48514 ( .A(x[485]), .B(y[8185]), .Z(n48155) );
  AND U48515 ( .A(x[499]), .B(y[8171]), .Z(n48154) );
  XOR U48516 ( .A(n48155), .B(n48154), .Z(n48152) );
  XNOR U48517 ( .A(n48153), .B(n48152), .Z(n48029) );
  AND U48518 ( .A(x[484]), .B(y[8186]), .Z(n48099) );
  AND U48519 ( .A(x[483]), .B(y[8187]), .Z(n48101) );
  AND U48520 ( .A(x[498]), .B(y[8172]), .Z(n48100) );
  XOR U48521 ( .A(n48101), .B(n48100), .Z(n48098) );
  XOR U48522 ( .A(n48099), .B(n48098), .Z(n48026) );
  NAND U48523 ( .A(n47885), .B(n47884), .Z(n47889) );
  NAND U48524 ( .A(n47887), .B(n47886), .Z(n47888) );
  AND U48525 ( .A(n47889), .B(n47888), .Z(n48027) );
  XOR U48526 ( .A(n48029), .B(n48028), .Z(n48022) );
  XOR U48527 ( .A(n48023), .B(n48022), .Z(n48021) );
  NAND U48528 ( .A(n47891), .B(n47890), .Z(n47895) );
  NAND U48529 ( .A(n47893), .B(n47892), .Z(n47894) );
  NAND U48530 ( .A(n47895), .B(n47894), .Z(n48020) );
  XOR U48531 ( .A(n48021), .B(n48020), .Z(n48011) );
  NAND U48532 ( .A(n47897), .B(n47896), .Z(n47901) );
  NAND U48533 ( .A(n47899), .B(n47898), .Z(n47900) );
  AND U48534 ( .A(n47901), .B(n47900), .Z(n48008) );
  XOR U48535 ( .A(n48009), .B(n48008), .Z(n48005) );
  AND U48536 ( .A(x[487]), .B(y[8183]), .Z(n48096) );
  NAND U48537 ( .A(n47902), .B(n48096), .Z(n47906) );
  NAND U48538 ( .A(n47904), .B(n47903), .Z(n47905) );
  AND U48539 ( .A(n47906), .B(n47905), .Z(n48035) );
  AND U48540 ( .A(y[8169]), .B(x[501]), .Z(n47908) );
  AND U48541 ( .A(y[8168]), .B(x[502]), .Z(n47907) );
  XOR U48542 ( .A(n47908), .B(n47907), .Z(n48095) );
  XOR U48543 ( .A(n48096), .B(n48095), .Z(n48033) );
  AND U48544 ( .A(x[497]), .B(y[8173]), .Z(n48064) );
  AND U48545 ( .A(x[482]), .B(y[8188]), .Z(n48066) );
  AND U48546 ( .A(x[506]), .B(y[8164]), .Z(n48065) );
  XOR U48547 ( .A(n48066), .B(n48065), .Z(n48063) );
  XNOR U48548 ( .A(n48064), .B(n48063), .Z(n48032) );
  XNOR U48549 ( .A(n48035), .B(n48034), .Z(n48015) );
  NAND U48550 ( .A(n47909), .B(n48054), .Z(n47913) );
  NAND U48551 ( .A(n47911), .B(n47910), .Z(n47912) );
  NAND U48552 ( .A(n47913), .B(n47912), .Z(n48017) );
  NAND U48553 ( .A(n47915), .B(n47914), .Z(n47919) );
  NAND U48554 ( .A(n47917), .B(n47916), .Z(n47918) );
  AND U48555 ( .A(n47919), .B(n47918), .Z(n48041) );
  AND U48556 ( .A(x[480]), .B(y[8190]), .Z(n48090) );
  AND U48557 ( .A(x[509]), .B(y[8161]), .Z(n48105) );
  XOR U48558 ( .A(o[510]), .B(n48105), .Z(n48092) );
  AND U48559 ( .A(x[510]), .B(y[8160]), .Z(n48091) );
  XOR U48560 ( .A(n48092), .B(n48091), .Z(n48089) );
  XOR U48561 ( .A(n48090), .B(n48089), .Z(n48039) );
  AND U48562 ( .A(x[500]), .B(y[8170]), .Z(n48172) );
  XOR U48563 ( .A(n48173), .B(n48172), .Z(n48171) );
  AND U48564 ( .A(x[488]), .B(y[8182]), .Z(n48170) );
  XNOR U48565 ( .A(n48171), .B(n48170), .Z(n48038) );
  XNOR U48566 ( .A(n48041), .B(n48040), .Z(n48016) );
  XOR U48567 ( .A(n48017), .B(n48016), .Z(n48014) );
  NAND U48568 ( .A(n47921), .B(n47920), .Z(n47925) );
  NAND U48569 ( .A(n47923), .B(n47922), .Z(n47924) );
  NAND U48570 ( .A(n47925), .B(n47924), .Z(n48230) );
  XOR U48571 ( .A(n48231), .B(n48230), .Z(n48229) );
  AND U48572 ( .A(n47927), .B(n47926), .Z(n47931) );
  NAND U48573 ( .A(n47929), .B(n47928), .Z(n47930) );
  NANDN U48574 ( .A(n47931), .B(n47930), .Z(n48046) );
  NANDN U48575 ( .A(n47935), .B(n48097), .Z(n47939) );
  NANDN U48576 ( .A(n47937), .B(n47936), .Z(n47938) );
  AND U48577 ( .A(n47939), .B(n47938), .Z(n48189) );
  AND U48578 ( .A(x[503]), .B(y[8167]), .Z(n48053) );
  AND U48579 ( .A(y[8166]), .B(x[504]), .Z(n47941) );
  AND U48580 ( .A(y[8165]), .B(x[505]), .Z(n47940) );
  XOR U48581 ( .A(n47941), .B(n47940), .Z(n48052) );
  XOR U48582 ( .A(n48053), .B(n48052), .Z(n48191) );
  AND U48583 ( .A(n47942), .B(o[509]), .Z(n48058) );
  AND U48584 ( .A(x[508]), .B(y[8162]), .Z(n48060) );
  AND U48585 ( .A(x[496]), .B(y[8174]), .Z(n48059) );
  XOR U48586 ( .A(n48060), .B(n48059), .Z(n48057) );
  XNOR U48587 ( .A(n48058), .B(n48057), .Z(n48190) );
  XNOR U48588 ( .A(n48189), .B(n48188), .Z(n48048) );
  XOR U48589 ( .A(n48049), .B(n48048), .Z(n48047) );
  XOR U48590 ( .A(n48046), .B(n48047), .Z(n48228) );
  XOR U48591 ( .A(n48229), .B(n48228), .Z(n48004) );
  XOR U48592 ( .A(n48002), .B(n48003), .Z(n48240) );
  NANDN U48593 ( .A(n47944), .B(n47943), .Z(n47948) );
  NANDN U48594 ( .A(n47946), .B(n47945), .Z(n47947) );
  AND U48595 ( .A(n47948), .B(n47947), .Z(n48243) );
  NANDN U48596 ( .A(n47950), .B(n47949), .Z(n47954) );
  NANDN U48597 ( .A(n47952), .B(n47951), .Z(n47953) );
  NAND U48598 ( .A(n47954), .B(n47953), .Z(n48242) );
  XOR U48599 ( .A(n48243), .B(n48242), .Z(n48241) );
  XOR U48600 ( .A(n48240), .B(n48241), .Z(n48263) );
  NANDN U48601 ( .A(n47956), .B(n47955), .Z(n47960) );
  NANDN U48602 ( .A(n47958), .B(n47957), .Z(n47959) );
  NAND U48603 ( .A(n47960), .B(n47959), .Z(n48264) );
  NAND U48604 ( .A(n47966), .B(n47965), .Z(n47970) );
  NAND U48605 ( .A(n47968), .B(n47967), .Z(n47969) );
  AND U48606 ( .A(n47970), .B(n47969), .Z(n48213) );
  NAND U48607 ( .A(n47972), .B(n47971), .Z(n47976) );
  NANDN U48608 ( .A(n47974), .B(n47973), .Z(n47975) );
  AND U48609 ( .A(n47976), .B(n47975), .Z(n48212) );
  XOR U48610 ( .A(n48213), .B(n48212), .Z(n48211) );
  NANDN U48611 ( .A(n47978), .B(n47977), .Z(n47982) );
  OR U48612 ( .A(n47980), .B(n47979), .Z(n47981) );
  NAND U48613 ( .A(n47982), .B(n47981), .Z(n48210) );
  XOR U48614 ( .A(n48211), .B(n48210), .Z(n48225) );
  NAND U48615 ( .A(n47987), .B(n48104), .Z(n47991) );
  NAND U48616 ( .A(n47989), .B(n47988), .Z(n47990) );
  AND U48617 ( .A(n47991), .B(n47990), .Z(n48207) );
  NAND U48618 ( .A(n47993), .B(n47992), .Z(n47997) );
  NAND U48619 ( .A(n47995), .B(n47994), .Z(n47996) );
  NAND U48620 ( .A(n47997), .B(n47996), .Z(n48182) );
  AND U48621 ( .A(y[8178]), .B(x[492]), .Z(n47998) );
  XOR U48622 ( .A(n47999), .B(n47998), .Z(n48160) );
  XOR U48623 ( .A(n48161), .B(n48160), .Z(n48103) );
  AND U48624 ( .A(y[8181]), .B(x[489]), .Z(n48001) );
  XOR U48625 ( .A(n48001), .B(n48000), .Z(n48102) );
  XOR U48626 ( .A(n48103), .B(n48102), .Z(n48185) );
  AND U48627 ( .A(x[507]), .B(y[8163]), .Z(n48169) );
  AND U48628 ( .A(x[481]), .B(y[8189]), .Z(n48168) );
  XOR U48629 ( .A(n48169), .B(n48168), .Z(n48166) );
  XOR U48630 ( .A(n48167), .B(n48166), .Z(n48184) );
  XNOR U48631 ( .A(n48185), .B(n48184), .Z(n48183) );
  XOR U48632 ( .A(n48182), .B(n48183), .Z(n48206) );
  XOR U48633 ( .A(n48207), .B(n48206), .Z(n48205) );
  XNOR U48634 ( .A(n48204), .B(n48205), .Z(n48224) );
  XNOR U48635 ( .A(n48222), .B(n48223), .Z(n48265) );
  XOR U48636 ( .A(n48264), .B(n48265), .Z(n48262) );
  XNOR U48637 ( .A(n48275), .B(n48274), .Z(n48256) );
  XNOR U48638 ( .A(n48257), .B(n48256), .Z(N1023) );
  NANDN U48639 ( .A(n48003), .B(n48002), .Z(n48007) );
  NANDN U48640 ( .A(n48005), .B(n48004), .Z(n48006) );
  AND U48641 ( .A(n48007), .B(n48006), .Z(n48273) );
  NAND U48642 ( .A(n48009), .B(n48008), .Z(n48013) );
  NANDN U48643 ( .A(n48011), .B(n48010), .Z(n48012) );
  AND U48644 ( .A(n48013), .B(n48012), .Z(n48255) );
  NANDN U48645 ( .A(n48015), .B(n48014), .Z(n48019) );
  NAND U48646 ( .A(n48017), .B(n48016), .Z(n48018) );
  AND U48647 ( .A(n48019), .B(n48018), .Z(n48239) );
  NAND U48648 ( .A(n48021), .B(n48020), .Z(n48025) );
  NAND U48649 ( .A(n48023), .B(n48022), .Z(n48024) );
  AND U48650 ( .A(n48025), .B(n48024), .Z(n48221) );
  ANDN U48651 ( .B(n48027), .A(n48026), .Z(n48031) );
  ANDN U48652 ( .B(n48029), .A(n48028), .Z(n48030) );
  NOR U48653 ( .A(n48031), .B(n48030), .Z(n48203) );
  NANDN U48654 ( .A(n48033), .B(n48032), .Z(n48037) );
  ANDN U48655 ( .B(n48035), .A(n48034), .Z(n48036) );
  ANDN U48656 ( .B(n48037), .A(n48036), .Z(n48045) );
  NANDN U48657 ( .A(n48039), .B(n48038), .Z(n48043) );
  AND U48658 ( .A(n48041), .B(n48040), .Z(n48042) );
  ANDN U48659 ( .B(n48043), .A(n48042), .Z(n48044) );
  XNOR U48660 ( .A(n48045), .B(n48044), .Z(n48201) );
  NAND U48661 ( .A(n48047), .B(n48046), .Z(n48051) );
  NAND U48662 ( .A(n48049), .B(n48048), .Z(n48050) );
  AND U48663 ( .A(n48051), .B(n48050), .Z(n48199) );
  NAND U48664 ( .A(n48053), .B(n48052), .Z(n48056) );
  AND U48665 ( .A(x[505]), .B(y[8166]), .Z(n48106) );
  NAND U48666 ( .A(n48054), .B(n48106), .Z(n48055) );
  AND U48667 ( .A(n48056), .B(n48055), .Z(n48088) );
  NAND U48668 ( .A(n48058), .B(n48057), .Z(n48062) );
  NAND U48669 ( .A(n48060), .B(n48059), .Z(n48061) );
  AND U48670 ( .A(n48062), .B(n48061), .Z(n48070) );
  NAND U48671 ( .A(n48064), .B(n48063), .Z(n48068) );
  NAND U48672 ( .A(n48066), .B(n48065), .Z(n48067) );
  NAND U48673 ( .A(n48068), .B(n48067), .Z(n48069) );
  XNOR U48674 ( .A(n48070), .B(n48069), .Z(n48086) );
  AND U48675 ( .A(y[8190]), .B(x[481]), .Z(n48072) );
  NAND U48676 ( .A(y[8163]), .B(x[508]), .Z(n48071) );
  XNOR U48677 ( .A(n48072), .B(n48071), .Z(n48076) );
  AND U48678 ( .A(y[8179]), .B(x[492]), .Z(n48074) );
  NAND U48679 ( .A(y[8191]), .B(x[480]), .Z(n48073) );
  XNOR U48680 ( .A(n48074), .B(n48073), .Z(n48075) );
  XOR U48681 ( .A(n48076), .B(n48075), .Z(n48084) );
  AND U48682 ( .A(y[8189]), .B(x[482]), .Z(n48078) );
  NAND U48683 ( .A(y[8183]), .B(x[488]), .Z(n48077) );
  XNOR U48684 ( .A(n48078), .B(n48077), .Z(n48082) );
  AND U48685 ( .A(y[8160]), .B(x[511]), .Z(n48080) );
  NAND U48686 ( .A(y[8172]), .B(x[499]), .Z(n48079) );
  XNOR U48687 ( .A(n48080), .B(n48079), .Z(n48081) );
  XNOR U48688 ( .A(n48082), .B(n48081), .Z(n48083) );
  XNOR U48689 ( .A(n48084), .B(n48083), .Z(n48085) );
  XNOR U48690 ( .A(n48086), .B(n48085), .Z(n48087) );
  XNOR U48691 ( .A(n48088), .B(n48087), .Z(n48151) );
  NAND U48692 ( .A(n48090), .B(n48089), .Z(n48094) );
  NAND U48693 ( .A(n48092), .B(n48091), .Z(n48093) );
  AND U48694 ( .A(n48094), .B(n48093), .Z(n48149) );
  AND U48695 ( .A(x[502]), .B(y[8169]), .Z(n48107) );
  AND U48696 ( .A(x[490]), .B(y[8181]), .Z(n48127) );
  AND U48697 ( .A(n48105), .B(o[510]), .Z(n48112) );
  XOR U48698 ( .A(n48106), .B(o[511]), .Z(n48110) );
  XNOR U48699 ( .A(n48108), .B(n48107), .Z(n48109) );
  XNOR U48700 ( .A(n48110), .B(n48109), .Z(n48111) );
  AND U48701 ( .A(y[8182]), .B(x[489]), .Z(n48118) );
  AND U48702 ( .A(y[8180]), .B(x[491]), .Z(n48114) );
  NAND U48703 ( .A(y[8165]), .B(x[506]), .Z(n48113) );
  XNOR U48704 ( .A(n48114), .B(n48113), .Z(n48115) );
  XNOR U48705 ( .A(n48116), .B(n48115), .Z(n48117) );
  XNOR U48706 ( .A(n48118), .B(n48117), .Z(n48141) );
  AND U48707 ( .A(y[8186]), .B(x[485]), .Z(n48120) );
  NAND U48708 ( .A(y[8185]), .B(x[486]), .Z(n48119) );
  XNOR U48709 ( .A(n48120), .B(n48119), .Z(n48131) );
  AND U48710 ( .A(y[8188]), .B(x[483]), .Z(n48122) );
  NAND U48711 ( .A(y[8173]), .B(x[498]), .Z(n48121) );
  XNOR U48712 ( .A(n48122), .B(n48121), .Z(n48126) );
  AND U48713 ( .A(y[8162]), .B(x[509]), .Z(n48124) );
  NAND U48714 ( .A(y[8184]), .B(x[487]), .Z(n48123) );
  XNOR U48715 ( .A(n48124), .B(n48123), .Z(n48125) );
  XOR U48716 ( .A(n48126), .B(n48125), .Z(n48129) );
  XNOR U48717 ( .A(n48158), .B(n48127), .Z(n48128) );
  XNOR U48718 ( .A(n48129), .B(n48128), .Z(n48130) );
  XOR U48719 ( .A(n48131), .B(n48130), .Z(n48139) );
  AND U48720 ( .A(y[8164]), .B(x[507]), .Z(n48133) );
  NAND U48721 ( .A(y[8170]), .B(x[501]), .Z(n48132) );
  XNOR U48722 ( .A(n48133), .B(n48132), .Z(n48137) );
  AND U48723 ( .A(y[8168]), .B(x[503]), .Z(n48135) );
  NAND U48724 ( .A(y[8174]), .B(x[497]), .Z(n48134) );
  XNOR U48725 ( .A(n48135), .B(n48134), .Z(n48136) );
  XNOR U48726 ( .A(n48137), .B(n48136), .Z(n48138) );
  XNOR U48727 ( .A(n48139), .B(n48138), .Z(n48140) );
  AND U48728 ( .A(y[8161]), .B(x[510]), .Z(n48143) );
  NAND U48729 ( .A(y[8175]), .B(x[496]), .Z(n48142) );
  XNOR U48730 ( .A(n48143), .B(n48142), .Z(n48147) );
  AND U48731 ( .A(y[8177]), .B(x[494]), .Z(n48145) );
  NAND U48732 ( .A(y[8171]), .B(x[500]), .Z(n48144) );
  XNOR U48733 ( .A(n48145), .B(n48144), .Z(n48146) );
  XNOR U48734 ( .A(n48149), .B(n48148), .Z(n48150) );
  XOR U48735 ( .A(n48151), .B(n48150), .Z(n48181) );
  NAND U48736 ( .A(n48153), .B(n48152), .Z(n48157) );
  NAND U48737 ( .A(n48155), .B(n48154), .Z(n48156) );
  AND U48738 ( .A(n48157), .B(n48156), .Z(n48165) );
  NANDN U48739 ( .A(n48159), .B(n48158), .Z(n48163) );
  NAND U48740 ( .A(n48161), .B(n48160), .Z(n48162) );
  AND U48741 ( .A(n48163), .B(n48162), .Z(n48164) );
  XNOR U48742 ( .A(n48165), .B(n48164), .Z(n48179) );
  NAND U48743 ( .A(n48171), .B(n48170), .Z(n48175) );
  NAND U48744 ( .A(n48173), .B(n48172), .Z(n48174) );
  NAND U48745 ( .A(n48175), .B(n48174), .Z(n48176) );
  XNOR U48746 ( .A(n48177), .B(n48176), .Z(n48178) );
  XOR U48747 ( .A(n48179), .B(n48178), .Z(n48180) );
  XNOR U48748 ( .A(n48181), .B(n48180), .Z(n48197) );
  NANDN U48749 ( .A(n48183), .B(n48182), .Z(n48187) );
  NAND U48750 ( .A(n48185), .B(n48184), .Z(n48186) );
  AND U48751 ( .A(n48187), .B(n48186), .Z(n48195) );
  NAND U48752 ( .A(n48189), .B(n48188), .Z(n48193) );
  NANDN U48753 ( .A(n48191), .B(n48190), .Z(n48192) );
  NAND U48754 ( .A(n48193), .B(n48192), .Z(n48194) );
  XNOR U48755 ( .A(n48195), .B(n48194), .Z(n48196) );
  XNOR U48756 ( .A(n48197), .B(n48196), .Z(n48198) );
  XNOR U48757 ( .A(n48199), .B(n48198), .Z(n48200) );
  XOR U48758 ( .A(n48201), .B(n48200), .Z(n48202) );
  XNOR U48759 ( .A(n48203), .B(n48202), .Z(n48219) );
  NAND U48760 ( .A(n48205), .B(n48204), .Z(n48209) );
  NAND U48761 ( .A(n48207), .B(n48206), .Z(n48208) );
  AND U48762 ( .A(n48209), .B(n48208), .Z(n48217) );
  NAND U48763 ( .A(n48213), .B(n48212), .Z(n48214) );
  NAND U48764 ( .A(n48215), .B(n48214), .Z(n48216) );
  XNOR U48765 ( .A(n48217), .B(n48216), .Z(n48218) );
  XNOR U48766 ( .A(n48219), .B(n48218), .Z(n48220) );
  XNOR U48767 ( .A(n48221), .B(n48220), .Z(n48237) );
  NANDN U48768 ( .A(n48223), .B(n48222), .Z(n48227) );
  NANDN U48769 ( .A(n48225), .B(n48224), .Z(n48226) );
  AND U48770 ( .A(n48227), .B(n48226), .Z(n48235) );
  NAND U48771 ( .A(n48229), .B(n48228), .Z(n48233) );
  NAND U48772 ( .A(n48231), .B(n48230), .Z(n48232) );
  NAND U48773 ( .A(n48233), .B(n48232), .Z(n48234) );
  XNOR U48774 ( .A(n48235), .B(n48234), .Z(n48236) );
  XNOR U48775 ( .A(n48237), .B(n48236), .Z(n48238) );
  XNOR U48776 ( .A(n48239), .B(n48238), .Z(n48253) );
  NAND U48777 ( .A(n48245), .B(n48244), .Z(n48249) );
  NAND U48778 ( .A(n48247), .B(n48246), .Z(n48248) );
  NAND U48779 ( .A(n48249), .B(n48248), .Z(n48250) );
  XNOR U48780 ( .A(n48251), .B(n48250), .Z(n48252) );
  XNOR U48781 ( .A(n48253), .B(n48252), .Z(n48254) );
  XNOR U48782 ( .A(n48255), .B(n48254), .Z(n48271) );
  NAND U48783 ( .A(n48257), .B(n48256), .Z(n48261) );
  NANDN U48784 ( .A(n48259), .B(n48258), .Z(n48260) );
  AND U48785 ( .A(n48261), .B(n48260), .Z(n48269) );
  NANDN U48786 ( .A(n48263), .B(n48262), .Z(n48267) );
  NAND U48787 ( .A(n48265), .B(n48264), .Z(n48266) );
  NAND U48788 ( .A(n48267), .B(n48266), .Z(n48268) );
  XNOR U48789 ( .A(n48269), .B(n48268), .Z(n48270) );
  XNOR U48790 ( .A(n48271), .B(n48270), .Z(n48272) );
  XNOR U48791 ( .A(n48273), .B(n48272), .Z(n48281) );
  NAND U48792 ( .A(n48275), .B(n48274), .Z(n48279) );
  NANDN U48793 ( .A(n48277), .B(n48276), .Z(n48278) );
  NAND U48794 ( .A(n48279), .B(n48278), .Z(n48280) );
  XNOR U48795 ( .A(n48281), .B(n48280), .Z(N1024) );
endmodule

