
module mult_N64_CC8 ( clk, rst, a, b, c );
  input [63:0] a;
  input [7:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153;
  wire   [63:8] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[112]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[113]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[114]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[115]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[116]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[117]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[118]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[119]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U11 ( .A(n2068), .B(n2089), .Z(n2077) );
  XNOR U12 ( .A(n1998), .B(n2014), .Z(n2002) );
  XNOR U13 ( .A(n1975), .B(n1974), .Z(n1949) );
  XOR U14 ( .A(n887), .B(n914), .Z(n892) );
  XOR U15 ( .A(n963), .B(n990), .Z(n968) );
  XOR U16 ( .A(n1039), .B(n1066), .Z(n1044) );
  XOR U17 ( .A(n1115), .B(n1142), .Z(n1120) );
  XOR U18 ( .A(n1191), .B(n1218), .Z(n1196) );
  XOR U19 ( .A(n1267), .B(n1294), .Z(n1272) );
  XOR U20 ( .A(n1343), .B(n1370), .Z(n1348) );
  XOR U21 ( .A(n1419), .B(n1446), .Z(n1424) );
  XOR U22 ( .A(n1495), .B(n1522), .Z(n1500) );
  XOR U23 ( .A(n1571), .B(n1598), .Z(n1576) );
  XOR U24 ( .A(n1647), .B(n1674), .Z(n1652) );
  XOR U25 ( .A(n1723), .B(n1750), .Z(n1728) );
  XOR U26 ( .A(n1799), .B(n1826), .Z(n1804) );
  XOR U27 ( .A(n1875), .B(n1912), .Z(n1880) );
  XOR U28 ( .A(n1971), .B(n1976), .Z(n1948) );
  XNOR U29 ( .A(n2104), .B(n2112), .Z(n2100) );
  XNOR U30 ( .A(n2040), .B(n2048), .Z(n2036) );
  AND U31 ( .A(n117), .B(n116), .Z(n84) );
  XOR U32 ( .A(n925), .B(n952), .Z(n930) );
  XOR U33 ( .A(n1001), .B(n1028), .Z(n1006) );
  XOR U34 ( .A(n1077), .B(n1104), .Z(n1082) );
  XOR U35 ( .A(n1153), .B(n1180), .Z(n1158) );
  XOR U36 ( .A(n1229), .B(n1256), .Z(n1234) );
  XOR U37 ( .A(n1305), .B(n1332), .Z(n1310) );
  XOR U38 ( .A(n1381), .B(n1408), .Z(n1386) );
  XOR U39 ( .A(n1457), .B(n1484), .Z(n1462) );
  XOR U40 ( .A(n1533), .B(n1560), .Z(n1538) );
  XOR U41 ( .A(n1609), .B(n1636), .Z(n1614) );
  XOR U42 ( .A(n1685), .B(n1712), .Z(n1690) );
  XOR U43 ( .A(n1761), .B(n1788), .Z(n1766) );
  XOR U44 ( .A(n1837), .B(n1864), .Z(n1842) );
  XOR U45 ( .A(n1929), .B(n1943), .Z(n1934) );
  AND U46 ( .A(a[1]), .B(n2138), .Z(n2149) );
  XNOR U47 ( .A(n2077), .B(n2085), .Z(n2073) );
  XNOR U48 ( .A(n2002), .B(n2010), .Z(n1980) );
  AND U49 ( .A(n149), .B(n148), .Z(n116) );
  XOR U50 ( .A(n1992), .B(n2015), .Z(n1997) );
  XOR U51 ( .A(n1923), .B(n1952), .Z(n1928) );
  XOR U52 ( .A(n73), .B(n92), .Z(n83) );
  XOR U53 ( .A(n137), .B(n157), .Z(n147) );
  XOR U54 ( .A(n202), .B(n222), .Z(n212) );
  XOR U55 ( .A(n273), .B(n294), .Z(n283) );
  XOR U56 ( .A(n341), .B(n362), .Z(n351) );
  XOR U57 ( .A(n409), .B(n430), .Z(n419) );
  XOR U58 ( .A(n477), .B(n498), .Z(n487) );
  XOR U59 ( .A(n545), .B(n566), .Z(n555) );
  XOR U60 ( .A(n613), .B(n634), .Z(n623) );
  XOR U61 ( .A(n681), .B(n702), .Z(n691) );
  XOR U62 ( .A(n749), .B(n770), .Z(n759) );
  XOR U63 ( .A(n817), .B(n838), .Z(n827) );
  XOR U64 ( .A(n893), .B(n913), .Z(n902) );
  XOR U65 ( .A(n969), .B(n989), .Z(n978) );
  XOR U66 ( .A(n1045), .B(n1065), .Z(n1054) );
  XOR U67 ( .A(n1121), .B(n1141), .Z(n1130) );
  XOR U68 ( .A(n1197), .B(n1217), .Z(n1206) );
  XOR U69 ( .A(n1273), .B(n1293), .Z(n1282) );
  XOR U70 ( .A(n1349), .B(n1369), .Z(n1358) );
  XOR U71 ( .A(n1425), .B(n1445), .Z(n1434) );
  XOR U72 ( .A(n1501), .B(n1521), .Z(n1510) );
  XOR U73 ( .A(n1577), .B(n1597), .Z(n1586) );
  XOR U74 ( .A(n1653), .B(n1673), .Z(n1662) );
  XOR U75 ( .A(n1729), .B(n1749), .Z(n1738) );
  XOR U76 ( .A(n1805), .B(n1825), .Z(n1814) );
  XOR U77 ( .A(n1881), .B(n1911), .Z(n1890) );
  XNOR U78 ( .A(n1949), .B(n1947), .Z(n1937) );
  XNOR U79 ( .A(n2140), .B(n2141), .Z(n2135) );
  XNOR U80 ( .A(n2100), .B(n2099), .Z(n2088) );
  XNOR U81 ( .A(n2036), .B(n2035), .Z(n2013) );
  AND U82 ( .A(n182), .B(n181), .Z(n148) );
  XOR U83 ( .A(n2026), .B(n2054), .Z(n2031) );
  XOR U84 ( .A(n1965), .B(n1981), .Z(n1970) );
  XOR U85 ( .A(n105), .B(n124), .Z(n115) );
  XOR U86 ( .A(n170), .B(n189), .Z(n180) );
  XOR U87 ( .A(n235), .B(n260), .Z(n245) );
  XOR U88 ( .A(n307), .B(n328), .Z(n317) );
  XOR U89 ( .A(n375), .B(n396), .Z(n385) );
  XOR U90 ( .A(n443), .B(n464), .Z(n453) );
  XOR U91 ( .A(n511), .B(n532), .Z(n521) );
  XOR U92 ( .A(n579), .B(n600), .Z(n589) );
  XOR U93 ( .A(n647), .B(n668), .Z(n657) );
  XOR U94 ( .A(n715), .B(n736), .Z(n725) );
  XOR U95 ( .A(n783), .B(n804), .Z(n793) );
  XOR U96 ( .A(n851), .B(n872), .Z(n861) );
  XOR U97 ( .A(n931), .B(n951), .Z(n940) );
  XOR U98 ( .A(n1007), .B(n1027), .Z(n1016) );
  XOR U99 ( .A(n1083), .B(n1103), .Z(n1092) );
  XOR U100 ( .A(n1159), .B(n1179), .Z(n1168) );
  XOR U101 ( .A(n1235), .B(n1255), .Z(n1244) );
  XOR U102 ( .A(n1311), .B(n1331), .Z(n1320) );
  XOR U103 ( .A(n1387), .B(n1407), .Z(n1396) );
  XOR U104 ( .A(n1463), .B(n1483), .Z(n1472) );
  XOR U105 ( .A(n1539), .B(n1559), .Z(n1548) );
  XOR U106 ( .A(n1615), .B(n1635), .Z(n1624) );
  XOR U107 ( .A(n1691), .B(n1711), .Z(n1700) );
  XOR U108 ( .A(n1767), .B(n1787), .Z(n1776) );
  XOR U109 ( .A(n1843), .B(n1863), .Z(n1852) );
  XNOR U110 ( .A(n1935), .B(n1933), .Z(n1910) );
  XNOR U111 ( .A(n2121), .B(n2120), .Z(n2115) );
  XNOR U112 ( .A(n2073), .B(n2072), .Z(n2051) );
  XNOR U113 ( .A(n1980), .B(n1979), .Z(n1951) );
  XOR U114 ( .A(n2135), .B(n2142), .Z(n2130) );
  AND U115 ( .A(n214), .B(n213), .Z(n181) );
  NAND U116 ( .A(n85), .B(n84), .Z(n46) );
  XNOR U117 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U118 ( .A(n3), .B(n4), .Z(swire[8]) );
  XOR U119 ( .A(n5), .B(n6), .Z(swire[63]) );
  XOR U120 ( .A(n7), .B(n8), .Z(n6) );
  XOR U121 ( .A(n9), .B(n10), .Z(n8) );
  ANDN U122 ( .B(a[63]), .A(n11), .Z(n10) );
  AND U123 ( .A(b[1]), .B(a[62]), .Z(n9) );
  XOR U124 ( .A(n12), .B(n13), .Z(n7) );
  AND U125 ( .A(b[2]), .B(a[61]), .Z(n13) );
  AND U126 ( .A(b[3]), .B(a[60]), .Z(n12) );
  XOR U127 ( .A(n14), .B(n15), .Z(n5) );
  XOR U128 ( .A(n16), .B(n17), .Z(n15) );
  AND U129 ( .A(b[4]), .B(a[59]), .Z(n17) );
  AND U130 ( .A(b[5]), .B(a[58]), .Z(n16) );
  XOR U131 ( .A(n18), .B(n19), .Z(n14) );
  AND U132 ( .A(b[6]), .B(a[57]), .Z(n19) );
  AND U133 ( .A(b[7]), .B(a[56]), .Z(n18) );
  XOR U134 ( .A(n20), .B(n21), .Z(swire[62]) );
  XOR U135 ( .A(n22), .B(n23), .Z(n21) );
  XNOR U136 ( .A(n24), .B(n25), .Z(n23) );
  ANDN U137 ( .B(a[62]), .A(n11), .Z(n24) );
  XOR U138 ( .A(n26), .B(n27), .Z(n22) );
  XNOR U139 ( .A(n25), .B(n28), .Z(n27) );
  XNOR U140 ( .A(n29), .B(n30), .Z(n28) );
  AND U141 ( .A(b[3]), .B(a[59]), .Z(n29) );
  XOR U142 ( .A(n31), .B(n32), .Z(n25) );
  OR U143 ( .A(n33), .B(n34), .Z(n32) );
  XOR U144 ( .A(n35), .B(n36), .Z(n26) );
  XOR U145 ( .A(n37), .B(n38), .Z(n36) );
  AND U146 ( .A(b[4]), .B(a[58]), .Z(n38) );
  AND U147 ( .A(b[5]), .B(a[57]), .Z(n37) );
  XOR U148 ( .A(n39), .B(n40), .Z(n35) );
  AND U149 ( .A(b[6]), .B(a[56]), .Z(n40) );
  AND U150 ( .A(b[7]), .B(a[55]), .Z(n39) );
  XOR U151 ( .A(n41), .B(n42), .Z(n20) );
  XNOR U152 ( .A(n43), .B(n30), .Z(n42) );
  NANDN U153 ( .A(n44), .B(n45), .Z(n30) );
  AND U154 ( .A(b[2]), .B(a[60]), .Z(n43) );
  AND U155 ( .A(b[1]), .B(a[61]), .Z(n41) );
  XNOR U156 ( .A(n46), .B(n47), .Z(swire[61]) );
  XOR U157 ( .A(n45), .B(n48), .Z(n47) );
  XOR U158 ( .A(n44), .B(n46), .Z(n48) );
  NANDN U159 ( .A(n11), .B(a[61]), .Z(n44) );
  XOR U160 ( .A(n33), .B(n34), .Z(n45) );
  XOR U161 ( .A(n31), .B(n49), .Z(n34) );
  NAND U162 ( .A(b[1]), .B(a[60]), .Z(n49) );
  XOR U163 ( .A(n50), .B(n51), .Z(n33) );
  XOR U164 ( .A(n31), .B(n52), .Z(n51) );
  XOR U165 ( .A(n53), .B(n54), .Z(n52) );
  AND U166 ( .A(b[2]), .B(a[59]), .Z(n53) );
  ANDN U167 ( .B(n55), .A(n56), .Z(n31) );
  XOR U168 ( .A(n57), .B(n58), .Z(n50) );
  XNOR U169 ( .A(n54), .B(n59), .Z(n58) );
  XOR U170 ( .A(n60), .B(n61), .Z(n59) );
  XOR U171 ( .A(n62), .B(n63), .Z(n61) );
  XOR U172 ( .A(n64), .B(n65), .Z(n63) );
  XOR U173 ( .A(n66), .B(n67), .Z(n65) );
  AND U174 ( .A(b[5]), .B(a[56]), .Z(n66) );
  XOR U175 ( .A(n68), .B(n69), .Z(n64) );
  AND U176 ( .A(b[6]), .B(a[55]), .Z(n69) );
  AND U177 ( .A(b[7]), .B(a[54]), .Z(n68) );
  XOR U178 ( .A(n70), .B(n67), .Z(n60) );
  XOR U179 ( .A(n71), .B(n72), .Z(n67) );
  NOR U180 ( .A(n73), .B(n74), .Z(n71) );
  AND U181 ( .A(b[4]), .B(a[57]), .Z(n70) );
  XNOR U182 ( .A(n75), .B(n76), .Z(n54) );
  NANDN U183 ( .A(n77), .B(n78), .Z(n76) );
  XOR U184 ( .A(n79), .B(n62), .Z(n57) );
  XNOR U185 ( .A(n80), .B(n81), .Z(n62) );
  AND U186 ( .A(n82), .B(n83), .Z(n80) );
  AND U187 ( .A(b[3]), .B(a[58]), .Z(n79) );
  XNOR U188 ( .A(n84), .B(n85), .Z(swire[60]) );
  XOR U189 ( .A(n55), .B(n86), .Z(n85) );
  XOR U190 ( .A(n56), .B(n84), .Z(n86) );
  NANDN U191 ( .A(n11), .B(a[60]), .Z(n56) );
  XNOR U192 ( .A(n77), .B(n78), .Z(n55) );
  XOR U193 ( .A(n75), .B(n87), .Z(n78) );
  NAND U194 ( .A(b[1]), .B(a[59]), .Z(n87) );
  XOR U195 ( .A(n83), .B(n88), .Z(n77) );
  XOR U196 ( .A(n75), .B(n82), .Z(n88) );
  XNOR U197 ( .A(n89), .B(n81), .Z(n82) );
  AND U198 ( .A(b[2]), .B(a[58]), .Z(n89) );
  NANDN U199 ( .A(n90), .B(n91), .Z(n75) );
  XNOR U200 ( .A(n81), .B(n74), .Z(n92) );
  XOR U201 ( .A(n93), .B(n94), .Z(n74) );
  XOR U202 ( .A(n72), .B(n95), .Z(n94) );
  XOR U203 ( .A(n96), .B(n97), .Z(n95) );
  XNOR U204 ( .A(n98), .B(n99), .Z(n97) );
  AND U205 ( .A(b[5]), .B(a[55]), .Z(n98) );
  XOR U206 ( .A(n100), .B(n101), .Z(n96) );
  AND U207 ( .A(b[6]), .B(a[54]), .Z(n101) );
  AND U208 ( .A(b[7]), .B(a[53]), .Z(n100) );
  XOR U209 ( .A(n102), .B(n99), .Z(n93) );
  XOR U210 ( .A(n103), .B(n104), .Z(n99) );
  NOR U211 ( .A(n105), .B(n106), .Z(n103) );
  AND U212 ( .A(b[4]), .B(a[56]), .Z(n102) );
  XNOR U213 ( .A(n107), .B(n108), .Z(n81) );
  NANDN U214 ( .A(n109), .B(n110), .Z(n108) );
  XNOR U215 ( .A(n111), .B(n72), .Z(n73) );
  XNOR U216 ( .A(n112), .B(n113), .Z(n72) );
  AND U217 ( .A(n114), .B(n115), .Z(n112) );
  AND U218 ( .A(b[3]), .B(a[57]), .Z(n111) );
  XNOR U219 ( .A(n116), .B(n117), .Z(swire[59]) );
  XOR U220 ( .A(n91), .B(n118), .Z(n117) );
  XOR U221 ( .A(n90), .B(n116), .Z(n118) );
  NANDN U222 ( .A(n11), .B(a[59]), .Z(n90) );
  XNOR U223 ( .A(n109), .B(n110), .Z(n91) );
  XOR U224 ( .A(n107), .B(n119), .Z(n110) );
  NAND U225 ( .A(b[1]), .B(a[58]), .Z(n119) );
  XOR U226 ( .A(n115), .B(n120), .Z(n109) );
  XOR U227 ( .A(n107), .B(n114), .Z(n120) );
  XNOR U228 ( .A(n121), .B(n113), .Z(n114) );
  AND U229 ( .A(b[2]), .B(a[57]), .Z(n121) );
  NANDN U230 ( .A(n122), .B(n123), .Z(n107) );
  XNOR U231 ( .A(n113), .B(n106), .Z(n124) );
  XOR U232 ( .A(n125), .B(n126), .Z(n106) );
  XOR U233 ( .A(n104), .B(n127), .Z(n126) );
  XOR U234 ( .A(n128), .B(n129), .Z(n127) );
  XNOR U235 ( .A(n130), .B(n131), .Z(n129) );
  AND U236 ( .A(b[5]), .B(a[54]), .Z(n130) );
  XOR U237 ( .A(n132), .B(n133), .Z(n128) );
  AND U238 ( .A(b[6]), .B(a[53]), .Z(n133) );
  AND U239 ( .A(b[7]), .B(a[52]), .Z(n132) );
  XOR U240 ( .A(n134), .B(n131), .Z(n125) );
  XOR U241 ( .A(n135), .B(n136), .Z(n131) );
  NOR U242 ( .A(n137), .B(n138), .Z(n135) );
  AND U243 ( .A(b[4]), .B(a[55]), .Z(n134) );
  XNOR U244 ( .A(n139), .B(n140), .Z(n113) );
  NANDN U245 ( .A(n141), .B(n142), .Z(n140) );
  XNOR U246 ( .A(n143), .B(n104), .Z(n105) );
  XNOR U247 ( .A(n144), .B(n145), .Z(n104) );
  AND U248 ( .A(n146), .B(n147), .Z(n144) );
  AND U249 ( .A(b[3]), .B(a[56]), .Z(n143) );
  XNOR U250 ( .A(n148), .B(n149), .Z(swire[58]) );
  XOR U251 ( .A(n123), .B(n151), .Z(n149) );
  XNOR U252 ( .A(n122), .B(n150), .Z(n151) );
  IV U253 ( .A(n148), .Z(n150) );
  NANDN U254 ( .A(n11), .B(a[58]), .Z(n122) );
  XNOR U255 ( .A(n141), .B(n142), .Z(n123) );
  XOR U256 ( .A(n139), .B(n152), .Z(n142) );
  NAND U257 ( .A(b[1]), .B(a[57]), .Z(n152) );
  XOR U258 ( .A(n147), .B(n153), .Z(n141) );
  XOR U259 ( .A(n139), .B(n146), .Z(n153) );
  XNOR U260 ( .A(n154), .B(n145), .Z(n146) );
  AND U261 ( .A(b[2]), .B(a[56]), .Z(n154) );
  NANDN U262 ( .A(n155), .B(n156), .Z(n139) );
  XNOR U263 ( .A(n145), .B(n138), .Z(n157) );
  XOR U264 ( .A(n158), .B(n159), .Z(n138) );
  XOR U265 ( .A(n136), .B(n160), .Z(n159) );
  XOR U266 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U267 ( .A(n163), .B(n164), .Z(n162) );
  AND U268 ( .A(b[5]), .B(a[53]), .Z(n163) );
  XOR U269 ( .A(n165), .B(n166), .Z(n161) );
  AND U270 ( .A(b[6]), .B(a[52]), .Z(n166) );
  AND U271 ( .A(b[7]), .B(a[51]), .Z(n165) );
  XOR U272 ( .A(n167), .B(n164), .Z(n158) );
  XOR U273 ( .A(n168), .B(n169), .Z(n164) );
  NOR U274 ( .A(n170), .B(n171), .Z(n168) );
  AND U275 ( .A(b[4]), .B(a[54]), .Z(n167) );
  XNOR U276 ( .A(n172), .B(n173), .Z(n145) );
  NANDN U277 ( .A(n174), .B(n175), .Z(n173) );
  XNOR U278 ( .A(n176), .B(n136), .Z(n137) );
  XNOR U279 ( .A(n177), .B(n178), .Z(n136) );
  AND U280 ( .A(n179), .B(n180), .Z(n177) );
  AND U281 ( .A(b[3]), .B(a[55]), .Z(n176) );
  XNOR U282 ( .A(n181), .B(n182), .Z(swire[57]) );
  XOR U283 ( .A(n156), .B(n183), .Z(n182) );
  XOR U284 ( .A(n155), .B(n181), .Z(n183) );
  NANDN U285 ( .A(n11), .B(a[57]), .Z(n155) );
  XNOR U286 ( .A(n174), .B(n175), .Z(n156) );
  XOR U287 ( .A(n172), .B(n184), .Z(n175) );
  NAND U288 ( .A(b[1]), .B(a[56]), .Z(n184) );
  XOR U289 ( .A(n180), .B(n185), .Z(n174) );
  XOR U290 ( .A(n172), .B(n179), .Z(n185) );
  XNOR U291 ( .A(n186), .B(n178), .Z(n179) );
  AND U292 ( .A(b[2]), .B(a[55]), .Z(n186) );
  NANDN U293 ( .A(n187), .B(n188), .Z(n172) );
  XNOR U294 ( .A(n178), .B(n171), .Z(n189) );
  XOR U295 ( .A(n190), .B(n191), .Z(n171) );
  XOR U296 ( .A(n169), .B(n192), .Z(n191) );
  XOR U297 ( .A(n193), .B(n194), .Z(n192) );
  XNOR U298 ( .A(n195), .B(n196), .Z(n194) );
  AND U299 ( .A(b[5]), .B(a[52]), .Z(n195) );
  XOR U300 ( .A(n197), .B(n198), .Z(n193) );
  AND U301 ( .A(b[6]), .B(a[51]), .Z(n198) );
  AND U302 ( .A(b[7]), .B(a[50]), .Z(n197) );
  XOR U303 ( .A(n199), .B(n196), .Z(n190) );
  XOR U304 ( .A(n200), .B(n201), .Z(n196) );
  NOR U305 ( .A(n202), .B(n203), .Z(n200) );
  AND U306 ( .A(b[4]), .B(a[53]), .Z(n199) );
  XNOR U307 ( .A(n204), .B(n205), .Z(n178) );
  NANDN U308 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U309 ( .A(n208), .B(n169), .Z(n170) );
  XNOR U310 ( .A(n209), .B(n210), .Z(n169) );
  AND U311 ( .A(n211), .B(n212), .Z(n209) );
  AND U312 ( .A(b[3]), .B(a[54]), .Z(n208) );
  XNOR U313 ( .A(n213), .B(n214), .Z(swire[56]) );
  XOR U314 ( .A(n188), .B(n216), .Z(n214) );
  XNOR U315 ( .A(n187), .B(n215), .Z(n216) );
  IV U316 ( .A(n213), .Z(n215) );
  NANDN U317 ( .A(n11), .B(a[56]), .Z(n187) );
  XNOR U318 ( .A(n206), .B(n207), .Z(n188) );
  XOR U319 ( .A(n204), .B(n217), .Z(n207) );
  NAND U320 ( .A(b[1]), .B(a[55]), .Z(n217) );
  XOR U321 ( .A(n212), .B(n218), .Z(n206) );
  XOR U322 ( .A(n204), .B(n211), .Z(n218) );
  XNOR U323 ( .A(n219), .B(n210), .Z(n211) );
  AND U324 ( .A(b[2]), .B(a[54]), .Z(n219) );
  NANDN U325 ( .A(n220), .B(n221), .Z(n204) );
  XNOR U326 ( .A(n210), .B(n203), .Z(n222) );
  XOR U327 ( .A(n223), .B(n224), .Z(n203) );
  XOR U328 ( .A(n201), .B(n225), .Z(n224) );
  XOR U329 ( .A(n226), .B(n227), .Z(n225) );
  XNOR U330 ( .A(n228), .B(n229), .Z(n227) );
  AND U331 ( .A(b[5]), .B(a[51]), .Z(n228) );
  XOR U332 ( .A(n230), .B(n231), .Z(n226) );
  AND U333 ( .A(b[6]), .B(a[50]), .Z(n231) );
  AND U334 ( .A(b[7]), .B(a[49]), .Z(n230) );
  XOR U335 ( .A(n232), .B(n229), .Z(n223) );
  XOR U336 ( .A(n233), .B(n234), .Z(n229) );
  NOR U337 ( .A(n235), .B(n236), .Z(n233) );
  AND U338 ( .A(b[4]), .B(a[52]), .Z(n232) );
  XNOR U339 ( .A(n237), .B(n238), .Z(n210) );
  NANDN U340 ( .A(n239), .B(n240), .Z(n238) );
  XNOR U341 ( .A(n241), .B(n201), .Z(n202) );
  XNOR U342 ( .A(n242), .B(n243), .Z(n201) );
  AND U343 ( .A(n244), .B(n245), .Z(n242) );
  AND U344 ( .A(b[3]), .B(a[53]), .Z(n241) );
  XNOR U345 ( .A(n246), .B(n247), .Z(n213) );
  NOR U346 ( .A(n248), .B(n249), .Z(n246) );
  XOR U347 ( .A(n249), .B(n248), .Z(swire[55]) );
  XOR U348 ( .A(sreg[119]), .B(n247), .Z(n248) );
  XOR U349 ( .A(n221), .B(n250), .Z(n249) );
  XNOR U350 ( .A(n220), .B(n247), .Z(n250) );
  XOR U351 ( .A(n251), .B(n252), .Z(n247) );
  NOR U352 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U353 ( .A(n11), .B(a[55]), .Z(n220) );
  XNOR U354 ( .A(n239), .B(n240), .Z(n221) );
  XOR U355 ( .A(n237), .B(n255), .Z(n240) );
  NAND U356 ( .A(b[1]), .B(a[54]), .Z(n255) );
  XOR U357 ( .A(n245), .B(n256), .Z(n239) );
  XOR U358 ( .A(n237), .B(n244), .Z(n256) );
  XNOR U359 ( .A(n257), .B(n243), .Z(n244) );
  AND U360 ( .A(b[2]), .B(a[53]), .Z(n257) );
  NANDN U361 ( .A(n258), .B(n259), .Z(n237) );
  XNOR U362 ( .A(n243), .B(n236), .Z(n260) );
  XOR U363 ( .A(n261), .B(n262), .Z(n236) );
  XOR U364 ( .A(n234), .B(n263), .Z(n262) );
  XOR U365 ( .A(n264), .B(n265), .Z(n263) );
  XNOR U366 ( .A(n266), .B(n267), .Z(n265) );
  AND U367 ( .A(b[5]), .B(a[50]), .Z(n266) );
  XOR U368 ( .A(n268), .B(n269), .Z(n264) );
  AND U369 ( .A(b[6]), .B(a[49]), .Z(n269) );
  AND U370 ( .A(b[7]), .B(a[48]), .Z(n268) );
  XOR U371 ( .A(n270), .B(n267), .Z(n261) );
  XOR U372 ( .A(n271), .B(n272), .Z(n267) );
  NOR U373 ( .A(n273), .B(n274), .Z(n271) );
  AND U374 ( .A(b[4]), .B(a[51]), .Z(n270) );
  XNOR U375 ( .A(n275), .B(n276), .Z(n243) );
  NANDN U376 ( .A(n277), .B(n278), .Z(n276) );
  XNOR U377 ( .A(n279), .B(n234), .Z(n235) );
  XNOR U378 ( .A(n280), .B(n281), .Z(n234) );
  AND U379 ( .A(n282), .B(n283), .Z(n280) );
  AND U380 ( .A(b[3]), .B(a[52]), .Z(n279) );
  XOR U381 ( .A(n254), .B(n253), .Z(swire[54]) );
  XOR U382 ( .A(sreg[118]), .B(n252), .Z(n253) );
  XOR U383 ( .A(n259), .B(n284), .Z(n254) );
  XNOR U384 ( .A(n258), .B(n252), .Z(n284) );
  XOR U385 ( .A(n285), .B(n286), .Z(n252) );
  NOR U386 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U387 ( .A(n11), .B(a[54]), .Z(n258) );
  XNOR U388 ( .A(n277), .B(n278), .Z(n259) );
  XOR U389 ( .A(n275), .B(n289), .Z(n278) );
  NAND U390 ( .A(b[1]), .B(a[53]), .Z(n289) );
  XOR U391 ( .A(n283), .B(n290), .Z(n277) );
  XOR U392 ( .A(n275), .B(n282), .Z(n290) );
  XNOR U393 ( .A(n291), .B(n281), .Z(n282) );
  AND U394 ( .A(b[2]), .B(a[52]), .Z(n291) );
  NANDN U395 ( .A(n292), .B(n293), .Z(n275) );
  XNOR U396 ( .A(n281), .B(n274), .Z(n294) );
  XOR U397 ( .A(n295), .B(n296), .Z(n274) );
  XOR U398 ( .A(n272), .B(n297), .Z(n296) );
  XOR U399 ( .A(n298), .B(n299), .Z(n297) );
  XNOR U400 ( .A(n300), .B(n301), .Z(n299) );
  AND U401 ( .A(b[5]), .B(a[49]), .Z(n300) );
  XOR U402 ( .A(n302), .B(n303), .Z(n298) );
  AND U403 ( .A(b[6]), .B(a[48]), .Z(n303) );
  AND U404 ( .A(b[7]), .B(a[47]), .Z(n302) );
  XOR U405 ( .A(n304), .B(n301), .Z(n295) );
  XOR U406 ( .A(n305), .B(n306), .Z(n301) );
  NOR U407 ( .A(n307), .B(n308), .Z(n305) );
  AND U408 ( .A(b[4]), .B(a[50]), .Z(n304) );
  XNOR U409 ( .A(n309), .B(n310), .Z(n281) );
  NANDN U410 ( .A(n311), .B(n312), .Z(n310) );
  XNOR U411 ( .A(n313), .B(n272), .Z(n273) );
  XNOR U412 ( .A(n314), .B(n315), .Z(n272) );
  AND U413 ( .A(n316), .B(n317), .Z(n314) );
  AND U414 ( .A(b[3]), .B(a[51]), .Z(n313) );
  XOR U415 ( .A(n288), .B(n287), .Z(swire[53]) );
  XOR U416 ( .A(sreg[117]), .B(n286), .Z(n287) );
  XOR U417 ( .A(n293), .B(n318), .Z(n288) );
  XNOR U418 ( .A(n292), .B(n286), .Z(n318) );
  XOR U419 ( .A(n319), .B(n320), .Z(n286) );
  NOR U420 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U421 ( .A(n11), .B(a[53]), .Z(n292) );
  XNOR U422 ( .A(n311), .B(n312), .Z(n293) );
  XOR U423 ( .A(n309), .B(n323), .Z(n312) );
  NAND U424 ( .A(b[1]), .B(a[52]), .Z(n323) );
  XOR U425 ( .A(n317), .B(n324), .Z(n311) );
  XOR U426 ( .A(n309), .B(n316), .Z(n324) );
  XNOR U427 ( .A(n325), .B(n315), .Z(n316) );
  AND U428 ( .A(b[2]), .B(a[51]), .Z(n325) );
  NANDN U429 ( .A(n326), .B(n327), .Z(n309) );
  XNOR U430 ( .A(n315), .B(n308), .Z(n328) );
  XOR U431 ( .A(n329), .B(n330), .Z(n308) );
  XOR U432 ( .A(n306), .B(n331), .Z(n330) );
  XOR U433 ( .A(n332), .B(n333), .Z(n331) );
  XNOR U434 ( .A(n334), .B(n335), .Z(n333) );
  AND U435 ( .A(b[5]), .B(a[48]), .Z(n334) );
  XOR U436 ( .A(n336), .B(n337), .Z(n332) );
  AND U437 ( .A(b[6]), .B(a[47]), .Z(n337) );
  AND U438 ( .A(b[7]), .B(a[46]), .Z(n336) );
  XOR U439 ( .A(n338), .B(n335), .Z(n329) );
  XOR U440 ( .A(n339), .B(n340), .Z(n335) );
  NOR U441 ( .A(n341), .B(n342), .Z(n339) );
  AND U442 ( .A(b[4]), .B(a[49]), .Z(n338) );
  XNOR U443 ( .A(n343), .B(n344), .Z(n315) );
  NANDN U444 ( .A(n345), .B(n346), .Z(n344) );
  XNOR U445 ( .A(n347), .B(n306), .Z(n307) );
  XNOR U446 ( .A(n348), .B(n349), .Z(n306) );
  AND U447 ( .A(n350), .B(n351), .Z(n348) );
  AND U448 ( .A(b[3]), .B(a[50]), .Z(n347) );
  XOR U449 ( .A(n322), .B(n321), .Z(swire[52]) );
  XOR U450 ( .A(sreg[116]), .B(n320), .Z(n321) );
  XOR U451 ( .A(n327), .B(n352), .Z(n322) );
  XNOR U452 ( .A(n326), .B(n320), .Z(n352) );
  XOR U453 ( .A(n353), .B(n354), .Z(n320) );
  NOR U454 ( .A(n355), .B(n356), .Z(n353) );
  NANDN U455 ( .A(n11), .B(a[52]), .Z(n326) );
  XNOR U456 ( .A(n345), .B(n346), .Z(n327) );
  XOR U457 ( .A(n343), .B(n357), .Z(n346) );
  NAND U458 ( .A(b[1]), .B(a[51]), .Z(n357) );
  XOR U459 ( .A(n351), .B(n358), .Z(n345) );
  XOR U460 ( .A(n343), .B(n350), .Z(n358) );
  XNOR U461 ( .A(n359), .B(n349), .Z(n350) );
  AND U462 ( .A(b[2]), .B(a[50]), .Z(n359) );
  NANDN U463 ( .A(n360), .B(n361), .Z(n343) );
  XNOR U464 ( .A(n349), .B(n342), .Z(n362) );
  XOR U465 ( .A(n363), .B(n364), .Z(n342) );
  XOR U466 ( .A(n340), .B(n365), .Z(n364) );
  XOR U467 ( .A(n366), .B(n367), .Z(n365) );
  XNOR U468 ( .A(n368), .B(n369), .Z(n367) );
  AND U469 ( .A(b[5]), .B(a[47]), .Z(n368) );
  XOR U470 ( .A(n370), .B(n371), .Z(n366) );
  AND U471 ( .A(b[6]), .B(a[46]), .Z(n371) );
  AND U472 ( .A(b[7]), .B(a[45]), .Z(n370) );
  XOR U473 ( .A(n372), .B(n369), .Z(n363) );
  XOR U474 ( .A(n373), .B(n374), .Z(n369) );
  NOR U475 ( .A(n375), .B(n376), .Z(n373) );
  AND U476 ( .A(b[4]), .B(a[48]), .Z(n372) );
  XNOR U477 ( .A(n377), .B(n378), .Z(n349) );
  NANDN U478 ( .A(n379), .B(n380), .Z(n378) );
  XNOR U479 ( .A(n381), .B(n340), .Z(n341) );
  XNOR U480 ( .A(n382), .B(n383), .Z(n340) );
  AND U481 ( .A(n384), .B(n385), .Z(n382) );
  AND U482 ( .A(b[3]), .B(a[49]), .Z(n381) );
  XOR U483 ( .A(n356), .B(n355), .Z(swire[51]) );
  XOR U484 ( .A(sreg[115]), .B(n354), .Z(n355) );
  XOR U485 ( .A(n361), .B(n386), .Z(n356) );
  XNOR U486 ( .A(n360), .B(n354), .Z(n386) );
  XOR U487 ( .A(n387), .B(n388), .Z(n354) );
  NOR U488 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U489 ( .A(n11), .B(a[51]), .Z(n360) );
  XNOR U490 ( .A(n379), .B(n380), .Z(n361) );
  XOR U491 ( .A(n377), .B(n391), .Z(n380) );
  NAND U492 ( .A(b[1]), .B(a[50]), .Z(n391) );
  XOR U493 ( .A(n385), .B(n392), .Z(n379) );
  XOR U494 ( .A(n377), .B(n384), .Z(n392) );
  XNOR U495 ( .A(n393), .B(n383), .Z(n384) );
  AND U496 ( .A(b[2]), .B(a[49]), .Z(n393) );
  NANDN U497 ( .A(n394), .B(n395), .Z(n377) );
  XNOR U498 ( .A(n383), .B(n376), .Z(n396) );
  XOR U499 ( .A(n397), .B(n398), .Z(n376) );
  XOR U500 ( .A(n374), .B(n399), .Z(n398) );
  XOR U501 ( .A(n400), .B(n401), .Z(n399) );
  XNOR U502 ( .A(n402), .B(n403), .Z(n401) );
  AND U503 ( .A(b[5]), .B(a[46]), .Z(n402) );
  XOR U504 ( .A(n404), .B(n405), .Z(n400) );
  AND U505 ( .A(b[6]), .B(a[45]), .Z(n405) );
  AND U506 ( .A(b[7]), .B(a[44]), .Z(n404) );
  XOR U507 ( .A(n406), .B(n403), .Z(n397) );
  XOR U508 ( .A(n407), .B(n408), .Z(n403) );
  NOR U509 ( .A(n409), .B(n410), .Z(n407) );
  AND U510 ( .A(b[4]), .B(a[47]), .Z(n406) );
  XNOR U511 ( .A(n411), .B(n412), .Z(n383) );
  NANDN U512 ( .A(n413), .B(n414), .Z(n412) );
  XNOR U513 ( .A(n415), .B(n374), .Z(n375) );
  XNOR U514 ( .A(n416), .B(n417), .Z(n374) );
  AND U515 ( .A(n418), .B(n419), .Z(n416) );
  AND U516 ( .A(b[3]), .B(a[48]), .Z(n415) );
  XOR U517 ( .A(n390), .B(n389), .Z(swire[50]) );
  XOR U518 ( .A(sreg[114]), .B(n388), .Z(n389) );
  XOR U519 ( .A(n395), .B(n420), .Z(n390) );
  XNOR U520 ( .A(n394), .B(n388), .Z(n420) );
  XOR U521 ( .A(n421), .B(n422), .Z(n388) );
  NOR U522 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U523 ( .A(n11), .B(a[50]), .Z(n394) );
  XNOR U524 ( .A(n413), .B(n414), .Z(n395) );
  XOR U525 ( .A(n411), .B(n425), .Z(n414) );
  NAND U526 ( .A(b[1]), .B(a[49]), .Z(n425) );
  XOR U527 ( .A(n419), .B(n426), .Z(n413) );
  XOR U528 ( .A(n411), .B(n418), .Z(n426) );
  XNOR U529 ( .A(n427), .B(n417), .Z(n418) );
  AND U530 ( .A(b[2]), .B(a[48]), .Z(n427) );
  NANDN U531 ( .A(n428), .B(n429), .Z(n411) );
  XNOR U532 ( .A(n417), .B(n410), .Z(n430) );
  XOR U533 ( .A(n431), .B(n432), .Z(n410) );
  XOR U534 ( .A(n408), .B(n433), .Z(n432) );
  XOR U535 ( .A(n434), .B(n435), .Z(n433) );
  XNOR U536 ( .A(n436), .B(n437), .Z(n435) );
  AND U537 ( .A(b[5]), .B(a[45]), .Z(n436) );
  XOR U538 ( .A(n438), .B(n439), .Z(n434) );
  AND U539 ( .A(b[6]), .B(a[44]), .Z(n439) );
  AND U540 ( .A(b[7]), .B(a[43]), .Z(n438) );
  XOR U541 ( .A(n440), .B(n437), .Z(n431) );
  XOR U542 ( .A(n441), .B(n442), .Z(n437) );
  NOR U543 ( .A(n443), .B(n444), .Z(n441) );
  AND U544 ( .A(b[4]), .B(a[46]), .Z(n440) );
  XNOR U545 ( .A(n445), .B(n446), .Z(n417) );
  NANDN U546 ( .A(n447), .B(n448), .Z(n446) );
  XNOR U547 ( .A(n449), .B(n408), .Z(n409) );
  XNOR U548 ( .A(n450), .B(n451), .Z(n408) );
  AND U549 ( .A(n452), .B(n453), .Z(n450) );
  AND U550 ( .A(b[3]), .B(a[47]), .Z(n449) );
  XOR U551 ( .A(n424), .B(n423), .Z(swire[49]) );
  XOR U552 ( .A(sreg[113]), .B(n422), .Z(n423) );
  XOR U553 ( .A(n429), .B(n454), .Z(n424) );
  XNOR U554 ( .A(n428), .B(n422), .Z(n454) );
  XOR U555 ( .A(n455), .B(n456), .Z(n422) );
  NOR U556 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U557 ( .A(n11), .B(a[49]), .Z(n428) );
  XNOR U558 ( .A(n447), .B(n448), .Z(n429) );
  XOR U559 ( .A(n445), .B(n459), .Z(n448) );
  NAND U560 ( .A(b[1]), .B(a[48]), .Z(n459) );
  XOR U561 ( .A(n453), .B(n460), .Z(n447) );
  XOR U562 ( .A(n445), .B(n452), .Z(n460) );
  XNOR U563 ( .A(n461), .B(n451), .Z(n452) );
  AND U564 ( .A(b[2]), .B(a[47]), .Z(n461) );
  NANDN U565 ( .A(n462), .B(n463), .Z(n445) );
  XNOR U566 ( .A(n451), .B(n444), .Z(n464) );
  XOR U567 ( .A(n465), .B(n466), .Z(n444) );
  XOR U568 ( .A(n442), .B(n467), .Z(n466) );
  XOR U569 ( .A(n468), .B(n469), .Z(n467) );
  XNOR U570 ( .A(n470), .B(n471), .Z(n469) );
  AND U571 ( .A(b[5]), .B(a[44]), .Z(n470) );
  XOR U572 ( .A(n472), .B(n473), .Z(n468) );
  AND U573 ( .A(b[6]), .B(a[43]), .Z(n473) );
  AND U574 ( .A(b[7]), .B(a[42]), .Z(n472) );
  XOR U575 ( .A(n474), .B(n471), .Z(n465) );
  XOR U576 ( .A(n475), .B(n476), .Z(n471) );
  NOR U577 ( .A(n477), .B(n478), .Z(n475) );
  AND U578 ( .A(b[4]), .B(a[45]), .Z(n474) );
  XNOR U579 ( .A(n479), .B(n480), .Z(n451) );
  NANDN U580 ( .A(n481), .B(n482), .Z(n480) );
  XNOR U581 ( .A(n483), .B(n442), .Z(n443) );
  XNOR U582 ( .A(n484), .B(n485), .Z(n442) );
  AND U583 ( .A(n486), .B(n487), .Z(n484) );
  AND U584 ( .A(b[3]), .B(a[46]), .Z(n483) );
  XOR U585 ( .A(n458), .B(n457), .Z(swire[48]) );
  XOR U586 ( .A(sreg[112]), .B(n456), .Z(n457) );
  XOR U587 ( .A(n463), .B(n488), .Z(n458) );
  XNOR U588 ( .A(n462), .B(n456), .Z(n488) );
  XOR U589 ( .A(n489), .B(n490), .Z(n456) );
  NOR U590 ( .A(n491), .B(n492), .Z(n489) );
  NANDN U591 ( .A(n11), .B(a[48]), .Z(n462) );
  XNOR U592 ( .A(n481), .B(n482), .Z(n463) );
  XOR U593 ( .A(n479), .B(n493), .Z(n482) );
  NAND U594 ( .A(b[1]), .B(a[47]), .Z(n493) );
  XOR U595 ( .A(n487), .B(n494), .Z(n481) );
  XOR U596 ( .A(n479), .B(n486), .Z(n494) );
  XNOR U597 ( .A(n495), .B(n485), .Z(n486) );
  AND U598 ( .A(b[2]), .B(a[46]), .Z(n495) );
  NANDN U599 ( .A(n496), .B(n497), .Z(n479) );
  XNOR U600 ( .A(n485), .B(n478), .Z(n498) );
  XOR U601 ( .A(n499), .B(n500), .Z(n478) );
  XOR U602 ( .A(n476), .B(n501), .Z(n500) );
  XOR U603 ( .A(n502), .B(n503), .Z(n501) );
  XNOR U604 ( .A(n504), .B(n505), .Z(n503) );
  AND U605 ( .A(b[5]), .B(a[43]), .Z(n504) );
  XOR U606 ( .A(n506), .B(n507), .Z(n502) );
  AND U607 ( .A(b[6]), .B(a[42]), .Z(n507) );
  AND U608 ( .A(b[7]), .B(a[41]), .Z(n506) );
  XOR U609 ( .A(n508), .B(n505), .Z(n499) );
  XOR U610 ( .A(n509), .B(n510), .Z(n505) );
  NOR U611 ( .A(n511), .B(n512), .Z(n509) );
  AND U612 ( .A(b[4]), .B(a[44]), .Z(n508) );
  XNOR U613 ( .A(n513), .B(n514), .Z(n485) );
  NANDN U614 ( .A(n515), .B(n516), .Z(n514) );
  XNOR U615 ( .A(n517), .B(n476), .Z(n477) );
  XNOR U616 ( .A(n518), .B(n519), .Z(n476) );
  AND U617 ( .A(n520), .B(n521), .Z(n518) );
  AND U618 ( .A(b[3]), .B(a[45]), .Z(n517) );
  XOR U619 ( .A(n492), .B(n491), .Z(swire[47]) );
  XOR U620 ( .A(sreg[111]), .B(n490), .Z(n491) );
  XOR U621 ( .A(n497), .B(n522), .Z(n492) );
  XNOR U622 ( .A(n496), .B(n490), .Z(n522) );
  XOR U623 ( .A(n523), .B(n524), .Z(n490) );
  NOR U624 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U625 ( .A(n11), .B(a[47]), .Z(n496) );
  XNOR U626 ( .A(n515), .B(n516), .Z(n497) );
  XOR U627 ( .A(n513), .B(n527), .Z(n516) );
  NAND U628 ( .A(b[1]), .B(a[46]), .Z(n527) );
  XOR U629 ( .A(n521), .B(n528), .Z(n515) );
  XOR U630 ( .A(n513), .B(n520), .Z(n528) );
  XNOR U631 ( .A(n529), .B(n519), .Z(n520) );
  AND U632 ( .A(b[2]), .B(a[45]), .Z(n529) );
  NANDN U633 ( .A(n530), .B(n531), .Z(n513) );
  XNOR U634 ( .A(n519), .B(n512), .Z(n532) );
  XOR U635 ( .A(n533), .B(n534), .Z(n512) );
  XOR U636 ( .A(n510), .B(n535), .Z(n534) );
  XOR U637 ( .A(n536), .B(n537), .Z(n535) );
  XNOR U638 ( .A(n538), .B(n539), .Z(n537) );
  AND U639 ( .A(b[5]), .B(a[42]), .Z(n538) );
  XOR U640 ( .A(n540), .B(n541), .Z(n536) );
  AND U641 ( .A(b[6]), .B(a[41]), .Z(n541) );
  AND U642 ( .A(b[7]), .B(a[40]), .Z(n540) );
  XOR U643 ( .A(n542), .B(n539), .Z(n533) );
  XOR U644 ( .A(n543), .B(n544), .Z(n539) );
  NOR U645 ( .A(n545), .B(n546), .Z(n543) );
  AND U646 ( .A(b[4]), .B(a[43]), .Z(n542) );
  XNOR U647 ( .A(n547), .B(n548), .Z(n519) );
  NANDN U648 ( .A(n549), .B(n550), .Z(n548) );
  XNOR U649 ( .A(n551), .B(n510), .Z(n511) );
  XNOR U650 ( .A(n552), .B(n553), .Z(n510) );
  AND U651 ( .A(n554), .B(n555), .Z(n552) );
  AND U652 ( .A(b[3]), .B(a[44]), .Z(n551) );
  XOR U653 ( .A(n526), .B(n525), .Z(swire[46]) );
  XOR U654 ( .A(sreg[110]), .B(n524), .Z(n525) );
  XOR U655 ( .A(n531), .B(n556), .Z(n526) );
  XNOR U656 ( .A(n530), .B(n524), .Z(n556) );
  XOR U657 ( .A(n557), .B(n558), .Z(n524) );
  NOR U658 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U659 ( .A(n11), .B(a[46]), .Z(n530) );
  XNOR U660 ( .A(n549), .B(n550), .Z(n531) );
  XOR U661 ( .A(n547), .B(n561), .Z(n550) );
  NAND U662 ( .A(b[1]), .B(a[45]), .Z(n561) );
  XOR U663 ( .A(n555), .B(n562), .Z(n549) );
  XOR U664 ( .A(n547), .B(n554), .Z(n562) );
  XNOR U665 ( .A(n563), .B(n553), .Z(n554) );
  AND U666 ( .A(b[2]), .B(a[44]), .Z(n563) );
  NANDN U667 ( .A(n564), .B(n565), .Z(n547) );
  XNOR U668 ( .A(n553), .B(n546), .Z(n566) );
  XOR U669 ( .A(n567), .B(n568), .Z(n546) );
  XOR U670 ( .A(n544), .B(n569), .Z(n568) );
  XOR U671 ( .A(n570), .B(n571), .Z(n569) );
  XNOR U672 ( .A(n572), .B(n573), .Z(n571) );
  AND U673 ( .A(b[5]), .B(a[41]), .Z(n572) );
  XOR U674 ( .A(n574), .B(n575), .Z(n570) );
  AND U675 ( .A(b[6]), .B(a[40]), .Z(n575) );
  AND U676 ( .A(b[7]), .B(a[39]), .Z(n574) );
  XOR U677 ( .A(n576), .B(n573), .Z(n567) );
  XOR U678 ( .A(n577), .B(n578), .Z(n573) );
  NOR U679 ( .A(n579), .B(n580), .Z(n577) );
  AND U680 ( .A(b[4]), .B(a[42]), .Z(n576) );
  XNOR U681 ( .A(n581), .B(n582), .Z(n553) );
  NANDN U682 ( .A(n583), .B(n584), .Z(n582) );
  XNOR U683 ( .A(n585), .B(n544), .Z(n545) );
  XNOR U684 ( .A(n586), .B(n587), .Z(n544) );
  AND U685 ( .A(n588), .B(n589), .Z(n586) );
  AND U686 ( .A(b[3]), .B(a[43]), .Z(n585) );
  XOR U687 ( .A(n560), .B(n559), .Z(swire[45]) );
  XOR U688 ( .A(sreg[109]), .B(n558), .Z(n559) );
  XOR U689 ( .A(n565), .B(n590), .Z(n560) );
  XNOR U690 ( .A(n564), .B(n558), .Z(n590) );
  XOR U691 ( .A(n591), .B(n592), .Z(n558) );
  NOR U692 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U693 ( .A(n11), .B(a[45]), .Z(n564) );
  XNOR U694 ( .A(n583), .B(n584), .Z(n565) );
  XOR U695 ( .A(n581), .B(n595), .Z(n584) );
  NAND U696 ( .A(b[1]), .B(a[44]), .Z(n595) );
  XOR U697 ( .A(n589), .B(n596), .Z(n583) );
  XOR U698 ( .A(n581), .B(n588), .Z(n596) );
  XNOR U699 ( .A(n597), .B(n587), .Z(n588) );
  AND U700 ( .A(b[2]), .B(a[43]), .Z(n597) );
  NANDN U701 ( .A(n598), .B(n599), .Z(n581) );
  XNOR U702 ( .A(n587), .B(n580), .Z(n600) );
  XOR U703 ( .A(n601), .B(n602), .Z(n580) );
  XOR U704 ( .A(n578), .B(n603), .Z(n602) );
  XOR U705 ( .A(n604), .B(n605), .Z(n603) );
  XNOR U706 ( .A(n606), .B(n607), .Z(n605) );
  AND U707 ( .A(b[5]), .B(a[40]), .Z(n606) );
  XOR U708 ( .A(n608), .B(n609), .Z(n604) );
  AND U709 ( .A(b[6]), .B(a[39]), .Z(n609) );
  AND U710 ( .A(b[7]), .B(a[38]), .Z(n608) );
  XOR U711 ( .A(n610), .B(n607), .Z(n601) );
  XOR U712 ( .A(n611), .B(n612), .Z(n607) );
  NOR U713 ( .A(n613), .B(n614), .Z(n611) );
  AND U714 ( .A(b[4]), .B(a[41]), .Z(n610) );
  XNOR U715 ( .A(n615), .B(n616), .Z(n587) );
  NANDN U716 ( .A(n617), .B(n618), .Z(n616) );
  XNOR U717 ( .A(n619), .B(n578), .Z(n579) );
  XNOR U718 ( .A(n620), .B(n621), .Z(n578) );
  AND U719 ( .A(n622), .B(n623), .Z(n620) );
  AND U720 ( .A(b[3]), .B(a[42]), .Z(n619) );
  XOR U721 ( .A(n594), .B(n593), .Z(swire[44]) );
  XOR U722 ( .A(sreg[108]), .B(n592), .Z(n593) );
  XOR U723 ( .A(n599), .B(n624), .Z(n594) );
  XNOR U724 ( .A(n598), .B(n592), .Z(n624) );
  XOR U725 ( .A(n625), .B(n626), .Z(n592) );
  NOR U726 ( .A(n627), .B(n628), .Z(n625) );
  NANDN U727 ( .A(n11), .B(a[44]), .Z(n598) );
  XNOR U728 ( .A(n617), .B(n618), .Z(n599) );
  XOR U729 ( .A(n615), .B(n629), .Z(n618) );
  NAND U730 ( .A(b[1]), .B(a[43]), .Z(n629) );
  XOR U731 ( .A(n623), .B(n630), .Z(n617) );
  XOR U732 ( .A(n615), .B(n622), .Z(n630) );
  XNOR U733 ( .A(n631), .B(n621), .Z(n622) );
  AND U734 ( .A(b[2]), .B(a[42]), .Z(n631) );
  NANDN U735 ( .A(n632), .B(n633), .Z(n615) );
  XNOR U736 ( .A(n621), .B(n614), .Z(n634) );
  XOR U737 ( .A(n635), .B(n636), .Z(n614) );
  XOR U738 ( .A(n612), .B(n637), .Z(n636) );
  XOR U739 ( .A(n638), .B(n639), .Z(n637) );
  XNOR U740 ( .A(n640), .B(n641), .Z(n639) );
  AND U741 ( .A(b[5]), .B(a[39]), .Z(n640) );
  XOR U742 ( .A(n642), .B(n643), .Z(n638) );
  AND U743 ( .A(b[6]), .B(a[38]), .Z(n643) );
  AND U744 ( .A(b[7]), .B(a[37]), .Z(n642) );
  XOR U745 ( .A(n644), .B(n641), .Z(n635) );
  XOR U746 ( .A(n645), .B(n646), .Z(n641) );
  NOR U747 ( .A(n647), .B(n648), .Z(n645) );
  AND U748 ( .A(b[4]), .B(a[40]), .Z(n644) );
  XNOR U749 ( .A(n649), .B(n650), .Z(n621) );
  NANDN U750 ( .A(n651), .B(n652), .Z(n650) );
  XNOR U751 ( .A(n653), .B(n612), .Z(n613) );
  XNOR U752 ( .A(n654), .B(n655), .Z(n612) );
  AND U753 ( .A(n656), .B(n657), .Z(n654) );
  AND U754 ( .A(b[3]), .B(a[41]), .Z(n653) );
  XOR U755 ( .A(n628), .B(n627), .Z(swire[43]) );
  XOR U756 ( .A(sreg[107]), .B(n626), .Z(n627) );
  XOR U757 ( .A(n633), .B(n658), .Z(n628) );
  XNOR U758 ( .A(n632), .B(n626), .Z(n658) );
  XOR U759 ( .A(n659), .B(n660), .Z(n626) );
  NOR U760 ( .A(n661), .B(n662), .Z(n659) );
  NANDN U761 ( .A(n11), .B(a[43]), .Z(n632) );
  XNOR U762 ( .A(n651), .B(n652), .Z(n633) );
  XOR U763 ( .A(n649), .B(n663), .Z(n652) );
  NAND U764 ( .A(b[1]), .B(a[42]), .Z(n663) );
  XOR U765 ( .A(n657), .B(n664), .Z(n651) );
  XOR U766 ( .A(n649), .B(n656), .Z(n664) );
  XNOR U767 ( .A(n665), .B(n655), .Z(n656) );
  AND U768 ( .A(b[2]), .B(a[41]), .Z(n665) );
  NANDN U769 ( .A(n666), .B(n667), .Z(n649) );
  XNOR U770 ( .A(n655), .B(n648), .Z(n668) );
  XOR U771 ( .A(n669), .B(n670), .Z(n648) );
  XOR U772 ( .A(n646), .B(n671), .Z(n670) );
  XOR U773 ( .A(n672), .B(n673), .Z(n671) );
  XNOR U774 ( .A(n674), .B(n675), .Z(n673) );
  AND U775 ( .A(b[5]), .B(a[38]), .Z(n674) );
  XOR U776 ( .A(n676), .B(n677), .Z(n672) );
  AND U777 ( .A(b[6]), .B(a[37]), .Z(n677) );
  AND U778 ( .A(b[7]), .B(a[36]), .Z(n676) );
  XOR U779 ( .A(n678), .B(n675), .Z(n669) );
  XOR U780 ( .A(n679), .B(n680), .Z(n675) );
  NOR U781 ( .A(n681), .B(n682), .Z(n679) );
  AND U782 ( .A(b[4]), .B(a[39]), .Z(n678) );
  XNOR U783 ( .A(n683), .B(n684), .Z(n655) );
  NANDN U784 ( .A(n685), .B(n686), .Z(n684) );
  XNOR U785 ( .A(n687), .B(n646), .Z(n647) );
  XNOR U786 ( .A(n688), .B(n689), .Z(n646) );
  AND U787 ( .A(n690), .B(n691), .Z(n688) );
  AND U788 ( .A(b[3]), .B(a[40]), .Z(n687) );
  XOR U789 ( .A(n662), .B(n661), .Z(swire[42]) );
  XOR U790 ( .A(sreg[106]), .B(n660), .Z(n661) );
  XOR U791 ( .A(n667), .B(n692), .Z(n662) );
  XNOR U792 ( .A(n666), .B(n660), .Z(n692) );
  XOR U793 ( .A(n693), .B(n694), .Z(n660) );
  NOR U794 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U795 ( .A(n11), .B(a[42]), .Z(n666) );
  XNOR U796 ( .A(n685), .B(n686), .Z(n667) );
  XOR U797 ( .A(n683), .B(n697), .Z(n686) );
  NAND U798 ( .A(b[1]), .B(a[41]), .Z(n697) );
  XOR U799 ( .A(n691), .B(n698), .Z(n685) );
  XOR U800 ( .A(n683), .B(n690), .Z(n698) );
  XNOR U801 ( .A(n699), .B(n689), .Z(n690) );
  AND U802 ( .A(b[2]), .B(a[40]), .Z(n699) );
  NANDN U803 ( .A(n700), .B(n701), .Z(n683) );
  XNOR U804 ( .A(n689), .B(n682), .Z(n702) );
  XOR U805 ( .A(n703), .B(n704), .Z(n682) );
  XOR U806 ( .A(n680), .B(n705), .Z(n704) );
  XOR U807 ( .A(n706), .B(n707), .Z(n705) );
  XNOR U808 ( .A(n708), .B(n709), .Z(n707) );
  AND U809 ( .A(b[5]), .B(a[37]), .Z(n708) );
  XOR U810 ( .A(n710), .B(n711), .Z(n706) );
  AND U811 ( .A(b[6]), .B(a[36]), .Z(n711) );
  AND U812 ( .A(b[7]), .B(a[35]), .Z(n710) );
  XOR U813 ( .A(n712), .B(n709), .Z(n703) );
  XOR U814 ( .A(n713), .B(n714), .Z(n709) );
  NOR U815 ( .A(n715), .B(n716), .Z(n713) );
  AND U816 ( .A(b[4]), .B(a[38]), .Z(n712) );
  XNOR U817 ( .A(n717), .B(n718), .Z(n689) );
  NANDN U818 ( .A(n719), .B(n720), .Z(n718) );
  XNOR U819 ( .A(n721), .B(n680), .Z(n681) );
  XNOR U820 ( .A(n722), .B(n723), .Z(n680) );
  AND U821 ( .A(n724), .B(n725), .Z(n722) );
  AND U822 ( .A(b[3]), .B(a[39]), .Z(n721) );
  XOR U823 ( .A(n696), .B(n695), .Z(swire[41]) );
  XOR U824 ( .A(sreg[105]), .B(n694), .Z(n695) );
  XOR U825 ( .A(n701), .B(n726), .Z(n696) );
  XNOR U826 ( .A(n700), .B(n694), .Z(n726) );
  XOR U827 ( .A(n727), .B(n728), .Z(n694) );
  NOR U828 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U829 ( .A(n11), .B(a[41]), .Z(n700) );
  XNOR U830 ( .A(n719), .B(n720), .Z(n701) );
  XOR U831 ( .A(n717), .B(n731), .Z(n720) );
  NAND U832 ( .A(b[1]), .B(a[40]), .Z(n731) );
  XOR U833 ( .A(n725), .B(n732), .Z(n719) );
  XOR U834 ( .A(n717), .B(n724), .Z(n732) );
  XNOR U835 ( .A(n733), .B(n723), .Z(n724) );
  AND U836 ( .A(b[2]), .B(a[39]), .Z(n733) );
  NANDN U837 ( .A(n734), .B(n735), .Z(n717) );
  XNOR U838 ( .A(n723), .B(n716), .Z(n736) );
  XOR U839 ( .A(n737), .B(n738), .Z(n716) );
  XOR U840 ( .A(n714), .B(n739), .Z(n738) );
  XOR U841 ( .A(n740), .B(n741), .Z(n739) );
  XNOR U842 ( .A(n742), .B(n743), .Z(n741) );
  AND U843 ( .A(b[5]), .B(a[36]), .Z(n742) );
  XOR U844 ( .A(n744), .B(n745), .Z(n740) );
  AND U845 ( .A(b[6]), .B(a[35]), .Z(n745) );
  AND U846 ( .A(b[7]), .B(a[34]), .Z(n744) );
  XOR U847 ( .A(n746), .B(n743), .Z(n737) );
  XOR U848 ( .A(n747), .B(n748), .Z(n743) );
  NOR U849 ( .A(n749), .B(n750), .Z(n747) );
  AND U850 ( .A(b[4]), .B(a[37]), .Z(n746) );
  XNOR U851 ( .A(n751), .B(n752), .Z(n723) );
  NANDN U852 ( .A(n753), .B(n754), .Z(n752) );
  XNOR U853 ( .A(n755), .B(n714), .Z(n715) );
  XNOR U854 ( .A(n756), .B(n757), .Z(n714) );
  AND U855 ( .A(n758), .B(n759), .Z(n756) );
  AND U856 ( .A(b[3]), .B(a[38]), .Z(n755) );
  XOR U857 ( .A(n730), .B(n729), .Z(swire[40]) );
  XOR U858 ( .A(sreg[104]), .B(n728), .Z(n729) );
  XOR U859 ( .A(n735), .B(n760), .Z(n730) );
  XNOR U860 ( .A(n734), .B(n728), .Z(n760) );
  XOR U861 ( .A(n761), .B(n762), .Z(n728) );
  NOR U862 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U863 ( .A(n11), .B(a[40]), .Z(n734) );
  XNOR U864 ( .A(n753), .B(n754), .Z(n735) );
  XOR U865 ( .A(n751), .B(n765), .Z(n754) );
  NAND U866 ( .A(b[1]), .B(a[39]), .Z(n765) );
  XOR U867 ( .A(n759), .B(n766), .Z(n753) );
  XOR U868 ( .A(n751), .B(n758), .Z(n766) );
  XNOR U869 ( .A(n767), .B(n757), .Z(n758) );
  AND U870 ( .A(b[2]), .B(a[38]), .Z(n767) );
  NANDN U871 ( .A(n768), .B(n769), .Z(n751) );
  XNOR U872 ( .A(n757), .B(n750), .Z(n770) );
  XOR U873 ( .A(n771), .B(n772), .Z(n750) );
  XOR U874 ( .A(n748), .B(n773), .Z(n772) );
  XOR U875 ( .A(n774), .B(n775), .Z(n773) );
  XNOR U876 ( .A(n776), .B(n777), .Z(n775) );
  AND U877 ( .A(b[5]), .B(a[35]), .Z(n776) );
  XOR U878 ( .A(n778), .B(n779), .Z(n774) );
  AND U879 ( .A(b[6]), .B(a[34]), .Z(n779) );
  AND U880 ( .A(b[7]), .B(a[33]), .Z(n778) );
  XOR U881 ( .A(n780), .B(n777), .Z(n771) );
  XOR U882 ( .A(n781), .B(n782), .Z(n777) );
  NOR U883 ( .A(n783), .B(n784), .Z(n781) );
  AND U884 ( .A(b[4]), .B(a[36]), .Z(n780) );
  XNOR U885 ( .A(n785), .B(n786), .Z(n757) );
  NANDN U886 ( .A(n787), .B(n788), .Z(n786) );
  XNOR U887 ( .A(n789), .B(n748), .Z(n749) );
  XNOR U888 ( .A(n790), .B(n791), .Z(n748) );
  AND U889 ( .A(n792), .B(n793), .Z(n790) );
  AND U890 ( .A(b[3]), .B(a[37]), .Z(n789) );
  XOR U891 ( .A(n764), .B(n763), .Z(swire[39]) );
  XOR U892 ( .A(sreg[103]), .B(n762), .Z(n763) );
  XOR U893 ( .A(n769), .B(n794), .Z(n764) );
  XNOR U894 ( .A(n768), .B(n762), .Z(n794) );
  XOR U895 ( .A(n795), .B(n796), .Z(n762) );
  NOR U896 ( .A(n797), .B(n798), .Z(n795) );
  NANDN U897 ( .A(n11), .B(a[39]), .Z(n768) );
  XNOR U898 ( .A(n787), .B(n788), .Z(n769) );
  XOR U899 ( .A(n785), .B(n799), .Z(n788) );
  NAND U900 ( .A(b[1]), .B(a[38]), .Z(n799) );
  XOR U901 ( .A(n793), .B(n800), .Z(n787) );
  XOR U902 ( .A(n785), .B(n792), .Z(n800) );
  XNOR U903 ( .A(n801), .B(n791), .Z(n792) );
  AND U904 ( .A(b[2]), .B(a[37]), .Z(n801) );
  NANDN U905 ( .A(n802), .B(n803), .Z(n785) );
  XNOR U906 ( .A(n791), .B(n784), .Z(n804) );
  XOR U907 ( .A(n805), .B(n806), .Z(n784) );
  XOR U908 ( .A(n782), .B(n807), .Z(n806) );
  XOR U909 ( .A(n808), .B(n809), .Z(n807) );
  XNOR U910 ( .A(n810), .B(n811), .Z(n809) );
  AND U911 ( .A(b[5]), .B(a[34]), .Z(n810) );
  XOR U912 ( .A(n812), .B(n813), .Z(n808) );
  AND U913 ( .A(b[6]), .B(a[33]), .Z(n813) );
  AND U914 ( .A(b[7]), .B(a[32]), .Z(n812) );
  XOR U915 ( .A(n814), .B(n811), .Z(n805) );
  XOR U916 ( .A(n815), .B(n816), .Z(n811) );
  NOR U917 ( .A(n817), .B(n818), .Z(n815) );
  AND U918 ( .A(b[4]), .B(a[35]), .Z(n814) );
  XNOR U919 ( .A(n819), .B(n820), .Z(n791) );
  NANDN U920 ( .A(n821), .B(n822), .Z(n820) );
  XNOR U921 ( .A(n823), .B(n782), .Z(n783) );
  XNOR U922 ( .A(n824), .B(n825), .Z(n782) );
  AND U923 ( .A(n826), .B(n827), .Z(n824) );
  AND U924 ( .A(b[3]), .B(a[36]), .Z(n823) );
  XOR U925 ( .A(n798), .B(n797), .Z(swire[38]) );
  XOR U926 ( .A(sreg[102]), .B(n796), .Z(n797) );
  XOR U927 ( .A(n803), .B(n828), .Z(n798) );
  XNOR U928 ( .A(n802), .B(n796), .Z(n828) );
  XOR U929 ( .A(n829), .B(n830), .Z(n796) );
  NOR U930 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U931 ( .A(n11), .B(a[38]), .Z(n802) );
  XNOR U932 ( .A(n821), .B(n822), .Z(n803) );
  XOR U933 ( .A(n819), .B(n833), .Z(n822) );
  NAND U934 ( .A(b[1]), .B(a[37]), .Z(n833) );
  XOR U935 ( .A(n827), .B(n834), .Z(n821) );
  XOR U936 ( .A(n819), .B(n826), .Z(n834) );
  XNOR U937 ( .A(n835), .B(n825), .Z(n826) );
  AND U938 ( .A(b[2]), .B(a[36]), .Z(n835) );
  NANDN U939 ( .A(n836), .B(n837), .Z(n819) );
  XNOR U940 ( .A(n825), .B(n818), .Z(n838) );
  XOR U941 ( .A(n839), .B(n840), .Z(n818) );
  XOR U942 ( .A(n816), .B(n841), .Z(n840) );
  XOR U943 ( .A(n842), .B(n843), .Z(n841) );
  XNOR U944 ( .A(n844), .B(n845), .Z(n843) );
  AND U945 ( .A(b[5]), .B(a[33]), .Z(n844) );
  XOR U946 ( .A(n846), .B(n847), .Z(n842) );
  AND U947 ( .A(b[6]), .B(a[32]), .Z(n847) );
  AND U948 ( .A(b[7]), .B(a[31]), .Z(n846) );
  XOR U949 ( .A(n848), .B(n845), .Z(n839) );
  XOR U950 ( .A(n849), .B(n850), .Z(n845) );
  NOR U951 ( .A(n851), .B(n852), .Z(n849) );
  AND U952 ( .A(b[4]), .B(a[34]), .Z(n848) );
  XNOR U953 ( .A(n853), .B(n854), .Z(n825) );
  NANDN U954 ( .A(n855), .B(n856), .Z(n854) );
  XNOR U955 ( .A(n857), .B(n816), .Z(n817) );
  XNOR U956 ( .A(n858), .B(n859), .Z(n816) );
  AND U957 ( .A(n860), .B(n861), .Z(n858) );
  AND U958 ( .A(b[3]), .B(a[35]), .Z(n857) );
  XOR U959 ( .A(n832), .B(n831), .Z(swire[37]) );
  XOR U960 ( .A(sreg[101]), .B(n830), .Z(n831) );
  XOR U961 ( .A(n837), .B(n862), .Z(n832) );
  XNOR U962 ( .A(n836), .B(n830), .Z(n862) );
  XOR U963 ( .A(n863), .B(n864), .Z(n830) );
  NOR U964 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U965 ( .A(n11), .B(a[37]), .Z(n836) );
  XNOR U966 ( .A(n855), .B(n856), .Z(n837) );
  XOR U967 ( .A(n853), .B(n867), .Z(n856) );
  NAND U968 ( .A(b[1]), .B(a[36]), .Z(n867) );
  XOR U969 ( .A(n861), .B(n868), .Z(n855) );
  XOR U970 ( .A(n853), .B(n860), .Z(n868) );
  XNOR U971 ( .A(n869), .B(n859), .Z(n860) );
  AND U972 ( .A(b[2]), .B(a[35]), .Z(n869) );
  NANDN U973 ( .A(n870), .B(n871), .Z(n853) );
  XNOR U974 ( .A(n859), .B(n852), .Z(n872) );
  XOR U975 ( .A(n873), .B(n874), .Z(n852) );
  XOR U976 ( .A(n850), .B(n875), .Z(n874) );
  XOR U977 ( .A(n876), .B(n877), .Z(n875) );
  XOR U978 ( .A(n878), .B(n879), .Z(n877) );
  XOR U979 ( .A(n880), .B(n881), .Z(n879) );
  XOR U980 ( .A(n882), .B(n883), .Z(n881) );
  NAND U981 ( .A(b[6]), .B(a[31]), .Z(n883) );
  AND U982 ( .A(b[7]), .B(a[30]), .Z(n882) );
  XOR U983 ( .A(n884), .B(n880), .Z(n876) );
  XOR U984 ( .A(n885), .B(n886), .Z(n880) );
  NOR U985 ( .A(n887), .B(n888), .Z(n885) );
  AND U986 ( .A(b[5]), .B(a[32]), .Z(n884) );
  XOR U987 ( .A(n889), .B(n878), .Z(n873) );
  XOR U988 ( .A(n890), .B(n891), .Z(n878) );
  ANDN U989 ( .B(n892), .A(n893), .Z(n890) );
  AND U990 ( .A(b[4]), .B(a[33]), .Z(n889) );
  XNOR U991 ( .A(n894), .B(n895), .Z(n859) );
  NANDN U992 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U993 ( .A(n898), .B(n850), .Z(n851) );
  XNOR U994 ( .A(n899), .B(n900), .Z(n850) );
  AND U995 ( .A(n901), .B(n902), .Z(n899) );
  AND U996 ( .A(b[3]), .B(a[34]), .Z(n898) );
  XOR U997 ( .A(n866), .B(n865), .Z(swire[36]) );
  XOR U998 ( .A(sreg[100]), .B(n864), .Z(n865) );
  XOR U999 ( .A(n871), .B(n903), .Z(n866) );
  XNOR U1000 ( .A(n870), .B(n864), .Z(n903) );
  XOR U1001 ( .A(n904), .B(n905), .Z(n864) );
  NOR U1002 ( .A(n906), .B(n907), .Z(n904) );
  NANDN U1003 ( .A(n11), .B(a[36]), .Z(n870) );
  XNOR U1004 ( .A(n896), .B(n897), .Z(n871) );
  XOR U1005 ( .A(n894), .B(n908), .Z(n897) );
  NAND U1006 ( .A(b[1]), .B(a[35]), .Z(n908) );
  XOR U1007 ( .A(n902), .B(n909), .Z(n896) );
  XOR U1008 ( .A(n894), .B(n901), .Z(n909) );
  XNOR U1009 ( .A(n910), .B(n900), .Z(n901) );
  AND U1010 ( .A(b[2]), .B(a[34]), .Z(n910) );
  NANDN U1011 ( .A(n911), .B(n912), .Z(n894) );
  XOR U1012 ( .A(n900), .B(n892), .Z(n913) );
  XOR U1013 ( .A(n891), .B(n888), .Z(n914) );
  XOR U1014 ( .A(n915), .B(n916), .Z(n888) );
  XOR U1015 ( .A(n886), .B(n917), .Z(n916) );
  XOR U1016 ( .A(n918), .B(n919), .Z(n917) );
  XOR U1017 ( .A(n920), .B(n921), .Z(n919) );
  NAND U1018 ( .A(b[6]), .B(a[30]), .Z(n921) );
  AND U1019 ( .A(b[7]), .B(a[29]), .Z(n920) );
  XOR U1020 ( .A(n922), .B(n918), .Z(n915) );
  XOR U1021 ( .A(n923), .B(n924), .Z(n918) );
  NOR U1022 ( .A(n925), .B(n926), .Z(n923) );
  AND U1023 ( .A(b[5]), .B(a[31]), .Z(n922) );
  XNOR U1024 ( .A(n927), .B(n886), .Z(n887) );
  XOR U1025 ( .A(n928), .B(n929), .Z(n886) );
  ANDN U1026 ( .B(n930), .A(n931), .Z(n928) );
  AND U1027 ( .A(b[4]), .B(a[32]), .Z(n927) );
  XNOR U1028 ( .A(n932), .B(n933), .Z(n900) );
  NANDN U1029 ( .A(n934), .B(n935), .Z(n933) );
  XNOR U1030 ( .A(n936), .B(n891), .Z(n893) );
  XNOR U1031 ( .A(n937), .B(n938), .Z(n891) );
  AND U1032 ( .A(n939), .B(n940), .Z(n937) );
  AND U1033 ( .A(b[3]), .B(a[33]), .Z(n936) );
  XOR U1034 ( .A(n907), .B(n906), .Z(swire[35]) );
  XOR U1035 ( .A(sreg[99]), .B(n905), .Z(n906) );
  XOR U1036 ( .A(n912), .B(n941), .Z(n907) );
  XNOR U1037 ( .A(n911), .B(n905), .Z(n941) );
  XOR U1038 ( .A(n942), .B(n943), .Z(n905) );
  NOR U1039 ( .A(n944), .B(n945), .Z(n942) );
  NANDN U1040 ( .A(n11), .B(a[35]), .Z(n911) );
  XNOR U1041 ( .A(n934), .B(n935), .Z(n912) );
  XOR U1042 ( .A(n932), .B(n946), .Z(n935) );
  NAND U1043 ( .A(b[1]), .B(a[34]), .Z(n946) );
  XOR U1044 ( .A(n940), .B(n947), .Z(n934) );
  XOR U1045 ( .A(n932), .B(n939), .Z(n947) );
  XNOR U1046 ( .A(n948), .B(n938), .Z(n939) );
  AND U1047 ( .A(b[2]), .B(a[33]), .Z(n948) );
  NANDN U1048 ( .A(n949), .B(n950), .Z(n932) );
  XOR U1049 ( .A(n938), .B(n930), .Z(n951) );
  XOR U1050 ( .A(n929), .B(n926), .Z(n952) );
  XOR U1051 ( .A(n953), .B(n954), .Z(n926) );
  XOR U1052 ( .A(n924), .B(n955), .Z(n954) );
  XOR U1053 ( .A(n956), .B(n957), .Z(n955) );
  XOR U1054 ( .A(n958), .B(n959), .Z(n957) );
  NAND U1055 ( .A(b[6]), .B(a[29]), .Z(n959) );
  AND U1056 ( .A(b[7]), .B(a[28]), .Z(n958) );
  XOR U1057 ( .A(n960), .B(n956), .Z(n953) );
  XOR U1058 ( .A(n961), .B(n962), .Z(n956) );
  NOR U1059 ( .A(n963), .B(n964), .Z(n961) );
  AND U1060 ( .A(b[5]), .B(a[30]), .Z(n960) );
  XNOR U1061 ( .A(n965), .B(n924), .Z(n925) );
  XOR U1062 ( .A(n966), .B(n967), .Z(n924) );
  ANDN U1063 ( .B(n968), .A(n969), .Z(n966) );
  AND U1064 ( .A(b[4]), .B(a[31]), .Z(n965) );
  XNOR U1065 ( .A(n970), .B(n971), .Z(n938) );
  NANDN U1066 ( .A(n972), .B(n973), .Z(n971) );
  XNOR U1067 ( .A(n974), .B(n929), .Z(n931) );
  XNOR U1068 ( .A(n975), .B(n976), .Z(n929) );
  AND U1069 ( .A(n977), .B(n978), .Z(n975) );
  AND U1070 ( .A(b[3]), .B(a[32]), .Z(n974) );
  XOR U1071 ( .A(n945), .B(n944), .Z(swire[34]) );
  XOR U1072 ( .A(sreg[98]), .B(n943), .Z(n944) );
  XOR U1073 ( .A(n950), .B(n979), .Z(n945) );
  XNOR U1074 ( .A(n949), .B(n943), .Z(n979) );
  XOR U1075 ( .A(n980), .B(n981), .Z(n943) );
  NOR U1076 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1077 ( .A(n11), .B(a[34]), .Z(n949) );
  XNOR U1078 ( .A(n972), .B(n973), .Z(n950) );
  XOR U1079 ( .A(n970), .B(n984), .Z(n973) );
  NAND U1080 ( .A(b[1]), .B(a[33]), .Z(n984) );
  XOR U1081 ( .A(n978), .B(n985), .Z(n972) );
  XOR U1082 ( .A(n970), .B(n977), .Z(n985) );
  XNOR U1083 ( .A(n986), .B(n976), .Z(n977) );
  AND U1084 ( .A(b[2]), .B(a[32]), .Z(n986) );
  NANDN U1085 ( .A(n987), .B(n988), .Z(n970) );
  XOR U1086 ( .A(n976), .B(n968), .Z(n989) );
  XOR U1087 ( .A(n967), .B(n964), .Z(n990) );
  XOR U1088 ( .A(n991), .B(n992), .Z(n964) );
  XOR U1089 ( .A(n962), .B(n993), .Z(n992) );
  XOR U1090 ( .A(n994), .B(n995), .Z(n993) );
  XOR U1091 ( .A(n996), .B(n997), .Z(n995) );
  NAND U1092 ( .A(b[6]), .B(a[28]), .Z(n997) );
  AND U1093 ( .A(b[7]), .B(a[27]), .Z(n996) );
  XOR U1094 ( .A(n998), .B(n994), .Z(n991) );
  XOR U1095 ( .A(n999), .B(n1000), .Z(n994) );
  NOR U1096 ( .A(n1001), .B(n1002), .Z(n999) );
  AND U1097 ( .A(b[5]), .B(a[29]), .Z(n998) );
  XNOR U1098 ( .A(n1003), .B(n962), .Z(n963) );
  XOR U1099 ( .A(n1004), .B(n1005), .Z(n962) );
  ANDN U1100 ( .B(n1006), .A(n1007), .Z(n1004) );
  AND U1101 ( .A(b[4]), .B(a[30]), .Z(n1003) );
  XNOR U1102 ( .A(n1008), .B(n1009), .Z(n976) );
  NANDN U1103 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U1104 ( .A(n1012), .B(n967), .Z(n969) );
  XNOR U1105 ( .A(n1013), .B(n1014), .Z(n967) );
  AND U1106 ( .A(n1015), .B(n1016), .Z(n1013) );
  AND U1107 ( .A(b[3]), .B(a[31]), .Z(n1012) );
  XOR U1108 ( .A(n983), .B(n982), .Z(swire[33]) );
  XOR U1109 ( .A(sreg[97]), .B(n981), .Z(n982) );
  XOR U1110 ( .A(n988), .B(n1017), .Z(n983) );
  XNOR U1111 ( .A(n987), .B(n981), .Z(n1017) );
  XOR U1112 ( .A(n1018), .B(n1019), .Z(n981) );
  NOR U1113 ( .A(n1020), .B(n1021), .Z(n1018) );
  NANDN U1114 ( .A(n11), .B(a[33]), .Z(n987) );
  XNOR U1115 ( .A(n1010), .B(n1011), .Z(n988) );
  XOR U1116 ( .A(n1008), .B(n1022), .Z(n1011) );
  NAND U1117 ( .A(b[1]), .B(a[32]), .Z(n1022) );
  XOR U1118 ( .A(n1016), .B(n1023), .Z(n1010) );
  XOR U1119 ( .A(n1008), .B(n1015), .Z(n1023) );
  XNOR U1120 ( .A(n1024), .B(n1014), .Z(n1015) );
  AND U1121 ( .A(b[2]), .B(a[31]), .Z(n1024) );
  NANDN U1122 ( .A(n1025), .B(n1026), .Z(n1008) );
  XOR U1123 ( .A(n1014), .B(n1006), .Z(n1027) );
  XOR U1124 ( .A(n1005), .B(n1002), .Z(n1028) );
  XOR U1125 ( .A(n1029), .B(n1030), .Z(n1002) );
  XOR U1126 ( .A(n1000), .B(n1031), .Z(n1030) );
  XOR U1127 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR U1128 ( .A(n1034), .B(n1035), .Z(n1033) );
  NAND U1129 ( .A(b[6]), .B(a[27]), .Z(n1035) );
  AND U1130 ( .A(b[7]), .B(a[26]), .Z(n1034) );
  XOR U1131 ( .A(n1036), .B(n1032), .Z(n1029) );
  XOR U1132 ( .A(n1037), .B(n1038), .Z(n1032) );
  NOR U1133 ( .A(n1039), .B(n1040), .Z(n1037) );
  AND U1134 ( .A(b[5]), .B(a[28]), .Z(n1036) );
  XNOR U1135 ( .A(n1041), .B(n1000), .Z(n1001) );
  XOR U1136 ( .A(n1042), .B(n1043), .Z(n1000) );
  ANDN U1137 ( .B(n1044), .A(n1045), .Z(n1042) );
  AND U1138 ( .A(b[4]), .B(a[29]), .Z(n1041) );
  XNOR U1139 ( .A(n1046), .B(n1047), .Z(n1014) );
  NANDN U1140 ( .A(n1048), .B(n1049), .Z(n1047) );
  XNOR U1141 ( .A(n1050), .B(n1005), .Z(n1007) );
  XNOR U1142 ( .A(n1051), .B(n1052), .Z(n1005) );
  AND U1143 ( .A(n1053), .B(n1054), .Z(n1051) );
  AND U1144 ( .A(b[3]), .B(a[30]), .Z(n1050) );
  XOR U1145 ( .A(n1021), .B(n1020), .Z(swire[32]) );
  XOR U1146 ( .A(sreg[96]), .B(n1019), .Z(n1020) );
  XOR U1147 ( .A(n1026), .B(n1055), .Z(n1021) );
  XNOR U1148 ( .A(n1025), .B(n1019), .Z(n1055) );
  XOR U1149 ( .A(n1056), .B(n1057), .Z(n1019) );
  NOR U1150 ( .A(n1058), .B(n1059), .Z(n1056) );
  NANDN U1151 ( .A(n11), .B(a[32]), .Z(n1025) );
  XNOR U1152 ( .A(n1048), .B(n1049), .Z(n1026) );
  XOR U1153 ( .A(n1046), .B(n1060), .Z(n1049) );
  NAND U1154 ( .A(b[1]), .B(a[31]), .Z(n1060) );
  XOR U1155 ( .A(n1054), .B(n1061), .Z(n1048) );
  XOR U1156 ( .A(n1046), .B(n1053), .Z(n1061) );
  XNOR U1157 ( .A(n1062), .B(n1052), .Z(n1053) );
  AND U1158 ( .A(b[2]), .B(a[30]), .Z(n1062) );
  NANDN U1159 ( .A(n1063), .B(n1064), .Z(n1046) );
  XOR U1160 ( .A(n1052), .B(n1044), .Z(n1065) );
  XOR U1161 ( .A(n1043), .B(n1040), .Z(n1066) );
  XOR U1162 ( .A(n1067), .B(n1068), .Z(n1040) );
  XOR U1163 ( .A(n1038), .B(n1069), .Z(n1068) );
  XOR U1164 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U1165 ( .A(n1072), .B(n1073), .Z(n1071) );
  NAND U1166 ( .A(b[6]), .B(a[26]), .Z(n1073) );
  AND U1167 ( .A(b[7]), .B(a[25]), .Z(n1072) );
  XOR U1168 ( .A(n1074), .B(n1070), .Z(n1067) );
  XOR U1169 ( .A(n1075), .B(n1076), .Z(n1070) );
  NOR U1170 ( .A(n1077), .B(n1078), .Z(n1075) );
  AND U1171 ( .A(b[5]), .B(a[27]), .Z(n1074) );
  XNOR U1172 ( .A(n1079), .B(n1038), .Z(n1039) );
  XOR U1173 ( .A(n1080), .B(n1081), .Z(n1038) );
  ANDN U1174 ( .B(n1082), .A(n1083), .Z(n1080) );
  AND U1175 ( .A(b[4]), .B(a[28]), .Z(n1079) );
  XNOR U1176 ( .A(n1084), .B(n1085), .Z(n1052) );
  NANDN U1177 ( .A(n1086), .B(n1087), .Z(n1085) );
  XNOR U1178 ( .A(n1088), .B(n1043), .Z(n1045) );
  XNOR U1179 ( .A(n1089), .B(n1090), .Z(n1043) );
  AND U1180 ( .A(n1091), .B(n1092), .Z(n1089) );
  AND U1181 ( .A(b[3]), .B(a[29]), .Z(n1088) );
  XOR U1182 ( .A(n1059), .B(n1058), .Z(swire[31]) );
  XOR U1183 ( .A(sreg[95]), .B(n1057), .Z(n1058) );
  XOR U1184 ( .A(n1064), .B(n1093), .Z(n1059) );
  XNOR U1185 ( .A(n1063), .B(n1057), .Z(n1093) );
  XOR U1186 ( .A(n1094), .B(n1095), .Z(n1057) );
  NOR U1187 ( .A(n1096), .B(n1097), .Z(n1094) );
  NANDN U1188 ( .A(n11), .B(a[31]), .Z(n1063) );
  XNOR U1189 ( .A(n1086), .B(n1087), .Z(n1064) );
  XOR U1190 ( .A(n1084), .B(n1098), .Z(n1087) );
  NAND U1191 ( .A(b[1]), .B(a[30]), .Z(n1098) );
  XOR U1192 ( .A(n1092), .B(n1099), .Z(n1086) );
  XOR U1193 ( .A(n1084), .B(n1091), .Z(n1099) );
  XNOR U1194 ( .A(n1100), .B(n1090), .Z(n1091) );
  AND U1195 ( .A(b[2]), .B(a[29]), .Z(n1100) );
  NANDN U1196 ( .A(n1101), .B(n1102), .Z(n1084) );
  XOR U1197 ( .A(n1090), .B(n1082), .Z(n1103) );
  XOR U1198 ( .A(n1081), .B(n1078), .Z(n1104) );
  XOR U1199 ( .A(n1105), .B(n1106), .Z(n1078) );
  XOR U1200 ( .A(n1076), .B(n1107), .Z(n1106) );
  XOR U1201 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U1202 ( .A(n1110), .B(n1111), .Z(n1109) );
  NAND U1203 ( .A(b[6]), .B(a[25]), .Z(n1111) );
  AND U1204 ( .A(b[7]), .B(a[24]), .Z(n1110) );
  XOR U1205 ( .A(n1112), .B(n1108), .Z(n1105) );
  XOR U1206 ( .A(n1113), .B(n1114), .Z(n1108) );
  NOR U1207 ( .A(n1115), .B(n1116), .Z(n1113) );
  AND U1208 ( .A(b[5]), .B(a[26]), .Z(n1112) );
  XNOR U1209 ( .A(n1117), .B(n1076), .Z(n1077) );
  XOR U1210 ( .A(n1118), .B(n1119), .Z(n1076) );
  ANDN U1211 ( .B(n1120), .A(n1121), .Z(n1118) );
  AND U1212 ( .A(b[4]), .B(a[27]), .Z(n1117) );
  XNOR U1213 ( .A(n1122), .B(n1123), .Z(n1090) );
  NANDN U1214 ( .A(n1124), .B(n1125), .Z(n1123) );
  XNOR U1215 ( .A(n1126), .B(n1081), .Z(n1083) );
  XNOR U1216 ( .A(n1127), .B(n1128), .Z(n1081) );
  AND U1217 ( .A(n1129), .B(n1130), .Z(n1127) );
  AND U1218 ( .A(b[3]), .B(a[28]), .Z(n1126) );
  XOR U1219 ( .A(n1097), .B(n1096), .Z(swire[30]) );
  XOR U1220 ( .A(sreg[94]), .B(n1095), .Z(n1096) );
  XOR U1221 ( .A(n1102), .B(n1131), .Z(n1097) );
  XNOR U1222 ( .A(n1101), .B(n1095), .Z(n1131) );
  XOR U1223 ( .A(n1132), .B(n1133), .Z(n1095) );
  NOR U1224 ( .A(n1134), .B(n1135), .Z(n1132) );
  NANDN U1225 ( .A(n11), .B(a[30]), .Z(n1101) );
  XNOR U1226 ( .A(n1124), .B(n1125), .Z(n1102) );
  XOR U1227 ( .A(n1122), .B(n1136), .Z(n1125) );
  NAND U1228 ( .A(b[1]), .B(a[29]), .Z(n1136) );
  XOR U1229 ( .A(n1130), .B(n1137), .Z(n1124) );
  XOR U1230 ( .A(n1122), .B(n1129), .Z(n1137) );
  XNOR U1231 ( .A(n1138), .B(n1128), .Z(n1129) );
  AND U1232 ( .A(b[2]), .B(a[28]), .Z(n1138) );
  NANDN U1233 ( .A(n1139), .B(n1140), .Z(n1122) );
  XOR U1234 ( .A(n1128), .B(n1120), .Z(n1141) );
  XOR U1235 ( .A(n1119), .B(n1116), .Z(n1142) );
  XOR U1236 ( .A(n1143), .B(n1144), .Z(n1116) );
  XOR U1237 ( .A(n1114), .B(n1145), .Z(n1144) );
  XOR U1238 ( .A(n1146), .B(n1147), .Z(n1145) );
  XOR U1239 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1240 ( .A(b[6]), .B(a[24]), .Z(n1149) );
  AND U1241 ( .A(b[7]), .B(a[23]), .Z(n1148) );
  XOR U1242 ( .A(n1150), .B(n1146), .Z(n1143) );
  XOR U1243 ( .A(n1151), .B(n1152), .Z(n1146) );
  NOR U1244 ( .A(n1153), .B(n1154), .Z(n1151) );
  AND U1245 ( .A(b[5]), .B(a[25]), .Z(n1150) );
  XNOR U1246 ( .A(n1155), .B(n1114), .Z(n1115) );
  XOR U1247 ( .A(n1156), .B(n1157), .Z(n1114) );
  ANDN U1248 ( .B(n1158), .A(n1159), .Z(n1156) );
  AND U1249 ( .A(b[4]), .B(a[26]), .Z(n1155) );
  XNOR U1250 ( .A(n1160), .B(n1161), .Z(n1128) );
  NANDN U1251 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U1252 ( .A(n1164), .B(n1119), .Z(n1121) );
  XNOR U1253 ( .A(n1165), .B(n1166), .Z(n1119) );
  AND U1254 ( .A(n1167), .B(n1168), .Z(n1165) );
  AND U1255 ( .A(b[3]), .B(a[27]), .Z(n1164) );
  XOR U1256 ( .A(n1135), .B(n1134), .Z(swire[29]) );
  XOR U1257 ( .A(sreg[93]), .B(n1133), .Z(n1134) );
  XOR U1258 ( .A(n1140), .B(n1169), .Z(n1135) );
  XNOR U1259 ( .A(n1139), .B(n1133), .Z(n1169) );
  XOR U1260 ( .A(n1170), .B(n1171), .Z(n1133) );
  NOR U1261 ( .A(n1172), .B(n1173), .Z(n1170) );
  NANDN U1262 ( .A(n11), .B(a[29]), .Z(n1139) );
  XNOR U1263 ( .A(n1162), .B(n1163), .Z(n1140) );
  XOR U1264 ( .A(n1160), .B(n1174), .Z(n1163) );
  NAND U1265 ( .A(b[1]), .B(a[28]), .Z(n1174) );
  XOR U1266 ( .A(n1168), .B(n1175), .Z(n1162) );
  XOR U1267 ( .A(n1160), .B(n1167), .Z(n1175) );
  XNOR U1268 ( .A(n1176), .B(n1166), .Z(n1167) );
  AND U1269 ( .A(b[2]), .B(a[27]), .Z(n1176) );
  NANDN U1270 ( .A(n1177), .B(n1178), .Z(n1160) );
  XOR U1271 ( .A(n1166), .B(n1158), .Z(n1179) );
  XOR U1272 ( .A(n1157), .B(n1154), .Z(n1180) );
  XOR U1273 ( .A(n1181), .B(n1182), .Z(n1154) );
  XOR U1274 ( .A(n1152), .B(n1183), .Z(n1182) );
  XOR U1275 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U1276 ( .A(n1186), .B(n1187), .Z(n1185) );
  NAND U1277 ( .A(b[6]), .B(a[23]), .Z(n1187) );
  AND U1278 ( .A(b[7]), .B(a[22]), .Z(n1186) );
  XOR U1279 ( .A(n1188), .B(n1184), .Z(n1181) );
  XOR U1280 ( .A(n1189), .B(n1190), .Z(n1184) );
  NOR U1281 ( .A(n1191), .B(n1192), .Z(n1189) );
  AND U1282 ( .A(b[5]), .B(a[24]), .Z(n1188) );
  XNOR U1283 ( .A(n1193), .B(n1152), .Z(n1153) );
  XOR U1284 ( .A(n1194), .B(n1195), .Z(n1152) );
  ANDN U1285 ( .B(n1196), .A(n1197), .Z(n1194) );
  AND U1286 ( .A(b[4]), .B(a[25]), .Z(n1193) );
  XNOR U1287 ( .A(n1198), .B(n1199), .Z(n1166) );
  NANDN U1288 ( .A(n1200), .B(n1201), .Z(n1199) );
  XNOR U1289 ( .A(n1202), .B(n1157), .Z(n1159) );
  XNOR U1290 ( .A(n1203), .B(n1204), .Z(n1157) );
  AND U1291 ( .A(n1205), .B(n1206), .Z(n1203) );
  AND U1292 ( .A(b[3]), .B(a[26]), .Z(n1202) );
  XOR U1293 ( .A(n1173), .B(n1172), .Z(swire[28]) );
  XOR U1294 ( .A(sreg[92]), .B(n1171), .Z(n1172) );
  XOR U1295 ( .A(n1178), .B(n1207), .Z(n1173) );
  XNOR U1296 ( .A(n1177), .B(n1171), .Z(n1207) );
  XOR U1297 ( .A(n1208), .B(n1209), .Z(n1171) );
  NOR U1298 ( .A(n1210), .B(n1211), .Z(n1208) );
  NANDN U1299 ( .A(n11), .B(a[28]), .Z(n1177) );
  XNOR U1300 ( .A(n1200), .B(n1201), .Z(n1178) );
  XOR U1301 ( .A(n1198), .B(n1212), .Z(n1201) );
  NAND U1302 ( .A(b[1]), .B(a[27]), .Z(n1212) );
  XOR U1303 ( .A(n1206), .B(n1213), .Z(n1200) );
  XOR U1304 ( .A(n1198), .B(n1205), .Z(n1213) );
  XNOR U1305 ( .A(n1214), .B(n1204), .Z(n1205) );
  AND U1306 ( .A(b[2]), .B(a[26]), .Z(n1214) );
  NANDN U1307 ( .A(n1215), .B(n1216), .Z(n1198) );
  XOR U1308 ( .A(n1204), .B(n1196), .Z(n1217) );
  XOR U1309 ( .A(n1195), .B(n1192), .Z(n1218) );
  XOR U1310 ( .A(n1219), .B(n1220), .Z(n1192) );
  XOR U1311 ( .A(n1190), .B(n1221), .Z(n1220) );
  XOR U1312 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U1313 ( .A(n1224), .B(n1225), .Z(n1223) );
  NAND U1314 ( .A(b[6]), .B(a[22]), .Z(n1225) );
  AND U1315 ( .A(b[7]), .B(a[21]), .Z(n1224) );
  XOR U1316 ( .A(n1226), .B(n1222), .Z(n1219) );
  XOR U1317 ( .A(n1227), .B(n1228), .Z(n1222) );
  NOR U1318 ( .A(n1229), .B(n1230), .Z(n1227) );
  AND U1319 ( .A(b[5]), .B(a[23]), .Z(n1226) );
  XNOR U1320 ( .A(n1231), .B(n1190), .Z(n1191) );
  XOR U1321 ( .A(n1232), .B(n1233), .Z(n1190) );
  ANDN U1322 ( .B(n1234), .A(n1235), .Z(n1232) );
  AND U1323 ( .A(b[4]), .B(a[24]), .Z(n1231) );
  XNOR U1324 ( .A(n1236), .B(n1237), .Z(n1204) );
  NANDN U1325 ( .A(n1238), .B(n1239), .Z(n1237) );
  XNOR U1326 ( .A(n1240), .B(n1195), .Z(n1197) );
  XNOR U1327 ( .A(n1241), .B(n1242), .Z(n1195) );
  AND U1328 ( .A(n1243), .B(n1244), .Z(n1241) );
  AND U1329 ( .A(b[3]), .B(a[25]), .Z(n1240) );
  XOR U1330 ( .A(n1211), .B(n1210), .Z(swire[27]) );
  XOR U1331 ( .A(sreg[91]), .B(n1209), .Z(n1210) );
  XOR U1332 ( .A(n1216), .B(n1245), .Z(n1211) );
  XNOR U1333 ( .A(n1215), .B(n1209), .Z(n1245) );
  XOR U1334 ( .A(n1246), .B(n1247), .Z(n1209) );
  NOR U1335 ( .A(n1248), .B(n1249), .Z(n1246) );
  NANDN U1336 ( .A(n11), .B(a[27]), .Z(n1215) );
  XNOR U1337 ( .A(n1238), .B(n1239), .Z(n1216) );
  XOR U1338 ( .A(n1236), .B(n1250), .Z(n1239) );
  NAND U1339 ( .A(b[1]), .B(a[26]), .Z(n1250) );
  XOR U1340 ( .A(n1244), .B(n1251), .Z(n1238) );
  XOR U1341 ( .A(n1236), .B(n1243), .Z(n1251) );
  XNOR U1342 ( .A(n1252), .B(n1242), .Z(n1243) );
  AND U1343 ( .A(b[2]), .B(a[25]), .Z(n1252) );
  NANDN U1344 ( .A(n1253), .B(n1254), .Z(n1236) );
  XOR U1345 ( .A(n1242), .B(n1234), .Z(n1255) );
  XOR U1346 ( .A(n1233), .B(n1230), .Z(n1256) );
  XOR U1347 ( .A(n1257), .B(n1258), .Z(n1230) );
  XOR U1348 ( .A(n1228), .B(n1259), .Z(n1258) );
  XOR U1349 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U1350 ( .A(n1262), .B(n1263), .Z(n1261) );
  NAND U1351 ( .A(b[6]), .B(a[21]), .Z(n1263) );
  AND U1352 ( .A(b[7]), .B(a[20]), .Z(n1262) );
  XOR U1353 ( .A(n1264), .B(n1260), .Z(n1257) );
  XOR U1354 ( .A(n1265), .B(n1266), .Z(n1260) );
  NOR U1355 ( .A(n1267), .B(n1268), .Z(n1265) );
  AND U1356 ( .A(b[5]), .B(a[22]), .Z(n1264) );
  XNOR U1357 ( .A(n1269), .B(n1228), .Z(n1229) );
  XOR U1358 ( .A(n1270), .B(n1271), .Z(n1228) );
  ANDN U1359 ( .B(n1272), .A(n1273), .Z(n1270) );
  AND U1360 ( .A(b[4]), .B(a[23]), .Z(n1269) );
  XNOR U1361 ( .A(n1274), .B(n1275), .Z(n1242) );
  NANDN U1362 ( .A(n1276), .B(n1277), .Z(n1275) );
  XNOR U1363 ( .A(n1278), .B(n1233), .Z(n1235) );
  XNOR U1364 ( .A(n1279), .B(n1280), .Z(n1233) );
  AND U1365 ( .A(n1281), .B(n1282), .Z(n1279) );
  AND U1366 ( .A(b[3]), .B(a[24]), .Z(n1278) );
  XOR U1367 ( .A(n1249), .B(n1248), .Z(swire[26]) );
  XOR U1368 ( .A(sreg[90]), .B(n1247), .Z(n1248) );
  XOR U1369 ( .A(n1254), .B(n1283), .Z(n1249) );
  XNOR U1370 ( .A(n1253), .B(n1247), .Z(n1283) );
  XOR U1371 ( .A(n1284), .B(n1285), .Z(n1247) );
  NOR U1372 ( .A(n1286), .B(n1287), .Z(n1284) );
  NANDN U1373 ( .A(n11), .B(a[26]), .Z(n1253) );
  XNOR U1374 ( .A(n1276), .B(n1277), .Z(n1254) );
  XOR U1375 ( .A(n1274), .B(n1288), .Z(n1277) );
  NAND U1376 ( .A(b[1]), .B(a[25]), .Z(n1288) );
  XOR U1377 ( .A(n1282), .B(n1289), .Z(n1276) );
  XOR U1378 ( .A(n1274), .B(n1281), .Z(n1289) );
  XNOR U1379 ( .A(n1290), .B(n1280), .Z(n1281) );
  AND U1380 ( .A(b[2]), .B(a[24]), .Z(n1290) );
  NANDN U1381 ( .A(n1291), .B(n1292), .Z(n1274) );
  XOR U1382 ( .A(n1280), .B(n1272), .Z(n1293) );
  XOR U1383 ( .A(n1271), .B(n1268), .Z(n1294) );
  XOR U1384 ( .A(n1295), .B(n1296), .Z(n1268) );
  XOR U1385 ( .A(n1266), .B(n1297), .Z(n1296) );
  XOR U1386 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U1387 ( .A(n1300), .B(n1301), .Z(n1299) );
  NAND U1388 ( .A(b[6]), .B(a[20]), .Z(n1301) );
  AND U1389 ( .A(b[7]), .B(a[19]), .Z(n1300) );
  XOR U1390 ( .A(n1302), .B(n1298), .Z(n1295) );
  XOR U1391 ( .A(n1303), .B(n1304), .Z(n1298) );
  NOR U1392 ( .A(n1305), .B(n1306), .Z(n1303) );
  AND U1393 ( .A(b[5]), .B(a[21]), .Z(n1302) );
  XNOR U1394 ( .A(n1307), .B(n1266), .Z(n1267) );
  XOR U1395 ( .A(n1308), .B(n1309), .Z(n1266) );
  ANDN U1396 ( .B(n1310), .A(n1311), .Z(n1308) );
  AND U1397 ( .A(b[4]), .B(a[22]), .Z(n1307) );
  XNOR U1398 ( .A(n1312), .B(n1313), .Z(n1280) );
  NANDN U1399 ( .A(n1314), .B(n1315), .Z(n1313) );
  XNOR U1400 ( .A(n1316), .B(n1271), .Z(n1273) );
  XNOR U1401 ( .A(n1317), .B(n1318), .Z(n1271) );
  AND U1402 ( .A(n1319), .B(n1320), .Z(n1317) );
  AND U1403 ( .A(b[3]), .B(a[23]), .Z(n1316) );
  XOR U1404 ( .A(n1287), .B(n1286), .Z(swire[25]) );
  XOR U1405 ( .A(sreg[89]), .B(n1285), .Z(n1286) );
  XOR U1406 ( .A(n1292), .B(n1321), .Z(n1287) );
  XNOR U1407 ( .A(n1291), .B(n1285), .Z(n1321) );
  XOR U1408 ( .A(n1322), .B(n1323), .Z(n1285) );
  NOR U1409 ( .A(n1324), .B(n1325), .Z(n1322) );
  NANDN U1410 ( .A(n11), .B(a[25]), .Z(n1291) );
  XNOR U1411 ( .A(n1314), .B(n1315), .Z(n1292) );
  XOR U1412 ( .A(n1312), .B(n1326), .Z(n1315) );
  NAND U1413 ( .A(b[1]), .B(a[24]), .Z(n1326) );
  XOR U1414 ( .A(n1320), .B(n1327), .Z(n1314) );
  XOR U1415 ( .A(n1312), .B(n1319), .Z(n1327) );
  XNOR U1416 ( .A(n1328), .B(n1318), .Z(n1319) );
  AND U1417 ( .A(b[2]), .B(a[23]), .Z(n1328) );
  NANDN U1418 ( .A(n1329), .B(n1330), .Z(n1312) );
  XOR U1419 ( .A(n1318), .B(n1310), .Z(n1331) );
  XOR U1420 ( .A(n1309), .B(n1306), .Z(n1332) );
  XOR U1421 ( .A(n1333), .B(n1334), .Z(n1306) );
  XOR U1422 ( .A(n1304), .B(n1335), .Z(n1334) );
  XOR U1423 ( .A(n1336), .B(n1337), .Z(n1335) );
  XOR U1424 ( .A(n1338), .B(n1339), .Z(n1337) );
  NAND U1425 ( .A(b[6]), .B(a[19]), .Z(n1339) );
  AND U1426 ( .A(b[7]), .B(a[18]), .Z(n1338) );
  XOR U1427 ( .A(n1340), .B(n1336), .Z(n1333) );
  XOR U1428 ( .A(n1341), .B(n1342), .Z(n1336) );
  NOR U1429 ( .A(n1343), .B(n1344), .Z(n1341) );
  AND U1430 ( .A(b[5]), .B(a[20]), .Z(n1340) );
  XNOR U1431 ( .A(n1345), .B(n1304), .Z(n1305) );
  XOR U1432 ( .A(n1346), .B(n1347), .Z(n1304) );
  ANDN U1433 ( .B(n1348), .A(n1349), .Z(n1346) );
  AND U1434 ( .A(b[4]), .B(a[21]), .Z(n1345) );
  XNOR U1435 ( .A(n1350), .B(n1351), .Z(n1318) );
  NANDN U1436 ( .A(n1352), .B(n1353), .Z(n1351) );
  XNOR U1437 ( .A(n1354), .B(n1309), .Z(n1311) );
  XNOR U1438 ( .A(n1355), .B(n1356), .Z(n1309) );
  AND U1439 ( .A(n1357), .B(n1358), .Z(n1355) );
  AND U1440 ( .A(b[3]), .B(a[22]), .Z(n1354) );
  XOR U1441 ( .A(n1325), .B(n1324), .Z(swire[24]) );
  XOR U1442 ( .A(sreg[88]), .B(n1323), .Z(n1324) );
  XOR U1443 ( .A(n1330), .B(n1359), .Z(n1325) );
  XNOR U1444 ( .A(n1329), .B(n1323), .Z(n1359) );
  XOR U1445 ( .A(n1360), .B(n1361), .Z(n1323) );
  NOR U1446 ( .A(n1362), .B(n1363), .Z(n1360) );
  NANDN U1447 ( .A(n11), .B(a[24]), .Z(n1329) );
  XNOR U1448 ( .A(n1352), .B(n1353), .Z(n1330) );
  XOR U1449 ( .A(n1350), .B(n1364), .Z(n1353) );
  NAND U1450 ( .A(b[1]), .B(a[23]), .Z(n1364) );
  XOR U1451 ( .A(n1358), .B(n1365), .Z(n1352) );
  XOR U1452 ( .A(n1350), .B(n1357), .Z(n1365) );
  XNOR U1453 ( .A(n1366), .B(n1356), .Z(n1357) );
  AND U1454 ( .A(b[2]), .B(a[22]), .Z(n1366) );
  NANDN U1455 ( .A(n1367), .B(n1368), .Z(n1350) );
  XOR U1456 ( .A(n1356), .B(n1348), .Z(n1369) );
  XOR U1457 ( .A(n1347), .B(n1344), .Z(n1370) );
  XOR U1458 ( .A(n1371), .B(n1372), .Z(n1344) );
  XOR U1459 ( .A(n1342), .B(n1373), .Z(n1372) );
  XOR U1460 ( .A(n1374), .B(n1375), .Z(n1373) );
  XOR U1461 ( .A(n1376), .B(n1377), .Z(n1375) );
  NAND U1462 ( .A(b[6]), .B(a[18]), .Z(n1377) );
  AND U1463 ( .A(b[7]), .B(a[17]), .Z(n1376) );
  XOR U1464 ( .A(n1378), .B(n1374), .Z(n1371) );
  XOR U1465 ( .A(n1379), .B(n1380), .Z(n1374) );
  NOR U1466 ( .A(n1381), .B(n1382), .Z(n1379) );
  AND U1467 ( .A(b[5]), .B(a[19]), .Z(n1378) );
  XNOR U1468 ( .A(n1383), .B(n1342), .Z(n1343) );
  XOR U1469 ( .A(n1384), .B(n1385), .Z(n1342) );
  ANDN U1470 ( .B(n1386), .A(n1387), .Z(n1384) );
  AND U1471 ( .A(b[4]), .B(a[20]), .Z(n1383) );
  XNOR U1472 ( .A(n1388), .B(n1389), .Z(n1356) );
  NANDN U1473 ( .A(n1390), .B(n1391), .Z(n1389) );
  XNOR U1474 ( .A(n1392), .B(n1347), .Z(n1349) );
  XNOR U1475 ( .A(n1393), .B(n1394), .Z(n1347) );
  AND U1476 ( .A(n1395), .B(n1396), .Z(n1393) );
  AND U1477 ( .A(b[3]), .B(a[21]), .Z(n1392) );
  XOR U1478 ( .A(n1363), .B(n1362), .Z(swire[23]) );
  XOR U1479 ( .A(sreg[87]), .B(n1361), .Z(n1362) );
  XOR U1480 ( .A(n1368), .B(n1397), .Z(n1363) );
  XNOR U1481 ( .A(n1367), .B(n1361), .Z(n1397) );
  XOR U1482 ( .A(n1398), .B(n1399), .Z(n1361) );
  NOR U1483 ( .A(n1400), .B(n1401), .Z(n1398) );
  NANDN U1484 ( .A(n11), .B(a[23]), .Z(n1367) );
  XNOR U1485 ( .A(n1390), .B(n1391), .Z(n1368) );
  XOR U1486 ( .A(n1388), .B(n1402), .Z(n1391) );
  NAND U1487 ( .A(b[1]), .B(a[22]), .Z(n1402) );
  XOR U1488 ( .A(n1396), .B(n1403), .Z(n1390) );
  XOR U1489 ( .A(n1388), .B(n1395), .Z(n1403) );
  XNOR U1490 ( .A(n1404), .B(n1394), .Z(n1395) );
  AND U1491 ( .A(b[2]), .B(a[21]), .Z(n1404) );
  NANDN U1492 ( .A(n1405), .B(n1406), .Z(n1388) );
  XOR U1493 ( .A(n1394), .B(n1386), .Z(n1407) );
  XOR U1494 ( .A(n1385), .B(n1382), .Z(n1408) );
  XOR U1495 ( .A(n1409), .B(n1410), .Z(n1382) );
  XOR U1496 ( .A(n1380), .B(n1411), .Z(n1410) );
  XOR U1497 ( .A(n1412), .B(n1413), .Z(n1411) );
  XOR U1498 ( .A(n1414), .B(n1415), .Z(n1413) );
  NAND U1499 ( .A(b[6]), .B(a[17]), .Z(n1415) );
  AND U1500 ( .A(b[7]), .B(a[16]), .Z(n1414) );
  XOR U1501 ( .A(n1416), .B(n1412), .Z(n1409) );
  XOR U1502 ( .A(n1417), .B(n1418), .Z(n1412) );
  NOR U1503 ( .A(n1419), .B(n1420), .Z(n1417) );
  AND U1504 ( .A(b[5]), .B(a[18]), .Z(n1416) );
  XNOR U1505 ( .A(n1421), .B(n1380), .Z(n1381) );
  XOR U1506 ( .A(n1422), .B(n1423), .Z(n1380) );
  ANDN U1507 ( .B(n1424), .A(n1425), .Z(n1422) );
  AND U1508 ( .A(b[4]), .B(a[19]), .Z(n1421) );
  XNOR U1509 ( .A(n1426), .B(n1427), .Z(n1394) );
  NANDN U1510 ( .A(n1428), .B(n1429), .Z(n1427) );
  XNOR U1511 ( .A(n1430), .B(n1385), .Z(n1387) );
  XNOR U1512 ( .A(n1431), .B(n1432), .Z(n1385) );
  AND U1513 ( .A(n1433), .B(n1434), .Z(n1431) );
  AND U1514 ( .A(b[3]), .B(a[20]), .Z(n1430) );
  XOR U1515 ( .A(n1401), .B(n1400), .Z(swire[22]) );
  XOR U1516 ( .A(sreg[86]), .B(n1399), .Z(n1400) );
  XOR U1517 ( .A(n1406), .B(n1435), .Z(n1401) );
  XNOR U1518 ( .A(n1405), .B(n1399), .Z(n1435) );
  XOR U1519 ( .A(n1436), .B(n1437), .Z(n1399) );
  NOR U1520 ( .A(n1438), .B(n1439), .Z(n1436) );
  NANDN U1521 ( .A(n11), .B(a[22]), .Z(n1405) );
  XNOR U1522 ( .A(n1428), .B(n1429), .Z(n1406) );
  XOR U1523 ( .A(n1426), .B(n1440), .Z(n1429) );
  NAND U1524 ( .A(b[1]), .B(a[21]), .Z(n1440) );
  XOR U1525 ( .A(n1434), .B(n1441), .Z(n1428) );
  XOR U1526 ( .A(n1426), .B(n1433), .Z(n1441) );
  XNOR U1527 ( .A(n1442), .B(n1432), .Z(n1433) );
  AND U1528 ( .A(b[2]), .B(a[20]), .Z(n1442) );
  NANDN U1529 ( .A(n1443), .B(n1444), .Z(n1426) );
  XOR U1530 ( .A(n1432), .B(n1424), .Z(n1445) );
  XOR U1531 ( .A(n1423), .B(n1420), .Z(n1446) );
  XOR U1532 ( .A(n1447), .B(n1448), .Z(n1420) );
  XOR U1533 ( .A(n1418), .B(n1449), .Z(n1448) );
  XOR U1534 ( .A(n1450), .B(n1451), .Z(n1449) );
  XOR U1535 ( .A(n1452), .B(n1453), .Z(n1451) );
  NAND U1536 ( .A(b[6]), .B(a[16]), .Z(n1453) );
  AND U1537 ( .A(b[7]), .B(a[15]), .Z(n1452) );
  XOR U1538 ( .A(n1454), .B(n1450), .Z(n1447) );
  XOR U1539 ( .A(n1455), .B(n1456), .Z(n1450) );
  NOR U1540 ( .A(n1457), .B(n1458), .Z(n1455) );
  AND U1541 ( .A(b[5]), .B(a[17]), .Z(n1454) );
  XNOR U1542 ( .A(n1459), .B(n1418), .Z(n1419) );
  XOR U1543 ( .A(n1460), .B(n1461), .Z(n1418) );
  ANDN U1544 ( .B(n1462), .A(n1463), .Z(n1460) );
  AND U1545 ( .A(b[4]), .B(a[18]), .Z(n1459) );
  XNOR U1546 ( .A(n1464), .B(n1465), .Z(n1432) );
  NANDN U1547 ( .A(n1466), .B(n1467), .Z(n1465) );
  XNOR U1548 ( .A(n1468), .B(n1423), .Z(n1425) );
  XNOR U1549 ( .A(n1469), .B(n1470), .Z(n1423) );
  AND U1550 ( .A(n1471), .B(n1472), .Z(n1469) );
  AND U1551 ( .A(b[3]), .B(a[19]), .Z(n1468) );
  XOR U1552 ( .A(n1439), .B(n1438), .Z(swire[21]) );
  XOR U1553 ( .A(sreg[85]), .B(n1437), .Z(n1438) );
  XOR U1554 ( .A(n1444), .B(n1473), .Z(n1439) );
  XNOR U1555 ( .A(n1443), .B(n1437), .Z(n1473) );
  XOR U1556 ( .A(n1474), .B(n1475), .Z(n1437) );
  NOR U1557 ( .A(n1476), .B(n1477), .Z(n1474) );
  NANDN U1558 ( .A(n11), .B(a[21]), .Z(n1443) );
  XNOR U1559 ( .A(n1466), .B(n1467), .Z(n1444) );
  XOR U1560 ( .A(n1464), .B(n1478), .Z(n1467) );
  NAND U1561 ( .A(b[1]), .B(a[20]), .Z(n1478) );
  XOR U1562 ( .A(n1472), .B(n1479), .Z(n1466) );
  XOR U1563 ( .A(n1464), .B(n1471), .Z(n1479) );
  XNOR U1564 ( .A(n1480), .B(n1470), .Z(n1471) );
  AND U1565 ( .A(b[2]), .B(a[19]), .Z(n1480) );
  NANDN U1566 ( .A(n1481), .B(n1482), .Z(n1464) );
  XOR U1567 ( .A(n1470), .B(n1462), .Z(n1483) );
  XOR U1568 ( .A(n1461), .B(n1458), .Z(n1484) );
  XOR U1569 ( .A(n1485), .B(n1486), .Z(n1458) );
  XOR U1570 ( .A(n1456), .B(n1487), .Z(n1486) );
  XOR U1571 ( .A(n1488), .B(n1489), .Z(n1487) );
  XOR U1572 ( .A(n1490), .B(n1491), .Z(n1489) );
  NAND U1573 ( .A(b[6]), .B(a[15]), .Z(n1491) );
  AND U1574 ( .A(b[7]), .B(a[14]), .Z(n1490) );
  XOR U1575 ( .A(n1492), .B(n1488), .Z(n1485) );
  XOR U1576 ( .A(n1493), .B(n1494), .Z(n1488) );
  NOR U1577 ( .A(n1495), .B(n1496), .Z(n1493) );
  AND U1578 ( .A(b[5]), .B(a[16]), .Z(n1492) );
  XNOR U1579 ( .A(n1497), .B(n1456), .Z(n1457) );
  XOR U1580 ( .A(n1498), .B(n1499), .Z(n1456) );
  ANDN U1581 ( .B(n1500), .A(n1501), .Z(n1498) );
  AND U1582 ( .A(b[4]), .B(a[17]), .Z(n1497) );
  XNOR U1583 ( .A(n1502), .B(n1503), .Z(n1470) );
  NANDN U1584 ( .A(n1504), .B(n1505), .Z(n1503) );
  XNOR U1585 ( .A(n1506), .B(n1461), .Z(n1463) );
  XNOR U1586 ( .A(n1507), .B(n1508), .Z(n1461) );
  AND U1587 ( .A(n1509), .B(n1510), .Z(n1507) );
  AND U1588 ( .A(b[3]), .B(a[18]), .Z(n1506) );
  XOR U1589 ( .A(n1477), .B(n1476), .Z(swire[20]) );
  XOR U1590 ( .A(sreg[84]), .B(n1475), .Z(n1476) );
  XOR U1591 ( .A(n1482), .B(n1511), .Z(n1477) );
  XNOR U1592 ( .A(n1481), .B(n1475), .Z(n1511) );
  XOR U1593 ( .A(n1512), .B(n1513), .Z(n1475) );
  NOR U1594 ( .A(n1514), .B(n1515), .Z(n1512) );
  NANDN U1595 ( .A(n11), .B(a[20]), .Z(n1481) );
  XNOR U1596 ( .A(n1504), .B(n1505), .Z(n1482) );
  XOR U1597 ( .A(n1502), .B(n1516), .Z(n1505) );
  NAND U1598 ( .A(b[1]), .B(a[19]), .Z(n1516) );
  XOR U1599 ( .A(n1510), .B(n1517), .Z(n1504) );
  XOR U1600 ( .A(n1502), .B(n1509), .Z(n1517) );
  XNOR U1601 ( .A(n1518), .B(n1508), .Z(n1509) );
  AND U1602 ( .A(b[2]), .B(a[18]), .Z(n1518) );
  NANDN U1603 ( .A(n1519), .B(n1520), .Z(n1502) );
  XOR U1604 ( .A(n1508), .B(n1500), .Z(n1521) );
  XOR U1605 ( .A(n1499), .B(n1496), .Z(n1522) );
  XOR U1606 ( .A(n1523), .B(n1524), .Z(n1496) );
  XOR U1607 ( .A(n1494), .B(n1525), .Z(n1524) );
  XOR U1608 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U1609 ( .A(n1528), .B(n1529), .Z(n1527) );
  NAND U1610 ( .A(b[6]), .B(a[14]), .Z(n1529) );
  AND U1611 ( .A(b[7]), .B(a[13]), .Z(n1528) );
  XOR U1612 ( .A(n1530), .B(n1526), .Z(n1523) );
  XOR U1613 ( .A(n1531), .B(n1532), .Z(n1526) );
  NOR U1614 ( .A(n1533), .B(n1534), .Z(n1531) );
  AND U1615 ( .A(b[5]), .B(a[15]), .Z(n1530) );
  XNOR U1616 ( .A(n1535), .B(n1494), .Z(n1495) );
  XOR U1617 ( .A(n1536), .B(n1537), .Z(n1494) );
  ANDN U1618 ( .B(n1538), .A(n1539), .Z(n1536) );
  AND U1619 ( .A(b[4]), .B(a[16]), .Z(n1535) );
  XNOR U1620 ( .A(n1540), .B(n1541), .Z(n1508) );
  NANDN U1621 ( .A(n1542), .B(n1543), .Z(n1541) );
  XNOR U1622 ( .A(n1544), .B(n1499), .Z(n1501) );
  XNOR U1623 ( .A(n1545), .B(n1546), .Z(n1499) );
  AND U1624 ( .A(n1547), .B(n1548), .Z(n1545) );
  AND U1625 ( .A(b[3]), .B(a[17]), .Z(n1544) );
  XOR U1626 ( .A(n1515), .B(n1514), .Z(swire[19]) );
  XOR U1627 ( .A(sreg[83]), .B(n1513), .Z(n1514) );
  XOR U1628 ( .A(n1520), .B(n1549), .Z(n1515) );
  XNOR U1629 ( .A(n1519), .B(n1513), .Z(n1549) );
  XOR U1630 ( .A(n1550), .B(n1551), .Z(n1513) );
  NOR U1631 ( .A(n1552), .B(n1553), .Z(n1550) );
  NANDN U1632 ( .A(n11), .B(a[19]), .Z(n1519) );
  XNOR U1633 ( .A(n1542), .B(n1543), .Z(n1520) );
  XOR U1634 ( .A(n1540), .B(n1554), .Z(n1543) );
  NAND U1635 ( .A(b[1]), .B(a[18]), .Z(n1554) );
  XOR U1636 ( .A(n1548), .B(n1555), .Z(n1542) );
  XOR U1637 ( .A(n1540), .B(n1547), .Z(n1555) );
  XNOR U1638 ( .A(n1556), .B(n1546), .Z(n1547) );
  AND U1639 ( .A(b[2]), .B(a[17]), .Z(n1556) );
  NANDN U1640 ( .A(n1557), .B(n1558), .Z(n1540) );
  XOR U1641 ( .A(n1546), .B(n1538), .Z(n1559) );
  XOR U1642 ( .A(n1537), .B(n1534), .Z(n1560) );
  XOR U1643 ( .A(n1561), .B(n1562), .Z(n1534) );
  XOR U1644 ( .A(n1532), .B(n1563), .Z(n1562) );
  XOR U1645 ( .A(n1564), .B(n1565), .Z(n1563) );
  XOR U1646 ( .A(n1566), .B(n1567), .Z(n1565) );
  NAND U1647 ( .A(b[6]), .B(a[13]), .Z(n1567) );
  AND U1648 ( .A(b[7]), .B(a[12]), .Z(n1566) );
  XOR U1649 ( .A(n1568), .B(n1564), .Z(n1561) );
  XOR U1650 ( .A(n1569), .B(n1570), .Z(n1564) );
  NOR U1651 ( .A(n1571), .B(n1572), .Z(n1569) );
  AND U1652 ( .A(b[5]), .B(a[14]), .Z(n1568) );
  XNOR U1653 ( .A(n1573), .B(n1532), .Z(n1533) );
  XOR U1654 ( .A(n1574), .B(n1575), .Z(n1532) );
  ANDN U1655 ( .B(n1576), .A(n1577), .Z(n1574) );
  AND U1656 ( .A(b[4]), .B(a[15]), .Z(n1573) );
  XNOR U1657 ( .A(n1578), .B(n1579), .Z(n1546) );
  NANDN U1658 ( .A(n1580), .B(n1581), .Z(n1579) );
  XNOR U1659 ( .A(n1582), .B(n1537), .Z(n1539) );
  XNOR U1660 ( .A(n1583), .B(n1584), .Z(n1537) );
  AND U1661 ( .A(n1585), .B(n1586), .Z(n1583) );
  AND U1662 ( .A(b[3]), .B(a[16]), .Z(n1582) );
  XOR U1663 ( .A(n1553), .B(n1552), .Z(swire[18]) );
  XOR U1664 ( .A(sreg[82]), .B(n1551), .Z(n1552) );
  XOR U1665 ( .A(n1558), .B(n1587), .Z(n1553) );
  XNOR U1666 ( .A(n1557), .B(n1551), .Z(n1587) );
  XOR U1667 ( .A(n1588), .B(n1589), .Z(n1551) );
  NOR U1668 ( .A(n1590), .B(n1591), .Z(n1588) );
  NANDN U1669 ( .A(n11), .B(a[18]), .Z(n1557) );
  XNOR U1670 ( .A(n1580), .B(n1581), .Z(n1558) );
  XOR U1671 ( .A(n1578), .B(n1592), .Z(n1581) );
  NAND U1672 ( .A(b[1]), .B(a[17]), .Z(n1592) );
  XOR U1673 ( .A(n1586), .B(n1593), .Z(n1580) );
  XOR U1674 ( .A(n1578), .B(n1585), .Z(n1593) );
  XNOR U1675 ( .A(n1594), .B(n1584), .Z(n1585) );
  AND U1676 ( .A(b[2]), .B(a[16]), .Z(n1594) );
  NANDN U1677 ( .A(n1595), .B(n1596), .Z(n1578) );
  XOR U1678 ( .A(n1584), .B(n1576), .Z(n1597) );
  XOR U1679 ( .A(n1575), .B(n1572), .Z(n1598) );
  XOR U1680 ( .A(n1599), .B(n1600), .Z(n1572) );
  XOR U1681 ( .A(n1570), .B(n1601), .Z(n1600) );
  XOR U1682 ( .A(n1602), .B(n1603), .Z(n1601) );
  XOR U1683 ( .A(n1604), .B(n1605), .Z(n1603) );
  NAND U1684 ( .A(b[6]), .B(a[12]), .Z(n1605) );
  AND U1685 ( .A(b[7]), .B(a[11]), .Z(n1604) );
  XOR U1686 ( .A(n1606), .B(n1602), .Z(n1599) );
  XOR U1687 ( .A(n1607), .B(n1608), .Z(n1602) );
  NOR U1688 ( .A(n1609), .B(n1610), .Z(n1607) );
  AND U1689 ( .A(b[5]), .B(a[13]), .Z(n1606) );
  XNOR U1690 ( .A(n1611), .B(n1570), .Z(n1571) );
  XOR U1691 ( .A(n1612), .B(n1613), .Z(n1570) );
  ANDN U1692 ( .B(n1614), .A(n1615), .Z(n1612) );
  AND U1693 ( .A(b[4]), .B(a[14]), .Z(n1611) );
  XNOR U1694 ( .A(n1616), .B(n1617), .Z(n1584) );
  NANDN U1695 ( .A(n1618), .B(n1619), .Z(n1617) );
  XNOR U1696 ( .A(n1620), .B(n1575), .Z(n1577) );
  XNOR U1697 ( .A(n1621), .B(n1622), .Z(n1575) );
  AND U1698 ( .A(n1623), .B(n1624), .Z(n1621) );
  AND U1699 ( .A(b[3]), .B(a[15]), .Z(n1620) );
  XOR U1700 ( .A(n1591), .B(n1590), .Z(swire[17]) );
  XOR U1701 ( .A(sreg[81]), .B(n1589), .Z(n1590) );
  XOR U1702 ( .A(n1596), .B(n1625), .Z(n1591) );
  XNOR U1703 ( .A(n1595), .B(n1589), .Z(n1625) );
  XOR U1704 ( .A(n1626), .B(n1627), .Z(n1589) );
  NOR U1705 ( .A(n1628), .B(n1629), .Z(n1626) );
  NANDN U1706 ( .A(n11), .B(a[17]), .Z(n1595) );
  XNOR U1707 ( .A(n1618), .B(n1619), .Z(n1596) );
  XOR U1708 ( .A(n1616), .B(n1630), .Z(n1619) );
  NAND U1709 ( .A(b[1]), .B(a[16]), .Z(n1630) );
  XOR U1710 ( .A(n1624), .B(n1631), .Z(n1618) );
  XOR U1711 ( .A(n1616), .B(n1623), .Z(n1631) );
  XNOR U1712 ( .A(n1632), .B(n1622), .Z(n1623) );
  AND U1713 ( .A(b[2]), .B(a[15]), .Z(n1632) );
  NANDN U1714 ( .A(n1633), .B(n1634), .Z(n1616) );
  XOR U1715 ( .A(n1622), .B(n1614), .Z(n1635) );
  XOR U1716 ( .A(n1613), .B(n1610), .Z(n1636) );
  XOR U1717 ( .A(n1637), .B(n1638), .Z(n1610) );
  XOR U1718 ( .A(n1608), .B(n1639), .Z(n1638) );
  XOR U1719 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U1720 ( .A(n1642), .B(n1643), .Z(n1641) );
  NAND U1721 ( .A(b[6]), .B(a[11]), .Z(n1643) );
  AND U1722 ( .A(b[7]), .B(a[10]), .Z(n1642) );
  XOR U1723 ( .A(n1644), .B(n1640), .Z(n1637) );
  XOR U1724 ( .A(n1645), .B(n1646), .Z(n1640) );
  NOR U1725 ( .A(n1647), .B(n1648), .Z(n1645) );
  AND U1726 ( .A(b[5]), .B(a[12]), .Z(n1644) );
  XNOR U1727 ( .A(n1649), .B(n1608), .Z(n1609) );
  XOR U1728 ( .A(n1650), .B(n1651), .Z(n1608) );
  ANDN U1729 ( .B(n1652), .A(n1653), .Z(n1650) );
  AND U1730 ( .A(b[4]), .B(a[13]), .Z(n1649) );
  XNOR U1731 ( .A(n1654), .B(n1655), .Z(n1622) );
  NANDN U1732 ( .A(n1656), .B(n1657), .Z(n1655) );
  XNOR U1733 ( .A(n1658), .B(n1613), .Z(n1615) );
  XNOR U1734 ( .A(n1659), .B(n1660), .Z(n1613) );
  AND U1735 ( .A(n1661), .B(n1662), .Z(n1659) );
  AND U1736 ( .A(b[3]), .B(a[14]), .Z(n1658) );
  XOR U1737 ( .A(n1629), .B(n1628), .Z(swire[16]) );
  XOR U1738 ( .A(sreg[80]), .B(n1627), .Z(n1628) );
  XOR U1739 ( .A(n1634), .B(n1663), .Z(n1629) );
  XNOR U1740 ( .A(n1633), .B(n1627), .Z(n1663) );
  XOR U1741 ( .A(n1664), .B(n1665), .Z(n1627) );
  NOR U1742 ( .A(n1666), .B(n1667), .Z(n1664) );
  NANDN U1743 ( .A(n11), .B(a[16]), .Z(n1633) );
  XNOR U1744 ( .A(n1656), .B(n1657), .Z(n1634) );
  XOR U1745 ( .A(n1654), .B(n1668), .Z(n1657) );
  NAND U1746 ( .A(b[1]), .B(a[15]), .Z(n1668) );
  XOR U1747 ( .A(n1662), .B(n1669), .Z(n1656) );
  XOR U1748 ( .A(n1654), .B(n1661), .Z(n1669) );
  XNOR U1749 ( .A(n1670), .B(n1660), .Z(n1661) );
  AND U1750 ( .A(b[2]), .B(a[14]), .Z(n1670) );
  NANDN U1751 ( .A(n1671), .B(n1672), .Z(n1654) );
  XOR U1752 ( .A(n1660), .B(n1652), .Z(n1673) );
  XOR U1753 ( .A(n1651), .B(n1648), .Z(n1674) );
  XOR U1754 ( .A(n1675), .B(n1676), .Z(n1648) );
  XOR U1755 ( .A(n1646), .B(n1677), .Z(n1676) );
  XOR U1756 ( .A(n1678), .B(n1679), .Z(n1677) );
  XOR U1757 ( .A(n1680), .B(n1681), .Z(n1679) );
  NAND U1758 ( .A(b[6]), .B(a[10]), .Z(n1681) );
  AND U1759 ( .A(b[7]), .B(a[9]), .Z(n1680) );
  XOR U1760 ( .A(n1682), .B(n1678), .Z(n1675) );
  XOR U1761 ( .A(n1683), .B(n1684), .Z(n1678) );
  NOR U1762 ( .A(n1685), .B(n1686), .Z(n1683) );
  AND U1763 ( .A(b[5]), .B(a[11]), .Z(n1682) );
  XNOR U1764 ( .A(n1687), .B(n1646), .Z(n1647) );
  XOR U1765 ( .A(n1688), .B(n1689), .Z(n1646) );
  ANDN U1766 ( .B(n1690), .A(n1691), .Z(n1688) );
  AND U1767 ( .A(b[4]), .B(a[12]), .Z(n1687) );
  XNOR U1768 ( .A(n1692), .B(n1693), .Z(n1660) );
  NANDN U1769 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U1770 ( .A(n1696), .B(n1651), .Z(n1653) );
  XNOR U1771 ( .A(n1697), .B(n1698), .Z(n1651) );
  AND U1772 ( .A(n1699), .B(n1700), .Z(n1697) );
  AND U1773 ( .A(b[3]), .B(a[13]), .Z(n1696) );
  XOR U1774 ( .A(n1667), .B(n1666), .Z(swire[15]) );
  XOR U1775 ( .A(sreg[79]), .B(n1665), .Z(n1666) );
  XOR U1776 ( .A(n1672), .B(n1701), .Z(n1667) );
  XNOR U1777 ( .A(n1671), .B(n1665), .Z(n1701) );
  XOR U1778 ( .A(n1702), .B(n1703), .Z(n1665) );
  NOR U1779 ( .A(n1704), .B(n1705), .Z(n1702) );
  NANDN U1780 ( .A(n11), .B(a[15]), .Z(n1671) );
  XNOR U1781 ( .A(n1694), .B(n1695), .Z(n1672) );
  XOR U1782 ( .A(n1692), .B(n1706), .Z(n1695) );
  NAND U1783 ( .A(b[1]), .B(a[14]), .Z(n1706) );
  XOR U1784 ( .A(n1700), .B(n1707), .Z(n1694) );
  XOR U1785 ( .A(n1692), .B(n1699), .Z(n1707) );
  XNOR U1786 ( .A(n1708), .B(n1698), .Z(n1699) );
  AND U1787 ( .A(b[2]), .B(a[13]), .Z(n1708) );
  NANDN U1788 ( .A(n1709), .B(n1710), .Z(n1692) );
  XOR U1789 ( .A(n1698), .B(n1690), .Z(n1711) );
  XOR U1790 ( .A(n1689), .B(n1686), .Z(n1712) );
  XOR U1791 ( .A(n1713), .B(n1714), .Z(n1686) );
  XOR U1792 ( .A(n1684), .B(n1715), .Z(n1714) );
  XOR U1793 ( .A(n1716), .B(n1717), .Z(n1715) );
  XOR U1794 ( .A(n1718), .B(n1719), .Z(n1717) );
  NAND U1795 ( .A(b[6]), .B(a[9]), .Z(n1719) );
  AND U1796 ( .A(b[7]), .B(a[8]), .Z(n1718) );
  XOR U1797 ( .A(n1720), .B(n1716), .Z(n1713) );
  XOR U1798 ( .A(n1721), .B(n1722), .Z(n1716) );
  NOR U1799 ( .A(n1723), .B(n1724), .Z(n1721) );
  AND U1800 ( .A(b[5]), .B(a[10]), .Z(n1720) );
  XNOR U1801 ( .A(n1725), .B(n1684), .Z(n1685) );
  XOR U1802 ( .A(n1726), .B(n1727), .Z(n1684) );
  ANDN U1803 ( .B(n1728), .A(n1729), .Z(n1726) );
  AND U1804 ( .A(b[4]), .B(a[11]), .Z(n1725) );
  XNOR U1805 ( .A(n1730), .B(n1731), .Z(n1698) );
  NANDN U1806 ( .A(n1732), .B(n1733), .Z(n1731) );
  XNOR U1807 ( .A(n1734), .B(n1689), .Z(n1691) );
  XNOR U1808 ( .A(n1735), .B(n1736), .Z(n1689) );
  AND U1809 ( .A(n1737), .B(n1738), .Z(n1735) );
  AND U1810 ( .A(b[3]), .B(a[12]), .Z(n1734) );
  XOR U1811 ( .A(n1705), .B(n1704), .Z(swire[14]) );
  XOR U1812 ( .A(sreg[78]), .B(n1703), .Z(n1704) );
  XOR U1813 ( .A(n1710), .B(n1739), .Z(n1705) );
  XNOR U1814 ( .A(n1709), .B(n1703), .Z(n1739) );
  XOR U1815 ( .A(n1740), .B(n1741), .Z(n1703) );
  NOR U1816 ( .A(n1742), .B(n1743), .Z(n1740) );
  NANDN U1817 ( .A(n11), .B(a[14]), .Z(n1709) );
  XNOR U1818 ( .A(n1732), .B(n1733), .Z(n1710) );
  XOR U1819 ( .A(n1730), .B(n1744), .Z(n1733) );
  NAND U1820 ( .A(b[1]), .B(a[13]), .Z(n1744) );
  XOR U1821 ( .A(n1738), .B(n1745), .Z(n1732) );
  XOR U1822 ( .A(n1730), .B(n1737), .Z(n1745) );
  XNOR U1823 ( .A(n1746), .B(n1736), .Z(n1737) );
  AND U1824 ( .A(b[2]), .B(a[12]), .Z(n1746) );
  NANDN U1825 ( .A(n1747), .B(n1748), .Z(n1730) );
  XOR U1826 ( .A(n1736), .B(n1728), .Z(n1749) );
  XOR U1827 ( .A(n1727), .B(n1724), .Z(n1750) );
  XOR U1828 ( .A(n1751), .B(n1752), .Z(n1724) );
  XOR U1829 ( .A(n1722), .B(n1753), .Z(n1752) );
  XOR U1830 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U1831 ( .A(n1756), .B(n1757), .Z(n1755) );
  NAND U1832 ( .A(b[6]), .B(a[8]), .Z(n1757) );
  AND U1833 ( .A(a[7]), .B(b[7]), .Z(n1756) );
  XOR U1834 ( .A(n1758), .B(n1754), .Z(n1751) );
  XOR U1835 ( .A(n1759), .B(n1760), .Z(n1754) );
  NOR U1836 ( .A(n1761), .B(n1762), .Z(n1759) );
  AND U1837 ( .A(b[5]), .B(a[9]), .Z(n1758) );
  XNOR U1838 ( .A(n1763), .B(n1722), .Z(n1723) );
  XOR U1839 ( .A(n1764), .B(n1765), .Z(n1722) );
  ANDN U1840 ( .B(n1766), .A(n1767), .Z(n1764) );
  AND U1841 ( .A(b[4]), .B(a[10]), .Z(n1763) );
  XNOR U1842 ( .A(n1768), .B(n1769), .Z(n1736) );
  NANDN U1843 ( .A(n1770), .B(n1771), .Z(n1769) );
  XNOR U1844 ( .A(n1772), .B(n1727), .Z(n1729) );
  XNOR U1845 ( .A(n1773), .B(n1774), .Z(n1727) );
  AND U1846 ( .A(n1775), .B(n1776), .Z(n1773) );
  AND U1847 ( .A(b[3]), .B(a[11]), .Z(n1772) );
  XOR U1848 ( .A(n1743), .B(n1742), .Z(swire[13]) );
  XOR U1849 ( .A(sreg[77]), .B(n1741), .Z(n1742) );
  XOR U1850 ( .A(n1748), .B(n1777), .Z(n1743) );
  XNOR U1851 ( .A(n1747), .B(n1741), .Z(n1777) );
  XOR U1852 ( .A(n1778), .B(n1779), .Z(n1741) );
  NOR U1853 ( .A(n1780), .B(n1781), .Z(n1778) );
  NANDN U1854 ( .A(n11), .B(a[13]), .Z(n1747) );
  XNOR U1855 ( .A(n1770), .B(n1771), .Z(n1748) );
  XOR U1856 ( .A(n1768), .B(n1782), .Z(n1771) );
  NAND U1857 ( .A(b[1]), .B(a[12]), .Z(n1782) );
  XOR U1858 ( .A(n1776), .B(n1783), .Z(n1770) );
  XOR U1859 ( .A(n1768), .B(n1775), .Z(n1783) );
  XNOR U1860 ( .A(n1784), .B(n1774), .Z(n1775) );
  AND U1861 ( .A(b[2]), .B(a[11]), .Z(n1784) );
  NANDN U1862 ( .A(n1785), .B(n1786), .Z(n1768) );
  XOR U1863 ( .A(n1774), .B(n1766), .Z(n1787) );
  XOR U1864 ( .A(n1765), .B(n1762), .Z(n1788) );
  XOR U1865 ( .A(n1789), .B(n1790), .Z(n1762) );
  XOR U1866 ( .A(n1760), .B(n1791), .Z(n1790) );
  XOR U1867 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U1868 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1869 ( .A(a[7]), .B(b[6]), .Z(n1795) );
  AND U1870 ( .A(a[6]), .B(b[7]), .Z(n1794) );
  XOR U1871 ( .A(n1796), .B(n1792), .Z(n1789) );
  XOR U1872 ( .A(n1797), .B(n1798), .Z(n1792) );
  NOR U1873 ( .A(n1799), .B(n1800), .Z(n1797) );
  AND U1874 ( .A(b[5]), .B(a[8]), .Z(n1796) );
  XNOR U1875 ( .A(n1801), .B(n1760), .Z(n1761) );
  XOR U1876 ( .A(n1802), .B(n1803), .Z(n1760) );
  ANDN U1877 ( .B(n1804), .A(n1805), .Z(n1802) );
  AND U1878 ( .A(b[4]), .B(a[9]), .Z(n1801) );
  XNOR U1879 ( .A(n1806), .B(n1807), .Z(n1774) );
  NANDN U1880 ( .A(n1808), .B(n1809), .Z(n1807) );
  XNOR U1881 ( .A(n1810), .B(n1765), .Z(n1767) );
  XNOR U1882 ( .A(n1811), .B(n1812), .Z(n1765) );
  AND U1883 ( .A(n1813), .B(n1814), .Z(n1811) );
  AND U1884 ( .A(b[3]), .B(a[10]), .Z(n1810) );
  XOR U1885 ( .A(n1781), .B(n1780), .Z(swire[12]) );
  XOR U1886 ( .A(sreg[76]), .B(n1779), .Z(n1780) );
  XOR U1887 ( .A(n1786), .B(n1815), .Z(n1781) );
  XNOR U1888 ( .A(n1785), .B(n1779), .Z(n1815) );
  XOR U1889 ( .A(n1816), .B(n1817), .Z(n1779) );
  NOR U1890 ( .A(n1818), .B(n1819), .Z(n1816) );
  NANDN U1891 ( .A(n11), .B(a[12]), .Z(n1785) );
  XNOR U1892 ( .A(n1808), .B(n1809), .Z(n1786) );
  XOR U1893 ( .A(n1806), .B(n1820), .Z(n1809) );
  NAND U1894 ( .A(b[1]), .B(a[11]), .Z(n1820) );
  XOR U1895 ( .A(n1814), .B(n1821), .Z(n1808) );
  XOR U1896 ( .A(n1806), .B(n1813), .Z(n1821) );
  XNOR U1897 ( .A(n1822), .B(n1812), .Z(n1813) );
  AND U1898 ( .A(b[2]), .B(a[10]), .Z(n1822) );
  NANDN U1899 ( .A(n1823), .B(n1824), .Z(n1806) );
  XOR U1900 ( .A(n1812), .B(n1804), .Z(n1825) );
  XOR U1901 ( .A(n1803), .B(n1800), .Z(n1826) );
  XOR U1902 ( .A(n1827), .B(n1828), .Z(n1800) );
  XOR U1903 ( .A(n1798), .B(n1829), .Z(n1828) );
  XOR U1904 ( .A(n1830), .B(n1831), .Z(n1829) );
  XOR U1905 ( .A(n1832), .B(n1833), .Z(n1831) );
  NAND U1906 ( .A(b[6]), .B(a[6]), .Z(n1833) );
  AND U1907 ( .A(a[5]), .B(b[7]), .Z(n1832) );
  XOR U1908 ( .A(n1834), .B(n1830), .Z(n1827) );
  XOR U1909 ( .A(n1835), .B(n1836), .Z(n1830) );
  NOR U1910 ( .A(n1837), .B(n1838), .Z(n1835) );
  AND U1911 ( .A(a[7]), .B(b[5]), .Z(n1834) );
  XNOR U1912 ( .A(n1839), .B(n1798), .Z(n1799) );
  XOR U1913 ( .A(n1840), .B(n1841), .Z(n1798) );
  ANDN U1914 ( .B(n1842), .A(n1843), .Z(n1840) );
  AND U1915 ( .A(b[4]), .B(a[8]), .Z(n1839) );
  XNOR U1916 ( .A(n1844), .B(n1845), .Z(n1812) );
  NANDN U1917 ( .A(n1846), .B(n1847), .Z(n1845) );
  XNOR U1918 ( .A(n1848), .B(n1803), .Z(n1805) );
  XNOR U1919 ( .A(n1849), .B(n1850), .Z(n1803) );
  AND U1920 ( .A(n1851), .B(n1852), .Z(n1849) );
  AND U1921 ( .A(b[3]), .B(a[9]), .Z(n1848) );
  XOR U1922 ( .A(n1819), .B(n1818), .Z(swire[11]) );
  XOR U1923 ( .A(sreg[75]), .B(n1817), .Z(n1818) );
  XOR U1924 ( .A(n1824), .B(n1853), .Z(n1819) );
  XNOR U1925 ( .A(n1823), .B(n1817), .Z(n1853) );
  XOR U1926 ( .A(n1854), .B(n1855), .Z(n1817) );
  NOR U1927 ( .A(n1856), .B(n1857), .Z(n1854) );
  NANDN U1928 ( .A(n11), .B(a[11]), .Z(n1823) );
  XNOR U1929 ( .A(n1846), .B(n1847), .Z(n1824) );
  XOR U1930 ( .A(n1844), .B(n1858), .Z(n1847) );
  NAND U1931 ( .A(b[1]), .B(a[10]), .Z(n1858) );
  XOR U1932 ( .A(n1852), .B(n1859), .Z(n1846) );
  XOR U1933 ( .A(n1844), .B(n1851), .Z(n1859) );
  XNOR U1934 ( .A(n1860), .B(n1850), .Z(n1851) );
  AND U1935 ( .A(b[2]), .B(a[9]), .Z(n1860) );
  NANDN U1936 ( .A(n1861), .B(n1862), .Z(n1844) );
  XOR U1937 ( .A(n1850), .B(n1842), .Z(n1863) );
  XOR U1938 ( .A(n1841), .B(n1838), .Z(n1864) );
  XOR U1939 ( .A(n1865), .B(n1866), .Z(n1838) );
  XOR U1940 ( .A(n1836), .B(n1867), .Z(n1866) );
  XOR U1941 ( .A(n1868), .B(n1869), .Z(n1867) );
  XOR U1942 ( .A(n1870), .B(n1871), .Z(n1869) );
  NAND U1943 ( .A(a[5]), .B(b[6]), .Z(n1871) );
  AND U1944 ( .A(a[4]), .B(b[7]), .Z(n1870) );
  XOR U1945 ( .A(n1872), .B(n1868), .Z(n1865) );
  XOR U1946 ( .A(n1873), .B(n1874), .Z(n1868) );
  NOR U1947 ( .A(n1875), .B(n1876), .Z(n1873) );
  AND U1948 ( .A(b[5]), .B(a[6]), .Z(n1872) );
  XNOR U1949 ( .A(n1877), .B(n1836), .Z(n1837) );
  XOR U1950 ( .A(n1878), .B(n1879), .Z(n1836) );
  ANDN U1951 ( .B(n1880), .A(n1881), .Z(n1878) );
  AND U1952 ( .A(a[7]), .B(b[4]), .Z(n1877) );
  XNOR U1953 ( .A(n1882), .B(n1883), .Z(n1850) );
  NANDN U1954 ( .A(n1884), .B(n1885), .Z(n1883) );
  XNOR U1955 ( .A(n1886), .B(n1841), .Z(n1843) );
  XNOR U1956 ( .A(n1887), .B(n1888), .Z(n1841) );
  AND U1957 ( .A(n1889), .B(n1890), .Z(n1887) );
  AND U1958 ( .A(b[3]), .B(a[8]), .Z(n1886) );
  XOR U1959 ( .A(n1857), .B(n1856), .Z(swire[10]) );
  XOR U1960 ( .A(sreg[74]), .B(n1855), .Z(n1856) );
  XOR U1961 ( .A(n1862), .B(n1891), .Z(n1857) );
  XNOR U1962 ( .A(n1861), .B(n1855), .Z(n1891) );
  XOR U1963 ( .A(n1892), .B(n1893), .Z(n1855) );
  ANDN U1964 ( .B(n2), .A(n1), .Z(n1892) );
  XOR U1965 ( .A(sreg[73]), .B(n1893), .Z(n1) );
  XOR U1966 ( .A(n1894), .B(n1895), .Z(n2) );
  XNOR U1967 ( .A(n1896), .B(n1893), .Z(n1895) );
  XOR U1968 ( .A(n1897), .B(n1898), .Z(n1893) );
  ANDN U1969 ( .B(n3), .A(n4), .Z(n1897) );
  XOR U1970 ( .A(sreg[72]), .B(n1898), .Z(n4) );
  XOR U1971 ( .A(n1899), .B(n1900), .Z(n3) );
  XNOR U1972 ( .A(n1901), .B(n1898), .Z(n1900) );
  XOR U1973 ( .A(n1902), .B(n1903), .Z(n1898) );
  ANDN U1974 ( .B(n1904), .A(n1905), .Z(n1902) );
  NANDN U1975 ( .A(n11), .B(a[10]), .Z(n1861) );
  XNOR U1976 ( .A(n1884), .B(n1885), .Z(n1862) );
  XOR U1977 ( .A(n1882), .B(n1906), .Z(n1885) );
  NAND U1978 ( .A(b[1]), .B(a[9]), .Z(n1906) );
  XOR U1979 ( .A(n1890), .B(n1907), .Z(n1884) );
  XOR U1980 ( .A(n1882), .B(n1889), .Z(n1907) );
  XNOR U1981 ( .A(n1908), .B(n1888), .Z(n1889) );
  AND U1982 ( .A(b[2]), .B(a[8]), .Z(n1908) );
  OR U1983 ( .A(n1896), .B(n1894), .Z(n1882) );
  XOR U1984 ( .A(n1909), .B(n1910), .Z(n1894) );
  NANDN U1985 ( .A(n11), .B(a[9]), .Z(n1896) );
  XOR U1986 ( .A(n1888), .B(n1880), .Z(n1911) );
  XOR U1987 ( .A(n1879), .B(n1876), .Z(n1912) );
  XOR U1988 ( .A(n1913), .B(n1914), .Z(n1876) );
  XOR U1989 ( .A(n1874), .B(n1915), .Z(n1914) );
  XNOR U1990 ( .A(n1916), .B(n1917), .Z(n1915) );
  XOR U1991 ( .A(n1918), .B(n1919), .Z(n1917) );
  NAND U1992 ( .A(a[4]), .B(b[6]), .Z(n1919) );
  AND U1993 ( .A(a[3]), .B(b[7]), .Z(n1918) );
  XNOR U1994 ( .A(n1920), .B(n1916), .Z(n1913) );
  XOR U1995 ( .A(n1921), .B(n1922), .Z(n1916) );
  NOR U1996 ( .A(n1923), .B(n1924), .Z(n1921) );
  AND U1997 ( .A(a[5]), .B(b[5]), .Z(n1920) );
  XNOR U1998 ( .A(n1925), .B(n1874), .Z(n1875) );
  XNOR U1999 ( .A(n1926), .B(n1927), .Z(n1874) );
  ANDN U2000 ( .B(n1928), .A(n1929), .Z(n1926) );
  AND U2001 ( .A(b[4]), .B(a[6]), .Z(n1925) );
  XNOR U2002 ( .A(n1930), .B(n1931), .Z(n1888) );
  NANDN U2003 ( .A(n1910), .B(n1909), .Z(n1931) );
  XOR U2004 ( .A(n1930), .B(n1932), .Z(n1909) );
  NAND U2005 ( .A(b[1]), .B(a[8]), .Z(n1932) );
  XOR U2006 ( .A(n1930), .B(n1934), .Z(n1933) );
  OR U2007 ( .A(n1901), .B(n1899), .Z(n1930) );
  XOR U2008 ( .A(n1936), .B(n1937), .Z(n1899) );
  NANDN U2009 ( .A(n11), .B(a[8]), .Z(n1901) );
  XNOR U2010 ( .A(n1938), .B(n1879), .Z(n1881) );
  XNOR U2011 ( .A(n1939), .B(n1940), .Z(n1879) );
  ANDN U2012 ( .B(n1934), .A(n1935), .Z(n1939) );
  XOR U2013 ( .A(n1941), .B(n1940), .Z(n1935) );
  IV U2014 ( .A(n1942), .Z(n1940) );
  AND U2015 ( .A(a[7]), .B(b[2]), .Z(n1941) );
  XNOR U2016 ( .A(n1928), .B(n1942), .Z(n1943) );
  XOR U2017 ( .A(n1944), .B(n1945), .Z(n1942) );
  NANDN U2018 ( .A(n1937), .B(n1936), .Z(n1945) );
  XOR U2019 ( .A(n1944), .B(n1946), .Z(n1936) );
  NAND U2020 ( .A(a[7]), .B(b[1]), .Z(n1946) );
  XOR U2021 ( .A(n1944), .B(n1948), .Z(n1947) );
  OR U2022 ( .A(n1950), .B(n1951), .Z(n1944) );
  XOR U2023 ( .A(n1924), .B(n1953), .Z(n1952) );
  XOR U2024 ( .A(n1954), .B(n1955), .Z(n1924) );
  XNOR U2025 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U2026 ( .A(n1958), .B(n1959), .Z(n1956) );
  XOR U2027 ( .A(n1960), .B(n1961), .Z(n1959) );
  AND U2028 ( .A(a[2]), .B(b[7]), .Z(n1961) );
  AND U2029 ( .A(a[3]), .B(b[6]), .Z(n1960) );
  XNOR U2030 ( .A(n1962), .B(n1958), .Z(n1954) );
  XNOR U2031 ( .A(n1963), .B(n1964), .Z(n1958) );
  NOR U2032 ( .A(n1965), .B(n1966), .Z(n1963) );
  AND U2033 ( .A(a[4]), .B(b[5]), .Z(n1962) );
  XOR U2034 ( .A(n1967), .B(n1922), .Z(n1923) );
  IV U2035 ( .A(n1957), .Z(n1922) );
  XOR U2036 ( .A(n1968), .B(n1969), .Z(n1957) );
  ANDN U2037 ( .B(n1970), .A(n1971), .Z(n1968) );
  AND U2038 ( .A(a[5]), .B(b[4]), .Z(n1967) );
  XOR U2039 ( .A(n1972), .B(n1927), .Z(n1929) );
  IV U2040 ( .A(n1953), .Z(n1927) );
  XOR U2041 ( .A(n1973), .B(n1974), .Z(n1953) );
  ANDN U2042 ( .B(n1948), .A(n1949), .Z(n1973) );
  AND U2043 ( .A(b[2]), .B(a[6]), .Z(n1975) );
  XNOR U2044 ( .A(n1970), .B(n1974), .Z(n1976) );
  XOR U2045 ( .A(n1977), .B(n1978), .Z(n1974) );
  OR U2046 ( .A(n1979), .B(n1980), .Z(n1978) );
  XOR U2047 ( .A(n1966), .B(n1969), .Z(n1981) );
  XOR U2048 ( .A(n1982), .B(n1983), .Z(n1966) );
  XNOR U2049 ( .A(n1984), .B(n1964), .Z(n1983) );
  XOR U2050 ( .A(n1985), .B(n1986), .Z(n1984) );
  XOR U2051 ( .A(n1987), .B(n1988), .Z(n1986) );
  AND U2052 ( .A(a[2]), .B(b[6]), .Z(n1988) );
  AND U2053 ( .A(a[1]), .B(b[7]), .Z(n1987) );
  XOR U2054 ( .A(n1989), .B(n1985), .Z(n1982) );
  XOR U2055 ( .A(n1990), .B(n1991), .Z(n1985) );
  NOR U2056 ( .A(n1992), .B(n1993), .Z(n1990) );
  AND U2057 ( .A(a[3]), .B(b[5]), .Z(n1989) );
  XNOR U2058 ( .A(n1994), .B(n1964), .Z(n1965) );
  XOR U2059 ( .A(n1995), .B(n1996), .Z(n1964) );
  ANDN U2060 ( .B(n1997), .A(n1998), .Z(n1995) );
  AND U2061 ( .A(b[4]), .B(a[4]), .Z(n1994) );
  XNOR U2062 ( .A(n1999), .B(n1969), .Z(n1971) );
  XNOR U2063 ( .A(n2000), .B(n2001), .Z(n1969) );
  NOR U2064 ( .A(n2002), .B(n2003), .Z(n2000) );
  AND U2065 ( .A(a[5]), .B(b[3]), .Z(n1999) );
  AND U2066 ( .A(b[3]), .B(a[6]), .Z(n1972) );
  AND U2067 ( .A(a[7]), .B(b[3]), .Z(n1938) );
  XNOR U2068 ( .A(n1904), .B(n1905), .Z(c[63]) );
  XOR U2069 ( .A(sreg[71]), .B(n1903), .Z(n1905) );
  XOR U2070 ( .A(n1951), .B(n2004), .Z(n1904) );
  XNOR U2071 ( .A(n1950), .B(n1903), .Z(n2004) );
  XOR U2072 ( .A(n2005), .B(n2006), .Z(n1903) );
  ANDN U2073 ( .B(n2007), .A(n2008), .Z(n2005) );
  NANDN U2074 ( .A(n11), .B(a[7]), .Z(n1950) );
  XNOR U2075 ( .A(n1977), .B(n2009), .Z(n1979) );
  NAND U2076 ( .A(b[1]), .B(a[6]), .Z(n2009) );
  XNOR U2077 ( .A(n1977), .B(n2003), .Z(n2010) );
  XOR U2078 ( .A(n2011), .B(n2001), .Z(n2003) );
  AND U2079 ( .A(a[5]), .B(b[2]), .Z(n2011) );
  OR U2080 ( .A(n2012), .B(n2013), .Z(n1977) );
  XOR U2081 ( .A(n2001), .B(n1997), .Z(n2014) );
  XOR U2082 ( .A(n1996), .B(n1993), .Z(n2015) );
  XOR U2083 ( .A(n2016), .B(n2017), .Z(n1993) );
  XOR U2084 ( .A(n1991), .B(n2018), .Z(n2017) );
  XOR U2085 ( .A(n2019), .B(n2020), .Z(n2018) );
  XOR U2086 ( .A(n2021), .B(n2022), .Z(n2020) );
  NAND U2087 ( .A(a[1]), .B(b[6]), .Z(n2022) );
  AND U2088 ( .A(a[0]), .B(b[7]), .Z(n2021) );
  XOR U2089 ( .A(n2023), .B(n2019), .Z(n2016) );
  XOR U2090 ( .A(n2024), .B(n2025), .Z(n2019) );
  NOR U2091 ( .A(n2026), .B(n2027), .Z(n2024) );
  AND U2092 ( .A(a[2]), .B(b[5]), .Z(n2023) );
  XNOR U2093 ( .A(n2028), .B(n1991), .Z(n1992) );
  XOR U2094 ( .A(n2029), .B(n2030), .Z(n1991) );
  ANDN U2095 ( .B(n2031), .A(n2032), .Z(n2029) );
  AND U2096 ( .A(a[3]), .B(b[4]), .Z(n2028) );
  XNOR U2097 ( .A(n2033), .B(n2034), .Z(n2001) );
  OR U2098 ( .A(n2035), .B(n2036), .Z(n2034) );
  XNOR U2099 ( .A(n2037), .B(n1996), .Z(n1998) );
  XNOR U2100 ( .A(n2038), .B(n2039), .Z(n1996) );
  NOR U2101 ( .A(n2040), .B(n2041), .Z(n2038) );
  AND U2102 ( .A(b[3]), .B(a[4]), .Z(n2037) );
  XNOR U2103 ( .A(n2007), .B(n2008), .Z(c[62]) );
  XOR U2104 ( .A(sreg[70]), .B(n2006), .Z(n2008) );
  XOR U2105 ( .A(n2013), .B(n2042), .Z(n2007) );
  XNOR U2106 ( .A(n2012), .B(n2006), .Z(n2042) );
  XOR U2107 ( .A(n2043), .B(n2044), .Z(n2006) );
  ANDN U2108 ( .B(n2045), .A(n2046), .Z(n2043) );
  NANDN U2109 ( .A(n11), .B(a[6]), .Z(n2012) );
  XNOR U2110 ( .A(n2033), .B(n2047), .Z(n2035) );
  NAND U2111 ( .A(a[5]), .B(b[1]), .Z(n2047) );
  XNOR U2112 ( .A(n2033), .B(n2041), .Z(n2048) );
  XOR U2113 ( .A(n2049), .B(n2039), .Z(n2041) );
  AND U2114 ( .A(b[2]), .B(a[4]), .Z(n2049) );
  OR U2115 ( .A(n2050), .B(n2051), .Z(n2033) );
  XOR U2116 ( .A(n2052), .B(n2053), .Z(n2040) );
  XOR U2117 ( .A(n2039), .B(n2031), .Z(n2053) );
  XOR U2118 ( .A(n2030), .B(n2027), .Z(n2054) );
  XOR U2119 ( .A(n2055), .B(n2056), .Z(n2027) );
  XOR U2120 ( .A(n2025), .B(n2057), .Z(n2056) );
  XOR U2121 ( .A(n2058), .B(n2059), .Z(n2057) );
  AND U2122 ( .A(a[0]), .B(b[6]), .Z(n2058) );
  XNOR U2123 ( .A(n2060), .B(n2059), .Z(n2055) );
  XOR U2124 ( .A(n2061), .B(n2062), .Z(n2059) );
  NOR U2125 ( .A(n2063), .B(n2064), .Z(n2061) );
  AND U2126 ( .A(a[1]), .B(b[5]), .Z(n2060) );
  XNOR U2127 ( .A(n2065), .B(n2025), .Z(n2026) );
  XOR U2128 ( .A(n2066), .B(n2067), .Z(n2025) );
  NOR U2129 ( .A(n2068), .B(n2069), .Z(n2066) );
  AND U2130 ( .A(a[2]), .B(b[4]), .Z(n2065) );
  XNOR U2131 ( .A(n2070), .B(n2071), .Z(n2039) );
  OR U2132 ( .A(n2072), .B(n2073), .Z(n2071) );
  IV U2133 ( .A(n2032), .Z(n2052) );
  XNOR U2134 ( .A(n2074), .B(n2030), .Z(n2032) );
  XNOR U2135 ( .A(n2075), .B(n2076), .Z(n2030) );
  NOR U2136 ( .A(n2077), .B(n2078), .Z(n2075) );
  AND U2137 ( .A(a[3]), .B(b[3]), .Z(n2074) );
  XNOR U2138 ( .A(n2045), .B(n2046), .Z(c[61]) );
  XOR U2139 ( .A(sreg[69]), .B(n2044), .Z(n2046) );
  XOR U2140 ( .A(n2051), .B(n2079), .Z(n2045) );
  XNOR U2141 ( .A(n2050), .B(n2044), .Z(n2079) );
  XOR U2142 ( .A(n2080), .B(n2081), .Z(n2044) );
  ANDN U2143 ( .B(n2082), .A(n2083), .Z(n2080) );
  NANDN U2144 ( .A(n11), .B(a[5]), .Z(n2050) );
  XNOR U2145 ( .A(n2070), .B(n2084), .Z(n2072) );
  NAND U2146 ( .A(b[1]), .B(a[4]), .Z(n2084) );
  XNOR U2147 ( .A(n2070), .B(n2078), .Z(n2085) );
  XOR U2148 ( .A(n2086), .B(n2076), .Z(n2078) );
  AND U2149 ( .A(b[2]), .B(a[3]), .Z(n2086) );
  OR U2150 ( .A(n2087), .B(n2088), .Z(n2070) );
  XNOR U2151 ( .A(n2076), .B(n2069), .Z(n2089) );
  XOR U2152 ( .A(n2063), .B(n2090), .Z(n2069) );
  XNOR U2153 ( .A(n2067), .B(n2064), .Z(n2090) );
  XNOR U2154 ( .A(n2091), .B(n2062), .Z(n2064) );
  AND U2155 ( .A(a[0]), .B(b[5]), .Z(n2091) );
  XNOR U2156 ( .A(n2092), .B(n2062), .Z(n2063) );
  XOR U2157 ( .A(n2093), .B(n2094), .Z(n2062) );
  NOR U2158 ( .A(n2095), .B(n2096), .Z(n2093) );
  AND U2159 ( .A(a[1]), .B(b[4]), .Z(n2092) );
  XNOR U2160 ( .A(n2097), .B(n2098), .Z(n2076) );
  OR U2161 ( .A(n2099), .B(n2100), .Z(n2098) );
  XNOR U2162 ( .A(n2101), .B(n2067), .Z(n2068) );
  XNOR U2163 ( .A(n2102), .B(n2103), .Z(n2067) );
  NOR U2164 ( .A(n2104), .B(n2105), .Z(n2102) );
  AND U2165 ( .A(a[2]), .B(b[3]), .Z(n2101) );
  XNOR U2166 ( .A(n2082), .B(n2083), .Z(c[60]) );
  XOR U2167 ( .A(sreg[68]), .B(n2081), .Z(n2083) );
  XOR U2168 ( .A(n2088), .B(n2106), .Z(n2082) );
  XNOR U2169 ( .A(n2087), .B(n2081), .Z(n2106) );
  XOR U2170 ( .A(n2107), .B(n2108), .Z(n2081) );
  ANDN U2171 ( .B(n2109), .A(n2110), .Z(n2107) );
  NANDN U2172 ( .A(n11), .B(a[4]), .Z(n2087) );
  XNOR U2173 ( .A(n2097), .B(n2111), .Z(n2099) );
  NAND U2174 ( .A(a[3]), .B(b[1]), .Z(n2111) );
  XNOR U2175 ( .A(n2097), .B(n2105), .Z(n2112) );
  XOR U2176 ( .A(n2113), .B(n2103), .Z(n2105) );
  AND U2177 ( .A(b[2]), .B(a[2]), .Z(n2113) );
  OR U2178 ( .A(n2114), .B(n2115), .Z(n2097) );
  XOR U2179 ( .A(n2095), .B(n2116), .Z(n2104) );
  XOR U2180 ( .A(n2103), .B(n2096), .Z(n2116) );
  XNOR U2181 ( .A(n2117), .B(n2094), .Z(n2096) );
  AND U2182 ( .A(a[0]), .B(b[4]), .Z(n2117) );
  XOR U2183 ( .A(n2118), .B(n2119), .Z(n2103) );
  OR U2184 ( .A(n2120), .B(n2121), .Z(n2119) );
  XNOR U2185 ( .A(n2122), .B(n2094), .Z(n2095) );
  XOR U2186 ( .A(n2123), .B(n2124), .Z(n2094) );
  NOR U2187 ( .A(n2125), .B(n2126), .Z(n2123) );
  AND U2188 ( .A(a[1]), .B(b[3]), .Z(n2122) );
  XNOR U2189 ( .A(n2109), .B(n2110), .Z(c[59]) );
  XOR U2190 ( .A(sreg[67]), .B(n2108), .Z(n2110) );
  XOR U2191 ( .A(n2115), .B(n2127), .Z(n2109) );
  XNOR U2192 ( .A(n2114), .B(n2108), .Z(n2127) );
  XNOR U2193 ( .A(n2128), .B(n2129), .Z(n2108) );
  ANDN U2194 ( .B(n2130), .A(n2131), .Z(n2128) );
  NANDN U2195 ( .A(n11), .B(a[3]), .Z(n2114) );
  XOR U2196 ( .A(n2118), .B(n2132), .Z(n2120) );
  NAND U2197 ( .A(b[1]), .B(a[2]), .Z(n2132) );
  XOR U2198 ( .A(n2125), .B(n2133), .Z(n2121) );
  XNOR U2199 ( .A(n2118), .B(n2126), .Z(n2133) );
  XNOR U2200 ( .A(n2134), .B(n2124), .Z(n2126) );
  AND U2201 ( .A(b[2]), .B(a[1]), .Z(n2134) );
  NOR U2202 ( .A(n2135), .B(n2136), .Z(n2118) );
  XNOR U2203 ( .A(n2137), .B(n2124), .Z(n2125) );
  NAND U2204 ( .A(n2138), .B(n2139), .Z(n2124) );
  OR U2205 ( .A(n2140), .B(n2141), .Z(n2139) );
  AND U2206 ( .A(a[0]), .B(b[3]), .Z(n2137) );
  XNOR U2207 ( .A(n2130), .B(n2131), .Z(c[58]) );
  XNOR U2208 ( .A(sreg[66]), .B(n2129), .Z(n2131) );
  XNOR U2209 ( .A(n2136), .B(n2143), .Z(n2142) );
  IV U2210 ( .A(n2129), .Z(n2143) );
  XNOR U2211 ( .A(n2144), .B(n2145), .Z(n2129) );
  NAND U2212 ( .A(n2146), .B(n2147), .Z(n2145) );
  NANDN U2213 ( .A(n11), .B(a[2]), .Z(n2136) );
  XOR U2214 ( .A(n2148), .B(n2138), .Z(n2141) );
  AND U2215 ( .A(b[2]), .B(a[0]), .Z(n2148) );
  NAND U2216 ( .A(n2149), .B(b[1]), .Z(n2140) );
  NANDN U2217 ( .A(n2150), .B(n2151), .Z(n2138) );
  XOR U2218 ( .A(n2146), .B(n2147), .Z(c[57]) );
  XOR U2219 ( .A(sreg[65]), .B(n2144), .Z(n2147) );
  XNOR U2220 ( .A(n2144), .B(n2152), .Z(n2146) );
  XOR U2221 ( .A(n2150), .B(n2151), .Z(n2152) );
  AND U2222 ( .A(a[1]), .B(b[0]), .Z(n2151) );
  NAND U2223 ( .A(b[1]), .B(a[0]), .Z(n2150) );
  ANDN U2224 ( .B(sreg[64]), .A(n2153), .Z(n2144) );
  XNOR U2225 ( .A(sreg[64]), .B(n2153), .Z(c[56]) );
  NANDN U2226 ( .A(n11), .B(a[0]), .Z(n2153) );
  IV U2227 ( .A(b[0]), .Z(n11) );
endmodule

