
module matrixMult_N_M_1_N3_M8 ( clk, rst, x, y, o );
  input [23:0] x;
  input [71:0] y;
  output [23:0] o;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N25, N26, N27, N28, N29, N30,
         N31, N32, N41, N42, N43, N44, N45, N46, N47, N48, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522;

  DFF \oi_reg[0][7]  ( .D(N16), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N15), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N14), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N13), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N12), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N11), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N10), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N9), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][7]  ( .D(N32), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[1][6]  ( .D(N31), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[1][5]  ( .D(N30), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[1][4]  ( .D(N29), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[1][3]  ( .D(N28), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[1][2]  ( .D(N27), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[1][1]  ( .D(N26), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[1][0]  ( .D(N25), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[2][7]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[2][6]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[2][5]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[2][4]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[2][3]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[2][2]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[2][1]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[2][0]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[16]) );
  NAND U3 ( .A(n445), .B(n446), .Z(n1) );
  XOR U4 ( .A(n445), .B(n446), .Z(n2) );
  NANDN U5 ( .A(n444), .B(n2), .Z(n3) );
  NAND U6 ( .A(n1), .B(n3), .Z(n458) );
  NAND U7 ( .A(n317), .B(n318), .Z(n4) );
  XOR U8 ( .A(n317), .B(n318), .Z(n5) );
  NANDN U9 ( .A(n316), .B(n5), .Z(n6) );
  NAND U10 ( .A(n4), .B(n6), .Z(n330) );
  NAND U11 ( .A(n189), .B(n190), .Z(n7) );
  XOR U12 ( .A(n189), .B(n190), .Z(n8) );
  NANDN U13 ( .A(n188), .B(n8), .Z(n9) );
  NAND U14 ( .A(n7), .B(n9), .Z(n202) );
  XOR U15 ( .A(n507), .B(n506), .Z(n10) );
  XNOR U16 ( .A(n509), .B(n10), .Z(n479) );
  XOR U17 ( .A(n379), .B(n378), .Z(n11) );
  XNOR U18 ( .A(n381), .B(n11), .Z(n351) );
  XOR U19 ( .A(n251), .B(n250), .Z(n12) );
  XNOR U20 ( .A(n253), .B(n12), .Z(n223) );
  NAND U21 ( .A(n442), .B(n443), .Z(n13) );
  XOR U22 ( .A(n442), .B(n443), .Z(n14) );
  NANDN U23 ( .A(n441), .B(n14), .Z(n15) );
  NAND U24 ( .A(n13), .B(n15), .Z(n457) );
  NAND U25 ( .A(n314), .B(n315), .Z(n16) );
  XOR U26 ( .A(n314), .B(n315), .Z(n17) );
  NANDN U27 ( .A(n313), .B(n17), .Z(n18) );
  NAND U28 ( .A(n16), .B(n18), .Z(n329) );
  NAND U29 ( .A(n186), .B(n187), .Z(n19) );
  XOR U30 ( .A(n186), .B(n187), .Z(n20) );
  NANDN U31 ( .A(n185), .B(n20), .Z(n21) );
  NAND U32 ( .A(n19), .B(n21), .Z(n201) );
  NAND U33 ( .A(n467), .B(n468), .Z(n22) );
  XOR U34 ( .A(n467), .B(n468), .Z(n23) );
  NANDN U35 ( .A(n466), .B(n23), .Z(n24) );
  NAND U36 ( .A(n22), .B(n24), .Z(n513) );
  NAND U37 ( .A(n339), .B(n340), .Z(n25) );
  XOR U38 ( .A(n339), .B(n340), .Z(n26) );
  NANDN U39 ( .A(n338), .B(n26), .Z(n27) );
  NAND U40 ( .A(n25), .B(n27), .Z(n385) );
  NAND U41 ( .A(n211), .B(n212), .Z(n28) );
  XOR U42 ( .A(n211), .B(n212), .Z(n29) );
  NANDN U43 ( .A(n210), .B(n29), .Z(n30) );
  NAND U44 ( .A(n28), .B(n30), .Z(n257) );
  NAND U45 ( .A(n473), .B(n471), .Z(n31) );
  XOR U46 ( .A(n473), .B(n471), .Z(n32) );
  NANDN U47 ( .A(n472), .B(n32), .Z(n33) );
  NAND U48 ( .A(n31), .B(n33), .Z(n476) );
  NAND U49 ( .A(n345), .B(n343), .Z(n34) );
  XOR U50 ( .A(n345), .B(n343), .Z(n35) );
  NANDN U51 ( .A(n344), .B(n35), .Z(n36) );
  NAND U52 ( .A(n34), .B(n36), .Z(n348) );
  NAND U53 ( .A(n217), .B(n215), .Z(n37) );
  XOR U54 ( .A(n217), .B(n215), .Z(n38) );
  NANDN U55 ( .A(n216), .B(n38), .Z(n39) );
  NAND U56 ( .A(n37), .B(n39), .Z(n220) );
  NAND U57 ( .A(n433), .B(n434), .Z(n40) );
  XOR U58 ( .A(n433), .B(n434), .Z(n41) );
  NANDN U59 ( .A(n432), .B(n41), .Z(n42) );
  NAND U60 ( .A(n40), .B(n42), .Z(n452) );
  NAND U61 ( .A(n464), .B(n465), .Z(n43) );
  XOR U62 ( .A(n464), .B(n465), .Z(n44) );
  NANDN U63 ( .A(n463), .B(n44), .Z(n45) );
  NAND U64 ( .A(n43), .B(n45), .Z(n514) );
  NAND U65 ( .A(n305), .B(n306), .Z(n46) );
  XOR U66 ( .A(n305), .B(n306), .Z(n47) );
  NANDN U67 ( .A(n304), .B(n47), .Z(n48) );
  NAND U68 ( .A(n46), .B(n48), .Z(n324) );
  NAND U69 ( .A(n336), .B(n337), .Z(n49) );
  XOR U70 ( .A(n336), .B(n337), .Z(n50) );
  NANDN U71 ( .A(n335), .B(n50), .Z(n51) );
  NAND U72 ( .A(n49), .B(n51), .Z(n386) );
  NAND U73 ( .A(n177), .B(n178), .Z(n52) );
  XOR U74 ( .A(n177), .B(n178), .Z(n53) );
  NANDN U75 ( .A(n176), .B(n53), .Z(n54) );
  NAND U76 ( .A(n52), .B(n54), .Z(n196) );
  NAND U77 ( .A(n208), .B(n209), .Z(n55) );
  XOR U78 ( .A(n208), .B(n209), .Z(n56) );
  NANDN U79 ( .A(n207), .B(n56), .Z(n57) );
  NAND U80 ( .A(n55), .B(n57), .Z(n258) );
  XOR U81 ( .A(n479), .B(n478), .Z(n477) );
  XOR U82 ( .A(n351), .B(n350), .Z(n349) );
  XOR U83 ( .A(n223), .B(n222), .Z(n221) );
  NAND U84 ( .A(n428), .B(n426), .Z(n58) );
  XOR U85 ( .A(n428), .B(n426), .Z(n59) );
  NANDN U86 ( .A(n427), .B(n59), .Z(n60) );
  NAND U87 ( .A(n58), .B(n60), .Z(n434) );
  NAND U88 ( .A(n300), .B(n298), .Z(n61) );
  XOR U89 ( .A(n300), .B(n298), .Z(n62) );
  NANDN U90 ( .A(n299), .B(n62), .Z(n63) );
  NAND U91 ( .A(n61), .B(n63), .Z(n306) );
  NAND U92 ( .A(n172), .B(n170), .Z(n64) );
  XOR U93 ( .A(n172), .B(n170), .Z(n65) );
  NANDN U94 ( .A(n171), .B(n65), .Z(n66) );
  NAND U95 ( .A(n64), .B(n66), .Z(n178) );
  XOR U96 ( .A(n520), .B(n519), .Z(n518) );
  NANDN U97 ( .A(n511), .B(n512), .Z(n516) );
  XOR U98 ( .A(n392), .B(n391), .Z(n390) );
  NANDN U99 ( .A(n383), .B(n384), .Z(n388) );
  XOR U100 ( .A(n264), .B(n263), .Z(n262) );
  NANDN U101 ( .A(n255), .B(n256), .Z(n260) );
  NAND U102 ( .A(n406), .B(n404), .Z(n67) );
  XOR U103 ( .A(n406), .B(n404), .Z(n68) );
  NANDN U104 ( .A(n405), .B(n68), .Z(n69) );
  NAND U105 ( .A(n67), .B(n69), .Z(n420) );
  XOR U106 ( .A(n418), .B(n416), .Z(n70) );
  NANDN U107 ( .A(n417), .B(n70), .Z(n71) );
  NAND U108 ( .A(n418), .B(n416), .Z(n72) );
  AND U109 ( .A(n71), .B(n72), .Z(n436) );
  NAND U110 ( .A(n278), .B(n276), .Z(n73) );
  XOR U111 ( .A(n278), .B(n276), .Z(n74) );
  NANDN U112 ( .A(n277), .B(n74), .Z(n75) );
  NAND U113 ( .A(n73), .B(n75), .Z(n292) );
  XOR U114 ( .A(n290), .B(n288), .Z(n76) );
  NANDN U115 ( .A(n289), .B(n76), .Z(n77) );
  NAND U116 ( .A(n290), .B(n288), .Z(n78) );
  AND U117 ( .A(n77), .B(n78), .Z(n308) );
  NAND U118 ( .A(n150), .B(n148), .Z(n79) );
  XOR U119 ( .A(n150), .B(n148), .Z(n80) );
  NANDN U120 ( .A(n149), .B(n80), .Z(n81) );
  NAND U121 ( .A(n79), .B(n81), .Z(n164) );
  XOR U122 ( .A(n162), .B(n160), .Z(n82) );
  NANDN U123 ( .A(n161), .B(n82), .Z(n83) );
  NAND U124 ( .A(n162), .B(n160), .Z(n84) );
  AND U125 ( .A(n83), .B(n84), .Z(n180) );
  AND U126 ( .A(n522), .B(n521), .Z(n85) );
  NAND U127 ( .A(n516), .B(n515), .Z(n86) );
  XNOR U128 ( .A(n85), .B(n86), .Z(n87) );
  NAND U129 ( .A(n507), .B(n506), .Z(n88) );
  NAND U130 ( .A(n510), .B(n88), .Z(n89) );
  XNOR U131 ( .A(n87), .B(n89), .Z(n90) );
  NAND U132 ( .A(n479), .B(n478), .Z(n91) );
  NAND U133 ( .A(n480), .B(n481), .Z(n92) );
  AND U134 ( .A(n91), .B(n92), .Z(n93) );
  AND U135 ( .A(n505), .B(n504), .Z(n94) );
  XNOR U136 ( .A(n499), .B(n498), .Z(n95) );
  XNOR U137 ( .A(n94), .B(n95), .Z(n96) );
  XNOR U138 ( .A(n93), .B(n96), .Z(n97) );
  XNOR U139 ( .A(n90), .B(n97), .Z(n98) );
  NANDN U140 ( .A(n475), .B(n476), .Z(n99) );
  XNOR U141 ( .A(n475), .B(n476), .Z(n100) );
  NAND U142 ( .A(n477), .B(n100), .Z(n101) );
  AND U143 ( .A(n99), .B(n101), .Z(n102) );
  XNOR U144 ( .A(n98), .B(n102), .Z(N48) );
  AND U145 ( .A(n394), .B(n393), .Z(n103) );
  NAND U146 ( .A(n388), .B(n387), .Z(n104) );
  XNOR U147 ( .A(n103), .B(n104), .Z(n105) );
  NAND U148 ( .A(n379), .B(n378), .Z(n106) );
  NAND U149 ( .A(n382), .B(n106), .Z(n107) );
  XNOR U150 ( .A(n105), .B(n107), .Z(n108) );
  NAND U151 ( .A(n351), .B(n350), .Z(n109) );
  NAND U152 ( .A(n352), .B(n353), .Z(n110) );
  AND U153 ( .A(n109), .B(n110), .Z(n111) );
  AND U154 ( .A(n377), .B(n376), .Z(n112) );
  XNOR U155 ( .A(n371), .B(n370), .Z(n113) );
  XNOR U156 ( .A(n112), .B(n113), .Z(n114) );
  XNOR U157 ( .A(n111), .B(n114), .Z(n115) );
  XNOR U158 ( .A(n108), .B(n115), .Z(n116) );
  NANDN U159 ( .A(n347), .B(n348), .Z(n117) );
  XNOR U160 ( .A(n347), .B(n348), .Z(n118) );
  NAND U161 ( .A(n349), .B(n118), .Z(n119) );
  AND U162 ( .A(n117), .B(n119), .Z(n120) );
  XNOR U163 ( .A(n116), .B(n120), .Z(N32) );
  NAND U164 ( .A(n223), .B(n222), .Z(n121) );
  NAND U165 ( .A(n224), .B(n225), .Z(n122) );
  AND U166 ( .A(n121), .B(n122), .Z(n123) );
  AND U167 ( .A(n249), .B(n248), .Z(n124) );
  XNOR U168 ( .A(n243), .B(n242), .Z(n125) );
  XNOR U169 ( .A(n124), .B(n125), .Z(n126) );
  AND U170 ( .A(n266), .B(n265), .Z(n127) );
  NAND U171 ( .A(n260), .B(n259), .Z(n128) );
  XNOR U172 ( .A(n127), .B(n128), .Z(n129) );
  NAND U173 ( .A(n251), .B(n250), .Z(n130) );
  NAND U174 ( .A(n254), .B(n130), .Z(n131) );
  XNOR U175 ( .A(n129), .B(n131), .Z(n132) );
  XNOR U176 ( .A(n123), .B(n126), .Z(n133) );
  XNOR U177 ( .A(n132), .B(n133), .Z(n134) );
  NANDN U178 ( .A(n219), .B(n220), .Z(n135) );
  XNOR U179 ( .A(n219), .B(n220), .Z(n136) );
  NAND U180 ( .A(n221), .B(n136), .Z(n137) );
  AND U181 ( .A(n135), .B(n137), .Z(n138) );
  XNOR U182 ( .A(n134), .B(n138), .Z(N16) );
  AND U183 ( .A(x[16]), .B(y[48]), .Z(n139) );
  XOR U184 ( .A(n139), .B(o[0]), .Z(N9) );
  AND U185 ( .A(x[16]), .B(y[49]), .Z(n146) );
  XOR U186 ( .A(n146), .B(o[1]), .Z(n141) );
  NAND U187 ( .A(x[17]), .B(y[48]), .Z(n140) );
  XNOR U188 ( .A(n141), .B(n140), .Z(n143) );
  NAND U189 ( .A(n139), .B(o[0]), .Z(n142) );
  XNOR U190 ( .A(n143), .B(n142), .Z(N10) );
  NANDN U191 ( .A(n141), .B(n140), .Z(n145) );
  NAND U192 ( .A(n143), .B(n142), .Z(n144) );
  AND U193 ( .A(n145), .B(n144), .Z(n152) );
  AND U194 ( .A(x[16]), .B(y[50]), .Z(n157) );
  XNOR U195 ( .A(n157), .B(o[2]), .Z(n151) );
  XNOR U196 ( .A(n152), .B(n151), .Z(n154) );
  NAND U197 ( .A(y[49]), .B(x[17]), .Z(n149) );
  AND U198 ( .A(n146), .B(o[1]), .Z(n150) );
  AND U199 ( .A(y[48]), .B(x[18]), .Z(n148) );
  XNOR U200 ( .A(n150), .B(n148), .Z(n147) );
  XNOR U201 ( .A(n149), .B(n147), .Z(n153) );
  XNOR U202 ( .A(n154), .B(n153), .Z(N11) );
  NANDN U203 ( .A(n152), .B(n151), .Z(n156) );
  NAND U204 ( .A(n154), .B(n153), .Z(n155) );
  NAND U205 ( .A(n156), .B(n155), .Z(n163) );
  XNOR U206 ( .A(n164), .B(n163), .Z(n166) );
  NAND U207 ( .A(y[48]), .B(x[19]), .Z(n171) );
  AND U208 ( .A(n157), .B(o[2]), .Z(n172) );
  AND U209 ( .A(x[16]), .B(y[51]), .Z(n170) );
  XNOR U210 ( .A(n172), .B(n170), .Z(n158) );
  XNOR U211 ( .A(n171), .B(n158), .Z(n162) );
  NAND U212 ( .A(y[49]), .B(x[18]), .Z(n173) );
  XNOR U213 ( .A(o[3]), .B(n173), .Z(n161) );
  NAND U214 ( .A(x[17]), .B(y[50]), .Z(n160) );
  XOR U215 ( .A(n161), .B(n160), .Z(n159) );
  XNOR U216 ( .A(n162), .B(n159), .Z(n165) );
  XNOR U217 ( .A(n166), .B(n165), .Z(N12) );
  NANDN U218 ( .A(n164), .B(n163), .Z(n168) );
  NAND U219 ( .A(n166), .B(n165), .Z(n167) );
  NAND U220 ( .A(n168), .B(n167), .Z(n179) );
  XNOR U221 ( .A(n180), .B(n179), .Z(n182) );
  NAND U222 ( .A(y[50]), .B(x[18]), .Z(n188) );
  NAND U223 ( .A(y[49]), .B(x[19]), .Z(n191) );
  XNOR U224 ( .A(o[4]), .B(n191), .Z(n190) );
  AND U225 ( .A(x[17]), .B(y[51]), .Z(n189) );
  XNOR U226 ( .A(n190), .B(n189), .Z(n169) );
  XNOR U227 ( .A(n188), .B(n169), .Z(n176) );
  NAND U228 ( .A(y[48]), .B(x[20]), .Z(n186) );
  ANDN U229 ( .B(o[3]), .A(n173), .Z(n185) );
  NAND U230 ( .A(x[16]), .B(y[52]), .Z(n187) );
  XOR U231 ( .A(n185), .B(n187), .Z(n174) );
  XOR U232 ( .A(n186), .B(n174), .Z(n177) );
  XNOR U233 ( .A(n178), .B(n177), .Z(n175) );
  XNOR U234 ( .A(n176), .B(n175), .Z(n181) );
  XNOR U235 ( .A(n182), .B(n181), .Z(N13) );
  NANDN U236 ( .A(n180), .B(n179), .Z(n184) );
  NAND U237 ( .A(n182), .B(n181), .Z(n183) );
  NAND U238 ( .A(n184), .B(n183), .Z(n195) );
  XNOR U239 ( .A(n196), .B(n195), .Z(n198) );
  XNOR U240 ( .A(n201), .B(n202), .Z(n204) );
  NAND U241 ( .A(y[48]), .B(x[21]), .Z(n216) );
  ANDN U242 ( .B(o[4]), .A(n191), .Z(n217) );
  AND U243 ( .A(x[16]), .B(y[53]), .Z(n215) );
  XNOR U244 ( .A(n217), .B(n215), .Z(n192) );
  XOR U245 ( .A(n216), .B(n192), .Z(n209) );
  NAND U246 ( .A(x[17]), .B(y[52]), .Z(n210) );
  NAND U247 ( .A(y[49]), .B(x[20]), .Z(n213) );
  XNOR U248 ( .A(o[5]), .B(n213), .Z(n212) );
  AND U249 ( .A(y[50]), .B(x[19]), .Z(n211) );
  XNOR U250 ( .A(n212), .B(n211), .Z(n193) );
  XOR U251 ( .A(n210), .B(n193), .Z(n208) );
  NAND U252 ( .A(x[18]), .B(y[51]), .Z(n207) );
  XOR U253 ( .A(n208), .B(n207), .Z(n194) );
  XOR U254 ( .A(n209), .B(n194), .Z(n203) );
  XOR U255 ( .A(n204), .B(n203), .Z(n197) );
  XNOR U256 ( .A(n198), .B(n197), .Z(N14) );
  NANDN U257 ( .A(n196), .B(n195), .Z(n200) );
  NAND U258 ( .A(n198), .B(n197), .Z(n199) );
  NAND U259 ( .A(n200), .B(n199), .Z(n264) );
  NANDN U260 ( .A(n202), .B(n201), .Z(n206) );
  NAND U261 ( .A(n204), .B(n203), .Z(n205) );
  NAND U262 ( .A(n206), .B(n205), .Z(n263) );
  XOR U263 ( .A(n258), .B(n257), .Z(n256) );
  NAND U264 ( .A(y[48]), .B(x[22]), .Z(n245) );
  ANDN U265 ( .B(o[5]), .A(n213), .Z(n244) );
  NAND U266 ( .A(x[16]), .B(y[54]), .Z(n247) );
  XOR U267 ( .A(n244), .B(n247), .Z(n214) );
  XNOR U268 ( .A(n245), .B(n214), .Z(n219) );
  AND U269 ( .A(x[18]), .B(y[52]), .Z(n225) );
  AND U270 ( .A(y[51]), .B(x[19]), .Z(n224) );
  XOR U271 ( .A(n225), .B(n224), .Z(n222) );
  AND U272 ( .A(y[49]), .B(x[21]), .Z(n226) );
  XOR U273 ( .A(n226), .B(o[6]), .Z(n250) );
  NAND U274 ( .A(x[17]), .B(y[53]), .Z(n253) );
  AND U275 ( .A(y[50]), .B(x[20]), .Z(n251) );
  XNOR U276 ( .A(n221), .B(n220), .Z(n218) );
  XOR U277 ( .A(n219), .B(n218), .Z(n255) );
  XNOR U278 ( .A(n256), .B(n255), .Z(n261) );
  XNOR U279 ( .A(n262), .B(n261), .Z(N15) );
  AND U280 ( .A(x[23]), .B(y[48]), .Z(n235) );
  AND U281 ( .A(n226), .B(o[6]), .Z(n233) );
  AND U282 ( .A(x[20]), .B(y[51]), .Z(n231) );
  AND U283 ( .A(y[52]), .B(x[19]), .Z(n228) );
  NAND U284 ( .A(y[53]), .B(x[18]), .Z(n227) );
  XNOR U285 ( .A(n228), .B(n227), .Z(n229) );
  XNOR U286 ( .A(o[7]), .B(n229), .Z(n230) );
  XNOR U287 ( .A(n231), .B(n230), .Z(n232) );
  XNOR U288 ( .A(n233), .B(n232), .Z(n234) );
  XNOR U289 ( .A(n235), .B(n234), .Z(n243) );
  AND U290 ( .A(x[21]), .B(y[50]), .Z(n237) );
  NAND U291 ( .A(x[22]), .B(y[49]), .Z(n236) );
  XNOR U292 ( .A(n237), .B(n236), .Z(n241) );
  AND U293 ( .A(y[54]), .B(x[17]), .Z(n239) );
  NAND U294 ( .A(y[55]), .B(x[16]), .Z(n238) );
  XNOR U295 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U296 ( .A(n241), .B(n240), .Z(n242) );
  NANDN U297 ( .A(n245), .B(n244), .Z(n249) );
  ANDN U298 ( .B(n245), .A(n244), .Z(n246) );
  OR U299 ( .A(n247), .B(n246), .Z(n248) );
  NOR U300 ( .A(n251), .B(n250), .Z(n252) );
  OR U301 ( .A(n253), .B(n252), .Z(n254) );
  OR U302 ( .A(n258), .B(n257), .Z(n259) );
  NAND U303 ( .A(n262), .B(n261), .Z(n266) );
  NAND U304 ( .A(n264), .B(n263), .Z(n265) );
  AND U305 ( .A(x[16]), .B(y[56]), .Z(n267) );
  XOR U306 ( .A(n267), .B(o[8]), .Z(N25) );
  AND U307 ( .A(x[16]), .B(y[57]), .Z(n274) );
  XOR U308 ( .A(n274), .B(o[9]), .Z(n269) );
  NAND U309 ( .A(x[17]), .B(y[56]), .Z(n268) );
  XNOR U310 ( .A(n269), .B(n268), .Z(n271) );
  NAND U311 ( .A(n267), .B(o[8]), .Z(n270) );
  XNOR U312 ( .A(n271), .B(n270), .Z(N26) );
  NANDN U313 ( .A(n269), .B(n268), .Z(n273) );
  NAND U314 ( .A(n271), .B(n270), .Z(n272) );
  AND U315 ( .A(n273), .B(n272), .Z(n280) );
  AND U316 ( .A(x[16]), .B(y[58]), .Z(n285) );
  XNOR U317 ( .A(n285), .B(o[10]), .Z(n279) );
  XNOR U318 ( .A(n280), .B(n279), .Z(n282) );
  NAND U319 ( .A(x[17]), .B(y[57]), .Z(n277) );
  AND U320 ( .A(n274), .B(o[9]), .Z(n278) );
  AND U321 ( .A(x[18]), .B(y[56]), .Z(n276) );
  XNOR U322 ( .A(n278), .B(n276), .Z(n275) );
  XNOR U323 ( .A(n277), .B(n275), .Z(n281) );
  XNOR U324 ( .A(n282), .B(n281), .Z(N27) );
  NANDN U325 ( .A(n280), .B(n279), .Z(n284) );
  NAND U326 ( .A(n282), .B(n281), .Z(n283) );
  NAND U327 ( .A(n284), .B(n283), .Z(n291) );
  XNOR U328 ( .A(n292), .B(n291), .Z(n294) );
  NAND U329 ( .A(x[19]), .B(y[56]), .Z(n299) );
  AND U330 ( .A(n285), .B(o[10]), .Z(n300) );
  AND U331 ( .A(x[16]), .B(y[59]), .Z(n298) );
  XNOR U332 ( .A(n300), .B(n298), .Z(n286) );
  XNOR U333 ( .A(n299), .B(n286), .Z(n290) );
  NAND U334 ( .A(x[18]), .B(y[57]), .Z(n301) );
  XNOR U335 ( .A(o[11]), .B(n301), .Z(n289) );
  NAND U336 ( .A(x[17]), .B(y[58]), .Z(n288) );
  XOR U337 ( .A(n289), .B(n288), .Z(n287) );
  XNOR U338 ( .A(n290), .B(n287), .Z(n293) );
  XNOR U339 ( .A(n294), .B(n293), .Z(N28) );
  NANDN U340 ( .A(n292), .B(n291), .Z(n296) );
  NAND U341 ( .A(n294), .B(n293), .Z(n295) );
  NAND U342 ( .A(n296), .B(n295), .Z(n307) );
  XNOR U343 ( .A(n308), .B(n307), .Z(n310) );
  NAND U344 ( .A(x[18]), .B(y[58]), .Z(n316) );
  NAND U345 ( .A(x[19]), .B(y[57]), .Z(n319) );
  XNOR U346 ( .A(o[12]), .B(n319), .Z(n318) );
  AND U347 ( .A(x[17]), .B(y[59]), .Z(n317) );
  XNOR U348 ( .A(n318), .B(n317), .Z(n297) );
  XNOR U349 ( .A(n316), .B(n297), .Z(n304) );
  NAND U350 ( .A(x[20]), .B(y[56]), .Z(n314) );
  ANDN U351 ( .B(o[11]), .A(n301), .Z(n313) );
  NAND U352 ( .A(x[16]), .B(y[60]), .Z(n315) );
  XOR U353 ( .A(n313), .B(n315), .Z(n302) );
  XOR U354 ( .A(n314), .B(n302), .Z(n305) );
  XNOR U355 ( .A(n306), .B(n305), .Z(n303) );
  XNOR U356 ( .A(n304), .B(n303), .Z(n309) );
  XNOR U357 ( .A(n310), .B(n309), .Z(N29) );
  NANDN U358 ( .A(n308), .B(n307), .Z(n312) );
  NAND U359 ( .A(n310), .B(n309), .Z(n311) );
  NAND U360 ( .A(n312), .B(n311), .Z(n323) );
  XNOR U361 ( .A(n324), .B(n323), .Z(n326) );
  XNOR U362 ( .A(n329), .B(n330), .Z(n332) );
  NAND U363 ( .A(x[21]), .B(y[56]), .Z(n344) );
  ANDN U364 ( .B(o[12]), .A(n319), .Z(n345) );
  AND U365 ( .A(x[16]), .B(y[61]), .Z(n343) );
  XNOR U366 ( .A(n345), .B(n343), .Z(n320) );
  XOR U367 ( .A(n344), .B(n320), .Z(n337) );
  NAND U368 ( .A(x[17]), .B(y[60]), .Z(n338) );
  NAND U369 ( .A(x[20]), .B(y[57]), .Z(n341) );
  XNOR U370 ( .A(o[13]), .B(n341), .Z(n340) );
  AND U371 ( .A(x[19]), .B(y[58]), .Z(n339) );
  XNOR U372 ( .A(n340), .B(n339), .Z(n321) );
  XOR U373 ( .A(n338), .B(n321), .Z(n336) );
  NAND U374 ( .A(x[18]), .B(y[59]), .Z(n335) );
  XOR U375 ( .A(n336), .B(n335), .Z(n322) );
  XOR U376 ( .A(n337), .B(n322), .Z(n331) );
  XOR U377 ( .A(n332), .B(n331), .Z(n325) );
  XNOR U378 ( .A(n326), .B(n325), .Z(N30) );
  NANDN U379 ( .A(n324), .B(n323), .Z(n328) );
  NAND U380 ( .A(n326), .B(n325), .Z(n327) );
  NAND U381 ( .A(n328), .B(n327), .Z(n392) );
  NANDN U382 ( .A(n330), .B(n329), .Z(n334) );
  NAND U383 ( .A(n332), .B(n331), .Z(n333) );
  NAND U384 ( .A(n334), .B(n333), .Z(n391) );
  XOR U385 ( .A(n386), .B(n385), .Z(n384) );
  NAND U386 ( .A(x[22]), .B(y[56]), .Z(n373) );
  ANDN U387 ( .B(o[13]), .A(n341), .Z(n372) );
  NAND U388 ( .A(x[16]), .B(y[62]), .Z(n375) );
  XOR U389 ( .A(n372), .B(n375), .Z(n342) );
  XNOR U390 ( .A(n373), .B(n342), .Z(n347) );
  AND U391 ( .A(x[18]), .B(y[60]), .Z(n353) );
  AND U392 ( .A(x[19]), .B(y[59]), .Z(n352) );
  XOR U393 ( .A(n353), .B(n352), .Z(n350) );
  AND U394 ( .A(x[21]), .B(y[57]), .Z(n354) );
  XOR U395 ( .A(n354), .B(o[14]), .Z(n378) );
  NAND U396 ( .A(x[17]), .B(y[61]), .Z(n381) );
  AND U397 ( .A(x[20]), .B(y[58]), .Z(n379) );
  XNOR U398 ( .A(n349), .B(n348), .Z(n346) );
  XOR U399 ( .A(n347), .B(n346), .Z(n383) );
  XNOR U400 ( .A(n384), .B(n383), .Z(n389) );
  XNOR U401 ( .A(n390), .B(n389), .Z(N31) );
  AND U402 ( .A(y[63]), .B(x[16]), .Z(n363) );
  AND U403 ( .A(n354), .B(o[14]), .Z(n361) );
  AND U404 ( .A(y[59]), .B(x[20]), .Z(n359) );
  AND U405 ( .A(y[60]), .B(x[19]), .Z(n356) );
  NAND U406 ( .A(y[61]), .B(x[18]), .Z(n355) );
  XNOR U407 ( .A(n356), .B(n355), .Z(n357) );
  XNOR U408 ( .A(o[15]), .B(n357), .Z(n358) );
  XNOR U409 ( .A(n359), .B(n358), .Z(n360) );
  XNOR U410 ( .A(n361), .B(n360), .Z(n362) );
  XNOR U411 ( .A(n363), .B(n362), .Z(n371) );
  AND U412 ( .A(y[57]), .B(x[22]), .Z(n365) );
  NAND U413 ( .A(y[58]), .B(x[21]), .Z(n364) );
  XNOR U414 ( .A(n365), .B(n364), .Z(n369) );
  AND U415 ( .A(y[56]), .B(x[23]), .Z(n367) );
  NAND U416 ( .A(y[62]), .B(x[17]), .Z(n366) );
  XNOR U417 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U418 ( .A(n369), .B(n368), .Z(n370) );
  NANDN U419 ( .A(n373), .B(n372), .Z(n377) );
  ANDN U420 ( .B(n373), .A(n372), .Z(n374) );
  OR U421 ( .A(n375), .B(n374), .Z(n376) );
  NOR U422 ( .A(n379), .B(n378), .Z(n380) );
  OR U423 ( .A(n381), .B(n380), .Z(n382) );
  OR U424 ( .A(n386), .B(n385), .Z(n387) );
  NAND U425 ( .A(n390), .B(n389), .Z(n394) );
  NAND U426 ( .A(n392), .B(n391), .Z(n393) );
  AND U427 ( .A(x[16]), .B(y[64]), .Z(n395) );
  XOR U428 ( .A(n395), .B(o[16]), .Z(N41) );
  AND U429 ( .A(x[16]), .B(y[65]), .Z(n402) );
  XOR U430 ( .A(n402), .B(o[17]), .Z(n397) );
  NAND U431 ( .A(x[17]), .B(y[64]), .Z(n396) );
  XNOR U432 ( .A(n397), .B(n396), .Z(n399) );
  NAND U433 ( .A(n395), .B(o[16]), .Z(n398) );
  XNOR U434 ( .A(n399), .B(n398), .Z(N42) );
  NANDN U435 ( .A(n397), .B(n396), .Z(n401) );
  NAND U436 ( .A(n399), .B(n398), .Z(n400) );
  AND U437 ( .A(n401), .B(n400), .Z(n408) );
  AND U438 ( .A(x[16]), .B(y[66]), .Z(n413) );
  XNOR U439 ( .A(n413), .B(o[18]), .Z(n407) );
  XNOR U440 ( .A(n408), .B(n407), .Z(n410) );
  NAND U441 ( .A(x[17]), .B(y[65]), .Z(n405) );
  AND U442 ( .A(n402), .B(o[17]), .Z(n406) );
  AND U443 ( .A(x[18]), .B(y[64]), .Z(n404) );
  XNOR U444 ( .A(n406), .B(n404), .Z(n403) );
  XNOR U445 ( .A(n405), .B(n403), .Z(n409) );
  XNOR U446 ( .A(n410), .B(n409), .Z(N43) );
  NANDN U447 ( .A(n408), .B(n407), .Z(n412) );
  NAND U448 ( .A(n410), .B(n409), .Z(n411) );
  NAND U449 ( .A(n412), .B(n411), .Z(n419) );
  XNOR U450 ( .A(n420), .B(n419), .Z(n422) );
  NAND U451 ( .A(x[19]), .B(y[64]), .Z(n427) );
  AND U452 ( .A(n413), .B(o[18]), .Z(n428) );
  AND U453 ( .A(x[16]), .B(y[67]), .Z(n426) );
  XNOR U454 ( .A(n428), .B(n426), .Z(n414) );
  XNOR U455 ( .A(n427), .B(n414), .Z(n418) );
  NAND U456 ( .A(x[18]), .B(y[65]), .Z(n429) );
  XNOR U457 ( .A(o[19]), .B(n429), .Z(n417) );
  NAND U458 ( .A(x[17]), .B(y[66]), .Z(n416) );
  XOR U459 ( .A(n417), .B(n416), .Z(n415) );
  XNOR U460 ( .A(n418), .B(n415), .Z(n421) );
  XNOR U461 ( .A(n422), .B(n421), .Z(N44) );
  NANDN U462 ( .A(n420), .B(n419), .Z(n424) );
  NAND U463 ( .A(n422), .B(n421), .Z(n423) );
  NAND U464 ( .A(n424), .B(n423), .Z(n435) );
  XNOR U465 ( .A(n436), .B(n435), .Z(n438) );
  NAND U466 ( .A(x[18]), .B(y[66]), .Z(n444) );
  NAND U467 ( .A(x[19]), .B(y[65]), .Z(n447) );
  XNOR U468 ( .A(o[20]), .B(n447), .Z(n446) );
  AND U469 ( .A(x[17]), .B(y[67]), .Z(n445) );
  XNOR U470 ( .A(n446), .B(n445), .Z(n425) );
  XNOR U471 ( .A(n444), .B(n425), .Z(n432) );
  NAND U472 ( .A(x[20]), .B(y[64]), .Z(n442) );
  ANDN U473 ( .B(o[19]), .A(n429), .Z(n441) );
  NAND U474 ( .A(x[16]), .B(y[68]), .Z(n443) );
  XOR U475 ( .A(n441), .B(n443), .Z(n430) );
  XOR U476 ( .A(n442), .B(n430), .Z(n433) );
  XNOR U477 ( .A(n434), .B(n433), .Z(n431) );
  XNOR U478 ( .A(n432), .B(n431), .Z(n437) );
  XNOR U479 ( .A(n438), .B(n437), .Z(N45) );
  NANDN U480 ( .A(n436), .B(n435), .Z(n440) );
  NAND U481 ( .A(n438), .B(n437), .Z(n439) );
  NAND U482 ( .A(n440), .B(n439), .Z(n451) );
  XNOR U483 ( .A(n452), .B(n451), .Z(n454) );
  XNOR U484 ( .A(n457), .B(n458), .Z(n460) );
  NAND U485 ( .A(x[21]), .B(y[64]), .Z(n472) );
  ANDN U486 ( .B(o[20]), .A(n447), .Z(n473) );
  AND U487 ( .A(x[16]), .B(y[69]), .Z(n471) );
  XNOR U488 ( .A(n473), .B(n471), .Z(n448) );
  XOR U489 ( .A(n472), .B(n448), .Z(n465) );
  NAND U490 ( .A(x[17]), .B(y[68]), .Z(n466) );
  NAND U491 ( .A(x[20]), .B(y[65]), .Z(n469) );
  XNOR U492 ( .A(o[21]), .B(n469), .Z(n468) );
  AND U493 ( .A(x[19]), .B(y[66]), .Z(n467) );
  XNOR U494 ( .A(n468), .B(n467), .Z(n449) );
  XOR U495 ( .A(n466), .B(n449), .Z(n464) );
  NAND U496 ( .A(x[18]), .B(y[67]), .Z(n463) );
  XOR U497 ( .A(n464), .B(n463), .Z(n450) );
  XOR U498 ( .A(n465), .B(n450), .Z(n459) );
  XOR U499 ( .A(n460), .B(n459), .Z(n453) );
  XNOR U500 ( .A(n454), .B(n453), .Z(N46) );
  NANDN U501 ( .A(n452), .B(n451), .Z(n456) );
  NAND U502 ( .A(n454), .B(n453), .Z(n455) );
  NAND U503 ( .A(n456), .B(n455), .Z(n520) );
  NANDN U504 ( .A(n458), .B(n457), .Z(n462) );
  NAND U505 ( .A(n460), .B(n459), .Z(n461) );
  NAND U506 ( .A(n462), .B(n461), .Z(n519) );
  XOR U507 ( .A(n514), .B(n513), .Z(n512) );
  NAND U508 ( .A(x[22]), .B(y[64]), .Z(n501) );
  ANDN U509 ( .B(o[21]), .A(n469), .Z(n500) );
  NAND U510 ( .A(x[16]), .B(y[70]), .Z(n503) );
  XOR U511 ( .A(n500), .B(n503), .Z(n470) );
  XNOR U512 ( .A(n501), .B(n470), .Z(n475) );
  AND U513 ( .A(x[18]), .B(y[68]), .Z(n481) );
  AND U514 ( .A(x[19]), .B(y[67]), .Z(n480) );
  XOR U515 ( .A(n481), .B(n480), .Z(n478) );
  AND U516 ( .A(x[21]), .B(y[65]), .Z(n482) );
  XOR U517 ( .A(n482), .B(o[22]), .Z(n506) );
  NAND U518 ( .A(x[17]), .B(y[69]), .Z(n509) );
  AND U519 ( .A(x[20]), .B(y[66]), .Z(n507) );
  XNOR U520 ( .A(n477), .B(n476), .Z(n474) );
  XOR U521 ( .A(n475), .B(n474), .Z(n511) );
  XNOR U522 ( .A(n512), .B(n511), .Z(n517) );
  XNOR U523 ( .A(n518), .B(n517), .Z(N47) );
  AND U524 ( .A(y[71]), .B(x[16]), .Z(n491) );
  AND U525 ( .A(n482), .B(o[22]), .Z(n489) );
  AND U526 ( .A(y[67]), .B(x[20]), .Z(n487) );
  AND U527 ( .A(y[68]), .B(x[19]), .Z(n484) );
  NAND U528 ( .A(y[69]), .B(x[18]), .Z(n483) );
  XNOR U529 ( .A(n484), .B(n483), .Z(n485) );
  XNOR U530 ( .A(o[23]), .B(n485), .Z(n486) );
  XNOR U531 ( .A(n487), .B(n486), .Z(n488) );
  XNOR U532 ( .A(n489), .B(n488), .Z(n490) );
  XNOR U533 ( .A(n491), .B(n490), .Z(n499) );
  AND U534 ( .A(y[65]), .B(x[22]), .Z(n493) );
  NAND U535 ( .A(y[66]), .B(x[21]), .Z(n492) );
  XNOR U536 ( .A(n493), .B(n492), .Z(n497) );
  AND U537 ( .A(y[64]), .B(x[23]), .Z(n495) );
  NAND U538 ( .A(y[70]), .B(x[17]), .Z(n494) );
  XNOR U539 ( .A(n495), .B(n494), .Z(n496) );
  XNOR U540 ( .A(n497), .B(n496), .Z(n498) );
  NANDN U541 ( .A(n501), .B(n500), .Z(n505) );
  ANDN U542 ( .B(n501), .A(n500), .Z(n502) );
  OR U543 ( .A(n503), .B(n502), .Z(n504) );
  NOR U544 ( .A(n507), .B(n506), .Z(n508) );
  OR U545 ( .A(n509), .B(n508), .Z(n510) );
  OR U546 ( .A(n514), .B(n513), .Z(n515) );
  NAND U547 ( .A(n518), .B(n517), .Z(n522) );
  NAND U548 ( .A(n520), .B(n519), .Z(n521) );
endmodule

