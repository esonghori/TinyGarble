
module modexp_2N_NN_N4_CC16 ( clk, rst, m, e, n, c );
  input [3:0] m;
  input [3:0] e;
  input [3:0] n;
  output [3:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, \modmult_1/xreg[3] , \modmult_1/xreg[2] ,
         \modmult_1/xin[1] , \modmult_1/xin[0] , \modmult_1/zreg[4] ,
         \modmult_1/zreg[3] , \modmult_1/zreg[2] , \modmult_1/zreg[1] ,
         \modmult_1/zreg[0] , \modmult_1/zout[1][4] , n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392;
  wire   [1:0] start_in;
  wire   [1:0] start_reg;
  wire   [3:0] ereg;
  wire   [3:0] o;
  wire   [3:0] creg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \modmult_1/xreg_reg[2]  ( .D(\modmult_1/xin[0] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[2] ) );
  DFF \modmult_1/xreg_reg[3]  ( .D(\modmult_1/xin[1] ), .CLK(clk), .RST(rst), 
        .Q(\modmult_1/xreg[3] ) );
  DFF \modmult_1/zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[0] ) );
  DFF \modmult_1/zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[1] ) );
  DFF \modmult_1/zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[2] ) );
  DFF \modmult_1/zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(
        \modmult_1/zreg[3] ) );
  DFF \modmult_1/zreg_reg[4]  ( .D(\modmult_1/zout[1][4] ), .CLK(clk), .RST(
        rst), .Q(\modmult_1/zreg[4] ) );
  DFF mul_pow_reg ( .D(n47), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n46), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n45), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n44), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n43), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF first_one_reg ( .D(n42), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n41), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n40), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n39), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n38), .CLK(clk), .RST(rst), .Q(creg[3]) );
  NANDN U172 ( .A(n246), .B(n247), .Z(n129) );
  NANDN U173 ( .A(n259), .B(n260), .Z(n130) );
  AND U174 ( .A(n129), .B(n130), .Z(n131) );
  NAND U175 ( .A(n281), .B(n280), .Z(n132) );
  XNOR U176 ( .A(n279), .B(n132), .Z(n133) );
  XNOR U177 ( .A(n131), .B(n133), .Z(n321) );
  NAND U178 ( .A(n313), .B(n[1]), .Z(n134) );
  XOR U179 ( .A(n313), .B(n[1]), .Z(n135) );
  NAND U180 ( .A(n135), .B(n310), .Z(n136) );
  NAND U181 ( .A(n134), .B(n136), .Z(n316) );
  ANDN U182 ( .B(n292), .A(n211), .Z(n206) );
  NAND U183 ( .A(n239), .B(n[1]), .Z(n137) );
  XOR U184 ( .A(n239), .B(n[1]), .Z(n138) );
  NAND U185 ( .A(n138), .B(n221), .Z(n139) );
  NAND U186 ( .A(n137), .B(n139), .Z(n235) );
  OR U187 ( .A(n[1]), .B(n313), .Z(n140) );
  NANDN U188 ( .A(n297), .B(n140), .Z(n141) );
  NAND U189 ( .A(n298), .B(n141), .Z(n142) );
  NOR U190 ( .A(n321), .B(n305), .Z(n143) );
  OR U191 ( .A(n142), .B(n302), .Z(n144) );
  AND U192 ( .A(n143), .B(n144), .Z(n145) );
  NANDN U193 ( .A(n300), .B(n145), .Z(n318) );
  NANDN U194 ( .A(n270), .B(n[0]), .Z(n146) );
  NANDN U195 ( .A(n[1]), .B(n249), .Z(n147) );
  XNOR U196 ( .A(n[1]), .B(n249), .Z(n148) );
  NAND U197 ( .A(n148), .B(n146), .Z(n149) );
  NAND U198 ( .A(n147), .B(n149), .Z(n150) );
  NAND U199 ( .A(n150), .B(n255), .Z(n151) );
  XOR U200 ( .A(n150), .B(n255), .Z(n152) );
  NANDN U201 ( .A(n[2]), .B(n152), .Z(n153) );
  NAND U202 ( .A(n151), .B(n153), .Z(n154) );
  NANDN U203 ( .A(n247), .B(n[3]), .Z(n155) );
  NAND U204 ( .A(n154), .B(n155), .Z(n156) );
  NAND U205 ( .A(n253), .B(n156), .Z(n254) );
  AND U206 ( .A(n[0]), .B(n322), .Z(n157) );
  XOR U207 ( .A(n[1]), .B(n327), .Z(n158) );
  NAND U208 ( .A(n158), .B(n157), .Z(n159) );
  NAND U209 ( .A(n[1]), .B(n327), .Z(n160) );
  AND U210 ( .A(n159), .B(n160), .Z(n161) );
  XOR U211 ( .A(n331), .B(n161), .Z(n162) );
  NANDN U212 ( .A(n[2]), .B(n162), .Z(n163) );
  NAND U213 ( .A(n331), .B(n161), .Z(n164) );
  AND U214 ( .A(n163), .B(n164), .Z(n165) );
  NANDN U215 ( .A(n333), .B(n165), .Z(n166) );
  XNOR U216 ( .A(n333), .B(n165), .Z(n167) );
  NAND U217 ( .A(n167), .B(n[3]), .Z(n168) );
  NAND U218 ( .A(n166), .B(n168), .Z(n169) );
  AND U219 ( .A(n340), .B(n169), .Z(n170) );
  NANDN U220 ( .A(n321), .B(n170), .Z(n332) );
  NAND U221 ( .A(n254), .B(n[2]), .Z(n171) );
  AND U222 ( .A(n255), .B(n171), .Z(n257) );
  NAND U223 ( .A(n329), .B(n331), .Z(n172) );
  XOR U224 ( .A(n329), .B(n331), .Z(n173) );
  NAND U225 ( .A(n173), .B(n330), .Z(n174) );
  NAND U226 ( .A(n172), .B(n174), .Z(n334) );
  ANDN U227 ( .B(n[0]), .A(n245), .Z(n239) );
  OR U228 ( .A(n228), .B(n229), .Z(n175) );
  AND U229 ( .A(n230), .B(n175), .Z(n176) );
  XNOR U230 ( .A(n231), .B(n176), .Z(n177) );
  OR U231 ( .A(n176), .B(n243), .Z(n178) );
  NAND U232 ( .A(n177), .B(n178), .Z(n279) );
  ANDN U233 ( .B(n292), .A(n294), .Z(n287) );
  NAND U234 ( .A(n359), .B(start_reg[1]), .Z(n179) );
  AND U235 ( .A(init), .B(n179), .Z(n372) );
  XOR U236 ( .A(n327), .B(n325), .Z(n180) );
  NANDN U237 ( .A(n326), .B(n180), .Z(n181) );
  NAND U238 ( .A(n327), .B(n325), .Z(n182) );
  AND U239 ( .A(n181), .B(n182), .Z(n330) );
  NANDN U240 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  ANDN U241 ( .B(\modmult_1/zreg[2] ), .A(start_in[0]), .Z(n197) );
  NAND U242 ( .A(init), .B(start_reg[0]), .Z(n351) );
  NANDN U243 ( .A(n351), .B(creg[3]), .Z(n184) );
  NANDN U244 ( .A(start_in[0]), .B(\modmult_1/xreg[3] ), .Z(n183) );
  NAND U245 ( .A(n184), .B(n183), .Z(n185) );
  NANDN U246 ( .A(init), .B(m[3]), .Z(n362) );
  NANDN U247 ( .A(n185), .B(n362), .Z(n220) );
  ANDN U248 ( .B(init), .A(mul_pow), .Z(n353) );
  NANDN U249 ( .A(creg[3]), .B(n353), .Z(n187) );
  OR U250 ( .A(n353), .B(m[3]), .Z(n186) );
  NAND U251 ( .A(n187), .B(n186), .Z(n283) );
  IV U252 ( .A(n283), .Z(n266) );
  NAND U253 ( .A(creg[2]), .B(n353), .Z(n189) );
  NANDN U254 ( .A(n353), .B(m[2]), .Z(n188) );
  NAND U255 ( .A(n189), .B(n188), .Z(n288) );
  NAND U256 ( .A(creg[1]), .B(n353), .Z(n191) );
  NANDN U257 ( .A(n353), .B(m[1]), .Z(n190) );
  NAND U258 ( .A(n191), .B(n190), .Z(n292) );
  NANDN U259 ( .A(start_in[0]), .B(\modmult_1/zreg[0] ), .Z(n211) );
  NAND U260 ( .A(n288), .B(n206), .Z(n194) );
  ANDN U261 ( .B(\modmult_1/zreg[1] ), .A(start_in[0]), .Z(n209) );
  IV U262 ( .A(n288), .Z(n271) );
  NANDN U263 ( .A(n206), .B(n271), .Z(n192) );
  NAND U264 ( .A(n209), .B(n192), .Z(n193) );
  NAND U265 ( .A(n194), .B(n193), .Z(n196) );
  XOR U266 ( .A(n266), .B(n196), .Z(n198) );
  NAND U267 ( .A(n220), .B(n198), .Z(n195) );
  XNOR U268 ( .A(n197), .B(n195), .Z(n227) );
  NAND U269 ( .A(n266), .B(n196), .Z(n200) );
  NAND U270 ( .A(n198), .B(n197), .Z(n199) );
  NAND U271 ( .A(n200), .B(n199), .Z(n201) );
  AND U272 ( .A(n220), .B(n201), .Z(n205) );
  ANDN U273 ( .B(\modmult_1/zreg[3] ), .A(start_in[0]), .Z(n204) );
  NAND U274 ( .A(n205), .B(n204), .Z(n203) );
  NANDN U275 ( .A(start_in[0]), .B(\modmult_1/zreg[4] ), .Z(n202) );
  XOR U276 ( .A(n203), .B(n202), .Z(n232) );
  ANDN U277 ( .B(n227), .A(n[3]), .Z(n229) );
  XOR U278 ( .A(n205), .B(n204), .Z(n231) );
  NOR U279 ( .A(n229), .B(n231), .Z(n216) );
  XOR U280 ( .A(n288), .B(n206), .Z(n207) );
  NAND U281 ( .A(n220), .B(n207), .Z(n208) );
  XNOR U282 ( .A(n209), .B(n208), .Z(n238) );
  NANDN U283 ( .A(n238), .B(n[2]), .Z(n224) );
  ANDN U284 ( .B(n238), .A(n[2]), .Z(n222) );
  NAND U285 ( .A(n292), .B(n220), .Z(n210) );
  XOR U286 ( .A(n211), .B(n210), .Z(n242) );
  IV U287 ( .A(n242), .Z(n221) );
  OR U288 ( .A(n[1]), .B(n221), .Z(n212) );
  NANDN U289 ( .A(n222), .B(n212), .Z(n213) );
  NAND U290 ( .A(n224), .B(n213), .Z(n214) );
  NANDN U291 ( .A(n227), .B(n[3]), .Z(n230) );
  NANDN U292 ( .A(n214), .B(n230), .Z(n215) );
  AND U293 ( .A(n216), .B(n215), .Z(n217) );
  NANDN U294 ( .A(n232), .B(n217), .Z(n243) );
  NAND U295 ( .A(creg[0]), .B(n353), .Z(n219) );
  NANDN U296 ( .A(n353), .B(m[0]), .Z(n218) );
  NAND U297 ( .A(n219), .B(n218), .Z(n295) );
  AND U298 ( .A(n220), .B(n295), .Z(n245) );
  NANDN U299 ( .A(n222), .B(n235), .Z(n223) );
  AND U300 ( .A(n224), .B(n223), .Z(n228) );
  XNOR U301 ( .A(n[3]), .B(n228), .Z(n225) );
  NAND U302 ( .A(n243), .B(n225), .Z(n226) );
  XNOR U303 ( .A(n227), .B(n226), .Z(n247) );
  ANDN U304 ( .B(n279), .A(n232), .Z(n234) );
  NANDN U305 ( .A(n[3]), .B(n247), .Z(n233) );
  AND U306 ( .A(n234), .B(n233), .Z(n253) );
  XOR U307 ( .A(n[2]), .B(n235), .Z(n236) );
  AND U308 ( .A(n236), .B(n243), .Z(n237) );
  XOR U309 ( .A(n238), .B(n237), .Z(n255) );
  XOR U310 ( .A(n[1]), .B(n239), .Z(n240) );
  NAND U311 ( .A(n243), .B(n240), .Z(n241) );
  XNOR U312 ( .A(n242), .B(n241), .Z(n249) );
  NAND U313 ( .A(n243), .B(n[0]), .Z(n244) );
  XNOR U314 ( .A(n245), .B(n244), .Z(n270) );
  AND U315 ( .A(n[3]), .B(n254), .Z(n246) );
  XNOR U316 ( .A(n247), .B(n246), .Z(n260) );
  AND U317 ( .A(n[1]), .B(n254), .Z(n248) );
  NANDN U318 ( .A(n248), .B(n249), .Z(n251) );
  AND U319 ( .A(n[0]), .B(n254), .Z(n269) );
  ANDN U320 ( .B(n269), .A(n270), .Z(n268) );
  XNOR U321 ( .A(n249), .B(n248), .Z(n267) );
  NANDN U322 ( .A(n268), .B(n267), .Z(n250) );
  AND U323 ( .A(n251), .B(n250), .Z(n264) );
  NANDN U324 ( .A(n255), .B(n[2]), .Z(n252) );
  OR U325 ( .A(n253), .B(n252), .Z(n256) );
  ANDN U326 ( .B(n256), .A(n257), .Z(n265) );
  NANDN U327 ( .A(n264), .B(n265), .Z(n258) );
  ANDN U328 ( .B(n258), .A(n257), .Z(n259) );
  XNOR U329 ( .A(n260), .B(n259), .Z(n281) );
  NANDN U330 ( .A(n351), .B(creg[2]), .Z(n262) );
  NANDN U331 ( .A(start_in[0]), .B(\modmult_1/xreg[2] ), .Z(n261) );
  NAND U332 ( .A(n262), .B(n261), .Z(n263) );
  NANDN U333 ( .A(init), .B(m[2]), .Z(n366) );
  NANDN U334 ( .A(n263), .B(n366), .Z(n296) );
  XNOR U335 ( .A(n265), .B(n264), .Z(n286) );
  AND U336 ( .A(n286), .B(n266), .Z(n277) );
  XNOR U337 ( .A(n283), .B(n286), .Z(n275) );
  XNOR U338 ( .A(n268), .B(n267), .Z(n291) );
  NAND U339 ( .A(n288), .B(n291), .Z(n274) );
  XNOR U340 ( .A(n270), .B(n269), .Z(n294) );
  XNOR U341 ( .A(n271), .B(n291), .Z(n272) );
  NAND U342 ( .A(n287), .B(n272), .Z(n273) );
  AND U343 ( .A(n274), .B(n273), .Z(n282) );
  ANDN U344 ( .B(n275), .A(n282), .Z(n276) );
  OR U345 ( .A(n277), .B(n276), .Z(n278) );
  AND U346 ( .A(n296), .B(n278), .Z(n280) );
  XOR U347 ( .A(n281), .B(n280), .Z(n305) );
  XOR U348 ( .A(n283), .B(n282), .Z(n284) );
  NAND U349 ( .A(n296), .B(n284), .Z(n285) );
  XNOR U350 ( .A(n286), .B(n285), .Z(n309) );
  ANDN U351 ( .B(n309), .A(n[3]), .Z(n300) );
  XOR U352 ( .A(n288), .B(n287), .Z(n289) );
  NAND U353 ( .A(n296), .B(n289), .Z(n290) );
  XNOR U354 ( .A(n291), .B(n290), .Z(n320) );
  NANDN U355 ( .A(n320), .B(n[2]), .Z(n298) );
  ANDN U356 ( .B(n320), .A(n[2]), .Z(n297) );
  NAND U357 ( .A(n292), .B(n296), .Z(n293) );
  XNOR U358 ( .A(n294), .B(n293), .Z(n313) );
  ANDN U359 ( .B(n[3]), .A(n309), .Z(n302) );
  NAND U360 ( .A(n296), .B(n295), .Z(n315) );
  AND U361 ( .A(n[0]), .B(n315), .Z(n310) );
  NANDN U362 ( .A(n297), .B(n316), .Z(n299) );
  AND U363 ( .A(n299), .B(n298), .Z(n306) );
  OR U364 ( .A(n300), .B(n306), .Z(n301) );
  NANDN U365 ( .A(n302), .B(n301), .Z(n303) );
  AND U366 ( .A(n318), .B(n303), .Z(n304) );
  XNOR U367 ( .A(n305), .B(n304), .Z(n340) );
  XNOR U368 ( .A(n[3]), .B(n306), .Z(n307) );
  NAND U369 ( .A(n318), .B(n307), .Z(n308) );
  XNOR U370 ( .A(n309), .B(n308), .Z(n333) );
  XOR U371 ( .A(n[1]), .B(n310), .Z(n311) );
  NAND U372 ( .A(n318), .B(n311), .Z(n312) );
  XNOR U373 ( .A(n313), .B(n312), .Z(n327) );
  NAND U374 ( .A(n318), .B(n[0]), .Z(n314) );
  XNOR U375 ( .A(n315), .B(n314), .Z(n322) );
  XOR U376 ( .A(n[2]), .B(n316), .Z(n317) );
  NAND U377 ( .A(n318), .B(n317), .Z(n319) );
  XNOR U378 ( .A(n320), .B(n319), .Z(n331) );
  AND U379 ( .A(n[0]), .B(n332), .Z(n323) );
  XNOR U380 ( .A(n323), .B(n322), .Z(o[0]) );
  AND U381 ( .A(n[1]), .B(n332), .Z(n325) );
  NAND U382 ( .A(n323), .B(n322), .Z(n326) );
  XOR U383 ( .A(n327), .B(n326), .Z(n324) );
  XOR U384 ( .A(n325), .B(n324), .Z(o[1]) );
  NAND U385 ( .A(n[2]), .B(n332), .Z(n329) );
  XNOR U386 ( .A(n331), .B(n330), .Z(n328) );
  XNOR U387 ( .A(n329), .B(n328), .Z(o[2]) );
  XOR U388 ( .A(n333), .B(n334), .Z(n335) );
  AND U389 ( .A(n[3]), .B(n332), .Z(n336) );
  XNOR U390 ( .A(n335), .B(n336), .Z(o[3]) );
  OR U391 ( .A(n334), .B(n333), .Z(n338) );
  NAND U392 ( .A(n336), .B(n335), .Z(n337) );
  NAND U393 ( .A(n338), .B(n337), .Z(n339) );
  XNOR U394 ( .A(n340), .B(n339), .Z(\modmult_1/zout[1][4] ) );
  NANDN U395 ( .A(init), .B(e[3]), .Z(n381) );
  NAND U396 ( .A(ereg[3]), .B(init), .Z(n341) );
  AND U397 ( .A(n381), .B(n341), .Z(n357) );
  NAND U398 ( .A(creg[0]), .B(n357), .Z(n343) );
  NANDN U399 ( .A(n357), .B(o[0]), .Z(n342) );
  NAND U400 ( .A(n343), .B(n342), .Z(c[0]) );
  NAND U401 ( .A(creg[1]), .B(n357), .Z(n345) );
  NANDN U402 ( .A(n357), .B(o[1]), .Z(n344) );
  NAND U403 ( .A(n345), .B(n344), .Z(c[1]) );
  NAND U404 ( .A(creg[2]), .B(n357), .Z(n347) );
  NANDN U405 ( .A(n357), .B(o[2]), .Z(n346) );
  NAND U406 ( .A(n347), .B(n346), .Z(c[2]) );
  NAND U407 ( .A(creg[3]), .B(n357), .Z(n349) );
  NANDN U408 ( .A(n357), .B(o[3]), .Z(n348) );
  NAND U409 ( .A(n349), .B(n348), .Z(c[3]) );
  NANDN U410 ( .A(init), .B(m[0]), .Z(n376) );
  NANDN U411 ( .A(n351), .B(creg[0]), .Z(n350) );
  NAND U412 ( .A(n376), .B(n350), .Z(\modmult_1/xin[0] ) );
  NANDN U413 ( .A(init), .B(m[1]), .Z(n370) );
  NANDN U414 ( .A(n351), .B(creg[1]), .Z(n352) );
  NAND U415 ( .A(n370), .B(n352), .Z(\modmult_1/xin[1] ) );
  NANDN U416 ( .A(start_reg[1]), .B(init), .Z(n354) );
  ANDN U417 ( .B(n354), .A(n353), .Z(n387) );
  NANDN U418 ( .A(n387), .B(ereg[0]), .Z(n356) );
  NANDN U419 ( .A(init), .B(e[0]), .Z(n355) );
  NAND U420 ( .A(n356), .B(n355), .Z(n46) );
  NAND U421 ( .A(n357), .B(mul_pow), .Z(n358) );
  AND U422 ( .A(first_one), .B(n358), .Z(n359) );
  NAND U423 ( .A(creg[3]), .B(n372), .Z(n361) );
  AND U424 ( .A(init), .B(start_reg[1]), .Z(start_in[1]) );
  AND U425 ( .A(start_in[1]), .B(n359), .Z(n373) );
  NAND U426 ( .A(n373), .B(o[3]), .Z(n360) );
  AND U427 ( .A(n361), .B(n360), .Z(n363) );
  NAND U428 ( .A(n363), .B(n362), .Z(n38) );
  NAND U429 ( .A(o[2]), .B(n373), .Z(n365) );
  NAND U430 ( .A(n372), .B(creg[2]), .Z(n364) );
  AND U431 ( .A(n365), .B(n364), .Z(n367) );
  NAND U432 ( .A(n367), .B(n366), .Z(n39) );
  NAND U433 ( .A(creg[1]), .B(n372), .Z(n369) );
  NAND U434 ( .A(n373), .B(o[1]), .Z(n368) );
  AND U435 ( .A(n369), .B(n368), .Z(n371) );
  NAND U436 ( .A(n371), .B(n370), .Z(n40) );
  NAND U437 ( .A(creg[0]), .B(n372), .Z(n375) );
  NAND U438 ( .A(n373), .B(o[0]), .Z(n374) );
  AND U439 ( .A(n375), .B(n374), .Z(n377) );
  NAND U440 ( .A(n377), .B(n376), .Z(n41) );
  AND U441 ( .A(mul_pow), .B(start_in[1]), .Z(n390) );
  NAND U442 ( .A(ereg[3]), .B(n390), .Z(n378) );
  NANDN U443 ( .A(first_one), .B(n378), .Z(n42) );
  NAND U444 ( .A(ereg[2]), .B(n390), .Z(n380) );
  NANDN U445 ( .A(n387), .B(ereg[3]), .Z(n379) );
  AND U446 ( .A(n380), .B(n379), .Z(n382) );
  NAND U447 ( .A(n382), .B(n381), .Z(n43) );
  NANDN U448 ( .A(init), .B(e[2]), .Z(n384) );
  NANDN U449 ( .A(n387), .B(ereg[2]), .Z(n383) );
  AND U450 ( .A(n384), .B(n383), .Z(n386) );
  NAND U451 ( .A(n390), .B(ereg[1]), .Z(n385) );
  NAND U452 ( .A(n386), .B(n385), .Z(n44) );
  NANDN U453 ( .A(init), .B(e[1]), .Z(n389) );
  NANDN U454 ( .A(n387), .B(ereg[1]), .Z(n388) );
  AND U455 ( .A(n389), .B(n388), .Z(n392) );
  NAND U456 ( .A(n390), .B(ereg[0]), .Z(n391) );
  NAND U457 ( .A(n392), .B(n391), .Z(n45) );
  XOR U458 ( .A(mul_pow), .B(start_in[1]), .Z(n47) );
endmodule

