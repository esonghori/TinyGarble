
module matrixMult_N_M_3_N8_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014;

  DFF \o_reg[31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \o_reg[30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \o_reg[29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \o_reg[28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \o_reg[27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \o_reg[26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \o_reg[25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \o_reg[24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \o_reg[23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \o_reg[22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \o_reg[21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \o_reg[20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \o_reg[19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \o_reg[18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \o_reg[17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \o_reg[16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \o_reg[15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \o_reg[14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \o_reg[13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \o_reg[12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \o_reg[11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \o_reg[10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \o_reg[9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \o_reg[8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \o_reg[7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \o_reg[6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \o_reg[5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \o_reg[4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \o_reg[3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \o_reg[2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \o_reg[1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \o_reg[0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  XNOR U3 ( .A(n1768), .B(n1767), .Z(n1705) );
  NAND U4 ( .A(n2021), .B(n2020), .Z(n1) );
  NANDN U5 ( .A(n2023), .B(n2022), .Z(n2) );
  AND U6 ( .A(n1), .B(n2), .Z(n2096) );
  XNOR U7 ( .A(n2183), .B(n2182), .Z(n2143) );
  XNOR U8 ( .A(n2353), .B(n2352), .Z(n2355) );
  XNOR U9 ( .A(n2310), .B(n2309), .Z(n2252) );
  XNOR U10 ( .A(n2639), .B(n2638), .Z(n2664) );
  XNOR U11 ( .A(n2724), .B(n2723), .Z(n2722) );
  XNOR U12 ( .A(n1208), .B(n1207), .Z(n1189) );
  XNOR U13 ( .A(n1216), .B(n1215), .Z(n1254) );
  XNOR U14 ( .A(n1590), .B(n1589), .Z(n1557) );
  XNOR U15 ( .A(n1756), .B(n1755), .Z(n1707) );
  OR U16 ( .A(n1960), .B(n1961), .Z(n3) );
  NAND U17 ( .A(n1959), .B(n1958), .Z(n4) );
  AND U18 ( .A(n3), .B(n4), .Z(n2138) );
  NAND U19 ( .A(n2145), .B(n2144), .Z(n5) );
  NAND U20 ( .A(n2143), .B(n2142), .Z(n6) );
  NAND U21 ( .A(n5), .B(n6), .Z(n2248) );
  XNOR U22 ( .A(n2676), .B(n2675), .Z(n2677) );
  XNOR U23 ( .A(n2684), .B(n2683), .Z(n2701) );
  XNOR U24 ( .A(n2494), .B(n2493), .Z(n2388) );
  NAND U25 ( .A(n2254), .B(n2253), .Z(n7) );
  NAND U26 ( .A(n2251), .B(n2252), .Z(n8) );
  NAND U27 ( .A(n7), .B(n8), .Z(n2384) );
  XNOR U28 ( .A(n1943), .B(n1942), .Z(n2072) );
  NAND U29 ( .A(n2570), .B(n2571), .Z(n9) );
  XOR U30 ( .A(n2570), .B(n2571), .Z(n10) );
  NANDN U31 ( .A(n2569), .B(n10), .Z(n11) );
  NAND U32 ( .A(n9), .B(n11), .Z(n2749) );
  XOR U33 ( .A(n1168), .B(n1169), .Z(n12) );
  NANDN U34 ( .A(n1170), .B(n12), .Z(n13) );
  NAND U35 ( .A(n1168), .B(n1169), .Z(n14) );
  AND U36 ( .A(n13), .B(n14), .Z(n1286) );
  XNOR U37 ( .A(n3008), .B(n3007), .Z(n3000) );
  XNOR U38 ( .A(n1440), .B(n1439), .Z(n1496) );
  XNOR U39 ( .A(n1613), .B(n1612), .Z(n1576) );
  XNOR U40 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U41 ( .A(n1969), .B(n1968), .Z(n1974) );
  XNOR U42 ( .A(n1096), .B(n1095), .Z(n1112) );
  NAND U43 ( .A(n1015), .B(n1014), .Z(n15) );
  NANDN U44 ( .A(n1017), .B(n1016), .Z(n16) );
  AND U45 ( .A(n15), .B(n16), .Z(n1058) );
  XNOR U46 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U47 ( .A(n1240), .B(n1239), .Z(n1190) );
  XNOR U48 ( .A(n1706), .B(n1705), .Z(n1708) );
  XNOR U49 ( .A(n1748), .B(n1747), .Z(n1749) );
  XNOR U50 ( .A(n2199), .B(n2198), .Z(n2200) );
  NAND U51 ( .A(n2017), .B(n2016), .Z(n17) );
  NANDN U52 ( .A(n2019), .B(n2018), .Z(n18) );
  AND U53 ( .A(n17), .B(n18), .Z(n2097) );
  NAND U54 ( .A(n991), .B(n990), .Z(n19) );
  NANDN U55 ( .A(n993), .B(n992), .Z(n20) );
  AND U56 ( .A(n19), .B(n20), .Z(n1124) );
  XNOR U57 ( .A(n1257), .B(n1256), .Z(n1178) );
  XOR U58 ( .A(n1631), .B(n1630), .Z(n1634) );
  XNOR U59 ( .A(n1792), .B(n1791), .Z(n1778) );
  XNOR U60 ( .A(n2504), .B(n2503), .Z(n2505) );
  NAND U61 ( .A(n2103), .B(n2102), .Z(n21) );
  NAND U62 ( .A(n2101), .B(n2100), .Z(n22) );
  NAND U63 ( .A(n21), .B(n22), .Z(n2251) );
  XNOR U64 ( .A(n210), .B(n209), .Z(n212) );
  XNOR U65 ( .A(n2560), .B(n2559), .Z(n2678) );
  XOR U66 ( .A(n2564), .B(n2563), .Z(n2565) );
  XNOR U67 ( .A(n2388), .B(n2387), .Z(n2390) );
  NAND U68 ( .A(n2247), .B(n2248), .Z(n23) );
  NANDN U69 ( .A(n2250), .B(n2249), .Z(n24) );
  NAND U70 ( .A(n23), .B(n24), .Z(n2383) );
  XNOR U71 ( .A(n1647), .B(n1646), .Z(n1648) );
  XNOR U72 ( .A(n2211), .B(n2210), .Z(n2213) );
  XOR U73 ( .A(n2664), .B(n2663), .Z(n2666) );
  XNOR U74 ( .A(n2750), .B(n2749), .Z(n2748) );
  NAND U75 ( .A(n137), .B(n138), .Z(n25) );
  XOR U76 ( .A(n137), .B(n138), .Z(n26) );
  NANDN U77 ( .A(n136), .B(n26), .Z(n27) );
  NAND U78 ( .A(n25), .B(n27), .Z(n149) );
  XOR U79 ( .A(n206), .B(n205), .Z(n28) );
  NANDN U80 ( .A(n207), .B(n28), .Z(n29) );
  NAND U81 ( .A(n206), .B(n205), .Z(n30) );
  AND U82 ( .A(n29), .B(n30), .Z(n232) );
  NAND U83 ( .A(n330), .B(n331), .Z(n31) );
  XOR U84 ( .A(n330), .B(n331), .Z(n32) );
  NANDN U85 ( .A(n329), .B(n32), .Z(n33) );
  NAND U86 ( .A(n31), .B(n33), .Z(n383) );
  XOR U87 ( .A(n1518), .B(n1517), .Z(n34) );
  NANDN U88 ( .A(n1519), .B(n34), .Z(n35) );
  NAND U89 ( .A(n1518), .B(n1517), .Z(n36) );
  AND U90 ( .A(n35), .B(n36), .Z(n1652) );
  NAND U91 ( .A(n2069), .B(n2070), .Z(n37) );
  XOR U92 ( .A(n2069), .B(n2070), .Z(n38) );
  NANDN U93 ( .A(n2068), .B(n38), .Z(n39) );
  NAND U94 ( .A(n37), .B(n39), .Z(n2217) );
  XOR U95 ( .A(n2706), .B(n2707), .Z(n40) );
  NANDN U96 ( .A(n2708), .B(n40), .Z(n41) );
  NAND U97 ( .A(n2706), .B(n2707), .Z(n42) );
  AND U98 ( .A(n41), .B(n42), .Z(n2717) );
  XNOR U99 ( .A(n1878), .B(n1877), .Z(n1879) );
  XNOR U100 ( .A(n1686), .B(n1685), .Z(n1723) );
  XNOR U101 ( .A(n1601), .B(n1600), .Z(n1577) );
  XNOR U102 ( .A(n1973), .B(n1972), .Z(n1975) );
  XNOR U103 ( .A(n2181), .B(n2180), .Z(n2182) );
  OR U104 ( .A(n1009), .B(n1963), .Z(n43) );
  NAND U105 ( .A(n1011), .B(n1010), .Z(n44) );
  NAND U106 ( .A(n43), .B(n44), .Z(n1114) );
  XNOR U107 ( .A(n1607), .B(n1606), .Z(n1558) );
  XOR U108 ( .A(n1548), .B(n1547), .Z(n1623) );
  XNOR U109 ( .A(n1617), .B(n1616), .Z(n1619) );
  XNOR U110 ( .A(n1762), .B(n1761), .Z(n1750) );
  XNOR U111 ( .A(n2205), .B(n2204), .Z(n2206) );
  NAND U112 ( .A(n2155), .B(n2154), .Z(n45) );
  NAND U113 ( .A(n2153), .B(n2152), .Z(n46) );
  NAND U114 ( .A(n45), .B(n46), .Z(n2301) );
  XOR U115 ( .A(n2337), .B(n2336), .Z(n2266) );
  NAND U116 ( .A(n2188), .B(n2187), .Z(n47) );
  NAND U117 ( .A(n2186), .B(n2300), .Z(n48) );
  NAND U118 ( .A(n47), .B(n48), .Z(n2315) );
  XNOR U119 ( .A(n2193), .B(n2192), .Z(n2101) );
  XNOR U120 ( .A(n443), .B(n442), .Z(n444) );
  XNOR U121 ( .A(n536), .B(n535), .Z(n529) );
  XNOR U122 ( .A(n1178), .B(n1177), .Z(n1179) );
  XNOR U123 ( .A(n1289), .B(n1288), .Z(n1291) );
  XNOR U124 ( .A(n1325), .B(n1324), .Z(n1383) );
  XNOR U125 ( .A(n1536), .B(n1535), .Z(n1640) );
  XNOR U126 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U127 ( .A(n2262), .B(n2261), .Z(n49) );
  NAND U128 ( .A(n2259), .B(n2260), .Z(n50) );
  NAND U129 ( .A(n49), .B(n50), .Z(n2486) );
  NAND U130 ( .A(n2099), .B(n2098), .Z(n51) );
  NAND U131 ( .A(n2096), .B(n2097), .Z(n52) );
  NAND U132 ( .A(n51), .B(n52), .Z(n2253) );
  NAND U133 ( .A(n2141), .B(n2140), .Z(n53) );
  NAND U134 ( .A(n2139), .B(n2138), .Z(n54) );
  NAND U135 ( .A(n53), .B(n54), .Z(n2249) );
  XNOR U136 ( .A(n271), .B(n270), .Z(n272) );
  XNOR U137 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U138 ( .A(n1668), .B(n1667), .Z(n1656) );
  XNOR U139 ( .A(n1917), .B(n1916), .Z(n1923) );
  XNOR U140 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U141 ( .A(n2474), .B(n2473), .Z(n2476) );
  XOR U142 ( .A(n2776), .B(n2775), .Z(n2774) );
  XNOR U143 ( .A(n584), .B(n583), .Z(n586) );
  XOR U144 ( .A(n1275), .B(n1274), .Z(n1163) );
  XNOR U145 ( .A(n2678), .B(n2677), .Z(n2665) );
  XNOR U146 ( .A(n2734), .B(n2733), .Z(n2968) );
  NAND U147 ( .A(n126), .B(n125), .Z(n55) );
  NAND U148 ( .A(n124), .B(n131), .Z(n56) );
  NAND U149 ( .A(n55), .B(n56), .Z(n136) );
  XOR U150 ( .A(n179), .B(n178), .Z(n57) );
  NANDN U151 ( .A(n177), .B(n57), .Z(n58) );
  NAND U152 ( .A(n179), .B(n178), .Z(n59) );
  AND U153 ( .A(n58), .B(n59), .Z(n206) );
  NAND U154 ( .A(n283), .B(n284), .Z(n60) );
  XOR U155 ( .A(n283), .B(n284), .Z(n61) );
  NANDN U156 ( .A(n282), .B(n61), .Z(n62) );
  NAND U157 ( .A(n60), .B(n62), .Z(n330) );
  XOR U158 ( .A(n392), .B(n393), .Z(n63) );
  NANDN U159 ( .A(n394), .B(n63), .Z(n64) );
  NAND U160 ( .A(n392), .B(n393), .Z(n65) );
  AND U161 ( .A(n64), .B(n65), .Z(n510) );
  XOR U162 ( .A(n840), .B(n841), .Z(n66) );
  NANDN U163 ( .A(n842), .B(n66), .Z(n67) );
  NAND U164 ( .A(n840), .B(n841), .Z(n68) );
  AND U165 ( .A(n67), .B(n68), .Z(n941) );
  XNOR U166 ( .A(n1282), .B(n1281), .Z(n1285) );
  NAND U167 ( .A(n1653), .B(n1652), .Z(n69) );
  XOR U168 ( .A(n1653), .B(n1652), .Z(n70) );
  NANDN U169 ( .A(n1654), .B(n70), .Z(n71) );
  NAND U170 ( .A(n69), .B(n71), .Z(n1663) );
  NAND U171 ( .A(n2217), .B(n2216), .Z(n72) );
  XOR U172 ( .A(n2217), .B(n2216), .Z(n73) );
  NANDN U173 ( .A(n2218), .B(n73), .Z(n74) );
  NAND U174 ( .A(n72), .B(n74), .Z(n2227) );
  NAND U175 ( .A(n2544), .B(n2543), .Z(n75) );
  NAND U176 ( .A(n2542), .B(n2541), .Z(n76) );
  AND U177 ( .A(n75), .B(n76), .Z(n3002) );
  XNOR U178 ( .A(n1002), .B(n1001), .Z(n1014) );
  XNOR U179 ( .A(n1088), .B(n1087), .Z(n1090) );
  XNOR U180 ( .A(n1423), .B(n1422), .Z(n1440) );
  XNOR U181 ( .A(n1488), .B(n1487), .Z(n1489) );
  XNOR U182 ( .A(n1594), .B(n1593), .Z(n1596) );
  XNOR U183 ( .A(n1880), .B(n1879), .Z(n1820) );
  XNOR U184 ( .A(n1867), .B(n1868), .Z(n1844) );
  XNOR U185 ( .A(n2189), .B(o[26]), .Z(n2153) );
  XNOR U186 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U187 ( .A(n882), .B(n883), .Z(n77) );
  NANDN U188 ( .A(n1686), .B(n1082), .Z(n78) );
  NAND U189 ( .A(n77), .B(n78), .Z(n994) );
  XNOR U190 ( .A(n1084), .B(n1083), .Z(n1119) );
  XOR U191 ( .A(n1139), .B(n1138), .Z(n1059) );
  XNOR U192 ( .A(n1540), .B(n1539), .Z(n1542) );
  XOR U193 ( .A(n1560), .B(n1559), .Z(n1628) );
  XNOR U194 ( .A(n1579), .B(n1578), .Z(n1622) );
  XNOR U195 ( .A(n1534), .B(n1533), .Z(n1535) );
  XNOR U196 ( .A(n1712), .B(n1711), .Z(n1714) );
  NAND U197 ( .A(n2151), .B(n2150), .Z(n79) );
  NAND U198 ( .A(n2149), .B(n2335), .Z(n80) );
  NAND U199 ( .A(n79), .B(n80), .Z(n2302) );
  NAND U200 ( .A(n2113), .B(n2112), .Z(n81) );
  NAND U201 ( .A(n2111), .B(n2110), .Z(n82) );
  NAND U202 ( .A(n81), .B(n82), .Z(n2307) );
  NAND U203 ( .A(n2035), .B(n2034), .Z(n83) );
  NANDN U204 ( .A(n2037), .B(n2036), .Z(n84) );
  AND U205 ( .A(n83), .B(n84), .Z(n2102) );
  NAND U206 ( .A(n2028), .B(n2027), .Z(n85) );
  NAND U207 ( .A(n2026), .B(n2025), .Z(n86) );
  AND U208 ( .A(n85), .B(n86), .Z(n2144) );
  NAND U209 ( .A(n1963), .B(n1962), .Z(n87) );
  NANDN U210 ( .A(n1965), .B(n1964), .Z(n88) );
  AND U211 ( .A(n87), .B(n88), .Z(n2140) );
  XOR U212 ( .A(n546), .B(n547), .Z(n531) );
  NAND U213 ( .A(n987), .B(n986), .Z(n89) );
  NANDN U214 ( .A(n989), .B(n988), .Z(n90) );
  AND U215 ( .A(n89), .B(n90), .Z(n1125) );
  XOR U216 ( .A(n1251), .B(n1250), .Z(n1180) );
  XNOR U217 ( .A(n1192), .B(n1191), .Z(n1172) );
  XNOR U218 ( .A(n1384), .B(n1383), .Z(n1385) );
  XNOR U219 ( .A(n1637), .B(n1636), .Z(n1643) );
  XNOR U220 ( .A(n1915), .B(n1914), .Z(n1916) );
  XNOR U221 ( .A(n1850), .B(n1849), .Z(n1852) );
  XNOR U222 ( .A(n2201), .B(n2200), .Z(n2165) );
  XNOR U223 ( .A(n2207), .B(n2206), .Z(n2090) );
  XNOR U224 ( .A(n2242), .B(n2241), .Z(n2244) );
  XOR U225 ( .A(n2402), .B(n2401), .Z(n2506) );
  XNOR U226 ( .A(n2492), .B(n2491), .Z(n2493) );
  NAND U227 ( .A(n2255), .B(n2256), .Z(n91) );
  NANDN U228 ( .A(n2258), .B(n2257), .Z(n92) );
  NAND U229 ( .A(n91), .B(n92), .Z(n2487) );
  XNOR U230 ( .A(n196), .B(o[5]), .Z(n181) );
  XOR U231 ( .A(n481), .B(n480), .Z(n483) );
  XOR U232 ( .A(n1269), .B(n1268), .Z(n1273) );
  XOR U233 ( .A(n1411), .B(n1410), .Z(n1404) );
  XNOR U234 ( .A(n1666), .B(n1665), .Z(n1667) );
  XNOR U235 ( .A(n1947), .B(n1946), .Z(n1949) );
  XOR U236 ( .A(n2367), .B(n2366), .Z(n2230) );
  NAND U237 ( .A(n2327), .B(n2328), .Z(n93) );
  NANDN U238 ( .A(n2326), .B(n2325), .Z(n94) );
  NAND U239 ( .A(n93), .B(n94), .Z(n2475) );
  XOR U240 ( .A(n2380), .B(n2379), .Z(n2374) );
  XOR U241 ( .A(n2762), .B(n2761), .Z(n2760) );
  XNOR U242 ( .A(n2770), .B(n2769), .Z(n2767) );
  XOR U243 ( .A(n2782), .B(n2781), .Z(n2780) );
  XNOR U244 ( .A(n273), .B(n272), .Z(n277) );
  XOR U245 ( .A(n1799), .B(n1798), .Z(n1934) );
  XNOR U246 ( .A(n2072), .B(n2071), .Z(n2073) );
  XNOR U247 ( .A(n2682), .B(n2681), .Z(n2683) );
  XNOR U248 ( .A(n2990), .B(n2989), .Z(n2988) );
  XOR U249 ( .A(n2962), .B(n2961), .Z(n2960) );
  NAND U250 ( .A(n2386), .B(n2385), .Z(n95) );
  NAND U251 ( .A(n2384), .B(n2383), .Z(n96) );
  NAND U252 ( .A(n95), .B(n96), .Z(n2541) );
  XOR U253 ( .A(n149), .B(n150), .Z(n97) );
  NANDN U254 ( .A(n151), .B(n97), .Z(n98) );
  NAND U255 ( .A(n149), .B(n150), .Z(n99) );
  AND U256 ( .A(n98), .B(n99), .Z(n178) );
  XOR U257 ( .A(n232), .B(n233), .Z(n100) );
  NANDN U258 ( .A(n234), .B(n100), .Z(n101) );
  NAND U259 ( .A(n232), .B(n233), .Z(n102) );
  AND U260 ( .A(n101), .B(n102), .Z(n283) );
  NAND U261 ( .A(n383), .B(n384), .Z(n103) );
  XOR U262 ( .A(n383), .B(n384), .Z(n104) );
  NANDN U263 ( .A(n382), .B(n104), .Z(n105) );
  NAND U264 ( .A(n103), .B(n105), .Z(n392) );
  XOR U265 ( .A(n580), .B(n581), .Z(n106) );
  NANDN U266 ( .A(n582), .B(n106), .Z(n107) );
  NAND U267 ( .A(n580), .B(n581), .Z(n108) );
  AND U268 ( .A(n107), .B(n108), .Z(n598) );
  XOR U269 ( .A(n1036), .B(n1037), .Z(n109) );
  NANDN U270 ( .A(n1038), .B(n109), .Z(n110) );
  NAND U271 ( .A(n1036), .B(n1037), .Z(n111) );
  AND U272 ( .A(n110), .B(n111), .Z(n1155) );
  NAND U273 ( .A(n1286), .B(n1287), .Z(n112) );
  XOR U274 ( .A(n1286), .B(n1287), .Z(n113) );
  NAND U275 ( .A(n113), .B(n1285), .Z(n114) );
  NAND U276 ( .A(n112), .B(n114), .Z(n1518) );
  XOR U277 ( .A(n1663), .B(n1662), .Z(n115) );
  NANDN U278 ( .A(n1664), .B(n115), .Z(n116) );
  NAND U279 ( .A(n1663), .B(n1662), .Z(n117) );
  AND U280 ( .A(n116), .B(n117), .Z(n1927) );
  XOR U281 ( .A(n2227), .B(n2226), .Z(n118) );
  NANDN U282 ( .A(n2228), .B(n118), .Z(n119) );
  NAND U283 ( .A(n2227), .B(n2226), .Z(n120) );
  AND U284 ( .A(n119), .B(n120), .Z(n2534) );
  XNOR U285 ( .A(n2718), .B(n2717), .Z(n2715) );
  AND U286 ( .A(x[0]), .B(y[0]), .Z(n763) );
  XOR U287 ( .A(n763), .B(o[0]), .Z(N33) );
  NAND U288 ( .A(y[0]), .B(x[1]), .Z(n131) );
  AND U289 ( .A(x[0]), .B(y[1]), .Z(n123) );
  XNOR U290 ( .A(n123), .B(o[1]), .Z(n124) );
  XOR U291 ( .A(n131), .B(n124), .Z(n126) );
  NAND U292 ( .A(n763), .B(o[0]), .Z(n125) );
  XNOR U293 ( .A(n126), .B(n125), .Z(N34) );
  AND U294 ( .A(x[2]), .B(y[0]), .Z(n122) );
  NAND U295 ( .A(x[1]), .B(y[1]), .Z(n121) );
  XNOR U296 ( .A(n122), .B(n121), .Z(n132) );
  AND U297 ( .A(n123), .B(o[1]), .Z(n133) );
  XOR U298 ( .A(n132), .B(n133), .Z(n138) );
  AND U299 ( .A(x[0]), .B(y[2]), .Z(n130) );
  XOR U300 ( .A(o[2]), .B(n130), .Z(n137) );
  XOR U301 ( .A(n136), .B(n137), .Z(n127) );
  XNOR U302 ( .A(n138), .B(n127), .Z(N35) );
  AND U303 ( .A(y[2]), .B(x[1]), .Z(n248) );
  AND U304 ( .A(y[1]), .B(x[2]), .Z(n147) );
  XOR U305 ( .A(n147), .B(o[3]), .Z(n152) );
  XOR U306 ( .A(n248), .B(n152), .Z(n154) );
  AND U307 ( .A(y[3]), .B(x[0]), .Z(n129) );
  NAND U308 ( .A(y[0]), .B(x[3]), .Z(n128) );
  XNOR U309 ( .A(n129), .B(n128), .Z(n142) );
  AND U310 ( .A(o[2]), .B(n130), .Z(n141) );
  XOR U311 ( .A(n142), .B(n141), .Z(n153) );
  XNOR U312 ( .A(n154), .B(n153), .Z(n151) );
  NANDN U313 ( .A(n131), .B(n147), .Z(n135) );
  NAND U314 ( .A(n133), .B(n132), .Z(n134) );
  NAND U315 ( .A(n135), .B(n134), .Z(n150) );
  XOR U316 ( .A(n150), .B(n149), .Z(n139) );
  XNOR U317 ( .A(n151), .B(n139), .Z(N36) );
  AND U318 ( .A(x[3]), .B(y[3]), .Z(n140) );
  NAND U319 ( .A(n763), .B(n140), .Z(n144) );
  NAND U320 ( .A(n142), .B(n141), .Z(n143) );
  AND U321 ( .A(n144), .B(n143), .Z(n174) );
  AND U322 ( .A(x[4]), .B(y[0]), .Z(n146) );
  NAND U323 ( .A(y[4]), .B(x[0]), .Z(n145) );
  XNOR U324 ( .A(n146), .B(n145), .Z(n168) );
  AND U325 ( .A(n147), .B(o[3]), .Z(n167) );
  XOR U326 ( .A(n168), .B(n167), .Z(n172) );
  AND U327 ( .A(x[1]), .B(y[3]), .Z(n352) );
  NAND U328 ( .A(y[2]), .B(x[2]), .Z(n148) );
  XNOR U329 ( .A(n352), .B(n148), .Z(n164) );
  AND U330 ( .A(x[3]), .B(y[1]), .Z(n162) );
  XOR U331 ( .A(n162), .B(o[4]), .Z(n163) );
  XOR U332 ( .A(n164), .B(n163), .Z(n171) );
  XOR U333 ( .A(n172), .B(n171), .Z(n173) );
  XOR U334 ( .A(n174), .B(n173), .Z(n179) );
  NAND U335 ( .A(n248), .B(n152), .Z(n156) );
  NAND U336 ( .A(n154), .B(n153), .Z(n155) );
  NAND U337 ( .A(n156), .B(n155), .Z(n177) );
  XNOR U338 ( .A(n178), .B(n177), .Z(n157) );
  XNOR U339 ( .A(n179), .B(n157), .Z(N37) );
  AND U340 ( .A(x[2]), .B(y[3]), .Z(n258) );
  AND U341 ( .A(x[1]), .B(y[4]), .Z(n159) );
  NAND U342 ( .A(y[2]), .B(x[3]), .Z(n158) );
  XNOR U343 ( .A(n159), .B(n158), .Z(n182) );
  NAND U344 ( .A(y[1]), .B(x[4]), .Z(n196) );
  XOR U345 ( .A(n182), .B(n181), .Z(n185) );
  XOR U346 ( .A(n258), .B(n185), .Z(n187) );
  AND U347 ( .A(x[5]), .B(y[0]), .Z(n161) );
  NAND U348 ( .A(x[0]), .B(y[5]), .Z(n160) );
  XNOR U349 ( .A(n161), .B(n160), .Z(n191) );
  AND U350 ( .A(n162), .B(o[4]), .Z(n190) );
  XOR U351 ( .A(n191), .B(n190), .Z(n186) );
  XOR U352 ( .A(n187), .B(n186), .Z(n202) );
  NAND U353 ( .A(n258), .B(n248), .Z(n166) );
  NAND U354 ( .A(n164), .B(n163), .Z(n165) );
  NAND U355 ( .A(n166), .B(n165), .Z(n200) );
  AND U356 ( .A(y[4]), .B(x[4]), .Z(n965) );
  NAND U357 ( .A(n965), .B(n763), .Z(n170) );
  NAND U358 ( .A(n168), .B(n167), .Z(n169) );
  NAND U359 ( .A(n170), .B(n169), .Z(n199) );
  XOR U360 ( .A(n200), .B(n199), .Z(n201) );
  XNOR U361 ( .A(n202), .B(n201), .Z(n207) );
  NAND U362 ( .A(n172), .B(n171), .Z(n176) );
  NANDN U363 ( .A(n174), .B(n173), .Z(n175) );
  NAND U364 ( .A(n176), .B(n175), .Z(n205) );
  XOR U365 ( .A(n205), .B(n206), .Z(n180) );
  XNOR U366 ( .A(n207), .B(n180), .Z(N38) );
  AND U367 ( .A(x[3]), .B(y[4]), .Z(n259) );
  NAND U368 ( .A(n259), .B(n248), .Z(n184) );
  NAND U369 ( .A(n182), .B(n181), .Z(n183) );
  NAND U370 ( .A(n184), .B(n183), .Z(n236) );
  NAND U371 ( .A(n258), .B(n185), .Z(n189) );
  NAND U372 ( .A(n187), .B(n186), .Z(n188) );
  NAND U373 ( .A(n189), .B(n188), .Z(n235) );
  XOR U374 ( .A(n236), .B(n235), .Z(n238) );
  AND U375 ( .A(y[5]), .B(x[5]), .Z(n438) );
  NAND U376 ( .A(n763), .B(n438), .Z(n193) );
  NAND U377 ( .A(n191), .B(n190), .Z(n192) );
  AND U378 ( .A(n193), .B(n192), .Z(n210) );
  AND U379 ( .A(x[6]), .B(y[0]), .Z(n195) );
  NAND U380 ( .A(x[0]), .B(y[6]), .Z(n194) );
  XNOR U381 ( .A(n195), .B(n194), .Z(n217) );
  ANDN U382 ( .B(o[5]), .A(n196), .Z(n216) );
  XOR U383 ( .A(n217), .B(n216), .Z(n209) );
  AND U384 ( .A(y[4]), .B(x[2]), .Z(n729) );
  NAND U385 ( .A(y[3]), .B(x[3]), .Z(n197) );
  XNOR U386 ( .A(n729), .B(n197), .Z(n221) );
  AND U387 ( .A(x[4]), .B(y[2]), .Z(n565) );
  NAND U388 ( .A(x[1]), .B(y[5]), .Z(n198) );
  XNOR U389 ( .A(n565), .B(n198), .Z(n225) );
  AND U390 ( .A(y[1]), .B(x[5]), .Z(n231) );
  XOR U391 ( .A(o[6]), .B(n231), .Z(n224) );
  XOR U392 ( .A(n225), .B(n224), .Z(n220) );
  XOR U393 ( .A(n221), .B(n220), .Z(n211) );
  XOR U394 ( .A(n212), .B(n211), .Z(n237) );
  XOR U395 ( .A(n238), .B(n237), .Z(n234) );
  NAND U396 ( .A(n200), .B(n199), .Z(n204) );
  NAND U397 ( .A(n202), .B(n201), .Z(n203) );
  AND U398 ( .A(n204), .B(n203), .Z(n233) );
  XNOR U399 ( .A(n233), .B(n232), .Z(n208) );
  XNOR U400 ( .A(n234), .B(n208), .Z(N39) );
  NANDN U401 ( .A(n210), .B(n209), .Z(n214) );
  NAND U402 ( .A(n212), .B(n211), .Z(n213) );
  AND U403 ( .A(n214), .B(n213), .Z(n279) );
  AND U404 ( .A(x[5]), .B(y[2]), .Z(n339) );
  NAND U405 ( .A(x[1]), .B(y[6]), .Z(n215) );
  XNOR U406 ( .A(n339), .B(n215), .Z(n251) );
  AND U407 ( .A(y[1]), .B(x[6]), .Z(n255) );
  XOR U408 ( .A(o[7]), .B(n255), .Z(n250) );
  XOR U409 ( .A(n251), .B(n250), .Z(n271) );
  AND U410 ( .A(y[6]), .B(x[6]), .Z(n287) );
  NAND U411 ( .A(n763), .B(n287), .Z(n219) );
  NAND U412 ( .A(n217), .B(n216), .Z(n218) );
  AND U413 ( .A(n219), .B(n218), .Z(n270) );
  NAND U414 ( .A(n258), .B(n259), .Z(n223) );
  NAND U415 ( .A(n221), .B(n220), .Z(n222) );
  NAND U416 ( .A(n223), .B(n222), .Z(n273) );
  AND U417 ( .A(y[5]), .B(x[4]), .Z(n768) );
  NAND U418 ( .A(n768), .B(n248), .Z(n227) );
  NAND U419 ( .A(n225), .B(n224), .Z(n226) );
  AND U420 ( .A(n227), .B(n226), .Z(n245) );
  AND U421 ( .A(x[4]), .B(y[3]), .Z(n413) );
  NAND U422 ( .A(x[2]), .B(y[5]), .Z(n228) );
  XNOR U423 ( .A(n413), .B(n228), .Z(n260) );
  XNOR U424 ( .A(n260), .B(n259), .Z(n243) );
  AND U425 ( .A(x[7]), .B(y[0]), .Z(n230) );
  NAND U426 ( .A(y[7]), .B(x[0]), .Z(n229) );
  XNOR U427 ( .A(n230), .B(n229), .Z(n265) );
  AND U428 ( .A(o[6]), .B(n231), .Z(n264) );
  XNOR U429 ( .A(n265), .B(n264), .Z(n242) );
  XOR U430 ( .A(n243), .B(n242), .Z(n244) );
  XOR U431 ( .A(n245), .B(n244), .Z(n276) );
  XOR U432 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U433 ( .A(n279), .B(n278), .Z(n284) );
  NAND U434 ( .A(n236), .B(n235), .Z(n240) );
  NAND U435 ( .A(n238), .B(n237), .Z(n239) );
  AND U436 ( .A(n240), .B(n239), .Z(n282) );
  XOR U437 ( .A(n283), .B(n282), .Z(n241) );
  XNOR U438 ( .A(n284), .B(n241), .Z(N40) );
  NAND U439 ( .A(n243), .B(n242), .Z(n247) );
  NAND U440 ( .A(n245), .B(n244), .Z(n246) );
  AND U441 ( .A(n247), .B(n246), .Z(n320) );
  AND U442 ( .A(y[6]), .B(x[5]), .Z(n249) );
  NAND U443 ( .A(n249), .B(n248), .Z(n253) );
  NAND U444 ( .A(n251), .B(n250), .Z(n252) );
  NAND U445 ( .A(n253), .B(n252), .Z(n318) );
  AND U446 ( .A(x[1]), .B(y[7]), .Z(n758) );
  NAND U447 ( .A(y[3]), .B(x[5]), .Z(n254) );
  XNOR U448 ( .A(n758), .B(n254), .Z(n308) );
  AND U449 ( .A(o[7]), .B(n255), .Z(n307) );
  XOR U450 ( .A(n308), .B(n307), .Z(n293) );
  NAND U451 ( .A(y[5]), .B(x[3]), .Z(n1094) );
  AND U452 ( .A(y[2]), .B(x[6]), .Z(n257) );
  NAND U453 ( .A(x[2]), .B(y[6]), .Z(n256) );
  XNOR U454 ( .A(n257), .B(n256), .Z(n288) );
  XNOR U455 ( .A(n965), .B(n288), .Z(n291) );
  XOR U456 ( .A(n1094), .B(n291), .Z(n292) );
  XOR U457 ( .A(n293), .B(n292), .Z(n317) );
  XOR U458 ( .A(n318), .B(n317), .Z(n319) );
  XOR U459 ( .A(n320), .B(n319), .Z(n326) );
  NAND U460 ( .A(n768), .B(n258), .Z(n262) );
  NAND U461 ( .A(n260), .B(n259), .Z(n261) );
  NAND U462 ( .A(n262), .B(n261), .Z(n314) );
  AND U463 ( .A(x[7]), .B(y[7]), .Z(n263) );
  NAND U464 ( .A(n763), .B(n263), .Z(n267) );
  NAND U465 ( .A(n265), .B(n264), .Z(n266) );
  NAND U466 ( .A(n267), .B(n266), .Z(n312) );
  AND U467 ( .A(x[8]), .B(y[0]), .Z(n269) );
  NAND U468 ( .A(y[8]), .B(x[0]), .Z(n268) );
  XNOR U469 ( .A(n269), .B(n268), .Z(n298) );
  AND U470 ( .A(y[1]), .B(x[7]), .Z(n303) );
  XOR U471 ( .A(o[8]), .B(n303), .Z(n297) );
  XOR U472 ( .A(n298), .B(n297), .Z(n311) );
  XOR U473 ( .A(n312), .B(n311), .Z(n313) );
  XNOR U474 ( .A(n314), .B(n313), .Z(n324) );
  NANDN U475 ( .A(n271), .B(n270), .Z(n275) );
  NANDN U476 ( .A(n273), .B(n272), .Z(n274) );
  NAND U477 ( .A(n275), .B(n274), .Z(n323) );
  XOR U478 ( .A(n324), .B(n323), .Z(n325) );
  XOR U479 ( .A(n326), .B(n325), .Z(n331) );
  NAND U480 ( .A(n277), .B(n276), .Z(n281) );
  NAND U481 ( .A(n279), .B(n278), .Z(n280) );
  NAND U482 ( .A(n281), .B(n280), .Z(n329) );
  XOR U483 ( .A(n329), .B(n330), .Z(n285) );
  XNOR U484 ( .A(n331), .B(n285), .Z(N41) );
  AND U485 ( .A(x[2]), .B(y[2]), .Z(n286) );
  NAND U486 ( .A(n287), .B(n286), .Z(n290) );
  NAND U487 ( .A(n965), .B(n288), .Z(n289) );
  NAND U488 ( .A(n290), .B(n289), .Z(n334) );
  NAND U489 ( .A(n1094), .B(n291), .Z(n295) );
  NANDN U490 ( .A(n293), .B(n292), .Z(n294) );
  AND U491 ( .A(n295), .B(n294), .Z(n333) );
  XOR U492 ( .A(n334), .B(n333), .Z(n336) );
  AND U493 ( .A(x[8]), .B(y[8]), .Z(n296) );
  NAND U494 ( .A(n296), .B(n763), .Z(n300) );
  NAND U495 ( .A(n298), .B(n297), .Z(n299) );
  AND U496 ( .A(n300), .B(n299), .Z(n369) );
  AND U497 ( .A(x[5]), .B(y[4]), .Z(n302) );
  NAND U498 ( .A(y[2]), .B(x[7]), .Z(n301) );
  XNOR U499 ( .A(n302), .B(n301), .Z(n342) );
  AND U500 ( .A(o[8]), .B(n303), .Z(n341) );
  XNOR U501 ( .A(n342), .B(n341), .Z(n367) );
  AND U502 ( .A(x[9]), .B(y[0]), .Z(n305) );
  NAND U503 ( .A(y[9]), .B(x[0]), .Z(n304) );
  XNOR U504 ( .A(n305), .B(n304), .Z(n349) );
  AND U505 ( .A(y[1]), .B(x[8]), .Z(n358) );
  XOR U506 ( .A(o[9]), .B(n358), .Z(n348) );
  XNOR U507 ( .A(n349), .B(n348), .Z(n366) );
  XOR U508 ( .A(n367), .B(n366), .Z(n368) );
  XNOR U509 ( .A(n369), .B(n368), .Z(n363) );
  AND U510 ( .A(x[1]), .B(y[8]), .Z(n1082) );
  NAND U511 ( .A(y[3]), .B(x[6]), .Z(n306) );
  XNOR U512 ( .A(n1082), .B(n306), .Z(n353) );
  XNOR U513 ( .A(n768), .B(n353), .Z(n373) );
  NAND U514 ( .A(x[2]), .B(y[7]), .Z(n1009) );
  AND U515 ( .A(y[6]), .B(x[3]), .Z(n703) );
  XNOR U516 ( .A(n1009), .B(n703), .Z(n372) );
  XNOR U517 ( .A(n373), .B(n372), .Z(n361) );
  NAND U518 ( .A(x[5]), .B(y[7]), .Z(n545) );
  NANDN U519 ( .A(n545), .B(n352), .Z(n310) );
  NAND U520 ( .A(n308), .B(n307), .Z(n309) );
  NAND U521 ( .A(n310), .B(n309), .Z(n360) );
  XOR U522 ( .A(n361), .B(n360), .Z(n362) );
  XOR U523 ( .A(n363), .B(n362), .Z(n335) );
  XOR U524 ( .A(n336), .B(n335), .Z(n379) );
  NAND U525 ( .A(n312), .B(n311), .Z(n316) );
  NAND U526 ( .A(n314), .B(n313), .Z(n315) );
  NAND U527 ( .A(n316), .B(n315), .Z(n377) );
  NAND U528 ( .A(n318), .B(n317), .Z(n322) );
  NAND U529 ( .A(n320), .B(n319), .Z(n321) );
  NAND U530 ( .A(n322), .B(n321), .Z(n376) );
  XOR U531 ( .A(n377), .B(n376), .Z(n378) );
  XOR U532 ( .A(n379), .B(n378), .Z(n384) );
  NAND U533 ( .A(n324), .B(n323), .Z(n328) );
  NANDN U534 ( .A(n326), .B(n325), .Z(n327) );
  NAND U535 ( .A(n328), .B(n327), .Z(n382) );
  XOR U536 ( .A(n382), .B(n383), .Z(n332) );
  XNOR U537 ( .A(n384), .B(n332), .Z(N42) );
  NAND U538 ( .A(n334), .B(n333), .Z(n338) );
  NAND U539 ( .A(n336), .B(n335), .Z(n337) );
  AND U540 ( .A(n338), .B(n337), .Z(n389) );
  AND U541 ( .A(x[7]), .B(y[4]), .Z(n340) );
  NAND U542 ( .A(n340), .B(n339), .Z(n344) );
  NAND U543 ( .A(n342), .B(n341), .Z(n343) );
  AND U544 ( .A(n344), .B(n343), .Z(n445) );
  AND U545 ( .A(y[3]), .B(x[7]), .Z(n346) );
  NAND U546 ( .A(x[4]), .B(y[6]), .Z(n345) );
  XNOR U547 ( .A(n346), .B(n345), .Z(n415) );
  AND U548 ( .A(x[6]), .B(y[4]), .Z(n416) );
  XOR U549 ( .A(n415), .B(n416), .Z(n443) );
  AND U550 ( .A(x[8]), .B(y[2]), .Z(n627) );
  AND U551 ( .A(y[1]), .B(x[9]), .Z(n426) );
  XOR U552 ( .A(o[10]), .B(n426), .Z(n437) );
  XOR U553 ( .A(n627), .B(n437), .Z(n439) );
  XNOR U554 ( .A(n439), .B(n438), .Z(n442) );
  XNOR U555 ( .A(n445), .B(n444), .Z(n404) );
  AND U556 ( .A(y[9]), .B(x[9]), .Z(n347) );
  NAND U557 ( .A(n347), .B(n763), .Z(n351) );
  NAND U558 ( .A(n349), .B(n348), .Z(n350) );
  NAND U559 ( .A(n351), .B(n350), .Z(n402) );
  AND U560 ( .A(x[6]), .B(y[8]), .Z(n662) );
  NAND U561 ( .A(n662), .B(n352), .Z(n355) );
  NAND U562 ( .A(n768), .B(n353), .Z(n354) );
  NAND U563 ( .A(n355), .B(n354), .Z(n410) );
  AND U564 ( .A(x[10]), .B(y[0]), .Z(n357) );
  NAND U565 ( .A(y[10]), .B(x[0]), .Z(n356) );
  XNOR U566 ( .A(n357), .B(n356), .Z(n421) );
  AND U567 ( .A(o[9]), .B(n358), .Z(n420) );
  XOR U568 ( .A(n421), .B(n420), .Z(n408) );
  AND U569 ( .A(x[1]), .B(y[9]), .Z(n1305) );
  NAND U570 ( .A(y[7]), .B(x[3]), .Z(n359) );
  XNOR U571 ( .A(n1305), .B(n359), .Z(n433) );
  AND U572 ( .A(y[8]), .B(x[2]), .Z(n434) );
  XOR U573 ( .A(n433), .B(n434), .Z(n407) );
  XOR U574 ( .A(n408), .B(n407), .Z(n409) );
  XOR U575 ( .A(n410), .B(n409), .Z(n401) );
  XOR U576 ( .A(n402), .B(n401), .Z(n403) );
  XNOR U577 ( .A(n404), .B(n403), .Z(n387) );
  NAND U578 ( .A(n361), .B(n360), .Z(n365) );
  NAND U579 ( .A(n363), .B(n362), .Z(n364) );
  AND U580 ( .A(n365), .B(n364), .Z(n398) );
  NAND U581 ( .A(n367), .B(n366), .Z(n371) );
  NAND U582 ( .A(n369), .B(n368), .Z(n370) );
  AND U583 ( .A(n371), .B(n370), .Z(n395) );
  NAND U584 ( .A(n373), .B(n372), .Z(n375) );
  ANDN U585 ( .B(n1009), .A(n703), .Z(n374) );
  ANDN U586 ( .B(n375), .A(n374), .Z(n396) );
  XOR U587 ( .A(n395), .B(n396), .Z(n397) );
  XOR U588 ( .A(n398), .B(n397), .Z(n386) );
  XOR U589 ( .A(n387), .B(n386), .Z(n388) );
  XOR U590 ( .A(n389), .B(n388), .Z(n394) );
  NAND U591 ( .A(n377), .B(n376), .Z(n381) );
  NAND U592 ( .A(n379), .B(n378), .Z(n380) );
  NAND U593 ( .A(n381), .B(n380), .Z(n393) );
  XOR U594 ( .A(n393), .B(n392), .Z(n385) );
  XNOR U595 ( .A(n394), .B(n385), .Z(N43) );
  NAND U596 ( .A(n387), .B(n386), .Z(n391) );
  NAND U597 ( .A(n389), .B(n388), .Z(n390) );
  NAND U598 ( .A(n391), .B(n390), .Z(n511) );
  IV U599 ( .A(n511), .Z(n509) );
  NAND U600 ( .A(n396), .B(n395), .Z(n400) );
  NANDN U601 ( .A(n398), .B(n397), .Z(n399) );
  NAND U602 ( .A(n400), .B(n399), .Z(n506) );
  NAND U603 ( .A(n402), .B(n401), .Z(n406) );
  NAND U604 ( .A(n404), .B(n403), .Z(n405) );
  NAND U605 ( .A(n406), .B(n405), .Z(n504) );
  NAND U606 ( .A(n408), .B(n407), .Z(n412) );
  NAND U607 ( .A(n410), .B(n409), .Z(n411) );
  NAND U608 ( .A(n412), .B(n411), .Z(n500) );
  AND U609 ( .A(y[6]), .B(x[7]), .Z(n414) );
  NAND U610 ( .A(n414), .B(n413), .Z(n418) );
  NAND U611 ( .A(n416), .B(n415), .Z(n417) );
  NAND U612 ( .A(n418), .B(n417), .Z(n498) );
  AND U613 ( .A(y[10]), .B(x[10]), .Z(n419) );
  NAND U614 ( .A(n419), .B(n763), .Z(n423) );
  NAND U615 ( .A(n421), .B(n420), .Z(n422) );
  NAND U616 ( .A(n423), .B(n422), .Z(n494) );
  AND U617 ( .A(y[11]), .B(x[0]), .Z(n425) );
  NAND U618 ( .A(y[0]), .B(x[11]), .Z(n424) );
  XNOR U619 ( .A(n425), .B(n424), .Z(n471) );
  AND U620 ( .A(o[10]), .B(n426), .Z(n470) );
  XOR U621 ( .A(n471), .B(n470), .Z(n492) );
  AND U622 ( .A(x[1]), .B(y[10]), .Z(n428) );
  NAND U623 ( .A(x[6]), .B(y[5]), .Z(n427) );
  XNOR U624 ( .A(n428), .B(n427), .Z(n462) );
  AND U625 ( .A(y[1]), .B(x[10]), .Z(n479) );
  XOR U626 ( .A(o[11]), .B(n479), .Z(n461) );
  XOR U627 ( .A(n462), .B(n461), .Z(n491) );
  XOR U628 ( .A(n492), .B(n491), .Z(n493) );
  XOR U629 ( .A(n494), .B(n493), .Z(n497) );
  XOR U630 ( .A(n498), .B(n497), .Z(n499) );
  XNOR U631 ( .A(n500), .B(n499), .Z(n482) );
  AND U632 ( .A(x[3]), .B(y[8]), .Z(n1459) );
  AND U633 ( .A(x[2]), .B(y[9]), .Z(n430) );
  NAND U634 ( .A(x[5]), .B(y[6]), .Z(n429) );
  XNOR U635 ( .A(n430), .B(n429), .Z(n456) );
  AND U636 ( .A(y[7]), .B(x[4]), .Z(n455) );
  XNOR U637 ( .A(n456), .B(n455), .Z(n486) );
  XNOR U638 ( .A(n1459), .B(n486), .Z(n488) );
  AND U639 ( .A(x[9]), .B(y[2]), .Z(n432) );
  NAND U640 ( .A(y[4]), .B(x[7]), .Z(n431) );
  XNOR U641 ( .A(n432), .B(n431), .Z(n475) );
  AND U642 ( .A(x[8]), .B(y[3]), .Z(n474) );
  XNOR U643 ( .A(n475), .B(n474), .Z(n487) );
  XNOR U644 ( .A(n488), .B(n487), .Z(n452) );
  NAND U645 ( .A(x[3]), .B(y[9]), .Z(n536) );
  NANDN U646 ( .A(n536), .B(n758), .Z(n436) );
  NAND U647 ( .A(n434), .B(n433), .Z(n435) );
  NAND U648 ( .A(n436), .B(n435), .Z(n450) );
  NAND U649 ( .A(n627), .B(n437), .Z(n441) );
  NAND U650 ( .A(n439), .B(n438), .Z(n440) );
  NAND U651 ( .A(n441), .B(n440), .Z(n449) );
  XOR U652 ( .A(n450), .B(n449), .Z(n451) );
  XOR U653 ( .A(n452), .B(n451), .Z(n481) );
  NANDN U654 ( .A(n443), .B(n442), .Z(n447) );
  NAND U655 ( .A(n445), .B(n444), .Z(n446) );
  NAND U656 ( .A(n447), .B(n446), .Z(n480) );
  XOR U657 ( .A(n482), .B(n483), .Z(n503) );
  XOR U658 ( .A(n504), .B(n503), .Z(n505) );
  XOR U659 ( .A(n506), .B(n505), .Z(n512) );
  XNOR U660 ( .A(n510), .B(n512), .Z(n448) );
  XOR U661 ( .A(n509), .B(n448), .Z(N44) );
  NAND U662 ( .A(n450), .B(n449), .Z(n454) );
  NAND U663 ( .A(n452), .B(n451), .Z(n453) );
  NAND U664 ( .A(n454), .B(n453), .Z(n577) );
  AND U665 ( .A(y[6]), .B(x[2]), .Z(n1206) );
  AND U666 ( .A(y[9]), .B(x[5]), .Z(n1000) );
  NAND U667 ( .A(n1206), .B(n1000), .Z(n458) );
  NAND U668 ( .A(n456), .B(n455), .Z(n457) );
  NAND U669 ( .A(n458), .B(n457), .Z(n524) );
  AND U670 ( .A(y[10]), .B(x[6]), .Z(n460) );
  AND U671 ( .A(y[5]), .B(x[1]), .Z(n459) );
  NAND U672 ( .A(n460), .B(n459), .Z(n464) );
  NAND U673 ( .A(n462), .B(n461), .Z(n463) );
  NAND U674 ( .A(n464), .B(n463), .Z(n523) );
  XOR U675 ( .A(n524), .B(n523), .Z(n526) );
  AND U676 ( .A(y[3]), .B(x[9]), .Z(n1201) );
  AND U677 ( .A(x[10]), .B(y[2]), .Z(n1243) );
  NAND U678 ( .A(x[4]), .B(y[8]), .Z(n465) );
  XNOR U679 ( .A(n1243), .B(n465), .Z(n567) );
  XOR U680 ( .A(n1201), .B(n567), .Z(n546) );
  NAND U681 ( .A(y[5]), .B(x[7]), .Z(n544) );
  XOR U682 ( .A(n545), .B(n544), .Z(n547) );
  AND U683 ( .A(x[12]), .B(y[0]), .Z(n467) );
  NAND U684 ( .A(x[0]), .B(y[12]), .Z(n466) );
  XNOR U685 ( .A(n467), .B(n466), .Z(n561) );
  AND U686 ( .A(x[11]), .B(y[1]), .Z(n541) );
  XOR U687 ( .A(o[12]), .B(n541), .Z(n560) );
  XOR U688 ( .A(n561), .B(n560), .Z(n530) );
  AND U689 ( .A(y[4]), .B(x[8]), .Z(n469) );
  NAND U690 ( .A(x[2]), .B(y[10]), .Z(n468) );
  XNOR U691 ( .A(n469), .B(n468), .Z(n535) );
  XOR U692 ( .A(n530), .B(n529), .Z(n532) );
  XOR U693 ( .A(n531), .B(n532), .Z(n525) );
  XOR U694 ( .A(n526), .B(n525), .Z(n575) );
  AND U695 ( .A(x[11]), .B(y[11]), .Z(n1572) );
  NAND U696 ( .A(n1572), .B(n763), .Z(n473) );
  NAND U697 ( .A(n471), .B(n470), .Z(n472) );
  NAND U698 ( .A(n473), .B(n472), .Z(n553) );
  AND U699 ( .A(x[7]), .B(y[2]), .Z(n719) );
  AND U700 ( .A(y[4]), .B(x[9]), .Z(n543) );
  NAND U701 ( .A(n719), .B(n543), .Z(n477) );
  NAND U702 ( .A(n475), .B(n474), .Z(n476) );
  NAND U703 ( .A(n477), .B(n476), .Z(n551) );
  AND U704 ( .A(x[1]), .B(y[11]), .Z(n1238) );
  NAND U705 ( .A(x[6]), .B(y[6]), .Z(n478) );
  XNOR U706 ( .A(n1238), .B(n478), .Z(n557) );
  AND U707 ( .A(o[11]), .B(n479), .Z(n556) );
  XOR U708 ( .A(n557), .B(n556), .Z(n550) );
  XOR U709 ( .A(n551), .B(n550), .Z(n552) );
  XOR U710 ( .A(n553), .B(n552), .Z(n574) );
  XOR U711 ( .A(n575), .B(n574), .Z(n576) );
  XOR U712 ( .A(n577), .B(n576), .Z(n584) );
  NANDN U713 ( .A(n481), .B(n480), .Z(n485) );
  NANDN U714 ( .A(n483), .B(n482), .Z(n484) );
  NAND U715 ( .A(n485), .B(n484), .Z(n583) );
  NANDN U716 ( .A(n1459), .B(n486), .Z(n490) );
  NAND U717 ( .A(n488), .B(n487), .Z(n489) );
  NAND U718 ( .A(n490), .B(n489), .Z(n518) );
  NAND U719 ( .A(n492), .B(n491), .Z(n496) );
  NAND U720 ( .A(n494), .B(n493), .Z(n495) );
  AND U721 ( .A(n496), .B(n495), .Z(n517) );
  XOR U722 ( .A(n518), .B(n517), .Z(n520) );
  NAND U723 ( .A(n498), .B(n497), .Z(n502) );
  NAND U724 ( .A(n500), .B(n499), .Z(n501) );
  AND U725 ( .A(n502), .B(n501), .Z(n519) );
  XOR U726 ( .A(n520), .B(n519), .Z(n585) );
  XOR U727 ( .A(n586), .B(n585), .Z(n582) );
  NAND U728 ( .A(n504), .B(n503), .Z(n508) );
  NAND U729 ( .A(n506), .B(n505), .Z(n507) );
  NAND U730 ( .A(n508), .B(n507), .Z(n581) );
  NANDN U731 ( .A(n509), .B(n510), .Z(n515) );
  NOR U732 ( .A(n511), .B(n510), .Z(n513) );
  OR U733 ( .A(n513), .B(n512), .Z(n514) );
  AND U734 ( .A(n515), .B(n514), .Z(n580) );
  XOR U735 ( .A(n581), .B(n580), .Z(n516) );
  XNOR U736 ( .A(n582), .B(n516), .Z(N45) );
  NAND U737 ( .A(n518), .B(n517), .Z(n522) );
  NAND U738 ( .A(n520), .B(n519), .Z(n521) );
  NAND U739 ( .A(n522), .B(n521), .Z(n593) );
  NAND U740 ( .A(n524), .B(n523), .Z(n528) );
  NAND U741 ( .A(n526), .B(n525), .Z(n527) );
  NAND U742 ( .A(n528), .B(n527), .Z(n604) );
  NAND U743 ( .A(n530), .B(n529), .Z(n534) );
  NAND U744 ( .A(n532), .B(n531), .Z(n533) );
  NAND U745 ( .A(n534), .B(n533), .Z(n611) );
  AND U746 ( .A(y[10]), .B(x[8]), .Z(n1860) );
  NAND U747 ( .A(n1860), .B(n729), .Z(n538) );
  NANDN U748 ( .A(n536), .B(n535), .Z(n537) );
  NAND U749 ( .A(n538), .B(n537), .Z(n643) );
  AND U750 ( .A(x[1]), .B(y[12]), .Z(n540) );
  NAND U751 ( .A(x[7]), .B(y[6]), .Z(n539) );
  XNOR U752 ( .A(n540), .B(n539), .Z(n634) );
  AND U753 ( .A(o[12]), .B(n541), .Z(n633) );
  XOR U754 ( .A(n634), .B(n633), .Z(n641) );
  AND U755 ( .A(x[6]), .B(y[7]), .Z(n1611) );
  NAND U756 ( .A(y[11]), .B(x[2]), .Z(n542) );
  XNOR U757 ( .A(n543), .B(n542), .Z(n646) );
  XOR U758 ( .A(n1611), .B(n646), .Z(n640) );
  XOR U759 ( .A(n641), .B(n640), .Z(n642) );
  XOR U760 ( .A(n643), .B(n642), .Z(n610) );
  NAND U761 ( .A(n545), .B(n544), .Z(n549) );
  ANDN U762 ( .B(n547), .A(n546), .Z(n548) );
  ANDN U763 ( .B(n549), .A(n548), .Z(n609) );
  XOR U764 ( .A(n610), .B(n609), .Z(n612) );
  XOR U765 ( .A(n611), .B(n612), .Z(n603) );
  XOR U766 ( .A(n604), .B(n603), .Z(n606) );
  NAND U767 ( .A(n551), .B(n550), .Z(n555) );
  NAND U768 ( .A(n553), .B(n552), .Z(n554) );
  NAND U769 ( .A(n555), .B(n554), .Z(n618) );
  NAND U770 ( .A(x[6]), .B(y[11]), .Z(n1002) );
  AND U771 ( .A(y[6]), .B(x[1]), .Z(n632) );
  NANDN U772 ( .A(n1002), .B(n632), .Z(n559) );
  NAND U773 ( .A(n557), .B(n556), .Z(n558) );
  NAND U774 ( .A(n559), .B(n558), .Z(n624) );
  AND U775 ( .A(y[12]), .B(x[12]), .Z(n1866) );
  NAND U776 ( .A(n1866), .B(n763), .Z(n563) );
  NAND U777 ( .A(n561), .B(n560), .Z(n562) );
  NAND U778 ( .A(n563), .B(n562), .Z(n622) );
  AND U779 ( .A(y[3]), .B(x[10]), .Z(n1471) );
  AND U780 ( .A(y[2]), .B(x[11]), .Z(n1432) );
  NAND U781 ( .A(x[8]), .B(y[5]), .Z(n564) );
  XNOR U782 ( .A(n1432), .B(n564), .Z(n629) );
  XOR U783 ( .A(n1471), .B(n629), .Z(n621) );
  XOR U784 ( .A(n622), .B(n621), .Z(n623) );
  XOR U785 ( .A(n624), .B(n623), .Z(n616) );
  AND U786 ( .A(y[8]), .B(x[10]), .Z(n566) );
  NAND U787 ( .A(n566), .B(n565), .Z(n569) );
  NAND U788 ( .A(n567), .B(n1201), .Z(n568) );
  NAND U789 ( .A(n569), .B(n568), .Z(n666) );
  AND U790 ( .A(y[13]), .B(x[0]), .Z(n571) );
  NAND U791 ( .A(y[0]), .B(x[13]), .Z(n570) );
  XNOR U792 ( .A(n571), .B(n570), .Z(n658) );
  AND U793 ( .A(y[1]), .B(x[12]), .Z(n651) );
  XOR U794 ( .A(o[13]), .B(n651), .Z(n657) );
  XOR U795 ( .A(n658), .B(n657), .Z(n664) );
  AND U796 ( .A(x[5]), .B(y[8]), .Z(n573) );
  NAND U797 ( .A(y[10]), .B(x[3]), .Z(n572) );
  XNOR U798 ( .A(n573), .B(n572), .Z(n653) );
  AND U799 ( .A(y[9]), .B(x[4]), .Z(n654) );
  XOR U800 ( .A(n653), .B(n654), .Z(n663) );
  XOR U801 ( .A(n664), .B(n663), .Z(n665) );
  XOR U802 ( .A(n666), .B(n665), .Z(n615) );
  XOR U803 ( .A(n616), .B(n615), .Z(n617) );
  XOR U804 ( .A(n618), .B(n617), .Z(n605) );
  XNOR U805 ( .A(n606), .B(n605), .Z(n591) );
  NAND U806 ( .A(n575), .B(n574), .Z(n579) );
  NAND U807 ( .A(n577), .B(n576), .Z(n578) );
  AND U808 ( .A(n579), .B(n578), .Z(n590) );
  XOR U809 ( .A(n591), .B(n590), .Z(n592) );
  XOR U810 ( .A(n593), .B(n592), .Z(n599) );
  NANDN U811 ( .A(n584), .B(n583), .Z(n588) );
  NAND U812 ( .A(n586), .B(n585), .Z(n587) );
  AND U813 ( .A(n588), .B(n587), .Z(n597) );
  IV U814 ( .A(n597), .Z(n596) );
  XOR U815 ( .A(n598), .B(n596), .Z(n589) );
  XNOR U816 ( .A(n599), .B(n589), .Z(N46) );
  NAND U817 ( .A(n591), .B(n590), .Z(n595) );
  NAND U818 ( .A(n593), .B(n592), .Z(n594) );
  NAND U819 ( .A(n595), .B(n594), .Z(n752) );
  IV U820 ( .A(n752), .Z(n750) );
  OR U821 ( .A(n598), .B(n596), .Z(n602) );
  ANDN U822 ( .B(n598), .A(n597), .Z(n600) );
  OR U823 ( .A(n600), .B(n599), .Z(n601) );
  AND U824 ( .A(n602), .B(n601), .Z(n751) );
  NAND U825 ( .A(n604), .B(n603), .Z(n608) );
  NAND U826 ( .A(n606), .B(n605), .Z(n607) );
  NAND U827 ( .A(n608), .B(n607), .Z(n745) );
  NAND U828 ( .A(n610), .B(n609), .Z(n614) );
  NAND U829 ( .A(n612), .B(n611), .Z(n613) );
  NAND U830 ( .A(n614), .B(n613), .Z(n744) );
  XOR U831 ( .A(n745), .B(n744), .Z(n747) );
  NAND U832 ( .A(n616), .B(n615), .Z(n620) );
  NAND U833 ( .A(n618), .B(n617), .Z(n619) );
  NAND U834 ( .A(n620), .B(n619), .Z(n673) );
  NAND U835 ( .A(n622), .B(n621), .Z(n626) );
  NAND U836 ( .A(n624), .B(n623), .Z(n625) );
  AND U837 ( .A(n626), .B(n625), .Z(n679) );
  AND U838 ( .A(y[5]), .B(x[11]), .Z(n628) );
  NAND U839 ( .A(n628), .B(n627), .Z(n631) );
  NAND U840 ( .A(n629), .B(n1471), .Z(n630) );
  NAND U841 ( .A(n631), .B(n630), .Z(n683) );
  NAND U842 ( .A(y[12]), .B(x[7]), .Z(n1216) );
  NANDN U843 ( .A(n1216), .B(n632), .Z(n636) );
  NAND U844 ( .A(n634), .B(n633), .Z(n635) );
  NAND U845 ( .A(n636), .B(n635), .Z(n682) );
  XOR U846 ( .A(n683), .B(n682), .Z(n685) );
  AND U847 ( .A(y[10]), .B(x[4]), .Z(n1103) );
  AND U848 ( .A(y[11]), .B(x[3]), .Z(n638) );
  NAND U849 ( .A(x[8]), .B(y[6]), .Z(n637) );
  XNOR U850 ( .A(n638), .B(n637), .Z(n704) );
  XOR U851 ( .A(n1000), .B(n704), .Z(n688) );
  XOR U852 ( .A(n1103), .B(n688), .Z(n690) );
  AND U853 ( .A(y[5]), .B(x[9]), .Z(n1294) );
  AND U854 ( .A(x[10]), .B(y[4]), .Z(n1334) );
  AND U855 ( .A(x[2]), .B(y[12]), .Z(n639) );
  XOR U856 ( .A(n1334), .B(n639), .Z(n730) );
  XOR U857 ( .A(n1294), .B(n730), .Z(n689) );
  XOR U858 ( .A(n690), .B(n689), .Z(n684) );
  XNOR U859 ( .A(n685), .B(n684), .Z(n677) );
  NAND U860 ( .A(n641), .B(n640), .Z(n645) );
  NAND U861 ( .A(n643), .B(n642), .Z(n644) );
  AND U862 ( .A(n645), .B(n644), .Z(n676) );
  XOR U863 ( .A(n677), .B(n676), .Z(n678) );
  XNOR U864 ( .A(n679), .B(n678), .Z(n671) );
  AND U865 ( .A(y[11]), .B(x[9]), .Z(n1214) );
  NAND U866 ( .A(n1214), .B(n729), .Z(n648) );
  NAND U867 ( .A(n646), .B(n1611), .Z(n647) );
  NAND U868 ( .A(n648), .B(n647), .Z(n716) );
  AND U869 ( .A(x[14]), .B(y[0]), .Z(n650) );
  NAND U870 ( .A(y[14]), .B(x[0]), .Z(n649) );
  XNOR U871 ( .A(n650), .B(n649), .Z(n700) );
  AND U872 ( .A(o[13]), .B(n651), .Z(n699) );
  XOR U873 ( .A(n700), .B(n699), .Z(n714) );
  AND U874 ( .A(x[12]), .B(y[2]), .Z(n1300) );
  NAND U875 ( .A(y[7]), .B(x[7]), .Z(n652) );
  XNOR U876 ( .A(n1300), .B(n652), .Z(n720) );
  NAND U877 ( .A(x[13]), .B(y[1]), .Z(n728) );
  XNOR U878 ( .A(o[14]), .B(n728), .Z(n721) );
  XOR U879 ( .A(n720), .B(n721), .Z(n713) );
  XOR U880 ( .A(n714), .B(n713), .Z(n715) );
  XNOR U881 ( .A(n716), .B(n715), .Z(n739) );
  AND U882 ( .A(y[10]), .B(x[5]), .Z(n775) );
  NAND U883 ( .A(n1459), .B(n775), .Z(n656) );
  NAND U884 ( .A(n654), .B(n653), .Z(n655) );
  AND U885 ( .A(n656), .B(n655), .Z(n710) );
  AND U886 ( .A(x[13]), .B(y[13]), .Z(n2175) );
  NAND U887 ( .A(n2175), .B(n763), .Z(n660) );
  NAND U888 ( .A(n658), .B(n657), .Z(n659) );
  NAND U889 ( .A(n660), .B(n659), .Z(n708) );
  NAND U890 ( .A(y[3]), .B(x[11]), .Z(n661) );
  XNOR U891 ( .A(n662), .B(n661), .Z(n734) );
  AND U892 ( .A(y[13]), .B(x[1]), .Z(n735) );
  XOR U893 ( .A(n734), .B(n735), .Z(n707) );
  XOR U894 ( .A(n708), .B(n707), .Z(n709) );
  XOR U895 ( .A(n710), .B(n709), .Z(n738) );
  XOR U896 ( .A(n739), .B(n738), .Z(n741) );
  NAND U897 ( .A(n664), .B(n663), .Z(n668) );
  NAND U898 ( .A(n666), .B(n665), .Z(n667) );
  AND U899 ( .A(n668), .B(n667), .Z(n740) );
  XNOR U900 ( .A(n741), .B(n740), .Z(n670) );
  XOR U901 ( .A(n671), .B(n670), .Z(n672) );
  XOR U902 ( .A(n673), .B(n672), .Z(n746) );
  XOR U903 ( .A(n747), .B(n746), .Z(n753) );
  XNOR U904 ( .A(n751), .B(n753), .Z(n669) );
  XOR U905 ( .A(n750), .B(n669), .Z(N47) );
  NAND U906 ( .A(n671), .B(n670), .Z(n675) );
  NAND U907 ( .A(n673), .B(n672), .Z(n674) );
  AND U908 ( .A(n675), .B(n674), .Z(n846) );
  NAND U909 ( .A(n677), .B(n676), .Z(n681) );
  NAND U910 ( .A(n679), .B(n678), .Z(n680) );
  NAND U911 ( .A(n681), .B(n680), .Z(n819) );
  NAND U912 ( .A(n683), .B(n682), .Z(n687) );
  NAND U913 ( .A(n685), .B(n684), .Z(n686) );
  NAND U914 ( .A(n687), .B(n686), .Z(n837) );
  NAND U915 ( .A(n1103), .B(n688), .Z(n692) );
  NAND U916 ( .A(n690), .B(n689), .Z(n691) );
  NAND U917 ( .A(n692), .B(n691), .Z(n835) );
  AND U918 ( .A(x[4]), .B(y[11]), .Z(n694) );
  NAND U919 ( .A(x[10]), .B(y[5]), .Z(n693) );
  XNOR U920 ( .A(n694), .B(n693), .Z(n770) );
  AND U921 ( .A(x[7]), .B(y[8]), .Z(n769) );
  XNOR U922 ( .A(n770), .B(n769), .Z(n777) );
  NAND U923 ( .A(x[6]), .B(y[9]), .Z(n877) );
  XNOR U924 ( .A(n877), .B(n775), .Z(n776) );
  XNOR U925 ( .A(n777), .B(n776), .Z(n812) );
  AND U926 ( .A(x[2]), .B(y[13]), .Z(n696) );
  NAND U927 ( .A(x[9]), .B(y[6]), .Z(n695) );
  XNOR U928 ( .A(n696), .B(n695), .Z(n780) );
  AND U929 ( .A(x[3]), .B(y[12]), .Z(n781) );
  XOR U930 ( .A(n780), .B(n781), .Z(n810) );
  AND U931 ( .A(y[14]), .B(x[1]), .Z(n698) );
  NAND U932 ( .A(y[7]), .B(x[8]), .Z(n697) );
  XNOR U933 ( .A(n698), .B(n697), .Z(n759) );
  NAND U934 ( .A(y[1]), .B(x[14]), .Z(n786) );
  XOR U935 ( .A(o[15]), .B(n786), .Z(n760) );
  XNOR U936 ( .A(n759), .B(n760), .Z(n811) );
  XOR U937 ( .A(n810), .B(n811), .Z(n813) );
  XOR U938 ( .A(n812), .B(n813), .Z(n792) );
  AND U939 ( .A(x[14]), .B(y[14]), .Z(n2437) );
  NAND U940 ( .A(n2437), .B(n763), .Z(n702) );
  NAND U941 ( .A(n700), .B(n699), .Z(n701) );
  NAND U942 ( .A(n702), .B(n701), .Z(n790) );
  AND U943 ( .A(x[8]), .B(y[11]), .Z(n1079) );
  NAND U944 ( .A(n703), .B(n1079), .Z(n706) );
  NAND U945 ( .A(n704), .B(n1000), .Z(n705) );
  NAND U946 ( .A(n706), .B(n705), .Z(n789) );
  XOR U947 ( .A(n790), .B(n789), .Z(n791) );
  XOR U948 ( .A(n792), .B(n791), .Z(n834) );
  XOR U949 ( .A(n835), .B(n834), .Z(n836) );
  XNOR U950 ( .A(n837), .B(n836), .Z(n817) );
  NAND U951 ( .A(n708), .B(n707), .Z(n712) );
  NANDN U952 ( .A(n710), .B(n709), .Z(n711) );
  AND U953 ( .A(n712), .B(n711), .Z(n825) );
  NAND U954 ( .A(n714), .B(n713), .Z(n718) );
  NAND U955 ( .A(n716), .B(n715), .Z(n717) );
  NAND U956 ( .A(n718), .B(n717), .Z(n823) );
  NAND U957 ( .A(y[7]), .B(x[12]), .Z(n1208) );
  NANDN U958 ( .A(n1208), .B(n719), .Z(n723) );
  NAND U959 ( .A(n721), .B(n720), .Z(n722) );
  AND U960 ( .A(n723), .B(n722), .Z(n798) );
  AND U961 ( .A(y[4]), .B(x[11]), .Z(n725) );
  NAND U962 ( .A(y[2]), .B(x[13]), .Z(n724) );
  XNOR U963 ( .A(n725), .B(n724), .Z(n803) );
  AND U964 ( .A(y[3]), .B(x[12]), .Z(n802) );
  XNOR U965 ( .A(n803), .B(n802), .Z(n796) );
  AND U966 ( .A(x[15]), .B(y[0]), .Z(n727) );
  NAND U967 ( .A(y[15]), .B(x[0]), .Z(n726) );
  XNOR U968 ( .A(n727), .B(n726), .Z(n765) );
  ANDN U969 ( .B(o[14]), .A(n728), .Z(n764) );
  XNOR U970 ( .A(n765), .B(n764), .Z(n795) );
  XOR U971 ( .A(n796), .B(n795), .Z(n797) );
  XNOR U972 ( .A(n798), .B(n797), .Z(n831) );
  NAND U973 ( .A(y[12]), .B(x[10]), .Z(n1613) );
  NANDN U974 ( .A(n1613), .B(n729), .Z(n732) );
  NAND U975 ( .A(n1294), .B(n730), .Z(n731) );
  NAND U976 ( .A(n732), .B(n731), .Z(n829) );
  AND U977 ( .A(x[11]), .B(y[8]), .Z(n1102) );
  AND U978 ( .A(x[6]), .B(y[3]), .Z(n733) );
  NAND U979 ( .A(n1102), .B(n733), .Z(n737) );
  NAND U980 ( .A(n735), .B(n734), .Z(n736) );
  NAND U981 ( .A(n737), .B(n736), .Z(n828) );
  XOR U982 ( .A(n829), .B(n828), .Z(n830) );
  XOR U983 ( .A(n831), .B(n830), .Z(n822) );
  XOR U984 ( .A(n823), .B(n822), .Z(n824) );
  XOR U985 ( .A(n825), .B(n824), .Z(n816) );
  XOR U986 ( .A(n817), .B(n816), .Z(n818) );
  XNOR U987 ( .A(n819), .B(n818), .Z(n843) );
  NAND U988 ( .A(n739), .B(n738), .Z(n743) );
  NAND U989 ( .A(n741), .B(n740), .Z(n742) );
  AND U990 ( .A(n743), .B(n742), .Z(n844) );
  XOR U991 ( .A(n843), .B(n844), .Z(n845) );
  XOR U992 ( .A(n846), .B(n845), .Z(n842) );
  NAND U993 ( .A(n745), .B(n744), .Z(n749) );
  NAND U994 ( .A(n747), .B(n746), .Z(n748) );
  NAND U995 ( .A(n749), .B(n748), .Z(n841) );
  NANDN U996 ( .A(n750), .B(n751), .Z(n756) );
  NOR U997 ( .A(n752), .B(n751), .Z(n754) );
  OR U998 ( .A(n754), .B(n753), .Z(n755) );
  AND U999 ( .A(n756), .B(n755), .Z(n840) );
  XOR U1000 ( .A(n841), .B(n840), .Z(n757) );
  XNOR U1001 ( .A(n842), .B(n757), .Z(N48) );
  AND U1002 ( .A(x[8]), .B(y[14]), .Z(n1104) );
  NAND U1003 ( .A(n1104), .B(n758), .Z(n762) );
  NANDN U1004 ( .A(n760), .B(n759), .Z(n761) );
  AND U1005 ( .A(n762), .B(n761), .Z(n905) );
  AND U1006 ( .A(y[15]), .B(x[15]), .Z(n2886) );
  NAND U1007 ( .A(n2886), .B(n763), .Z(n767) );
  NAND U1008 ( .A(n765), .B(n764), .Z(n766) );
  NAND U1009 ( .A(n767), .B(n766), .Z(n904) );
  XNOR U1010 ( .A(n905), .B(n904), .Z(n907) );
  AND U1011 ( .A(y[11]), .B(x[10]), .Z(n1347) );
  NAND U1012 ( .A(n1347), .B(n768), .Z(n772) );
  NAND U1013 ( .A(n770), .B(n769), .Z(n771) );
  NAND U1014 ( .A(n772), .B(n771), .Z(n864) );
  AND U1015 ( .A(y[16]), .B(x[0]), .Z(n884) );
  NAND U1016 ( .A(y[0]), .B(x[16]), .Z(n885) );
  XNOR U1017 ( .A(n884), .B(n885), .Z(n886) );
  NAND U1018 ( .A(y[1]), .B(x[15]), .Z(n874) );
  XOR U1019 ( .A(o[16]), .B(n874), .Z(n887) );
  XNOR U1020 ( .A(n886), .B(n887), .Z(n863) );
  AND U1021 ( .A(y[9]), .B(x[7]), .Z(n774) );
  NAND U1022 ( .A(x[6]), .B(y[10]), .Z(n773) );
  XNOR U1023 ( .A(n774), .B(n773), .Z(n879) );
  AND U1024 ( .A(y[6]), .B(x[10]), .Z(n878) );
  XOR U1025 ( .A(n879), .B(n878), .Z(n862) );
  XOR U1026 ( .A(n863), .B(n862), .Z(n865) );
  XOR U1027 ( .A(n864), .B(n865), .Z(n906) );
  XNOR U1028 ( .A(n907), .B(n906), .Z(n859) );
  NANDN U1029 ( .A(n775), .B(n877), .Z(n779) );
  NAND U1030 ( .A(n777), .B(n776), .Z(n778) );
  NAND U1031 ( .A(n779), .B(n778), .Z(n857) );
  AND U1032 ( .A(y[13]), .B(x[9]), .Z(n1582) );
  NAND U1033 ( .A(n1582), .B(n1206), .Z(n783) );
  NAND U1034 ( .A(n781), .B(n780), .Z(n782) );
  AND U1035 ( .A(n783), .B(n782), .Z(n895) );
  AND U1036 ( .A(x[1]), .B(y[15]), .Z(n785) );
  NAND U1037 ( .A(y[8]), .B(x[8]), .Z(n784) );
  XNOR U1038 ( .A(n785), .B(n784), .Z(n883) );
  ANDN U1039 ( .B(o[15]), .A(n786), .Z(n882) );
  XOR U1040 ( .A(n883), .B(n882), .Z(n892) );
  AND U1041 ( .A(y[2]), .B(x[14]), .Z(n788) );
  NAND U1042 ( .A(x[11]), .B(y[5]), .Z(n787) );
  XNOR U1043 ( .A(n788), .B(n787), .Z(n916) );
  NAND U1044 ( .A(y[12]), .B(x[4]), .Z(n917) );
  XNOR U1045 ( .A(n916), .B(n917), .Z(n893) );
  XOR U1046 ( .A(n892), .B(n893), .Z(n894) );
  XOR U1047 ( .A(n895), .B(n894), .Z(n856) );
  XOR U1048 ( .A(n857), .B(n856), .Z(n858) );
  XOR U1049 ( .A(n859), .B(n858), .Z(n898) );
  NAND U1050 ( .A(n790), .B(n789), .Z(n794) );
  NAND U1051 ( .A(n792), .B(n791), .Z(n793) );
  AND U1052 ( .A(n794), .B(n793), .Z(n899) );
  XOR U1053 ( .A(n898), .B(n899), .Z(n901) );
  NAND U1054 ( .A(n796), .B(n795), .Z(n800) );
  NAND U1055 ( .A(n798), .B(n797), .Z(n799) );
  NAND U1056 ( .A(n800), .B(n799), .Z(n931) );
  AND U1057 ( .A(x[13]), .B(y[4]), .Z(n801) );
  NAND U1058 ( .A(n1432), .B(n801), .Z(n805) );
  NAND U1059 ( .A(n803), .B(n802), .Z(n804) );
  AND U1060 ( .A(n805), .B(n804), .Z(n912) );
  AND U1061 ( .A(x[9]), .B(y[7]), .Z(n807) );
  NAND U1062 ( .A(y[14]), .B(x[2]), .Z(n806) );
  XNOR U1063 ( .A(n807), .B(n806), .Z(n920) );
  NAND U1064 ( .A(x[3]), .B(y[13]), .Z(n921) );
  XNOR U1065 ( .A(n920), .B(n921), .Z(n910) );
  AND U1066 ( .A(y[4]), .B(x[12]), .Z(n1588) );
  AND U1067 ( .A(x[5]), .B(y[11]), .Z(n809) );
  NAND U1068 ( .A(y[3]), .B(x[13]), .Z(n808) );
  XOR U1069 ( .A(n809), .B(n808), .Z(n869) );
  XOR U1070 ( .A(n1588), .B(n869), .Z(n911) );
  XOR U1071 ( .A(n910), .B(n911), .Z(n913) );
  XNOR U1072 ( .A(n912), .B(n913), .Z(n929) );
  NAND U1073 ( .A(n811), .B(n810), .Z(n815) );
  NAND U1074 ( .A(n813), .B(n812), .Z(n814) );
  AND U1075 ( .A(n815), .B(n814), .Z(n928) );
  XOR U1076 ( .A(n929), .B(n928), .Z(n930) );
  XOR U1077 ( .A(n931), .B(n930), .Z(n900) );
  XNOR U1078 ( .A(n901), .B(n900), .Z(n935) );
  NAND U1079 ( .A(n817), .B(n816), .Z(n821) );
  NAND U1080 ( .A(n819), .B(n818), .Z(n820) );
  AND U1081 ( .A(n821), .B(n820), .Z(n934) );
  XOR U1082 ( .A(n935), .B(n934), .Z(n937) );
  NAND U1083 ( .A(n823), .B(n822), .Z(n827) );
  NANDN U1084 ( .A(n825), .B(n824), .Z(n826) );
  NAND U1085 ( .A(n827), .B(n826), .Z(n853) );
  NAND U1086 ( .A(n829), .B(n828), .Z(n833) );
  NAND U1087 ( .A(n831), .B(n830), .Z(n832) );
  NAND U1088 ( .A(n833), .B(n832), .Z(n850) );
  NAND U1089 ( .A(n835), .B(n834), .Z(n839) );
  NAND U1090 ( .A(n837), .B(n836), .Z(n838) );
  NAND U1091 ( .A(n839), .B(n838), .Z(n851) );
  XOR U1092 ( .A(n850), .B(n851), .Z(n852) );
  XOR U1093 ( .A(n853), .B(n852), .Z(n936) );
  XOR U1094 ( .A(n937), .B(n936), .Z(n943) );
  NAND U1095 ( .A(n844), .B(n843), .Z(n848) );
  NANDN U1096 ( .A(n846), .B(n845), .Z(n847) );
  AND U1097 ( .A(n848), .B(n847), .Z(n942) );
  IV U1098 ( .A(n942), .Z(n940) );
  XOR U1099 ( .A(n941), .B(n940), .Z(n849) );
  XNOR U1100 ( .A(n943), .B(n849), .Z(N49) );
  NAND U1101 ( .A(n851), .B(n850), .Z(n855) );
  NAND U1102 ( .A(n853), .B(n852), .Z(n854) );
  AND U1103 ( .A(n855), .B(n854), .Z(n1042) );
  NAND U1104 ( .A(n857), .B(n856), .Z(n861) );
  NAND U1105 ( .A(n859), .B(n858), .Z(n860) );
  NAND U1106 ( .A(n861), .B(n860), .Z(n957) );
  NAND U1107 ( .A(n863), .B(n862), .Z(n867) );
  NAND U1108 ( .A(n865), .B(n864), .Z(n866) );
  AND U1109 ( .A(n867), .B(n866), .Z(n1032) );
  AND U1110 ( .A(x[13]), .B(y[11]), .Z(n1874) );
  AND U1111 ( .A(x[5]), .B(y[3]), .Z(n868) );
  NAND U1112 ( .A(n1874), .B(n868), .Z(n871) );
  NANDN U1113 ( .A(n869), .B(n1588), .Z(n870) );
  AND U1114 ( .A(n871), .B(n870), .Z(n989) );
  AND U1115 ( .A(x[9]), .B(y[8]), .Z(n873) );
  NAND U1116 ( .A(x[1]), .B(y[16]), .Z(n872) );
  XNOR U1117 ( .A(n873), .B(n872), .Z(n1006) );
  ANDN U1118 ( .B(o[16]), .A(n874), .Z(n1005) );
  XOR U1119 ( .A(n1006), .B(n1005), .Z(n987) );
  AND U1120 ( .A(x[15]), .B(y[2]), .Z(n876) );
  NAND U1121 ( .A(x[12]), .B(y[5]), .Z(n875) );
  XNOR U1122 ( .A(n876), .B(n875), .Z(n962) );
  AND U1123 ( .A(x[14]), .B(y[3]), .Z(n961) );
  XOR U1124 ( .A(n962), .B(n961), .Z(n986) );
  XOR U1125 ( .A(n987), .B(n986), .Z(n988) );
  XNOR U1126 ( .A(n989), .B(n988), .Z(n1030) );
  AND U1127 ( .A(y[10]), .B(x[7]), .Z(n1015) );
  NANDN U1128 ( .A(n877), .B(n1015), .Z(n881) );
  NAND U1129 ( .A(n879), .B(n878), .Z(n880) );
  AND U1130 ( .A(n881), .B(n880), .Z(n995) );
  NAND U1131 ( .A(x[8]), .B(y[15]), .Z(n1686) );
  XNOR U1132 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U1133 ( .A(n885), .B(n884), .Z(n889) );
  NANDN U1134 ( .A(n887), .B(n886), .Z(n888) );
  AND U1135 ( .A(n889), .B(n888), .Z(n993) );
  AND U1136 ( .A(x[0]), .B(y[17]), .Z(n976) );
  AND U1137 ( .A(x[17]), .B(y[0]), .Z(n975) );
  XOR U1138 ( .A(n976), .B(n975), .Z(n978) );
  AND U1139 ( .A(y[1]), .B(x[16]), .Z(n972) );
  XOR U1140 ( .A(n972), .B(o[17]), .Z(n977) );
  XOR U1141 ( .A(n978), .B(n977), .Z(n991) );
  AND U1142 ( .A(x[10]), .B(y[7]), .Z(n891) );
  NAND U1143 ( .A(y[15]), .B(x[2]), .Z(n890) );
  XNOR U1144 ( .A(n891), .B(n890), .Z(n1011) );
  AND U1145 ( .A(x[3]), .B(y[14]), .Z(n1010) );
  XOR U1146 ( .A(n1011), .B(n1010), .Z(n990) );
  XOR U1147 ( .A(n991), .B(n990), .Z(n992) );
  XOR U1148 ( .A(n993), .B(n992), .Z(n997) );
  XOR U1149 ( .A(n996), .B(n997), .Z(n1031) );
  XOR U1150 ( .A(n1030), .B(n1031), .Z(n1033) );
  XNOR U1151 ( .A(n1032), .B(n1033), .Z(n955) );
  NAND U1152 ( .A(n893), .B(n892), .Z(n897) );
  NANDN U1153 ( .A(n895), .B(n894), .Z(n896) );
  AND U1154 ( .A(n897), .B(n896), .Z(n954) );
  XOR U1155 ( .A(n955), .B(n954), .Z(n956) );
  XNOR U1156 ( .A(n957), .B(n956), .Z(n1040) );
  NAND U1157 ( .A(n899), .B(n898), .Z(n903) );
  NAND U1158 ( .A(n901), .B(n900), .Z(n902) );
  AND U1159 ( .A(n903), .B(n902), .Z(n951) );
  NANDN U1160 ( .A(n905), .B(n904), .Z(n909) );
  NAND U1161 ( .A(n907), .B(n906), .Z(n908) );
  AND U1162 ( .A(n909), .B(n908), .Z(n1026) );
  NANDN U1163 ( .A(n911), .B(n910), .Z(n915) );
  OR U1164 ( .A(n913), .B(n912), .Z(n914) );
  AND U1165 ( .A(n915), .B(n914), .Z(n1025) );
  NAND U1166 ( .A(y[5]), .B(x[14]), .Z(n1240) );
  NANDN U1167 ( .A(n1240), .B(n1432), .Z(n919) );
  NANDN U1168 ( .A(n917), .B(n916), .Z(n918) );
  AND U1169 ( .A(n919), .B(n918), .Z(n1019) );
  AND U1170 ( .A(x[9]), .B(y[14]), .Z(n1855) );
  NANDN U1171 ( .A(n1009), .B(n1855), .Z(n923) );
  NANDN U1172 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1173 ( .A(n923), .B(n922), .Z(n1018) );
  XNOR U1174 ( .A(n1019), .B(n1018), .Z(n1020) );
  AND U1175 ( .A(y[9]), .B(x[8]), .Z(n925) );
  NAND U1176 ( .A(x[5]), .B(y[12]), .Z(n924) );
  XNOR U1177 ( .A(n925), .B(n924), .Z(n1001) );
  XOR U1178 ( .A(n1015), .B(n1014), .Z(n1016) );
  AND U1179 ( .A(x[4]), .B(y[13]), .Z(n927) );
  NAND U1180 ( .A(y[4]), .B(x[13]), .Z(n926) );
  XNOR U1181 ( .A(n927), .B(n926), .Z(n966) );
  NAND U1182 ( .A(y[6]), .B(x[11]), .Z(n967) );
  XOR U1183 ( .A(n966), .B(n967), .Z(n1017) );
  XOR U1184 ( .A(n1016), .B(n1017), .Z(n1021) );
  XNOR U1185 ( .A(n1020), .B(n1021), .Z(n1024) );
  XOR U1186 ( .A(n1025), .B(n1024), .Z(n1027) );
  XNOR U1187 ( .A(n1026), .B(n1027), .Z(n949) );
  NAND U1188 ( .A(n929), .B(n928), .Z(n933) );
  NAND U1189 ( .A(n931), .B(n930), .Z(n932) );
  NAND U1190 ( .A(n933), .B(n932), .Z(n948) );
  XOR U1191 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1192 ( .A(n951), .B(n950), .Z(n1039) );
  XOR U1193 ( .A(n1040), .B(n1039), .Z(n1041) );
  XOR U1194 ( .A(n1042), .B(n1041), .Z(n1038) );
  NAND U1195 ( .A(n935), .B(n934), .Z(n939) );
  NAND U1196 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1197 ( .A(n939), .B(n938), .Z(n1037) );
  NANDN U1198 ( .A(n940), .B(n941), .Z(n946) );
  NOR U1199 ( .A(n942), .B(n941), .Z(n944) );
  OR U1200 ( .A(n944), .B(n943), .Z(n945) );
  AND U1201 ( .A(n946), .B(n945), .Z(n1036) );
  XOR U1202 ( .A(n1037), .B(n1036), .Z(n947) );
  XNOR U1203 ( .A(n1038), .B(n947), .Z(N50) );
  NAND U1204 ( .A(n949), .B(n948), .Z(n953) );
  NANDN U1205 ( .A(n951), .B(n950), .Z(n952) );
  AND U1206 ( .A(n953), .B(n952), .Z(n1151) );
  NAND U1207 ( .A(n955), .B(n954), .Z(n959) );
  NAND U1208 ( .A(n957), .B(n956), .Z(n958) );
  AND U1209 ( .A(n959), .B(n958), .Z(n1148) );
  AND U1210 ( .A(y[5]), .B(x[15]), .Z(n960) );
  NAND U1211 ( .A(n960), .B(n1300), .Z(n964) );
  NAND U1212 ( .A(n962), .B(n961), .Z(n963) );
  NAND U1213 ( .A(n964), .B(n963), .Z(n1130) );
  NAND U1214 ( .A(n2175), .B(n965), .Z(n969) );
  NANDN U1215 ( .A(n967), .B(n966), .Z(n968) );
  NAND U1216 ( .A(n969), .B(n968), .Z(n1120) );
  AND U1217 ( .A(x[1]), .B(y[17]), .Z(n971) );
  NAND U1218 ( .A(x[10]), .B(y[8]), .Z(n970) );
  XNOR U1219 ( .A(n971), .B(n970), .Z(n1083) );
  NAND U1220 ( .A(n972), .B(o[17]), .Z(n1084) );
  AND U1221 ( .A(x[15]), .B(y[3]), .Z(n974) );
  NAND U1222 ( .A(x[9]), .B(y[9]), .Z(n973) );
  XNOR U1223 ( .A(n974), .B(n973), .Z(n1075) );
  AND U1224 ( .A(x[14]), .B(y[4]), .Z(n1074) );
  XOR U1225 ( .A(n1075), .B(n1074), .Z(n1118) );
  XOR U1226 ( .A(n1119), .B(n1118), .Z(n1121) );
  XOR U1227 ( .A(n1120), .B(n1121), .Z(n1131) );
  XOR U1228 ( .A(n1130), .B(n1131), .Z(n1133) );
  NAND U1229 ( .A(n976), .B(n975), .Z(n980) );
  NAND U1230 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1231 ( .A(n980), .B(n979), .Z(n1142) );
  AND U1232 ( .A(y[2]), .B(x[16]), .Z(n982) );
  NAND U1233 ( .A(y[7]), .B(x[11]), .Z(n981) );
  XNOR U1234 ( .A(n982), .B(n981), .Z(n1071) );
  AND U1235 ( .A(y[16]), .B(x[2]), .Z(n1070) );
  XOR U1236 ( .A(n1071), .B(n1070), .Z(n1143) );
  XOR U1237 ( .A(n1142), .B(n1143), .Z(n1145) );
  AND U1238 ( .A(x[5]), .B(y[13]), .Z(n1222) );
  NAND U1239 ( .A(x[6]), .B(y[12]), .Z(n983) );
  XNOR U1240 ( .A(n1222), .B(n983), .Z(n1067) );
  AND U1241 ( .A(x[4]), .B(y[14]), .Z(n985) );
  NAND U1242 ( .A(x[8]), .B(y[10]), .Z(n984) );
  XNOR U1243 ( .A(n985), .B(n984), .Z(n1105) );
  AND U1244 ( .A(x[7]), .B(y[11]), .Z(n1106) );
  XOR U1245 ( .A(n1105), .B(n1106), .Z(n1066) );
  XOR U1246 ( .A(n1067), .B(n1066), .Z(n1144) );
  XOR U1247 ( .A(n1145), .B(n1144), .Z(n1132) );
  XOR U1248 ( .A(n1133), .B(n1132), .Z(n1053) );
  XOR U1249 ( .A(n1125), .B(n1124), .Z(n1127) );
  NANDN U1250 ( .A(n995), .B(n994), .Z(n999) );
  NANDN U1251 ( .A(n997), .B(n996), .Z(n998) );
  AND U1252 ( .A(n999), .B(n998), .Z(n1126) );
  XOR U1253 ( .A(n1127), .B(n1126), .Z(n1052) );
  XNOR U1254 ( .A(n1053), .B(n1052), .Z(n1055) );
  AND U1255 ( .A(y[12]), .B(x[8]), .Z(n1340) );
  NAND U1256 ( .A(n1340), .B(n1000), .Z(n1004) );
  NANDN U1257 ( .A(n1002), .B(n1001), .Z(n1003) );
  NAND U1258 ( .A(n1004), .B(n1003), .Z(n1137) );
  NAND U1259 ( .A(y[16]), .B(x[9]), .Z(n1962) );
  NANDN U1260 ( .A(n1962), .B(n1082), .Z(n1008) );
  NAND U1261 ( .A(n1006), .B(n1005), .Z(n1007) );
  NAND U1262 ( .A(n1008), .B(n1007), .Z(n1136) );
  XOR U1263 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U1264 ( .A(y[15]), .B(x[10]), .Z(n1963) );
  AND U1265 ( .A(y[18]), .B(x[0]), .Z(n1087) );
  NAND U1266 ( .A(y[0]), .B(x[18]), .Z(n1088) );
  AND U1267 ( .A(x[17]), .B(y[1]), .Z(n1109) );
  XOR U1268 ( .A(o[18]), .B(n1109), .Z(n1089) );
  XOR U1269 ( .A(n1090), .B(n1089), .Z(n1113) );
  AND U1270 ( .A(y[15]), .B(x[3]), .Z(n1013) );
  NAND U1271 ( .A(y[5]), .B(x[13]), .Z(n1012) );
  XNOR U1272 ( .A(n1013), .B(n1012), .Z(n1095) );
  NAND U1273 ( .A(y[6]), .B(x[12]), .Z(n1096) );
  XOR U1274 ( .A(n1113), .B(n1112), .Z(n1115) );
  XNOR U1275 ( .A(n1114), .B(n1115), .Z(n1139) );
  XOR U1276 ( .A(n1059), .B(n1058), .Z(n1061) );
  NANDN U1277 ( .A(n1019), .B(n1018), .Z(n1023) );
  NANDN U1278 ( .A(n1021), .B(n1020), .Z(n1022) );
  AND U1279 ( .A(n1023), .B(n1022), .Z(n1060) );
  XOR U1280 ( .A(n1061), .B(n1060), .Z(n1054) );
  XOR U1281 ( .A(n1055), .B(n1054), .Z(n1049) );
  NANDN U1282 ( .A(n1025), .B(n1024), .Z(n1029) );
  OR U1283 ( .A(n1027), .B(n1026), .Z(n1028) );
  AND U1284 ( .A(n1029), .B(n1028), .Z(n1047) );
  NANDN U1285 ( .A(n1031), .B(n1030), .Z(n1035) );
  OR U1286 ( .A(n1033), .B(n1032), .Z(n1034) );
  NAND U1287 ( .A(n1035), .B(n1034), .Z(n1046) );
  XNOR U1288 ( .A(n1047), .B(n1046), .Z(n1048) );
  XNOR U1289 ( .A(n1049), .B(n1048), .Z(n1149) );
  XOR U1290 ( .A(n1148), .B(n1149), .Z(n1150) );
  XOR U1291 ( .A(n1151), .B(n1150), .Z(n1157) );
  NAND U1292 ( .A(n1040), .B(n1039), .Z(n1044) );
  NANDN U1293 ( .A(n1042), .B(n1041), .Z(n1043) );
  AND U1294 ( .A(n1044), .B(n1043), .Z(n1156) );
  IV U1295 ( .A(n1156), .Z(n1154) );
  XOR U1296 ( .A(n1155), .B(n1154), .Z(n1045) );
  XNOR U1297 ( .A(n1157), .B(n1045), .Z(N51) );
  NANDN U1298 ( .A(n1047), .B(n1046), .Z(n1051) );
  NANDN U1299 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1300 ( .A(n1051), .B(n1050), .Z(n1165) );
  NANDN U1301 ( .A(n1053), .B(n1052), .Z(n1057) );
  NAND U1302 ( .A(n1055), .B(n1054), .Z(n1056) );
  AND U1303 ( .A(n1057), .B(n1056), .Z(n1162) );
  NAND U1304 ( .A(n1059), .B(n1058), .Z(n1063) );
  NAND U1305 ( .A(n1061), .B(n1060), .Z(n1062) );
  NAND U1306 ( .A(n1063), .B(n1062), .Z(n1262) );
  AND U1307 ( .A(x[6]), .B(y[13]), .Z(n1065) );
  AND U1308 ( .A(y[12]), .B(x[5]), .Z(n1064) );
  NAND U1309 ( .A(n1065), .B(n1064), .Z(n1069) );
  NAND U1310 ( .A(n1067), .B(n1066), .Z(n1068) );
  NAND U1311 ( .A(n1069), .B(n1068), .Z(n1173) );
  AND U1312 ( .A(x[16]), .B(y[7]), .Z(n1587) );
  NAND U1313 ( .A(n1587), .B(n1432), .Z(n1073) );
  NAND U1314 ( .A(n1071), .B(n1070), .Z(n1072) );
  NAND U1315 ( .A(n1073), .B(n1072), .Z(n1171) );
  AND U1316 ( .A(y[9]), .B(x[15]), .Z(n1887) );
  NAND U1317 ( .A(n1887), .B(n1201), .Z(n1077) );
  NAND U1318 ( .A(n1075), .B(n1074), .Z(n1076) );
  AND U1319 ( .A(n1077), .B(n1076), .Z(n1192) );
  NAND U1320 ( .A(x[1]), .B(y[18]), .Z(n1078) );
  XNOR U1321 ( .A(n1079), .B(n1078), .Z(n1239) );
  AND U1322 ( .A(y[17]), .B(x[2]), .Z(n1081) );
  NAND U1323 ( .A(y[6]), .B(x[13]), .Z(n1080) );
  XNOR U1324 ( .A(n1081), .B(n1080), .Z(n1207) );
  XOR U1325 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U1326 ( .A(n1171), .B(n1172), .Z(n1174) );
  XNOR U1327 ( .A(n1173), .B(n1174), .Z(n1261) );
  AND U1328 ( .A(y[17]), .B(x[10]), .Z(n2326) );
  IV U1329 ( .A(n2326), .Z(n2146) );
  NANDN U1330 ( .A(n2146), .B(n1082), .Z(n1086) );
  NANDN U1331 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U1332 ( .A(n1086), .B(n1085), .Z(n1251) );
  NANDN U1333 ( .A(n1088), .B(n1087), .Z(n1092) );
  NAND U1334 ( .A(n1090), .B(n1089), .Z(n1091) );
  AND U1335 ( .A(n1092), .B(n1091), .Z(n1249) );
  AND U1336 ( .A(y[3]), .B(x[16]), .Z(n1826) );
  NAND U1337 ( .A(x[9]), .B(y[10]), .Z(n1093) );
  XNOR U1338 ( .A(n1826), .B(n1093), .Z(n1202) );
  AND U1339 ( .A(y[4]), .B(x[15]), .Z(n1203) );
  XOR U1340 ( .A(n1202), .B(n1203), .Z(n1248) );
  AND U1341 ( .A(x[13]), .B(y[15]), .Z(n2467) );
  NANDN U1342 ( .A(n1094), .B(n2467), .Z(n1098) );
  NANDN U1343 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1344 ( .A(n1098), .B(n1097), .Z(n1257) );
  AND U1345 ( .A(x[10]), .B(y[9]), .Z(n1100) );
  NAND U1346 ( .A(y[2]), .B(x[17]), .Z(n1099) );
  XNOR U1347 ( .A(n1100), .B(n1099), .Z(n1245) );
  AND U1348 ( .A(y[1]), .B(x[18]), .Z(n1221) );
  XOR U1349 ( .A(o[19]), .B(n1221), .Z(n1244) );
  XOR U1350 ( .A(n1245), .B(n1244), .Z(n1255) );
  NAND U1351 ( .A(x[3]), .B(y[16]), .Z(n1101) );
  XNOR U1352 ( .A(n1102), .B(n1101), .Z(n1215) );
  XOR U1353 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U1354 ( .A(n1104), .B(n1103), .Z(n1108) );
  NAND U1355 ( .A(n1106), .B(n1105), .Z(n1107) );
  AND U1356 ( .A(n1108), .B(n1107), .Z(n1198) );
  AND U1357 ( .A(x[0]), .B(y[19]), .Z(n1226) );
  AND U1358 ( .A(y[0]), .B(x[19]), .Z(n1227) );
  XOR U1359 ( .A(n1226), .B(n1227), .Z(n1229) );
  AND U1360 ( .A(o[18]), .B(n1109), .Z(n1228) );
  XOR U1361 ( .A(n1229), .B(n1228), .Z(n1196) );
  AND U1362 ( .A(y[15]), .B(x[4]), .Z(n1354) );
  AND U1363 ( .A(y[14]), .B(x[5]), .Z(n1111) );
  NAND U1364 ( .A(y[13]), .B(x[6]), .Z(n1110) );
  XNOR U1365 ( .A(n1111), .B(n1110), .Z(n1223) );
  XOR U1366 ( .A(n1354), .B(n1223), .Z(n1195) );
  XOR U1367 ( .A(n1196), .B(n1195), .Z(n1197) );
  XOR U1368 ( .A(n1198), .B(n1197), .Z(n1177) );
  XNOR U1369 ( .A(n1180), .B(n1179), .Z(n1185) );
  NAND U1370 ( .A(n1113), .B(n1112), .Z(n1117) );
  NAND U1371 ( .A(n1115), .B(n1114), .Z(n1116) );
  NAND U1372 ( .A(n1117), .B(n1116), .Z(n1184) );
  NAND U1373 ( .A(n1119), .B(n1118), .Z(n1123) );
  NAND U1374 ( .A(n1121), .B(n1120), .Z(n1122) );
  NAND U1375 ( .A(n1123), .B(n1122), .Z(n1183) );
  XNOR U1376 ( .A(n1184), .B(n1183), .Z(n1186) );
  XOR U1377 ( .A(n1185), .B(n1186), .Z(n1260) );
  XOR U1378 ( .A(n1261), .B(n1260), .Z(n1263) );
  XOR U1379 ( .A(n1262), .B(n1263), .Z(n1275) );
  NAND U1380 ( .A(n1125), .B(n1124), .Z(n1129) );
  NAND U1381 ( .A(n1127), .B(n1126), .Z(n1128) );
  AND U1382 ( .A(n1129), .B(n1128), .Z(n1272) );
  NAND U1383 ( .A(n1131), .B(n1130), .Z(n1135) );
  NAND U1384 ( .A(n1133), .B(n1132), .Z(n1134) );
  NAND U1385 ( .A(n1135), .B(n1134), .Z(n1268) );
  NAND U1386 ( .A(n1137), .B(n1136), .Z(n1141) );
  NANDN U1387 ( .A(n1139), .B(n1138), .Z(n1140) );
  NAND U1388 ( .A(n1141), .B(n1140), .Z(n1267) );
  NAND U1389 ( .A(n1143), .B(n1142), .Z(n1147) );
  NAND U1390 ( .A(n1145), .B(n1144), .Z(n1146) );
  NAND U1391 ( .A(n1147), .B(n1146), .Z(n1266) );
  XNOR U1392 ( .A(n1267), .B(n1266), .Z(n1269) );
  XNOR U1393 ( .A(n1272), .B(n1273), .Z(n1274) );
  XNOR U1394 ( .A(n1162), .B(n1163), .Z(n1164) );
  XOR U1395 ( .A(n1165), .B(n1164), .Z(n1170) );
  NAND U1396 ( .A(n1149), .B(n1148), .Z(n1153) );
  NAND U1397 ( .A(n1151), .B(n1150), .Z(n1152) );
  NAND U1398 ( .A(n1153), .B(n1152), .Z(n1169) );
  NANDN U1399 ( .A(n1154), .B(n1155), .Z(n1160) );
  NOR U1400 ( .A(n1156), .B(n1155), .Z(n1158) );
  OR U1401 ( .A(n1158), .B(n1157), .Z(n1159) );
  AND U1402 ( .A(n1160), .B(n1159), .Z(n1168) );
  XOR U1403 ( .A(n1169), .B(n1168), .Z(n1161) );
  XNOR U1404 ( .A(n1170), .B(n1161), .Z(N52) );
  NANDN U1405 ( .A(n1163), .B(n1162), .Z(n1167) );
  NANDN U1406 ( .A(n1165), .B(n1164), .Z(n1166) );
  AND U1407 ( .A(n1167), .B(n1166), .Z(n1287) );
  NAND U1408 ( .A(n1172), .B(n1171), .Z(n1176) );
  NAND U1409 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U1410 ( .A(n1176), .B(n1175), .Z(n1397) );
  NANDN U1411 ( .A(n1178), .B(n1177), .Z(n1182) );
  NAND U1412 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U1413 ( .A(n1182), .B(n1181), .Z(n1395) );
  NAND U1414 ( .A(n1184), .B(n1183), .Z(n1188) );
  NANDN U1415 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1416 ( .A(n1188), .B(n1187), .Z(n1396) );
  XOR U1417 ( .A(n1395), .B(n1396), .Z(n1398) );
  XNOR U1418 ( .A(n1397), .B(n1398), .Z(n1390) );
  NAND U1419 ( .A(n1190), .B(n1189), .Z(n1194) );
  NANDN U1420 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U1421 ( .A(n1194), .B(n1193), .Z(n1289) );
  NAND U1422 ( .A(n1196), .B(n1195), .Z(n1200) );
  NANDN U1423 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U1424 ( .A(n1200), .B(n1199), .Z(n1288) );
  AND U1425 ( .A(y[10]), .B(x[16]), .Z(n2111) );
  NAND U1426 ( .A(n2111), .B(n1201), .Z(n1205) );
  NAND U1427 ( .A(n1203), .B(n1202), .Z(n1204) );
  NAND U1428 ( .A(n1205), .B(n1204), .Z(n1329) );
  AND U1429 ( .A(x[13]), .B(y[17]), .Z(n2578) );
  NAND U1430 ( .A(n2578), .B(n1206), .Z(n1210) );
  NANDN U1431 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1432 ( .A(n1210), .B(n1209), .Z(n1374) );
  AND U1433 ( .A(x[16]), .B(y[4]), .Z(n1212) );
  NAND U1434 ( .A(x[10]), .B(y[10]), .Z(n1211) );
  XNOR U1435 ( .A(n1212), .B(n1211), .Z(n1335) );
  AND U1436 ( .A(y[18]), .B(x[2]), .Z(n1336) );
  XOR U1437 ( .A(n1335), .B(n1336), .Z(n1372) );
  NAND U1438 ( .A(x[15]), .B(y[5]), .Z(n1213) );
  XNOR U1439 ( .A(n1214), .B(n1213), .Z(n1295) );
  AND U1440 ( .A(y[6]), .B(x[14]), .Z(n1296) );
  XOR U1441 ( .A(n1295), .B(n1296), .Z(n1371) );
  XOR U1442 ( .A(n1372), .B(n1371), .Z(n1373) );
  XOR U1443 ( .A(n1374), .B(n1373), .Z(n1328) );
  XOR U1444 ( .A(n1329), .B(n1328), .Z(n1331) );
  NAND U1445 ( .A(y[16]), .B(x[11]), .Z(n2327) );
  NANDN U1446 ( .A(n2327), .B(n1459), .Z(n1218) );
  NANDN U1447 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U1448 ( .A(n1218), .B(n1217), .Z(n1380) );
  AND U1449 ( .A(y[19]), .B(x[1]), .Z(n1220) );
  NAND U1450 ( .A(y[9]), .B(x[11]), .Z(n1219) );
  XNOR U1451 ( .A(n1220), .B(n1219), .Z(n1307) );
  AND U1452 ( .A(y[1]), .B(x[19]), .Z(n1299) );
  XOR U1453 ( .A(o[20]), .B(n1299), .Z(n1306) );
  XOR U1454 ( .A(n1307), .B(n1306), .Z(n1378) );
  AND U1455 ( .A(x[0]), .B(y[20]), .Z(n1359) );
  AND U1456 ( .A(y[0]), .B(x[20]), .Z(n1360) );
  XOR U1457 ( .A(n1359), .B(n1360), .Z(n1362) );
  AND U1458 ( .A(o[19]), .B(n1221), .Z(n1361) );
  XOR U1459 ( .A(n1362), .B(n1361), .Z(n1377) );
  XOR U1460 ( .A(n1378), .B(n1377), .Z(n1379) );
  XOR U1461 ( .A(n1380), .B(n1379), .Z(n1330) );
  XOR U1462 ( .A(n1331), .B(n1330), .Z(n1290) );
  XOR U1463 ( .A(n1291), .B(n1290), .Z(n1386) );
  NAND U1464 ( .A(x[6]), .B(y[14]), .Z(n1311) );
  NANDN U1465 ( .A(n1311), .B(n1222), .Z(n1225) );
  NAND U1466 ( .A(n1223), .B(n1354), .Z(n1224) );
  NAND U1467 ( .A(n1225), .B(n1224), .Z(n1319) );
  NAND U1468 ( .A(n1227), .B(n1226), .Z(n1231) );
  NAND U1469 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U1470 ( .A(n1231), .B(n1230), .Z(n1317) );
  AND U1471 ( .A(y[2]), .B(x[18]), .Z(n1233) );
  NAND U1472 ( .A(x[12]), .B(y[8]), .Z(n1232) );
  XNOR U1473 ( .A(n1233), .B(n1232), .Z(n1301) );
  AND U1474 ( .A(x[17]), .B(y[3]), .Z(n1302) );
  XOR U1475 ( .A(n1301), .B(n1302), .Z(n1316) );
  XOR U1476 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U1477 ( .A(n1319), .B(n1318), .Z(n1323) );
  AND U1478 ( .A(y[17]), .B(x[3]), .Z(n1235) );
  NAND U1479 ( .A(y[7]), .B(x[13]), .Z(n1234) );
  XNOR U1480 ( .A(n1235), .B(n1234), .Z(n1341) );
  XNOR U1481 ( .A(n1341), .B(n1340), .Z(n1313) );
  AND U1482 ( .A(y[15]), .B(x[5]), .Z(n1237) );
  NAND U1483 ( .A(x[4]), .B(y[16]), .Z(n1236) );
  XNOR U1484 ( .A(n1237), .B(n1236), .Z(n1356) );
  AND U1485 ( .A(x[7]), .B(y[13]), .Z(n1355) );
  XNOR U1486 ( .A(n1356), .B(n1355), .Z(n1310) );
  XOR U1487 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U1488 ( .A(n1313), .B(n1312), .Z(n1367) );
  AND U1489 ( .A(y[18]), .B(x[8]), .Z(n2423) );
  NAND U1490 ( .A(n2423), .B(n1238), .Z(n1242) );
  NANDN U1491 ( .A(n1240), .B(n1239), .Z(n1241) );
  NAND U1492 ( .A(n1242), .B(n1241), .Z(n1366) );
  AND U1493 ( .A(x[17]), .B(y[9]), .Z(n2114) );
  NAND U1494 ( .A(n2114), .B(n1243), .Z(n1247) );
  NAND U1495 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U1496 ( .A(n1247), .B(n1246), .Z(n1365) );
  XOR U1497 ( .A(n1366), .B(n1365), .Z(n1368) );
  XNOR U1498 ( .A(n1367), .B(n1368), .Z(n1322) );
  XOR U1499 ( .A(n1323), .B(n1322), .Z(n1324) );
  NANDN U1500 ( .A(n1249), .B(n1248), .Z(n1253) );
  NANDN U1501 ( .A(n1251), .B(n1250), .Z(n1252) );
  NAND U1502 ( .A(n1253), .B(n1252), .Z(n1325) );
  NAND U1503 ( .A(n1255), .B(n1254), .Z(n1259) );
  NANDN U1504 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U1505 ( .A(n1259), .B(n1258), .Z(n1384) );
  XOR U1506 ( .A(n1386), .B(n1385), .Z(n1389) );
  XOR U1507 ( .A(n1390), .B(n1389), .Z(n1392) );
  NAND U1508 ( .A(n1261), .B(n1260), .Z(n1265) );
  NAND U1509 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U1510 ( .A(n1265), .B(n1264), .Z(n1391) );
  XOR U1511 ( .A(n1392), .B(n1391), .Z(n1282) );
  NAND U1512 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U1513 ( .A(n1269), .B(n1268), .Z(n1270) );
  AND U1514 ( .A(n1271), .B(n1270), .Z(n1280) );
  NANDN U1515 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U1516 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U1517 ( .A(n1277), .B(n1276), .Z(n1279) );
  XOR U1518 ( .A(n1280), .B(n1279), .Z(n1281) );
  XNOR U1519 ( .A(n1286), .B(n1285), .Z(n1278) );
  XOR U1520 ( .A(n1287), .B(n1278), .Z(N53) );
  NAND U1521 ( .A(n1280), .B(n1279), .Z(n1284) );
  NANDN U1522 ( .A(n1282), .B(n1281), .Z(n1283) );
  NAND U1523 ( .A(n1284), .B(n1283), .Z(n1517) );
  NANDN U1524 ( .A(n1289), .B(n1288), .Z(n1293) );
  NAND U1525 ( .A(n1291), .B(n1290), .Z(n1292) );
  AND U1526 ( .A(n1293), .B(n1292), .Z(n1411) );
  AND U1527 ( .A(y[11]), .B(x[15]), .Z(n2105) );
  NAND U1528 ( .A(n2105), .B(n1294), .Z(n1298) );
  NAND U1529 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U1530 ( .A(n1298), .B(n1297), .Z(n1445) );
  AND U1531 ( .A(x[0]), .B(y[21]), .Z(n1466) );
  AND U1532 ( .A(y[0]), .B(x[21]), .Z(n1465) );
  XOR U1533 ( .A(n1466), .B(n1465), .Z(n1468) );
  AND U1534 ( .A(n1299), .B(o[20]), .Z(n1467) );
  XOR U1535 ( .A(n1468), .B(n1467), .Z(n1444) );
  AND U1536 ( .A(y[16]), .B(x[5]), .Z(n1450) );
  AND U1537 ( .A(y[5]), .B(x[16]), .Z(n1449) );
  XOR U1538 ( .A(n1450), .B(n1449), .Z(n1452) );
  AND U1539 ( .A(y[6]), .B(x[15]), .Z(n1451) );
  XOR U1540 ( .A(n1452), .B(n1451), .Z(n1443) );
  XOR U1541 ( .A(n1444), .B(n1443), .Z(n1446) );
  XOR U1542 ( .A(n1445), .B(n1446), .Z(n1490) );
  AND U1543 ( .A(y[8]), .B(x[18]), .Z(n2116) );
  NAND U1544 ( .A(n2116), .B(n1300), .Z(n1304) );
  NAND U1545 ( .A(n1302), .B(n1301), .Z(n1303) );
  AND U1546 ( .A(n1304), .B(n1303), .Z(n1488) );
  AND U1547 ( .A(x[11]), .B(y[19]), .Z(n2916) );
  NAND U1548 ( .A(n2916), .B(n1305), .Z(n1309) );
  NAND U1549 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U1550 ( .A(n1309), .B(n1308), .Z(n1487) );
  XNOR U1551 ( .A(n1490), .B(n1489), .Z(n1482) );
  NAND U1552 ( .A(n1311), .B(n1310), .Z(n1315) );
  NAND U1553 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1554 ( .A(n1315), .B(n1314), .Z(n1481) );
  XOR U1555 ( .A(n1482), .B(n1481), .Z(n1484) );
  NAND U1556 ( .A(n1317), .B(n1316), .Z(n1321) );
  NAND U1557 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U1558 ( .A(n1321), .B(n1320), .Z(n1483) );
  XOR U1559 ( .A(n1484), .B(n1483), .Z(n1409) );
  NAND U1560 ( .A(n1323), .B(n1322), .Z(n1327) );
  NANDN U1561 ( .A(n1325), .B(n1324), .Z(n1326) );
  AND U1562 ( .A(n1327), .B(n1326), .Z(n1408) );
  NAND U1563 ( .A(n1329), .B(n1328), .Z(n1333) );
  NAND U1564 ( .A(n1331), .B(n1330), .Z(n1332) );
  NAND U1565 ( .A(n1333), .B(n1332), .Z(n1508) );
  NAND U1566 ( .A(n2111), .B(n1334), .Z(n1338) );
  NAND U1567 ( .A(n1336), .B(n1335), .Z(n1337) );
  NAND U1568 ( .A(n1338), .B(n1337), .Z(n1415) );
  AND U1569 ( .A(x[3]), .B(y[7]), .Z(n1339) );
  NAND U1570 ( .A(n2578), .B(n1339), .Z(n1343) );
  NAND U1571 ( .A(n1341), .B(n1340), .Z(n1342) );
  NAND U1572 ( .A(n1343), .B(n1342), .Z(n1502) );
  AND U1573 ( .A(y[2]), .B(x[19]), .Z(n1345) );
  NAND U1574 ( .A(y[10]), .B(x[11]), .Z(n1344) );
  XNOR U1575 ( .A(n1345), .B(n1344), .Z(n1434) );
  AND U1576 ( .A(y[1]), .B(x[20]), .Z(n1464) );
  XOR U1577 ( .A(n1464), .B(o[21]), .Z(n1433) );
  XOR U1578 ( .A(n1434), .B(n1433), .Z(n1500) );
  NAND U1579 ( .A(y[3]), .B(x[18]), .Z(n1346) );
  XNOR U1580 ( .A(n1347), .B(n1346), .Z(n1473) );
  AND U1581 ( .A(x[1]), .B(y[20]), .Z(n1472) );
  XOR U1582 ( .A(n1473), .B(n1472), .Z(n1499) );
  XOR U1583 ( .A(n1500), .B(n1499), .Z(n1501) );
  XOR U1584 ( .A(n1502), .B(n1501), .Z(n1414) );
  XOR U1585 ( .A(n1415), .B(n1414), .Z(n1417) );
  AND U1586 ( .A(x[7]), .B(y[14]), .Z(n1684) );
  AND U1587 ( .A(y[15]), .B(x[6]), .Z(n1349) );
  AND U1588 ( .A(y[7]), .B(x[14]), .Z(n1348) );
  XOR U1589 ( .A(n1349), .B(n1348), .Z(n1476) );
  XOR U1590 ( .A(n1684), .B(n1476), .Z(n1423) );
  NAND U1591 ( .A(y[12]), .B(x[9]), .Z(n1421) );
  NAND U1592 ( .A(x[8]), .B(y[13]), .Z(n1420) );
  XOR U1593 ( .A(n1421), .B(n1420), .Z(n1422) );
  AND U1594 ( .A(x[12]), .B(y[9]), .Z(n1351) );
  NAND U1595 ( .A(y[4]), .B(x[17]), .Z(n1350) );
  XNOR U1596 ( .A(n1351), .B(n1350), .Z(n1427) );
  AND U1597 ( .A(x[2]), .B(y[19]), .Z(n1426) );
  XOR U1598 ( .A(n1427), .B(n1426), .Z(n1438) );
  AND U1599 ( .A(y[18]), .B(x[3]), .Z(n1353) );
  NAND U1600 ( .A(y[8]), .B(x[13]), .Z(n1352) );
  XNOR U1601 ( .A(n1353), .B(n1352), .Z(n1461) );
  AND U1602 ( .A(y[17]), .B(x[4]), .Z(n1460) );
  XOR U1603 ( .A(n1461), .B(n1460), .Z(n1437) );
  XOR U1604 ( .A(n1438), .B(n1437), .Z(n1439) );
  NAND U1605 ( .A(n1450), .B(n1354), .Z(n1358) );
  NAND U1606 ( .A(n1356), .B(n1355), .Z(n1357) );
  NAND U1607 ( .A(n1358), .B(n1357), .Z(n1494) );
  NAND U1608 ( .A(n1360), .B(n1359), .Z(n1364) );
  NAND U1609 ( .A(n1362), .B(n1361), .Z(n1363) );
  NAND U1610 ( .A(n1364), .B(n1363), .Z(n1493) );
  XOR U1611 ( .A(n1494), .B(n1493), .Z(n1495) );
  XOR U1612 ( .A(n1496), .B(n1495), .Z(n1416) );
  XOR U1613 ( .A(n1417), .B(n1416), .Z(n1506) );
  NAND U1614 ( .A(n1366), .B(n1365), .Z(n1370) );
  NAND U1615 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U1616 ( .A(n1370), .B(n1369), .Z(n1513) );
  NAND U1617 ( .A(n1372), .B(n1371), .Z(n1376) );
  NAND U1618 ( .A(n1374), .B(n1373), .Z(n1375) );
  NAND U1619 ( .A(n1376), .B(n1375), .Z(n1512) );
  NAND U1620 ( .A(n1378), .B(n1377), .Z(n1382) );
  NAND U1621 ( .A(n1380), .B(n1379), .Z(n1381) );
  NAND U1622 ( .A(n1382), .B(n1381), .Z(n1511) );
  XOR U1623 ( .A(n1512), .B(n1511), .Z(n1514) );
  XOR U1624 ( .A(n1513), .B(n1514), .Z(n1505) );
  XOR U1625 ( .A(n1506), .B(n1505), .Z(n1507) );
  XNOR U1626 ( .A(n1508), .B(n1507), .Z(n1403) );
  NANDN U1627 ( .A(n1384), .B(n1383), .Z(n1388) );
  NANDN U1628 ( .A(n1386), .B(n1385), .Z(n1387) );
  NAND U1629 ( .A(n1388), .B(n1387), .Z(n1402) );
  XOR U1630 ( .A(n1403), .B(n1402), .Z(n1405) );
  XNOR U1631 ( .A(n1404), .B(n1405), .Z(n1523) );
  NAND U1632 ( .A(n1390), .B(n1389), .Z(n1394) );
  NAND U1633 ( .A(n1392), .B(n1391), .Z(n1393) );
  NAND U1634 ( .A(n1394), .B(n1393), .Z(n1520) );
  NAND U1635 ( .A(n1396), .B(n1395), .Z(n1400) );
  NAND U1636 ( .A(n1398), .B(n1397), .Z(n1399) );
  AND U1637 ( .A(n1400), .B(n1399), .Z(n1521) );
  XOR U1638 ( .A(n1520), .B(n1521), .Z(n1522) );
  XOR U1639 ( .A(n1523), .B(n1522), .Z(n1519) );
  XNOR U1640 ( .A(n1518), .B(n1519), .Z(n1401) );
  XNOR U1641 ( .A(n1517), .B(n1401), .Z(N54) );
  NAND U1642 ( .A(n1403), .B(n1402), .Z(n1407) );
  NAND U1643 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U1644 ( .A(n1407), .B(n1406), .Z(n1649) );
  NANDN U1645 ( .A(n1409), .B(n1408), .Z(n1413) );
  NANDN U1646 ( .A(n1411), .B(n1410), .Z(n1412) );
  AND U1647 ( .A(n1413), .B(n1412), .Z(n1647) );
  NAND U1648 ( .A(n1415), .B(n1414), .Z(n1419) );
  NAND U1649 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U1650 ( .A(n1419), .B(n1418), .Z(n1637) );
  NAND U1651 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U1652 ( .A(n1423), .B(n1422), .Z(n1424) );
  AND U1653 ( .A(n1425), .B(n1424), .Z(n1631) );
  NAND U1654 ( .A(n2114), .B(n1588), .Z(n1429) );
  NAND U1655 ( .A(n1427), .B(n1426), .Z(n1428) );
  AND U1656 ( .A(n1429), .B(n1428), .Z(n1560) );
  AND U1657 ( .A(x[5]), .B(y[17]), .Z(n1604) );
  NAND U1658 ( .A(y[5]), .B(x[17]), .Z(n1605) );
  NAND U1659 ( .A(y[6]), .B(x[16]), .Z(n1607) );
  AND U1660 ( .A(x[18]), .B(y[4]), .Z(n1431) );
  NAND U1661 ( .A(x[12]), .B(y[10]), .Z(n1430) );
  XNOR U1662 ( .A(n1431), .B(n1430), .Z(n1589) );
  NAND U1663 ( .A(y[18]), .B(x[4]), .Z(n1590) );
  XOR U1664 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1665 ( .A(y[10]), .B(x[19]), .Z(n2642) );
  NAND U1666 ( .A(n2642), .B(n1432), .Z(n1436) );
  NAND U1667 ( .A(n1434), .B(n1433), .Z(n1435) );
  AND U1668 ( .A(n1436), .B(n1435), .Z(n1629) );
  XOR U1669 ( .A(n1628), .B(n1629), .Z(n1630) );
  NAND U1670 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1671 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1672 ( .A(n1442), .B(n1441), .Z(n1617) );
  NAND U1673 ( .A(n1444), .B(n1443), .Z(n1448) );
  NAND U1674 ( .A(n1446), .B(n1445), .Z(n1447) );
  NAND U1675 ( .A(n1448), .B(n1447), .Z(n1616) );
  NAND U1676 ( .A(n1450), .B(n1449), .Z(n1454) );
  AND U1677 ( .A(n1452), .B(n1451), .Z(n1453) );
  ANDN U1678 ( .B(n1454), .A(n1453), .Z(n1579) );
  AND U1679 ( .A(y[2]), .B(x[20]), .Z(n1456) );
  NAND U1680 ( .A(y[9]), .B(x[13]), .Z(n1455) );
  XNOR U1681 ( .A(n1456), .B(n1455), .Z(n1600) );
  NAND U1682 ( .A(x[2]), .B(y[20]), .Z(n1601) );
  AND U1683 ( .A(x[15]), .B(y[7]), .Z(n1458) );
  NAND U1684 ( .A(x[6]), .B(y[16]), .Z(n1457) );
  XNOR U1685 ( .A(n1458), .B(n1457), .Z(n1612) );
  XOR U1686 ( .A(n1577), .B(n1576), .Z(n1578) );
  AND U1687 ( .A(x[13]), .B(y[18]), .Z(n2917) );
  NAND U1688 ( .A(n1459), .B(n2917), .Z(n1463) );
  NAND U1689 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1690 ( .A(n1463), .B(n1462), .Z(n1548) );
  AND U1691 ( .A(y[21]), .B(x[1]), .Z(n1571) );
  XOR U1692 ( .A(n1572), .B(n1571), .Z(n1570) );
  AND U1693 ( .A(n1464), .B(o[21]), .Z(n1569) );
  XOR U1694 ( .A(n1570), .B(n1569), .Z(n1546) );
  AND U1695 ( .A(x[14]), .B(y[8]), .Z(n1563) );
  AND U1696 ( .A(x[3]), .B(y[19]), .Z(n1564) );
  XOR U1697 ( .A(n1563), .B(n1564), .Z(n1565) );
  AND U1698 ( .A(x[19]), .B(y[3]), .Z(n1566) );
  XOR U1699 ( .A(n1565), .B(n1566), .Z(n1545) );
  XOR U1700 ( .A(n1546), .B(n1545), .Z(n1547) );
  XNOR U1701 ( .A(n1622), .B(n1623), .Z(n1625) );
  NAND U1702 ( .A(n1466), .B(n1465), .Z(n1470) );
  NAND U1703 ( .A(n1468), .B(n1467), .Z(n1469) );
  AND U1704 ( .A(n1470), .B(n1469), .Z(n1540) );
  AND U1705 ( .A(x[18]), .B(y[11]), .Z(n2645) );
  NAND U1706 ( .A(n2645), .B(n1471), .Z(n1475) );
  NAND U1707 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U1708 ( .A(n1475), .B(n1474), .Z(n1539) );
  AND U1709 ( .A(x[14]), .B(y[15]), .Z(n2612) );
  NAND U1710 ( .A(n2612), .B(n1611), .Z(n1478) );
  NAND U1711 ( .A(n1684), .B(n1476), .Z(n1477) );
  NAND U1712 ( .A(n1478), .B(n1477), .Z(n1553) );
  AND U1713 ( .A(x[0]), .B(y[22]), .Z(n1593) );
  NAND U1714 ( .A(y[0]), .B(x[22]), .Z(n1594) );
  AND U1715 ( .A(y[1]), .B(x[21]), .Z(n1610) );
  XOR U1716 ( .A(o[22]), .B(n1610), .Z(n1595) );
  XOR U1717 ( .A(n1596), .B(n1595), .Z(n1552) );
  AND U1718 ( .A(y[15]), .B(x[7]), .Z(n1480) );
  NAND U1719 ( .A(y[14]), .B(x[8]), .Z(n1479) );
  XNOR U1720 ( .A(n1480), .B(n1479), .Z(n1583) );
  XOR U1721 ( .A(n1583), .B(n1582), .Z(n1551) );
  XOR U1722 ( .A(n1552), .B(n1551), .Z(n1554) );
  XOR U1723 ( .A(n1553), .B(n1554), .Z(n1541) );
  XOR U1724 ( .A(n1542), .B(n1541), .Z(n1624) );
  XOR U1725 ( .A(n1625), .B(n1624), .Z(n1618) );
  XOR U1726 ( .A(n1619), .B(n1618), .Z(n1635) );
  XOR U1727 ( .A(n1634), .B(n1635), .Z(n1636) );
  NAND U1728 ( .A(n1482), .B(n1481), .Z(n1486) );
  NAND U1729 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1730 ( .A(n1486), .B(n1485), .Z(n1641) );
  NANDN U1731 ( .A(n1488), .B(n1487), .Z(n1492) );
  NAND U1732 ( .A(n1490), .B(n1489), .Z(n1491) );
  AND U1733 ( .A(n1492), .B(n1491), .Z(n1536) );
  NAND U1734 ( .A(n1494), .B(n1493), .Z(n1498) );
  NAND U1735 ( .A(n1496), .B(n1495), .Z(n1497) );
  AND U1736 ( .A(n1498), .B(n1497), .Z(n1534) );
  NAND U1737 ( .A(n1500), .B(n1499), .Z(n1504) );
  NAND U1738 ( .A(n1502), .B(n1501), .Z(n1503) );
  NAND U1739 ( .A(n1504), .B(n1503), .Z(n1533) );
  XOR U1740 ( .A(n1641), .B(n1640), .Z(n1642) );
  XOR U1741 ( .A(n1643), .B(n1642), .Z(n1530) );
  NAND U1742 ( .A(n1506), .B(n1505), .Z(n1510) );
  NAND U1743 ( .A(n1508), .B(n1507), .Z(n1509) );
  NAND U1744 ( .A(n1510), .B(n1509), .Z(n1528) );
  NAND U1745 ( .A(n1512), .B(n1511), .Z(n1516) );
  NAND U1746 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U1747 ( .A(n1516), .B(n1515), .Z(n1527) );
  XOR U1748 ( .A(n1528), .B(n1527), .Z(n1529) );
  XOR U1749 ( .A(n1530), .B(n1529), .Z(n1646) );
  XNOR U1750 ( .A(n1649), .B(n1648), .Z(n1654) );
  NAND U1751 ( .A(n1521), .B(n1520), .Z(n1525) );
  NAND U1752 ( .A(n1523), .B(n1522), .Z(n1524) );
  NAND U1753 ( .A(n1525), .B(n1524), .Z(n1653) );
  XOR U1754 ( .A(n1652), .B(n1653), .Z(n1526) );
  XNOR U1755 ( .A(n1654), .B(n1526), .Z(N55) );
  NAND U1756 ( .A(n1528), .B(n1527), .Z(n1532) );
  NAND U1757 ( .A(n1530), .B(n1529), .Z(n1531) );
  AND U1758 ( .A(n1532), .B(n1531), .Z(n1659) );
  NANDN U1759 ( .A(n1534), .B(n1533), .Z(n1538) );
  NANDN U1760 ( .A(n1536), .B(n1535), .Z(n1537) );
  NAND U1761 ( .A(n1538), .B(n1537), .Z(n1779) );
  NANDN U1762 ( .A(n1540), .B(n1539), .Z(n1544) );
  NAND U1763 ( .A(n1542), .B(n1541), .Z(n1543) );
  NAND U1764 ( .A(n1544), .B(n1543), .Z(n1773) );
  NAND U1765 ( .A(n1546), .B(n1545), .Z(n1550) );
  NANDN U1766 ( .A(n1548), .B(n1547), .Z(n1549) );
  NAND U1767 ( .A(n1550), .B(n1549), .Z(n1772) );
  NAND U1768 ( .A(n1552), .B(n1551), .Z(n1556) );
  NAND U1769 ( .A(n1554), .B(n1553), .Z(n1555) );
  NAND U1770 ( .A(n1556), .B(n1555), .Z(n1771) );
  XOR U1771 ( .A(n1772), .B(n1771), .Z(n1774) );
  XOR U1772 ( .A(n1773), .B(n1774), .Z(n1791) );
  NAND U1773 ( .A(n1558), .B(n1557), .Z(n1562) );
  NANDN U1774 ( .A(n1560), .B(n1559), .Z(n1561) );
  NAND U1775 ( .A(n1562), .B(n1561), .Z(n1789) );
  NAND U1776 ( .A(n1564), .B(n1563), .Z(n1568) );
  NAND U1777 ( .A(n1566), .B(n1565), .Z(n1567) );
  NAND U1778 ( .A(n1568), .B(n1567), .Z(n1718) );
  AND U1779 ( .A(n1570), .B(n1569), .Z(n1574) );
  NAND U1780 ( .A(n1572), .B(n1571), .Z(n1573) );
  NANDN U1781 ( .A(n1574), .B(n1573), .Z(n1717) );
  XOR U1782 ( .A(n1718), .B(n1717), .Z(n1720) );
  NAND U1783 ( .A(x[7]), .B(y[16]), .Z(n1575) );
  XNOR U1784 ( .A(n1855), .B(n1575), .Z(n1685) );
  AND U1785 ( .A(y[13]), .B(x[10]), .Z(n1724) );
  XOR U1786 ( .A(n1723), .B(n1724), .Z(n1726) );
  AND U1787 ( .A(x[6]), .B(y[17]), .Z(n1676) );
  AND U1788 ( .A(y[8]), .B(x[15]), .Z(n1677) );
  XOR U1789 ( .A(n1676), .B(n1677), .Z(n1678) );
  AND U1790 ( .A(y[12]), .B(x[11]), .Z(n1679) );
  XOR U1791 ( .A(n1678), .B(n1679), .Z(n1725) );
  XOR U1792 ( .A(n1726), .B(n1725), .Z(n1719) );
  XOR U1793 ( .A(n1720), .B(n1719), .Z(n1790) );
  XNOR U1794 ( .A(n1789), .B(n1790), .Z(n1792) );
  NAND U1795 ( .A(n1577), .B(n1576), .Z(n1581) );
  NANDN U1796 ( .A(n1579), .B(n1578), .Z(n1580) );
  AND U1797 ( .A(n1581), .B(n1580), .Z(n1712) );
  NANDN U1798 ( .A(n1686), .B(n1684), .Z(n1585) );
  NAND U1799 ( .A(n1583), .B(n1582), .Z(n1584) );
  AND U1800 ( .A(n1585), .B(n1584), .Z(n1762) );
  AND U1801 ( .A(x[0]), .B(y[23]), .Z(n1695) );
  AND U1802 ( .A(x[23]), .B(y[0]), .Z(n1696) );
  XOR U1803 ( .A(n1695), .B(n1696), .Z(n1698) );
  AND U1804 ( .A(y[1]), .B(x[22]), .Z(n1675) );
  XOR U1805 ( .A(o[23]), .B(n1675), .Z(n1697) );
  XOR U1806 ( .A(n1698), .B(n1697), .Z(n1760) );
  NAND U1807 ( .A(y[3]), .B(x[20]), .Z(n1586) );
  XNOR U1808 ( .A(n1587), .B(n1586), .Z(n1671) );
  AND U1809 ( .A(y[4]), .B(x[19]), .Z(n1672) );
  XOR U1810 ( .A(n1671), .B(n1672), .Z(n1759) );
  XOR U1811 ( .A(n1760), .B(n1759), .Z(n1761) );
  AND U1812 ( .A(y[10]), .B(x[18]), .Z(n2447) );
  NAND U1813 ( .A(n2447), .B(n1588), .Z(n1592) );
  NANDN U1814 ( .A(n1590), .B(n1589), .Z(n1591) );
  AND U1815 ( .A(n1592), .B(n1591), .Z(n1748) );
  NANDN U1816 ( .A(n1594), .B(n1593), .Z(n1598) );
  NAND U1817 ( .A(n1596), .B(n1595), .Z(n1597) );
  NAND U1818 ( .A(n1598), .B(n1597), .Z(n1747) );
  XOR U1819 ( .A(n1750), .B(n1749), .Z(n1711) );
  AND U1820 ( .A(x[20]), .B(y[9]), .Z(n2623) );
  AND U1821 ( .A(x[13]), .B(y[2]), .Z(n1599) );
  NAND U1822 ( .A(n2623), .B(n1599), .Z(n1603) );
  NANDN U1823 ( .A(n1601), .B(n1600), .Z(n1602) );
  AND U1824 ( .A(n1603), .B(n1602), .Z(n1706) );
  NANDN U1825 ( .A(n1605), .B(n1604), .Z(n1609) );
  NANDN U1826 ( .A(n1607), .B(n1606), .Z(n1608) );
  AND U1827 ( .A(n1609), .B(n1608), .Z(n1768) );
  AND U1828 ( .A(x[13]), .B(y[10]), .Z(n1741) );
  AND U1829 ( .A(y[21]), .B(x[2]), .Z(n1742) );
  XOR U1830 ( .A(n1741), .B(n1742), .Z(n1743) );
  AND U1831 ( .A(x[21]), .B(y[2]), .Z(n1744) );
  XOR U1832 ( .A(n1743), .B(n1744), .Z(n1766) );
  AND U1833 ( .A(y[11]), .B(x[12]), .Z(n1689) );
  AND U1834 ( .A(y[22]), .B(x[1]), .Z(n1690) );
  XOR U1835 ( .A(n1689), .B(n1690), .Z(n1692) );
  AND U1836 ( .A(o[22]), .B(n1610), .Z(n1691) );
  XOR U1837 ( .A(n1692), .B(n1691), .Z(n1765) );
  XOR U1838 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U1839 ( .A(y[16]), .B(x[15]), .Z(n2865) );
  NAND U1840 ( .A(n2865), .B(n1611), .Z(n1615) );
  NANDN U1841 ( .A(n1613), .B(n1612), .Z(n1614) );
  AND U1842 ( .A(n1615), .B(n1614), .Z(n1756) );
  AND U1843 ( .A(x[14]), .B(y[9]), .Z(n1735) );
  AND U1844 ( .A(x[3]), .B(y[20]), .Z(n1736) );
  XOR U1845 ( .A(n1735), .B(n1736), .Z(n1737) );
  AND U1846 ( .A(x[4]), .B(y[19]), .Z(n1738) );
  XOR U1847 ( .A(n1737), .B(n1738), .Z(n1754) );
  AND U1848 ( .A(y[18]), .B(x[5]), .Z(n1729) );
  AND U1849 ( .A(y[5]), .B(x[18]), .Z(n1730) );
  XOR U1850 ( .A(n1729), .B(n1730), .Z(n1731) );
  AND U1851 ( .A(y[6]), .B(x[17]), .Z(n1732) );
  XOR U1852 ( .A(n1731), .B(n1732), .Z(n1753) );
  XOR U1853 ( .A(n1754), .B(n1753), .Z(n1755) );
  XOR U1854 ( .A(n1708), .B(n1707), .Z(n1713) );
  XOR U1855 ( .A(n1714), .B(n1713), .Z(n1777) );
  XOR U1856 ( .A(n1778), .B(n1777), .Z(n1780) );
  XOR U1857 ( .A(n1779), .B(n1780), .Z(n1668) );
  NANDN U1858 ( .A(n1617), .B(n1616), .Z(n1621) );
  NAND U1859 ( .A(n1619), .B(n1618), .Z(n1620) );
  NAND U1860 ( .A(n1621), .B(n1620), .Z(n1785) );
  NANDN U1861 ( .A(n1623), .B(n1622), .Z(n1627) );
  NAND U1862 ( .A(n1625), .B(n1624), .Z(n1626) );
  NAND U1863 ( .A(n1627), .B(n1626), .Z(n1783) );
  NAND U1864 ( .A(n1629), .B(n1628), .Z(n1633) );
  NANDN U1865 ( .A(n1631), .B(n1630), .Z(n1632) );
  AND U1866 ( .A(n1633), .B(n1632), .Z(n1784) );
  XOR U1867 ( .A(n1783), .B(n1784), .Z(n1786) );
  XOR U1868 ( .A(n1785), .B(n1786), .Z(n1666) );
  NAND U1869 ( .A(n1635), .B(n1634), .Z(n1639) );
  NANDN U1870 ( .A(n1637), .B(n1636), .Z(n1638) );
  AND U1871 ( .A(n1639), .B(n1638), .Z(n1665) );
  NAND U1872 ( .A(n1641), .B(n1640), .Z(n1645) );
  NAND U1873 ( .A(n1643), .B(n1642), .Z(n1644) );
  AND U1874 ( .A(n1645), .B(n1644), .Z(n1657) );
  XOR U1875 ( .A(n1656), .B(n1657), .Z(n1658) );
  XOR U1876 ( .A(n1659), .B(n1658), .Z(n1664) );
  NANDN U1877 ( .A(n1647), .B(n1646), .Z(n1651) );
  NAND U1878 ( .A(n1649), .B(n1648), .Z(n1650) );
  NAND U1879 ( .A(n1651), .B(n1650), .Z(n1662) );
  XOR U1880 ( .A(n1662), .B(n1663), .Z(n1655) );
  XNOR U1881 ( .A(n1664), .B(n1655), .Z(N56) );
  NAND U1882 ( .A(n1657), .B(n1656), .Z(n1661) );
  NAND U1883 ( .A(n1659), .B(n1658), .Z(n1660) );
  NAND U1884 ( .A(n1661), .B(n1660), .Z(n1928) );
  IV U1885 ( .A(n1928), .Z(n1926) );
  NANDN U1886 ( .A(n1666), .B(n1665), .Z(n1670) );
  NANDN U1887 ( .A(n1668), .B(n1667), .Z(n1669) );
  AND U1888 ( .A(n1670), .B(n1669), .Z(n1935) );
  AND U1889 ( .A(x[20]), .B(y[7]), .Z(n2197) );
  NAND U1890 ( .A(n2197), .B(n1826), .Z(n1674) );
  NAND U1891 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U1892 ( .A(n1674), .B(n1673), .Z(n1846) );
  AND U1893 ( .A(x[22]), .B(y[2]), .Z(n1865) );
  XOR U1894 ( .A(n1866), .B(n1865), .Z(n1868) );
  NAND U1895 ( .A(y[22]), .B(x[2]), .Z(n1867) );
  AND U1896 ( .A(y[23]), .B(x[1]), .Z(n1873) );
  XOR U1897 ( .A(n1874), .B(n1873), .Z(n1872) );
  AND U1898 ( .A(o[23]), .B(n1675), .Z(n1871) );
  XOR U1899 ( .A(n1872), .B(n1871), .Z(n1843) );
  XOR U1900 ( .A(n1844), .B(n1843), .Z(n1845) );
  XOR U1901 ( .A(n1846), .B(n1845), .Z(n1903) );
  NAND U1902 ( .A(n1677), .B(n1676), .Z(n1681) );
  NAND U1903 ( .A(n1679), .B(n1678), .Z(n1680) );
  NAND U1904 ( .A(n1681), .B(n1680), .Z(n1840) );
  AND U1905 ( .A(y[3]), .B(x[21]), .Z(n1683) );
  NAND U1906 ( .A(x[16]), .B(y[8]), .Z(n1682) );
  XNOR U1907 ( .A(n1683), .B(n1682), .Z(n1827) );
  AND U1908 ( .A(x[5]), .B(y[19]), .Z(n1828) );
  XOR U1909 ( .A(n1827), .B(n1828), .Z(n1838) );
  AND U1910 ( .A(y[18]), .B(x[6]), .Z(n2186) );
  AND U1911 ( .A(x[20]), .B(y[4]), .Z(n2029) );
  XOR U1912 ( .A(n2186), .B(n2029), .Z(n1833) );
  AND U1913 ( .A(y[5]), .B(x[19]), .Z(n1834) );
  XOR U1914 ( .A(n1833), .B(n1834), .Z(n1837) );
  XOR U1915 ( .A(n1838), .B(n1837), .Z(n1839) );
  XOR U1916 ( .A(n1840), .B(n1839), .Z(n1817) );
  NANDN U1917 ( .A(n1962), .B(n1684), .Z(n1688) );
  NANDN U1918 ( .A(n1686), .B(n1685), .Z(n1687) );
  NAND U1919 ( .A(n1688), .B(n1687), .Z(n1815) );
  NAND U1920 ( .A(n1690), .B(n1689), .Z(n1694) );
  NAND U1921 ( .A(n1692), .B(n1691), .Z(n1693) );
  NAND U1922 ( .A(n1694), .B(n1693), .Z(n1814) );
  XOR U1923 ( .A(n1815), .B(n1814), .Z(n1816) );
  XOR U1924 ( .A(n1817), .B(n1816), .Z(n1902) );
  XOR U1925 ( .A(n1903), .B(n1902), .Z(n1905) );
  NAND U1926 ( .A(n1696), .B(n1695), .Z(n1700) );
  NAND U1927 ( .A(n1698), .B(n1697), .Z(n1699) );
  NAND U1928 ( .A(n1700), .B(n1699), .Z(n1897) );
  AND U1929 ( .A(x[3]), .B(y[21]), .Z(n1886) );
  XOR U1930 ( .A(n1887), .B(n1886), .Z(n1885) );
  AND U1931 ( .A(x[4]), .B(y[20]), .Z(n1884) );
  XOR U1932 ( .A(n1885), .B(n1884), .Z(n1896) );
  XOR U1933 ( .A(n1897), .B(n1896), .Z(n1899) );
  AND U1934 ( .A(x[10]), .B(y[14]), .Z(n1702) );
  NAND U1935 ( .A(x[9]), .B(y[15]), .Z(n1701) );
  XNOR U1936 ( .A(n1702), .B(n1701), .Z(n1857) );
  AND U1937 ( .A(y[10]), .B(x[14]), .Z(n1704) );
  NAND U1938 ( .A(x[8]), .B(y[16]), .Z(n1703) );
  XNOR U1939 ( .A(n1704), .B(n1703), .Z(n1861) );
  AND U1940 ( .A(x[11]), .B(y[13]), .Z(n1862) );
  XOR U1941 ( .A(n1861), .B(n1862), .Z(n1856) );
  XOR U1942 ( .A(n1857), .B(n1856), .Z(n1898) );
  XOR U1943 ( .A(n1899), .B(n1898), .Z(n1904) );
  XOR U1944 ( .A(n1905), .B(n1904), .Z(n1915) );
  NANDN U1945 ( .A(n1706), .B(n1705), .Z(n1710) );
  NAND U1946 ( .A(n1708), .B(n1707), .Z(n1709) );
  AND U1947 ( .A(n1710), .B(n1709), .Z(n1914) );
  NANDN U1948 ( .A(n1712), .B(n1711), .Z(n1716) );
  NAND U1949 ( .A(n1714), .B(n1713), .Z(n1715) );
  NAND U1950 ( .A(n1716), .B(n1715), .Z(n1917) );
  NAND U1951 ( .A(n1718), .B(n1717), .Z(n1722) );
  NAND U1952 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U1953 ( .A(n1722), .B(n1721), .Z(n1911) );
  NAND U1954 ( .A(n1724), .B(n1723), .Z(n1728) );
  NAND U1955 ( .A(n1726), .B(n1725), .Z(n1727) );
  NAND U1956 ( .A(n1728), .B(n1727), .Z(n1909) );
  NAND U1957 ( .A(n1730), .B(n1729), .Z(n1734) );
  NAND U1958 ( .A(n1732), .B(n1731), .Z(n1733) );
  NAND U1959 ( .A(n1734), .B(n1733), .Z(n1823) );
  AND U1960 ( .A(x[0]), .B(y[24]), .Z(n1890) );
  AND U1961 ( .A(x[24]), .B(y[0]), .Z(n1891) );
  XOR U1962 ( .A(n1890), .B(n1891), .Z(n1892) );
  NAND U1963 ( .A(x[23]), .B(y[1]), .Z(n1883) );
  XNOR U1964 ( .A(o[24]), .B(n1883), .Z(n1893) );
  XOR U1965 ( .A(n1892), .B(n1893), .Z(n1821) );
  AND U1966 ( .A(x[7]), .B(y[17]), .Z(n1877) );
  NAND U1967 ( .A(y[6]), .B(x[18]), .Z(n1878) );
  NAND U1968 ( .A(x[17]), .B(y[7]), .Z(n1880) );
  XOR U1969 ( .A(n1821), .B(n1820), .Z(n1822) );
  XOR U1970 ( .A(n1823), .B(n1822), .Z(n1811) );
  NAND U1971 ( .A(n1736), .B(n1735), .Z(n1740) );
  NAND U1972 ( .A(n1738), .B(n1737), .Z(n1739) );
  NAND U1973 ( .A(n1740), .B(n1739), .Z(n1809) );
  NAND U1974 ( .A(n1742), .B(n1741), .Z(n1746) );
  NAND U1975 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U1976 ( .A(n1746), .B(n1745), .Z(n1808) );
  XOR U1977 ( .A(n1809), .B(n1808), .Z(n1810) );
  XOR U1978 ( .A(n1811), .B(n1810), .Z(n1908) );
  XOR U1979 ( .A(n1909), .B(n1908), .Z(n1910) );
  XNOR U1980 ( .A(n1911), .B(n1910), .Z(n1851) );
  NANDN U1981 ( .A(n1748), .B(n1747), .Z(n1752) );
  NAND U1982 ( .A(n1750), .B(n1749), .Z(n1751) );
  AND U1983 ( .A(n1752), .B(n1751), .Z(n1805) );
  NAND U1984 ( .A(n1754), .B(n1753), .Z(n1758) );
  NANDN U1985 ( .A(n1756), .B(n1755), .Z(n1757) );
  AND U1986 ( .A(n1758), .B(n1757), .Z(n1802) );
  NAND U1987 ( .A(n1760), .B(n1759), .Z(n1764) );
  NANDN U1988 ( .A(n1762), .B(n1761), .Z(n1763) );
  NAND U1989 ( .A(n1764), .B(n1763), .Z(n1803) );
  XOR U1990 ( .A(n1805), .B(n1804), .Z(n1849) );
  NAND U1991 ( .A(n1766), .B(n1765), .Z(n1770) );
  NANDN U1992 ( .A(n1768), .B(n1767), .Z(n1769) );
  NAND U1993 ( .A(n1770), .B(n1769), .Z(n1850) );
  XOR U1994 ( .A(n1851), .B(n1852), .Z(n1921) );
  NAND U1995 ( .A(n1772), .B(n1771), .Z(n1776) );
  NAND U1996 ( .A(n1774), .B(n1773), .Z(n1775) );
  AND U1997 ( .A(n1776), .B(n1775), .Z(n1920) );
  XOR U1998 ( .A(n1921), .B(n1920), .Z(n1922) );
  XNOR U1999 ( .A(n1923), .B(n1922), .Z(n1933) );
  NAND U2000 ( .A(n1778), .B(n1777), .Z(n1782) );
  NAND U2001 ( .A(n1780), .B(n1779), .Z(n1781) );
  NAND U2002 ( .A(n1782), .B(n1781), .Z(n1798) );
  NAND U2003 ( .A(n1784), .B(n1783), .Z(n1788) );
  NAND U2004 ( .A(n1786), .B(n1785), .Z(n1787) );
  NAND U2005 ( .A(n1788), .B(n1787), .Z(n1797) );
  NAND U2006 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U2007 ( .A(n1792), .B(n1791), .Z(n1793) );
  NAND U2008 ( .A(n1794), .B(n1793), .Z(n1796) );
  XNOR U2009 ( .A(n1797), .B(n1796), .Z(n1799) );
  XOR U2010 ( .A(n1933), .B(n1934), .Z(n1936) );
  XNOR U2011 ( .A(n1935), .B(n1936), .Z(n1929) );
  XNOR U2012 ( .A(n1927), .B(n1929), .Z(n1795) );
  XOR U2013 ( .A(n1926), .B(n1795), .Z(N57) );
  NAND U2014 ( .A(n1797), .B(n1796), .Z(n1801) );
  NANDN U2015 ( .A(n1799), .B(n1798), .Z(n1800) );
  AND U2016 ( .A(n1801), .B(n1800), .Z(n2074) );
  NANDN U2017 ( .A(n1803), .B(n1802), .Z(n1807) );
  NAND U2018 ( .A(n1805), .B(n1804), .Z(n1806) );
  AND U2019 ( .A(n1807), .B(n1806), .Z(n1947) );
  NAND U2020 ( .A(n1809), .B(n1808), .Z(n1813) );
  NAND U2021 ( .A(n1811), .B(n1810), .Z(n1812) );
  NAND U2022 ( .A(n1813), .B(n1812), .Z(n1953) );
  NAND U2023 ( .A(n1815), .B(n1814), .Z(n1819) );
  NAND U2024 ( .A(n1817), .B(n1816), .Z(n1818) );
  NAND U2025 ( .A(n1819), .B(n1818), .Z(n1952) );
  XOR U2026 ( .A(n1953), .B(n1952), .Z(n1955) );
  NAND U2027 ( .A(n1821), .B(n1820), .Z(n1825) );
  NAND U2028 ( .A(n1823), .B(n1822), .Z(n1824) );
  AND U2029 ( .A(n1825), .B(n1824), .Z(n1981) );
  AND U2030 ( .A(y[8]), .B(x[21]), .Z(n2923) );
  NAND U2031 ( .A(n2923), .B(n1826), .Z(n1830) );
  NAND U2032 ( .A(n1828), .B(n1827), .Z(n1829) );
  NAND U2033 ( .A(n1830), .B(n1829), .Z(n2047) );
  NAND U2034 ( .A(x[22]), .B(y[3]), .Z(n2022) );
  NAND U2035 ( .A(x[5]), .B(y[20]), .Z(n2020) );
  NAND U2036 ( .A(x[17]), .B(y[8]), .Z(n2021) );
  XNOR U2037 ( .A(n2020), .B(n2021), .Z(n2023) );
  XOR U2038 ( .A(n2022), .B(n2023), .Z(n2044) );
  AND U2039 ( .A(y[4]), .B(x[21]), .Z(n1832) );
  NAND U2040 ( .A(x[20]), .B(y[5]), .Z(n1831) );
  XNOR U2041 ( .A(n1832), .B(n1831), .Z(n2031) );
  AND U2042 ( .A(y[6]), .B(x[19]), .Z(n2030) );
  XOR U2043 ( .A(n2031), .B(n2030), .Z(n2045) );
  XOR U2044 ( .A(n2044), .B(n2045), .Z(n2046) );
  XNOR U2045 ( .A(n2047), .B(n2046), .Z(n1979) );
  NAND U2046 ( .A(n2029), .B(n2186), .Z(n1836) );
  NAND U2047 ( .A(n1834), .B(n1833), .Z(n1835) );
  AND U2048 ( .A(n1836), .B(n1835), .Z(n2053) );
  NAND U2049 ( .A(y[10]), .B(x[15]), .Z(n2036) );
  NAND U2050 ( .A(x[18]), .B(y[7]), .Z(n2034) );
  NAND U2051 ( .A(x[6]), .B(y[19]), .Z(n2035) );
  XNOR U2052 ( .A(n2034), .B(n2035), .Z(n2037) );
  XOR U2053 ( .A(n2036), .B(n2037), .Z(n2051) );
  NAND U2054 ( .A(x[23]), .B(y[2]), .Z(n2018) );
  NAND U2055 ( .A(y[21]), .B(x[4]), .Z(n2016) );
  NAND U2056 ( .A(y[9]), .B(x[16]), .Z(n2017) );
  XNOR U2057 ( .A(n2016), .B(n2017), .Z(n2019) );
  XOR U2058 ( .A(n2018), .B(n2019), .Z(n2050) );
  XOR U2059 ( .A(n2051), .B(n2050), .Z(n2052) );
  XOR U2060 ( .A(n2053), .B(n2052), .Z(n1978) );
  XOR U2061 ( .A(n1979), .B(n1978), .Z(n1980) );
  XNOR U2062 ( .A(n1981), .B(n1980), .Z(n1993) );
  NAND U2063 ( .A(n1838), .B(n1837), .Z(n1842) );
  NAND U2064 ( .A(n1840), .B(n1839), .Z(n1841) );
  NAND U2065 ( .A(n1842), .B(n1841), .Z(n1991) );
  NAND U2066 ( .A(n1844), .B(n1843), .Z(n1848) );
  NAND U2067 ( .A(n1846), .B(n1845), .Z(n1847) );
  NAND U2068 ( .A(n1848), .B(n1847), .Z(n1990) );
  XOR U2069 ( .A(n1991), .B(n1990), .Z(n1992) );
  XOR U2070 ( .A(n1993), .B(n1992), .Z(n1954) );
  XNOR U2071 ( .A(n1955), .B(n1954), .Z(n1946) );
  NANDN U2072 ( .A(n1850), .B(n1849), .Z(n1854) );
  NAND U2073 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U2074 ( .A(n1854), .B(n1853), .Z(n1948) );
  XOR U2075 ( .A(n1949), .B(n1948), .Z(n1943) );
  NANDN U2076 ( .A(n1963), .B(n1855), .Z(n1859) );
  NAND U2077 ( .A(n1857), .B(n1856), .Z(n1858) );
  NAND U2078 ( .A(n1859), .B(n1858), .Z(n1985) );
  AND U2079 ( .A(y[16]), .B(x[14]), .Z(n2894) );
  NAND U2080 ( .A(n2894), .B(n1860), .Z(n1864) );
  NAND U2081 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U2082 ( .A(n1864), .B(n1863), .Z(n2012) );
  NAND U2083 ( .A(x[11]), .B(y[14]), .Z(n2027) );
  NAND U2084 ( .A(y[13]), .B(x[12]), .Z(n2025) );
  NAND U2085 ( .A(y[18]), .B(x[7]), .Z(n2026) );
  XOR U2086 ( .A(n2025), .B(n2026), .Z(n2028) );
  XNOR U2087 ( .A(n2027), .B(n2028), .Z(n2011) );
  NAND U2088 ( .A(x[24]), .B(y[1]), .Z(n2024) );
  XNOR U2089 ( .A(o[25]), .B(n2024), .Z(n1999) );
  AND U2090 ( .A(x[1]), .B(y[24]), .Z(n1998) );
  XOR U2091 ( .A(n1999), .B(n1998), .Z(n2001) );
  AND U2092 ( .A(x[13]), .B(y[12]), .Z(n2000) );
  XOR U2093 ( .A(n2001), .B(n2000), .Z(n2010) );
  XOR U2094 ( .A(n2011), .B(n2010), .Z(n2013) );
  XOR U2095 ( .A(n2012), .B(n2013), .Z(n1984) );
  XOR U2096 ( .A(n1985), .B(n1984), .Z(n1987) );
  NAND U2097 ( .A(n1866), .B(n1865), .Z(n1870) );
  ANDN U2098 ( .B(n1868), .A(n1867), .Z(n1869) );
  ANDN U2099 ( .B(n1870), .A(n1869), .Z(n1973) );
  AND U2100 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U2101 ( .A(n1874), .B(n1873), .Z(n1875) );
  NANDN U2102 ( .A(n1876), .B(n1875), .Z(n1972) );
  NANDN U2103 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2104 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U2105 ( .A(n1882), .B(n1881), .Z(n1969) );
  NAND U2106 ( .A(x[8]), .B(y[17]), .Z(n1964) );
  XNOR U2107 ( .A(n1962), .B(n1963), .Z(n1965) );
  XOR U2108 ( .A(n1964), .B(n1965), .Z(n1967) );
  ANDN U2109 ( .B(o[24]), .A(n1883), .Z(n1960) );
  NAND U2110 ( .A(y[0]), .B(x[25]), .Z(n1958) );
  NAND U2111 ( .A(x[0]), .B(y[25]), .Z(n1959) );
  XNOR U2112 ( .A(n1958), .B(n1959), .Z(n1961) );
  XNOR U2113 ( .A(n1960), .B(n1961), .Z(n1966) );
  XOR U2114 ( .A(n1967), .B(n1966), .Z(n1968) );
  XOR U2115 ( .A(n1975), .B(n1974), .Z(n1986) );
  XNOR U2116 ( .A(n1987), .B(n1986), .Z(n2065) );
  AND U2117 ( .A(n1885), .B(n1884), .Z(n1889) );
  NAND U2118 ( .A(n1887), .B(n1886), .Z(n1888) );
  NANDN U2119 ( .A(n1889), .B(n1888), .Z(n2041) );
  NAND U2120 ( .A(n1891), .B(n1890), .Z(n1895) );
  NAND U2121 ( .A(n1893), .B(n1892), .Z(n1894) );
  NAND U2122 ( .A(n1895), .B(n1894), .Z(n2039) );
  AND U2123 ( .A(x[14]), .B(y[11]), .Z(n2005) );
  AND U2124 ( .A(y[23]), .B(x[2]), .Z(n2004) );
  XOR U2125 ( .A(n2005), .B(n2004), .Z(n2007) );
  AND U2126 ( .A(x[3]), .B(y[22]), .Z(n2006) );
  XOR U2127 ( .A(n2007), .B(n2006), .Z(n2038) );
  XOR U2128 ( .A(n2039), .B(n2038), .Z(n2040) );
  XNOR U2129 ( .A(n2041), .B(n2040), .Z(n2063) );
  NAND U2130 ( .A(n1897), .B(n1896), .Z(n1901) );
  NAND U2131 ( .A(n1899), .B(n1898), .Z(n1900) );
  AND U2132 ( .A(n1901), .B(n1900), .Z(n2062) );
  XOR U2133 ( .A(n2063), .B(n2062), .Z(n2064) );
  XOR U2134 ( .A(n2065), .B(n2064), .Z(n2056) );
  NAND U2135 ( .A(n1903), .B(n1902), .Z(n1907) );
  NAND U2136 ( .A(n1905), .B(n1904), .Z(n1906) );
  AND U2137 ( .A(n1907), .B(n1906), .Z(n2057) );
  XOR U2138 ( .A(n2056), .B(n2057), .Z(n2059) );
  NAND U2139 ( .A(n1909), .B(n1908), .Z(n1913) );
  NAND U2140 ( .A(n1911), .B(n1910), .Z(n1912) );
  AND U2141 ( .A(n1913), .B(n1912), .Z(n2058) );
  XOR U2142 ( .A(n2059), .B(n2058), .Z(n1941) );
  NANDN U2143 ( .A(n1915), .B(n1914), .Z(n1919) );
  NANDN U2144 ( .A(n1917), .B(n1916), .Z(n1918) );
  AND U2145 ( .A(n1919), .B(n1918), .Z(n1940) );
  NAND U2146 ( .A(n1921), .B(n1920), .Z(n1925) );
  NAND U2147 ( .A(n1923), .B(n1922), .Z(n1924) );
  NAND U2148 ( .A(n1925), .B(n1924), .Z(n2071) );
  XNOR U2149 ( .A(n2074), .B(n2073), .Z(n2070) );
  NANDN U2150 ( .A(n1926), .B(n1927), .Z(n1932) );
  NOR U2151 ( .A(n1928), .B(n1927), .Z(n1930) );
  OR U2152 ( .A(n1930), .B(n1929), .Z(n1931) );
  AND U2153 ( .A(n1932), .B(n1931), .Z(n2069) );
  NANDN U2154 ( .A(n1934), .B(n1933), .Z(n1938) );
  NANDN U2155 ( .A(n1936), .B(n1935), .Z(n1937) );
  AND U2156 ( .A(n1938), .B(n1937), .Z(n2068) );
  XOR U2157 ( .A(n2069), .B(n2068), .Z(n1939) );
  XNOR U2158 ( .A(n2070), .B(n1939), .Z(N58) );
  NANDN U2159 ( .A(n1941), .B(n1940), .Z(n1945) );
  NANDN U2160 ( .A(n1943), .B(n1942), .Z(n1944) );
  AND U2161 ( .A(n1945), .B(n1944), .Z(n2211) );
  NANDN U2162 ( .A(n1947), .B(n1946), .Z(n1951) );
  NAND U2163 ( .A(n1949), .B(n1948), .Z(n1950) );
  AND U2164 ( .A(n1951), .B(n1950), .Z(n2210) );
  NAND U2165 ( .A(n1953), .B(n1952), .Z(n1957) );
  NAND U2166 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U2167 ( .A(n1957), .B(n1956), .Z(n2087) );
  AND U2168 ( .A(x[2]), .B(y[24]), .Z(n2104) );
  XOR U2169 ( .A(n2105), .B(n2104), .Z(n2107) );
  AND U2170 ( .A(x[24]), .B(y[2]), .Z(n2106) );
  XOR U2171 ( .A(n2107), .B(n2106), .Z(n2139) );
  XOR U2172 ( .A(n2139), .B(n2138), .Z(n2141) );
  XOR U2173 ( .A(n2141), .B(n2140), .Z(n2199) );
  NAND U2174 ( .A(n1967), .B(n1966), .Z(n1971) );
  NANDN U2175 ( .A(n1969), .B(n1968), .Z(n1970) );
  AND U2176 ( .A(n1971), .B(n1970), .Z(n2198) );
  NANDN U2177 ( .A(n1973), .B(n1972), .Z(n1977) );
  NAND U2178 ( .A(n1975), .B(n1974), .Z(n1976) );
  NAND U2179 ( .A(n1977), .B(n1976), .Z(n2201) );
  NAND U2180 ( .A(n1979), .B(n1978), .Z(n1983) );
  NAND U2181 ( .A(n1981), .B(n1980), .Z(n1982) );
  NAND U2182 ( .A(n1983), .B(n1982), .Z(n2163) );
  NAND U2183 ( .A(n1985), .B(n1984), .Z(n1989) );
  NAND U2184 ( .A(n1987), .B(n1986), .Z(n1988) );
  AND U2185 ( .A(n1989), .B(n1988), .Z(n2162) );
  XOR U2186 ( .A(n2163), .B(n2162), .Z(n2164) );
  XNOR U2187 ( .A(n2165), .B(n2164), .Z(n2085) );
  NAND U2188 ( .A(n1991), .B(n1990), .Z(n1995) );
  NAND U2189 ( .A(n1993), .B(n1992), .Z(n1994) );
  NAND U2190 ( .A(n1995), .B(n1994), .Z(n2093) );
  AND U2191 ( .A(x[12]), .B(y[14]), .Z(n2335) );
  AND U2192 ( .A(y[21]), .B(x[5]), .Z(n2149) );
  XOR U2193 ( .A(n2335), .B(n2149), .Z(n2151) );
  AND U2194 ( .A(y[16]), .B(x[10]), .Z(n2150) );
  XOR U2195 ( .A(n2151), .B(n2150), .Z(n2171) );
  AND U2196 ( .A(x[7]), .B(y[19]), .Z(n2169) );
  AND U2197 ( .A(y[20]), .B(x[6]), .Z(n1997) );
  NAND U2198 ( .A(x[8]), .B(y[18]), .Z(n1996) );
  XNOR U2199 ( .A(n1997), .B(n1996), .Z(n2188) );
  AND U2200 ( .A(y[17]), .B(x[9]), .Z(n2187) );
  XOR U2201 ( .A(n2188), .B(n2187), .Z(n2168) );
  XOR U2202 ( .A(n2169), .B(n2168), .Z(n2170) );
  XOR U2203 ( .A(n2171), .B(n2170), .Z(n2128) );
  NAND U2204 ( .A(n1999), .B(n1998), .Z(n2003) );
  NAND U2205 ( .A(n2001), .B(n2000), .Z(n2002) );
  NAND U2206 ( .A(n2003), .B(n2002), .Z(n2127) );
  NAND U2207 ( .A(n2005), .B(n2004), .Z(n2009) );
  NAND U2208 ( .A(n2007), .B(n2006), .Z(n2008) );
  NAND U2209 ( .A(n2009), .B(n2008), .Z(n2126) );
  XOR U2210 ( .A(n2127), .B(n2126), .Z(n2129) );
  XNOR U2211 ( .A(n2128), .B(n2129), .Z(n2157) );
  NAND U2212 ( .A(n2011), .B(n2010), .Z(n2015) );
  NAND U2213 ( .A(n2013), .B(n2012), .Z(n2014) );
  AND U2214 ( .A(n2015), .B(n2014), .Z(n2156) );
  XOR U2215 ( .A(n2157), .B(n2156), .Z(n2159) );
  XOR U2216 ( .A(n2097), .B(n2096), .Z(n2099) );
  ANDN U2217 ( .B(o[25]), .A(n2024), .Z(n2180) );
  NAND U2218 ( .A(y[12]), .B(x[14]), .Z(n2181) );
  NAND U2219 ( .A(x[1]), .B(y[25]), .Z(n2183) );
  NAND U2220 ( .A(y[1]), .B(x[25]), .Z(n2189) );
  AND U2221 ( .A(y[0]), .B(x[26]), .Z(n2152) );
  XOR U2222 ( .A(n2153), .B(n2152), .Z(n2155) );
  AND U2223 ( .A(y[26]), .B(x[0]), .Z(n2154) );
  XOR U2224 ( .A(n2155), .B(n2154), .Z(n2142) );
  XOR U2225 ( .A(n2143), .B(n2142), .Z(n2145) );
  XOR U2226 ( .A(n2145), .B(n2144), .Z(n2098) );
  XNOR U2227 ( .A(n2099), .B(n2098), .Z(n2135) );
  AND U2228 ( .A(y[5]), .B(x[21]), .Z(n2174) );
  NAND U2229 ( .A(n2029), .B(n2174), .Z(n2033) );
  NAND U2230 ( .A(n2031), .B(n2030), .Z(n2032) );
  NAND U2231 ( .A(n2033), .B(n2032), .Z(n2122) );
  XOR U2232 ( .A(n2175), .B(n2174), .Z(n2176) );
  NAND U2233 ( .A(y[6]), .B(x[20]), .Z(n2177) );
  XNOR U2234 ( .A(n2176), .B(n2177), .Z(n2121) );
  AND U2235 ( .A(x[23]), .B(y[3]), .Z(n2110) );
  XOR U2236 ( .A(n2111), .B(n2110), .Z(n2113) );
  AND U2237 ( .A(x[22]), .B(y[4]), .Z(n2112) );
  XOR U2238 ( .A(n2113), .B(n2112), .Z(n2120) );
  XOR U2239 ( .A(n2121), .B(n2120), .Z(n2123) );
  XNOR U2240 ( .A(n2122), .B(n2123), .Z(n2133) );
  AND U2241 ( .A(x[3]), .B(y[23]), .Z(n2190) );
  NAND U2242 ( .A(x[11]), .B(y[15]), .Z(n2191) );
  NAND U2243 ( .A(x[19]), .B(y[7]), .Z(n2193) );
  NAND U2244 ( .A(y[22]), .B(x[4]), .Z(n2115) );
  XNOR U2245 ( .A(n2114), .B(n2115), .Z(n2117) );
  XOR U2246 ( .A(n2117), .B(n2116), .Z(n2100) );
  XOR U2247 ( .A(n2101), .B(n2100), .Z(n2103) );
  XNOR U2248 ( .A(n2103), .B(n2102), .Z(n2132) );
  XOR U2249 ( .A(n2133), .B(n2132), .Z(n2134) );
  XOR U2250 ( .A(n2135), .B(n2134), .Z(n2158) );
  XNOR U2251 ( .A(n2159), .B(n2158), .Z(n2091) );
  NAND U2252 ( .A(n2039), .B(n2038), .Z(n2043) );
  NAND U2253 ( .A(n2041), .B(n2040), .Z(n2042) );
  AND U2254 ( .A(n2043), .B(n2042), .Z(n2207) );
  NAND U2255 ( .A(n2045), .B(n2044), .Z(n2049) );
  NAND U2256 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2257 ( .A(n2049), .B(n2048), .Z(n2205) );
  NAND U2258 ( .A(n2051), .B(n2050), .Z(n2055) );
  NANDN U2259 ( .A(n2053), .B(n2052), .Z(n2054) );
  NAND U2260 ( .A(n2055), .B(n2054), .Z(n2204) );
  XOR U2261 ( .A(n2091), .B(n2090), .Z(n2092) );
  XOR U2262 ( .A(n2093), .B(n2092), .Z(n2084) );
  XOR U2263 ( .A(n2085), .B(n2084), .Z(n2086) );
  XOR U2264 ( .A(n2087), .B(n2086), .Z(n2081) );
  NAND U2265 ( .A(n2057), .B(n2056), .Z(n2061) );
  NAND U2266 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2267 ( .A(n2061), .B(n2060), .Z(n2078) );
  NAND U2268 ( .A(n2063), .B(n2062), .Z(n2067) );
  NAND U2269 ( .A(n2065), .B(n2064), .Z(n2066) );
  AND U2270 ( .A(n2067), .B(n2066), .Z(n2079) );
  XOR U2271 ( .A(n2078), .B(n2079), .Z(n2080) );
  XOR U2272 ( .A(n2081), .B(n2080), .Z(n2212) );
  XNOR U2273 ( .A(n2213), .B(n2212), .Z(n2218) );
  NANDN U2274 ( .A(n2072), .B(n2071), .Z(n2076) );
  NAND U2275 ( .A(n2074), .B(n2073), .Z(n2075) );
  AND U2276 ( .A(n2076), .B(n2075), .Z(n2216) );
  XOR U2277 ( .A(n2217), .B(n2216), .Z(n2077) );
  XNOR U2278 ( .A(n2218), .B(n2077), .Z(N59) );
  NAND U2279 ( .A(n2079), .B(n2078), .Z(n2083) );
  NAND U2280 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U2281 ( .A(n2083), .B(n2082), .Z(n2223) );
  NAND U2282 ( .A(n2085), .B(n2084), .Z(n2089) );
  NAND U2283 ( .A(n2087), .B(n2086), .Z(n2088) );
  AND U2284 ( .A(n2089), .B(n2088), .Z(n2221) );
  NAND U2285 ( .A(n2091), .B(n2090), .Z(n2095) );
  NAND U2286 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2287 ( .A(n2095), .B(n2094), .Z(n2231) );
  AND U2288 ( .A(n2105), .B(n2104), .Z(n2109) );
  NAND U2289 ( .A(n2107), .B(n2106), .Z(n2108) );
  NANDN U2290 ( .A(n2109), .B(n2108), .Z(n2308) );
  XOR U2291 ( .A(n2308), .B(n2307), .Z(n2309) );
  NANDN U2292 ( .A(n2115), .B(n2114), .Z(n2119) );
  NAND U2293 ( .A(n2117), .B(n2116), .Z(n2118) );
  NAND U2294 ( .A(n2119), .B(n2118), .Z(n2321) );
  AND U2295 ( .A(x[0]), .B(y[27]), .Z(n2287) );
  AND U2296 ( .A(y[0]), .B(x[27]), .Z(n2286) );
  XOR U2297 ( .A(n2287), .B(n2286), .Z(n2289) );
  AND U2298 ( .A(y[1]), .B(x[26]), .Z(n2298) );
  XOR U2299 ( .A(n2298), .B(o[27]), .Z(n2288) );
  XOR U2300 ( .A(n2289), .B(n2288), .Z(n2320) );
  AND U2301 ( .A(y[18]), .B(x[9]), .Z(n2293) );
  AND U2302 ( .A(y[6]), .B(x[21]), .Z(n2292) );
  XOR U2303 ( .A(n2293), .B(n2292), .Z(n2295) );
  AND U2304 ( .A(y[9]), .B(x[18]), .Z(n2294) );
  XOR U2305 ( .A(n2295), .B(n2294), .Z(n2319) );
  XOR U2306 ( .A(n2320), .B(n2319), .Z(n2322) );
  XNOR U2307 ( .A(n2321), .B(n2322), .Z(n2310) );
  XOR U2308 ( .A(n2251), .B(n2252), .Z(n2254) );
  XOR U2309 ( .A(n2253), .B(n2254), .Z(n2367) );
  NAND U2310 ( .A(n2121), .B(n2120), .Z(n2125) );
  NAND U2311 ( .A(n2123), .B(n2122), .Z(n2124) );
  AND U2312 ( .A(n2125), .B(n2124), .Z(n2365) );
  NAND U2313 ( .A(n2127), .B(n2126), .Z(n2131) );
  NAND U2314 ( .A(n2129), .B(n2128), .Z(n2130) );
  AND U2315 ( .A(n2131), .B(n2130), .Z(n2364) );
  XOR U2316 ( .A(n2365), .B(n2364), .Z(n2366) );
  NAND U2317 ( .A(n2133), .B(n2132), .Z(n2137) );
  NAND U2318 ( .A(n2135), .B(n2134), .Z(n2136) );
  AND U2319 ( .A(n2137), .B(n2136), .Z(n2352) );
  AND U2320 ( .A(y[8]), .B(x[19]), .Z(n2275) );
  AND U2321 ( .A(y[2]), .B(x[25]), .Z(n2274) );
  XOR U2322 ( .A(n2275), .B(n2274), .Z(n2277) );
  AND U2323 ( .A(x[6]), .B(y[21]), .Z(n2276) );
  XOR U2324 ( .A(n2277), .B(n2276), .Z(n2264) );
  AND U2325 ( .A(y[12]), .B(x[15]), .Z(n2341) );
  AND U2326 ( .A(x[2]), .B(y[25]), .Z(n2340) );
  XOR U2327 ( .A(n2341), .B(n2340), .Z(n2343) );
  AND U2328 ( .A(x[3]), .B(y[24]), .Z(n2342) );
  XOR U2329 ( .A(n2343), .B(n2342), .Z(n2263) );
  XOR U2330 ( .A(n2264), .B(n2263), .Z(n2265) );
  NAND U2331 ( .A(y[11]), .B(x[16]), .Z(n2325) );
  XOR U2332 ( .A(n2325), .B(n2146), .Z(n2328) );
  XOR U2333 ( .A(n2327), .B(n2328), .Z(n2337) );
  AND U2334 ( .A(y[15]), .B(x[12]), .Z(n2148) );
  AND U2335 ( .A(y[14]), .B(x[13]), .Z(n2147) );
  XOR U2336 ( .A(n2148), .B(n2147), .Z(n2336) );
  XNOR U2337 ( .A(n2265), .B(n2266), .Z(n2304) );
  XOR U2338 ( .A(n2302), .B(n2301), .Z(n2303) );
  XOR U2339 ( .A(n2304), .B(n2303), .Z(n2247) );
  XNOR U2340 ( .A(n2248), .B(n2247), .Z(n2250) );
  XOR U2341 ( .A(n2249), .B(n2250), .Z(n2353) );
  NAND U2342 ( .A(n2157), .B(n2156), .Z(n2161) );
  NAND U2343 ( .A(n2159), .B(n2158), .Z(n2160) );
  AND U2344 ( .A(n2161), .B(n2160), .Z(n2354) );
  XOR U2345 ( .A(n2355), .B(n2354), .Z(n2229) );
  XNOR U2346 ( .A(n2230), .B(n2229), .Z(n2232) );
  XOR U2347 ( .A(n2231), .B(n2232), .Z(n2237) );
  NAND U2348 ( .A(n2163), .B(n2162), .Z(n2167) );
  NAND U2349 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2350 ( .A(n2167), .B(n2166), .Z(n2236) );
  NAND U2351 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2352 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2353 ( .A(n2173), .B(n2172), .Z(n2360) );
  AND U2354 ( .A(n2175), .B(n2174), .Z(n2179) );
  NANDN U2355 ( .A(n2177), .B(n2176), .Z(n2178) );
  NANDN U2356 ( .A(n2179), .B(n2178), .Z(n2255) );
  NANDN U2357 ( .A(n2181), .B(n2180), .Z(n2185) );
  NANDN U2358 ( .A(n2183), .B(n2182), .Z(n2184) );
  NAND U2359 ( .A(n2185), .B(n2184), .Z(n2256) );
  XOR U2360 ( .A(n2255), .B(n2256), .Z(n2257) );
  AND U2361 ( .A(y[20]), .B(x[8]), .Z(n2300) );
  AND U2362 ( .A(x[14]), .B(y[13]), .Z(n2347) );
  AND U2363 ( .A(y[26]), .B(x[1]), .Z(n2346) );
  XOR U2364 ( .A(n2347), .B(n2346), .Z(n2349) );
  ANDN U2365 ( .B(o[26]), .A(n2189), .Z(n2348) );
  XOR U2366 ( .A(n2349), .B(n2348), .Z(n2314) );
  AND U2367 ( .A(x[17]), .B(y[10]), .Z(n2281) );
  AND U2368 ( .A(y[23]), .B(x[4]), .Z(n2280) );
  XOR U2369 ( .A(n2281), .B(n2280), .Z(n2283) );
  AND U2370 ( .A(y[22]), .B(x[5]), .Z(n2282) );
  XOR U2371 ( .A(n2283), .B(n2282), .Z(n2313) );
  XOR U2372 ( .A(n2314), .B(n2313), .Z(n2316) );
  XNOR U2373 ( .A(n2315), .B(n2316), .Z(n2258) );
  XNOR U2374 ( .A(n2257), .B(n2258), .Z(n2358) );
  NANDN U2375 ( .A(n2191), .B(n2190), .Z(n2195) );
  NANDN U2376 ( .A(n2193), .B(n2192), .Z(n2194) );
  NAND U2377 ( .A(n2195), .B(n2194), .Z(n2262) );
  NAND U2378 ( .A(y[3]), .B(x[24]), .Z(n2196) );
  XNOR U2379 ( .A(n2197), .B(n2196), .Z(n2271) );
  AND U2380 ( .A(x[7]), .B(y[20]), .Z(n2270) );
  XOR U2381 ( .A(n2271), .B(n2270), .Z(n2260) );
  AND U2382 ( .A(x[8]), .B(y[19]), .Z(n2330) );
  AND U2383 ( .A(x[23]), .B(y[4]), .Z(n2329) );
  XOR U2384 ( .A(n2330), .B(n2329), .Z(n2332) );
  AND U2385 ( .A(y[5]), .B(x[22]), .Z(n2331) );
  XOR U2386 ( .A(n2332), .B(n2331), .Z(n2259) );
  XOR U2387 ( .A(n2260), .B(n2259), .Z(n2261) );
  XNOR U2388 ( .A(n2262), .B(n2261), .Z(n2359) );
  XNOR U2389 ( .A(n2358), .B(n2359), .Z(n2361) );
  XOR U2390 ( .A(n2360), .B(n2361), .Z(n2242) );
  NANDN U2391 ( .A(n2199), .B(n2198), .Z(n2203) );
  NANDN U2392 ( .A(n2201), .B(n2200), .Z(n2202) );
  NAND U2393 ( .A(n2203), .B(n2202), .Z(n2241) );
  NANDN U2394 ( .A(n2205), .B(n2204), .Z(n2209) );
  NANDN U2395 ( .A(n2207), .B(n2206), .Z(n2208) );
  AND U2396 ( .A(n2209), .B(n2208), .Z(n2243) );
  XOR U2397 ( .A(n2244), .B(n2243), .Z(n2235) );
  XOR U2398 ( .A(n2236), .B(n2235), .Z(n2238) );
  XOR U2399 ( .A(n2237), .B(n2238), .Z(n2220) );
  XOR U2400 ( .A(n2221), .B(n2220), .Z(n2222) );
  XOR U2401 ( .A(n2223), .B(n2222), .Z(n2228) );
  NANDN U2402 ( .A(n2211), .B(n2210), .Z(n2215) );
  NAND U2403 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2404 ( .A(n2215), .B(n2214), .Z(n2226) );
  XOR U2405 ( .A(n2226), .B(n2227), .Z(n2219) );
  XNOR U2406 ( .A(n2228), .B(n2219), .Z(N60) );
  NAND U2407 ( .A(n2221), .B(n2220), .Z(n2225) );
  NAND U2408 ( .A(n2223), .B(n2222), .Z(n2224) );
  NAND U2409 ( .A(n2225), .B(n2224), .Z(n2535) );
  IV U2410 ( .A(n2535), .Z(n2533) );
  NAND U2411 ( .A(n2230), .B(n2229), .Z(n2234) );
  NANDN U2412 ( .A(n2232), .B(n2231), .Z(n2233) );
  NAND U2413 ( .A(n2234), .B(n2233), .Z(n2528) );
  NAND U2414 ( .A(n2236), .B(n2235), .Z(n2240) );
  NAND U2415 ( .A(n2238), .B(n2237), .Z(n2239) );
  AND U2416 ( .A(n2240), .B(n2239), .Z(n2527) );
  XOR U2417 ( .A(n2528), .B(n2527), .Z(n2530) );
  NANDN U2418 ( .A(n2242), .B(n2241), .Z(n2246) );
  NAND U2419 ( .A(n2244), .B(n2243), .Z(n2245) );
  AND U2420 ( .A(n2246), .B(n2245), .Z(n2372) );
  XOR U2421 ( .A(n2383), .B(n2384), .Z(n2386) );
  NAND U2422 ( .A(n2264), .B(n2263), .Z(n2268) );
  NANDN U2423 ( .A(n2266), .B(n2265), .Z(n2267) );
  NAND U2424 ( .A(n2268), .B(n2267), .Z(n2485) );
  XOR U2425 ( .A(n2486), .B(n2485), .Z(n2488) );
  XOR U2426 ( .A(n2487), .B(n2488), .Z(n2387) );
  AND U2427 ( .A(x[24]), .B(y[7]), .Z(n2878) );
  AND U2428 ( .A(x[20]), .B(y[3]), .Z(n2269) );
  NAND U2429 ( .A(n2878), .B(n2269), .Z(n2273) );
  NAND U2430 ( .A(n2271), .B(n2270), .Z(n2272) );
  NAND U2431 ( .A(n2273), .B(n2272), .Z(n2523) );
  AND U2432 ( .A(y[3]), .B(x[25]), .Z(n2436) );
  XOR U2433 ( .A(n2437), .B(n2436), .Z(n2435) );
  AND U2434 ( .A(y[27]), .B(x[1]), .Z(n2434) );
  XOR U2435 ( .A(n2435), .B(n2434), .Z(n2522) );
  AND U2436 ( .A(y[12]), .B(x[16]), .Z(n2429) );
  AND U2437 ( .A(x[24]), .B(y[4]), .Z(n2428) );
  XOR U2438 ( .A(n2429), .B(n2428), .Z(n2431) );
  AND U2439 ( .A(y[26]), .B(x[2]), .Z(n2430) );
  XOR U2440 ( .A(n2431), .B(n2430), .Z(n2521) );
  XOR U2441 ( .A(n2522), .B(n2521), .Z(n2524) );
  XOR U2442 ( .A(n2523), .B(n2524), .Z(n2494) );
  NAND U2443 ( .A(n2275), .B(n2274), .Z(n2279) );
  NAND U2444 ( .A(n2277), .B(n2276), .Z(n2278) );
  NAND U2445 ( .A(n2279), .B(n2278), .Z(n2517) );
  AND U2446 ( .A(x[3]), .B(y[25]), .Z(n2468) );
  XOR U2447 ( .A(n2468), .B(n2467), .Z(n2470) );
  AND U2448 ( .A(y[5]), .B(x[23]), .Z(n2469) );
  XOR U2449 ( .A(n2470), .B(n2469), .Z(n2516) );
  AND U2450 ( .A(y[23]), .B(x[5]), .Z(n2452) );
  AND U2451 ( .A(x[21]), .B(y[7]), .Z(n2451) );
  XOR U2452 ( .A(n2452), .B(n2451), .Z(n2454) );
  AND U2453 ( .A(x[20]), .B(y[8]), .Z(n2453) );
  XOR U2454 ( .A(n2454), .B(n2453), .Z(n2515) );
  XOR U2455 ( .A(n2516), .B(n2515), .Z(n2518) );
  XOR U2456 ( .A(n2517), .B(n2518), .Z(n2492) );
  NAND U2457 ( .A(n2281), .B(n2280), .Z(n2285) );
  NAND U2458 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U2459 ( .A(n2285), .B(n2284), .Z(n2510) );
  NAND U2460 ( .A(n2287), .B(n2286), .Z(n2291) );
  NAND U2461 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2462 ( .A(n2291), .B(n2290), .Z(n2509) );
  XOR U2463 ( .A(n2510), .B(n2509), .Z(n2512) );
  NAND U2464 ( .A(n2293), .B(n2292), .Z(n2297) );
  NAND U2465 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2466 ( .A(n2297), .B(n2296), .Z(n2407) );
  AND U2467 ( .A(n2298), .B(o[27]), .Z(n2420) );
  AND U2468 ( .A(x[0]), .B(y[28]), .Z(n2418) );
  AND U2469 ( .A(y[0]), .B(x[28]), .Z(n2417) );
  XOR U2470 ( .A(n2418), .B(n2417), .Z(n2419) );
  XOR U2471 ( .A(n2420), .B(n2419), .Z(n2406) );
  NAND U2472 ( .A(x[10]), .B(y[18]), .Z(n2299) );
  XNOR U2473 ( .A(n2300), .B(n2299), .Z(n2425) );
  AND U2474 ( .A(y[19]), .B(x[9]), .Z(n2424) );
  XOR U2475 ( .A(n2425), .B(n2424), .Z(n2405) );
  XOR U2476 ( .A(n2406), .B(n2405), .Z(n2408) );
  XOR U2477 ( .A(n2407), .B(n2408), .Z(n2511) );
  XNOR U2478 ( .A(n2512), .B(n2511), .Z(n2491) );
  NAND U2479 ( .A(n2302), .B(n2301), .Z(n2306) );
  NAND U2480 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U2481 ( .A(n2306), .B(n2305), .Z(n2393) );
  NAND U2482 ( .A(n2308), .B(n2307), .Z(n2312) );
  NANDN U2483 ( .A(n2310), .B(n2309), .Z(n2311) );
  NAND U2484 ( .A(n2312), .B(n2311), .Z(n2499) );
  NAND U2485 ( .A(n2314), .B(n2313), .Z(n2318) );
  NAND U2486 ( .A(n2316), .B(n2315), .Z(n2317) );
  NAND U2487 ( .A(n2318), .B(n2317), .Z(n2498) );
  NAND U2488 ( .A(n2320), .B(n2319), .Z(n2324) );
  NAND U2489 ( .A(n2322), .B(n2321), .Z(n2323) );
  NAND U2490 ( .A(n2324), .B(n2323), .Z(n2497) );
  XOR U2491 ( .A(n2498), .B(n2497), .Z(n2500) );
  XOR U2492 ( .A(n2499), .B(n2500), .Z(n2394) );
  XOR U2493 ( .A(n2393), .B(n2394), .Z(n2396) );
  AND U2494 ( .A(x[7]), .B(y[21]), .Z(n2441) );
  AND U2495 ( .A(y[16]), .B(x[12]), .Z(n2440) );
  XOR U2496 ( .A(n2441), .B(n2440), .Z(n2443) );
  AND U2497 ( .A(x[11]), .B(y[17]), .Z(n2442) );
  XOR U2498 ( .A(n2443), .B(n2442), .Z(n2474) );
  AND U2499 ( .A(y[1]), .B(x[27]), .Z(n2457) );
  XOR U2500 ( .A(o[28]), .B(n2457), .Z(n2462) );
  AND U2501 ( .A(x[26]), .B(y[2]), .Z(n2461) );
  XOR U2502 ( .A(n2462), .B(n2461), .Z(n2464) );
  AND U2503 ( .A(y[13]), .B(x[15]), .Z(n2463) );
  XNOR U2504 ( .A(n2464), .B(n2463), .Z(n2473) );
  XOR U2505 ( .A(n2475), .B(n2476), .Z(n2504) );
  NAND U2506 ( .A(n2330), .B(n2329), .Z(n2334) );
  NAND U2507 ( .A(n2332), .B(n2331), .Z(n2333) );
  NAND U2508 ( .A(n2334), .B(n2333), .Z(n2481) );
  AND U2509 ( .A(x[17]), .B(y[11]), .Z(n2412) );
  AND U2510 ( .A(y[6]), .B(x[22]), .Z(n2411) );
  XOR U2511 ( .A(n2412), .B(n2411), .Z(n2414) );
  AND U2512 ( .A(y[24]), .B(x[4]), .Z(n2413) );
  XOR U2513 ( .A(n2414), .B(n2413), .Z(n2480) );
  AND U2514 ( .A(y[22]), .B(x[6]), .Z(n2598) );
  AND U2515 ( .A(y[9]), .B(x[19]), .Z(n2446) );
  XOR U2516 ( .A(n2598), .B(n2446), .Z(n2448) );
  XOR U2517 ( .A(n2448), .B(n2447), .Z(n2479) );
  XOR U2518 ( .A(n2480), .B(n2479), .Z(n2482) );
  XOR U2519 ( .A(n2481), .B(n2482), .Z(n2503) );
  NAND U2520 ( .A(n2467), .B(n2335), .Z(n2339) );
  NANDN U2521 ( .A(n2337), .B(n2336), .Z(n2338) );
  NAND U2522 ( .A(n2339), .B(n2338), .Z(n2401) );
  NAND U2523 ( .A(n2341), .B(n2340), .Z(n2345) );
  NAND U2524 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U2525 ( .A(n2345), .B(n2344), .Z(n2400) );
  NAND U2526 ( .A(n2347), .B(n2346), .Z(n2351) );
  NAND U2527 ( .A(n2349), .B(n2348), .Z(n2350) );
  NAND U2528 ( .A(n2351), .B(n2350), .Z(n2399) );
  XNOR U2529 ( .A(n2400), .B(n2399), .Z(n2402) );
  XNOR U2530 ( .A(n2505), .B(n2506), .Z(n2395) );
  XOR U2531 ( .A(n2396), .B(n2395), .Z(n2389) );
  XOR U2532 ( .A(n2390), .B(n2389), .Z(n2385) );
  XOR U2533 ( .A(n2386), .B(n2385), .Z(n2371) );
  XOR U2534 ( .A(n2372), .B(n2371), .Z(n2373) );
  NANDN U2535 ( .A(n2353), .B(n2352), .Z(n2357) );
  NAND U2536 ( .A(n2355), .B(n2354), .Z(n2356) );
  NAND U2537 ( .A(n2357), .B(n2356), .Z(n2379) );
  NANDN U2538 ( .A(n2359), .B(n2358), .Z(n2363) );
  NAND U2539 ( .A(n2361), .B(n2360), .Z(n2362) );
  NAND U2540 ( .A(n2363), .B(n2362), .Z(n2377) );
  NAND U2541 ( .A(n2365), .B(n2364), .Z(n2369) );
  NANDN U2542 ( .A(n2367), .B(n2366), .Z(n2368) );
  AND U2543 ( .A(n2369), .B(n2368), .Z(n2378) );
  XNOR U2544 ( .A(n2377), .B(n2378), .Z(n2380) );
  XNOR U2545 ( .A(n2373), .B(n2374), .Z(n2529) );
  XOR U2546 ( .A(n2530), .B(n2529), .Z(n2536) );
  XNOR U2547 ( .A(n2534), .B(n2536), .Z(n2370) );
  XOR U2548 ( .A(n2533), .B(n2370), .Z(N61) );
  NAND U2549 ( .A(n2372), .B(n2371), .Z(n2376) );
  NANDN U2550 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U2551 ( .A(n2376), .B(n2375), .Z(n2711) );
  NAND U2552 ( .A(n2378), .B(n2377), .Z(n2382) );
  NANDN U2553 ( .A(n2380), .B(n2379), .Z(n2381) );
  NAND U2554 ( .A(n2382), .B(n2381), .Z(n2709) );
  NANDN U2555 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U2556 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U2557 ( .A(n2392), .B(n2391), .Z(n2542) );
  XOR U2558 ( .A(n2541), .B(n2542), .Z(n2544) );
  NAND U2559 ( .A(n2394), .B(n2393), .Z(n2398) );
  NAND U2560 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U2561 ( .A(n2398), .B(n2397), .Z(n2700) );
  NAND U2562 ( .A(n2400), .B(n2399), .Z(n2404) );
  NANDN U2563 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U2564 ( .A(n2404), .B(n2403), .Z(n2548) );
  NAND U2565 ( .A(n2406), .B(n2405), .Z(n2410) );
  NAND U2566 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U2567 ( .A(n2410), .B(n2409), .Z(n2546) );
  NAND U2568 ( .A(n2412), .B(n2411), .Z(n2416) );
  NAND U2569 ( .A(n2414), .B(n2413), .Z(n2415) );
  NAND U2570 ( .A(n2416), .B(n2415), .Z(n2583) );
  NAND U2571 ( .A(n2418), .B(n2417), .Z(n2422) );
  NAND U2572 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U2573 ( .A(n2422), .B(n2421), .Z(n2582) );
  XOR U2574 ( .A(n2583), .B(n2582), .Z(n2585) );
  AND U2575 ( .A(x[10]), .B(y[20]), .Z(n2581) );
  NAND U2576 ( .A(n2581), .B(n2423), .Z(n2427) );
  NAND U2577 ( .A(n2425), .B(n2424), .Z(n2426) );
  NAND U2578 ( .A(n2427), .B(n2426), .Z(n2553) );
  AND U2579 ( .A(y[17]), .B(x[12]), .Z(n2918) );
  AND U2580 ( .A(y[28]), .B(x[1]), .Z(n2617) );
  XOR U2581 ( .A(n2918), .B(n2617), .Z(n2619) );
  AND U2582 ( .A(x[22]), .B(y[7]), .Z(n2618) );
  XOR U2583 ( .A(n2619), .B(n2618), .Z(n2552) );
  AND U2584 ( .A(y[14]), .B(x[15]), .Z(n2622) );
  XOR U2585 ( .A(n2923), .B(n2622), .Z(n2624) );
  XOR U2586 ( .A(n2624), .B(n2623), .Z(n2551) );
  XOR U2587 ( .A(n2552), .B(n2551), .Z(n2554) );
  XOR U2588 ( .A(n2553), .B(n2554), .Z(n2584) );
  XNOR U2589 ( .A(n2585), .B(n2584), .Z(n2545) );
  XOR U2590 ( .A(n2546), .B(n2545), .Z(n2547) );
  XOR U2591 ( .A(n2548), .B(n2547), .Z(n2684) );
  NAND U2592 ( .A(n2429), .B(n2428), .Z(n2433) );
  NAND U2593 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U2594 ( .A(n2433), .B(n2432), .Z(n2558) );
  AND U2595 ( .A(n2435), .B(n2434), .Z(n2439) );
  NAND U2596 ( .A(n2437), .B(n2436), .Z(n2438) );
  NANDN U2597 ( .A(n2439), .B(n2438), .Z(n2557) );
  XOR U2598 ( .A(n2558), .B(n2557), .Z(n2559) );
  NAND U2599 ( .A(n2441), .B(n2440), .Z(n2445) );
  NAND U2600 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U2601 ( .A(n2445), .B(n2444), .Z(n2632) );
  AND U2602 ( .A(x[3]), .B(y[26]), .Z(n2808) );
  AND U2603 ( .A(y[12]), .B(x[17]), .Z(n2595) );
  XOR U2604 ( .A(n2808), .B(n2595), .Z(n2594) );
  AND U2605 ( .A(y[18]), .B(x[11]), .Z(n2593) );
  XOR U2606 ( .A(n2594), .B(n2593), .Z(n2631) );
  AND U2607 ( .A(x[13]), .B(y[16]), .Z(n2589) );
  AND U2608 ( .A(x[24]), .B(y[5]), .Z(n2588) );
  XOR U2609 ( .A(n2589), .B(n2588), .Z(n2590) );
  AND U2610 ( .A(x[23]), .B(y[6]), .Z(n2818) );
  XOR U2611 ( .A(n2590), .B(n2818), .Z(n2630) );
  XOR U2612 ( .A(n2631), .B(n2630), .Z(n2633) );
  XNOR U2613 ( .A(n2632), .B(n2633), .Z(n2560) );
  NAND U2614 ( .A(n2598), .B(n2446), .Z(n2450) );
  NAND U2615 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U2616 ( .A(n2450), .B(n2449), .Z(n2566) );
  AND U2617 ( .A(x[26]), .B(y[3]), .Z(n2611) );
  XOR U2618 ( .A(n2612), .B(n2611), .Z(n2614) );
  AND U2619 ( .A(y[4]), .B(x[25]), .Z(n2613) );
  XOR U2620 ( .A(n2614), .B(n2613), .Z(n2564) );
  AND U2621 ( .A(y[1]), .B(x[28]), .Z(n2627) );
  XOR U2622 ( .A(o[29]), .B(n2627), .Z(n2575) );
  AND U2623 ( .A(x[0]), .B(y[29]), .Z(n2573) );
  AND U2624 ( .A(x[29]), .B(y[0]), .Z(n2572) );
  XOR U2625 ( .A(n2573), .B(n2572), .Z(n2574) );
  XNOR U2626 ( .A(n2575), .B(n2574), .Z(n2563) );
  XOR U2627 ( .A(n2566), .B(n2565), .Z(n2675) );
  NAND U2628 ( .A(n2452), .B(n2451), .Z(n2456) );
  NAND U2629 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U2630 ( .A(n2456), .B(n2455), .Z(n2607) );
  AND U2631 ( .A(x[2]), .B(y[27]), .Z(n2643) );
  XOR U2632 ( .A(n2643), .B(n2642), .Z(n2644) );
  XOR U2633 ( .A(n2645), .B(n2644), .Z(n2606) );
  AND U2634 ( .A(n2457), .B(o[28]), .Z(n2660) );
  AND U2635 ( .A(y[13]), .B(x[16]), .Z(n2658) );
  AND U2636 ( .A(x[27]), .B(y[2]), .Z(n2657) );
  XOR U2637 ( .A(n2658), .B(n2657), .Z(n2659) );
  XOR U2638 ( .A(n2660), .B(n2659), .Z(n2605) );
  XOR U2639 ( .A(n2606), .B(n2605), .Z(n2608) );
  XOR U2640 ( .A(n2607), .B(n2608), .Z(n2676) );
  AND U2641 ( .A(y[23]), .B(x[6]), .Z(n2459) );
  NAND U2642 ( .A(x[7]), .B(y[22]), .Z(n2458) );
  XNOR U2643 ( .A(n2459), .B(n2458), .Z(n2600) );
  AND U2644 ( .A(x[8]), .B(y[21]), .Z(n2599) );
  XNOR U2645 ( .A(n2600), .B(n2599), .Z(n2570) );
  AND U2646 ( .A(y[20]), .B(x[9]), .Z(n2569) );
  IV U2647 ( .A(n2569), .Z(n2795) );
  XOR U2648 ( .A(n2570), .B(n2795), .Z(n2460) );
  AND U2649 ( .A(x[5]), .B(y[24]), .Z(n2813) );
  AND U2650 ( .A(y[25]), .B(x[4]), .Z(n2653) );
  AND U2651 ( .A(x[10]), .B(y[19]), .Z(n2652) );
  XOR U2652 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U2653 ( .A(n2813), .B(n2654), .Z(n2571) );
  XNOR U2654 ( .A(n2460), .B(n2571), .Z(n2638) );
  NAND U2655 ( .A(n2462), .B(n2461), .Z(n2466) );
  NAND U2656 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U2657 ( .A(n2466), .B(n2465), .Z(n2637) );
  NAND U2658 ( .A(n2468), .B(n2467), .Z(n2472) );
  NAND U2659 ( .A(n2470), .B(n2469), .Z(n2471) );
  NAND U2660 ( .A(n2472), .B(n2471), .Z(n2636) );
  XNOR U2661 ( .A(n2637), .B(n2636), .Z(n2639) );
  NANDN U2662 ( .A(n2474), .B(n2473), .Z(n2478) );
  NAND U2663 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U2664 ( .A(n2478), .B(n2477), .Z(n2663) );
  XNOR U2665 ( .A(n2665), .B(n2666), .Z(n2682) );
  NAND U2666 ( .A(n2480), .B(n2479), .Z(n2484) );
  NAND U2667 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U2668 ( .A(n2484), .B(n2483), .Z(n2681) );
  XOR U2669 ( .A(n2700), .B(n2701), .Z(n2703) );
  NAND U2670 ( .A(n2486), .B(n2485), .Z(n2490) );
  NAND U2671 ( .A(n2488), .B(n2487), .Z(n2489) );
  NAND U2672 ( .A(n2490), .B(n2489), .Z(n2694) );
  NANDN U2673 ( .A(n2492), .B(n2491), .Z(n2496) );
  NANDN U2674 ( .A(n2494), .B(n2493), .Z(n2495) );
  AND U2675 ( .A(n2496), .B(n2495), .Z(n2695) );
  XOR U2676 ( .A(n2694), .B(n2695), .Z(n2697) );
  NAND U2677 ( .A(n2498), .B(n2497), .Z(n2502) );
  NAND U2678 ( .A(n2500), .B(n2499), .Z(n2501) );
  NAND U2679 ( .A(n2502), .B(n2501), .Z(n2690) );
  NANDN U2680 ( .A(n2504), .B(n2503), .Z(n2508) );
  NANDN U2681 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2682 ( .A(n2508), .B(n2507), .Z(n2688) );
  NAND U2683 ( .A(n2510), .B(n2509), .Z(n2514) );
  NAND U2684 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U2685 ( .A(n2514), .B(n2513), .Z(n2671) );
  NAND U2686 ( .A(n2516), .B(n2515), .Z(n2520) );
  NAND U2687 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U2688 ( .A(n2520), .B(n2519), .Z(n2670) );
  NAND U2689 ( .A(n2522), .B(n2521), .Z(n2526) );
  NAND U2690 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U2691 ( .A(n2526), .B(n2525), .Z(n2669) );
  XOR U2692 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U2693 ( .A(n2671), .B(n2672), .Z(n2689) );
  XOR U2694 ( .A(n2688), .B(n2689), .Z(n2691) );
  XOR U2695 ( .A(n2690), .B(n2691), .Z(n2696) );
  XOR U2696 ( .A(n2697), .B(n2696), .Z(n2702) );
  XOR U2697 ( .A(n2703), .B(n2702), .Z(n2543) );
  XOR U2698 ( .A(n2544), .B(n2543), .Z(n2710) );
  XNOR U2699 ( .A(n2709), .B(n2710), .Z(n2712) );
  XOR U2700 ( .A(n2711), .B(n2712), .Z(n2708) );
  NAND U2701 ( .A(n2528), .B(n2527), .Z(n2532) );
  NAND U2702 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U2703 ( .A(n2532), .B(n2531), .Z(n2707) );
  NANDN U2704 ( .A(n2533), .B(n2534), .Z(n2539) );
  NOR U2705 ( .A(n2535), .B(n2534), .Z(n2537) );
  OR U2706 ( .A(n2537), .B(n2536), .Z(n2538) );
  AND U2707 ( .A(n2539), .B(n2538), .Z(n2706) );
  XOR U2708 ( .A(n2707), .B(n2706), .Z(n2540) );
  XNOR U2709 ( .A(n2708), .B(n2540), .Z(N62) );
  NAND U2710 ( .A(n2546), .B(n2545), .Z(n2550) );
  NAND U2711 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U2712 ( .A(n2550), .B(n2549), .Z(n2959) );
  NAND U2713 ( .A(n2552), .B(n2551), .Z(n2556) );
  NAND U2714 ( .A(n2554), .B(n2553), .Z(n2555) );
  AND U2715 ( .A(n2556), .B(n2555), .Z(n2744) );
  NAND U2716 ( .A(n2558), .B(n2557), .Z(n2562) );
  NANDN U2717 ( .A(n2560), .B(n2559), .Z(n2561) );
  AND U2718 ( .A(n2562), .B(n2561), .Z(n2743) );
  XOR U2719 ( .A(n2744), .B(n2743), .Z(n2742) );
  NANDN U2720 ( .A(n2564), .B(n2563), .Z(n2568) );
  OR U2721 ( .A(n2566), .B(n2565), .Z(n2567) );
  NAND U2722 ( .A(n2568), .B(n2567), .Z(n2741) );
  XOR U2723 ( .A(n2742), .B(n2741), .Z(n2962) );
  NAND U2724 ( .A(n2573), .B(n2572), .Z(n2577) );
  NAND U2725 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U2726 ( .A(n2577), .B(n2576), .Z(n2787) );
  AND U2727 ( .A(x[12]), .B(y[18]), .Z(n2579) );
  XOR U2728 ( .A(n2579), .B(n2578), .Z(n2915) );
  XOR U2729 ( .A(n2916), .B(n2915), .Z(n2794) );
  AND U2730 ( .A(x[9]), .B(y[21]), .Z(n2580) );
  XOR U2731 ( .A(n2581), .B(n2580), .Z(n2793) );
  XOR U2732 ( .A(n2794), .B(n2793), .Z(n2790) );
  AND U2733 ( .A(x[27]), .B(y[3]), .Z(n2888) );
  AND U2734 ( .A(x[1]), .B(y[29]), .Z(n2887) );
  XOR U2735 ( .A(n2888), .B(n2887), .Z(n2885) );
  XOR U2736 ( .A(n2886), .B(n2885), .Z(n2789) );
  XOR U2737 ( .A(n2790), .B(n2789), .Z(n2788) );
  XOR U2738 ( .A(n2787), .B(n2788), .Z(n2750) );
  NAND U2739 ( .A(n2583), .B(n2582), .Z(n2587) );
  NAND U2740 ( .A(n2585), .B(n2584), .Z(n2586) );
  AND U2741 ( .A(n2587), .B(n2586), .Z(n2747) );
  XNOR U2742 ( .A(n2748), .B(n2747), .Z(n2961) );
  XNOR U2743 ( .A(n2959), .B(n2960), .Z(n3008) );
  NAND U2744 ( .A(n2589), .B(n2588), .Z(n2592) );
  NAND U2745 ( .A(n2590), .B(n2818), .Z(n2591) );
  NAND U2746 ( .A(n2592), .B(n2591), .Z(n2736) );
  NAND U2747 ( .A(n2594), .B(n2593), .Z(n2597) );
  AND U2748 ( .A(n2808), .B(n2595), .Z(n2596) );
  ANDN U2749 ( .B(n2597), .A(n2596), .Z(n2768) );
  AND U2750 ( .A(x[0]), .B(y[30]), .Z(n2799) );
  AND U2751 ( .A(y[1]), .B(x[29]), .Z(n2876) );
  XOR U2752 ( .A(o[30]), .B(n2876), .Z(n2801) );
  AND U2753 ( .A(y[0]), .B(x[30]), .Z(n2800) );
  XOR U2754 ( .A(n2801), .B(n2800), .Z(n2798) );
  XOR U2755 ( .A(n2799), .B(n2798), .Z(n2770) );
  AND U2756 ( .A(x[20]), .B(y[10]), .Z(n2893) );
  XOR U2757 ( .A(n2894), .B(n2893), .Z(n2892) );
  AND U2758 ( .A(y[22]), .B(x[8]), .Z(n2891) );
  XNOR U2759 ( .A(n2892), .B(n2891), .Z(n2769) );
  XNOR U2760 ( .A(n2768), .B(n2767), .Z(n2735) );
  XOR U2761 ( .A(n2736), .B(n2735), .Z(n2733) );
  AND U2762 ( .A(y[23]), .B(x[7]), .Z(n2922) );
  NAND U2763 ( .A(n2598), .B(n2922), .Z(n2602) );
  NAND U2764 ( .A(n2600), .B(n2599), .Z(n2601) );
  AND U2765 ( .A(n2602), .B(n2601), .Z(n2779) );
  AND U2766 ( .A(x[22]), .B(y[8]), .Z(n2604) );
  AND U2767 ( .A(x[21]), .B(y[9]), .Z(n2603) );
  XOR U2768 ( .A(n2604), .B(n2603), .Z(n2921) );
  XOR U2769 ( .A(n2922), .B(n2921), .Z(n2782) );
  AND U2770 ( .A(x[17]), .B(y[13]), .Z(n2936) );
  AND U2771 ( .A(x[2]), .B(y[28]), .Z(n2938) );
  AND U2772 ( .A(y[4]), .B(x[26]), .Z(n2937) );
  XOR U2773 ( .A(n2938), .B(n2937), .Z(n2935) );
  XNOR U2774 ( .A(n2936), .B(n2935), .Z(n2781) );
  XNOR U2775 ( .A(n2779), .B(n2780), .Z(n2734) );
  NAND U2776 ( .A(n2606), .B(n2605), .Z(n2610) );
  NAND U2777 ( .A(n2608), .B(n2607), .Z(n2609) );
  NAND U2778 ( .A(n2610), .B(n2609), .Z(n2967) );
  XOR U2779 ( .A(n2968), .B(n2967), .Z(n2965) );
  AND U2780 ( .A(n2612), .B(n2611), .Z(n2616) );
  NAND U2781 ( .A(n2614), .B(n2613), .Z(n2615) );
  NANDN U2782 ( .A(n2616), .B(n2615), .Z(n2759) );
  AND U2783 ( .A(n2918), .B(n2617), .Z(n2621) );
  NAND U2784 ( .A(n2619), .B(n2618), .Z(n2620) );
  NANDN U2785 ( .A(n2621), .B(n2620), .Z(n2761) );
  NAND U2786 ( .A(n2923), .B(n2622), .Z(n2626) );
  NAND U2787 ( .A(n2624), .B(n2623), .Z(n2625) );
  AND U2788 ( .A(n2626), .B(n2625), .Z(n2773) );
  AND U2789 ( .A(n2627), .B(o[29]), .Z(n2930) );
  AND U2790 ( .A(y[2]), .B(x[28]), .Z(n2932) );
  AND U2791 ( .A(x[16]), .B(y[14]), .Z(n2931) );
  XOR U2792 ( .A(n2932), .B(n2931), .Z(n2929) );
  XOR U2793 ( .A(n2930), .B(n2929), .Z(n2776) );
  AND U2794 ( .A(y[5]), .B(x[25]), .Z(n2817) );
  AND U2795 ( .A(y[7]), .B(x[23]), .Z(n2629) );
  AND U2796 ( .A(y[6]), .B(x[24]), .Z(n2628) );
  XOR U2797 ( .A(n2629), .B(n2628), .Z(n2816) );
  XNOR U2798 ( .A(n2817), .B(n2816), .Z(n2775) );
  XNOR U2799 ( .A(n2773), .B(n2774), .Z(n2762) );
  XOR U2800 ( .A(n2759), .B(n2760), .Z(n2966) );
  XNOR U2801 ( .A(n2965), .B(n2966), .Z(n2724) );
  NAND U2802 ( .A(n2631), .B(n2630), .Z(n2635) );
  NAND U2803 ( .A(n2633), .B(n2632), .Z(n2634) );
  NAND U2804 ( .A(n2635), .B(n2634), .Z(n2730) );
  NAND U2805 ( .A(n2637), .B(n2636), .Z(n2641) );
  NANDN U2806 ( .A(n2639), .B(n2638), .Z(n2640) );
  NAND U2807 ( .A(n2641), .B(n2640), .Z(n2729) );
  XOR U2808 ( .A(n2730), .B(n2729), .Z(n2728) );
  NAND U2809 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U2810 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U2811 ( .A(n2647), .B(n2646), .Z(n2841) );
  AND U2812 ( .A(x[4]), .B(y[26]), .Z(n2649) );
  NAND U2813 ( .A(y[27]), .B(x[3]), .Z(n2648) );
  XNOR U2814 ( .A(n2649), .B(n2648), .Z(n2807) );
  AND U2815 ( .A(y[12]), .B(x[18]), .Z(n2806) );
  XOR U2816 ( .A(n2807), .B(n2806), .Z(n2844) );
  AND U2817 ( .A(y[25]), .B(x[5]), .Z(n2651) );
  NAND U2818 ( .A(y[24]), .B(x[6]), .Z(n2650) );
  XNOR U2819 ( .A(n2651), .B(n2650), .Z(n2812) );
  AND U2820 ( .A(y[11]), .B(x[19]), .Z(n2811) );
  XOR U2821 ( .A(n2812), .B(n2811), .Z(n2843) );
  XOR U2822 ( .A(n2844), .B(n2843), .Z(n2842) );
  XOR U2823 ( .A(n2841), .B(n2842), .Z(n2756) );
  NAND U2824 ( .A(n2653), .B(n2652), .Z(n2656) );
  NAND U2825 ( .A(n2813), .B(n2654), .Z(n2655) );
  NAND U2826 ( .A(n2656), .B(n2655), .Z(n2755) );
  XOR U2827 ( .A(n2756), .B(n2755), .Z(n2754) );
  NAND U2828 ( .A(n2658), .B(n2657), .Z(n2662) );
  NAND U2829 ( .A(n2660), .B(n2659), .Z(n2661) );
  NAND U2830 ( .A(n2662), .B(n2661), .Z(n2753) );
  XOR U2831 ( .A(n2754), .B(n2753), .Z(n2727) );
  XNOR U2832 ( .A(n2728), .B(n2727), .Z(n2723) );
  NANDN U2833 ( .A(n2664), .B(n2663), .Z(n2668) );
  NANDN U2834 ( .A(n2666), .B(n2665), .Z(n2667) );
  NAND U2835 ( .A(n2668), .B(n2667), .Z(n2721) );
  XOR U2836 ( .A(n2722), .B(n2721), .Z(n2990) );
  NAND U2837 ( .A(n2670), .B(n2669), .Z(n2674) );
  NAND U2838 ( .A(n2672), .B(n2671), .Z(n2673) );
  NAND U2839 ( .A(n2674), .B(n2673), .Z(n2989) );
  NANDN U2840 ( .A(n2676), .B(n2675), .Z(n2680) );
  NANDN U2841 ( .A(n2678), .B(n2677), .Z(n2679) );
  AND U2842 ( .A(n2680), .B(n2679), .Z(n2987) );
  XOR U2843 ( .A(n2988), .B(n2987), .Z(n3006) );
  IV U2844 ( .A(n3006), .Z(n2687) );
  NANDN U2845 ( .A(n2682), .B(n2681), .Z(n2686) );
  NANDN U2846 ( .A(n2684), .B(n2683), .Z(n2685) );
  AND U2847 ( .A(n2686), .B(n2685), .Z(n3005) );
  XOR U2848 ( .A(n2687), .B(n3005), .Z(n3007) );
  NAND U2849 ( .A(n2689), .B(n2688), .Z(n2693) );
  NAND U2850 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U2851 ( .A(n2693), .B(n2692), .Z(n2982) );
  NAND U2852 ( .A(n2695), .B(n2694), .Z(n2699) );
  NAND U2853 ( .A(n2697), .B(n2696), .Z(n2698) );
  AND U2854 ( .A(n2699), .B(n2698), .Z(n2984) );
  NAND U2855 ( .A(n2701), .B(n2700), .Z(n2705) );
  NAND U2856 ( .A(n2703), .B(n2702), .Z(n2704) );
  AND U2857 ( .A(n2705), .B(n2704), .Z(n2983) );
  XOR U2858 ( .A(n2984), .B(n2983), .Z(n2981) );
  XOR U2859 ( .A(n2982), .B(n2981), .Z(n2999) );
  XOR U2860 ( .A(n3000), .B(n2999), .Z(n3001) );
  XOR U2861 ( .A(n3002), .B(n3001), .Z(n2716) );
  NAND U2862 ( .A(n2710), .B(n2709), .Z(n2714) );
  NANDN U2863 ( .A(n2712), .B(n2711), .Z(n2713) );
  NAND U2864 ( .A(n2714), .B(n2713), .Z(n2718) );
  XNOR U2865 ( .A(n2716), .B(n2715), .Z(N63) );
  NAND U2866 ( .A(n2716), .B(n2715), .Z(n2720) );
  NANDN U2867 ( .A(n2718), .B(n2717), .Z(n2719) );
  AND U2868 ( .A(n2720), .B(n2719), .Z(n2998) );
  NAND U2869 ( .A(n2722), .B(n2721), .Z(n2726) );
  NANDN U2870 ( .A(n2724), .B(n2723), .Z(n2725) );
  AND U2871 ( .A(n2726), .B(n2725), .Z(n2980) );
  NAND U2872 ( .A(n2728), .B(n2727), .Z(n2732) );
  NAND U2873 ( .A(n2730), .B(n2729), .Z(n2731) );
  AND U2874 ( .A(n2732), .B(n2731), .Z(n2740) );
  NANDN U2875 ( .A(n2734), .B(n2733), .Z(n2738) );
  NAND U2876 ( .A(n2736), .B(n2735), .Z(n2737) );
  NAND U2877 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U2878 ( .A(n2740), .B(n2739), .Z(n2978) );
  NAND U2879 ( .A(n2742), .B(n2741), .Z(n2746) );
  NAND U2880 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U2881 ( .A(n2746), .B(n2745), .Z(n2976) );
  NAND U2882 ( .A(n2748), .B(n2747), .Z(n2752) );
  NANDN U2883 ( .A(n2750), .B(n2749), .Z(n2751) );
  AND U2884 ( .A(n2752), .B(n2751), .Z(n2958) );
  NAND U2885 ( .A(n2754), .B(n2753), .Z(n2758) );
  NAND U2886 ( .A(n2756), .B(n2755), .Z(n2757) );
  AND U2887 ( .A(n2758), .B(n2757), .Z(n2766) );
  NANDN U2888 ( .A(n2760), .B(n2759), .Z(n2764) );
  NANDN U2889 ( .A(n2762), .B(n2761), .Z(n2763) );
  NAND U2890 ( .A(n2764), .B(n2763), .Z(n2765) );
  XNOR U2891 ( .A(n2766), .B(n2765), .Z(n2956) );
  NAND U2892 ( .A(n2768), .B(n2767), .Z(n2772) );
  NANDN U2893 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U2894 ( .A(n2772), .B(n2771), .Z(n2954) );
  NANDN U2895 ( .A(n2774), .B(n2773), .Z(n2778) );
  NANDN U2896 ( .A(n2776), .B(n2775), .Z(n2777) );
  AND U2897 ( .A(n2778), .B(n2777), .Z(n2786) );
  NANDN U2898 ( .A(n2780), .B(n2779), .Z(n2784) );
  NANDN U2899 ( .A(n2782), .B(n2781), .Z(n2783) );
  NAND U2900 ( .A(n2784), .B(n2783), .Z(n2785) );
  XNOR U2901 ( .A(n2786), .B(n2785), .Z(n2952) );
  NAND U2902 ( .A(n2788), .B(n2787), .Z(n2792) );
  NAND U2903 ( .A(n2790), .B(n2789), .Z(n2791) );
  AND U2904 ( .A(n2792), .B(n2791), .Z(n2950) );
  NAND U2905 ( .A(n2794), .B(n2793), .Z(n2797) );
  AND U2906 ( .A(y[21]), .B(x[10]), .Z(n2866) );
  NANDN U2907 ( .A(n2795), .B(n2866), .Z(n2796) );
  AND U2908 ( .A(n2797), .B(n2796), .Z(n2805) );
  NAND U2909 ( .A(n2799), .B(n2798), .Z(n2803) );
  NAND U2910 ( .A(n2801), .B(n2800), .Z(n2802) );
  NAND U2911 ( .A(n2803), .B(n2802), .Z(n2804) );
  XNOR U2912 ( .A(n2805), .B(n2804), .Z(n2948) );
  NAND U2913 ( .A(n2807), .B(n2806), .Z(n2810) );
  AND U2914 ( .A(y[27]), .B(x[4]), .Z(n2877) );
  NAND U2915 ( .A(n2808), .B(n2877), .Z(n2809) );
  AND U2916 ( .A(n2810), .B(n2809), .Z(n2840) );
  NAND U2917 ( .A(n2812), .B(n2811), .Z(n2815) );
  AND U2918 ( .A(x[6]), .B(y[25]), .Z(n2867) );
  NAND U2919 ( .A(n2813), .B(n2867), .Z(n2814) );
  AND U2920 ( .A(n2815), .B(n2814), .Z(n2822) );
  NAND U2921 ( .A(n2817), .B(n2816), .Z(n2820) );
  NAND U2922 ( .A(n2818), .B(n2878), .Z(n2819) );
  NAND U2923 ( .A(n2820), .B(n2819), .Z(n2821) );
  XNOR U2924 ( .A(n2822), .B(n2821), .Z(n2838) );
  AND U2925 ( .A(x[18]), .B(y[13]), .Z(n2824) );
  NAND U2926 ( .A(x[5]), .B(y[26]), .Z(n2823) );
  XNOR U2927 ( .A(n2824), .B(n2823), .Z(n2828) );
  AND U2928 ( .A(y[24]), .B(x[7]), .Z(n2826) );
  NAND U2929 ( .A(x[26]), .B(y[5]), .Z(n2825) );
  XNOR U2930 ( .A(n2826), .B(n2825), .Z(n2827) );
  XOR U2931 ( .A(n2828), .B(n2827), .Z(n2836) );
  AND U2932 ( .A(x[31]), .B(y[0]), .Z(n2830) );
  NAND U2933 ( .A(y[28]), .B(x[3]), .Z(n2829) );
  XNOR U2934 ( .A(n2830), .B(n2829), .Z(n2834) );
  AND U2935 ( .A(y[29]), .B(x[2]), .Z(n2832) );
  NAND U2936 ( .A(y[14]), .B(x[17]), .Z(n2831) );
  XNOR U2937 ( .A(n2832), .B(n2831), .Z(n2833) );
  XNOR U2938 ( .A(n2834), .B(n2833), .Z(n2835) );
  XNOR U2939 ( .A(n2836), .B(n2835), .Z(n2837) );
  XNOR U2940 ( .A(n2838), .B(n2837), .Z(n2839) );
  XNOR U2941 ( .A(n2840), .B(n2839), .Z(n2914) );
  NAND U2942 ( .A(n2842), .B(n2841), .Z(n2846) );
  AND U2943 ( .A(n2844), .B(n2843), .Z(n2845) );
  ANDN U2944 ( .B(n2846), .A(n2845), .Z(n2912) );
  AND U2945 ( .A(y[17]), .B(x[14]), .Z(n2848) );
  NAND U2946 ( .A(x[25]), .B(y[6]), .Z(n2847) );
  XNOR U2947 ( .A(n2848), .B(n2847), .Z(n2864) );
  AND U2948 ( .A(y[19]), .B(x[12]), .Z(n2850) );
  NAND U2949 ( .A(y[20]), .B(x[11]), .Z(n2849) );
  XNOR U2950 ( .A(n2850), .B(n2849), .Z(n2854) );
  AND U2951 ( .A(y[2]), .B(x[29]), .Z(n2852) );
  NAND U2952 ( .A(x[30]), .B(y[1]), .Z(n2851) );
  XNOR U2953 ( .A(n2852), .B(n2851), .Z(n2853) );
  XOR U2954 ( .A(n2854), .B(n2853), .Z(n2862) );
  AND U2955 ( .A(y[15]), .B(x[16]), .Z(n2856) );
  NAND U2956 ( .A(y[11]), .B(x[20]), .Z(n2855) );
  XNOR U2957 ( .A(n2856), .B(n2855), .Z(n2860) );
  AND U2958 ( .A(x[1]), .B(y[30]), .Z(n2858) );
  NAND U2959 ( .A(y[31]), .B(x[0]), .Z(n2857) );
  XNOR U2960 ( .A(n2858), .B(n2857), .Z(n2859) );
  XNOR U2961 ( .A(n2860), .B(n2859), .Z(n2861) );
  XNOR U2962 ( .A(n2862), .B(n2861), .Z(n2863) );
  XOR U2963 ( .A(n2864), .B(n2863), .Z(n2875) );
  XOR U2964 ( .A(n2866), .B(n2865), .Z(n2869) );
  XNOR U2965 ( .A(n2867), .B(n2917), .Z(n2868) );
  XNOR U2966 ( .A(n2869), .B(n2868), .Z(n2873) );
  AND U2967 ( .A(x[28]), .B(y[3]), .Z(n2871) );
  NAND U2968 ( .A(x[9]), .B(y[22]), .Z(n2870) );
  XNOR U2969 ( .A(n2871), .B(n2870), .Z(n2872) );
  XNOR U2970 ( .A(n2873), .B(n2872), .Z(n2874) );
  XNOR U2971 ( .A(n2875), .B(n2874), .Z(n2910) );
  AND U2972 ( .A(x[19]), .B(y[12]), .Z(n2884) );
  AND U2973 ( .A(n2876), .B(o[30]), .Z(n2882) );
  XOR U2974 ( .A(n2877), .B(o[31]), .Z(n2880) );
  AND U2975 ( .A(y[9]), .B(x[22]), .Z(n2924) );
  XNOR U2976 ( .A(n2924), .B(n2878), .Z(n2879) );
  XNOR U2977 ( .A(n2880), .B(n2879), .Z(n2881) );
  XNOR U2978 ( .A(n2882), .B(n2881), .Z(n2883) );
  XNOR U2979 ( .A(n2884), .B(n2883), .Z(n2900) );
  NAND U2980 ( .A(n2886), .B(n2885), .Z(n2890) );
  NAND U2981 ( .A(n2888), .B(n2887), .Z(n2889) );
  AND U2982 ( .A(n2890), .B(n2889), .Z(n2898) );
  NAND U2983 ( .A(n2892), .B(n2891), .Z(n2896) );
  NAND U2984 ( .A(n2894), .B(n2893), .Z(n2895) );
  NAND U2985 ( .A(n2896), .B(n2895), .Z(n2897) );
  XNOR U2986 ( .A(n2898), .B(n2897), .Z(n2899) );
  XOR U2987 ( .A(n2900), .B(n2899), .Z(n2908) );
  AND U2988 ( .A(x[27]), .B(y[4]), .Z(n2902) );
  NAND U2989 ( .A(y[8]), .B(x[23]), .Z(n2901) );
  XNOR U2990 ( .A(n2902), .B(n2901), .Z(n2906) );
  AND U2991 ( .A(y[23]), .B(x[8]), .Z(n2904) );
  NAND U2992 ( .A(x[21]), .B(y[10]), .Z(n2903) );
  XNOR U2993 ( .A(n2904), .B(n2903), .Z(n2905) );
  XNOR U2994 ( .A(n2906), .B(n2905), .Z(n2907) );
  XNOR U2995 ( .A(n2908), .B(n2907), .Z(n2909) );
  XNOR U2996 ( .A(n2910), .B(n2909), .Z(n2911) );
  XNOR U2997 ( .A(n2912), .B(n2911), .Z(n2913) );
  XOR U2998 ( .A(n2914), .B(n2913), .Z(n2946) );
  NAND U2999 ( .A(n2916), .B(n2915), .Z(n2920) );
  NAND U3000 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3001 ( .A(n2920), .B(n2919), .Z(n2928) );
  NAND U3002 ( .A(n2922), .B(n2921), .Z(n2926) );
  NAND U3003 ( .A(n2924), .B(n2923), .Z(n2925) );
  NAND U3004 ( .A(n2926), .B(n2925), .Z(n2927) );
  XNOR U3005 ( .A(n2928), .B(n2927), .Z(n2944) );
  NAND U3006 ( .A(n2930), .B(n2929), .Z(n2934) );
  NAND U3007 ( .A(n2932), .B(n2931), .Z(n2933) );
  AND U3008 ( .A(n2934), .B(n2933), .Z(n2942) );
  NAND U3009 ( .A(n2936), .B(n2935), .Z(n2940) );
  NAND U3010 ( .A(n2938), .B(n2937), .Z(n2939) );
  NAND U3011 ( .A(n2940), .B(n2939), .Z(n2941) );
  XNOR U3012 ( .A(n2942), .B(n2941), .Z(n2943) );
  XNOR U3013 ( .A(n2944), .B(n2943), .Z(n2945) );
  XNOR U3014 ( .A(n2946), .B(n2945), .Z(n2947) );
  XNOR U3015 ( .A(n2948), .B(n2947), .Z(n2949) );
  XNOR U3016 ( .A(n2950), .B(n2949), .Z(n2951) );
  XNOR U3017 ( .A(n2952), .B(n2951), .Z(n2953) );
  XNOR U3018 ( .A(n2954), .B(n2953), .Z(n2955) );
  XNOR U3019 ( .A(n2956), .B(n2955), .Z(n2957) );
  XNOR U3020 ( .A(n2958), .B(n2957), .Z(n2974) );
  NANDN U3021 ( .A(n2960), .B(n2959), .Z(n2964) );
  NANDN U3022 ( .A(n2962), .B(n2961), .Z(n2963) );
  AND U3023 ( .A(n2964), .B(n2963), .Z(n2972) );
  NANDN U3024 ( .A(n2966), .B(n2965), .Z(n2970) );
  NAND U3025 ( .A(n2968), .B(n2967), .Z(n2969) );
  NAND U3026 ( .A(n2970), .B(n2969), .Z(n2971) );
  XNOR U3027 ( .A(n2972), .B(n2971), .Z(n2973) );
  XNOR U3028 ( .A(n2974), .B(n2973), .Z(n2975) );
  XNOR U3029 ( .A(n2976), .B(n2975), .Z(n2977) );
  XNOR U3030 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U3031 ( .A(n2980), .B(n2979), .Z(n2996) );
  NAND U3032 ( .A(n2982), .B(n2981), .Z(n2986) );
  NAND U3033 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U3034 ( .A(n2986), .B(n2985), .Z(n2994) );
  NAND U3035 ( .A(n2988), .B(n2987), .Z(n2992) );
  NANDN U3036 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U3037 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U3038 ( .A(n2994), .B(n2993), .Z(n2995) );
  XNOR U3039 ( .A(n2996), .B(n2995), .Z(n2997) );
  XNOR U3040 ( .A(n2998), .B(n2997), .Z(n3014) );
  AND U3041 ( .A(n3000), .B(n2999), .Z(n3004) );
  AND U3042 ( .A(n3002), .B(n3001), .Z(n3003) );
  NOR U3043 ( .A(n3004), .B(n3003), .Z(n3012) );
  NANDN U3044 ( .A(n3006), .B(n3005), .Z(n3010) );
  NANDN U3045 ( .A(n3008), .B(n3007), .Z(n3009) );
  AND U3046 ( .A(n3010), .B(n3009), .Z(n3011) );
  XNOR U3047 ( .A(n3012), .B(n3011), .Z(n3013) );
  XNOR U3048 ( .A(n3014), .B(n3013), .Z(N64) );
endmodule

