
module stackMachine_N64 ( clk, rst, x, opcode, o );
  input [63:0] x;
  input [2:0] opcode;
  output [63:0] o;
  input clk, rst;
  wire   \stack[7][63] , \stack[7][62] , \stack[7][61] , \stack[7][60] ,
         \stack[7][59] , \stack[7][58] , \stack[7][57] , \stack[7][56] ,
         \stack[7][55] , \stack[7][54] , \stack[7][53] , \stack[7][52] ,
         \stack[7][51] , \stack[7][50] , \stack[7][49] , \stack[7][48] ,
         \stack[7][47] , \stack[7][46] , \stack[7][45] , \stack[7][44] ,
         \stack[7][43] , \stack[7][42] , \stack[7][41] , \stack[7][40] ,
         \stack[7][39] , \stack[7][38] , \stack[7][37] , \stack[7][36] ,
         \stack[7][35] , \stack[7][34] , \stack[7][33] , \stack[7][32] ,
         \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][63] , \stack[6][62] , \stack[6][61] , \stack[6][60] ,
         \stack[6][59] , \stack[6][58] , \stack[6][57] , \stack[6][56] ,
         \stack[6][55] , \stack[6][54] , \stack[6][53] , \stack[6][52] ,
         \stack[6][51] , \stack[6][50] , \stack[6][49] , \stack[6][48] ,
         \stack[6][47] , \stack[6][46] , \stack[6][45] , \stack[6][44] ,
         \stack[6][43] , \stack[6][42] , \stack[6][41] , \stack[6][40] ,
         \stack[6][39] , \stack[6][38] , \stack[6][37] , \stack[6][36] ,
         \stack[6][35] , \stack[6][34] , \stack[6][33] , \stack[6][32] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][63] , \stack[5][62] , \stack[5][61] , \stack[5][60] ,
         \stack[5][59] , \stack[5][58] , \stack[5][57] , \stack[5][56] ,
         \stack[5][55] , \stack[5][54] , \stack[5][53] , \stack[5][52] ,
         \stack[5][51] , \stack[5][50] , \stack[5][49] , \stack[5][48] ,
         \stack[5][47] , \stack[5][46] , \stack[5][45] , \stack[5][44] ,
         \stack[5][43] , \stack[5][42] , \stack[5][41] , \stack[5][40] ,
         \stack[5][39] , \stack[5][38] , \stack[5][37] , \stack[5][36] ,
         \stack[5][35] , \stack[5][34] , \stack[5][33] , \stack[5][32] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][63] , \stack[4][62] , \stack[4][61] , \stack[4][60] ,
         \stack[4][59] , \stack[4][58] , \stack[4][57] , \stack[4][56] ,
         \stack[4][55] , \stack[4][54] , \stack[4][53] , \stack[4][52] ,
         \stack[4][51] , \stack[4][50] , \stack[4][49] , \stack[4][48] ,
         \stack[4][47] , \stack[4][46] , \stack[4][45] , \stack[4][44] ,
         \stack[4][43] , \stack[4][42] , \stack[4][41] , \stack[4][40] ,
         \stack[4][39] , \stack[4][38] , \stack[4][37] , \stack[4][36] ,
         \stack[4][35] , \stack[4][34] , \stack[4][33] , \stack[4][32] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][63] , \stack[3][62] , \stack[3][61] , \stack[3][60] ,
         \stack[3][59] , \stack[3][58] , \stack[3][57] , \stack[3][56] ,
         \stack[3][55] , \stack[3][54] , \stack[3][53] , \stack[3][52] ,
         \stack[3][51] , \stack[3][50] , \stack[3][49] , \stack[3][48] ,
         \stack[3][47] , \stack[3][46] , \stack[3][45] , \stack[3][44] ,
         \stack[3][43] , \stack[3][42] , \stack[3][41] , \stack[3][40] ,
         \stack[3][39] , \stack[3][38] , \stack[3][37] , \stack[3][36] ,
         \stack[3][35] , \stack[3][34] , \stack[3][33] , \stack[3][32] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][63] , \stack[2][62] , \stack[2][61] , \stack[2][60] ,
         \stack[2][59] , \stack[2][58] , \stack[2][57] , \stack[2][56] ,
         \stack[2][55] , \stack[2][54] , \stack[2][53] , \stack[2][52] ,
         \stack[2][51] , \stack[2][50] , \stack[2][49] , \stack[2][48] ,
         \stack[2][47] , \stack[2][46] , \stack[2][45] , \stack[2][44] ,
         \stack[2][43] , \stack[2][42] , \stack[2][41] , \stack[2][40] ,
         \stack[2][39] , \stack[2][38] , \stack[2][37] , \stack[2][36] ,
         \stack[2][35] , \stack[2][34] , \stack[2][33] , \stack[2][32] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][63] , \stack[1][62] , \stack[1][61] , \stack[1][60] ,
         \stack[1][59] , \stack[1][58] , \stack[1][57] , \stack[1][56] ,
         \stack[1][55] , \stack[1][54] , \stack[1][53] , \stack[1][52] ,
         \stack[1][51] , \stack[1][50] , \stack[1][49] , \stack[1][48] ,
         \stack[1][47] , \stack[1][46] , \stack[1][45] , \stack[1][44] ,
         \stack[1][43] , \stack[1][42] , \stack[1][41] , \stack[1][40] ,
         \stack[1][39] , \stack[1][38] , \stack[1][37] , \stack[1][36] ,
         \stack[1][35] , \stack[1][34] , \stack[1][33] , \stack[1][32] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \stack[0][63] , \stack[0][62] , \stack[0][61] , \stack[0][60] ,
         \stack[0][59] , \stack[0][58] , \stack[0][57] , \stack[0][56] ,
         \stack[0][55] , \stack[0][54] , \stack[0][53] , \stack[0][52] ,
         \stack[0][51] , \stack[0][50] , \stack[0][49] , \stack[0][48] ,
         \stack[0][47] , \stack[0][46] , \stack[0][45] , \stack[0][44] ,
         \stack[0][43] , \stack[0][42] , \stack[0][41] , \stack[0][40] ,
         \stack[0][39] , \stack[0][38] , \stack[0][37] , \stack[0][36] ,
         \stack[0][35] , \stack[0][34] , \stack[0][33] , \stack[0][32] ,
         \stack[0][31] , \stack[0][30] , \stack[0][29] , \stack[0][28] ,
         \stack[0][27] , \stack[0][26] , \stack[0][25] , \stack[0][24] ,
         \stack[0][23] , \stack[0][22] , \stack[0][21] , \stack[0][20] ,
         \stack[0][19] , \stack[0][18] , \stack[0][17] , \stack[0][16] ,
         \stack[0][15] , \stack[0][14] , \stack[0][13] , \stack[0][12] ,
         \stack[0][11] , \stack[0][10] , \stack[0][9] , \stack[0][8] ,
         \stack[0][7] , \stack[0][6] , \stack[0][5] , \stack[0][4] ,
         \stack[0][3] , \stack[0][2] , \stack[0][1] , \stack[0][0] , n3941,
         n3948, n3955, n3964, n3973, n3982, n3991, n4000, n4009, n4018, n4027,
         n4036, n4045, n4054, n4063, n4072, n4081, n4090, n4099, n4108, n4117,
         n4126, n4135, n4144, n4153, n4162, n4171, n4180, n4189, n4198, n4207,
         n4216, n4225, n4234, n4243, n4252, n4261, n4270, n4279, n4288, n4297,
         n4306, n4315, n4324, n4333, n4342, n4351, n4360, n4369, n4378, n4387,
         n4396, n4405, n4414, n4423, n4432, n4441, n4450, n4459, n4468, n4477,
         n4486, n4495, n4504, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855;

  DFF \stack_reg[0][0]  ( .D(n4963), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][0] ) );
  DFF \stack_reg[1][0]  ( .D(n4899), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][0] ) );
  DFF \stack_reg[0][63]  ( .D(n4900), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][63] ) );
  DFF \stack_reg[1][63]  ( .D(n4836), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][63] ) );
  DFF \stack_reg[0][1]  ( .D(n4962), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][1] ) );
  DFF \stack_reg[1][1]  ( .D(n4898), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][1] ) );
  DFF \stack_reg[2][1]  ( .D(n4834), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][1] ) );
  DFF \stack_reg[3][1]  ( .D(n4770), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][1] ) );
  DFF \stack_reg[4][1]  ( .D(n4706), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][1] ) );
  DFF \stack_reg[5][1]  ( .D(n4642), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][1] ) );
  DFF \stack_reg[6][1]  ( .D(n4578), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][1] ) );
  DFF \stack_reg[7][1]  ( .D(n4504), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][1] ) );
  DFF \stack_reg[0][2]  ( .D(n4961), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][2] ) );
  DFF \stack_reg[1][2]  ( .D(n4897), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][2] ) );
  DFF \stack_reg[2][2]  ( .D(n4833), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][2] ) );
  DFF \stack_reg[3][2]  ( .D(n4769), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][2] ) );
  DFF \stack_reg[4][2]  ( .D(n4705), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][2] ) );
  DFF \stack_reg[5][2]  ( .D(n4641), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][2] ) );
  DFF \stack_reg[6][2]  ( .D(n4577), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][2] ) );
  DFF \stack_reg[7][2]  ( .D(n4495), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][2] ) );
  DFF \stack_reg[0][3]  ( .D(n4960), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][3] ) );
  DFF \stack_reg[1][3]  ( .D(n4896), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][3] ) );
  DFF \stack_reg[2][3]  ( .D(n4832), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][3] ) );
  DFF \stack_reg[3][3]  ( .D(n4768), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][3] ) );
  DFF \stack_reg[4][3]  ( .D(n4704), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][3] ) );
  DFF \stack_reg[5][3]  ( .D(n4640), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][3] ) );
  DFF \stack_reg[6][3]  ( .D(n4576), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][3] ) );
  DFF \stack_reg[7][3]  ( .D(n4486), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][3] ) );
  DFF \stack_reg[0][4]  ( .D(n4959), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][4] ) );
  DFF \stack_reg[1][4]  ( .D(n4895), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][4] ) );
  DFF \stack_reg[2][4]  ( .D(n4831), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][4] ) );
  DFF \stack_reg[3][4]  ( .D(n4767), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][4] ) );
  DFF \stack_reg[4][4]  ( .D(n4703), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][4] ) );
  DFF \stack_reg[5][4]  ( .D(n4639), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][4] ) );
  DFF \stack_reg[6][4]  ( .D(n4575), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][4] ) );
  DFF \stack_reg[7][4]  ( .D(n4477), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][4] ) );
  DFF \stack_reg[0][5]  ( .D(n4958), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][5] ) );
  DFF \stack_reg[1][5]  ( .D(n4894), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][5] ) );
  DFF \stack_reg[2][5]  ( .D(n4830), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][5] ) );
  DFF \stack_reg[3][5]  ( .D(n4766), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][5] ) );
  DFF \stack_reg[4][5]  ( .D(n4702), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][5] ) );
  DFF \stack_reg[5][5]  ( .D(n4638), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][5] ) );
  DFF \stack_reg[6][5]  ( .D(n4574), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][5] ) );
  DFF \stack_reg[7][5]  ( .D(n4468), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][5] ) );
  DFF \stack_reg[0][6]  ( .D(n4957), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][6] ) );
  DFF \stack_reg[1][6]  ( .D(n4893), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][6] ) );
  DFF \stack_reg[2][6]  ( .D(n4829), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][6] ) );
  DFF \stack_reg[3][6]  ( .D(n4765), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][6] ) );
  DFF \stack_reg[4][6]  ( .D(n4701), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][6] ) );
  DFF \stack_reg[5][6]  ( .D(n4637), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][6] ) );
  DFF \stack_reg[6][6]  ( .D(n4573), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][6] ) );
  DFF \stack_reg[7][6]  ( .D(n4459), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][6] ) );
  DFF \stack_reg[0][7]  ( .D(n4956), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][7] ) );
  DFF \stack_reg[1][7]  ( .D(n4892), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][7] ) );
  DFF \stack_reg[2][7]  ( .D(n4828), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][7] ) );
  DFF \stack_reg[3][7]  ( .D(n4764), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][7] ) );
  DFF \stack_reg[4][7]  ( .D(n4700), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][7] ) );
  DFF \stack_reg[5][7]  ( .D(n4636), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][7] ) );
  DFF \stack_reg[6][7]  ( .D(n4572), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][7] ) );
  DFF \stack_reg[7][7]  ( .D(n4450), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][7] ) );
  DFF \stack_reg[0][8]  ( .D(n4955), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][8] ) );
  DFF \stack_reg[1][8]  ( .D(n4891), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][8] ) );
  DFF \stack_reg[2][8]  ( .D(n4827), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][8] ) );
  DFF \stack_reg[3][8]  ( .D(n4763), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][8] ) );
  DFF \stack_reg[4][8]  ( .D(n4699), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][8] ) );
  DFF \stack_reg[5][8]  ( .D(n4635), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][8] ) );
  DFF \stack_reg[6][8]  ( .D(n4571), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][8] ) );
  DFF \stack_reg[7][8]  ( .D(n4441), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][8] ) );
  DFF \stack_reg[0][9]  ( .D(n4954), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][9] ) );
  DFF \stack_reg[1][9]  ( .D(n4890), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][9] ) );
  DFF \stack_reg[2][9]  ( .D(n4826), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][9] ) );
  DFF \stack_reg[3][9]  ( .D(n4762), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][9] ) );
  DFF \stack_reg[4][9]  ( .D(n4698), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][9] ) );
  DFF \stack_reg[5][9]  ( .D(n4634), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][9] ) );
  DFF \stack_reg[6][9]  ( .D(n4570), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][9] ) );
  DFF \stack_reg[7][9]  ( .D(n4432), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][9] ) );
  DFF \stack_reg[0][10]  ( .D(n4953), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][10] ) );
  DFF \stack_reg[1][10]  ( .D(n4889), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][10] ) );
  DFF \stack_reg[2][10]  ( .D(n4825), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][10] ) );
  DFF \stack_reg[3][10]  ( .D(n4761), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][10] ) );
  DFF \stack_reg[4][10]  ( .D(n4697), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][10] ) );
  DFF \stack_reg[5][10]  ( .D(n4633), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][10] ) );
  DFF \stack_reg[6][10]  ( .D(n4569), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][10] ) );
  DFF \stack_reg[7][10]  ( .D(n4423), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][10] ) );
  DFF \stack_reg[0][11]  ( .D(n4952), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][11] ) );
  DFF \stack_reg[1][11]  ( .D(n4888), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][11] ) );
  DFF \stack_reg[2][11]  ( .D(n4824), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][11] ) );
  DFF \stack_reg[3][11]  ( .D(n4760), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][11] ) );
  DFF \stack_reg[4][11]  ( .D(n4696), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][11] ) );
  DFF \stack_reg[5][11]  ( .D(n4632), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][11] ) );
  DFF \stack_reg[6][11]  ( .D(n4568), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][11] ) );
  DFF \stack_reg[7][11]  ( .D(n4414), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][11] ) );
  DFF \stack_reg[0][12]  ( .D(n4951), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][12] ) );
  DFF \stack_reg[1][12]  ( .D(n4887), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][12] ) );
  DFF \stack_reg[2][12]  ( .D(n4823), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][12] ) );
  DFF \stack_reg[3][12]  ( .D(n4759), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][12] ) );
  DFF \stack_reg[4][12]  ( .D(n4695), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][12] ) );
  DFF \stack_reg[5][12]  ( .D(n4631), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][12] ) );
  DFF \stack_reg[6][12]  ( .D(n4567), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][12] ) );
  DFF \stack_reg[7][12]  ( .D(n4405), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][12] ) );
  DFF \stack_reg[0][13]  ( .D(n4950), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][13] ) );
  DFF \stack_reg[1][13]  ( .D(n4886), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][13] ) );
  DFF \stack_reg[2][13]  ( .D(n4822), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][13] ) );
  DFF \stack_reg[3][13]  ( .D(n4758), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][13] ) );
  DFF \stack_reg[4][13]  ( .D(n4694), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][13] ) );
  DFF \stack_reg[5][13]  ( .D(n4630), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][13] ) );
  DFF \stack_reg[6][13]  ( .D(n4566), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][13] ) );
  DFF \stack_reg[7][13]  ( .D(n4396), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][13] ) );
  DFF \stack_reg[0][14]  ( .D(n4949), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][14] ) );
  DFF \stack_reg[1][14]  ( .D(n4885), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][14] ) );
  DFF \stack_reg[2][14]  ( .D(n4821), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][14] ) );
  DFF \stack_reg[3][14]  ( .D(n4757), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][14] ) );
  DFF \stack_reg[4][14]  ( .D(n4693), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][14] ) );
  DFF \stack_reg[5][14]  ( .D(n4629), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][14] ) );
  DFF \stack_reg[6][14]  ( .D(n4565), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][14] ) );
  DFF \stack_reg[7][14]  ( .D(n4387), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][14] ) );
  DFF \stack_reg[0][15]  ( .D(n4948), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][15] ) );
  DFF \stack_reg[1][15]  ( .D(n4884), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][15] ) );
  DFF \stack_reg[2][15]  ( .D(n4820), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][15] ) );
  DFF \stack_reg[3][15]  ( .D(n4756), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][15] ) );
  DFF \stack_reg[4][15]  ( .D(n4692), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][15] ) );
  DFF \stack_reg[5][15]  ( .D(n4628), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][15] ) );
  DFF \stack_reg[6][15]  ( .D(n4564), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][15] ) );
  DFF \stack_reg[7][15]  ( .D(n4378), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][15] ) );
  DFF \stack_reg[0][16]  ( .D(n4947), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][16] ) );
  DFF \stack_reg[1][16]  ( .D(n4883), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][16] ) );
  DFF \stack_reg[2][16]  ( .D(n4819), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][16] ) );
  DFF \stack_reg[3][16]  ( .D(n4755), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][16] ) );
  DFF \stack_reg[4][16]  ( .D(n4691), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][16] ) );
  DFF \stack_reg[5][16]  ( .D(n4627), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][16] ) );
  DFF \stack_reg[6][16]  ( .D(n4563), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][16] ) );
  DFF \stack_reg[7][16]  ( .D(n4369), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][16] ) );
  DFF \stack_reg[0][17]  ( .D(n4946), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][17] ) );
  DFF \stack_reg[1][17]  ( .D(n4882), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][17] ) );
  DFF \stack_reg[2][17]  ( .D(n4818), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][17] ) );
  DFF \stack_reg[3][17]  ( .D(n4754), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][17] ) );
  DFF \stack_reg[4][17]  ( .D(n4690), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][17] ) );
  DFF \stack_reg[5][17]  ( .D(n4626), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][17] ) );
  DFF \stack_reg[6][17]  ( .D(n4562), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][17] ) );
  DFF \stack_reg[7][17]  ( .D(n4360), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][17] ) );
  DFF \stack_reg[0][18]  ( .D(n4945), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][18] ) );
  DFF \stack_reg[1][18]  ( .D(n4881), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][18] ) );
  DFF \stack_reg[2][18]  ( .D(n4817), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][18] ) );
  DFF \stack_reg[3][18]  ( .D(n4753), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][18] ) );
  DFF \stack_reg[4][18]  ( .D(n4689), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][18] ) );
  DFF \stack_reg[5][18]  ( .D(n4625), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][18] ) );
  DFF \stack_reg[6][18]  ( .D(n4561), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][18] ) );
  DFF \stack_reg[7][18]  ( .D(n4351), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][18] ) );
  DFF \stack_reg[0][19]  ( .D(n4944), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][19] ) );
  DFF \stack_reg[1][19]  ( .D(n4880), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][19] ) );
  DFF \stack_reg[2][19]  ( .D(n4816), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][19] ) );
  DFF \stack_reg[3][19]  ( .D(n4752), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][19] ) );
  DFF \stack_reg[4][19]  ( .D(n4688), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][19] ) );
  DFF \stack_reg[5][19]  ( .D(n4624), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][19] ) );
  DFF \stack_reg[6][19]  ( .D(n4560), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][19] ) );
  DFF \stack_reg[7][19]  ( .D(n4342), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][19] ) );
  DFF \stack_reg[0][20]  ( .D(n4943), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][20] ) );
  DFF \stack_reg[1][20]  ( .D(n4879), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][20] ) );
  DFF \stack_reg[2][20]  ( .D(n4815), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][20] ) );
  DFF \stack_reg[3][20]  ( .D(n4751), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][20] ) );
  DFF \stack_reg[4][20]  ( .D(n4687), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][20] ) );
  DFF \stack_reg[5][20]  ( .D(n4623), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][20] ) );
  DFF \stack_reg[6][20]  ( .D(n4559), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][20] ) );
  DFF \stack_reg[7][20]  ( .D(n4333), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][20] ) );
  DFF \stack_reg[0][21]  ( .D(n4942), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][21] ) );
  DFF \stack_reg[1][21]  ( .D(n4878), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][21] ) );
  DFF \stack_reg[2][21]  ( .D(n4814), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][21] ) );
  DFF \stack_reg[3][21]  ( .D(n4750), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][21] ) );
  DFF \stack_reg[4][21]  ( .D(n4686), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][21] ) );
  DFF \stack_reg[5][21]  ( .D(n4622), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][21] ) );
  DFF \stack_reg[6][21]  ( .D(n4558), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][21] ) );
  DFF \stack_reg[7][21]  ( .D(n4324), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][21] ) );
  DFF \stack_reg[0][22]  ( .D(n4941), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][22] ) );
  DFF \stack_reg[1][22]  ( .D(n4877), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][22] ) );
  DFF \stack_reg[2][22]  ( .D(n4813), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][22] ) );
  DFF \stack_reg[3][22]  ( .D(n4749), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][22] ) );
  DFF \stack_reg[4][22]  ( .D(n4685), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][22] ) );
  DFF \stack_reg[5][22]  ( .D(n4621), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][22] ) );
  DFF \stack_reg[6][22]  ( .D(n4557), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][22] ) );
  DFF \stack_reg[7][22]  ( .D(n4315), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][22] ) );
  DFF \stack_reg[0][23]  ( .D(n4940), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][23] ) );
  DFF \stack_reg[1][23]  ( .D(n4876), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][23] ) );
  DFF \stack_reg[2][23]  ( .D(n4812), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][23] ) );
  DFF \stack_reg[3][23]  ( .D(n4748), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][23] ) );
  DFF \stack_reg[4][23]  ( .D(n4684), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][23] ) );
  DFF \stack_reg[5][23]  ( .D(n4620), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][23] ) );
  DFF \stack_reg[6][23]  ( .D(n4556), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][23] ) );
  DFF \stack_reg[7][23]  ( .D(n4306), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][23] ) );
  DFF \stack_reg[0][24]  ( .D(n4939), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][24] ) );
  DFF \stack_reg[1][24]  ( .D(n4875), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][24] ) );
  DFF \stack_reg[2][24]  ( .D(n4811), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][24] ) );
  DFF \stack_reg[3][24]  ( .D(n4747), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][24] ) );
  DFF \stack_reg[4][24]  ( .D(n4683), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][24] ) );
  DFF \stack_reg[5][24]  ( .D(n4619), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][24] ) );
  DFF \stack_reg[6][24]  ( .D(n4555), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][24] ) );
  DFF \stack_reg[7][24]  ( .D(n4297), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][24] ) );
  DFF \stack_reg[0][25]  ( .D(n4938), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][25] ) );
  DFF \stack_reg[1][25]  ( .D(n4874), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][25] ) );
  DFF \stack_reg[2][25]  ( .D(n4810), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][25] ) );
  DFF \stack_reg[3][25]  ( .D(n4746), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][25] ) );
  DFF \stack_reg[4][25]  ( .D(n4682), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][25] ) );
  DFF \stack_reg[5][25]  ( .D(n4618), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][25] ) );
  DFF \stack_reg[6][25]  ( .D(n4554), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][25] ) );
  DFF \stack_reg[7][25]  ( .D(n4288), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][25] ) );
  DFF \stack_reg[0][26]  ( .D(n4937), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][26] ) );
  DFF \stack_reg[1][26]  ( .D(n4873), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][26] ) );
  DFF \stack_reg[2][26]  ( .D(n4809), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][26] ) );
  DFF \stack_reg[3][26]  ( .D(n4745), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][26] ) );
  DFF \stack_reg[4][26]  ( .D(n4681), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][26] ) );
  DFF \stack_reg[5][26]  ( .D(n4617), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][26] ) );
  DFF \stack_reg[6][26]  ( .D(n4553), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][26] ) );
  DFF \stack_reg[7][26]  ( .D(n4279), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][26] ) );
  DFF \stack_reg[0][27]  ( .D(n4936), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][27] ) );
  DFF \stack_reg[1][27]  ( .D(n4872), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][27] ) );
  DFF \stack_reg[2][27]  ( .D(n4808), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][27] ) );
  DFF \stack_reg[3][27]  ( .D(n4744), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][27] ) );
  DFF \stack_reg[4][27]  ( .D(n4680), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][27] ) );
  DFF \stack_reg[5][27]  ( .D(n4616), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][27] ) );
  DFF \stack_reg[6][27]  ( .D(n4552), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][27] ) );
  DFF \stack_reg[7][27]  ( .D(n4270), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][27] ) );
  DFF \stack_reg[0][28]  ( .D(n4935), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][28] ) );
  DFF \stack_reg[1][28]  ( .D(n4871), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][28] ) );
  DFF \stack_reg[2][28]  ( .D(n4807), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][28] ) );
  DFF \stack_reg[3][28]  ( .D(n4743), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][28] ) );
  DFF \stack_reg[4][28]  ( .D(n4679), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][28] ) );
  DFF \stack_reg[5][28]  ( .D(n4615), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][28] ) );
  DFF \stack_reg[6][28]  ( .D(n4551), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][28] ) );
  DFF \stack_reg[7][28]  ( .D(n4261), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][28] ) );
  DFF \stack_reg[0][29]  ( .D(n4934), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][29] ) );
  DFF \stack_reg[1][29]  ( .D(n4870), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][29] ) );
  DFF \stack_reg[2][29]  ( .D(n4806), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][29] ) );
  DFF \stack_reg[3][29]  ( .D(n4742), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][29] ) );
  DFF \stack_reg[4][29]  ( .D(n4678), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][29] ) );
  DFF \stack_reg[5][29]  ( .D(n4614), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][29] ) );
  DFF \stack_reg[6][29]  ( .D(n4550), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][29] ) );
  DFF \stack_reg[7][29]  ( .D(n4252), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][29] ) );
  DFF \stack_reg[0][30]  ( .D(n4933), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][30] ) );
  DFF \stack_reg[1][30]  ( .D(n4869), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][30] ) );
  DFF \stack_reg[2][30]  ( .D(n4805), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][30] ) );
  DFF \stack_reg[3][30]  ( .D(n4741), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][30] ) );
  DFF \stack_reg[4][30]  ( .D(n4677), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][30] ) );
  DFF \stack_reg[5][30]  ( .D(n4613), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][30] ) );
  DFF \stack_reg[6][30]  ( .D(n4549), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][30] ) );
  DFF \stack_reg[7][30]  ( .D(n4243), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][30] ) );
  DFF \stack_reg[0][31]  ( .D(n4932), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][31] ) );
  DFF \stack_reg[1][31]  ( .D(n4868), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][31] ) );
  DFF \stack_reg[2][31]  ( .D(n4804), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][31] ) );
  DFF \stack_reg[3][31]  ( .D(n4740), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][31] ) );
  DFF \stack_reg[4][31]  ( .D(n4676), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][31] ) );
  DFF \stack_reg[5][31]  ( .D(n4612), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][31] ) );
  DFF \stack_reg[6][31]  ( .D(n4548), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][31] ) );
  DFF \stack_reg[7][31]  ( .D(n4234), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][31] ) );
  DFF \stack_reg[0][32]  ( .D(n4931), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][32] ) );
  DFF \stack_reg[1][32]  ( .D(n4867), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][32] ) );
  DFF \stack_reg[2][32]  ( .D(n4803), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][32] ) );
  DFF \stack_reg[3][32]  ( .D(n4739), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][32] ) );
  DFF \stack_reg[4][32]  ( .D(n4675), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][32] ) );
  DFF \stack_reg[5][32]  ( .D(n4611), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][32] ) );
  DFF \stack_reg[6][32]  ( .D(n4547), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][32] ) );
  DFF \stack_reg[7][32]  ( .D(n4225), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][32] ) );
  DFF \stack_reg[0][33]  ( .D(n4930), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][33] ) );
  DFF \stack_reg[1][33]  ( .D(n4866), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][33] ) );
  DFF \stack_reg[2][33]  ( .D(n4802), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][33] ) );
  DFF \stack_reg[3][33]  ( .D(n4738), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][33] ) );
  DFF \stack_reg[4][33]  ( .D(n4674), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][33] ) );
  DFF \stack_reg[5][33]  ( .D(n4610), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][33] ) );
  DFF \stack_reg[6][33]  ( .D(n4546), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][33] ) );
  DFF \stack_reg[7][33]  ( .D(n4216), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][33] ) );
  DFF \stack_reg[0][34]  ( .D(n4929), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][34] ) );
  DFF \stack_reg[1][34]  ( .D(n4865), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][34] ) );
  DFF \stack_reg[2][34]  ( .D(n4801), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][34] ) );
  DFF \stack_reg[3][34]  ( .D(n4737), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][34] ) );
  DFF \stack_reg[4][34]  ( .D(n4673), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][34] ) );
  DFF \stack_reg[5][34]  ( .D(n4609), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][34] ) );
  DFF \stack_reg[6][34]  ( .D(n4545), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][34] ) );
  DFF \stack_reg[7][34]  ( .D(n4207), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][34] ) );
  DFF \stack_reg[0][35]  ( .D(n4928), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][35] ) );
  DFF \stack_reg[1][35]  ( .D(n4864), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][35] ) );
  DFF \stack_reg[2][35]  ( .D(n4800), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][35] ) );
  DFF \stack_reg[3][35]  ( .D(n4736), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][35] ) );
  DFF \stack_reg[4][35]  ( .D(n4672), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][35] ) );
  DFF \stack_reg[5][35]  ( .D(n4608), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][35] ) );
  DFF \stack_reg[6][35]  ( .D(n4544), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][35] ) );
  DFF \stack_reg[7][35]  ( .D(n4198), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][35] ) );
  DFF \stack_reg[0][36]  ( .D(n4927), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][36] ) );
  DFF \stack_reg[1][36]  ( .D(n4863), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][36] ) );
  DFF \stack_reg[2][36]  ( .D(n4799), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][36] ) );
  DFF \stack_reg[3][36]  ( .D(n4735), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][36] ) );
  DFF \stack_reg[4][36]  ( .D(n4671), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][36] ) );
  DFF \stack_reg[5][36]  ( .D(n4607), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][36] ) );
  DFF \stack_reg[6][36]  ( .D(n4543), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][36] ) );
  DFF \stack_reg[7][36]  ( .D(n4189), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][36] ) );
  DFF \stack_reg[0][37]  ( .D(n4926), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][37] ) );
  DFF \stack_reg[1][37]  ( .D(n4862), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][37] ) );
  DFF \stack_reg[2][37]  ( .D(n4798), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][37] ) );
  DFF \stack_reg[3][37]  ( .D(n4734), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][37] ) );
  DFF \stack_reg[4][37]  ( .D(n4670), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][37] ) );
  DFF \stack_reg[5][37]  ( .D(n4606), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][37] ) );
  DFF \stack_reg[6][37]  ( .D(n4542), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][37] ) );
  DFF \stack_reg[7][37]  ( .D(n4180), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][37] ) );
  DFF \stack_reg[0][38]  ( .D(n4925), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][38] ) );
  DFF \stack_reg[1][38]  ( .D(n4861), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][38] ) );
  DFF \stack_reg[2][38]  ( .D(n4797), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][38] ) );
  DFF \stack_reg[3][38]  ( .D(n4733), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][38] ) );
  DFF \stack_reg[4][38]  ( .D(n4669), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][38] ) );
  DFF \stack_reg[5][38]  ( .D(n4605), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][38] ) );
  DFF \stack_reg[6][38]  ( .D(n4541), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][38] ) );
  DFF \stack_reg[7][38]  ( .D(n4171), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][38] ) );
  DFF \stack_reg[0][39]  ( .D(n4924), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][39] ) );
  DFF \stack_reg[1][39]  ( .D(n4860), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][39] ) );
  DFF \stack_reg[2][39]  ( .D(n4796), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][39] ) );
  DFF \stack_reg[3][39]  ( .D(n4732), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][39] ) );
  DFF \stack_reg[4][39]  ( .D(n4668), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][39] ) );
  DFF \stack_reg[5][39]  ( .D(n4604), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][39] ) );
  DFF \stack_reg[6][39]  ( .D(n4540), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][39] ) );
  DFF \stack_reg[7][39]  ( .D(n4162), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][39] ) );
  DFF \stack_reg[0][40]  ( .D(n4923), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][40] ) );
  DFF \stack_reg[1][40]  ( .D(n4859), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][40] ) );
  DFF \stack_reg[2][40]  ( .D(n4795), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][40] ) );
  DFF \stack_reg[3][40]  ( .D(n4731), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][40] ) );
  DFF \stack_reg[4][40]  ( .D(n4667), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][40] ) );
  DFF \stack_reg[5][40]  ( .D(n4603), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][40] ) );
  DFF \stack_reg[6][40]  ( .D(n4539), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][40] ) );
  DFF \stack_reg[7][40]  ( .D(n4153), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][40] ) );
  DFF \stack_reg[0][41]  ( .D(n4922), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][41] ) );
  DFF \stack_reg[1][41]  ( .D(n4858), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][41] ) );
  DFF \stack_reg[2][41]  ( .D(n4794), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][41] ) );
  DFF \stack_reg[3][41]  ( .D(n4730), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][41] ) );
  DFF \stack_reg[4][41]  ( .D(n4666), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][41] ) );
  DFF \stack_reg[5][41]  ( .D(n4602), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][41] ) );
  DFF \stack_reg[6][41]  ( .D(n4538), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][41] ) );
  DFF \stack_reg[7][41]  ( .D(n4144), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][41] ) );
  DFF \stack_reg[0][42]  ( .D(n4921), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][42] ) );
  DFF \stack_reg[1][42]  ( .D(n4857), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][42] ) );
  DFF \stack_reg[2][42]  ( .D(n4793), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][42] ) );
  DFF \stack_reg[3][42]  ( .D(n4729), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][42] ) );
  DFF \stack_reg[4][42]  ( .D(n4665), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][42] ) );
  DFF \stack_reg[5][42]  ( .D(n4601), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][42] ) );
  DFF \stack_reg[6][42]  ( .D(n4537), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][42] ) );
  DFF \stack_reg[7][42]  ( .D(n4135), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][42] ) );
  DFF \stack_reg[0][43]  ( .D(n4920), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][43] ) );
  DFF \stack_reg[1][43]  ( .D(n4856), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][43] ) );
  DFF \stack_reg[2][43]  ( .D(n4792), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][43] ) );
  DFF \stack_reg[3][43]  ( .D(n4728), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][43] ) );
  DFF \stack_reg[4][43]  ( .D(n4664), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][43] ) );
  DFF \stack_reg[5][43]  ( .D(n4600), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][43] ) );
  DFF \stack_reg[6][43]  ( .D(n4536), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][43] ) );
  DFF \stack_reg[7][43]  ( .D(n4126), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][43] ) );
  DFF \stack_reg[0][44]  ( .D(n4919), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][44] ) );
  DFF \stack_reg[1][44]  ( .D(n4855), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][44] ) );
  DFF \stack_reg[2][44]  ( .D(n4791), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][44] ) );
  DFF \stack_reg[3][44]  ( .D(n4727), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][44] ) );
  DFF \stack_reg[4][44]  ( .D(n4663), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][44] ) );
  DFF \stack_reg[5][44]  ( .D(n4599), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][44] ) );
  DFF \stack_reg[6][44]  ( .D(n4535), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][44] ) );
  DFF \stack_reg[7][44]  ( .D(n4117), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][44] ) );
  DFF \stack_reg[0][45]  ( .D(n4918), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][45] ) );
  DFF \stack_reg[1][45]  ( .D(n4854), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][45] ) );
  DFF \stack_reg[2][45]  ( .D(n4790), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][45] ) );
  DFF \stack_reg[3][45]  ( .D(n4726), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][45] ) );
  DFF \stack_reg[4][45]  ( .D(n4662), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][45] ) );
  DFF \stack_reg[5][45]  ( .D(n4598), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][45] ) );
  DFF \stack_reg[6][45]  ( .D(n4534), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][45] ) );
  DFF \stack_reg[7][45]  ( .D(n4108), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][45] ) );
  DFF \stack_reg[0][46]  ( .D(n4917), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][46] ) );
  DFF \stack_reg[1][46]  ( .D(n4853), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][46] ) );
  DFF \stack_reg[2][46]  ( .D(n4789), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][46] ) );
  DFF \stack_reg[3][46]  ( .D(n4725), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][46] ) );
  DFF \stack_reg[4][46]  ( .D(n4661), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][46] ) );
  DFF \stack_reg[5][46]  ( .D(n4597), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][46] ) );
  DFF \stack_reg[6][46]  ( .D(n4533), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][46] ) );
  DFF \stack_reg[7][46]  ( .D(n4099), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][46] ) );
  DFF \stack_reg[0][47]  ( .D(n4916), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][47] ) );
  DFF \stack_reg[1][47]  ( .D(n4852), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][47] ) );
  DFF \stack_reg[2][47]  ( .D(n4788), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][47] ) );
  DFF \stack_reg[3][47]  ( .D(n4724), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][47] ) );
  DFF \stack_reg[4][47]  ( .D(n4660), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][47] ) );
  DFF \stack_reg[5][47]  ( .D(n4596), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][47] ) );
  DFF \stack_reg[6][47]  ( .D(n4532), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][47] ) );
  DFF \stack_reg[7][47]  ( .D(n4090), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][47] ) );
  DFF \stack_reg[0][48]  ( .D(n4915), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][48] ) );
  DFF \stack_reg[1][48]  ( .D(n4851), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][48] ) );
  DFF \stack_reg[2][48]  ( .D(n4787), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][48] ) );
  DFF \stack_reg[3][48]  ( .D(n4723), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][48] ) );
  DFF \stack_reg[4][48]  ( .D(n4659), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][48] ) );
  DFF \stack_reg[5][48]  ( .D(n4595), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][48] ) );
  DFF \stack_reg[6][48]  ( .D(n4531), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][48] ) );
  DFF \stack_reg[7][48]  ( .D(n4081), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][48] ) );
  DFF \stack_reg[0][49]  ( .D(n4914), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][49] ) );
  DFF \stack_reg[1][49]  ( .D(n4850), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][49] ) );
  DFF \stack_reg[2][49]  ( .D(n4786), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][49] ) );
  DFF \stack_reg[3][49]  ( .D(n4722), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][49] ) );
  DFF \stack_reg[4][49]  ( .D(n4658), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][49] ) );
  DFF \stack_reg[5][49]  ( .D(n4594), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][49] ) );
  DFF \stack_reg[6][49]  ( .D(n4530), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][49] ) );
  DFF \stack_reg[7][49]  ( .D(n4072), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][49] ) );
  DFF \stack_reg[0][50]  ( .D(n4913), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][50] ) );
  DFF \stack_reg[1][50]  ( .D(n4849), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][50] ) );
  DFF \stack_reg[2][50]  ( .D(n4785), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][50] ) );
  DFF \stack_reg[3][50]  ( .D(n4721), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][50] ) );
  DFF \stack_reg[4][50]  ( .D(n4657), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][50] ) );
  DFF \stack_reg[5][50]  ( .D(n4593), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][50] ) );
  DFF \stack_reg[6][50]  ( .D(n4529), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][50] ) );
  DFF \stack_reg[7][50]  ( .D(n4063), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][50] ) );
  DFF \stack_reg[0][51]  ( .D(n4912), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][51] ) );
  DFF \stack_reg[1][51]  ( .D(n4848), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][51] ) );
  DFF \stack_reg[2][51]  ( .D(n4784), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][51] ) );
  DFF \stack_reg[3][51]  ( .D(n4720), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][51] ) );
  DFF \stack_reg[4][51]  ( .D(n4656), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][51] ) );
  DFF \stack_reg[5][51]  ( .D(n4592), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][51] ) );
  DFF \stack_reg[6][51]  ( .D(n4528), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][51] ) );
  DFF \stack_reg[7][51]  ( .D(n4054), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][51] ) );
  DFF \stack_reg[0][52]  ( .D(n4911), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][52] ) );
  DFF \stack_reg[1][52]  ( .D(n4847), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][52] ) );
  DFF \stack_reg[2][52]  ( .D(n4783), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][52] ) );
  DFF \stack_reg[3][52]  ( .D(n4719), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][52] ) );
  DFF \stack_reg[4][52]  ( .D(n4655), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][52] ) );
  DFF \stack_reg[5][52]  ( .D(n4591), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][52] ) );
  DFF \stack_reg[6][52]  ( .D(n4527), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][52] ) );
  DFF \stack_reg[7][52]  ( .D(n4045), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][52] ) );
  DFF \stack_reg[0][53]  ( .D(n4910), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][53] ) );
  DFF \stack_reg[1][53]  ( .D(n4846), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][53] ) );
  DFF \stack_reg[2][53]  ( .D(n4782), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][53] ) );
  DFF \stack_reg[3][53]  ( .D(n4718), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][53] ) );
  DFF \stack_reg[4][53]  ( .D(n4654), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][53] ) );
  DFF \stack_reg[5][53]  ( .D(n4590), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][53] ) );
  DFF \stack_reg[6][53]  ( .D(n4526), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][53] ) );
  DFF \stack_reg[7][53]  ( .D(n4036), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][53] ) );
  DFF \stack_reg[0][54]  ( .D(n4909), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][54] ) );
  DFF \stack_reg[1][54]  ( .D(n4845), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][54] ) );
  DFF \stack_reg[2][54]  ( .D(n4781), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][54] ) );
  DFF \stack_reg[3][54]  ( .D(n4717), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][54] ) );
  DFF \stack_reg[4][54]  ( .D(n4653), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][54] ) );
  DFF \stack_reg[5][54]  ( .D(n4589), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][54] ) );
  DFF \stack_reg[6][54]  ( .D(n4525), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][54] ) );
  DFF \stack_reg[7][54]  ( .D(n4027), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][54] ) );
  DFF \stack_reg[0][55]  ( .D(n4908), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][55] ) );
  DFF \stack_reg[1][55]  ( .D(n4844), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][55] ) );
  DFF \stack_reg[2][55]  ( .D(n4780), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][55] ) );
  DFF \stack_reg[3][55]  ( .D(n4716), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][55] ) );
  DFF \stack_reg[4][55]  ( .D(n4652), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][55] ) );
  DFF \stack_reg[5][55]  ( .D(n4588), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][55] ) );
  DFF \stack_reg[6][55]  ( .D(n4524), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][55] ) );
  DFF \stack_reg[7][55]  ( .D(n4018), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][55] ) );
  DFF \stack_reg[0][56]  ( .D(n4907), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][56] ) );
  DFF \stack_reg[1][56]  ( .D(n4843), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][56] ) );
  DFF \stack_reg[2][56]  ( .D(n4779), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][56] ) );
  DFF \stack_reg[3][56]  ( .D(n4715), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][56] ) );
  DFF \stack_reg[4][56]  ( .D(n4651), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][56] ) );
  DFF \stack_reg[5][56]  ( .D(n4587), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][56] ) );
  DFF \stack_reg[6][56]  ( .D(n4523), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][56] ) );
  DFF \stack_reg[7][56]  ( .D(n4009), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][56] ) );
  DFF \stack_reg[0][57]  ( .D(n4906), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][57] ) );
  DFF \stack_reg[1][57]  ( .D(n4842), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][57] ) );
  DFF \stack_reg[2][57]  ( .D(n4778), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][57] ) );
  DFF \stack_reg[3][57]  ( .D(n4714), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][57] ) );
  DFF \stack_reg[4][57]  ( .D(n4650), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][57] ) );
  DFF \stack_reg[5][57]  ( .D(n4586), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][57] ) );
  DFF \stack_reg[6][57]  ( .D(n4522), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][57] ) );
  DFF \stack_reg[7][57]  ( .D(n4000), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][57] ) );
  DFF \stack_reg[0][58]  ( .D(n4905), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][58] ) );
  DFF \stack_reg[1][58]  ( .D(n4841), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][58] ) );
  DFF \stack_reg[2][58]  ( .D(n4777), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][58] ) );
  DFF \stack_reg[3][58]  ( .D(n4713), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][58] ) );
  DFF \stack_reg[4][58]  ( .D(n4649), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][58] ) );
  DFF \stack_reg[5][58]  ( .D(n4585), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][58] ) );
  DFF \stack_reg[6][58]  ( .D(n4521), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][58] ) );
  DFF \stack_reg[7][58]  ( .D(n3991), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][58] ) );
  DFF \stack_reg[0][59]  ( .D(n4904), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][59] ) );
  DFF \stack_reg[1][59]  ( .D(n4840), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][59] ) );
  DFF \stack_reg[2][59]  ( .D(n4776), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][59] ) );
  DFF \stack_reg[3][59]  ( .D(n4712), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][59] ) );
  DFF \stack_reg[4][59]  ( .D(n4648), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][59] ) );
  DFF \stack_reg[5][59]  ( .D(n4584), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][59] ) );
  DFF \stack_reg[6][59]  ( .D(n4520), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][59] ) );
  DFF \stack_reg[7][59]  ( .D(n3982), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][59] ) );
  DFF \stack_reg[0][60]  ( .D(n4903), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][60] ) );
  DFF \stack_reg[1][60]  ( .D(n4839), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][60] ) );
  DFF \stack_reg[2][60]  ( .D(n4775), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][60] ) );
  DFF \stack_reg[3][60]  ( .D(n4711), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][60] ) );
  DFF \stack_reg[4][60]  ( .D(n4647), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][60] ) );
  DFF \stack_reg[5][60]  ( .D(n4583), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][60] ) );
  DFF \stack_reg[6][60]  ( .D(n4519), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][60] ) );
  DFF \stack_reg[7][60]  ( .D(n3973), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][60] ) );
  DFF \stack_reg[0][61]  ( .D(n4902), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][61] ) );
  DFF \stack_reg[1][61]  ( .D(n4838), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][61] ) );
  DFF \stack_reg[2][61]  ( .D(n4774), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][61] ) );
  DFF \stack_reg[3][61]  ( .D(n4710), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][61] ) );
  DFF \stack_reg[4][61]  ( .D(n4646), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][61] ) );
  DFF \stack_reg[5][61]  ( .D(n4582), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][61] ) );
  DFF \stack_reg[6][61]  ( .D(n4518), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][61] ) );
  DFF \stack_reg[7][61]  ( .D(n3964), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][61] ) );
  DFF \stack_reg[0][62]  ( .D(n4901), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][62] ) );
  DFF \stack_reg[1][62]  ( .D(n4837), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][62] ) );
  DFF \stack_reg[2][62]  ( .D(n4773), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][62] ) );
  DFF \stack_reg[3][62]  ( .D(n4709), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][62] ) );
  DFF \stack_reg[4][62]  ( .D(n4645), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][62] ) );
  DFF \stack_reg[5][62]  ( .D(n4581), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][62] ) );
  DFF \stack_reg[6][62]  ( .D(n4517), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][62] ) );
  DFF \stack_reg[7][62]  ( .D(n3955), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][62] ) );
  DFF \stack_reg[2][63]  ( .D(n4772), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][63] ) );
  DFF \stack_reg[3][63]  ( .D(n4708), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][63] ) );
  DFF \stack_reg[4][63]  ( .D(n4644), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][63] ) );
  DFF \stack_reg[5][63]  ( .D(n4580), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][63] ) );
  DFF \stack_reg[6][63]  ( .D(n4516), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][63] ) );
  DFF \stack_reg[7][63]  ( .D(n3948), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][63] ) );
  DFF \stack_reg[2][0]  ( .D(n4835), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][0] ) );
  DFF \stack_reg[3][0]  ( .D(n4771), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][0] ) );
  DFF \stack_reg[4][0]  ( .D(n4707), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][0] ) );
  DFF \stack_reg[5][0]  ( .D(n4643), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][0] ) );
  DFF \stack_reg[6][0]  ( .D(n4579), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][0] ) );
  DFF \stack_reg[7][0]  ( .D(n3941), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][0] ) );
  NAND U5024 ( .A(n15958), .B(n15957), .Z(n15953) );
  NANDN U5025 ( .A(n8997), .B(n8999), .Z(n11216) );
  NANDN U5026 ( .A(n9025), .B(n9027), .Z(n12575) );
  NANDN U5027 ( .A(n9053), .B(n9055), .Z(n13822) );
  NANDN U5028 ( .A(n7772), .B(n7774), .Z(n8571) );
  NAND U5029 ( .A(n15181), .B(n15180), .Z(n15176) );
  NAND U5030 ( .A(n14047), .B(n14046), .Z(n14042) );
  NAND U5031 ( .A(n12800), .B(n12799), .Z(n12795) );
  NAND U5032 ( .A(n11441), .B(n11440), .Z(n11436) );
  NAND U5033 ( .A(n9971), .B(n9970), .Z(n9966) );
  NANDN U5034 ( .A(n8930), .B(n8932), .Z(n9339) );
  NANDN U5035 ( .A(n8594), .B(n8596), .Z(n9002) );
  NANDN U5036 ( .A(n8622), .B(n8624), .Z(n9030) );
  NANDN U5037 ( .A(n8650), .B(n8652), .Z(n9058) );
  NANDN U5038 ( .A(n8566), .B(n8568), .Z(n8973) );
  NANDN U5039 ( .A(n7099), .B(n7101), .Z(n7763) );
  NANDN U5040 ( .A(n7083), .B(n7085), .Z(n7819) );
  NANDN U5041 ( .A(n7067), .B(n7069), .Z(n7875) );
  NANDN U5042 ( .A(n7051), .B(n7053), .Z(n7931) );
  NAND U5043 ( .A(n15965), .B(n15964), .Z(n15960) );
  NAND U5044 ( .A(n15447), .B(n15446), .Z(n15442) );
  NAND U5045 ( .A(n14628), .B(n14627), .Z(n14623) );
  NAND U5046 ( .A(n13438), .B(n13437), .Z(n13433) );
  NAND U5047 ( .A(n12135), .B(n12134), .Z(n12130) );
  NAND U5048 ( .A(n10720), .B(n10719), .Z(n10715) );
  XOR U5049 ( .A(n7501), .B(n9580), .Z(n7518) );
  NANDN U5050 ( .A(n8608), .B(n8610), .Z(n9016) );
  NANDN U5051 ( .A(n8636), .B(n8638), .Z(n9044) );
  NANDN U5052 ( .A(n8982), .B(n8984), .Z(n10495) );
  NANDN U5053 ( .A(n7744), .B(n7746), .Z(n8557) );
  NANDN U5054 ( .A(n8498), .B(n8499), .Z(n8497) );
  NANDN U5055 ( .A(n7091), .B(n7093), .Z(n7791) );
  NANDN U5056 ( .A(n7075), .B(n7077), .Z(n7847) );
  NANDN U5057 ( .A(n7059), .B(n7061), .Z(n7903) );
  NANDN U5058 ( .A(n7043), .B(n7045), .Z(n7959) );
  NAND U5059 ( .A(n16203), .B(n16202), .Z(n16198) );
  NAND U5060 ( .A(n15454), .B(n15453), .Z(n15449) );
  NAND U5061 ( .A(n14908), .B(n14907), .Z(n14903) );
  NAND U5062 ( .A(n14348), .B(n14347), .Z(n14343) );
  NAND U5063 ( .A(n13746), .B(n13745), .Z(n13741) );
  NAND U5064 ( .A(n13129), .B(n13128), .Z(n13124) );
  NAND U5065 ( .A(n12471), .B(n12470), .Z(n12466) );
  NAND U5066 ( .A(n11798), .B(n11797), .Z(n11793) );
  NAND U5067 ( .A(n11084), .B(n11083), .Z(n11079) );
  NAND U5068 ( .A(n10356), .B(n10355), .Z(n10351) );
  NAND U5069 ( .A(n9586), .B(n9585), .Z(n9581) );
  NANDN U5070 ( .A(n9067), .B(n9069), .Z(n14403) );
  NANDN U5071 ( .A(n9095), .B(n9097), .Z(n15481) );
  NANDN U5072 ( .A(n9123), .B(n9125), .Z(n16447) );
  NANDN U5073 ( .A(n9151), .B(n9153), .Z(n17301) );
  NANDN U5074 ( .A(n9179), .B(n9181), .Z(n18043) );
  NANDN U5075 ( .A(n9207), .B(n9209), .Z(n18673) );
  NANDN U5076 ( .A(n9235), .B(n9237), .Z(n19191) );
  NANDN U5077 ( .A(n9263), .B(n9265), .Z(n19597) );
  NANDN U5078 ( .A(n9291), .B(n9293), .Z(n19891) );
  NANDN U5079 ( .A(n9319), .B(n9321), .Z(n20073) );
  NANDN U5080 ( .A(n8664), .B(n8666), .Z(n9072) );
  NANDN U5081 ( .A(n8692), .B(n8694), .Z(n9100) );
  NANDN U5082 ( .A(n8720), .B(n8722), .Z(n9128) );
  NANDN U5083 ( .A(n8748), .B(n8750), .Z(n9156) );
  NANDN U5084 ( .A(n8776), .B(n8778), .Z(n9184) );
  NANDN U5085 ( .A(n8804), .B(n8806), .Z(n9212) );
  NANDN U5086 ( .A(n8832), .B(n8834), .Z(n9240) );
  NANDN U5087 ( .A(n8860), .B(n8862), .Z(n9268) );
  NANDN U5088 ( .A(n8888), .B(n8890), .Z(n9296) );
  NANDN U5089 ( .A(n8916), .B(n8918), .Z(n9324) );
  NANDN U5090 ( .A(n7800), .B(n7802), .Z(n8585) );
  NANDN U5091 ( .A(n7856), .B(n7858), .Z(n8613) );
  NANDN U5092 ( .A(n7912), .B(n7914), .Z(n8641) );
  NANDN U5093 ( .A(n7968), .B(n7970), .Z(n8669) );
  NANDN U5094 ( .A(n8024), .B(n8026), .Z(n8697) );
  NANDN U5095 ( .A(n8080), .B(n8082), .Z(n8725) );
  NANDN U5096 ( .A(n8136), .B(n8138), .Z(n8753) );
  NANDN U5097 ( .A(n8192), .B(n8194), .Z(n8781) );
  NANDN U5098 ( .A(n8248), .B(n8250), .Z(n8809) );
  NANDN U5099 ( .A(n8304), .B(n8306), .Z(n8837) );
  NANDN U5100 ( .A(n8360), .B(n8362), .Z(n8865) );
  NANDN U5101 ( .A(n8416), .B(n8418), .Z(n8893) );
  NANDN U5102 ( .A(n8502), .B(n8504), .Z(n8935) );
  NANDN U5103 ( .A(n8552), .B(n8554), .Z(n8959) );
  NANDN U5104 ( .A(n7027), .B(n7029), .Z(n8015) );
  NANDN U5105 ( .A(n7011), .B(n7013), .Z(n8071) );
  NANDN U5106 ( .A(n6995), .B(n6997), .Z(n8127) );
  NANDN U5107 ( .A(n6979), .B(n6981), .Z(n8183) );
  NANDN U5108 ( .A(n6963), .B(n6965), .Z(n8239) );
  NANDN U5109 ( .A(n6947), .B(n6949), .Z(n8295) );
  NANDN U5110 ( .A(n6931), .B(n6933), .Z(n8351) );
  NANDN U5111 ( .A(n6915), .B(n6917), .Z(n8407) );
  NANDN U5112 ( .A(n6903), .B(n6905), .Z(n8493) );
  NANDN U5113 ( .A(n6605), .B(n6607), .Z(n6697) );
  NANDN U5114 ( .A(n6509), .B(n6511), .Z(n6709) );
  NANDN U5115 ( .A(n6413), .B(n6415), .Z(n6721) );
  NANDN U5116 ( .A(n6317), .B(n6319), .Z(n6733) );
  NANDN U5117 ( .A(n6221), .B(n6223), .Z(n6745) );
  NANDN U5118 ( .A(n6125), .B(n6127), .Z(n6757) );
  NANDN U5119 ( .A(n6029), .B(n6031), .Z(n6769) );
  NANDN U5120 ( .A(n5933), .B(n5935), .Z(n6781) );
  NANDN U5121 ( .A(n5837), .B(n5839), .Z(n6793) );
  NANDN U5122 ( .A(n5741), .B(n5743), .Z(n6805) );
  NANDN U5123 ( .A(n5645), .B(n5647), .Z(n6817) );
  NANDN U5124 ( .A(n5549), .B(n5551), .Z(n6829) );
  NAND U5125 ( .A(n15706), .B(n15705), .Z(n15701) );
  NAND U5126 ( .A(n14915), .B(n14914), .Z(n14910) );
  NAND U5127 ( .A(n14341), .B(n14340), .Z(n14336) );
  NAND U5128 ( .A(n13753), .B(n13752), .Z(n13748) );
  NAND U5129 ( .A(n13122), .B(n13121), .Z(n13117) );
  NAND U5130 ( .A(n12478), .B(n12477), .Z(n12473) );
  NAND U5131 ( .A(n11791), .B(n11790), .Z(n11786) );
  NAND U5132 ( .A(n11091), .B(n11090), .Z(n11086) );
  NAND U5133 ( .A(n10349), .B(n10348), .Z(n10344) );
  NAND U5134 ( .A(n9593), .B(n9592), .Z(n9588) );
  NAND U5135 ( .A(n7504), .B(n7503), .Z(n7499) );
  NANDN U5136 ( .A(n9081), .B(n9083), .Z(n14956) );
  NANDN U5137 ( .A(n9109), .B(n9111), .Z(n15978) );
  NANDN U5138 ( .A(n9137), .B(n9139), .Z(n16888) );
  NANDN U5139 ( .A(n9165), .B(n9167), .Z(n17686) );
  NANDN U5140 ( .A(n9193), .B(n9195), .Z(n18372) );
  NANDN U5141 ( .A(n9221), .B(n9223), .Z(n18946) );
  NANDN U5142 ( .A(n9249), .B(n9251), .Z(n19408) );
  NANDN U5143 ( .A(n9277), .B(n9279), .Z(n19758) );
  NANDN U5144 ( .A(n9305), .B(n9307), .Z(n19996) );
  NANDN U5145 ( .A(n8678), .B(n8680), .Z(n9086) );
  NANDN U5146 ( .A(n8706), .B(n8708), .Z(n9114) );
  NANDN U5147 ( .A(n8734), .B(n8736), .Z(n9142) );
  NANDN U5148 ( .A(n8762), .B(n8764), .Z(n9170) );
  NANDN U5149 ( .A(n8790), .B(n8792), .Z(n9198) );
  NANDN U5150 ( .A(n8818), .B(n8820), .Z(n9226) );
  NANDN U5151 ( .A(n8846), .B(n8848), .Z(n9254) );
  NANDN U5152 ( .A(n8874), .B(n8876), .Z(n9282) );
  NANDN U5153 ( .A(n8902), .B(n8904), .Z(n9310) );
  NANDN U5154 ( .A(n7134), .B(n7133), .Z(n7136) );
  NANDN U5155 ( .A(n7828), .B(n7830), .Z(n8599) );
  NANDN U5156 ( .A(n7884), .B(n7886), .Z(n8627) );
  NANDN U5157 ( .A(n7940), .B(n7942), .Z(n8655) );
  NANDN U5158 ( .A(n7996), .B(n7998), .Z(n8683) );
  NANDN U5159 ( .A(n8052), .B(n8054), .Z(n8711) );
  NANDN U5160 ( .A(n8108), .B(n8110), .Z(n8739) );
  NANDN U5161 ( .A(n8164), .B(n8166), .Z(n8767) );
  NANDN U5162 ( .A(n8220), .B(n8222), .Z(n8795) );
  NANDN U5163 ( .A(n8276), .B(n8278), .Z(n8823) );
  NANDN U5164 ( .A(n8332), .B(n8334), .Z(n8851) );
  NANDN U5165 ( .A(n8388), .B(n8390), .Z(n8879) );
  NANDN U5166 ( .A(n8444), .B(n8446), .Z(n8907) );
  NANDN U5167 ( .A(n8470), .B(n8471), .Z(n8469) );
  NANDN U5168 ( .A(n8968), .B(n8970), .Z(n9746) );
  NANDN U5169 ( .A(n7107), .B(n7109), .Z(n7735) );
  NANDN U5170 ( .A(n7035), .B(n7037), .Z(n7987) );
  NANDN U5171 ( .A(n7019), .B(n7021), .Z(n8043) );
  NANDN U5172 ( .A(n7003), .B(n7005), .Z(n8099) );
  NANDN U5173 ( .A(n6987), .B(n6989), .Z(n8155) );
  NANDN U5174 ( .A(n6971), .B(n6973), .Z(n8211) );
  NANDN U5175 ( .A(n6955), .B(n6957), .Z(n8267) );
  NANDN U5176 ( .A(n6939), .B(n6941), .Z(n8323) );
  NANDN U5177 ( .A(n6923), .B(n6925), .Z(n8379) );
  NANDN U5178 ( .A(n6907), .B(n6909), .Z(n8435) );
  NANDN U5179 ( .A(n6899), .B(n6901), .Z(n8521) );
  NANDN U5180 ( .A(n6557), .B(n6559), .Z(n6703) );
  NANDN U5181 ( .A(n6461), .B(n6463), .Z(n6715) );
  NANDN U5182 ( .A(n6365), .B(n6367), .Z(n6727) );
  NANDN U5183 ( .A(n6269), .B(n6271), .Z(n6739) );
  NANDN U5184 ( .A(n6173), .B(n6175), .Z(n6751) );
  NANDN U5185 ( .A(n6077), .B(n6079), .Z(n6763) );
  NANDN U5186 ( .A(n5981), .B(n5983), .Z(n6775) );
  NANDN U5187 ( .A(n5885), .B(n5887), .Z(n6787) );
  NANDN U5188 ( .A(n5789), .B(n5791), .Z(n6799) );
  NANDN U5189 ( .A(n5693), .B(n5695), .Z(n6811) );
  NANDN U5190 ( .A(n5597), .B(n5599), .Z(n6823) );
  NANDN U5191 ( .A(n5501), .B(n5503), .Z(n6835) );
  NAND U5192 ( .A(n5392), .B(n5394), .Z(n20384) );
  XNOR U5193 ( .A(n5383), .B(n5384), .Z(n5382) );
  NANDN U5194 ( .A(n4964), .B(n4965), .Z(o[9]) );
  OR U5195 ( .A(n4966), .B(n4967), .Z(n4965) );
  NANDN U5196 ( .A(n4968), .B(n4969), .Z(o[8]) );
  OR U5197 ( .A(n4970), .B(n4967), .Z(n4969) );
  NANDN U5198 ( .A(n4971), .B(n4972), .Z(o[7]) );
  OR U5199 ( .A(n4973), .B(n4967), .Z(n4972) );
  NANDN U5200 ( .A(n4974), .B(n4975), .Z(o[6]) );
  OR U5201 ( .A(n4976), .B(n4967), .Z(n4975) );
  NANDN U5202 ( .A(n4977), .B(n4978), .Z(o[63]) );
  OR U5203 ( .A(n4979), .B(n4967), .Z(n4978) );
  NANDN U5204 ( .A(n4980), .B(n4981), .Z(o[62]) );
  OR U5205 ( .A(n4982), .B(n4967), .Z(n4981) );
  NANDN U5206 ( .A(n4983), .B(n4984), .Z(o[61]) );
  OR U5207 ( .A(n4985), .B(n4967), .Z(n4984) );
  NANDN U5208 ( .A(n4986), .B(n4987), .Z(o[60]) );
  OR U5209 ( .A(n4988), .B(n4967), .Z(n4987) );
  NANDN U5210 ( .A(n4989), .B(n4990), .Z(o[5]) );
  OR U5211 ( .A(n4991), .B(n4967), .Z(n4990) );
  NANDN U5212 ( .A(n4992), .B(n4993), .Z(o[59]) );
  OR U5213 ( .A(n4994), .B(n4967), .Z(n4993) );
  NANDN U5214 ( .A(n4995), .B(n4996), .Z(o[58]) );
  OR U5215 ( .A(n4997), .B(n4967), .Z(n4996) );
  NANDN U5216 ( .A(n4998), .B(n4999), .Z(o[57]) );
  OR U5217 ( .A(n5000), .B(n4967), .Z(n4999) );
  NANDN U5218 ( .A(n5001), .B(n5002), .Z(o[56]) );
  OR U5219 ( .A(n5003), .B(n4967), .Z(n5002) );
  NANDN U5220 ( .A(n5004), .B(n5005), .Z(o[55]) );
  OR U5221 ( .A(n5006), .B(n4967), .Z(n5005) );
  NANDN U5222 ( .A(n5007), .B(n5008), .Z(o[54]) );
  OR U5223 ( .A(n5009), .B(n4967), .Z(n5008) );
  NANDN U5224 ( .A(n5010), .B(n5011), .Z(o[53]) );
  OR U5225 ( .A(n5012), .B(n4967), .Z(n5011) );
  NANDN U5226 ( .A(n5013), .B(n5014), .Z(o[52]) );
  OR U5227 ( .A(n5015), .B(n4967), .Z(n5014) );
  NANDN U5228 ( .A(n5016), .B(n5017), .Z(o[51]) );
  OR U5229 ( .A(n5018), .B(n4967), .Z(n5017) );
  NANDN U5230 ( .A(n5019), .B(n5020), .Z(o[50]) );
  OR U5231 ( .A(n5021), .B(n4967), .Z(n5020) );
  NANDN U5232 ( .A(n5022), .B(n5023), .Z(o[4]) );
  OR U5233 ( .A(n5024), .B(n4967), .Z(n5023) );
  NANDN U5234 ( .A(n5025), .B(n5026), .Z(o[49]) );
  OR U5235 ( .A(n5027), .B(n4967), .Z(n5026) );
  NANDN U5236 ( .A(n5028), .B(n5029), .Z(o[48]) );
  OR U5237 ( .A(n5030), .B(n4967), .Z(n5029) );
  NANDN U5238 ( .A(n5031), .B(n5032), .Z(o[47]) );
  OR U5239 ( .A(n5033), .B(n4967), .Z(n5032) );
  NANDN U5240 ( .A(n5034), .B(n5035), .Z(o[46]) );
  OR U5241 ( .A(n5036), .B(n4967), .Z(n5035) );
  NANDN U5242 ( .A(n5037), .B(n5038), .Z(o[45]) );
  OR U5243 ( .A(n5039), .B(n4967), .Z(n5038) );
  NANDN U5244 ( .A(n5040), .B(n5041), .Z(o[44]) );
  OR U5245 ( .A(n5042), .B(n4967), .Z(n5041) );
  NANDN U5246 ( .A(n5043), .B(n5044), .Z(o[43]) );
  OR U5247 ( .A(n5045), .B(n4967), .Z(n5044) );
  NANDN U5248 ( .A(n5046), .B(n5047), .Z(o[42]) );
  OR U5249 ( .A(n5048), .B(n4967), .Z(n5047) );
  NANDN U5250 ( .A(n5049), .B(n5050), .Z(o[41]) );
  OR U5251 ( .A(n5051), .B(n4967), .Z(n5050) );
  NANDN U5252 ( .A(n5052), .B(n5053), .Z(o[40]) );
  OR U5253 ( .A(n5054), .B(n4967), .Z(n5053) );
  NANDN U5254 ( .A(n5055), .B(n5056), .Z(o[3]) );
  OR U5255 ( .A(n5057), .B(n4967), .Z(n5056) );
  NANDN U5256 ( .A(n5058), .B(n5059), .Z(o[39]) );
  OR U5257 ( .A(n5060), .B(n4967), .Z(n5059) );
  NANDN U5258 ( .A(n5061), .B(n5062), .Z(o[38]) );
  OR U5259 ( .A(n5063), .B(n4967), .Z(n5062) );
  NANDN U5260 ( .A(n5064), .B(n5065), .Z(o[37]) );
  OR U5261 ( .A(n5066), .B(n4967), .Z(n5065) );
  NANDN U5262 ( .A(n5067), .B(n5068), .Z(o[36]) );
  OR U5263 ( .A(n5069), .B(n4967), .Z(n5068) );
  NANDN U5264 ( .A(n5070), .B(n5071), .Z(o[35]) );
  OR U5265 ( .A(n5072), .B(n4967), .Z(n5071) );
  NANDN U5266 ( .A(n5073), .B(n5074), .Z(o[34]) );
  OR U5267 ( .A(n5075), .B(n4967), .Z(n5074) );
  NANDN U5268 ( .A(n5076), .B(n5077), .Z(o[33]) );
  OR U5269 ( .A(n5078), .B(n4967), .Z(n5077) );
  NANDN U5270 ( .A(n5079), .B(n5080), .Z(o[32]) );
  OR U5271 ( .A(n5081), .B(n4967), .Z(n5080) );
  NANDN U5272 ( .A(n5082), .B(n5083), .Z(o[31]) );
  OR U5273 ( .A(n5084), .B(n4967), .Z(n5083) );
  NANDN U5274 ( .A(n5085), .B(n5086), .Z(o[30]) );
  OR U5275 ( .A(n5087), .B(n4967), .Z(n5086) );
  NANDN U5276 ( .A(n5088), .B(n5089), .Z(o[2]) );
  OR U5277 ( .A(n5090), .B(n4967), .Z(n5089) );
  NANDN U5278 ( .A(n5091), .B(n5092), .Z(o[29]) );
  OR U5279 ( .A(n5093), .B(n4967), .Z(n5092) );
  NANDN U5280 ( .A(n5094), .B(n5095), .Z(o[28]) );
  OR U5281 ( .A(n5096), .B(n4967), .Z(n5095) );
  NANDN U5282 ( .A(n5097), .B(n5098), .Z(o[27]) );
  OR U5283 ( .A(n5099), .B(n4967), .Z(n5098) );
  NANDN U5284 ( .A(n5100), .B(n5101), .Z(o[26]) );
  OR U5285 ( .A(n5102), .B(n4967), .Z(n5101) );
  NANDN U5286 ( .A(n5103), .B(n5104), .Z(o[25]) );
  OR U5287 ( .A(n5105), .B(n4967), .Z(n5104) );
  NANDN U5288 ( .A(n5106), .B(n5107), .Z(o[24]) );
  OR U5289 ( .A(n5108), .B(n4967), .Z(n5107) );
  NANDN U5290 ( .A(n5109), .B(n5110), .Z(o[23]) );
  OR U5291 ( .A(n5111), .B(n4967), .Z(n5110) );
  NANDN U5292 ( .A(n5112), .B(n5113), .Z(o[22]) );
  OR U5293 ( .A(n5114), .B(n4967), .Z(n5113) );
  NANDN U5294 ( .A(n5115), .B(n5116), .Z(o[21]) );
  OR U5295 ( .A(n5117), .B(n4967), .Z(n5116) );
  NANDN U5296 ( .A(n5118), .B(n5119), .Z(o[20]) );
  OR U5297 ( .A(n5120), .B(n4967), .Z(n5119) );
  NANDN U5298 ( .A(n5121), .B(n5122), .Z(o[1]) );
  OR U5299 ( .A(n5123), .B(n4967), .Z(n5122) );
  NANDN U5300 ( .A(n5124), .B(n5125), .Z(o[19]) );
  OR U5301 ( .A(n5126), .B(n4967), .Z(n5125) );
  NANDN U5302 ( .A(n5127), .B(n5128), .Z(o[18]) );
  OR U5303 ( .A(n5129), .B(n4967), .Z(n5128) );
  NANDN U5304 ( .A(n5130), .B(n5131), .Z(o[17]) );
  OR U5305 ( .A(n5132), .B(n4967), .Z(n5131) );
  NANDN U5306 ( .A(n5133), .B(n5134), .Z(o[16]) );
  OR U5307 ( .A(n5135), .B(n4967), .Z(n5134) );
  NANDN U5308 ( .A(n5136), .B(n5137), .Z(o[15]) );
  OR U5309 ( .A(n5138), .B(n4967), .Z(n5137) );
  NANDN U5310 ( .A(n5139), .B(n5140), .Z(o[14]) );
  OR U5311 ( .A(n5141), .B(n4967), .Z(n5140) );
  NANDN U5312 ( .A(n5142), .B(n5143), .Z(o[13]) );
  OR U5313 ( .A(n5144), .B(n4967), .Z(n5143) );
  NANDN U5314 ( .A(n5145), .B(n5146), .Z(o[12]) );
  OR U5315 ( .A(n5147), .B(n4967), .Z(n5146) );
  NANDN U5316 ( .A(n5148), .B(n5149), .Z(o[11]) );
  OR U5317 ( .A(n5150), .B(n4967), .Z(n5149) );
  NANDN U5318 ( .A(n5151), .B(n5152), .Z(o[10]) );
  OR U5319 ( .A(n5153), .B(n4967), .Z(n5152) );
  NANDN U5320 ( .A(n5154), .B(n5155), .Z(o[0]) );
  OR U5321 ( .A(n5156), .B(n4967), .Z(n5155) );
  NAND U5322 ( .A(n5157), .B(n5158), .Z(n4963) );
  OR U5323 ( .A(n5159), .B(n5160), .Z(n5158) );
  ANDN U5324 ( .B(n5161), .A(n5154), .Z(n5157) );
  AND U5325 ( .A(x[0]), .B(n4967), .Z(n5154) );
  NANDN U5326 ( .A(n5156), .B(n5162), .Z(n5161) );
  AND U5327 ( .A(n5163), .B(n5164), .Z(n5156) );
  AND U5328 ( .A(n5165), .B(n5166), .Z(n5164) );
  NAND U5329 ( .A(n5167), .B(n5168), .Z(n5166) );
  ANDN U5330 ( .B(\stack[0][0] ), .A(n5169), .Z(n5167) );
  AND U5331 ( .A(n5170), .B(n5171), .Z(n5165) );
  NANDN U5332 ( .A(n5169), .B(n5172), .Z(n5171) );
  NOR U5333 ( .A(n5160), .B(n5173), .Z(n5172) );
  NAND U5334 ( .A(n5174), .B(n5175), .Z(n5170) );
  NANDN U5335 ( .A(\stack[0][0] ), .B(n5169), .Z(n5174) );
  AND U5336 ( .A(n5176), .B(n5177), .Z(n5163) );
  NANDN U5337 ( .A(n5160), .B(n5178), .Z(n5177) );
  XNOR U5338 ( .A(n5179), .B(n5180), .Z(n5176) );
  XOR U5339 ( .A(n5181), .B(n5182), .Z(n5180) );
  NAND U5340 ( .A(n5183), .B(n5184), .Z(n4962) );
  NANDN U5341 ( .A(n5159), .B(\stack[0][1] ), .Z(n5184) );
  ANDN U5342 ( .B(n5185), .A(n5121), .Z(n5183) );
  AND U5343 ( .A(x[1]), .B(n4967), .Z(n5121) );
  NANDN U5344 ( .A(n5123), .B(n5162), .Z(n5185) );
  AND U5345 ( .A(n5186), .B(n5187), .Z(n5123) );
  AND U5346 ( .A(n5188), .B(n5189), .Z(n5187) );
  NAND U5347 ( .A(n5190), .B(n5168), .Z(n5189) );
  XOR U5348 ( .A(n5191), .B(n5192), .Z(n5190) );
  AND U5349 ( .A(n5193), .B(n5194), .Z(n5188) );
  NANDN U5350 ( .A(n5195), .B(n5196), .Z(n5194) );
  ANDN U5351 ( .B(\stack[0][1] ), .A(n5173), .Z(n5196) );
  NAND U5352 ( .A(n5197), .B(n5175), .Z(n5193) );
  OR U5353 ( .A(\stack[0][1] ), .B(\stack[1][1] ), .Z(n5197) );
  AND U5354 ( .A(n5198), .B(n5199), .Z(n5186) );
  NAND U5355 ( .A(\stack[0][1] ), .B(n5178), .Z(n5199) );
  XOR U5356 ( .A(n5200), .B(n5201), .Z(n5198) );
  XNOR U5357 ( .A(n5202), .B(n5203), .Z(n5201) );
  NAND U5358 ( .A(n5204), .B(n5205), .Z(n4961) );
  OR U5359 ( .A(n5159), .B(n5206), .Z(n5205) );
  ANDN U5360 ( .B(n5207), .A(n5088), .Z(n5204) );
  AND U5361 ( .A(x[2]), .B(n4967), .Z(n5088) );
  NANDN U5362 ( .A(n5090), .B(n5162), .Z(n5207) );
  AND U5363 ( .A(n5208), .B(n5209), .Z(n5090) );
  AND U5364 ( .A(n5210), .B(n5211), .Z(n5209) );
  NAND U5365 ( .A(n5212), .B(n5168), .Z(n5211) );
  XNOR U5366 ( .A(n5213), .B(n5214), .Z(n5212) );
  XNOR U5367 ( .A(n5215), .B(n5216), .Z(n5214) );
  AND U5368 ( .A(n5217), .B(n5218), .Z(n5210) );
  NANDN U5369 ( .A(n5219), .B(n5220), .Z(n5218) );
  NOR U5370 ( .A(n5206), .B(n5173), .Z(n5220) );
  NAND U5371 ( .A(n5221), .B(n5175), .Z(n5217) );
  NANDN U5372 ( .A(\stack[0][2] ), .B(n5219), .Z(n5221) );
  AND U5373 ( .A(n5222), .B(n5223), .Z(n5208) );
  NANDN U5374 ( .A(n5206), .B(n5178), .Z(n5223) );
  XOR U5375 ( .A(n5224), .B(n5225), .Z(n5222) );
  XNOR U5376 ( .A(n5226), .B(n5227), .Z(n5225) );
  NAND U5377 ( .A(n5228), .B(n5229), .Z(n4960) );
  OR U5378 ( .A(n5159), .B(n5230), .Z(n5229) );
  ANDN U5379 ( .B(n5231), .A(n5055), .Z(n5228) );
  AND U5380 ( .A(x[3]), .B(n4967), .Z(n5055) );
  NANDN U5381 ( .A(n5057), .B(n5162), .Z(n5231) );
  AND U5382 ( .A(n5232), .B(n5233), .Z(n5057) );
  AND U5383 ( .A(n5234), .B(n5235), .Z(n5233) );
  NAND U5384 ( .A(n5236), .B(n5168), .Z(n5235) );
  XNOR U5385 ( .A(n5237), .B(n5238), .Z(n5236) );
  XNOR U5386 ( .A(n5239), .B(n5240), .Z(n5238) );
  AND U5387 ( .A(n5241), .B(n5242), .Z(n5234) );
  NANDN U5388 ( .A(n5243), .B(n5244), .Z(n5242) );
  NOR U5389 ( .A(n5230), .B(n5173), .Z(n5244) );
  NAND U5390 ( .A(n5245), .B(n5175), .Z(n5241) );
  NANDN U5391 ( .A(\stack[0][3] ), .B(n5243), .Z(n5245) );
  AND U5392 ( .A(n5246), .B(n5247), .Z(n5232) );
  NANDN U5393 ( .A(n5230), .B(n5178), .Z(n5247) );
  XOR U5394 ( .A(n5248), .B(n5249), .Z(n5246) );
  XNOR U5395 ( .A(n5250), .B(n5251), .Z(n5249) );
  NAND U5396 ( .A(n5252), .B(n5253), .Z(n4959) );
  OR U5397 ( .A(n5159), .B(n5254), .Z(n5253) );
  ANDN U5398 ( .B(n5255), .A(n5022), .Z(n5252) );
  AND U5399 ( .A(x[4]), .B(n4967), .Z(n5022) );
  NANDN U5400 ( .A(n5024), .B(n5162), .Z(n5255) );
  AND U5401 ( .A(n5256), .B(n5257), .Z(n5024) );
  AND U5402 ( .A(n5258), .B(n5259), .Z(n5257) );
  NAND U5403 ( .A(n5260), .B(n5168), .Z(n5259) );
  XNOR U5404 ( .A(n5261), .B(n5262), .Z(n5260) );
  XNOR U5405 ( .A(n5263), .B(n5264), .Z(n5262) );
  AND U5406 ( .A(n5265), .B(n5266), .Z(n5258) );
  NANDN U5407 ( .A(n5267), .B(n5268), .Z(n5266) );
  NOR U5408 ( .A(n5254), .B(n5173), .Z(n5268) );
  NAND U5409 ( .A(n5269), .B(n5175), .Z(n5265) );
  NANDN U5410 ( .A(\stack[0][4] ), .B(n5267), .Z(n5269) );
  AND U5411 ( .A(n5270), .B(n5271), .Z(n5256) );
  NANDN U5412 ( .A(n5254), .B(n5178), .Z(n5271) );
  XOR U5413 ( .A(n5272), .B(n5273), .Z(n5270) );
  XNOR U5414 ( .A(n5274), .B(n5275), .Z(n5273) );
  NAND U5415 ( .A(n5276), .B(n5277), .Z(n4958) );
  OR U5416 ( .A(n5159), .B(n5278), .Z(n5277) );
  ANDN U5417 ( .B(n5279), .A(n4989), .Z(n5276) );
  AND U5418 ( .A(x[5]), .B(n4967), .Z(n4989) );
  NANDN U5419 ( .A(n4991), .B(n5162), .Z(n5279) );
  AND U5420 ( .A(n5280), .B(n5281), .Z(n4991) );
  AND U5421 ( .A(n5282), .B(n5283), .Z(n5281) );
  NAND U5422 ( .A(n5284), .B(n5168), .Z(n5283) );
  XNOR U5423 ( .A(n5285), .B(n5286), .Z(n5284) );
  XOR U5424 ( .A(n5287), .B(n5288), .Z(n5286) );
  AND U5425 ( .A(n5289), .B(n5290), .Z(n5282) );
  NANDN U5426 ( .A(n5278), .B(n5291), .Z(n5290) );
  NOR U5427 ( .A(n5292), .B(n5173), .Z(n5291) );
  NAND U5428 ( .A(n5293), .B(n5175), .Z(n5289) );
  NANDN U5429 ( .A(\stack[0][5] ), .B(n5292), .Z(n5293) );
  AND U5430 ( .A(n5294), .B(n5295), .Z(n5280) );
  NANDN U5431 ( .A(n5278), .B(n5178), .Z(n5295) );
  XOR U5432 ( .A(n5296), .B(n5297), .Z(n5294) );
  XNOR U5433 ( .A(n5298), .B(n5299), .Z(n5297) );
  NAND U5434 ( .A(n5300), .B(n5301), .Z(n4957) );
  OR U5435 ( .A(n5159), .B(n5302), .Z(n5301) );
  ANDN U5436 ( .B(n5303), .A(n4974), .Z(n5300) );
  AND U5437 ( .A(x[6]), .B(n4967), .Z(n4974) );
  NANDN U5438 ( .A(n4976), .B(n5162), .Z(n5303) );
  AND U5439 ( .A(n5304), .B(n5305), .Z(n4976) );
  AND U5440 ( .A(n5306), .B(n5307), .Z(n5305) );
  NAND U5441 ( .A(n5308), .B(n5168), .Z(n5307) );
  XNOR U5442 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U5443 ( .A(n5311), .B(n5312), .Z(n5310) );
  AND U5444 ( .A(n5313), .B(n5314), .Z(n5306) );
  NANDN U5445 ( .A(n5302), .B(n5315), .Z(n5314) );
  NOR U5446 ( .A(n5316), .B(n5173), .Z(n5315) );
  NAND U5447 ( .A(n5317), .B(n5175), .Z(n5313) );
  NANDN U5448 ( .A(\stack[0][6] ), .B(n5316), .Z(n5317) );
  AND U5449 ( .A(n5318), .B(n5319), .Z(n5304) );
  NANDN U5450 ( .A(n5302), .B(n5178), .Z(n5319) );
  XOR U5451 ( .A(n5320), .B(n5321), .Z(n5318) );
  XNOR U5452 ( .A(n5322), .B(n5323), .Z(n5321) );
  NAND U5453 ( .A(n5324), .B(n5325), .Z(n4956) );
  OR U5454 ( .A(n5159), .B(n5326), .Z(n5325) );
  ANDN U5455 ( .B(n5327), .A(n4971), .Z(n5324) );
  AND U5456 ( .A(x[7]), .B(n4967), .Z(n4971) );
  NANDN U5457 ( .A(n4973), .B(n5162), .Z(n5327) );
  AND U5458 ( .A(n5328), .B(n5329), .Z(n4973) );
  AND U5459 ( .A(n5330), .B(n5331), .Z(n5329) );
  NAND U5460 ( .A(n5332), .B(n5168), .Z(n5331) );
  XNOR U5461 ( .A(n5333), .B(n5334), .Z(n5332) );
  XOR U5462 ( .A(n5335), .B(n5336), .Z(n5334) );
  AND U5463 ( .A(n5337), .B(n5338), .Z(n5330) );
  NANDN U5464 ( .A(n5326), .B(n5339), .Z(n5338) );
  NOR U5465 ( .A(n5340), .B(n5173), .Z(n5339) );
  NAND U5466 ( .A(n5341), .B(n5175), .Z(n5337) );
  NANDN U5467 ( .A(\stack[0][7] ), .B(n5340), .Z(n5341) );
  AND U5468 ( .A(n5342), .B(n5343), .Z(n5328) );
  NANDN U5469 ( .A(n5326), .B(n5178), .Z(n5343) );
  XOR U5470 ( .A(n5344), .B(n5345), .Z(n5342) );
  XNOR U5471 ( .A(n5346), .B(n5347), .Z(n5345) );
  NAND U5472 ( .A(n5348), .B(n5349), .Z(n4955) );
  OR U5473 ( .A(n5159), .B(n5350), .Z(n5349) );
  ANDN U5474 ( .B(n5351), .A(n4968), .Z(n5348) );
  AND U5475 ( .A(x[8]), .B(n4967), .Z(n4968) );
  NANDN U5476 ( .A(n4970), .B(n5162), .Z(n5351) );
  AND U5477 ( .A(n5352), .B(n5353), .Z(n4970) );
  AND U5478 ( .A(n5354), .B(n5355), .Z(n5353) );
  NAND U5479 ( .A(n5356), .B(n5168), .Z(n5355) );
  XNOR U5480 ( .A(n5357), .B(n5358), .Z(n5356) );
  XNOR U5481 ( .A(n5359), .B(n5360), .Z(n5358) );
  AND U5482 ( .A(n5361), .B(n5362), .Z(n5354) );
  NANDN U5483 ( .A(n5350), .B(n5363), .Z(n5362) );
  NOR U5484 ( .A(n5364), .B(n5173), .Z(n5363) );
  NAND U5485 ( .A(n5365), .B(n5175), .Z(n5361) );
  NANDN U5486 ( .A(\stack[0][8] ), .B(n5364), .Z(n5365) );
  AND U5487 ( .A(n5366), .B(n5367), .Z(n5352) );
  NANDN U5488 ( .A(n5350), .B(n5178), .Z(n5367) );
  XOR U5489 ( .A(n5368), .B(n5369), .Z(n5366) );
  XNOR U5490 ( .A(n5370), .B(n5371), .Z(n5369) );
  NAND U5491 ( .A(n5372), .B(n5373), .Z(n4954) );
  OR U5492 ( .A(n5159), .B(n5374), .Z(n5373) );
  ANDN U5493 ( .B(n5375), .A(n4964), .Z(n5372) );
  AND U5494 ( .A(x[9]), .B(n4967), .Z(n4964) );
  NANDN U5495 ( .A(n4966), .B(n5162), .Z(n5375) );
  AND U5496 ( .A(n5376), .B(n5377), .Z(n4966) );
  AND U5497 ( .A(n5378), .B(n5379), .Z(n5377) );
  NAND U5498 ( .A(n5380), .B(n5168), .Z(n5379) );
  XNOR U5499 ( .A(n5381), .B(n5382), .Z(n5380) );
  AND U5500 ( .A(n5385), .B(n5386), .Z(n5378) );
  NANDN U5501 ( .A(n5387), .B(n5388), .Z(n5386) );
  NOR U5502 ( .A(n5374), .B(n5173), .Z(n5388) );
  NAND U5503 ( .A(n5389), .B(n5175), .Z(n5385) );
  NANDN U5504 ( .A(\stack[0][9] ), .B(n5387), .Z(n5389) );
  AND U5505 ( .A(n5390), .B(n5391), .Z(n5376) );
  NANDN U5506 ( .A(n5374), .B(n5178), .Z(n5391) );
  XNOR U5507 ( .A(n5392), .B(n5393), .Z(n5390) );
  XNOR U5508 ( .A(n5394), .B(n5395), .Z(n5393) );
  NAND U5509 ( .A(n5396), .B(n5397), .Z(n4953) );
  OR U5510 ( .A(n5159), .B(n5398), .Z(n5397) );
  ANDN U5511 ( .B(n5399), .A(n5151), .Z(n5396) );
  AND U5512 ( .A(x[10]), .B(n4967), .Z(n5151) );
  NANDN U5513 ( .A(n5153), .B(n5162), .Z(n5399) );
  AND U5514 ( .A(n5400), .B(n5401), .Z(n5153) );
  AND U5515 ( .A(n5402), .B(n5403), .Z(n5401) );
  NAND U5516 ( .A(n5404), .B(n5168), .Z(n5403) );
  XNOR U5517 ( .A(n5405), .B(n5406), .Z(n5404) );
  XNOR U5518 ( .A(n5407), .B(n5408), .Z(n5406) );
  AND U5519 ( .A(n5409), .B(n5410), .Z(n5402) );
  NANDN U5520 ( .A(n5411), .B(n5412), .Z(n5410) );
  NOR U5521 ( .A(n5398), .B(n5173), .Z(n5412) );
  NAND U5522 ( .A(n5413), .B(n5175), .Z(n5409) );
  NANDN U5523 ( .A(\stack[0][10] ), .B(n5411), .Z(n5413) );
  AND U5524 ( .A(n5414), .B(n5415), .Z(n5400) );
  NANDN U5525 ( .A(n5398), .B(n5178), .Z(n5415) );
  XOR U5526 ( .A(n5416), .B(n5417), .Z(n5414) );
  XNOR U5527 ( .A(n5418), .B(n5419), .Z(n5417) );
  NAND U5528 ( .A(n5420), .B(n5421), .Z(n4952) );
  OR U5529 ( .A(n5159), .B(n5422), .Z(n5421) );
  ANDN U5530 ( .B(n5423), .A(n5148), .Z(n5420) );
  AND U5531 ( .A(x[11]), .B(n4967), .Z(n5148) );
  NANDN U5532 ( .A(n5150), .B(n5162), .Z(n5423) );
  AND U5533 ( .A(n5424), .B(n5425), .Z(n5150) );
  AND U5534 ( .A(n5426), .B(n5427), .Z(n5425) );
  NAND U5535 ( .A(n5428), .B(n5168), .Z(n5427) );
  XNOR U5536 ( .A(n5429), .B(n5430), .Z(n5428) );
  XOR U5537 ( .A(n5431), .B(n5432), .Z(n5430) );
  AND U5538 ( .A(n5433), .B(n5434), .Z(n5426) );
  NANDN U5539 ( .A(n5435), .B(n5436), .Z(n5434) );
  NOR U5540 ( .A(n5422), .B(n5173), .Z(n5436) );
  NAND U5541 ( .A(n5437), .B(n5175), .Z(n5433) );
  NANDN U5542 ( .A(\stack[0][11] ), .B(n5435), .Z(n5437) );
  AND U5543 ( .A(n5438), .B(n5439), .Z(n5424) );
  NANDN U5544 ( .A(n5422), .B(n5178), .Z(n5439) );
  XOR U5545 ( .A(n5440), .B(n5441), .Z(n5438) );
  XNOR U5546 ( .A(n5442), .B(n5443), .Z(n5441) );
  NAND U5547 ( .A(n5444), .B(n5445), .Z(n4951) );
  OR U5548 ( .A(n5159), .B(n5446), .Z(n5445) );
  ANDN U5549 ( .B(n5447), .A(n5145), .Z(n5444) );
  AND U5550 ( .A(x[12]), .B(n4967), .Z(n5145) );
  NANDN U5551 ( .A(n5147), .B(n5162), .Z(n5447) );
  AND U5552 ( .A(n5448), .B(n5449), .Z(n5147) );
  AND U5553 ( .A(n5450), .B(n5451), .Z(n5449) );
  NAND U5554 ( .A(n5452), .B(n5168), .Z(n5451) );
  XOR U5555 ( .A(n5453), .B(n5454), .Z(n5452) );
  XNOR U5556 ( .A(n5455), .B(n5456), .Z(n5454) );
  AND U5557 ( .A(n5457), .B(n5458), .Z(n5450) );
  NANDN U5558 ( .A(n5459), .B(n5460), .Z(n5458) );
  NOR U5559 ( .A(n5446), .B(n5173), .Z(n5460) );
  NAND U5560 ( .A(n5461), .B(n5175), .Z(n5457) );
  NANDN U5561 ( .A(\stack[0][12] ), .B(n5459), .Z(n5461) );
  AND U5562 ( .A(n5462), .B(n5463), .Z(n5448) );
  NANDN U5563 ( .A(n5446), .B(n5178), .Z(n5463) );
  XOR U5564 ( .A(n5464), .B(n5465), .Z(n5462) );
  XNOR U5565 ( .A(n5466), .B(n5467), .Z(n5465) );
  NAND U5566 ( .A(n5468), .B(n5469), .Z(n4950) );
  OR U5567 ( .A(n5159), .B(n5470), .Z(n5469) );
  ANDN U5568 ( .B(n5471), .A(n5142), .Z(n5468) );
  AND U5569 ( .A(x[13]), .B(n4967), .Z(n5142) );
  NANDN U5570 ( .A(n5144), .B(n5162), .Z(n5471) );
  AND U5571 ( .A(n5472), .B(n5473), .Z(n5144) );
  AND U5572 ( .A(n5474), .B(n5475), .Z(n5473) );
  NAND U5573 ( .A(n5476), .B(n5168), .Z(n5475) );
  XOR U5574 ( .A(n5477), .B(n5478), .Z(n5476) );
  XNOR U5575 ( .A(n5479), .B(n5480), .Z(n5478) );
  AND U5576 ( .A(n5481), .B(n5482), .Z(n5474) );
  NANDN U5577 ( .A(n5483), .B(n5484), .Z(n5482) );
  NOR U5578 ( .A(n5470), .B(n5173), .Z(n5484) );
  NAND U5579 ( .A(n5485), .B(n5175), .Z(n5481) );
  NANDN U5580 ( .A(\stack[0][13] ), .B(n5483), .Z(n5485) );
  AND U5581 ( .A(n5486), .B(n5487), .Z(n5472) );
  NANDN U5582 ( .A(n5470), .B(n5178), .Z(n5487) );
  XOR U5583 ( .A(n5488), .B(n5489), .Z(n5486) );
  XNOR U5584 ( .A(n5490), .B(n5491), .Z(n5489) );
  NAND U5585 ( .A(n5492), .B(n5493), .Z(n4949) );
  OR U5586 ( .A(n5159), .B(n5494), .Z(n5493) );
  ANDN U5587 ( .B(n5495), .A(n5139), .Z(n5492) );
  AND U5588 ( .A(x[14]), .B(n4967), .Z(n5139) );
  NANDN U5589 ( .A(n5141), .B(n5162), .Z(n5495) );
  AND U5590 ( .A(n5496), .B(n5497), .Z(n5141) );
  AND U5591 ( .A(n5498), .B(n5499), .Z(n5497) );
  NAND U5592 ( .A(n5500), .B(n5168), .Z(n5499) );
  XOR U5593 ( .A(n5501), .B(n5502), .Z(n5500) );
  XNOR U5594 ( .A(n5503), .B(n5504), .Z(n5502) );
  AND U5595 ( .A(n5505), .B(n5506), .Z(n5498) );
  NANDN U5596 ( .A(n5507), .B(n5508), .Z(n5506) );
  NOR U5597 ( .A(n5494), .B(n5173), .Z(n5508) );
  NAND U5598 ( .A(n5509), .B(n5175), .Z(n5505) );
  NANDN U5599 ( .A(\stack[0][14] ), .B(n5507), .Z(n5509) );
  AND U5600 ( .A(n5510), .B(n5511), .Z(n5496) );
  NANDN U5601 ( .A(n5494), .B(n5178), .Z(n5511) );
  XOR U5602 ( .A(n5512), .B(n5513), .Z(n5510) );
  XNOR U5603 ( .A(n5514), .B(n5515), .Z(n5513) );
  NAND U5604 ( .A(n5516), .B(n5517), .Z(n4948) );
  OR U5605 ( .A(n5159), .B(n5518), .Z(n5517) );
  ANDN U5606 ( .B(n5519), .A(n5136), .Z(n5516) );
  AND U5607 ( .A(x[15]), .B(n4967), .Z(n5136) );
  NANDN U5608 ( .A(n5138), .B(n5162), .Z(n5519) );
  AND U5609 ( .A(n5520), .B(n5521), .Z(n5138) );
  AND U5610 ( .A(n5522), .B(n5523), .Z(n5521) );
  NAND U5611 ( .A(n5524), .B(n5168), .Z(n5523) );
  XOR U5612 ( .A(n5525), .B(n5526), .Z(n5524) );
  XNOR U5613 ( .A(n5527), .B(n5528), .Z(n5526) );
  AND U5614 ( .A(n5529), .B(n5530), .Z(n5522) );
  NANDN U5615 ( .A(n5531), .B(n5532), .Z(n5530) );
  NOR U5616 ( .A(n5518), .B(n5173), .Z(n5532) );
  NAND U5617 ( .A(n5533), .B(n5175), .Z(n5529) );
  NANDN U5618 ( .A(\stack[0][15] ), .B(n5531), .Z(n5533) );
  AND U5619 ( .A(n5534), .B(n5535), .Z(n5520) );
  NANDN U5620 ( .A(n5518), .B(n5178), .Z(n5535) );
  XOR U5621 ( .A(n5536), .B(n5537), .Z(n5534) );
  XNOR U5622 ( .A(n5538), .B(n5539), .Z(n5537) );
  NAND U5623 ( .A(n5540), .B(n5541), .Z(n4947) );
  OR U5624 ( .A(n5159), .B(n5542), .Z(n5541) );
  ANDN U5625 ( .B(n5543), .A(n5133), .Z(n5540) );
  AND U5626 ( .A(x[16]), .B(n4967), .Z(n5133) );
  NANDN U5627 ( .A(n5135), .B(n5162), .Z(n5543) );
  AND U5628 ( .A(n5544), .B(n5545), .Z(n5135) );
  AND U5629 ( .A(n5546), .B(n5547), .Z(n5545) );
  NAND U5630 ( .A(n5548), .B(n5168), .Z(n5547) );
  XOR U5631 ( .A(n5549), .B(n5550), .Z(n5548) );
  XNOR U5632 ( .A(n5551), .B(n5552), .Z(n5550) );
  AND U5633 ( .A(n5553), .B(n5554), .Z(n5546) );
  NANDN U5634 ( .A(n5555), .B(n5556), .Z(n5554) );
  NOR U5635 ( .A(n5542), .B(n5173), .Z(n5556) );
  NAND U5636 ( .A(n5557), .B(n5175), .Z(n5553) );
  NANDN U5637 ( .A(\stack[0][16] ), .B(n5555), .Z(n5557) );
  AND U5638 ( .A(n5558), .B(n5559), .Z(n5544) );
  NANDN U5639 ( .A(n5542), .B(n5178), .Z(n5559) );
  XOR U5640 ( .A(n5560), .B(n5561), .Z(n5558) );
  XNOR U5641 ( .A(n5562), .B(n5563), .Z(n5561) );
  NAND U5642 ( .A(n5564), .B(n5565), .Z(n4946) );
  OR U5643 ( .A(n5159), .B(n5566), .Z(n5565) );
  ANDN U5644 ( .B(n5567), .A(n5130), .Z(n5564) );
  AND U5645 ( .A(x[17]), .B(n4967), .Z(n5130) );
  NANDN U5646 ( .A(n5132), .B(n5162), .Z(n5567) );
  AND U5647 ( .A(n5568), .B(n5569), .Z(n5132) );
  AND U5648 ( .A(n5570), .B(n5571), .Z(n5569) );
  NAND U5649 ( .A(n5572), .B(n5168), .Z(n5571) );
  XOR U5650 ( .A(n5573), .B(n5574), .Z(n5572) );
  XNOR U5651 ( .A(n5575), .B(n5576), .Z(n5574) );
  AND U5652 ( .A(n5577), .B(n5578), .Z(n5570) );
  NANDN U5653 ( .A(n5579), .B(n5580), .Z(n5578) );
  NOR U5654 ( .A(n5566), .B(n5173), .Z(n5580) );
  NAND U5655 ( .A(n5581), .B(n5175), .Z(n5577) );
  NANDN U5656 ( .A(\stack[0][17] ), .B(n5579), .Z(n5581) );
  AND U5657 ( .A(n5582), .B(n5583), .Z(n5568) );
  NANDN U5658 ( .A(n5566), .B(n5178), .Z(n5583) );
  XOR U5659 ( .A(n5584), .B(n5585), .Z(n5582) );
  XNOR U5660 ( .A(n5586), .B(n5587), .Z(n5585) );
  NAND U5661 ( .A(n5588), .B(n5589), .Z(n4945) );
  OR U5662 ( .A(n5159), .B(n5590), .Z(n5589) );
  ANDN U5663 ( .B(n5591), .A(n5127), .Z(n5588) );
  AND U5664 ( .A(x[18]), .B(n4967), .Z(n5127) );
  NANDN U5665 ( .A(n5129), .B(n5162), .Z(n5591) );
  AND U5666 ( .A(n5592), .B(n5593), .Z(n5129) );
  AND U5667 ( .A(n5594), .B(n5595), .Z(n5593) );
  NAND U5668 ( .A(n5596), .B(n5168), .Z(n5595) );
  XOR U5669 ( .A(n5597), .B(n5598), .Z(n5596) );
  XNOR U5670 ( .A(n5599), .B(n5600), .Z(n5598) );
  AND U5671 ( .A(n5601), .B(n5602), .Z(n5594) );
  NANDN U5672 ( .A(n5603), .B(n5604), .Z(n5602) );
  NOR U5673 ( .A(n5590), .B(n5173), .Z(n5604) );
  NAND U5674 ( .A(n5605), .B(n5175), .Z(n5601) );
  NANDN U5675 ( .A(\stack[0][18] ), .B(n5603), .Z(n5605) );
  AND U5676 ( .A(n5606), .B(n5607), .Z(n5592) );
  NANDN U5677 ( .A(n5590), .B(n5178), .Z(n5607) );
  XOR U5678 ( .A(n5608), .B(n5609), .Z(n5606) );
  XNOR U5679 ( .A(n5610), .B(n5611), .Z(n5609) );
  NAND U5680 ( .A(n5612), .B(n5613), .Z(n4944) );
  OR U5681 ( .A(n5159), .B(n5614), .Z(n5613) );
  ANDN U5682 ( .B(n5615), .A(n5124), .Z(n5612) );
  AND U5683 ( .A(x[19]), .B(n4967), .Z(n5124) );
  NANDN U5684 ( .A(n5126), .B(n5162), .Z(n5615) );
  AND U5685 ( .A(n5616), .B(n5617), .Z(n5126) );
  AND U5686 ( .A(n5618), .B(n5619), .Z(n5617) );
  NAND U5687 ( .A(n5620), .B(n5168), .Z(n5619) );
  XOR U5688 ( .A(n5621), .B(n5622), .Z(n5620) );
  XNOR U5689 ( .A(n5623), .B(n5624), .Z(n5622) );
  AND U5690 ( .A(n5625), .B(n5626), .Z(n5618) );
  NANDN U5691 ( .A(n5627), .B(n5628), .Z(n5626) );
  NOR U5692 ( .A(n5614), .B(n5173), .Z(n5628) );
  NAND U5693 ( .A(n5629), .B(n5175), .Z(n5625) );
  NANDN U5694 ( .A(\stack[0][19] ), .B(n5627), .Z(n5629) );
  AND U5695 ( .A(n5630), .B(n5631), .Z(n5616) );
  NANDN U5696 ( .A(n5614), .B(n5178), .Z(n5631) );
  XOR U5697 ( .A(n5632), .B(n5633), .Z(n5630) );
  XNOR U5698 ( .A(n5634), .B(n5635), .Z(n5633) );
  NAND U5699 ( .A(n5636), .B(n5637), .Z(n4943) );
  OR U5700 ( .A(n5159), .B(n5638), .Z(n5637) );
  ANDN U5701 ( .B(n5639), .A(n5118), .Z(n5636) );
  AND U5702 ( .A(x[20]), .B(n4967), .Z(n5118) );
  NANDN U5703 ( .A(n5120), .B(n5162), .Z(n5639) );
  AND U5704 ( .A(n5640), .B(n5641), .Z(n5120) );
  AND U5705 ( .A(n5642), .B(n5643), .Z(n5641) );
  NAND U5706 ( .A(n5644), .B(n5168), .Z(n5643) );
  XOR U5707 ( .A(n5645), .B(n5646), .Z(n5644) );
  XNOR U5708 ( .A(n5647), .B(n5648), .Z(n5646) );
  AND U5709 ( .A(n5649), .B(n5650), .Z(n5642) );
  NANDN U5710 ( .A(n5651), .B(n5652), .Z(n5650) );
  NOR U5711 ( .A(n5638), .B(n5173), .Z(n5652) );
  NAND U5712 ( .A(n5653), .B(n5175), .Z(n5649) );
  NANDN U5713 ( .A(\stack[0][20] ), .B(n5651), .Z(n5653) );
  AND U5714 ( .A(n5654), .B(n5655), .Z(n5640) );
  NANDN U5715 ( .A(n5638), .B(n5178), .Z(n5655) );
  XOR U5716 ( .A(n5656), .B(n5657), .Z(n5654) );
  XNOR U5717 ( .A(n5658), .B(n5659), .Z(n5657) );
  NAND U5718 ( .A(n5660), .B(n5661), .Z(n4942) );
  OR U5719 ( .A(n5159), .B(n5662), .Z(n5661) );
  ANDN U5720 ( .B(n5663), .A(n5115), .Z(n5660) );
  AND U5721 ( .A(x[21]), .B(n4967), .Z(n5115) );
  NANDN U5722 ( .A(n5117), .B(n5162), .Z(n5663) );
  AND U5723 ( .A(n5664), .B(n5665), .Z(n5117) );
  AND U5724 ( .A(n5666), .B(n5667), .Z(n5665) );
  NAND U5725 ( .A(n5668), .B(n5168), .Z(n5667) );
  XOR U5726 ( .A(n5669), .B(n5670), .Z(n5668) );
  XNOR U5727 ( .A(n5671), .B(n5672), .Z(n5670) );
  AND U5728 ( .A(n5673), .B(n5674), .Z(n5666) );
  NANDN U5729 ( .A(n5675), .B(n5676), .Z(n5674) );
  NOR U5730 ( .A(n5662), .B(n5173), .Z(n5676) );
  NAND U5731 ( .A(n5677), .B(n5175), .Z(n5673) );
  NANDN U5732 ( .A(\stack[0][21] ), .B(n5675), .Z(n5677) );
  AND U5733 ( .A(n5678), .B(n5679), .Z(n5664) );
  NANDN U5734 ( .A(n5662), .B(n5178), .Z(n5679) );
  XOR U5735 ( .A(n5680), .B(n5681), .Z(n5678) );
  XNOR U5736 ( .A(n5682), .B(n5683), .Z(n5681) );
  NAND U5737 ( .A(n5684), .B(n5685), .Z(n4941) );
  OR U5738 ( .A(n5159), .B(n5686), .Z(n5685) );
  ANDN U5739 ( .B(n5687), .A(n5112), .Z(n5684) );
  AND U5740 ( .A(x[22]), .B(n4967), .Z(n5112) );
  NANDN U5741 ( .A(n5114), .B(n5162), .Z(n5687) );
  AND U5742 ( .A(n5688), .B(n5689), .Z(n5114) );
  AND U5743 ( .A(n5690), .B(n5691), .Z(n5689) );
  NAND U5744 ( .A(n5692), .B(n5168), .Z(n5691) );
  XOR U5745 ( .A(n5693), .B(n5694), .Z(n5692) );
  XNOR U5746 ( .A(n5695), .B(n5696), .Z(n5694) );
  AND U5747 ( .A(n5697), .B(n5698), .Z(n5690) );
  NANDN U5748 ( .A(n5699), .B(n5700), .Z(n5698) );
  NOR U5749 ( .A(n5686), .B(n5173), .Z(n5700) );
  NAND U5750 ( .A(n5701), .B(n5175), .Z(n5697) );
  NANDN U5751 ( .A(\stack[0][22] ), .B(n5699), .Z(n5701) );
  AND U5752 ( .A(n5702), .B(n5703), .Z(n5688) );
  NANDN U5753 ( .A(n5686), .B(n5178), .Z(n5703) );
  XOR U5754 ( .A(n5704), .B(n5705), .Z(n5702) );
  XNOR U5755 ( .A(n5706), .B(n5707), .Z(n5705) );
  NAND U5756 ( .A(n5708), .B(n5709), .Z(n4940) );
  OR U5757 ( .A(n5159), .B(n5710), .Z(n5709) );
  ANDN U5758 ( .B(n5711), .A(n5109), .Z(n5708) );
  AND U5759 ( .A(x[23]), .B(n4967), .Z(n5109) );
  NANDN U5760 ( .A(n5111), .B(n5162), .Z(n5711) );
  AND U5761 ( .A(n5712), .B(n5713), .Z(n5111) );
  AND U5762 ( .A(n5714), .B(n5715), .Z(n5713) );
  NAND U5763 ( .A(n5716), .B(n5168), .Z(n5715) );
  XOR U5764 ( .A(n5717), .B(n5718), .Z(n5716) );
  XNOR U5765 ( .A(n5719), .B(n5720), .Z(n5718) );
  AND U5766 ( .A(n5721), .B(n5722), .Z(n5714) );
  NANDN U5767 ( .A(n5723), .B(n5724), .Z(n5722) );
  NOR U5768 ( .A(n5710), .B(n5173), .Z(n5724) );
  NAND U5769 ( .A(n5725), .B(n5175), .Z(n5721) );
  NANDN U5770 ( .A(\stack[0][23] ), .B(n5723), .Z(n5725) );
  AND U5771 ( .A(n5726), .B(n5727), .Z(n5712) );
  NANDN U5772 ( .A(n5710), .B(n5178), .Z(n5727) );
  XOR U5773 ( .A(n5728), .B(n5729), .Z(n5726) );
  XNOR U5774 ( .A(n5730), .B(n5731), .Z(n5729) );
  NAND U5775 ( .A(n5732), .B(n5733), .Z(n4939) );
  OR U5776 ( .A(n5159), .B(n5734), .Z(n5733) );
  ANDN U5777 ( .B(n5735), .A(n5106), .Z(n5732) );
  AND U5778 ( .A(x[24]), .B(n4967), .Z(n5106) );
  NANDN U5779 ( .A(n5108), .B(n5162), .Z(n5735) );
  AND U5780 ( .A(n5736), .B(n5737), .Z(n5108) );
  AND U5781 ( .A(n5738), .B(n5739), .Z(n5737) );
  NAND U5782 ( .A(n5740), .B(n5168), .Z(n5739) );
  XOR U5783 ( .A(n5741), .B(n5742), .Z(n5740) );
  XNOR U5784 ( .A(n5743), .B(n5744), .Z(n5742) );
  AND U5785 ( .A(n5745), .B(n5746), .Z(n5738) );
  NANDN U5786 ( .A(n5747), .B(n5748), .Z(n5746) );
  NOR U5787 ( .A(n5734), .B(n5173), .Z(n5748) );
  NAND U5788 ( .A(n5749), .B(n5175), .Z(n5745) );
  NANDN U5789 ( .A(\stack[0][24] ), .B(n5747), .Z(n5749) );
  AND U5790 ( .A(n5750), .B(n5751), .Z(n5736) );
  NANDN U5791 ( .A(n5734), .B(n5178), .Z(n5751) );
  XOR U5792 ( .A(n5752), .B(n5753), .Z(n5750) );
  XNOR U5793 ( .A(n5754), .B(n5755), .Z(n5753) );
  NAND U5794 ( .A(n5756), .B(n5757), .Z(n4938) );
  OR U5795 ( .A(n5159), .B(n5758), .Z(n5757) );
  ANDN U5796 ( .B(n5759), .A(n5103), .Z(n5756) );
  AND U5797 ( .A(x[25]), .B(n4967), .Z(n5103) );
  NANDN U5798 ( .A(n5105), .B(n5162), .Z(n5759) );
  AND U5799 ( .A(n5760), .B(n5761), .Z(n5105) );
  AND U5800 ( .A(n5762), .B(n5763), .Z(n5761) );
  NAND U5801 ( .A(n5764), .B(n5168), .Z(n5763) );
  XOR U5802 ( .A(n5765), .B(n5766), .Z(n5764) );
  XNOR U5803 ( .A(n5767), .B(n5768), .Z(n5766) );
  AND U5804 ( .A(n5769), .B(n5770), .Z(n5762) );
  NANDN U5805 ( .A(n5771), .B(n5772), .Z(n5770) );
  NOR U5806 ( .A(n5758), .B(n5173), .Z(n5772) );
  NAND U5807 ( .A(n5773), .B(n5175), .Z(n5769) );
  NANDN U5808 ( .A(\stack[0][25] ), .B(n5771), .Z(n5773) );
  AND U5809 ( .A(n5774), .B(n5775), .Z(n5760) );
  NANDN U5810 ( .A(n5758), .B(n5178), .Z(n5775) );
  XOR U5811 ( .A(n5776), .B(n5777), .Z(n5774) );
  XNOR U5812 ( .A(n5778), .B(n5779), .Z(n5777) );
  NAND U5813 ( .A(n5780), .B(n5781), .Z(n4937) );
  OR U5814 ( .A(n5159), .B(n5782), .Z(n5781) );
  ANDN U5815 ( .B(n5783), .A(n5100), .Z(n5780) );
  AND U5816 ( .A(x[26]), .B(n4967), .Z(n5100) );
  NANDN U5817 ( .A(n5102), .B(n5162), .Z(n5783) );
  AND U5818 ( .A(n5784), .B(n5785), .Z(n5102) );
  AND U5819 ( .A(n5786), .B(n5787), .Z(n5785) );
  NAND U5820 ( .A(n5788), .B(n5168), .Z(n5787) );
  XOR U5821 ( .A(n5789), .B(n5790), .Z(n5788) );
  XNOR U5822 ( .A(n5791), .B(n5792), .Z(n5790) );
  AND U5823 ( .A(n5793), .B(n5794), .Z(n5786) );
  NANDN U5824 ( .A(n5795), .B(n5796), .Z(n5794) );
  NOR U5825 ( .A(n5782), .B(n5173), .Z(n5796) );
  NAND U5826 ( .A(n5797), .B(n5175), .Z(n5793) );
  NANDN U5827 ( .A(\stack[0][26] ), .B(n5795), .Z(n5797) );
  AND U5828 ( .A(n5798), .B(n5799), .Z(n5784) );
  NANDN U5829 ( .A(n5782), .B(n5178), .Z(n5799) );
  XOR U5830 ( .A(n5800), .B(n5801), .Z(n5798) );
  XNOR U5831 ( .A(n5802), .B(n5803), .Z(n5801) );
  NAND U5832 ( .A(n5804), .B(n5805), .Z(n4936) );
  OR U5833 ( .A(n5159), .B(n5806), .Z(n5805) );
  ANDN U5834 ( .B(n5807), .A(n5097), .Z(n5804) );
  AND U5835 ( .A(x[27]), .B(n4967), .Z(n5097) );
  NANDN U5836 ( .A(n5099), .B(n5162), .Z(n5807) );
  AND U5837 ( .A(n5808), .B(n5809), .Z(n5099) );
  AND U5838 ( .A(n5810), .B(n5811), .Z(n5809) );
  NAND U5839 ( .A(n5812), .B(n5168), .Z(n5811) );
  XOR U5840 ( .A(n5813), .B(n5814), .Z(n5812) );
  XNOR U5841 ( .A(n5815), .B(n5816), .Z(n5814) );
  AND U5842 ( .A(n5817), .B(n5818), .Z(n5810) );
  NANDN U5843 ( .A(n5819), .B(n5820), .Z(n5818) );
  NOR U5844 ( .A(n5806), .B(n5173), .Z(n5820) );
  NAND U5845 ( .A(n5821), .B(n5175), .Z(n5817) );
  NANDN U5846 ( .A(\stack[0][27] ), .B(n5819), .Z(n5821) );
  AND U5847 ( .A(n5822), .B(n5823), .Z(n5808) );
  NANDN U5848 ( .A(n5806), .B(n5178), .Z(n5823) );
  XOR U5849 ( .A(n5824), .B(n5825), .Z(n5822) );
  XNOR U5850 ( .A(n5826), .B(n5827), .Z(n5825) );
  NAND U5851 ( .A(n5828), .B(n5829), .Z(n4935) );
  OR U5852 ( .A(n5159), .B(n5830), .Z(n5829) );
  ANDN U5853 ( .B(n5831), .A(n5094), .Z(n5828) );
  AND U5854 ( .A(x[28]), .B(n4967), .Z(n5094) );
  NANDN U5855 ( .A(n5096), .B(n5162), .Z(n5831) );
  AND U5856 ( .A(n5832), .B(n5833), .Z(n5096) );
  AND U5857 ( .A(n5834), .B(n5835), .Z(n5833) );
  NAND U5858 ( .A(n5836), .B(n5168), .Z(n5835) );
  XOR U5859 ( .A(n5837), .B(n5838), .Z(n5836) );
  XNOR U5860 ( .A(n5839), .B(n5840), .Z(n5838) );
  AND U5861 ( .A(n5841), .B(n5842), .Z(n5834) );
  NANDN U5862 ( .A(n5843), .B(n5844), .Z(n5842) );
  NOR U5863 ( .A(n5830), .B(n5173), .Z(n5844) );
  NAND U5864 ( .A(n5845), .B(n5175), .Z(n5841) );
  NANDN U5865 ( .A(\stack[0][28] ), .B(n5843), .Z(n5845) );
  AND U5866 ( .A(n5846), .B(n5847), .Z(n5832) );
  NANDN U5867 ( .A(n5830), .B(n5178), .Z(n5847) );
  XOR U5868 ( .A(n5848), .B(n5849), .Z(n5846) );
  XNOR U5869 ( .A(n5850), .B(n5851), .Z(n5849) );
  NAND U5870 ( .A(n5852), .B(n5853), .Z(n4934) );
  OR U5871 ( .A(n5159), .B(n5854), .Z(n5853) );
  ANDN U5872 ( .B(n5855), .A(n5091), .Z(n5852) );
  AND U5873 ( .A(x[29]), .B(n4967), .Z(n5091) );
  NANDN U5874 ( .A(n5093), .B(n5162), .Z(n5855) );
  AND U5875 ( .A(n5856), .B(n5857), .Z(n5093) );
  AND U5876 ( .A(n5858), .B(n5859), .Z(n5857) );
  NAND U5877 ( .A(n5860), .B(n5168), .Z(n5859) );
  XOR U5878 ( .A(n5861), .B(n5862), .Z(n5860) );
  XNOR U5879 ( .A(n5863), .B(n5864), .Z(n5862) );
  AND U5880 ( .A(n5865), .B(n5866), .Z(n5858) );
  NANDN U5881 ( .A(n5867), .B(n5868), .Z(n5866) );
  NOR U5882 ( .A(n5854), .B(n5173), .Z(n5868) );
  NAND U5883 ( .A(n5869), .B(n5175), .Z(n5865) );
  NANDN U5884 ( .A(\stack[0][29] ), .B(n5867), .Z(n5869) );
  AND U5885 ( .A(n5870), .B(n5871), .Z(n5856) );
  NANDN U5886 ( .A(n5854), .B(n5178), .Z(n5871) );
  XOR U5887 ( .A(n5872), .B(n5873), .Z(n5870) );
  XNOR U5888 ( .A(n5874), .B(n5875), .Z(n5873) );
  NAND U5889 ( .A(n5876), .B(n5877), .Z(n4933) );
  OR U5890 ( .A(n5159), .B(n5878), .Z(n5877) );
  ANDN U5891 ( .B(n5879), .A(n5085), .Z(n5876) );
  AND U5892 ( .A(x[30]), .B(n4967), .Z(n5085) );
  NANDN U5893 ( .A(n5087), .B(n5162), .Z(n5879) );
  AND U5894 ( .A(n5880), .B(n5881), .Z(n5087) );
  AND U5895 ( .A(n5882), .B(n5883), .Z(n5881) );
  NAND U5896 ( .A(n5884), .B(n5168), .Z(n5883) );
  XOR U5897 ( .A(n5885), .B(n5886), .Z(n5884) );
  XNOR U5898 ( .A(n5887), .B(n5888), .Z(n5886) );
  AND U5899 ( .A(n5889), .B(n5890), .Z(n5882) );
  NANDN U5900 ( .A(n5891), .B(n5892), .Z(n5890) );
  NOR U5901 ( .A(n5878), .B(n5173), .Z(n5892) );
  NAND U5902 ( .A(n5893), .B(n5175), .Z(n5889) );
  NANDN U5903 ( .A(\stack[0][30] ), .B(n5891), .Z(n5893) );
  AND U5904 ( .A(n5894), .B(n5895), .Z(n5880) );
  NANDN U5905 ( .A(n5878), .B(n5178), .Z(n5895) );
  XOR U5906 ( .A(n5896), .B(n5897), .Z(n5894) );
  XNOR U5907 ( .A(n5898), .B(n5899), .Z(n5897) );
  NAND U5908 ( .A(n5900), .B(n5901), .Z(n4932) );
  OR U5909 ( .A(n5159), .B(n5902), .Z(n5901) );
  ANDN U5910 ( .B(n5903), .A(n5082), .Z(n5900) );
  AND U5911 ( .A(x[31]), .B(n4967), .Z(n5082) );
  NANDN U5912 ( .A(n5084), .B(n5162), .Z(n5903) );
  AND U5913 ( .A(n5904), .B(n5905), .Z(n5084) );
  AND U5914 ( .A(n5906), .B(n5907), .Z(n5905) );
  NAND U5915 ( .A(n5908), .B(n5168), .Z(n5907) );
  XOR U5916 ( .A(n5909), .B(n5910), .Z(n5908) );
  XNOR U5917 ( .A(n5911), .B(n5912), .Z(n5910) );
  AND U5918 ( .A(n5913), .B(n5914), .Z(n5906) );
  NANDN U5919 ( .A(n5915), .B(n5916), .Z(n5914) );
  NOR U5920 ( .A(n5902), .B(n5173), .Z(n5916) );
  NAND U5921 ( .A(n5917), .B(n5175), .Z(n5913) );
  NANDN U5922 ( .A(\stack[0][31] ), .B(n5915), .Z(n5917) );
  AND U5923 ( .A(n5918), .B(n5919), .Z(n5904) );
  NANDN U5924 ( .A(n5902), .B(n5178), .Z(n5919) );
  XOR U5925 ( .A(n5920), .B(n5921), .Z(n5918) );
  XNOR U5926 ( .A(n5922), .B(n5923), .Z(n5921) );
  NAND U5927 ( .A(n5924), .B(n5925), .Z(n4931) );
  OR U5928 ( .A(n5159), .B(n5926), .Z(n5925) );
  ANDN U5929 ( .B(n5927), .A(n5079), .Z(n5924) );
  AND U5930 ( .A(x[32]), .B(n4967), .Z(n5079) );
  NANDN U5931 ( .A(n5081), .B(n5162), .Z(n5927) );
  AND U5932 ( .A(n5928), .B(n5929), .Z(n5081) );
  AND U5933 ( .A(n5930), .B(n5931), .Z(n5929) );
  NAND U5934 ( .A(n5932), .B(n5168), .Z(n5931) );
  XOR U5935 ( .A(n5933), .B(n5934), .Z(n5932) );
  XNOR U5936 ( .A(n5935), .B(n5936), .Z(n5934) );
  AND U5937 ( .A(n5937), .B(n5938), .Z(n5930) );
  NANDN U5938 ( .A(n5926), .B(n5939), .Z(n5938) );
  NOR U5939 ( .A(n5940), .B(n5173), .Z(n5939) );
  NAND U5940 ( .A(n5941), .B(n5175), .Z(n5937) );
  NANDN U5941 ( .A(\stack[0][32] ), .B(n5940), .Z(n5941) );
  AND U5942 ( .A(n5942), .B(n5943), .Z(n5928) );
  NANDN U5943 ( .A(n5926), .B(n5178), .Z(n5943) );
  XOR U5944 ( .A(n5944), .B(n5945), .Z(n5942) );
  XNOR U5945 ( .A(n5946), .B(n5947), .Z(n5945) );
  NAND U5946 ( .A(n5948), .B(n5949), .Z(n4930) );
  OR U5947 ( .A(n5159), .B(n5950), .Z(n5949) );
  ANDN U5948 ( .B(n5951), .A(n5076), .Z(n5948) );
  AND U5949 ( .A(x[33]), .B(n4967), .Z(n5076) );
  NANDN U5950 ( .A(n5078), .B(n5162), .Z(n5951) );
  AND U5951 ( .A(n5952), .B(n5953), .Z(n5078) );
  AND U5952 ( .A(n5954), .B(n5955), .Z(n5953) );
  NAND U5953 ( .A(n5956), .B(n5168), .Z(n5955) );
  XOR U5954 ( .A(n5957), .B(n5958), .Z(n5956) );
  XNOR U5955 ( .A(n5959), .B(n5960), .Z(n5958) );
  AND U5956 ( .A(n5961), .B(n5962), .Z(n5954) );
  NANDN U5957 ( .A(n5950), .B(n5963), .Z(n5962) );
  NOR U5958 ( .A(n5964), .B(n5173), .Z(n5963) );
  NAND U5959 ( .A(n5965), .B(n5175), .Z(n5961) );
  NANDN U5960 ( .A(\stack[0][33] ), .B(n5964), .Z(n5965) );
  AND U5961 ( .A(n5966), .B(n5967), .Z(n5952) );
  NANDN U5962 ( .A(n5950), .B(n5178), .Z(n5967) );
  XOR U5963 ( .A(n5968), .B(n5969), .Z(n5966) );
  XNOR U5964 ( .A(n5970), .B(n5971), .Z(n5969) );
  NAND U5965 ( .A(n5972), .B(n5973), .Z(n4929) );
  OR U5966 ( .A(n5159), .B(n5974), .Z(n5973) );
  ANDN U5967 ( .B(n5975), .A(n5073), .Z(n5972) );
  AND U5968 ( .A(x[34]), .B(n4967), .Z(n5073) );
  NANDN U5969 ( .A(n5075), .B(n5162), .Z(n5975) );
  AND U5970 ( .A(n5976), .B(n5977), .Z(n5075) );
  AND U5971 ( .A(n5978), .B(n5979), .Z(n5977) );
  NAND U5972 ( .A(n5980), .B(n5168), .Z(n5979) );
  XOR U5973 ( .A(n5981), .B(n5982), .Z(n5980) );
  XNOR U5974 ( .A(n5983), .B(n5984), .Z(n5982) );
  AND U5975 ( .A(n5985), .B(n5986), .Z(n5978) );
  NANDN U5976 ( .A(n5974), .B(n5987), .Z(n5986) );
  NOR U5977 ( .A(n5988), .B(n5173), .Z(n5987) );
  NAND U5978 ( .A(n5989), .B(n5175), .Z(n5985) );
  NANDN U5979 ( .A(\stack[0][34] ), .B(n5988), .Z(n5989) );
  AND U5980 ( .A(n5990), .B(n5991), .Z(n5976) );
  NANDN U5981 ( .A(n5974), .B(n5178), .Z(n5991) );
  XOR U5982 ( .A(n5992), .B(n5993), .Z(n5990) );
  XNOR U5983 ( .A(n5994), .B(n5995), .Z(n5993) );
  NAND U5984 ( .A(n5996), .B(n5997), .Z(n4928) );
  OR U5985 ( .A(n5159), .B(n5998), .Z(n5997) );
  ANDN U5986 ( .B(n5999), .A(n5070), .Z(n5996) );
  AND U5987 ( .A(x[35]), .B(n4967), .Z(n5070) );
  NANDN U5988 ( .A(n5072), .B(n5162), .Z(n5999) );
  AND U5989 ( .A(n6000), .B(n6001), .Z(n5072) );
  AND U5990 ( .A(n6002), .B(n6003), .Z(n6001) );
  NAND U5991 ( .A(n6004), .B(n5168), .Z(n6003) );
  XOR U5992 ( .A(n6005), .B(n6006), .Z(n6004) );
  XNOR U5993 ( .A(n6007), .B(n6008), .Z(n6006) );
  AND U5994 ( .A(n6009), .B(n6010), .Z(n6002) );
  NANDN U5995 ( .A(n5998), .B(n6011), .Z(n6010) );
  NOR U5996 ( .A(n6012), .B(n5173), .Z(n6011) );
  NAND U5997 ( .A(n6013), .B(n5175), .Z(n6009) );
  NANDN U5998 ( .A(\stack[0][35] ), .B(n6012), .Z(n6013) );
  AND U5999 ( .A(n6014), .B(n6015), .Z(n6000) );
  NANDN U6000 ( .A(n5998), .B(n5178), .Z(n6015) );
  XOR U6001 ( .A(n6016), .B(n6017), .Z(n6014) );
  XNOR U6002 ( .A(n6018), .B(n6019), .Z(n6017) );
  NAND U6003 ( .A(n6020), .B(n6021), .Z(n4927) );
  OR U6004 ( .A(n5159), .B(n6022), .Z(n6021) );
  ANDN U6005 ( .B(n6023), .A(n5067), .Z(n6020) );
  AND U6006 ( .A(x[36]), .B(n4967), .Z(n5067) );
  NANDN U6007 ( .A(n5069), .B(n5162), .Z(n6023) );
  AND U6008 ( .A(n6024), .B(n6025), .Z(n5069) );
  AND U6009 ( .A(n6026), .B(n6027), .Z(n6025) );
  NAND U6010 ( .A(n6028), .B(n5168), .Z(n6027) );
  XOR U6011 ( .A(n6029), .B(n6030), .Z(n6028) );
  XNOR U6012 ( .A(n6031), .B(n6032), .Z(n6030) );
  AND U6013 ( .A(n6033), .B(n6034), .Z(n6026) );
  NANDN U6014 ( .A(n6022), .B(n6035), .Z(n6034) );
  NOR U6015 ( .A(n6036), .B(n5173), .Z(n6035) );
  NAND U6016 ( .A(n6037), .B(n5175), .Z(n6033) );
  NANDN U6017 ( .A(\stack[0][36] ), .B(n6036), .Z(n6037) );
  AND U6018 ( .A(n6038), .B(n6039), .Z(n6024) );
  NANDN U6019 ( .A(n6022), .B(n5178), .Z(n6039) );
  XOR U6020 ( .A(n6040), .B(n6041), .Z(n6038) );
  XNOR U6021 ( .A(n6042), .B(n6043), .Z(n6041) );
  NAND U6022 ( .A(n6044), .B(n6045), .Z(n4926) );
  OR U6023 ( .A(n5159), .B(n6046), .Z(n6045) );
  ANDN U6024 ( .B(n6047), .A(n5064), .Z(n6044) );
  AND U6025 ( .A(x[37]), .B(n4967), .Z(n5064) );
  NANDN U6026 ( .A(n5066), .B(n5162), .Z(n6047) );
  AND U6027 ( .A(n6048), .B(n6049), .Z(n5066) );
  AND U6028 ( .A(n6050), .B(n6051), .Z(n6049) );
  NAND U6029 ( .A(n6052), .B(n5168), .Z(n6051) );
  XOR U6030 ( .A(n6053), .B(n6054), .Z(n6052) );
  XNOR U6031 ( .A(n6055), .B(n6056), .Z(n6054) );
  AND U6032 ( .A(n6057), .B(n6058), .Z(n6050) );
  NANDN U6033 ( .A(n6046), .B(n6059), .Z(n6058) );
  NOR U6034 ( .A(n6060), .B(n5173), .Z(n6059) );
  NAND U6035 ( .A(n6061), .B(n5175), .Z(n6057) );
  NANDN U6036 ( .A(\stack[0][37] ), .B(n6060), .Z(n6061) );
  AND U6037 ( .A(n6062), .B(n6063), .Z(n6048) );
  NANDN U6038 ( .A(n6046), .B(n5178), .Z(n6063) );
  XOR U6039 ( .A(n6064), .B(n6065), .Z(n6062) );
  XNOR U6040 ( .A(n6066), .B(n6067), .Z(n6065) );
  NAND U6041 ( .A(n6068), .B(n6069), .Z(n4925) );
  OR U6042 ( .A(n5159), .B(n6070), .Z(n6069) );
  ANDN U6043 ( .B(n6071), .A(n5061), .Z(n6068) );
  AND U6044 ( .A(x[38]), .B(n4967), .Z(n5061) );
  NANDN U6045 ( .A(n5063), .B(n5162), .Z(n6071) );
  AND U6046 ( .A(n6072), .B(n6073), .Z(n5063) );
  AND U6047 ( .A(n6074), .B(n6075), .Z(n6073) );
  NAND U6048 ( .A(n6076), .B(n5168), .Z(n6075) );
  XOR U6049 ( .A(n6077), .B(n6078), .Z(n6076) );
  XNOR U6050 ( .A(n6079), .B(n6080), .Z(n6078) );
  AND U6051 ( .A(n6081), .B(n6082), .Z(n6074) );
  NANDN U6052 ( .A(n6070), .B(n6083), .Z(n6082) );
  NOR U6053 ( .A(n6084), .B(n5173), .Z(n6083) );
  NAND U6054 ( .A(n6085), .B(n5175), .Z(n6081) );
  NANDN U6055 ( .A(\stack[0][38] ), .B(n6084), .Z(n6085) );
  AND U6056 ( .A(n6086), .B(n6087), .Z(n6072) );
  NANDN U6057 ( .A(n6070), .B(n5178), .Z(n6087) );
  XOR U6058 ( .A(n6088), .B(n6089), .Z(n6086) );
  XNOR U6059 ( .A(n6090), .B(n6091), .Z(n6089) );
  NAND U6060 ( .A(n6092), .B(n6093), .Z(n4924) );
  OR U6061 ( .A(n5159), .B(n6094), .Z(n6093) );
  ANDN U6062 ( .B(n6095), .A(n5058), .Z(n6092) );
  AND U6063 ( .A(x[39]), .B(n4967), .Z(n5058) );
  NANDN U6064 ( .A(n5060), .B(n5162), .Z(n6095) );
  AND U6065 ( .A(n6096), .B(n6097), .Z(n5060) );
  AND U6066 ( .A(n6098), .B(n6099), .Z(n6097) );
  NAND U6067 ( .A(n6100), .B(n5168), .Z(n6099) );
  XOR U6068 ( .A(n6101), .B(n6102), .Z(n6100) );
  XNOR U6069 ( .A(n6103), .B(n6104), .Z(n6102) );
  AND U6070 ( .A(n6105), .B(n6106), .Z(n6098) );
  NANDN U6071 ( .A(n6094), .B(n6107), .Z(n6106) );
  NOR U6072 ( .A(n6108), .B(n5173), .Z(n6107) );
  NAND U6073 ( .A(n6109), .B(n5175), .Z(n6105) );
  NANDN U6074 ( .A(\stack[0][39] ), .B(n6108), .Z(n6109) );
  AND U6075 ( .A(n6110), .B(n6111), .Z(n6096) );
  NANDN U6076 ( .A(n6094), .B(n5178), .Z(n6111) );
  XOR U6077 ( .A(n6112), .B(n6113), .Z(n6110) );
  XNOR U6078 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U6079 ( .A(n6116), .B(n6117), .Z(n4923) );
  OR U6080 ( .A(n5159), .B(n6118), .Z(n6117) );
  ANDN U6081 ( .B(n6119), .A(n5052), .Z(n6116) );
  AND U6082 ( .A(x[40]), .B(n4967), .Z(n5052) );
  NANDN U6083 ( .A(n5054), .B(n5162), .Z(n6119) );
  AND U6084 ( .A(n6120), .B(n6121), .Z(n5054) );
  AND U6085 ( .A(n6122), .B(n6123), .Z(n6121) );
  NAND U6086 ( .A(n6124), .B(n5168), .Z(n6123) );
  XOR U6087 ( .A(n6125), .B(n6126), .Z(n6124) );
  XNOR U6088 ( .A(n6127), .B(n6128), .Z(n6126) );
  AND U6089 ( .A(n6129), .B(n6130), .Z(n6122) );
  NANDN U6090 ( .A(n6118), .B(n6131), .Z(n6130) );
  NOR U6091 ( .A(n6132), .B(n5173), .Z(n6131) );
  NAND U6092 ( .A(n6133), .B(n5175), .Z(n6129) );
  NANDN U6093 ( .A(\stack[0][40] ), .B(n6132), .Z(n6133) );
  AND U6094 ( .A(n6134), .B(n6135), .Z(n6120) );
  NANDN U6095 ( .A(n6118), .B(n5178), .Z(n6135) );
  XOR U6096 ( .A(n6136), .B(n6137), .Z(n6134) );
  XNOR U6097 ( .A(n6138), .B(n6139), .Z(n6137) );
  NAND U6098 ( .A(n6140), .B(n6141), .Z(n4922) );
  OR U6099 ( .A(n5159), .B(n6142), .Z(n6141) );
  ANDN U6100 ( .B(n6143), .A(n5049), .Z(n6140) );
  AND U6101 ( .A(x[41]), .B(n4967), .Z(n5049) );
  NANDN U6102 ( .A(n5051), .B(n5162), .Z(n6143) );
  AND U6103 ( .A(n6144), .B(n6145), .Z(n5051) );
  AND U6104 ( .A(n6146), .B(n6147), .Z(n6145) );
  NAND U6105 ( .A(n6148), .B(n5168), .Z(n6147) );
  XOR U6106 ( .A(n6149), .B(n6150), .Z(n6148) );
  XNOR U6107 ( .A(n6151), .B(n6152), .Z(n6150) );
  AND U6108 ( .A(n6153), .B(n6154), .Z(n6146) );
  NANDN U6109 ( .A(n6142), .B(n6155), .Z(n6154) );
  NOR U6110 ( .A(n6156), .B(n5173), .Z(n6155) );
  NAND U6111 ( .A(n6157), .B(n5175), .Z(n6153) );
  NANDN U6112 ( .A(\stack[0][41] ), .B(n6156), .Z(n6157) );
  AND U6113 ( .A(n6158), .B(n6159), .Z(n6144) );
  NANDN U6114 ( .A(n6142), .B(n5178), .Z(n6159) );
  XOR U6115 ( .A(n6160), .B(n6161), .Z(n6158) );
  XNOR U6116 ( .A(n6162), .B(n6163), .Z(n6161) );
  NAND U6117 ( .A(n6164), .B(n6165), .Z(n4921) );
  OR U6118 ( .A(n5159), .B(n6166), .Z(n6165) );
  ANDN U6119 ( .B(n6167), .A(n5046), .Z(n6164) );
  AND U6120 ( .A(x[42]), .B(n4967), .Z(n5046) );
  NANDN U6121 ( .A(n5048), .B(n5162), .Z(n6167) );
  AND U6122 ( .A(n6168), .B(n6169), .Z(n5048) );
  AND U6123 ( .A(n6170), .B(n6171), .Z(n6169) );
  NAND U6124 ( .A(n6172), .B(n5168), .Z(n6171) );
  XOR U6125 ( .A(n6173), .B(n6174), .Z(n6172) );
  XNOR U6126 ( .A(n6175), .B(n6176), .Z(n6174) );
  AND U6127 ( .A(n6177), .B(n6178), .Z(n6170) );
  NANDN U6128 ( .A(n6166), .B(n6179), .Z(n6178) );
  NOR U6129 ( .A(n6180), .B(n5173), .Z(n6179) );
  NAND U6130 ( .A(n6181), .B(n5175), .Z(n6177) );
  NANDN U6131 ( .A(\stack[0][42] ), .B(n6180), .Z(n6181) );
  AND U6132 ( .A(n6182), .B(n6183), .Z(n6168) );
  NANDN U6133 ( .A(n6166), .B(n5178), .Z(n6183) );
  XOR U6134 ( .A(n6184), .B(n6185), .Z(n6182) );
  XNOR U6135 ( .A(n6186), .B(n6187), .Z(n6185) );
  NAND U6136 ( .A(n6188), .B(n6189), .Z(n4920) );
  OR U6137 ( .A(n5159), .B(n6190), .Z(n6189) );
  ANDN U6138 ( .B(n6191), .A(n5043), .Z(n6188) );
  AND U6139 ( .A(x[43]), .B(n4967), .Z(n5043) );
  NANDN U6140 ( .A(n5045), .B(n5162), .Z(n6191) );
  AND U6141 ( .A(n6192), .B(n6193), .Z(n5045) );
  AND U6142 ( .A(n6194), .B(n6195), .Z(n6193) );
  NAND U6143 ( .A(n6196), .B(n5168), .Z(n6195) );
  XOR U6144 ( .A(n6197), .B(n6198), .Z(n6196) );
  XNOR U6145 ( .A(n6199), .B(n6200), .Z(n6198) );
  AND U6146 ( .A(n6201), .B(n6202), .Z(n6194) );
  NANDN U6147 ( .A(n6190), .B(n6203), .Z(n6202) );
  NOR U6148 ( .A(n6204), .B(n5173), .Z(n6203) );
  NAND U6149 ( .A(n6205), .B(n5175), .Z(n6201) );
  NANDN U6150 ( .A(\stack[0][43] ), .B(n6204), .Z(n6205) );
  AND U6151 ( .A(n6206), .B(n6207), .Z(n6192) );
  NANDN U6152 ( .A(n6190), .B(n5178), .Z(n6207) );
  XOR U6153 ( .A(n6208), .B(n6209), .Z(n6206) );
  XNOR U6154 ( .A(n6210), .B(n6211), .Z(n6209) );
  NAND U6155 ( .A(n6212), .B(n6213), .Z(n4919) );
  OR U6156 ( .A(n5159), .B(n6214), .Z(n6213) );
  ANDN U6157 ( .B(n6215), .A(n5040), .Z(n6212) );
  AND U6158 ( .A(x[44]), .B(n4967), .Z(n5040) );
  NANDN U6159 ( .A(n5042), .B(n5162), .Z(n6215) );
  AND U6160 ( .A(n6216), .B(n6217), .Z(n5042) );
  AND U6161 ( .A(n6218), .B(n6219), .Z(n6217) );
  NAND U6162 ( .A(n6220), .B(n5168), .Z(n6219) );
  XOR U6163 ( .A(n6221), .B(n6222), .Z(n6220) );
  XNOR U6164 ( .A(n6223), .B(n6224), .Z(n6222) );
  AND U6165 ( .A(n6225), .B(n6226), .Z(n6218) );
  NANDN U6166 ( .A(n6214), .B(n6227), .Z(n6226) );
  NOR U6167 ( .A(n6228), .B(n5173), .Z(n6227) );
  NAND U6168 ( .A(n6229), .B(n5175), .Z(n6225) );
  NANDN U6169 ( .A(\stack[0][44] ), .B(n6228), .Z(n6229) );
  AND U6170 ( .A(n6230), .B(n6231), .Z(n6216) );
  NANDN U6171 ( .A(n6214), .B(n5178), .Z(n6231) );
  XOR U6172 ( .A(n6232), .B(n6233), .Z(n6230) );
  XNOR U6173 ( .A(n6234), .B(n6235), .Z(n6233) );
  NAND U6174 ( .A(n6236), .B(n6237), .Z(n4918) );
  OR U6175 ( .A(n5159), .B(n6238), .Z(n6237) );
  ANDN U6176 ( .B(n6239), .A(n5037), .Z(n6236) );
  AND U6177 ( .A(x[45]), .B(n4967), .Z(n5037) );
  NANDN U6178 ( .A(n5039), .B(n5162), .Z(n6239) );
  AND U6179 ( .A(n6240), .B(n6241), .Z(n5039) );
  AND U6180 ( .A(n6242), .B(n6243), .Z(n6241) );
  NAND U6181 ( .A(n6244), .B(n5168), .Z(n6243) );
  XOR U6182 ( .A(n6245), .B(n6246), .Z(n6244) );
  XNOR U6183 ( .A(n6247), .B(n6248), .Z(n6246) );
  AND U6184 ( .A(n6249), .B(n6250), .Z(n6242) );
  NANDN U6185 ( .A(n6238), .B(n6251), .Z(n6250) );
  NOR U6186 ( .A(n6252), .B(n5173), .Z(n6251) );
  NAND U6187 ( .A(n6253), .B(n5175), .Z(n6249) );
  NANDN U6188 ( .A(\stack[0][45] ), .B(n6252), .Z(n6253) );
  AND U6189 ( .A(n6254), .B(n6255), .Z(n6240) );
  NANDN U6190 ( .A(n6238), .B(n5178), .Z(n6255) );
  XOR U6191 ( .A(n6256), .B(n6257), .Z(n6254) );
  XNOR U6192 ( .A(n6258), .B(n6259), .Z(n6257) );
  NAND U6193 ( .A(n6260), .B(n6261), .Z(n4917) );
  OR U6194 ( .A(n5159), .B(n6262), .Z(n6261) );
  ANDN U6195 ( .B(n6263), .A(n5034), .Z(n6260) );
  AND U6196 ( .A(x[46]), .B(n4967), .Z(n5034) );
  NANDN U6197 ( .A(n5036), .B(n5162), .Z(n6263) );
  AND U6198 ( .A(n6264), .B(n6265), .Z(n5036) );
  AND U6199 ( .A(n6266), .B(n6267), .Z(n6265) );
  NAND U6200 ( .A(n6268), .B(n5168), .Z(n6267) );
  XOR U6201 ( .A(n6269), .B(n6270), .Z(n6268) );
  XNOR U6202 ( .A(n6271), .B(n6272), .Z(n6270) );
  AND U6203 ( .A(n6273), .B(n6274), .Z(n6266) );
  NANDN U6204 ( .A(n6262), .B(n6275), .Z(n6274) );
  NOR U6205 ( .A(n6276), .B(n5173), .Z(n6275) );
  NAND U6206 ( .A(n6277), .B(n5175), .Z(n6273) );
  NANDN U6207 ( .A(\stack[0][46] ), .B(n6276), .Z(n6277) );
  AND U6208 ( .A(n6278), .B(n6279), .Z(n6264) );
  NANDN U6209 ( .A(n6262), .B(n5178), .Z(n6279) );
  XOR U6210 ( .A(n6280), .B(n6281), .Z(n6278) );
  XNOR U6211 ( .A(n6282), .B(n6283), .Z(n6281) );
  NAND U6212 ( .A(n6284), .B(n6285), .Z(n4916) );
  OR U6213 ( .A(n5159), .B(n6286), .Z(n6285) );
  ANDN U6214 ( .B(n6287), .A(n5031), .Z(n6284) );
  AND U6215 ( .A(x[47]), .B(n4967), .Z(n5031) );
  NANDN U6216 ( .A(n5033), .B(n5162), .Z(n6287) );
  AND U6217 ( .A(n6288), .B(n6289), .Z(n5033) );
  AND U6218 ( .A(n6290), .B(n6291), .Z(n6289) );
  NAND U6219 ( .A(n6292), .B(n5168), .Z(n6291) );
  XOR U6220 ( .A(n6293), .B(n6294), .Z(n6292) );
  XNOR U6221 ( .A(n6295), .B(n6296), .Z(n6294) );
  AND U6222 ( .A(n6297), .B(n6298), .Z(n6290) );
  NANDN U6223 ( .A(n6286), .B(n6299), .Z(n6298) );
  NOR U6224 ( .A(n6300), .B(n5173), .Z(n6299) );
  NAND U6225 ( .A(n6301), .B(n5175), .Z(n6297) );
  NANDN U6226 ( .A(\stack[0][47] ), .B(n6300), .Z(n6301) );
  AND U6227 ( .A(n6302), .B(n6303), .Z(n6288) );
  NANDN U6228 ( .A(n6286), .B(n5178), .Z(n6303) );
  XOR U6229 ( .A(n6304), .B(n6305), .Z(n6302) );
  XNOR U6230 ( .A(n6306), .B(n6307), .Z(n6305) );
  NAND U6231 ( .A(n6308), .B(n6309), .Z(n4915) );
  OR U6232 ( .A(n5159), .B(n6310), .Z(n6309) );
  ANDN U6233 ( .B(n6311), .A(n5028), .Z(n6308) );
  AND U6234 ( .A(x[48]), .B(n4967), .Z(n5028) );
  NANDN U6235 ( .A(n5030), .B(n5162), .Z(n6311) );
  AND U6236 ( .A(n6312), .B(n6313), .Z(n5030) );
  AND U6237 ( .A(n6314), .B(n6315), .Z(n6313) );
  NAND U6238 ( .A(n6316), .B(n5168), .Z(n6315) );
  XOR U6239 ( .A(n6317), .B(n6318), .Z(n6316) );
  XNOR U6240 ( .A(n6319), .B(n6320), .Z(n6318) );
  AND U6241 ( .A(n6321), .B(n6322), .Z(n6314) );
  NANDN U6242 ( .A(n6310), .B(n6323), .Z(n6322) );
  NOR U6243 ( .A(n6324), .B(n5173), .Z(n6323) );
  NAND U6244 ( .A(n6325), .B(n5175), .Z(n6321) );
  NANDN U6245 ( .A(\stack[0][48] ), .B(n6324), .Z(n6325) );
  AND U6246 ( .A(n6326), .B(n6327), .Z(n6312) );
  NANDN U6247 ( .A(n6310), .B(n5178), .Z(n6327) );
  XOR U6248 ( .A(n6328), .B(n6329), .Z(n6326) );
  XNOR U6249 ( .A(n6330), .B(n6331), .Z(n6329) );
  NAND U6250 ( .A(n6332), .B(n6333), .Z(n4914) );
  OR U6251 ( .A(n5159), .B(n6334), .Z(n6333) );
  ANDN U6252 ( .B(n6335), .A(n5025), .Z(n6332) );
  AND U6253 ( .A(x[49]), .B(n4967), .Z(n5025) );
  NANDN U6254 ( .A(n5027), .B(n5162), .Z(n6335) );
  AND U6255 ( .A(n6336), .B(n6337), .Z(n5027) );
  AND U6256 ( .A(n6338), .B(n6339), .Z(n6337) );
  NAND U6257 ( .A(n6340), .B(n5168), .Z(n6339) );
  XOR U6258 ( .A(n6341), .B(n6342), .Z(n6340) );
  XNOR U6259 ( .A(n6343), .B(n6344), .Z(n6342) );
  AND U6260 ( .A(n6345), .B(n6346), .Z(n6338) );
  NANDN U6261 ( .A(n6334), .B(n6347), .Z(n6346) );
  NOR U6262 ( .A(n6348), .B(n5173), .Z(n6347) );
  NAND U6263 ( .A(n6349), .B(n5175), .Z(n6345) );
  NANDN U6264 ( .A(\stack[0][49] ), .B(n6348), .Z(n6349) );
  AND U6265 ( .A(n6350), .B(n6351), .Z(n6336) );
  NANDN U6266 ( .A(n6334), .B(n5178), .Z(n6351) );
  XOR U6267 ( .A(n6352), .B(n6353), .Z(n6350) );
  XNOR U6268 ( .A(n6354), .B(n6355), .Z(n6353) );
  NAND U6269 ( .A(n6356), .B(n6357), .Z(n4913) );
  OR U6270 ( .A(n5159), .B(n6358), .Z(n6357) );
  ANDN U6271 ( .B(n6359), .A(n5019), .Z(n6356) );
  AND U6272 ( .A(x[50]), .B(n4967), .Z(n5019) );
  NANDN U6273 ( .A(n5021), .B(n5162), .Z(n6359) );
  AND U6274 ( .A(n6360), .B(n6361), .Z(n5021) );
  AND U6275 ( .A(n6362), .B(n6363), .Z(n6361) );
  NAND U6276 ( .A(n6364), .B(n5168), .Z(n6363) );
  XOR U6277 ( .A(n6365), .B(n6366), .Z(n6364) );
  XNOR U6278 ( .A(n6367), .B(n6368), .Z(n6366) );
  AND U6279 ( .A(n6369), .B(n6370), .Z(n6362) );
  NANDN U6280 ( .A(n6358), .B(n6371), .Z(n6370) );
  NOR U6281 ( .A(n6372), .B(n5173), .Z(n6371) );
  NAND U6282 ( .A(n6373), .B(n5175), .Z(n6369) );
  NANDN U6283 ( .A(\stack[0][50] ), .B(n6372), .Z(n6373) );
  AND U6284 ( .A(n6374), .B(n6375), .Z(n6360) );
  NANDN U6285 ( .A(n6358), .B(n5178), .Z(n6375) );
  XOR U6286 ( .A(n6376), .B(n6377), .Z(n6374) );
  XNOR U6287 ( .A(n6378), .B(n6379), .Z(n6377) );
  NAND U6288 ( .A(n6380), .B(n6381), .Z(n4912) );
  OR U6289 ( .A(n5159), .B(n6382), .Z(n6381) );
  ANDN U6290 ( .B(n6383), .A(n5016), .Z(n6380) );
  AND U6291 ( .A(x[51]), .B(n4967), .Z(n5016) );
  NANDN U6292 ( .A(n5018), .B(n5162), .Z(n6383) );
  AND U6293 ( .A(n6384), .B(n6385), .Z(n5018) );
  AND U6294 ( .A(n6386), .B(n6387), .Z(n6385) );
  NAND U6295 ( .A(n6388), .B(n5168), .Z(n6387) );
  XOR U6296 ( .A(n6389), .B(n6390), .Z(n6388) );
  XNOR U6297 ( .A(n6391), .B(n6392), .Z(n6390) );
  AND U6298 ( .A(n6393), .B(n6394), .Z(n6386) );
  NANDN U6299 ( .A(n6382), .B(n6395), .Z(n6394) );
  NOR U6300 ( .A(n6396), .B(n5173), .Z(n6395) );
  NAND U6301 ( .A(n6397), .B(n5175), .Z(n6393) );
  NANDN U6302 ( .A(\stack[0][51] ), .B(n6396), .Z(n6397) );
  AND U6303 ( .A(n6398), .B(n6399), .Z(n6384) );
  NANDN U6304 ( .A(n6382), .B(n5178), .Z(n6399) );
  XOR U6305 ( .A(n6400), .B(n6401), .Z(n6398) );
  XNOR U6306 ( .A(n6402), .B(n6403), .Z(n6401) );
  NAND U6307 ( .A(n6404), .B(n6405), .Z(n4911) );
  OR U6308 ( .A(n5159), .B(n6406), .Z(n6405) );
  ANDN U6309 ( .B(n6407), .A(n5013), .Z(n6404) );
  AND U6310 ( .A(x[52]), .B(n4967), .Z(n5013) );
  NANDN U6311 ( .A(n5015), .B(n5162), .Z(n6407) );
  AND U6312 ( .A(n6408), .B(n6409), .Z(n5015) );
  AND U6313 ( .A(n6410), .B(n6411), .Z(n6409) );
  NAND U6314 ( .A(n6412), .B(n5168), .Z(n6411) );
  XOR U6315 ( .A(n6413), .B(n6414), .Z(n6412) );
  XNOR U6316 ( .A(n6415), .B(n6416), .Z(n6414) );
  AND U6317 ( .A(n6417), .B(n6418), .Z(n6410) );
  NANDN U6318 ( .A(n6406), .B(n6419), .Z(n6418) );
  NOR U6319 ( .A(n6420), .B(n5173), .Z(n6419) );
  NAND U6320 ( .A(n6421), .B(n5175), .Z(n6417) );
  NANDN U6321 ( .A(\stack[0][52] ), .B(n6420), .Z(n6421) );
  AND U6322 ( .A(n6422), .B(n6423), .Z(n6408) );
  NANDN U6323 ( .A(n6406), .B(n5178), .Z(n6423) );
  XOR U6324 ( .A(n6424), .B(n6425), .Z(n6422) );
  XNOR U6325 ( .A(n6426), .B(n6427), .Z(n6425) );
  NAND U6326 ( .A(n6428), .B(n6429), .Z(n4910) );
  OR U6327 ( .A(n5159), .B(n6430), .Z(n6429) );
  ANDN U6328 ( .B(n6431), .A(n5010), .Z(n6428) );
  AND U6329 ( .A(x[53]), .B(n4967), .Z(n5010) );
  NANDN U6330 ( .A(n5012), .B(n5162), .Z(n6431) );
  AND U6331 ( .A(n6432), .B(n6433), .Z(n5012) );
  AND U6332 ( .A(n6434), .B(n6435), .Z(n6433) );
  NAND U6333 ( .A(n6436), .B(n5168), .Z(n6435) );
  XOR U6334 ( .A(n6437), .B(n6438), .Z(n6436) );
  XNOR U6335 ( .A(n6439), .B(n6440), .Z(n6438) );
  AND U6336 ( .A(n6441), .B(n6442), .Z(n6434) );
  NANDN U6337 ( .A(n6430), .B(n6443), .Z(n6442) );
  NOR U6338 ( .A(n6444), .B(n5173), .Z(n6443) );
  NAND U6339 ( .A(n6445), .B(n5175), .Z(n6441) );
  NANDN U6340 ( .A(\stack[0][53] ), .B(n6444), .Z(n6445) );
  AND U6341 ( .A(n6446), .B(n6447), .Z(n6432) );
  NANDN U6342 ( .A(n6430), .B(n5178), .Z(n6447) );
  XOR U6343 ( .A(n6448), .B(n6449), .Z(n6446) );
  XNOR U6344 ( .A(n6450), .B(n6451), .Z(n6449) );
  NAND U6345 ( .A(n6452), .B(n6453), .Z(n4909) );
  OR U6346 ( .A(n5159), .B(n6454), .Z(n6453) );
  ANDN U6347 ( .B(n6455), .A(n5007), .Z(n6452) );
  AND U6348 ( .A(x[54]), .B(n4967), .Z(n5007) );
  NANDN U6349 ( .A(n5009), .B(n5162), .Z(n6455) );
  AND U6350 ( .A(n6456), .B(n6457), .Z(n5009) );
  AND U6351 ( .A(n6458), .B(n6459), .Z(n6457) );
  NAND U6352 ( .A(n6460), .B(n5168), .Z(n6459) );
  XOR U6353 ( .A(n6461), .B(n6462), .Z(n6460) );
  XNOR U6354 ( .A(n6463), .B(n6464), .Z(n6462) );
  AND U6355 ( .A(n6465), .B(n6466), .Z(n6458) );
  NANDN U6356 ( .A(n6454), .B(n6467), .Z(n6466) );
  NOR U6357 ( .A(n6468), .B(n5173), .Z(n6467) );
  NAND U6358 ( .A(n6469), .B(n5175), .Z(n6465) );
  NANDN U6359 ( .A(\stack[0][54] ), .B(n6468), .Z(n6469) );
  AND U6360 ( .A(n6470), .B(n6471), .Z(n6456) );
  NANDN U6361 ( .A(n6454), .B(n5178), .Z(n6471) );
  XOR U6362 ( .A(n6472), .B(n6473), .Z(n6470) );
  XNOR U6363 ( .A(n6474), .B(n6475), .Z(n6473) );
  NAND U6364 ( .A(n6476), .B(n6477), .Z(n4908) );
  OR U6365 ( .A(n5159), .B(n6478), .Z(n6477) );
  ANDN U6366 ( .B(n6479), .A(n5004), .Z(n6476) );
  AND U6367 ( .A(x[55]), .B(n4967), .Z(n5004) );
  NANDN U6368 ( .A(n5006), .B(n5162), .Z(n6479) );
  AND U6369 ( .A(n6480), .B(n6481), .Z(n5006) );
  AND U6370 ( .A(n6482), .B(n6483), .Z(n6481) );
  NAND U6371 ( .A(n6484), .B(n5168), .Z(n6483) );
  XOR U6372 ( .A(n6485), .B(n6486), .Z(n6484) );
  XNOR U6373 ( .A(n6487), .B(n6488), .Z(n6486) );
  AND U6374 ( .A(n6489), .B(n6490), .Z(n6482) );
  NANDN U6375 ( .A(n6478), .B(n6491), .Z(n6490) );
  NOR U6376 ( .A(n6492), .B(n5173), .Z(n6491) );
  NAND U6377 ( .A(n6493), .B(n5175), .Z(n6489) );
  NANDN U6378 ( .A(\stack[0][55] ), .B(n6492), .Z(n6493) );
  AND U6379 ( .A(n6494), .B(n6495), .Z(n6480) );
  NANDN U6380 ( .A(n6478), .B(n5178), .Z(n6495) );
  XOR U6381 ( .A(n6496), .B(n6497), .Z(n6494) );
  XNOR U6382 ( .A(n6498), .B(n6499), .Z(n6497) );
  NAND U6383 ( .A(n6500), .B(n6501), .Z(n4907) );
  OR U6384 ( .A(n5159), .B(n6502), .Z(n6501) );
  ANDN U6385 ( .B(n6503), .A(n5001), .Z(n6500) );
  AND U6386 ( .A(x[56]), .B(n4967), .Z(n5001) );
  NANDN U6387 ( .A(n5003), .B(n5162), .Z(n6503) );
  AND U6388 ( .A(n6504), .B(n6505), .Z(n5003) );
  AND U6389 ( .A(n6506), .B(n6507), .Z(n6505) );
  NAND U6390 ( .A(n6508), .B(n5168), .Z(n6507) );
  XOR U6391 ( .A(n6509), .B(n6510), .Z(n6508) );
  XNOR U6392 ( .A(n6511), .B(n6512), .Z(n6510) );
  AND U6393 ( .A(n6513), .B(n6514), .Z(n6506) );
  NANDN U6394 ( .A(n6502), .B(n6515), .Z(n6514) );
  NOR U6395 ( .A(n6516), .B(n5173), .Z(n6515) );
  NAND U6396 ( .A(n6517), .B(n5175), .Z(n6513) );
  NANDN U6397 ( .A(\stack[0][56] ), .B(n6516), .Z(n6517) );
  AND U6398 ( .A(n6518), .B(n6519), .Z(n6504) );
  NANDN U6399 ( .A(n6502), .B(n5178), .Z(n6519) );
  XOR U6400 ( .A(n6520), .B(n6521), .Z(n6518) );
  XNOR U6401 ( .A(n6522), .B(n6523), .Z(n6521) );
  NAND U6402 ( .A(n6524), .B(n6525), .Z(n4906) );
  OR U6403 ( .A(n5159), .B(n6526), .Z(n6525) );
  ANDN U6404 ( .B(n6527), .A(n4998), .Z(n6524) );
  AND U6405 ( .A(x[57]), .B(n4967), .Z(n4998) );
  NANDN U6406 ( .A(n5000), .B(n5162), .Z(n6527) );
  AND U6407 ( .A(n6528), .B(n6529), .Z(n5000) );
  AND U6408 ( .A(n6530), .B(n6531), .Z(n6529) );
  NAND U6409 ( .A(n6532), .B(n5168), .Z(n6531) );
  XOR U6410 ( .A(n6533), .B(n6534), .Z(n6532) );
  XNOR U6411 ( .A(n6535), .B(n6536), .Z(n6534) );
  AND U6412 ( .A(n6537), .B(n6538), .Z(n6530) );
  NANDN U6413 ( .A(n6526), .B(n6539), .Z(n6538) );
  NOR U6414 ( .A(n6540), .B(n5173), .Z(n6539) );
  NAND U6415 ( .A(n6541), .B(n5175), .Z(n6537) );
  NANDN U6416 ( .A(\stack[0][57] ), .B(n6540), .Z(n6541) );
  AND U6417 ( .A(n6542), .B(n6543), .Z(n6528) );
  NANDN U6418 ( .A(n6526), .B(n5178), .Z(n6543) );
  XOR U6419 ( .A(n6544), .B(n6545), .Z(n6542) );
  XNOR U6420 ( .A(n6546), .B(n6547), .Z(n6545) );
  NAND U6421 ( .A(n6548), .B(n6549), .Z(n4905) );
  OR U6422 ( .A(n5159), .B(n6550), .Z(n6549) );
  ANDN U6423 ( .B(n6551), .A(n4995), .Z(n6548) );
  AND U6424 ( .A(x[58]), .B(n4967), .Z(n4995) );
  NANDN U6425 ( .A(n4997), .B(n5162), .Z(n6551) );
  AND U6426 ( .A(n6552), .B(n6553), .Z(n4997) );
  AND U6427 ( .A(n6554), .B(n6555), .Z(n6553) );
  NAND U6428 ( .A(n6556), .B(n5168), .Z(n6555) );
  XOR U6429 ( .A(n6557), .B(n6558), .Z(n6556) );
  XNOR U6430 ( .A(n6559), .B(n6560), .Z(n6558) );
  AND U6431 ( .A(n6561), .B(n6562), .Z(n6554) );
  NANDN U6432 ( .A(n6550), .B(n6563), .Z(n6562) );
  NOR U6433 ( .A(n6564), .B(n5173), .Z(n6563) );
  NAND U6434 ( .A(n6565), .B(n5175), .Z(n6561) );
  NANDN U6435 ( .A(\stack[0][58] ), .B(n6564), .Z(n6565) );
  AND U6436 ( .A(n6566), .B(n6567), .Z(n6552) );
  NANDN U6437 ( .A(n6550), .B(n5178), .Z(n6567) );
  XOR U6438 ( .A(n6568), .B(n6569), .Z(n6566) );
  XNOR U6439 ( .A(n6570), .B(n6571), .Z(n6569) );
  NAND U6440 ( .A(n6572), .B(n6573), .Z(n4904) );
  OR U6441 ( .A(n5159), .B(n6574), .Z(n6573) );
  ANDN U6442 ( .B(n6575), .A(n4992), .Z(n6572) );
  AND U6443 ( .A(x[59]), .B(n4967), .Z(n4992) );
  NANDN U6444 ( .A(n4994), .B(n5162), .Z(n6575) );
  AND U6445 ( .A(n6576), .B(n6577), .Z(n4994) );
  AND U6446 ( .A(n6578), .B(n6579), .Z(n6577) );
  NAND U6447 ( .A(n6580), .B(n5168), .Z(n6579) );
  XOR U6448 ( .A(n6581), .B(n6582), .Z(n6580) );
  XNOR U6449 ( .A(n6583), .B(n6584), .Z(n6582) );
  AND U6450 ( .A(n6585), .B(n6586), .Z(n6578) );
  NANDN U6451 ( .A(n6574), .B(n6587), .Z(n6586) );
  NOR U6452 ( .A(n6588), .B(n5173), .Z(n6587) );
  NAND U6453 ( .A(n6589), .B(n5175), .Z(n6585) );
  NANDN U6454 ( .A(\stack[0][59] ), .B(n6588), .Z(n6589) );
  AND U6455 ( .A(n6590), .B(n6591), .Z(n6576) );
  NANDN U6456 ( .A(n6574), .B(n5178), .Z(n6591) );
  XOR U6457 ( .A(n6592), .B(n6593), .Z(n6590) );
  XNOR U6458 ( .A(n6594), .B(n6595), .Z(n6593) );
  NAND U6459 ( .A(n6596), .B(n6597), .Z(n4903) );
  OR U6460 ( .A(n5159), .B(n6598), .Z(n6597) );
  ANDN U6461 ( .B(n6599), .A(n4986), .Z(n6596) );
  AND U6462 ( .A(x[60]), .B(n4967), .Z(n4986) );
  NANDN U6463 ( .A(n4988), .B(n5162), .Z(n6599) );
  AND U6464 ( .A(n6600), .B(n6601), .Z(n4988) );
  AND U6465 ( .A(n6602), .B(n6603), .Z(n6601) );
  NAND U6466 ( .A(n6604), .B(n5168), .Z(n6603) );
  XOR U6467 ( .A(n6605), .B(n6606), .Z(n6604) );
  XNOR U6468 ( .A(n6607), .B(n6608), .Z(n6606) );
  AND U6469 ( .A(n6609), .B(n6610), .Z(n6602) );
  NANDN U6470 ( .A(n6598), .B(n6611), .Z(n6610) );
  NOR U6471 ( .A(n6612), .B(n5173), .Z(n6611) );
  NAND U6472 ( .A(n6613), .B(n5175), .Z(n6609) );
  NANDN U6473 ( .A(\stack[0][60] ), .B(n6612), .Z(n6613) );
  AND U6474 ( .A(n6614), .B(n6615), .Z(n6600) );
  NANDN U6475 ( .A(n6598), .B(n5178), .Z(n6615) );
  XOR U6476 ( .A(n6616), .B(n6617), .Z(n6614) );
  XNOR U6477 ( .A(n6618), .B(n6619), .Z(n6617) );
  NAND U6478 ( .A(n6620), .B(n6621), .Z(n4902) );
  OR U6479 ( .A(n5159), .B(n6622), .Z(n6621) );
  ANDN U6480 ( .B(n6623), .A(n4983), .Z(n6620) );
  AND U6481 ( .A(x[61]), .B(n4967), .Z(n4983) );
  NANDN U6482 ( .A(n4985), .B(n5162), .Z(n6623) );
  AND U6483 ( .A(n6624), .B(n6625), .Z(n4985) );
  AND U6484 ( .A(n6626), .B(n6627), .Z(n6625) );
  NAND U6485 ( .A(n6628), .B(n5168), .Z(n6627) );
  XOR U6486 ( .A(n6629), .B(n6630), .Z(n6628) );
  XNOR U6487 ( .A(n6631), .B(n6632), .Z(n6630) );
  AND U6488 ( .A(n6633), .B(n6634), .Z(n6626) );
  NANDN U6489 ( .A(n6622), .B(n6635), .Z(n6634) );
  NOR U6490 ( .A(n6636), .B(n5173), .Z(n6635) );
  NAND U6491 ( .A(n6637), .B(n5175), .Z(n6633) );
  NANDN U6492 ( .A(\stack[0][61] ), .B(n6636), .Z(n6637) );
  AND U6493 ( .A(n6638), .B(n6639), .Z(n6624) );
  NANDN U6494 ( .A(n6622), .B(n5178), .Z(n6639) );
  XOR U6495 ( .A(n6640), .B(n6641), .Z(n6638) );
  XNOR U6496 ( .A(n6642), .B(n6643), .Z(n6641) );
  NAND U6497 ( .A(n6644), .B(n6645), .Z(n4901) );
  OR U6498 ( .A(n5159), .B(n6646), .Z(n6645) );
  ANDN U6499 ( .B(n6647), .A(n4980), .Z(n6644) );
  AND U6500 ( .A(x[62]), .B(n4967), .Z(n4980) );
  NANDN U6501 ( .A(n4982), .B(n5162), .Z(n6647) );
  AND U6502 ( .A(n6648), .B(n6649), .Z(n4982) );
  AND U6503 ( .A(n6650), .B(n6651), .Z(n6649) );
  NAND U6504 ( .A(n6652), .B(n5168), .Z(n6651) );
  XOR U6505 ( .A(n6653), .B(n6654), .Z(n6652) );
  XNOR U6506 ( .A(n6655), .B(n6656), .Z(n6654) );
  AND U6507 ( .A(n6657), .B(n6658), .Z(n6650) );
  NANDN U6508 ( .A(n6659), .B(n6660), .Z(n6658) );
  NOR U6509 ( .A(n6646), .B(n5173), .Z(n6660) );
  NAND U6510 ( .A(n6661), .B(n5175), .Z(n6657) );
  NANDN U6511 ( .A(\stack[0][62] ), .B(n6659), .Z(n6661) );
  AND U6512 ( .A(n6662), .B(n6663), .Z(n6648) );
  NANDN U6513 ( .A(n6646), .B(n5178), .Z(n6663) );
  XOR U6514 ( .A(n6664), .B(n6665), .Z(n6662) );
  XOR U6515 ( .A(n6666), .B(n6667), .Z(n6665) );
  NAND U6516 ( .A(n6668), .B(n6669), .Z(n4900) );
  OR U6517 ( .A(n5159), .B(n6670), .Z(n6669) );
  NANDN U6518 ( .A(n6671), .B(n6672), .Z(n5159) );
  NOR U6519 ( .A(n4967), .B(n6673), .Z(n6672) );
  ANDN U6520 ( .B(n6674), .A(n4977), .Z(n6668) );
  AND U6521 ( .A(x[63]), .B(n4967), .Z(n4977) );
  NANDN U6522 ( .A(n4979), .B(n5162), .Z(n6674) );
  OR U6523 ( .A(n6673), .B(n6671), .Z(n5162) );
  AND U6524 ( .A(n6675), .B(n6676), .Z(n4979) );
  AND U6525 ( .A(n6677), .B(n6678), .Z(n6676) );
  NAND U6526 ( .A(n6679), .B(n5168), .Z(n6678) );
  AND U6527 ( .A(n6680), .B(n6681), .Z(n6679) );
  NANDN U6528 ( .A(n6682), .B(n6683), .Z(n6681) );
  XNOR U6529 ( .A(n6684), .B(n6670), .Z(n6683) );
  NAND U6530 ( .A(n6685), .B(n6682), .Z(n6680) );
  XNOR U6531 ( .A(n6686), .B(n6687), .Z(n6682) );
  XOR U6532 ( .A(n6688), .B(n6689), .Z(n6687) );
  NANDN U6533 ( .A(n5195), .B(\stack[0][62] ), .Z(n6689) );
  AND U6534 ( .A(n6690), .B(n6691), .Z(n6688) );
  NAND U6535 ( .A(n6692), .B(n6656), .Z(n6691) );
  NAND U6536 ( .A(n6693), .B(n6694), .Z(n6656) );
  NANDN U6537 ( .A(n6632), .B(n6695), .Z(n6694) );
  OR U6538 ( .A(n6631), .B(n6629), .Z(n6695) );
  AND U6539 ( .A(n6696), .B(n6697), .Z(n6632) );
  NAND U6540 ( .A(n6698), .B(n6608), .Z(n6696) );
  NAND U6541 ( .A(n6699), .B(n6700), .Z(n6608) );
  NANDN U6542 ( .A(n6584), .B(n6701), .Z(n6700) );
  OR U6543 ( .A(n6583), .B(n6581), .Z(n6701) );
  AND U6544 ( .A(n6702), .B(n6703), .Z(n6584) );
  NAND U6545 ( .A(n6704), .B(n6560), .Z(n6702) );
  NAND U6546 ( .A(n6705), .B(n6706), .Z(n6560) );
  NANDN U6547 ( .A(n6536), .B(n6707), .Z(n6706) );
  OR U6548 ( .A(n6535), .B(n6533), .Z(n6707) );
  AND U6549 ( .A(n6708), .B(n6709), .Z(n6536) );
  NAND U6550 ( .A(n6710), .B(n6512), .Z(n6708) );
  NAND U6551 ( .A(n6711), .B(n6712), .Z(n6512) );
  NANDN U6552 ( .A(n6488), .B(n6713), .Z(n6712) );
  OR U6553 ( .A(n6487), .B(n6485), .Z(n6713) );
  AND U6554 ( .A(n6714), .B(n6715), .Z(n6488) );
  NAND U6555 ( .A(n6716), .B(n6464), .Z(n6714) );
  NAND U6556 ( .A(n6717), .B(n6718), .Z(n6464) );
  NANDN U6557 ( .A(n6440), .B(n6719), .Z(n6718) );
  OR U6558 ( .A(n6439), .B(n6437), .Z(n6719) );
  AND U6559 ( .A(n6720), .B(n6721), .Z(n6440) );
  NAND U6560 ( .A(n6722), .B(n6416), .Z(n6720) );
  NAND U6561 ( .A(n6723), .B(n6724), .Z(n6416) );
  NANDN U6562 ( .A(n6392), .B(n6725), .Z(n6724) );
  OR U6563 ( .A(n6391), .B(n6389), .Z(n6725) );
  AND U6564 ( .A(n6726), .B(n6727), .Z(n6392) );
  NAND U6565 ( .A(n6728), .B(n6368), .Z(n6726) );
  NAND U6566 ( .A(n6729), .B(n6730), .Z(n6368) );
  NANDN U6567 ( .A(n6344), .B(n6731), .Z(n6730) );
  OR U6568 ( .A(n6343), .B(n6341), .Z(n6731) );
  AND U6569 ( .A(n6732), .B(n6733), .Z(n6344) );
  NAND U6570 ( .A(n6734), .B(n6320), .Z(n6732) );
  NAND U6571 ( .A(n6735), .B(n6736), .Z(n6320) );
  NANDN U6572 ( .A(n6296), .B(n6737), .Z(n6736) );
  OR U6573 ( .A(n6295), .B(n6293), .Z(n6737) );
  AND U6574 ( .A(n6738), .B(n6739), .Z(n6296) );
  NAND U6575 ( .A(n6740), .B(n6272), .Z(n6738) );
  NAND U6576 ( .A(n6741), .B(n6742), .Z(n6272) );
  NANDN U6577 ( .A(n6248), .B(n6743), .Z(n6742) );
  OR U6578 ( .A(n6247), .B(n6245), .Z(n6743) );
  AND U6579 ( .A(n6744), .B(n6745), .Z(n6248) );
  NAND U6580 ( .A(n6746), .B(n6224), .Z(n6744) );
  NAND U6581 ( .A(n6747), .B(n6748), .Z(n6224) );
  NANDN U6582 ( .A(n6200), .B(n6749), .Z(n6748) );
  OR U6583 ( .A(n6199), .B(n6197), .Z(n6749) );
  AND U6584 ( .A(n6750), .B(n6751), .Z(n6200) );
  NAND U6585 ( .A(n6752), .B(n6176), .Z(n6750) );
  NAND U6586 ( .A(n6753), .B(n6754), .Z(n6176) );
  NANDN U6587 ( .A(n6152), .B(n6755), .Z(n6754) );
  OR U6588 ( .A(n6151), .B(n6149), .Z(n6755) );
  AND U6589 ( .A(n6756), .B(n6757), .Z(n6152) );
  NAND U6590 ( .A(n6758), .B(n6128), .Z(n6756) );
  NAND U6591 ( .A(n6759), .B(n6760), .Z(n6128) );
  NANDN U6592 ( .A(n6104), .B(n6761), .Z(n6760) );
  OR U6593 ( .A(n6103), .B(n6101), .Z(n6761) );
  AND U6594 ( .A(n6762), .B(n6763), .Z(n6104) );
  NAND U6595 ( .A(n6764), .B(n6080), .Z(n6762) );
  NAND U6596 ( .A(n6765), .B(n6766), .Z(n6080) );
  NANDN U6597 ( .A(n6056), .B(n6767), .Z(n6766) );
  OR U6598 ( .A(n6055), .B(n6053), .Z(n6767) );
  AND U6599 ( .A(n6768), .B(n6769), .Z(n6056) );
  NAND U6600 ( .A(n6770), .B(n6032), .Z(n6768) );
  NAND U6601 ( .A(n6771), .B(n6772), .Z(n6032) );
  NANDN U6602 ( .A(n6008), .B(n6773), .Z(n6772) );
  OR U6603 ( .A(n6007), .B(n6005), .Z(n6773) );
  AND U6604 ( .A(n6774), .B(n6775), .Z(n6008) );
  NAND U6605 ( .A(n6776), .B(n5984), .Z(n6774) );
  NAND U6606 ( .A(n6777), .B(n6778), .Z(n5984) );
  NANDN U6607 ( .A(n5960), .B(n6779), .Z(n6778) );
  OR U6608 ( .A(n5959), .B(n5957), .Z(n6779) );
  AND U6609 ( .A(n6780), .B(n6781), .Z(n5960) );
  NAND U6610 ( .A(n6782), .B(n5936), .Z(n6780) );
  NAND U6611 ( .A(n6783), .B(n6784), .Z(n5936) );
  NANDN U6612 ( .A(n5912), .B(n6785), .Z(n6784) );
  OR U6613 ( .A(n5911), .B(n5909), .Z(n6785) );
  AND U6614 ( .A(n6786), .B(n6787), .Z(n5912) );
  NAND U6615 ( .A(n6788), .B(n5888), .Z(n6786) );
  NAND U6616 ( .A(n6789), .B(n6790), .Z(n5888) );
  NANDN U6617 ( .A(n5864), .B(n6791), .Z(n6790) );
  OR U6618 ( .A(n5863), .B(n5861), .Z(n6791) );
  AND U6619 ( .A(n6792), .B(n6793), .Z(n5864) );
  NAND U6620 ( .A(n6794), .B(n5840), .Z(n6792) );
  NAND U6621 ( .A(n6795), .B(n6796), .Z(n5840) );
  NANDN U6622 ( .A(n5816), .B(n6797), .Z(n6796) );
  OR U6623 ( .A(n5815), .B(n5813), .Z(n6797) );
  AND U6624 ( .A(n6798), .B(n6799), .Z(n5816) );
  NAND U6625 ( .A(n6800), .B(n5792), .Z(n6798) );
  NAND U6626 ( .A(n6801), .B(n6802), .Z(n5792) );
  NANDN U6627 ( .A(n5768), .B(n6803), .Z(n6802) );
  OR U6628 ( .A(n5767), .B(n5765), .Z(n6803) );
  AND U6629 ( .A(n6804), .B(n6805), .Z(n5768) );
  NAND U6630 ( .A(n6806), .B(n5744), .Z(n6804) );
  NAND U6631 ( .A(n6807), .B(n6808), .Z(n5744) );
  NANDN U6632 ( .A(n5720), .B(n6809), .Z(n6808) );
  OR U6633 ( .A(n5719), .B(n5717), .Z(n6809) );
  AND U6634 ( .A(n6810), .B(n6811), .Z(n5720) );
  NAND U6635 ( .A(n6812), .B(n5696), .Z(n6810) );
  NAND U6636 ( .A(n6813), .B(n6814), .Z(n5696) );
  NANDN U6637 ( .A(n5672), .B(n6815), .Z(n6814) );
  OR U6638 ( .A(n5671), .B(n5669), .Z(n6815) );
  AND U6639 ( .A(n6816), .B(n6817), .Z(n5672) );
  NAND U6640 ( .A(n6818), .B(n5648), .Z(n6816) );
  NAND U6641 ( .A(n6819), .B(n6820), .Z(n5648) );
  NANDN U6642 ( .A(n5624), .B(n6821), .Z(n6820) );
  OR U6643 ( .A(n5623), .B(n5621), .Z(n6821) );
  AND U6644 ( .A(n6822), .B(n6823), .Z(n5624) );
  NAND U6645 ( .A(n6824), .B(n5600), .Z(n6822) );
  NAND U6646 ( .A(n6825), .B(n6826), .Z(n5600) );
  NANDN U6647 ( .A(n5576), .B(n6827), .Z(n6826) );
  OR U6648 ( .A(n5575), .B(n5573), .Z(n6827) );
  AND U6649 ( .A(n6828), .B(n6829), .Z(n5576) );
  NAND U6650 ( .A(n6830), .B(n5552), .Z(n6828) );
  NAND U6651 ( .A(n6831), .B(n6832), .Z(n5552) );
  NANDN U6652 ( .A(n5528), .B(n6833), .Z(n6832) );
  OR U6653 ( .A(n5527), .B(n5525), .Z(n6833) );
  AND U6654 ( .A(n6834), .B(n6835), .Z(n5528) );
  NAND U6655 ( .A(n6836), .B(n5504), .Z(n6834) );
  NAND U6656 ( .A(n6837), .B(n6838), .Z(n5504) );
  NANDN U6657 ( .A(n5480), .B(n6839), .Z(n6838) );
  OR U6658 ( .A(n5479), .B(n5477), .Z(n6839) );
  AND U6659 ( .A(n6840), .B(n6841), .Z(n5480) );
  OR U6660 ( .A(n5453), .B(n5455), .Z(n6841) );
  NANDN U6661 ( .A(n5456), .B(n6842), .Z(n6840) );
  NAND U6662 ( .A(n5453), .B(n5455), .Z(n6842) );
  AND U6663 ( .A(n6843), .B(n6844), .Z(n5455) );
  OR U6664 ( .A(n5429), .B(n5431), .Z(n6844) );
  NANDN U6665 ( .A(n5432), .B(n6845), .Z(n6843) );
  NAND U6666 ( .A(n5429), .B(n5431), .Z(n6845) );
  AND U6667 ( .A(n6846), .B(n6847), .Z(n5431) );
  NANDN U6668 ( .A(n5408), .B(n6848), .Z(n6847) );
  NANDN U6669 ( .A(n5405), .B(n5407), .Z(n6848) );
  NANDN U6670 ( .A(n5398), .B(\stack[1][0] ), .Z(n5408) );
  NANDN U6671 ( .A(n5407), .B(n5405), .Z(n6846) );
  XNOR U6672 ( .A(n6849), .B(n6850), .Z(n5405) );
  XNOR U6673 ( .A(n6851), .B(n6852), .Z(n6850) );
  AND U6674 ( .A(n6853), .B(n6854), .Z(n5407) );
  NANDN U6675 ( .A(n5381), .B(n5384), .Z(n6854) );
  NANDN U6676 ( .A(n5383), .B(n6855), .Z(n6853) );
  NANDN U6677 ( .A(n5384), .B(n5381), .Z(n6855) );
  XOR U6678 ( .A(n6856), .B(n6857), .Z(n5381) );
  XNOR U6679 ( .A(n6858), .B(n6859), .Z(n6857) );
  NAND U6680 ( .A(n6860), .B(n6861), .Z(n5384) );
  NANDN U6681 ( .A(n5360), .B(n6862), .Z(n6861) );
  NANDN U6682 ( .A(n5357), .B(n5359), .Z(n6862) );
  NANDN U6683 ( .A(n5169), .B(\stack[0][8] ), .Z(n5360) );
  NANDN U6684 ( .A(n5359), .B(n5357), .Z(n6860) );
  XNOR U6685 ( .A(n6863), .B(n6864), .Z(n5357) );
  XNOR U6686 ( .A(n6865), .B(n6866), .Z(n6864) );
  AND U6687 ( .A(n6867), .B(n6868), .Z(n5359) );
  OR U6688 ( .A(n5333), .B(n5335), .Z(n6868) );
  NANDN U6689 ( .A(n5336), .B(n6869), .Z(n6867) );
  NAND U6690 ( .A(n5333), .B(n5335), .Z(n6869) );
  AND U6691 ( .A(n6870), .B(n6871), .Z(n5335) );
  NANDN U6692 ( .A(n5312), .B(n6872), .Z(n6871) );
  NANDN U6693 ( .A(n5309), .B(n5311), .Z(n6872) );
  NANDN U6694 ( .A(n5169), .B(\stack[0][6] ), .Z(n5312) );
  NANDN U6695 ( .A(n5311), .B(n5309), .Z(n6870) );
  XNOR U6696 ( .A(n6873), .B(n6874), .Z(n5309) );
  XNOR U6697 ( .A(n6875), .B(n6876), .Z(n6874) );
  AND U6698 ( .A(n6877), .B(n6878), .Z(n5311) );
  OR U6699 ( .A(n5285), .B(n5287), .Z(n6878) );
  NANDN U6700 ( .A(n5288), .B(n6879), .Z(n6877) );
  NAND U6701 ( .A(n5285), .B(n5287), .Z(n6879) );
  AND U6702 ( .A(n6880), .B(n6881), .Z(n5287) );
  NANDN U6703 ( .A(n5264), .B(n6882), .Z(n6881) );
  NANDN U6704 ( .A(n5261), .B(n5263), .Z(n6882) );
  NANDN U6705 ( .A(n5169), .B(\stack[0][4] ), .Z(n5264) );
  NANDN U6706 ( .A(n5263), .B(n5261), .Z(n6880) );
  XNOR U6707 ( .A(n6883), .B(n6884), .Z(n5261) );
  XNOR U6708 ( .A(n6885), .B(n6886), .Z(n6884) );
  AND U6709 ( .A(n6887), .B(n6888), .Z(n5263) );
  NANDN U6710 ( .A(n5237), .B(n5239), .Z(n6888) );
  NANDN U6711 ( .A(n5240), .B(n6889), .Z(n6887) );
  NANDN U6712 ( .A(n5239), .B(n5237), .Z(n6889) );
  XNOR U6713 ( .A(n6890), .B(n6891), .Z(n5237) );
  XNOR U6714 ( .A(n6892), .B(n6893), .Z(n6891) );
  ANDN U6715 ( .B(\stack[1][0] ), .A(n5230), .Z(n5239) );
  AND U6716 ( .A(n6894), .B(n6895), .Z(n5240) );
  NANDN U6717 ( .A(n5213), .B(n5215), .Z(n6895) );
  NANDN U6718 ( .A(n5216), .B(n6896), .Z(n6894) );
  NANDN U6719 ( .A(n5215), .B(n5213), .Z(n6896) );
  XNOR U6720 ( .A(n6897), .B(n6898), .Z(n5213) );
  NANDN U6721 ( .A(n5160), .B(\stack[1][2] ), .Z(n6898) );
  NOR U6722 ( .A(n5191), .B(n5192), .Z(n5215) );
  NANDN U6723 ( .A(n5169), .B(\stack[0][1] ), .Z(n5192) );
  NANDN U6724 ( .A(n5195), .B(\stack[0][0] ), .Z(n5191) );
  NANDN U6725 ( .A(n5169), .B(\stack[0][2] ), .Z(n5216) );
  XOR U6726 ( .A(n6899), .B(n6900), .Z(n5285) );
  XNOR U6727 ( .A(n6901), .B(n6902), .Z(n6900) );
  NANDN U6728 ( .A(n5278), .B(\stack[1][0] ), .Z(n5288) );
  XOR U6729 ( .A(n6903), .B(n6904), .Z(n5333) );
  XNOR U6730 ( .A(n6905), .B(n6906), .Z(n6904) );
  NANDN U6731 ( .A(n5326), .B(\stack[1][0] ), .Z(n5336) );
  NANDN U6732 ( .A(n5169), .B(\stack[0][9] ), .Z(n5383) );
  XOR U6733 ( .A(n6907), .B(n6908), .Z(n5429) );
  XNOR U6734 ( .A(n6909), .B(n6910), .Z(n6908) );
  NANDN U6735 ( .A(n5169), .B(\stack[0][11] ), .Z(n5432) );
  XOR U6736 ( .A(n6911), .B(n6912), .Z(n5453) );
  XNOR U6737 ( .A(n6913), .B(n6914), .Z(n6912) );
  NANDN U6738 ( .A(n5446), .B(\stack[1][0] ), .Z(n5456) );
  NAND U6739 ( .A(n5477), .B(n5479), .Z(n6837) );
  AND U6740 ( .A(\stack[1][0] ), .B(\stack[0][13] ), .Z(n5479) );
  XNOR U6741 ( .A(n6915), .B(n6916), .Z(n5477) );
  XNOR U6742 ( .A(n6917), .B(n6918), .Z(n6916) );
  NANDN U6743 ( .A(n5503), .B(n5501), .Z(n6836) );
  XOR U6744 ( .A(n6919), .B(n6920), .Z(n5501) );
  XNOR U6745 ( .A(n6921), .B(n6922), .Z(n6920) );
  ANDN U6746 ( .B(\stack[1][0] ), .A(n5494), .Z(n5503) );
  NAND U6747 ( .A(n5525), .B(n5527), .Z(n6831) );
  AND U6748 ( .A(\stack[1][0] ), .B(\stack[0][15] ), .Z(n5527) );
  XNOR U6749 ( .A(n6923), .B(n6924), .Z(n5525) );
  XNOR U6750 ( .A(n6925), .B(n6926), .Z(n6924) );
  NANDN U6751 ( .A(n5551), .B(n5549), .Z(n6830) );
  XOR U6752 ( .A(n6927), .B(n6928), .Z(n5549) );
  XNOR U6753 ( .A(n6929), .B(n6930), .Z(n6928) );
  ANDN U6754 ( .B(\stack[1][0] ), .A(n5542), .Z(n5551) );
  NAND U6755 ( .A(n5573), .B(n5575), .Z(n6825) );
  AND U6756 ( .A(\stack[1][0] ), .B(\stack[0][17] ), .Z(n5575) );
  XNOR U6757 ( .A(n6931), .B(n6932), .Z(n5573) );
  XNOR U6758 ( .A(n6933), .B(n6934), .Z(n6932) );
  NANDN U6759 ( .A(n5599), .B(n5597), .Z(n6824) );
  XOR U6760 ( .A(n6935), .B(n6936), .Z(n5597) );
  XNOR U6761 ( .A(n6937), .B(n6938), .Z(n6936) );
  ANDN U6762 ( .B(\stack[1][0] ), .A(n5590), .Z(n5599) );
  NAND U6763 ( .A(n5621), .B(n5623), .Z(n6819) );
  AND U6764 ( .A(\stack[1][0] ), .B(\stack[0][19] ), .Z(n5623) );
  XNOR U6765 ( .A(n6939), .B(n6940), .Z(n5621) );
  XNOR U6766 ( .A(n6941), .B(n6942), .Z(n6940) );
  NANDN U6767 ( .A(n5647), .B(n5645), .Z(n6818) );
  XOR U6768 ( .A(n6943), .B(n6944), .Z(n5645) );
  XNOR U6769 ( .A(n6945), .B(n6946), .Z(n6944) );
  ANDN U6770 ( .B(\stack[1][0] ), .A(n5638), .Z(n5647) );
  NAND U6771 ( .A(n5669), .B(n5671), .Z(n6813) );
  AND U6772 ( .A(\stack[1][0] ), .B(\stack[0][21] ), .Z(n5671) );
  XNOR U6773 ( .A(n6947), .B(n6948), .Z(n5669) );
  XNOR U6774 ( .A(n6949), .B(n6950), .Z(n6948) );
  NANDN U6775 ( .A(n5695), .B(n5693), .Z(n6812) );
  XOR U6776 ( .A(n6951), .B(n6952), .Z(n5693) );
  XNOR U6777 ( .A(n6953), .B(n6954), .Z(n6952) );
  ANDN U6778 ( .B(\stack[1][0] ), .A(n5686), .Z(n5695) );
  NAND U6779 ( .A(n5717), .B(n5719), .Z(n6807) );
  AND U6780 ( .A(\stack[1][0] ), .B(\stack[0][23] ), .Z(n5719) );
  XNOR U6781 ( .A(n6955), .B(n6956), .Z(n5717) );
  XNOR U6782 ( .A(n6957), .B(n6958), .Z(n6956) );
  NANDN U6783 ( .A(n5743), .B(n5741), .Z(n6806) );
  XOR U6784 ( .A(n6959), .B(n6960), .Z(n5741) );
  XNOR U6785 ( .A(n6961), .B(n6962), .Z(n6960) );
  ANDN U6786 ( .B(\stack[1][0] ), .A(n5734), .Z(n5743) );
  NAND U6787 ( .A(n5765), .B(n5767), .Z(n6801) );
  AND U6788 ( .A(\stack[1][0] ), .B(\stack[0][25] ), .Z(n5767) );
  XNOR U6789 ( .A(n6963), .B(n6964), .Z(n5765) );
  XNOR U6790 ( .A(n6965), .B(n6966), .Z(n6964) );
  NANDN U6791 ( .A(n5791), .B(n5789), .Z(n6800) );
  XOR U6792 ( .A(n6967), .B(n6968), .Z(n5789) );
  XNOR U6793 ( .A(n6969), .B(n6970), .Z(n6968) );
  ANDN U6794 ( .B(\stack[1][0] ), .A(n5782), .Z(n5791) );
  NAND U6795 ( .A(n5813), .B(n5815), .Z(n6795) );
  AND U6796 ( .A(\stack[1][0] ), .B(\stack[0][27] ), .Z(n5815) );
  XNOR U6797 ( .A(n6971), .B(n6972), .Z(n5813) );
  XNOR U6798 ( .A(n6973), .B(n6974), .Z(n6972) );
  NANDN U6799 ( .A(n5839), .B(n5837), .Z(n6794) );
  XOR U6800 ( .A(n6975), .B(n6976), .Z(n5837) );
  XNOR U6801 ( .A(n6977), .B(n6978), .Z(n6976) );
  ANDN U6802 ( .B(\stack[1][0] ), .A(n5830), .Z(n5839) );
  NAND U6803 ( .A(n5861), .B(n5863), .Z(n6789) );
  AND U6804 ( .A(\stack[1][0] ), .B(\stack[0][29] ), .Z(n5863) );
  XNOR U6805 ( .A(n6979), .B(n6980), .Z(n5861) );
  XNOR U6806 ( .A(n6981), .B(n6982), .Z(n6980) );
  NANDN U6807 ( .A(n5887), .B(n5885), .Z(n6788) );
  XOR U6808 ( .A(n6983), .B(n6984), .Z(n5885) );
  XNOR U6809 ( .A(n6985), .B(n6986), .Z(n6984) );
  ANDN U6810 ( .B(\stack[1][0] ), .A(n5878), .Z(n5887) );
  NAND U6811 ( .A(n5909), .B(n5911), .Z(n6783) );
  AND U6812 ( .A(\stack[1][0] ), .B(\stack[0][31] ), .Z(n5911) );
  XNOR U6813 ( .A(n6987), .B(n6988), .Z(n5909) );
  XNOR U6814 ( .A(n6989), .B(n6990), .Z(n6988) );
  NANDN U6815 ( .A(n5935), .B(n5933), .Z(n6782) );
  XOR U6816 ( .A(n6991), .B(n6992), .Z(n5933) );
  XNOR U6817 ( .A(n6993), .B(n6994), .Z(n6992) );
  ANDN U6818 ( .B(\stack[1][0] ), .A(n5926), .Z(n5935) );
  NAND U6819 ( .A(n5957), .B(n5959), .Z(n6777) );
  AND U6820 ( .A(\stack[1][0] ), .B(\stack[0][33] ), .Z(n5959) );
  XNOR U6821 ( .A(n6995), .B(n6996), .Z(n5957) );
  XNOR U6822 ( .A(n6997), .B(n6998), .Z(n6996) );
  NANDN U6823 ( .A(n5983), .B(n5981), .Z(n6776) );
  XOR U6824 ( .A(n6999), .B(n7000), .Z(n5981) );
  XNOR U6825 ( .A(n7001), .B(n7002), .Z(n7000) );
  ANDN U6826 ( .B(\stack[1][0] ), .A(n5974), .Z(n5983) );
  NAND U6827 ( .A(n6005), .B(n6007), .Z(n6771) );
  AND U6828 ( .A(\stack[1][0] ), .B(\stack[0][35] ), .Z(n6007) );
  XNOR U6829 ( .A(n7003), .B(n7004), .Z(n6005) );
  XNOR U6830 ( .A(n7005), .B(n7006), .Z(n7004) );
  NANDN U6831 ( .A(n6031), .B(n6029), .Z(n6770) );
  XOR U6832 ( .A(n7007), .B(n7008), .Z(n6029) );
  XNOR U6833 ( .A(n7009), .B(n7010), .Z(n7008) );
  ANDN U6834 ( .B(\stack[1][0] ), .A(n6022), .Z(n6031) );
  NAND U6835 ( .A(n6053), .B(n6055), .Z(n6765) );
  AND U6836 ( .A(\stack[1][0] ), .B(\stack[0][37] ), .Z(n6055) );
  XNOR U6837 ( .A(n7011), .B(n7012), .Z(n6053) );
  XNOR U6838 ( .A(n7013), .B(n7014), .Z(n7012) );
  NANDN U6839 ( .A(n6079), .B(n6077), .Z(n6764) );
  XOR U6840 ( .A(n7015), .B(n7016), .Z(n6077) );
  XNOR U6841 ( .A(n7017), .B(n7018), .Z(n7016) );
  ANDN U6842 ( .B(\stack[1][0] ), .A(n6070), .Z(n6079) );
  NAND U6843 ( .A(n6101), .B(n6103), .Z(n6759) );
  AND U6844 ( .A(\stack[1][0] ), .B(\stack[0][39] ), .Z(n6103) );
  XNOR U6845 ( .A(n7019), .B(n7020), .Z(n6101) );
  XNOR U6846 ( .A(n7021), .B(n7022), .Z(n7020) );
  NANDN U6847 ( .A(n6127), .B(n6125), .Z(n6758) );
  XOR U6848 ( .A(n7023), .B(n7024), .Z(n6125) );
  XNOR U6849 ( .A(n7025), .B(n7026), .Z(n7024) );
  ANDN U6850 ( .B(\stack[1][0] ), .A(n6118), .Z(n6127) );
  NAND U6851 ( .A(n6149), .B(n6151), .Z(n6753) );
  AND U6852 ( .A(\stack[1][0] ), .B(\stack[0][41] ), .Z(n6151) );
  XNOR U6853 ( .A(n7027), .B(n7028), .Z(n6149) );
  XNOR U6854 ( .A(n7029), .B(n7030), .Z(n7028) );
  NANDN U6855 ( .A(n6175), .B(n6173), .Z(n6752) );
  XOR U6856 ( .A(n7031), .B(n7032), .Z(n6173) );
  XNOR U6857 ( .A(n7033), .B(n7034), .Z(n7032) );
  ANDN U6858 ( .B(\stack[1][0] ), .A(n6166), .Z(n6175) );
  NAND U6859 ( .A(n6197), .B(n6199), .Z(n6747) );
  AND U6860 ( .A(\stack[1][0] ), .B(\stack[0][43] ), .Z(n6199) );
  XNOR U6861 ( .A(n7035), .B(n7036), .Z(n6197) );
  XNOR U6862 ( .A(n7037), .B(n7038), .Z(n7036) );
  NANDN U6863 ( .A(n6223), .B(n6221), .Z(n6746) );
  XOR U6864 ( .A(n7039), .B(n7040), .Z(n6221) );
  XNOR U6865 ( .A(n7041), .B(n7042), .Z(n7040) );
  ANDN U6866 ( .B(\stack[1][0] ), .A(n6214), .Z(n6223) );
  NAND U6867 ( .A(n6245), .B(n6247), .Z(n6741) );
  AND U6868 ( .A(\stack[1][0] ), .B(\stack[0][45] ), .Z(n6247) );
  XNOR U6869 ( .A(n7043), .B(n7044), .Z(n6245) );
  XNOR U6870 ( .A(n7045), .B(n7046), .Z(n7044) );
  NANDN U6871 ( .A(n6271), .B(n6269), .Z(n6740) );
  XOR U6872 ( .A(n7047), .B(n7048), .Z(n6269) );
  XNOR U6873 ( .A(n7049), .B(n7050), .Z(n7048) );
  ANDN U6874 ( .B(\stack[1][0] ), .A(n6262), .Z(n6271) );
  NAND U6875 ( .A(n6293), .B(n6295), .Z(n6735) );
  AND U6876 ( .A(\stack[1][0] ), .B(\stack[0][47] ), .Z(n6295) );
  XNOR U6877 ( .A(n7051), .B(n7052), .Z(n6293) );
  XNOR U6878 ( .A(n7053), .B(n7054), .Z(n7052) );
  NANDN U6879 ( .A(n6319), .B(n6317), .Z(n6734) );
  XOR U6880 ( .A(n7055), .B(n7056), .Z(n6317) );
  XNOR U6881 ( .A(n7057), .B(n7058), .Z(n7056) );
  ANDN U6882 ( .B(\stack[1][0] ), .A(n6310), .Z(n6319) );
  NAND U6883 ( .A(n6341), .B(n6343), .Z(n6729) );
  AND U6884 ( .A(\stack[1][0] ), .B(\stack[0][49] ), .Z(n6343) );
  XNOR U6885 ( .A(n7059), .B(n7060), .Z(n6341) );
  XNOR U6886 ( .A(n7061), .B(n7062), .Z(n7060) );
  NANDN U6887 ( .A(n6367), .B(n6365), .Z(n6728) );
  XOR U6888 ( .A(n7063), .B(n7064), .Z(n6365) );
  XNOR U6889 ( .A(n7065), .B(n7066), .Z(n7064) );
  ANDN U6890 ( .B(\stack[1][0] ), .A(n6358), .Z(n6367) );
  NAND U6891 ( .A(n6389), .B(n6391), .Z(n6723) );
  AND U6892 ( .A(\stack[1][0] ), .B(\stack[0][51] ), .Z(n6391) );
  XNOR U6893 ( .A(n7067), .B(n7068), .Z(n6389) );
  XNOR U6894 ( .A(n7069), .B(n7070), .Z(n7068) );
  NANDN U6895 ( .A(n6415), .B(n6413), .Z(n6722) );
  XOR U6896 ( .A(n7071), .B(n7072), .Z(n6413) );
  XNOR U6897 ( .A(n7073), .B(n7074), .Z(n7072) );
  ANDN U6898 ( .B(\stack[1][0] ), .A(n6406), .Z(n6415) );
  NAND U6899 ( .A(n6437), .B(n6439), .Z(n6717) );
  AND U6900 ( .A(\stack[1][0] ), .B(\stack[0][53] ), .Z(n6439) );
  XNOR U6901 ( .A(n7075), .B(n7076), .Z(n6437) );
  XNOR U6902 ( .A(n7077), .B(n7078), .Z(n7076) );
  NANDN U6903 ( .A(n6463), .B(n6461), .Z(n6716) );
  XOR U6904 ( .A(n7079), .B(n7080), .Z(n6461) );
  XNOR U6905 ( .A(n7081), .B(n7082), .Z(n7080) );
  ANDN U6906 ( .B(\stack[1][0] ), .A(n6454), .Z(n6463) );
  NAND U6907 ( .A(n6485), .B(n6487), .Z(n6711) );
  AND U6908 ( .A(\stack[1][0] ), .B(\stack[0][55] ), .Z(n6487) );
  XNOR U6909 ( .A(n7083), .B(n7084), .Z(n6485) );
  XNOR U6910 ( .A(n7085), .B(n7086), .Z(n7084) );
  NANDN U6911 ( .A(n6511), .B(n6509), .Z(n6710) );
  XOR U6912 ( .A(n7087), .B(n7088), .Z(n6509) );
  XNOR U6913 ( .A(n7089), .B(n7090), .Z(n7088) );
  ANDN U6914 ( .B(\stack[1][0] ), .A(n6502), .Z(n6511) );
  NAND U6915 ( .A(n6533), .B(n6535), .Z(n6705) );
  AND U6916 ( .A(\stack[1][0] ), .B(\stack[0][57] ), .Z(n6535) );
  XNOR U6917 ( .A(n7091), .B(n7092), .Z(n6533) );
  XNOR U6918 ( .A(n7093), .B(n7094), .Z(n7092) );
  NANDN U6919 ( .A(n6559), .B(n6557), .Z(n6704) );
  XOR U6920 ( .A(n7095), .B(n7096), .Z(n6557) );
  XNOR U6921 ( .A(n7097), .B(n7098), .Z(n7096) );
  ANDN U6922 ( .B(\stack[1][0] ), .A(n6550), .Z(n6559) );
  NAND U6923 ( .A(n6581), .B(n6583), .Z(n6699) );
  AND U6924 ( .A(\stack[1][0] ), .B(\stack[0][59] ), .Z(n6583) );
  XNOR U6925 ( .A(n7099), .B(n7100), .Z(n6581) );
  XNOR U6926 ( .A(n7101), .B(n7102), .Z(n7100) );
  NANDN U6927 ( .A(n6607), .B(n6605), .Z(n6698) );
  XOR U6928 ( .A(n7103), .B(n7104), .Z(n6605) );
  XNOR U6929 ( .A(n7105), .B(n7106), .Z(n7104) );
  ANDN U6930 ( .B(\stack[1][0] ), .A(n6598), .Z(n6607) );
  NAND U6931 ( .A(n6629), .B(n6631), .Z(n6693) );
  AND U6932 ( .A(\stack[1][0] ), .B(\stack[0][61] ), .Z(n6631) );
  XNOR U6933 ( .A(n7107), .B(n7108), .Z(n6629) );
  XNOR U6934 ( .A(n7109), .B(n7110), .Z(n7108) );
  NANDN U6935 ( .A(n6655), .B(n6653), .Z(n6692) );
  AND U6936 ( .A(n7111), .B(n7112), .Z(n6690) );
  NANDN U6937 ( .A(n6670), .B(n5169), .Z(n7112) );
  NANDN U6938 ( .A(n6653), .B(n6655), .Z(n7111) );
  AND U6939 ( .A(\stack[1][0] ), .B(\stack[0][62] ), .Z(n6655) );
  XOR U6940 ( .A(n7113), .B(n7114), .Z(n6653) );
  XNOR U6941 ( .A(n7115), .B(n7116), .Z(n7114) );
  XOR U6942 ( .A(n7117), .B(n7118), .Z(n6686) );
  XOR U6943 ( .A(n7119), .B(n7120), .Z(n7118) );
  XOR U6944 ( .A(n7121), .B(n7122), .Z(n7120) );
  XOR U6945 ( .A(n7123), .B(n7124), .Z(n7122) );
  XOR U6946 ( .A(n7125), .B(n7126), .Z(n7124) );
  XOR U6947 ( .A(n7127), .B(n7128), .Z(n7126) );
  XOR U6948 ( .A(n7129), .B(n7130), .Z(n7128) );
  AND U6949 ( .A(n7131), .B(n7132), .Z(n7130) );
  NANDN U6950 ( .A(n7133), .B(n7134), .Z(n7132) );
  NANDN U6951 ( .A(n7135), .B(n7136), .Z(n7131) );
  ANDN U6952 ( .B(\stack[1][2] ), .A(n6622), .Z(n7129) );
  XOR U6953 ( .A(n7137), .B(n7138), .Z(n7127) );
  XOR U6954 ( .A(n7139), .B(n7140), .Z(n7138) );
  XOR U6955 ( .A(n7141), .B(n7142), .Z(n7140) );
  XOR U6956 ( .A(n7143), .B(n7144), .Z(n7142) );
  AND U6957 ( .A(n7145), .B(n7146), .Z(n7144) );
  NANDN U6958 ( .A(n7147), .B(n7148), .Z(n7146) );
  NANDN U6959 ( .A(n7149), .B(n7150), .Z(n7145) );
  OR U6960 ( .A(n7148), .B(n7151), .Z(n7150) );
  ANDN U6961 ( .B(\stack[1][6] ), .A(n6526), .Z(n7143) );
  XOR U6962 ( .A(n7152), .B(n7153), .Z(n7141) );
  XOR U6963 ( .A(n7154), .B(n7155), .Z(n7153) );
  XOR U6964 ( .A(n7156), .B(n7157), .Z(n7155) );
  XOR U6965 ( .A(n7158), .B(n7159), .Z(n7157) );
  AND U6966 ( .A(n7160), .B(n7161), .Z(n7159) );
  NANDN U6967 ( .A(n7162), .B(n7163), .Z(n7161) );
  NANDN U6968 ( .A(n7164), .B(n7165), .Z(n7160) );
  NANDN U6969 ( .A(n7163), .B(n7162), .Z(n7165) );
  ANDN U6970 ( .B(\stack[1][10] ), .A(n6430), .Z(n7158) );
  XOR U6971 ( .A(n7166), .B(n7167), .Z(n7156) );
  XOR U6972 ( .A(n7168), .B(n7169), .Z(n7167) );
  XOR U6973 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U6974 ( .A(n7172), .B(n7173), .Z(n7171) );
  AND U6975 ( .A(n7174), .B(n7175), .Z(n7173) );
  NANDN U6976 ( .A(n7176), .B(n7177), .Z(n7175) );
  NANDN U6977 ( .A(n7178), .B(n7179), .Z(n7174) );
  NANDN U6978 ( .A(n7177), .B(n7176), .Z(n7179) );
  ANDN U6979 ( .B(\stack[1][14] ), .A(n6334), .Z(n7172) );
  XOR U6980 ( .A(n7180), .B(n7181), .Z(n7170) );
  XOR U6981 ( .A(n7182), .B(n7183), .Z(n7181) );
  XOR U6982 ( .A(n7184), .B(n7185), .Z(n7183) );
  XOR U6983 ( .A(n7186), .B(n7187), .Z(n7185) );
  AND U6984 ( .A(n7188), .B(n7189), .Z(n7187) );
  NANDN U6985 ( .A(n7190), .B(n7191), .Z(n7189) );
  NANDN U6986 ( .A(n7192), .B(n7193), .Z(n7188) );
  NANDN U6987 ( .A(n7191), .B(n7190), .Z(n7193) );
  ANDN U6988 ( .B(\stack[1][18] ), .A(n6238), .Z(n7186) );
  XOR U6989 ( .A(n7194), .B(n7195), .Z(n7184) );
  XOR U6990 ( .A(n7196), .B(n7197), .Z(n7195) );
  XOR U6991 ( .A(n7198), .B(n7199), .Z(n7197) );
  XOR U6992 ( .A(n7200), .B(n7201), .Z(n7199) );
  AND U6993 ( .A(n7202), .B(n7203), .Z(n7201) );
  NANDN U6994 ( .A(n7204), .B(n7205), .Z(n7203) );
  NANDN U6995 ( .A(n7206), .B(n7207), .Z(n7202) );
  NANDN U6996 ( .A(n7205), .B(n7204), .Z(n7207) );
  ANDN U6997 ( .B(\stack[1][22] ), .A(n6142), .Z(n7200) );
  XOR U6998 ( .A(n7208), .B(n7209), .Z(n7198) );
  XOR U6999 ( .A(n7210), .B(n7211), .Z(n7209) );
  XOR U7000 ( .A(n7212), .B(n7213), .Z(n7211) );
  XOR U7001 ( .A(n7214), .B(n7215), .Z(n7213) );
  AND U7002 ( .A(n7216), .B(n7217), .Z(n7215) );
  NANDN U7003 ( .A(n7218), .B(n7219), .Z(n7217) );
  NANDN U7004 ( .A(n7220), .B(n7221), .Z(n7216) );
  NANDN U7005 ( .A(n7219), .B(n7218), .Z(n7221) );
  ANDN U7006 ( .B(\stack[1][26] ), .A(n6046), .Z(n7214) );
  XOR U7007 ( .A(n7222), .B(n7223), .Z(n7212) );
  XOR U7008 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U7009 ( .A(n7226), .B(n7227), .Z(n7225) );
  XOR U7010 ( .A(n7228), .B(n7229), .Z(n7227) );
  AND U7011 ( .A(n7230), .B(n7231), .Z(n7229) );
  NANDN U7012 ( .A(n7232), .B(n7233), .Z(n7231) );
  NANDN U7013 ( .A(n7234), .B(n7235), .Z(n7230) );
  NANDN U7014 ( .A(n7233), .B(n7232), .Z(n7235) );
  ANDN U7015 ( .B(\stack[1][30] ), .A(n5950), .Z(n7228) );
  XOR U7016 ( .A(n7236), .B(n7237), .Z(n7226) );
  XOR U7017 ( .A(n7238), .B(n7239), .Z(n7237) );
  XOR U7018 ( .A(n7240), .B(n7241), .Z(n7239) );
  AND U7019 ( .A(n7242), .B(n7243), .Z(n7241) );
  NANDN U7020 ( .A(n7244), .B(n7245), .Z(n7243) );
  NANDN U7021 ( .A(n7246), .B(n7247), .Z(n7242) );
  NANDN U7022 ( .A(n7245), .B(n7244), .Z(n7247) );
  ANDN U7023 ( .B(\stack[1][34] ), .A(n5854), .Z(n7240) );
  XOR U7024 ( .A(n7248), .B(n7249), .Z(n7238) );
  XOR U7025 ( .A(n7250), .B(n7251), .Z(n7249) );
  XOR U7026 ( .A(n7252), .B(n7253), .Z(n7251) );
  ANDN U7027 ( .B(\stack[1][38] ), .A(n5758), .Z(n7253) );
  AND U7028 ( .A(n7254), .B(n7255), .Z(n7252) );
  NANDN U7029 ( .A(n7256), .B(n7257), .Z(n7255) );
  NANDN U7030 ( .A(n7258), .B(n7259), .Z(n7254) );
  NANDN U7031 ( .A(n7260), .B(n7261), .Z(n7259) );
  XOR U7032 ( .A(n7262), .B(n7263), .Z(n7250) );
  XOR U7033 ( .A(n7264), .B(n7265), .Z(n7263) );
  XOR U7034 ( .A(n7266), .B(n7267), .Z(n7265) );
  AND U7035 ( .A(n7268), .B(n7269), .Z(n7267) );
  NANDN U7036 ( .A(n7270), .B(n7271), .Z(n7269) );
  NANDN U7037 ( .A(n7272), .B(n7273), .Z(n7268) );
  OR U7038 ( .A(n7271), .B(n7274), .Z(n7273) );
  ANDN U7039 ( .B(\stack[1][41] ), .A(n5686), .Z(n7266) );
  XOR U7040 ( .A(n7275), .B(n7276), .Z(n7264) );
  XOR U7041 ( .A(n7277), .B(n7278), .Z(n7276) );
  XOR U7042 ( .A(n7279), .B(n7280), .Z(n7278) );
  AND U7043 ( .A(n7281), .B(n7282), .Z(n7280) );
  NANDN U7044 ( .A(n7283), .B(n7284), .Z(n7282) );
  NANDN U7045 ( .A(n7285), .B(n7286), .Z(n7281) );
  NANDN U7046 ( .A(n7284), .B(n7283), .Z(n7286) );
  ANDN U7047 ( .B(\stack[1][44] ), .A(n5614), .Z(n7279) );
  XOR U7048 ( .A(n7287), .B(n7288), .Z(n7277) );
  XOR U7049 ( .A(n7289), .B(n7290), .Z(n7288) );
  XOR U7050 ( .A(n7291), .B(n7292), .Z(n7290) );
  AND U7051 ( .A(n7293), .B(n7294), .Z(n7292) );
  NANDN U7052 ( .A(n7295), .B(n7296), .Z(n7294) );
  NANDN U7053 ( .A(n7297), .B(n7298), .Z(n7293) );
  OR U7054 ( .A(n7296), .B(n7299), .Z(n7298) );
  ANDN U7055 ( .B(\stack[1][47] ), .A(n5542), .Z(n7291) );
  XOR U7056 ( .A(n7300), .B(n7301), .Z(n7289) );
  XOR U7057 ( .A(n7302), .B(n7303), .Z(n7301) );
  XOR U7058 ( .A(n7304), .B(n7305), .Z(n7303) );
  AND U7059 ( .A(n7306), .B(n7307), .Z(n7305) );
  NANDN U7060 ( .A(n7308), .B(n7309), .Z(n7307) );
  NANDN U7061 ( .A(n7310), .B(n7311), .Z(n7306) );
  NANDN U7062 ( .A(n7309), .B(n7308), .Z(n7311) );
  ANDN U7063 ( .B(\stack[1][50] ), .A(n5470), .Z(n7304) );
  XOR U7064 ( .A(n7312), .B(n7313), .Z(n7302) );
  XOR U7065 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U7066 ( .A(n7316), .B(n7317), .Z(n7315) );
  AND U7067 ( .A(n7318), .B(n7319), .Z(n7317) );
  NANDN U7068 ( .A(n7320), .B(n7321), .Z(n7319) );
  NANDN U7069 ( .A(n7322), .B(n7323), .Z(n7318) );
  OR U7070 ( .A(n7321), .B(n7324), .Z(n7323) );
  ANDN U7071 ( .B(\stack[1][53] ), .A(n5398), .Z(n7316) );
  XOR U7072 ( .A(n7325), .B(n7326), .Z(n7314) );
  XOR U7073 ( .A(n7327), .B(n7328), .Z(n7326) );
  XOR U7074 ( .A(n7329), .B(n7330), .Z(n7328) );
  AND U7075 ( .A(n7331), .B(n7332), .Z(n7330) );
  NANDN U7076 ( .A(n5160), .B(n7333), .Z(n7332) );
  NOR U7077 ( .A(n6659), .B(n7334), .Z(n7333) );
  NANDN U7078 ( .A(n6684), .B(n5160), .Z(n7331) );
  XOR U7079 ( .A(n7335), .B(n7336), .Z(n7329) );
  AND U7080 ( .A(n7337), .B(n7338), .Z(n7336) );
  NANDN U7081 ( .A(n7339), .B(n7340), .Z(n7338) );
  NANDN U7082 ( .A(n7341), .B(n7342), .Z(n7337) );
  NANDN U7083 ( .A(n7340), .B(n7339), .Z(n7342) );
  ANDN U7084 ( .B(\stack[0][7] ), .A(n6516), .Z(n7335) );
  XOR U7085 ( .A(n7343), .B(n7344), .Z(n7327) );
  ANDN U7086 ( .B(\stack[0][1] ), .A(n6659), .Z(n7344) );
  AND U7087 ( .A(n7345), .B(n7346), .Z(n7343) );
  NANDN U7088 ( .A(n7347), .B(n7348), .Z(n7346) );
  NANDN U7089 ( .A(n7349), .B(n7350), .Z(n7345) );
  OR U7090 ( .A(n7348), .B(n7351), .Z(n7350) );
  XOR U7091 ( .A(n7352), .B(n7353), .Z(n7325) );
  XOR U7092 ( .A(n7354), .B(n7355), .Z(n7353) );
  ANDN U7093 ( .B(\stack[0][4] ), .A(n6588), .Z(n7355) );
  AND U7094 ( .A(n7356), .B(n7357), .Z(n7354) );
  NAND U7095 ( .A(n7358), .B(n7359), .Z(n7357) );
  NANDN U7096 ( .A(n7360), .B(n7361), .Z(n7356) );
  OR U7097 ( .A(n7358), .B(n7359), .Z(n7361) );
  XOR U7098 ( .A(n7362), .B(n7363), .Z(n7352) );
  ANDN U7099 ( .B(\stack[0][3] ), .A(n6612), .Z(n7363) );
  ANDN U7100 ( .B(\stack[0][2] ), .A(n6636), .Z(n7362) );
  XOR U7101 ( .A(n7364), .B(n7365), .Z(n7312) );
  XOR U7102 ( .A(n7366), .B(n7367), .Z(n7365) );
  AND U7103 ( .A(n7368), .B(n7369), .Z(n7367) );
  NANDN U7104 ( .A(n7370), .B(n7371), .Z(n7369) );
  NANDN U7105 ( .A(n7372), .B(n7373), .Z(n7368) );
  OR U7106 ( .A(n7371), .B(n7374), .Z(n7373) );
  ANDN U7107 ( .B(\stack[0][6] ), .A(n6540), .Z(n7366) );
  XOR U7108 ( .A(n7375), .B(n7376), .Z(n7364) );
  AND U7109 ( .A(n7377), .B(n7378), .Z(n7376) );
  NANDN U7110 ( .A(n7379), .B(n7380), .Z(n7378) );
  NANDN U7111 ( .A(n7381), .B(n7382), .Z(n7377) );
  NANDN U7112 ( .A(n7380), .B(n7379), .Z(n7382) );
  ANDN U7113 ( .B(\stack[0][5] ), .A(n6564), .Z(n7375) );
  XOR U7114 ( .A(n7383), .B(n7384), .Z(n7300) );
  XOR U7115 ( .A(n7385), .B(n7386), .Z(n7384) );
  AND U7116 ( .A(n7387), .B(n7388), .Z(n7386) );
  NANDN U7117 ( .A(n7389), .B(n7390), .Z(n7388) );
  NANDN U7118 ( .A(n7391), .B(n7392), .Z(n7387) );
  NANDN U7119 ( .A(n7390), .B(n7389), .Z(n7392) );
  ANDN U7120 ( .B(\stack[0][9] ), .A(n6468), .Z(n7385) );
  XOR U7121 ( .A(n7393), .B(n7394), .Z(n7383) );
  AND U7122 ( .A(n7395), .B(n7396), .Z(n7394) );
  NANDN U7123 ( .A(n7397), .B(n7398), .Z(n7396) );
  NANDN U7124 ( .A(n7399), .B(n7400), .Z(n7395) );
  OR U7125 ( .A(n7398), .B(n7401), .Z(n7400) );
  ANDN U7126 ( .B(\stack[0][8] ), .A(n6492), .Z(n7393) );
  XOR U7127 ( .A(n7402), .B(n7403), .Z(n7287) );
  XOR U7128 ( .A(n7404), .B(n7405), .Z(n7403) );
  AND U7129 ( .A(n7406), .B(n7407), .Z(n7405) );
  NANDN U7130 ( .A(n7408), .B(n7409), .Z(n7407) );
  NANDN U7131 ( .A(n7410), .B(n7411), .Z(n7406) );
  OR U7132 ( .A(n7409), .B(n7412), .Z(n7411) );
  ANDN U7133 ( .B(\stack[1][51] ), .A(n5446), .Z(n7404) );
  XOR U7134 ( .A(n7413), .B(n7414), .Z(n7402) );
  AND U7135 ( .A(n7415), .B(n7416), .Z(n7414) );
  NANDN U7136 ( .A(n7417), .B(n7418), .Z(n7416) );
  NANDN U7137 ( .A(n7419), .B(n7420), .Z(n7415) );
  NANDN U7138 ( .A(n7418), .B(n7417), .Z(n7420) );
  ANDN U7139 ( .B(\stack[1][52] ), .A(n5422), .Z(n7413) );
  XOR U7140 ( .A(n7421), .B(n7422), .Z(n7275) );
  XOR U7141 ( .A(n7423), .B(n7424), .Z(n7422) );
  AND U7142 ( .A(n7425), .B(n7426), .Z(n7424) );
  NANDN U7143 ( .A(n7427), .B(n7428), .Z(n7426) );
  NANDN U7144 ( .A(n7429), .B(n7430), .Z(n7425) );
  NANDN U7145 ( .A(n7428), .B(n7427), .Z(n7430) );
  ANDN U7146 ( .B(\stack[1][48] ), .A(n5518), .Z(n7423) );
  XOR U7147 ( .A(n7431), .B(n7432), .Z(n7421) );
  AND U7148 ( .A(n7433), .B(n7434), .Z(n7432) );
  NANDN U7149 ( .A(n7435), .B(n7436), .Z(n7434) );
  NANDN U7150 ( .A(n7437), .B(n7438), .Z(n7433) );
  OR U7151 ( .A(n7436), .B(n7439), .Z(n7438) );
  ANDN U7152 ( .B(\stack[1][49] ), .A(n5494), .Z(n7431) );
  XOR U7153 ( .A(n7440), .B(n7441), .Z(n7262) );
  XOR U7154 ( .A(n7442), .B(n7443), .Z(n7441) );
  AND U7155 ( .A(n7444), .B(n7445), .Z(n7443) );
  NANDN U7156 ( .A(n7446), .B(n7447), .Z(n7445) );
  NANDN U7157 ( .A(n7448), .B(n7449), .Z(n7444) );
  OR U7158 ( .A(n7447), .B(n7450), .Z(n7449) );
  ANDN U7159 ( .B(\stack[1][45] ), .A(n5590), .Z(n7442) );
  XOR U7160 ( .A(n7451), .B(n7452), .Z(n7440) );
  AND U7161 ( .A(n7453), .B(n7454), .Z(n7452) );
  NANDN U7162 ( .A(n7455), .B(n7456), .Z(n7454) );
  NANDN U7163 ( .A(n7457), .B(n7458), .Z(n7453) );
  NANDN U7164 ( .A(n7456), .B(n7455), .Z(n7458) );
  ANDN U7165 ( .B(\stack[1][46] ), .A(n5566), .Z(n7451) );
  XOR U7166 ( .A(n7459), .B(n7460), .Z(n7248) );
  XOR U7167 ( .A(n7461), .B(n7462), .Z(n7460) );
  AND U7168 ( .A(n7463), .B(n7464), .Z(n7462) );
  NANDN U7169 ( .A(n7465), .B(n7466), .Z(n7464) );
  NANDN U7170 ( .A(n7467), .B(n7468), .Z(n7463) );
  NANDN U7171 ( .A(n7466), .B(n7465), .Z(n7468) );
  ANDN U7172 ( .B(\stack[1][42] ), .A(n5662), .Z(n7461) );
  XOR U7173 ( .A(n7469), .B(n7470), .Z(n7459) );
  AND U7174 ( .A(n7471), .B(n7472), .Z(n7470) );
  NANDN U7175 ( .A(n7473), .B(n7474), .Z(n7472) );
  NANDN U7176 ( .A(n7475), .B(n7476), .Z(n7471) );
  OR U7177 ( .A(n7474), .B(n7477), .Z(n7476) );
  ANDN U7178 ( .B(\stack[1][43] ), .A(n5638), .Z(n7469) );
  XOR U7179 ( .A(n7478), .B(n7479), .Z(n7236) );
  XOR U7180 ( .A(n7480), .B(n7481), .Z(n7479) );
  AND U7181 ( .A(n7482), .B(n7483), .Z(n7481) );
  NANDN U7182 ( .A(n7484), .B(n7485), .Z(n7483) );
  NANDN U7183 ( .A(n7486), .B(n7487), .Z(n7482) );
  OR U7184 ( .A(n7485), .B(n7488), .Z(n7487) );
  ANDN U7185 ( .B(\stack[1][39] ), .A(n5734), .Z(n7480) );
  XOR U7186 ( .A(n7489), .B(n7490), .Z(n7478) );
  AND U7187 ( .A(n7491), .B(n7492), .Z(n7490) );
  NANDN U7188 ( .A(n7493), .B(n7494), .Z(n7492) );
  NANDN U7189 ( .A(n7495), .B(n7496), .Z(n7491) );
  NANDN U7190 ( .A(n7494), .B(n7493), .Z(n7496) );
  ANDN U7191 ( .B(\stack[1][40] ), .A(n5710), .Z(n7489) );
  XOR U7192 ( .A(n7497), .B(n7498), .Z(n7224) );
  AND U7193 ( .A(n7499), .B(n7500), .Z(n7498) );
  NANDN U7194 ( .A(n7501), .B(n7502), .Z(n7500) );
  OR U7195 ( .A(n7503), .B(n7504), .Z(n7502) );
  AND U7196 ( .A(n7505), .B(n7506), .Z(n7497) );
  NANDN U7197 ( .A(n7507), .B(n7508), .Z(n7506) );
  NANDN U7198 ( .A(n7509), .B(n7510), .Z(n7505) );
  OR U7199 ( .A(n7508), .B(n7511), .Z(n7510) );
  XOR U7200 ( .A(n7512), .B(n7513), .Z(n7222) );
  XOR U7201 ( .A(n7514), .B(n7515), .Z(n7513) );
  ANDN U7202 ( .B(\stack[1][35] ), .A(n5830), .Z(n7515) );
  AND U7203 ( .A(n7516), .B(n7517), .Z(n7514) );
  NANDN U7204 ( .A(n7518), .B(n7519), .Z(n7517) );
  NANDN U7205 ( .A(n7520), .B(n7521), .Z(n7516) );
  NANDN U7206 ( .A(n7519), .B(n7518), .Z(n7521) );
  XOR U7207 ( .A(n7522), .B(n7523), .Z(n7512) );
  ANDN U7208 ( .B(\stack[1][36] ), .A(n5806), .Z(n7523) );
  ANDN U7209 ( .B(\stack[1][37] ), .A(n5782), .Z(n7522) );
  XOR U7210 ( .A(n7524), .B(n7525), .Z(n7210) );
  AND U7211 ( .A(n7526), .B(n7527), .Z(n7525) );
  NANDN U7212 ( .A(n7528), .B(n7529), .Z(n7527) );
  NANDN U7213 ( .A(n7530), .B(n7531), .Z(n7526) );
  OR U7214 ( .A(n7529), .B(n7532), .Z(n7531) );
  ANDN U7215 ( .B(\stack[1][31] ), .A(n5926), .Z(n7524) );
  XOR U7216 ( .A(n7533), .B(n7534), .Z(n7208) );
  XOR U7217 ( .A(n7535), .B(n7536), .Z(n7534) );
  AND U7218 ( .A(n7537), .B(n7538), .Z(n7536) );
  NANDN U7219 ( .A(n7539), .B(n7540), .Z(n7538) );
  NANDN U7220 ( .A(n7541), .B(n7542), .Z(n7537) );
  NANDN U7221 ( .A(n7540), .B(n7539), .Z(n7542) );
  ANDN U7222 ( .B(\stack[1][32] ), .A(n5902), .Z(n7535) );
  XOR U7223 ( .A(n7543), .B(n7544), .Z(n7533) );
  AND U7224 ( .A(n7545), .B(n7546), .Z(n7544) );
  NANDN U7225 ( .A(n7547), .B(n7548), .Z(n7546) );
  NANDN U7226 ( .A(n7549), .B(n7550), .Z(n7545) );
  OR U7227 ( .A(n7548), .B(n7551), .Z(n7550) );
  ANDN U7228 ( .B(\stack[1][33] ), .A(n5878), .Z(n7543) );
  XOR U7229 ( .A(n7552), .B(n7553), .Z(n7196) );
  AND U7230 ( .A(n7554), .B(n7555), .Z(n7553) );
  NANDN U7231 ( .A(n7556), .B(n7557), .Z(n7555) );
  NANDN U7232 ( .A(n7558), .B(n7559), .Z(n7554) );
  OR U7233 ( .A(n7557), .B(n7560), .Z(n7559) );
  ANDN U7234 ( .B(\stack[1][27] ), .A(n6022), .Z(n7552) );
  XOR U7235 ( .A(n7561), .B(n7562), .Z(n7194) );
  XOR U7236 ( .A(n7563), .B(n7564), .Z(n7562) );
  AND U7237 ( .A(n7565), .B(n7566), .Z(n7564) );
  NANDN U7238 ( .A(n7567), .B(n7568), .Z(n7566) );
  NANDN U7239 ( .A(n7569), .B(n7570), .Z(n7565) );
  NANDN U7240 ( .A(n7568), .B(n7567), .Z(n7570) );
  ANDN U7241 ( .B(\stack[1][28] ), .A(n5998), .Z(n7563) );
  XOR U7242 ( .A(n7571), .B(n7572), .Z(n7561) );
  AND U7243 ( .A(n7573), .B(n7574), .Z(n7572) );
  NANDN U7244 ( .A(n7575), .B(n7576), .Z(n7574) );
  NANDN U7245 ( .A(n7577), .B(n7578), .Z(n7573) );
  OR U7246 ( .A(n7576), .B(n7579), .Z(n7578) );
  ANDN U7247 ( .B(\stack[1][29] ), .A(n5974), .Z(n7571) );
  XOR U7248 ( .A(n7580), .B(n7581), .Z(n7182) );
  AND U7249 ( .A(n7582), .B(n7583), .Z(n7581) );
  NANDN U7250 ( .A(n7584), .B(n7585), .Z(n7583) );
  NANDN U7251 ( .A(n7586), .B(n7587), .Z(n7582) );
  OR U7252 ( .A(n7585), .B(n7588), .Z(n7587) );
  ANDN U7253 ( .B(\stack[1][23] ), .A(n6118), .Z(n7580) );
  XOR U7254 ( .A(n7589), .B(n7590), .Z(n7180) );
  XOR U7255 ( .A(n7591), .B(n7592), .Z(n7590) );
  AND U7256 ( .A(n7593), .B(n7594), .Z(n7592) );
  NANDN U7257 ( .A(n7595), .B(n7596), .Z(n7594) );
  NANDN U7258 ( .A(n7597), .B(n7598), .Z(n7593) );
  NANDN U7259 ( .A(n7596), .B(n7595), .Z(n7598) );
  ANDN U7260 ( .B(\stack[1][24] ), .A(n6094), .Z(n7591) );
  XOR U7261 ( .A(n7599), .B(n7600), .Z(n7589) );
  AND U7262 ( .A(n7601), .B(n7602), .Z(n7600) );
  NANDN U7263 ( .A(n7603), .B(n7604), .Z(n7602) );
  NANDN U7264 ( .A(n7605), .B(n7606), .Z(n7601) );
  OR U7265 ( .A(n7604), .B(n7607), .Z(n7606) );
  ANDN U7266 ( .B(\stack[1][25] ), .A(n6070), .Z(n7599) );
  XOR U7267 ( .A(n7608), .B(n7609), .Z(n7168) );
  AND U7268 ( .A(n7610), .B(n7611), .Z(n7609) );
  NANDN U7269 ( .A(n7612), .B(n7613), .Z(n7611) );
  NANDN U7270 ( .A(n7614), .B(n7615), .Z(n7610) );
  OR U7271 ( .A(n7613), .B(n7616), .Z(n7615) );
  ANDN U7272 ( .B(\stack[1][19] ), .A(n6214), .Z(n7608) );
  XOR U7273 ( .A(n7617), .B(n7618), .Z(n7166) );
  XOR U7274 ( .A(n7619), .B(n7620), .Z(n7618) );
  AND U7275 ( .A(n7621), .B(n7622), .Z(n7620) );
  NANDN U7276 ( .A(n7623), .B(n7624), .Z(n7622) );
  NANDN U7277 ( .A(n7625), .B(n7626), .Z(n7621) );
  NANDN U7278 ( .A(n7624), .B(n7623), .Z(n7626) );
  ANDN U7279 ( .B(\stack[1][20] ), .A(n6190), .Z(n7619) );
  XOR U7280 ( .A(n7627), .B(n7628), .Z(n7617) );
  AND U7281 ( .A(n7629), .B(n7630), .Z(n7628) );
  NANDN U7282 ( .A(n7631), .B(n7632), .Z(n7630) );
  NANDN U7283 ( .A(n7633), .B(n7634), .Z(n7629) );
  OR U7284 ( .A(n7632), .B(n7635), .Z(n7634) );
  ANDN U7285 ( .B(\stack[1][21] ), .A(n6166), .Z(n7627) );
  XOR U7286 ( .A(n7636), .B(n7637), .Z(n7154) );
  AND U7287 ( .A(n7638), .B(n7639), .Z(n7637) );
  NANDN U7288 ( .A(n7640), .B(n7641), .Z(n7639) );
  NANDN U7289 ( .A(n7642), .B(n7643), .Z(n7638) );
  OR U7290 ( .A(n7641), .B(n7644), .Z(n7643) );
  ANDN U7291 ( .B(\stack[1][15] ), .A(n6310), .Z(n7636) );
  XOR U7292 ( .A(n7645), .B(n7646), .Z(n7152) );
  XOR U7293 ( .A(n7647), .B(n7648), .Z(n7646) );
  AND U7294 ( .A(n7649), .B(n7650), .Z(n7648) );
  NANDN U7295 ( .A(n7651), .B(n7652), .Z(n7650) );
  NANDN U7296 ( .A(n7653), .B(n7654), .Z(n7649) );
  NANDN U7297 ( .A(n7652), .B(n7651), .Z(n7654) );
  ANDN U7298 ( .B(\stack[1][16] ), .A(n6286), .Z(n7647) );
  XOR U7299 ( .A(n7655), .B(n7656), .Z(n7645) );
  AND U7300 ( .A(n7657), .B(n7658), .Z(n7656) );
  NANDN U7301 ( .A(n7659), .B(n7660), .Z(n7658) );
  NANDN U7302 ( .A(n7661), .B(n7662), .Z(n7657) );
  OR U7303 ( .A(n7660), .B(n7663), .Z(n7662) );
  ANDN U7304 ( .B(\stack[1][17] ), .A(n6262), .Z(n7655) );
  XOR U7305 ( .A(n7664), .B(n7665), .Z(n7139) );
  AND U7306 ( .A(n7666), .B(n7667), .Z(n7665) );
  NANDN U7307 ( .A(n7668), .B(n7669), .Z(n7667) );
  NANDN U7308 ( .A(n7670), .B(n7671), .Z(n7666) );
  OR U7309 ( .A(n7669), .B(n7672), .Z(n7671) );
  ANDN U7310 ( .B(\stack[1][11] ), .A(n6406), .Z(n7664) );
  XOR U7311 ( .A(n7673), .B(n7674), .Z(n7137) );
  XOR U7312 ( .A(n7675), .B(n7676), .Z(n7674) );
  AND U7313 ( .A(n7677), .B(n7678), .Z(n7676) );
  NANDN U7314 ( .A(n7679), .B(n7680), .Z(n7678) );
  NANDN U7315 ( .A(n7681), .B(n7682), .Z(n7677) );
  NANDN U7316 ( .A(n7680), .B(n7679), .Z(n7682) );
  ANDN U7317 ( .B(\stack[1][12] ), .A(n6382), .Z(n7675) );
  XOR U7318 ( .A(n7683), .B(n7684), .Z(n7673) );
  AND U7319 ( .A(n7685), .B(n7686), .Z(n7684) );
  NANDN U7320 ( .A(n7687), .B(n7688), .Z(n7686) );
  NANDN U7321 ( .A(n7689), .B(n7690), .Z(n7685) );
  OR U7322 ( .A(n7688), .B(n7691), .Z(n7690) );
  ANDN U7323 ( .B(\stack[1][13] ), .A(n6358), .Z(n7683) );
  XOR U7324 ( .A(n7692), .B(n7693), .Z(n7125) );
  AND U7325 ( .A(n7694), .B(n7695), .Z(n7693) );
  NANDN U7326 ( .A(n7696), .B(n7697), .Z(n7695) );
  NANDN U7327 ( .A(n7698), .B(n7699), .Z(n7694) );
  OR U7328 ( .A(n7697), .B(n7700), .Z(n7699) );
  ANDN U7329 ( .B(\stack[1][7] ), .A(n6502), .Z(n7692) );
  XOR U7330 ( .A(n7701), .B(n7702), .Z(n7123) );
  XOR U7331 ( .A(n7703), .B(n7704), .Z(n7702) );
  AND U7332 ( .A(n7705), .B(n7706), .Z(n7704) );
  NANDN U7333 ( .A(n7707), .B(n7708), .Z(n7706) );
  NANDN U7334 ( .A(n7709), .B(n7710), .Z(n7705) );
  NANDN U7335 ( .A(n7708), .B(n7707), .Z(n7710) );
  ANDN U7336 ( .B(\stack[1][8] ), .A(n6478), .Z(n7703) );
  XOR U7337 ( .A(n7711), .B(n7712), .Z(n7701) );
  AND U7338 ( .A(n7713), .B(n7714), .Z(n7712) );
  NANDN U7339 ( .A(n7715), .B(n7716), .Z(n7714) );
  NANDN U7340 ( .A(n7717), .B(n7718), .Z(n7713) );
  OR U7341 ( .A(n7716), .B(n7719), .Z(n7718) );
  ANDN U7342 ( .B(\stack[1][9] ), .A(n6454), .Z(n7711) );
  AND U7343 ( .A(n7720), .B(n7721), .Z(n7121) );
  NANDN U7344 ( .A(n7113), .B(n7115), .Z(n7721) );
  NANDN U7345 ( .A(n7116), .B(n7722), .Z(n7720) );
  NANDN U7346 ( .A(n7115), .B(n7113), .Z(n7722) );
  XOR U7347 ( .A(n7133), .B(n7723), .Z(n7113) );
  XNOR U7348 ( .A(n7134), .B(n7135), .Z(n7723) );
  AND U7349 ( .A(n7724), .B(n7725), .Z(n7135) );
  NAND U7350 ( .A(n7726), .B(n7727), .Z(n7725) );
  NANDN U7351 ( .A(n7728), .B(n7729), .Z(n7724) );
  OR U7352 ( .A(n7726), .B(n7727), .Z(n7729) );
  AND U7353 ( .A(\stack[1][2] ), .B(\stack[0][60] ), .Z(n7134) );
  XOR U7354 ( .A(n7730), .B(n7731), .Z(n7133) );
  XNOR U7355 ( .A(n7732), .B(n7733), .Z(n7731) );
  ANDN U7356 ( .B(\stack[0][61] ), .A(n5195), .Z(n7115) );
  AND U7357 ( .A(n7734), .B(n7735), .Z(n7116) );
  NANDN U7358 ( .A(n7110), .B(n7736), .Z(n7734) );
  NANDN U7359 ( .A(n7109), .B(n7107), .Z(n7736) );
  XNOR U7360 ( .A(n7726), .B(n7737), .Z(n7107) );
  XNOR U7361 ( .A(n7727), .B(n7728), .Z(n7737) );
  AND U7362 ( .A(n7738), .B(n7739), .Z(n7728) );
  NANDN U7363 ( .A(n7740), .B(n7741), .Z(n7739) );
  NANDN U7364 ( .A(n7742), .B(n7743), .Z(n7738) );
  NANDN U7365 ( .A(n7741), .B(n7740), .Z(n7743) );
  ANDN U7366 ( .B(\stack[0][59] ), .A(n5219), .Z(n7727) );
  XNOR U7367 ( .A(n7744), .B(n7745), .Z(n7726) );
  XNOR U7368 ( .A(n7746), .B(n7747), .Z(n7745) );
  ANDN U7369 ( .B(\stack[1][1] ), .A(n6598), .Z(n7109) );
  AND U7370 ( .A(n7748), .B(n7749), .Z(n7110) );
  NANDN U7371 ( .A(n7103), .B(n7105), .Z(n7749) );
  NANDN U7372 ( .A(n7106), .B(n7750), .Z(n7748) );
  NANDN U7373 ( .A(n7105), .B(n7103), .Z(n7750) );
  XOR U7374 ( .A(n7740), .B(n7751), .Z(n7103) );
  XNOR U7375 ( .A(n7741), .B(n7742), .Z(n7751) );
  AND U7376 ( .A(n7752), .B(n7753), .Z(n7742) );
  NAND U7377 ( .A(n7754), .B(n7755), .Z(n7753) );
  NANDN U7378 ( .A(n7756), .B(n7757), .Z(n7752) );
  OR U7379 ( .A(n7754), .B(n7755), .Z(n7757) );
  ANDN U7380 ( .B(\stack[0][58] ), .A(n5219), .Z(n7741) );
  XOR U7381 ( .A(n7758), .B(n7759), .Z(n7740) );
  XNOR U7382 ( .A(n7760), .B(n7761), .Z(n7759) );
  ANDN U7383 ( .B(\stack[0][59] ), .A(n5195), .Z(n7105) );
  AND U7384 ( .A(n7762), .B(n7763), .Z(n7106) );
  NANDN U7385 ( .A(n7102), .B(n7764), .Z(n7762) );
  NANDN U7386 ( .A(n7101), .B(n7099), .Z(n7764) );
  XNOR U7387 ( .A(n7754), .B(n7765), .Z(n7099) );
  XNOR U7388 ( .A(n7755), .B(n7756), .Z(n7765) );
  AND U7389 ( .A(n7766), .B(n7767), .Z(n7756) );
  NANDN U7390 ( .A(n7768), .B(n7769), .Z(n7767) );
  NANDN U7391 ( .A(n7770), .B(n7771), .Z(n7766) );
  NANDN U7392 ( .A(n7769), .B(n7768), .Z(n7771) );
  ANDN U7393 ( .B(\stack[0][57] ), .A(n5219), .Z(n7755) );
  XNOR U7394 ( .A(n7772), .B(n7773), .Z(n7754) );
  XNOR U7395 ( .A(n7774), .B(n7775), .Z(n7773) );
  ANDN U7396 ( .B(\stack[1][1] ), .A(n6550), .Z(n7101) );
  AND U7397 ( .A(n7776), .B(n7777), .Z(n7102) );
  NANDN U7398 ( .A(n7095), .B(n7097), .Z(n7777) );
  NANDN U7399 ( .A(n7098), .B(n7778), .Z(n7776) );
  NANDN U7400 ( .A(n7097), .B(n7095), .Z(n7778) );
  XOR U7401 ( .A(n7768), .B(n7779), .Z(n7095) );
  XNOR U7402 ( .A(n7769), .B(n7770), .Z(n7779) );
  AND U7403 ( .A(n7780), .B(n7781), .Z(n7770) );
  NAND U7404 ( .A(n7782), .B(n7783), .Z(n7781) );
  NANDN U7405 ( .A(n7784), .B(n7785), .Z(n7780) );
  OR U7406 ( .A(n7782), .B(n7783), .Z(n7785) );
  ANDN U7407 ( .B(\stack[0][56] ), .A(n5219), .Z(n7769) );
  XOR U7408 ( .A(n7786), .B(n7787), .Z(n7768) );
  XNOR U7409 ( .A(n7788), .B(n7789), .Z(n7787) );
  ANDN U7410 ( .B(\stack[0][57] ), .A(n5195), .Z(n7097) );
  AND U7411 ( .A(n7790), .B(n7791), .Z(n7098) );
  NANDN U7412 ( .A(n7094), .B(n7792), .Z(n7790) );
  NANDN U7413 ( .A(n7093), .B(n7091), .Z(n7792) );
  XNOR U7414 ( .A(n7782), .B(n7793), .Z(n7091) );
  XNOR U7415 ( .A(n7783), .B(n7784), .Z(n7793) );
  AND U7416 ( .A(n7794), .B(n7795), .Z(n7784) );
  NANDN U7417 ( .A(n7796), .B(n7797), .Z(n7795) );
  NANDN U7418 ( .A(n7798), .B(n7799), .Z(n7794) );
  NANDN U7419 ( .A(n7797), .B(n7796), .Z(n7799) );
  ANDN U7420 ( .B(\stack[0][55] ), .A(n5219), .Z(n7783) );
  XNOR U7421 ( .A(n7800), .B(n7801), .Z(n7782) );
  XNOR U7422 ( .A(n7802), .B(n7803), .Z(n7801) );
  ANDN U7423 ( .B(\stack[1][1] ), .A(n6502), .Z(n7093) );
  AND U7424 ( .A(n7804), .B(n7805), .Z(n7094) );
  NANDN U7425 ( .A(n7087), .B(n7089), .Z(n7805) );
  NANDN U7426 ( .A(n7090), .B(n7806), .Z(n7804) );
  NANDN U7427 ( .A(n7089), .B(n7087), .Z(n7806) );
  XOR U7428 ( .A(n7796), .B(n7807), .Z(n7087) );
  XNOR U7429 ( .A(n7797), .B(n7798), .Z(n7807) );
  AND U7430 ( .A(n7808), .B(n7809), .Z(n7798) );
  NAND U7431 ( .A(n7810), .B(n7811), .Z(n7809) );
  NANDN U7432 ( .A(n7812), .B(n7813), .Z(n7808) );
  OR U7433 ( .A(n7810), .B(n7811), .Z(n7813) );
  ANDN U7434 ( .B(\stack[0][54] ), .A(n5219), .Z(n7797) );
  XOR U7435 ( .A(n7814), .B(n7815), .Z(n7796) );
  XNOR U7436 ( .A(n7816), .B(n7817), .Z(n7815) );
  ANDN U7437 ( .B(\stack[0][55] ), .A(n5195), .Z(n7089) );
  AND U7438 ( .A(n7818), .B(n7819), .Z(n7090) );
  NANDN U7439 ( .A(n7086), .B(n7820), .Z(n7818) );
  NANDN U7440 ( .A(n7085), .B(n7083), .Z(n7820) );
  XNOR U7441 ( .A(n7810), .B(n7821), .Z(n7083) );
  XNOR U7442 ( .A(n7811), .B(n7812), .Z(n7821) );
  AND U7443 ( .A(n7822), .B(n7823), .Z(n7812) );
  NANDN U7444 ( .A(n7824), .B(n7825), .Z(n7823) );
  NANDN U7445 ( .A(n7826), .B(n7827), .Z(n7822) );
  NANDN U7446 ( .A(n7825), .B(n7824), .Z(n7827) );
  ANDN U7447 ( .B(\stack[0][53] ), .A(n5219), .Z(n7811) );
  XNOR U7448 ( .A(n7828), .B(n7829), .Z(n7810) );
  XNOR U7449 ( .A(n7830), .B(n7831), .Z(n7829) );
  ANDN U7450 ( .B(\stack[1][1] ), .A(n6454), .Z(n7085) );
  AND U7451 ( .A(n7832), .B(n7833), .Z(n7086) );
  NANDN U7452 ( .A(n7079), .B(n7081), .Z(n7833) );
  NANDN U7453 ( .A(n7082), .B(n7834), .Z(n7832) );
  NANDN U7454 ( .A(n7081), .B(n7079), .Z(n7834) );
  XOR U7455 ( .A(n7824), .B(n7835), .Z(n7079) );
  XNOR U7456 ( .A(n7825), .B(n7826), .Z(n7835) );
  AND U7457 ( .A(n7836), .B(n7837), .Z(n7826) );
  NAND U7458 ( .A(n7838), .B(n7839), .Z(n7837) );
  NANDN U7459 ( .A(n7840), .B(n7841), .Z(n7836) );
  OR U7460 ( .A(n7838), .B(n7839), .Z(n7841) );
  ANDN U7461 ( .B(\stack[0][52] ), .A(n5219), .Z(n7825) );
  XOR U7462 ( .A(n7842), .B(n7843), .Z(n7824) );
  XNOR U7463 ( .A(n7844), .B(n7845), .Z(n7843) );
  ANDN U7464 ( .B(\stack[0][53] ), .A(n5195), .Z(n7081) );
  AND U7465 ( .A(n7846), .B(n7847), .Z(n7082) );
  NANDN U7466 ( .A(n7078), .B(n7848), .Z(n7846) );
  NANDN U7467 ( .A(n7077), .B(n7075), .Z(n7848) );
  XNOR U7468 ( .A(n7838), .B(n7849), .Z(n7075) );
  XNOR U7469 ( .A(n7839), .B(n7840), .Z(n7849) );
  AND U7470 ( .A(n7850), .B(n7851), .Z(n7840) );
  NANDN U7471 ( .A(n7852), .B(n7853), .Z(n7851) );
  NANDN U7472 ( .A(n7854), .B(n7855), .Z(n7850) );
  NANDN U7473 ( .A(n7853), .B(n7852), .Z(n7855) );
  ANDN U7474 ( .B(\stack[0][51] ), .A(n5219), .Z(n7839) );
  XNOR U7475 ( .A(n7856), .B(n7857), .Z(n7838) );
  XNOR U7476 ( .A(n7858), .B(n7859), .Z(n7857) );
  ANDN U7477 ( .B(\stack[1][1] ), .A(n6406), .Z(n7077) );
  AND U7478 ( .A(n7860), .B(n7861), .Z(n7078) );
  NANDN U7479 ( .A(n7071), .B(n7073), .Z(n7861) );
  NANDN U7480 ( .A(n7074), .B(n7862), .Z(n7860) );
  NANDN U7481 ( .A(n7073), .B(n7071), .Z(n7862) );
  XOR U7482 ( .A(n7852), .B(n7863), .Z(n7071) );
  XNOR U7483 ( .A(n7853), .B(n7854), .Z(n7863) );
  AND U7484 ( .A(n7864), .B(n7865), .Z(n7854) );
  NAND U7485 ( .A(n7866), .B(n7867), .Z(n7865) );
  NANDN U7486 ( .A(n7868), .B(n7869), .Z(n7864) );
  OR U7487 ( .A(n7866), .B(n7867), .Z(n7869) );
  ANDN U7488 ( .B(\stack[0][50] ), .A(n5219), .Z(n7853) );
  XOR U7489 ( .A(n7870), .B(n7871), .Z(n7852) );
  XNOR U7490 ( .A(n7872), .B(n7873), .Z(n7871) );
  ANDN U7491 ( .B(\stack[0][51] ), .A(n5195), .Z(n7073) );
  AND U7492 ( .A(n7874), .B(n7875), .Z(n7074) );
  NANDN U7493 ( .A(n7070), .B(n7876), .Z(n7874) );
  NANDN U7494 ( .A(n7069), .B(n7067), .Z(n7876) );
  XNOR U7495 ( .A(n7866), .B(n7877), .Z(n7067) );
  XNOR U7496 ( .A(n7867), .B(n7868), .Z(n7877) );
  AND U7497 ( .A(n7878), .B(n7879), .Z(n7868) );
  NANDN U7498 ( .A(n7880), .B(n7881), .Z(n7879) );
  NANDN U7499 ( .A(n7882), .B(n7883), .Z(n7878) );
  NANDN U7500 ( .A(n7881), .B(n7880), .Z(n7883) );
  ANDN U7501 ( .B(\stack[0][49] ), .A(n5219), .Z(n7867) );
  XNOR U7502 ( .A(n7884), .B(n7885), .Z(n7866) );
  XNOR U7503 ( .A(n7886), .B(n7887), .Z(n7885) );
  ANDN U7504 ( .B(\stack[1][1] ), .A(n6358), .Z(n7069) );
  AND U7505 ( .A(n7888), .B(n7889), .Z(n7070) );
  NANDN U7506 ( .A(n7063), .B(n7065), .Z(n7889) );
  NANDN U7507 ( .A(n7066), .B(n7890), .Z(n7888) );
  NANDN U7508 ( .A(n7065), .B(n7063), .Z(n7890) );
  XOR U7509 ( .A(n7880), .B(n7891), .Z(n7063) );
  XNOR U7510 ( .A(n7881), .B(n7882), .Z(n7891) );
  AND U7511 ( .A(n7892), .B(n7893), .Z(n7882) );
  NAND U7512 ( .A(n7894), .B(n7895), .Z(n7893) );
  NANDN U7513 ( .A(n7896), .B(n7897), .Z(n7892) );
  OR U7514 ( .A(n7894), .B(n7895), .Z(n7897) );
  ANDN U7515 ( .B(\stack[0][48] ), .A(n5219), .Z(n7881) );
  XOR U7516 ( .A(n7898), .B(n7899), .Z(n7880) );
  XNOR U7517 ( .A(n7900), .B(n7901), .Z(n7899) );
  ANDN U7518 ( .B(\stack[0][49] ), .A(n5195), .Z(n7065) );
  AND U7519 ( .A(n7902), .B(n7903), .Z(n7066) );
  NANDN U7520 ( .A(n7062), .B(n7904), .Z(n7902) );
  NANDN U7521 ( .A(n7061), .B(n7059), .Z(n7904) );
  XNOR U7522 ( .A(n7894), .B(n7905), .Z(n7059) );
  XNOR U7523 ( .A(n7895), .B(n7896), .Z(n7905) );
  AND U7524 ( .A(n7906), .B(n7907), .Z(n7896) );
  NANDN U7525 ( .A(n7908), .B(n7909), .Z(n7907) );
  NANDN U7526 ( .A(n7910), .B(n7911), .Z(n7906) );
  NANDN U7527 ( .A(n7909), .B(n7908), .Z(n7911) );
  ANDN U7528 ( .B(\stack[0][47] ), .A(n5219), .Z(n7895) );
  XNOR U7529 ( .A(n7912), .B(n7913), .Z(n7894) );
  XNOR U7530 ( .A(n7914), .B(n7915), .Z(n7913) );
  ANDN U7531 ( .B(\stack[1][1] ), .A(n6310), .Z(n7061) );
  AND U7532 ( .A(n7916), .B(n7917), .Z(n7062) );
  NANDN U7533 ( .A(n7055), .B(n7057), .Z(n7917) );
  NANDN U7534 ( .A(n7058), .B(n7918), .Z(n7916) );
  NANDN U7535 ( .A(n7057), .B(n7055), .Z(n7918) );
  XOR U7536 ( .A(n7908), .B(n7919), .Z(n7055) );
  XNOR U7537 ( .A(n7909), .B(n7910), .Z(n7919) );
  AND U7538 ( .A(n7920), .B(n7921), .Z(n7910) );
  NAND U7539 ( .A(n7922), .B(n7923), .Z(n7921) );
  NANDN U7540 ( .A(n7924), .B(n7925), .Z(n7920) );
  OR U7541 ( .A(n7922), .B(n7923), .Z(n7925) );
  ANDN U7542 ( .B(\stack[0][46] ), .A(n5219), .Z(n7909) );
  XOR U7543 ( .A(n7926), .B(n7927), .Z(n7908) );
  XNOR U7544 ( .A(n7928), .B(n7929), .Z(n7927) );
  ANDN U7545 ( .B(\stack[0][47] ), .A(n5195), .Z(n7057) );
  AND U7546 ( .A(n7930), .B(n7931), .Z(n7058) );
  NANDN U7547 ( .A(n7054), .B(n7932), .Z(n7930) );
  NANDN U7548 ( .A(n7053), .B(n7051), .Z(n7932) );
  XNOR U7549 ( .A(n7922), .B(n7933), .Z(n7051) );
  XNOR U7550 ( .A(n7923), .B(n7924), .Z(n7933) );
  AND U7551 ( .A(n7934), .B(n7935), .Z(n7924) );
  NANDN U7552 ( .A(n7936), .B(n7937), .Z(n7935) );
  NANDN U7553 ( .A(n7938), .B(n7939), .Z(n7934) );
  NANDN U7554 ( .A(n7937), .B(n7936), .Z(n7939) );
  ANDN U7555 ( .B(\stack[0][45] ), .A(n5219), .Z(n7923) );
  XNOR U7556 ( .A(n7940), .B(n7941), .Z(n7922) );
  XNOR U7557 ( .A(n7942), .B(n7943), .Z(n7941) );
  ANDN U7558 ( .B(\stack[1][1] ), .A(n6262), .Z(n7053) );
  AND U7559 ( .A(n7944), .B(n7945), .Z(n7054) );
  NANDN U7560 ( .A(n7047), .B(n7049), .Z(n7945) );
  NANDN U7561 ( .A(n7050), .B(n7946), .Z(n7944) );
  NANDN U7562 ( .A(n7049), .B(n7047), .Z(n7946) );
  XOR U7563 ( .A(n7936), .B(n7947), .Z(n7047) );
  XNOR U7564 ( .A(n7937), .B(n7938), .Z(n7947) );
  AND U7565 ( .A(n7948), .B(n7949), .Z(n7938) );
  NAND U7566 ( .A(n7950), .B(n7951), .Z(n7949) );
  NANDN U7567 ( .A(n7952), .B(n7953), .Z(n7948) );
  OR U7568 ( .A(n7950), .B(n7951), .Z(n7953) );
  ANDN U7569 ( .B(\stack[0][44] ), .A(n5219), .Z(n7937) );
  XOR U7570 ( .A(n7954), .B(n7955), .Z(n7936) );
  XNOR U7571 ( .A(n7956), .B(n7957), .Z(n7955) );
  ANDN U7572 ( .B(\stack[0][45] ), .A(n5195), .Z(n7049) );
  AND U7573 ( .A(n7958), .B(n7959), .Z(n7050) );
  NANDN U7574 ( .A(n7046), .B(n7960), .Z(n7958) );
  NANDN U7575 ( .A(n7045), .B(n7043), .Z(n7960) );
  XNOR U7576 ( .A(n7950), .B(n7961), .Z(n7043) );
  XNOR U7577 ( .A(n7951), .B(n7952), .Z(n7961) );
  AND U7578 ( .A(n7962), .B(n7963), .Z(n7952) );
  NANDN U7579 ( .A(n7964), .B(n7965), .Z(n7963) );
  NANDN U7580 ( .A(n7966), .B(n7967), .Z(n7962) );
  NANDN U7581 ( .A(n7965), .B(n7964), .Z(n7967) );
  ANDN U7582 ( .B(\stack[0][43] ), .A(n5219), .Z(n7951) );
  XNOR U7583 ( .A(n7968), .B(n7969), .Z(n7950) );
  XNOR U7584 ( .A(n7970), .B(n7971), .Z(n7969) );
  ANDN U7585 ( .B(\stack[1][1] ), .A(n6214), .Z(n7045) );
  AND U7586 ( .A(n7972), .B(n7973), .Z(n7046) );
  NANDN U7587 ( .A(n7039), .B(n7041), .Z(n7973) );
  NANDN U7588 ( .A(n7042), .B(n7974), .Z(n7972) );
  NANDN U7589 ( .A(n7041), .B(n7039), .Z(n7974) );
  XOR U7590 ( .A(n7964), .B(n7975), .Z(n7039) );
  XNOR U7591 ( .A(n7965), .B(n7966), .Z(n7975) );
  AND U7592 ( .A(n7976), .B(n7977), .Z(n7966) );
  NAND U7593 ( .A(n7978), .B(n7979), .Z(n7977) );
  NANDN U7594 ( .A(n7980), .B(n7981), .Z(n7976) );
  OR U7595 ( .A(n7978), .B(n7979), .Z(n7981) );
  ANDN U7596 ( .B(\stack[0][42] ), .A(n5219), .Z(n7965) );
  XOR U7597 ( .A(n7982), .B(n7983), .Z(n7964) );
  XNOR U7598 ( .A(n7984), .B(n7985), .Z(n7983) );
  ANDN U7599 ( .B(\stack[0][43] ), .A(n5195), .Z(n7041) );
  AND U7600 ( .A(n7986), .B(n7987), .Z(n7042) );
  NANDN U7601 ( .A(n7038), .B(n7988), .Z(n7986) );
  NANDN U7602 ( .A(n7037), .B(n7035), .Z(n7988) );
  XNOR U7603 ( .A(n7978), .B(n7989), .Z(n7035) );
  XNOR U7604 ( .A(n7979), .B(n7980), .Z(n7989) );
  AND U7605 ( .A(n7990), .B(n7991), .Z(n7980) );
  NANDN U7606 ( .A(n7992), .B(n7993), .Z(n7991) );
  NANDN U7607 ( .A(n7994), .B(n7995), .Z(n7990) );
  NANDN U7608 ( .A(n7993), .B(n7992), .Z(n7995) );
  ANDN U7609 ( .B(\stack[0][41] ), .A(n5219), .Z(n7979) );
  XNOR U7610 ( .A(n7996), .B(n7997), .Z(n7978) );
  XNOR U7611 ( .A(n7998), .B(n7999), .Z(n7997) );
  ANDN U7612 ( .B(\stack[1][1] ), .A(n6166), .Z(n7037) );
  AND U7613 ( .A(n8000), .B(n8001), .Z(n7038) );
  NANDN U7614 ( .A(n7031), .B(n7033), .Z(n8001) );
  NANDN U7615 ( .A(n7034), .B(n8002), .Z(n8000) );
  NANDN U7616 ( .A(n7033), .B(n7031), .Z(n8002) );
  XOR U7617 ( .A(n7992), .B(n8003), .Z(n7031) );
  XNOR U7618 ( .A(n7993), .B(n7994), .Z(n8003) );
  AND U7619 ( .A(n8004), .B(n8005), .Z(n7994) );
  NAND U7620 ( .A(n8006), .B(n8007), .Z(n8005) );
  NANDN U7621 ( .A(n8008), .B(n8009), .Z(n8004) );
  OR U7622 ( .A(n8006), .B(n8007), .Z(n8009) );
  ANDN U7623 ( .B(\stack[0][40] ), .A(n5219), .Z(n7993) );
  XOR U7624 ( .A(n8010), .B(n8011), .Z(n7992) );
  XNOR U7625 ( .A(n8012), .B(n8013), .Z(n8011) );
  ANDN U7626 ( .B(\stack[0][41] ), .A(n5195), .Z(n7033) );
  AND U7627 ( .A(n8014), .B(n8015), .Z(n7034) );
  NANDN U7628 ( .A(n7030), .B(n8016), .Z(n8014) );
  NANDN U7629 ( .A(n7029), .B(n7027), .Z(n8016) );
  XNOR U7630 ( .A(n8006), .B(n8017), .Z(n7027) );
  XNOR U7631 ( .A(n8007), .B(n8008), .Z(n8017) );
  AND U7632 ( .A(n8018), .B(n8019), .Z(n8008) );
  NANDN U7633 ( .A(n8020), .B(n8021), .Z(n8019) );
  NANDN U7634 ( .A(n8022), .B(n8023), .Z(n8018) );
  NANDN U7635 ( .A(n8021), .B(n8020), .Z(n8023) );
  ANDN U7636 ( .B(\stack[0][39] ), .A(n5219), .Z(n8007) );
  XNOR U7637 ( .A(n8024), .B(n8025), .Z(n8006) );
  XNOR U7638 ( .A(n8026), .B(n8027), .Z(n8025) );
  ANDN U7639 ( .B(\stack[1][1] ), .A(n6118), .Z(n7029) );
  AND U7640 ( .A(n8028), .B(n8029), .Z(n7030) );
  NANDN U7641 ( .A(n7023), .B(n7025), .Z(n8029) );
  NANDN U7642 ( .A(n7026), .B(n8030), .Z(n8028) );
  NANDN U7643 ( .A(n7025), .B(n7023), .Z(n8030) );
  XOR U7644 ( .A(n8020), .B(n8031), .Z(n7023) );
  XNOR U7645 ( .A(n8021), .B(n8022), .Z(n8031) );
  AND U7646 ( .A(n8032), .B(n8033), .Z(n8022) );
  NAND U7647 ( .A(n8034), .B(n8035), .Z(n8033) );
  NANDN U7648 ( .A(n8036), .B(n8037), .Z(n8032) );
  OR U7649 ( .A(n8034), .B(n8035), .Z(n8037) );
  ANDN U7650 ( .B(\stack[0][38] ), .A(n5219), .Z(n8021) );
  XOR U7651 ( .A(n8038), .B(n8039), .Z(n8020) );
  XNOR U7652 ( .A(n8040), .B(n8041), .Z(n8039) );
  ANDN U7653 ( .B(\stack[0][39] ), .A(n5195), .Z(n7025) );
  AND U7654 ( .A(n8042), .B(n8043), .Z(n7026) );
  NANDN U7655 ( .A(n7022), .B(n8044), .Z(n8042) );
  NANDN U7656 ( .A(n7021), .B(n7019), .Z(n8044) );
  XNOR U7657 ( .A(n8034), .B(n8045), .Z(n7019) );
  XNOR U7658 ( .A(n8035), .B(n8036), .Z(n8045) );
  AND U7659 ( .A(n8046), .B(n8047), .Z(n8036) );
  NANDN U7660 ( .A(n8048), .B(n8049), .Z(n8047) );
  NANDN U7661 ( .A(n8050), .B(n8051), .Z(n8046) );
  NANDN U7662 ( .A(n8049), .B(n8048), .Z(n8051) );
  ANDN U7663 ( .B(\stack[0][37] ), .A(n5219), .Z(n8035) );
  XNOR U7664 ( .A(n8052), .B(n8053), .Z(n8034) );
  XNOR U7665 ( .A(n8054), .B(n8055), .Z(n8053) );
  ANDN U7666 ( .B(\stack[1][1] ), .A(n6070), .Z(n7021) );
  AND U7667 ( .A(n8056), .B(n8057), .Z(n7022) );
  NANDN U7668 ( .A(n7015), .B(n7017), .Z(n8057) );
  NANDN U7669 ( .A(n7018), .B(n8058), .Z(n8056) );
  NANDN U7670 ( .A(n7017), .B(n7015), .Z(n8058) );
  XOR U7671 ( .A(n8048), .B(n8059), .Z(n7015) );
  XNOR U7672 ( .A(n8049), .B(n8050), .Z(n8059) );
  AND U7673 ( .A(n8060), .B(n8061), .Z(n8050) );
  NAND U7674 ( .A(n8062), .B(n8063), .Z(n8061) );
  NANDN U7675 ( .A(n8064), .B(n8065), .Z(n8060) );
  OR U7676 ( .A(n8062), .B(n8063), .Z(n8065) );
  ANDN U7677 ( .B(\stack[0][36] ), .A(n5219), .Z(n8049) );
  XOR U7678 ( .A(n8066), .B(n8067), .Z(n8048) );
  XNOR U7679 ( .A(n8068), .B(n8069), .Z(n8067) );
  ANDN U7680 ( .B(\stack[0][37] ), .A(n5195), .Z(n7017) );
  AND U7681 ( .A(n8070), .B(n8071), .Z(n7018) );
  NANDN U7682 ( .A(n7014), .B(n8072), .Z(n8070) );
  NANDN U7683 ( .A(n7013), .B(n7011), .Z(n8072) );
  XNOR U7684 ( .A(n8062), .B(n8073), .Z(n7011) );
  XNOR U7685 ( .A(n8063), .B(n8064), .Z(n8073) );
  AND U7686 ( .A(n8074), .B(n8075), .Z(n8064) );
  NANDN U7687 ( .A(n8076), .B(n8077), .Z(n8075) );
  NANDN U7688 ( .A(n8078), .B(n8079), .Z(n8074) );
  NANDN U7689 ( .A(n8077), .B(n8076), .Z(n8079) );
  ANDN U7690 ( .B(\stack[0][35] ), .A(n5219), .Z(n8063) );
  XNOR U7691 ( .A(n8080), .B(n8081), .Z(n8062) );
  XNOR U7692 ( .A(n8082), .B(n8083), .Z(n8081) );
  ANDN U7693 ( .B(\stack[1][1] ), .A(n6022), .Z(n7013) );
  AND U7694 ( .A(n8084), .B(n8085), .Z(n7014) );
  NANDN U7695 ( .A(n7007), .B(n7009), .Z(n8085) );
  NANDN U7696 ( .A(n7010), .B(n8086), .Z(n8084) );
  NANDN U7697 ( .A(n7009), .B(n7007), .Z(n8086) );
  XOR U7698 ( .A(n8076), .B(n8087), .Z(n7007) );
  XNOR U7699 ( .A(n8077), .B(n8078), .Z(n8087) );
  AND U7700 ( .A(n8088), .B(n8089), .Z(n8078) );
  NAND U7701 ( .A(n8090), .B(n8091), .Z(n8089) );
  NANDN U7702 ( .A(n8092), .B(n8093), .Z(n8088) );
  OR U7703 ( .A(n8090), .B(n8091), .Z(n8093) );
  ANDN U7704 ( .B(\stack[0][34] ), .A(n5219), .Z(n8077) );
  XOR U7705 ( .A(n8094), .B(n8095), .Z(n8076) );
  XNOR U7706 ( .A(n8096), .B(n8097), .Z(n8095) );
  ANDN U7707 ( .B(\stack[0][35] ), .A(n5195), .Z(n7009) );
  AND U7708 ( .A(n8098), .B(n8099), .Z(n7010) );
  NANDN U7709 ( .A(n7006), .B(n8100), .Z(n8098) );
  NANDN U7710 ( .A(n7005), .B(n7003), .Z(n8100) );
  XNOR U7711 ( .A(n8090), .B(n8101), .Z(n7003) );
  XNOR U7712 ( .A(n8091), .B(n8092), .Z(n8101) );
  AND U7713 ( .A(n8102), .B(n8103), .Z(n8092) );
  NANDN U7714 ( .A(n8104), .B(n8105), .Z(n8103) );
  NANDN U7715 ( .A(n8106), .B(n8107), .Z(n8102) );
  NANDN U7716 ( .A(n8105), .B(n8104), .Z(n8107) );
  ANDN U7717 ( .B(\stack[0][33] ), .A(n5219), .Z(n8091) );
  XNOR U7718 ( .A(n8108), .B(n8109), .Z(n8090) );
  XNOR U7719 ( .A(n8110), .B(n8111), .Z(n8109) );
  ANDN U7720 ( .B(\stack[1][1] ), .A(n5974), .Z(n7005) );
  AND U7721 ( .A(n8112), .B(n8113), .Z(n7006) );
  NANDN U7722 ( .A(n6999), .B(n7001), .Z(n8113) );
  NANDN U7723 ( .A(n7002), .B(n8114), .Z(n8112) );
  NANDN U7724 ( .A(n7001), .B(n6999), .Z(n8114) );
  XOR U7725 ( .A(n8104), .B(n8115), .Z(n6999) );
  XNOR U7726 ( .A(n8105), .B(n8106), .Z(n8115) );
  AND U7727 ( .A(n8116), .B(n8117), .Z(n8106) );
  NAND U7728 ( .A(n8118), .B(n8119), .Z(n8117) );
  NANDN U7729 ( .A(n8120), .B(n8121), .Z(n8116) );
  OR U7730 ( .A(n8118), .B(n8119), .Z(n8121) );
  ANDN U7731 ( .B(\stack[0][32] ), .A(n5219), .Z(n8105) );
  XOR U7732 ( .A(n8122), .B(n8123), .Z(n8104) );
  XNOR U7733 ( .A(n8124), .B(n8125), .Z(n8123) );
  ANDN U7734 ( .B(\stack[0][33] ), .A(n5195), .Z(n7001) );
  AND U7735 ( .A(n8126), .B(n8127), .Z(n7002) );
  NANDN U7736 ( .A(n6998), .B(n8128), .Z(n8126) );
  NANDN U7737 ( .A(n6997), .B(n6995), .Z(n8128) );
  XNOR U7738 ( .A(n8118), .B(n8129), .Z(n6995) );
  XNOR U7739 ( .A(n8119), .B(n8120), .Z(n8129) );
  AND U7740 ( .A(n8130), .B(n8131), .Z(n8120) );
  NANDN U7741 ( .A(n8132), .B(n8133), .Z(n8131) );
  NANDN U7742 ( .A(n8134), .B(n8135), .Z(n8130) );
  NANDN U7743 ( .A(n8133), .B(n8132), .Z(n8135) );
  ANDN U7744 ( .B(\stack[0][31] ), .A(n5219), .Z(n8119) );
  XNOR U7745 ( .A(n8136), .B(n8137), .Z(n8118) );
  XNOR U7746 ( .A(n8138), .B(n8139), .Z(n8137) );
  ANDN U7747 ( .B(\stack[1][1] ), .A(n5926), .Z(n6997) );
  AND U7748 ( .A(n8140), .B(n8141), .Z(n6998) );
  NANDN U7749 ( .A(n6991), .B(n6993), .Z(n8141) );
  NANDN U7750 ( .A(n6994), .B(n8142), .Z(n8140) );
  NANDN U7751 ( .A(n6993), .B(n6991), .Z(n8142) );
  XOR U7752 ( .A(n8132), .B(n8143), .Z(n6991) );
  XNOR U7753 ( .A(n8133), .B(n8134), .Z(n8143) );
  AND U7754 ( .A(n8144), .B(n8145), .Z(n8134) );
  NAND U7755 ( .A(n8146), .B(n8147), .Z(n8145) );
  NANDN U7756 ( .A(n8148), .B(n8149), .Z(n8144) );
  OR U7757 ( .A(n8146), .B(n8147), .Z(n8149) );
  ANDN U7758 ( .B(\stack[0][30] ), .A(n5219), .Z(n8133) );
  XOR U7759 ( .A(n8150), .B(n8151), .Z(n8132) );
  XNOR U7760 ( .A(n8152), .B(n8153), .Z(n8151) );
  ANDN U7761 ( .B(\stack[0][31] ), .A(n5195), .Z(n6993) );
  AND U7762 ( .A(n8154), .B(n8155), .Z(n6994) );
  NANDN U7763 ( .A(n6990), .B(n8156), .Z(n8154) );
  NANDN U7764 ( .A(n6989), .B(n6987), .Z(n8156) );
  XNOR U7765 ( .A(n8146), .B(n8157), .Z(n6987) );
  XNOR U7766 ( .A(n8147), .B(n8148), .Z(n8157) );
  AND U7767 ( .A(n8158), .B(n8159), .Z(n8148) );
  NANDN U7768 ( .A(n8160), .B(n8161), .Z(n8159) );
  NANDN U7769 ( .A(n8162), .B(n8163), .Z(n8158) );
  NANDN U7770 ( .A(n8161), .B(n8160), .Z(n8163) );
  ANDN U7771 ( .B(\stack[0][29] ), .A(n5219), .Z(n8147) );
  XNOR U7772 ( .A(n8164), .B(n8165), .Z(n8146) );
  XNOR U7773 ( .A(n8166), .B(n8167), .Z(n8165) );
  ANDN U7774 ( .B(\stack[1][1] ), .A(n5878), .Z(n6989) );
  AND U7775 ( .A(n8168), .B(n8169), .Z(n6990) );
  NANDN U7776 ( .A(n6983), .B(n6985), .Z(n8169) );
  NANDN U7777 ( .A(n6986), .B(n8170), .Z(n8168) );
  NANDN U7778 ( .A(n6985), .B(n6983), .Z(n8170) );
  XOR U7779 ( .A(n8160), .B(n8171), .Z(n6983) );
  XNOR U7780 ( .A(n8161), .B(n8162), .Z(n8171) );
  AND U7781 ( .A(n8172), .B(n8173), .Z(n8162) );
  NAND U7782 ( .A(n8174), .B(n8175), .Z(n8173) );
  NANDN U7783 ( .A(n8176), .B(n8177), .Z(n8172) );
  OR U7784 ( .A(n8174), .B(n8175), .Z(n8177) );
  ANDN U7785 ( .B(\stack[0][28] ), .A(n5219), .Z(n8161) );
  XOR U7786 ( .A(n8178), .B(n8179), .Z(n8160) );
  XNOR U7787 ( .A(n8180), .B(n8181), .Z(n8179) );
  ANDN U7788 ( .B(\stack[0][29] ), .A(n5195), .Z(n6985) );
  AND U7789 ( .A(n8182), .B(n8183), .Z(n6986) );
  NANDN U7790 ( .A(n6982), .B(n8184), .Z(n8182) );
  NANDN U7791 ( .A(n6981), .B(n6979), .Z(n8184) );
  XNOR U7792 ( .A(n8174), .B(n8185), .Z(n6979) );
  XNOR U7793 ( .A(n8175), .B(n8176), .Z(n8185) );
  AND U7794 ( .A(n8186), .B(n8187), .Z(n8176) );
  NANDN U7795 ( .A(n8188), .B(n8189), .Z(n8187) );
  NANDN U7796 ( .A(n8190), .B(n8191), .Z(n8186) );
  NANDN U7797 ( .A(n8189), .B(n8188), .Z(n8191) );
  ANDN U7798 ( .B(\stack[0][27] ), .A(n5219), .Z(n8175) );
  XNOR U7799 ( .A(n8192), .B(n8193), .Z(n8174) );
  XNOR U7800 ( .A(n8194), .B(n8195), .Z(n8193) );
  ANDN U7801 ( .B(\stack[1][1] ), .A(n5830), .Z(n6981) );
  AND U7802 ( .A(n8196), .B(n8197), .Z(n6982) );
  NANDN U7803 ( .A(n6975), .B(n6977), .Z(n8197) );
  NANDN U7804 ( .A(n6978), .B(n8198), .Z(n8196) );
  NANDN U7805 ( .A(n6977), .B(n6975), .Z(n8198) );
  XOR U7806 ( .A(n8188), .B(n8199), .Z(n6975) );
  XNOR U7807 ( .A(n8189), .B(n8190), .Z(n8199) );
  AND U7808 ( .A(n8200), .B(n8201), .Z(n8190) );
  NAND U7809 ( .A(n8202), .B(n8203), .Z(n8201) );
  NANDN U7810 ( .A(n8204), .B(n8205), .Z(n8200) );
  OR U7811 ( .A(n8202), .B(n8203), .Z(n8205) );
  ANDN U7812 ( .B(\stack[0][26] ), .A(n5219), .Z(n8189) );
  XOR U7813 ( .A(n8206), .B(n8207), .Z(n8188) );
  XNOR U7814 ( .A(n8208), .B(n8209), .Z(n8207) );
  ANDN U7815 ( .B(\stack[0][27] ), .A(n5195), .Z(n6977) );
  AND U7816 ( .A(n8210), .B(n8211), .Z(n6978) );
  NANDN U7817 ( .A(n6974), .B(n8212), .Z(n8210) );
  NANDN U7818 ( .A(n6973), .B(n6971), .Z(n8212) );
  XNOR U7819 ( .A(n8202), .B(n8213), .Z(n6971) );
  XNOR U7820 ( .A(n8203), .B(n8204), .Z(n8213) );
  AND U7821 ( .A(n8214), .B(n8215), .Z(n8204) );
  NANDN U7822 ( .A(n8216), .B(n8217), .Z(n8215) );
  NANDN U7823 ( .A(n8218), .B(n8219), .Z(n8214) );
  NANDN U7824 ( .A(n8217), .B(n8216), .Z(n8219) );
  ANDN U7825 ( .B(\stack[0][25] ), .A(n5219), .Z(n8203) );
  XNOR U7826 ( .A(n8220), .B(n8221), .Z(n8202) );
  XNOR U7827 ( .A(n8222), .B(n8223), .Z(n8221) );
  ANDN U7828 ( .B(\stack[1][1] ), .A(n5782), .Z(n6973) );
  AND U7829 ( .A(n8224), .B(n8225), .Z(n6974) );
  NANDN U7830 ( .A(n6967), .B(n6969), .Z(n8225) );
  NANDN U7831 ( .A(n6970), .B(n8226), .Z(n8224) );
  NANDN U7832 ( .A(n6969), .B(n6967), .Z(n8226) );
  XOR U7833 ( .A(n8216), .B(n8227), .Z(n6967) );
  XNOR U7834 ( .A(n8217), .B(n8218), .Z(n8227) );
  AND U7835 ( .A(n8228), .B(n8229), .Z(n8218) );
  NAND U7836 ( .A(n8230), .B(n8231), .Z(n8229) );
  NANDN U7837 ( .A(n8232), .B(n8233), .Z(n8228) );
  OR U7838 ( .A(n8230), .B(n8231), .Z(n8233) );
  ANDN U7839 ( .B(\stack[0][24] ), .A(n5219), .Z(n8217) );
  XOR U7840 ( .A(n8234), .B(n8235), .Z(n8216) );
  XNOR U7841 ( .A(n8236), .B(n8237), .Z(n8235) );
  ANDN U7842 ( .B(\stack[0][25] ), .A(n5195), .Z(n6969) );
  AND U7843 ( .A(n8238), .B(n8239), .Z(n6970) );
  NANDN U7844 ( .A(n6966), .B(n8240), .Z(n8238) );
  NANDN U7845 ( .A(n6965), .B(n6963), .Z(n8240) );
  XNOR U7846 ( .A(n8230), .B(n8241), .Z(n6963) );
  XNOR U7847 ( .A(n8231), .B(n8232), .Z(n8241) );
  AND U7848 ( .A(n8242), .B(n8243), .Z(n8232) );
  NANDN U7849 ( .A(n8244), .B(n8245), .Z(n8243) );
  NANDN U7850 ( .A(n8246), .B(n8247), .Z(n8242) );
  NANDN U7851 ( .A(n8245), .B(n8244), .Z(n8247) );
  ANDN U7852 ( .B(\stack[0][23] ), .A(n5219), .Z(n8231) );
  XNOR U7853 ( .A(n8248), .B(n8249), .Z(n8230) );
  XNOR U7854 ( .A(n8250), .B(n8251), .Z(n8249) );
  ANDN U7855 ( .B(\stack[1][1] ), .A(n5734), .Z(n6965) );
  AND U7856 ( .A(n8252), .B(n8253), .Z(n6966) );
  NANDN U7857 ( .A(n6959), .B(n6961), .Z(n8253) );
  NANDN U7858 ( .A(n6962), .B(n8254), .Z(n8252) );
  NANDN U7859 ( .A(n6961), .B(n6959), .Z(n8254) );
  XOR U7860 ( .A(n8244), .B(n8255), .Z(n6959) );
  XNOR U7861 ( .A(n8245), .B(n8246), .Z(n8255) );
  AND U7862 ( .A(n8256), .B(n8257), .Z(n8246) );
  NAND U7863 ( .A(n8258), .B(n8259), .Z(n8257) );
  NANDN U7864 ( .A(n8260), .B(n8261), .Z(n8256) );
  OR U7865 ( .A(n8258), .B(n8259), .Z(n8261) );
  ANDN U7866 ( .B(\stack[0][22] ), .A(n5219), .Z(n8245) );
  XOR U7867 ( .A(n8262), .B(n8263), .Z(n8244) );
  XNOR U7868 ( .A(n8264), .B(n8265), .Z(n8263) );
  ANDN U7869 ( .B(\stack[0][23] ), .A(n5195), .Z(n6961) );
  AND U7870 ( .A(n8266), .B(n8267), .Z(n6962) );
  NANDN U7871 ( .A(n6958), .B(n8268), .Z(n8266) );
  NANDN U7872 ( .A(n6957), .B(n6955), .Z(n8268) );
  XNOR U7873 ( .A(n8258), .B(n8269), .Z(n6955) );
  XNOR U7874 ( .A(n8259), .B(n8260), .Z(n8269) );
  AND U7875 ( .A(n8270), .B(n8271), .Z(n8260) );
  NANDN U7876 ( .A(n8272), .B(n8273), .Z(n8271) );
  NANDN U7877 ( .A(n8274), .B(n8275), .Z(n8270) );
  NANDN U7878 ( .A(n8273), .B(n8272), .Z(n8275) );
  ANDN U7879 ( .B(\stack[0][21] ), .A(n5219), .Z(n8259) );
  XNOR U7880 ( .A(n8276), .B(n8277), .Z(n8258) );
  XNOR U7881 ( .A(n8278), .B(n8279), .Z(n8277) );
  ANDN U7882 ( .B(\stack[1][1] ), .A(n5686), .Z(n6957) );
  AND U7883 ( .A(n8280), .B(n8281), .Z(n6958) );
  NANDN U7884 ( .A(n6951), .B(n6953), .Z(n8281) );
  NANDN U7885 ( .A(n6954), .B(n8282), .Z(n8280) );
  NANDN U7886 ( .A(n6953), .B(n6951), .Z(n8282) );
  XOR U7887 ( .A(n8272), .B(n8283), .Z(n6951) );
  XNOR U7888 ( .A(n8273), .B(n8274), .Z(n8283) );
  AND U7889 ( .A(n8284), .B(n8285), .Z(n8274) );
  NAND U7890 ( .A(n8286), .B(n8287), .Z(n8285) );
  NANDN U7891 ( .A(n8288), .B(n8289), .Z(n8284) );
  OR U7892 ( .A(n8286), .B(n8287), .Z(n8289) );
  ANDN U7893 ( .B(\stack[0][20] ), .A(n5219), .Z(n8273) );
  XOR U7894 ( .A(n8290), .B(n8291), .Z(n8272) );
  XNOR U7895 ( .A(n8292), .B(n8293), .Z(n8291) );
  ANDN U7896 ( .B(\stack[0][21] ), .A(n5195), .Z(n6953) );
  AND U7897 ( .A(n8294), .B(n8295), .Z(n6954) );
  NANDN U7898 ( .A(n6950), .B(n8296), .Z(n8294) );
  NANDN U7899 ( .A(n6949), .B(n6947), .Z(n8296) );
  XNOR U7900 ( .A(n8286), .B(n8297), .Z(n6947) );
  XNOR U7901 ( .A(n8287), .B(n8288), .Z(n8297) );
  AND U7902 ( .A(n8298), .B(n8299), .Z(n8288) );
  NANDN U7903 ( .A(n8300), .B(n8301), .Z(n8299) );
  NANDN U7904 ( .A(n8302), .B(n8303), .Z(n8298) );
  NANDN U7905 ( .A(n8301), .B(n8300), .Z(n8303) );
  ANDN U7906 ( .B(\stack[0][19] ), .A(n5219), .Z(n8287) );
  XNOR U7907 ( .A(n8304), .B(n8305), .Z(n8286) );
  XNOR U7908 ( .A(n8306), .B(n8307), .Z(n8305) );
  ANDN U7909 ( .B(\stack[1][1] ), .A(n5638), .Z(n6949) );
  AND U7910 ( .A(n8308), .B(n8309), .Z(n6950) );
  NANDN U7911 ( .A(n6943), .B(n6945), .Z(n8309) );
  NANDN U7912 ( .A(n6946), .B(n8310), .Z(n8308) );
  NANDN U7913 ( .A(n6945), .B(n6943), .Z(n8310) );
  XOR U7914 ( .A(n8300), .B(n8311), .Z(n6943) );
  XNOR U7915 ( .A(n8301), .B(n8302), .Z(n8311) );
  AND U7916 ( .A(n8312), .B(n8313), .Z(n8302) );
  NAND U7917 ( .A(n8314), .B(n8315), .Z(n8313) );
  NANDN U7918 ( .A(n8316), .B(n8317), .Z(n8312) );
  OR U7919 ( .A(n8314), .B(n8315), .Z(n8317) );
  ANDN U7920 ( .B(\stack[0][18] ), .A(n5219), .Z(n8301) );
  XOR U7921 ( .A(n8318), .B(n8319), .Z(n8300) );
  XNOR U7922 ( .A(n8320), .B(n8321), .Z(n8319) );
  ANDN U7923 ( .B(\stack[0][19] ), .A(n5195), .Z(n6945) );
  AND U7924 ( .A(n8322), .B(n8323), .Z(n6946) );
  NANDN U7925 ( .A(n6942), .B(n8324), .Z(n8322) );
  NANDN U7926 ( .A(n6941), .B(n6939), .Z(n8324) );
  XNOR U7927 ( .A(n8314), .B(n8325), .Z(n6939) );
  XNOR U7928 ( .A(n8315), .B(n8316), .Z(n8325) );
  AND U7929 ( .A(n8326), .B(n8327), .Z(n8316) );
  NANDN U7930 ( .A(n8328), .B(n8329), .Z(n8327) );
  NANDN U7931 ( .A(n8330), .B(n8331), .Z(n8326) );
  NANDN U7932 ( .A(n8329), .B(n8328), .Z(n8331) );
  ANDN U7933 ( .B(\stack[0][17] ), .A(n5219), .Z(n8315) );
  XNOR U7934 ( .A(n8332), .B(n8333), .Z(n8314) );
  XNOR U7935 ( .A(n8334), .B(n8335), .Z(n8333) );
  ANDN U7936 ( .B(\stack[1][1] ), .A(n5590), .Z(n6941) );
  AND U7937 ( .A(n8336), .B(n8337), .Z(n6942) );
  NANDN U7938 ( .A(n6935), .B(n6937), .Z(n8337) );
  NANDN U7939 ( .A(n6938), .B(n8338), .Z(n8336) );
  NANDN U7940 ( .A(n6937), .B(n6935), .Z(n8338) );
  XOR U7941 ( .A(n8328), .B(n8339), .Z(n6935) );
  XNOR U7942 ( .A(n8329), .B(n8330), .Z(n8339) );
  AND U7943 ( .A(n8340), .B(n8341), .Z(n8330) );
  NAND U7944 ( .A(n8342), .B(n8343), .Z(n8341) );
  NANDN U7945 ( .A(n8344), .B(n8345), .Z(n8340) );
  OR U7946 ( .A(n8342), .B(n8343), .Z(n8345) );
  ANDN U7947 ( .B(\stack[0][16] ), .A(n5219), .Z(n8329) );
  XOR U7948 ( .A(n8346), .B(n8347), .Z(n8328) );
  XNOR U7949 ( .A(n8348), .B(n8349), .Z(n8347) );
  ANDN U7950 ( .B(\stack[0][17] ), .A(n5195), .Z(n6937) );
  AND U7951 ( .A(n8350), .B(n8351), .Z(n6938) );
  NANDN U7952 ( .A(n6934), .B(n8352), .Z(n8350) );
  NANDN U7953 ( .A(n6933), .B(n6931), .Z(n8352) );
  XNOR U7954 ( .A(n8342), .B(n8353), .Z(n6931) );
  XNOR U7955 ( .A(n8343), .B(n8344), .Z(n8353) );
  AND U7956 ( .A(n8354), .B(n8355), .Z(n8344) );
  NANDN U7957 ( .A(n8356), .B(n8357), .Z(n8355) );
  NANDN U7958 ( .A(n8358), .B(n8359), .Z(n8354) );
  NANDN U7959 ( .A(n8357), .B(n8356), .Z(n8359) );
  ANDN U7960 ( .B(\stack[0][15] ), .A(n5219), .Z(n8343) );
  XNOR U7961 ( .A(n8360), .B(n8361), .Z(n8342) );
  XNOR U7962 ( .A(n8362), .B(n8363), .Z(n8361) );
  ANDN U7963 ( .B(\stack[1][1] ), .A(n5542), .Z(n6933) );
  AND U7964 ( .A(n8364), .B(n8365), .Z(n6934) );
  NANDN U7965 ( .A(n6927), .B(n6929), .Z(n8365) );
  NANDN U7966 ( .A(n6930), .B(n8366), .Z(n8364) );
  NANDN U7967 ( .A(n6929), .B(n6927), .Z(n8366) );
  XOR U7968 ( .A(n8356), .B(n8367), .Z(n6927) );
  XNOR U7969 ( .A(n8357), .B(n8358), .Z(n8367) );
  AND U7970 ( .A(n8368), .B(n8369), .Z(n8358) );
  NAND U7971 ( .A(n8370), .B(n8371), .Z(n8369) );
  NANDN U7972 ( .A(n8372), .B(n8373), .Z(n8368) );
  OR U7973 ( .A(n8370), .B(n8371), .Z(n8373) );
  ANDN U7974 ( .B(\stack[0][14] ), .A(n5219), .Z(n8357) );
  XOR U7975 ( .A(n8374), .B(n8375), .Z(n8356) );
  XNOR U7976 ( .A(n8376), .B(n8377), .Z(n8375) );
  ANDN U7977 ( .B(\stack[0][15] ), .A(n5195), .Z(n6929) );
  AND U7978 ( .A(n8378), .B(n8379), .Z(n6930) );
  NANDN U7979 ( .A(n6926), .B(n8380), .Z(n8378) );
  NANDN U7980 ( .A(n6925), .B(n6923), .Z(n8380) );
  XNOR U7981 ( .A(n8370), .B(n8381), .Z(n6923) );
  XNOR U7982 ( .A(n8371), .B(n8372), .Z(n8381) );
  AND U7983 ( .A(n8382), .B(n8383), .Z(n8372) );
  NANDN U7984 ( .A(n8384), .B(n8385), .Z(n8383) );
  NANDN U7985 ( .A(n8386), .B(n8387), .Z(n8382) );
  NANDN U7986 ( .A(n8385), .B(n8384), .Z(n8387) );
  ANDN U7987 ( .B(\stack[0][13] ), .A(n5219), .Z(n8371) );
  XNOR U7988 ( .A(n8388), .B(n8389), .Z(n8370) );
  XNOR U7989 ( .A(n8390), .B(n8391), .Z(n8389) );
  ANDN U7990 ( .B(\stack[1][1] ), .A(n5494), .Z(n6925) );
  AND U7991 ( .A(n8392), .B(n8393), .Z(n6926) );
  NANDN U7992 ( .A(n6919), .B(n6921), .Z(n8393) );
  NANDN U7993 ( .A(n6922), .B(n8394), .Z(n8392) );
  NANDN U7994 ( .A(n6921), .B(n6919), .Z(n8394) );
  XOR U7995 ( .A(n8384), .B(n8395), .Z(n6919) );
  XNOR U7996 ( .A(n8385), .B(n8386), .Z(n8395) );
  AND U7997 ( .A(n8396), .B(n8397), .Z(n8386) );
  NAND U7998 ( .A(n8398), .B(n8399), .Z(n8397) );
  NANDN U7999 ( .A(n8400), .B(n8401), .Z(n8396) );
  OR U8000 ( .A(n8398), .B(n8399), .Z(n8401) );
  ANDN U8001 ( .B(\stack[0][12] ), .A(n5219), .Z(n8385) );
  XOR U8002 ( .A(n8402), .B(n8403), .Z(n8384) );
  XNOR U8003 ( .A(n8404), .B(n8405), .Z(n8403) );
  ANDN U8004 ( .B(\stack[0][13] ), .A(n5195), .Z(n6921) );
  AND U8005 ( .A(n8406), .B(n8407), .Z(n6922) );
  NANDN U8006 ( .A(n6918), .B(n8408), .Z(n8406) );
  NANDN U8007 ( .A(n6917), .B(n6915), .Z(n8408) );
  XNOR U8008 ( .A(n8398), .B(n8409), .Z(n6915) );
  XNOR U8009 ( .A(n8399), .B(n8400), .Z(n8409) );
  AND U8010 ( .A(n8410), .B(n8411), .Z(n8400) );
  NANDN U8011 ( .A(n8412), .B(n8413), .Z(n8411) );
  NANDN U8012 ( .A(n8414), .B(n8415), .Z(n8410) );
  NANDN U8013 ( .A(n8413), .B(n8412), .Z(n8415) );
  ANDN U8014 ( .B(\stack[0][11] ), .A(n5219), .Z(n8399) );
  XNOR U8015 ( .A(n8416), .B(n8417), .Z(n8398) );
  XNOR U8016 ( .A(n8418), .B(n8419), .Z(n8417) );
  ANDN U8017 ( .B(\stack[1][1] ), .A(n5446), .Z(n6917) );
  AND U8018 ( .A(n8420), .B(n8421), .Z(n6918) );
  NANDN U8019 ( .A(n6911), .B(n6913), .Z(n8421) );
  NANDN U8020 ( .A(n6914), .B(n8422), .Z(n8420) );
  NANDN U8021 ( .A(n6913), .B(n6911), .Z(n8422) );
  XOR U8022 ( .A(n8412), .B(n8423), .Z(n6911) );
  XNOR U8023 ( .A(n8413), .B(n8414), .Z(n8423) );
  AND U8024 ( .A(n8424), .B(n8425), .Z(n8414) );
  NAND U8025 ( .A(n8426), .B(n8427), .Z(n8425) );
  NANDN U8026 ( .A(n8428), .B(n8429), .Z(n8424) );
  OR U8027 ( .A(n8426), .B(n8427), .Z(n8429) );
  ANDN U8028 ( .B(\stack[0][10] ), .A(n5219), .Z(n8413) );
  XOR U8029 ( .A(n8430), .B(n8431), .Z(n8412) );
  XNOR U8030 ( .A(n8432), .B(n8433), .Z(n8431) );
  ANDN U8031 ( .B(\stack[0][11] ), .A(n5195), .Z(n6913) );
  AND U8032 ( .A(n8434), .B(n8435), .Z(n6914) );
  NANDN U8033 ( .A(n6910), .B(n8436), .Z(n8434) );
  NANDN U8034 ( .A(n6909), .B(n6907), .Z(n8436) );
  XNOR U8035 ( .A(n8426), .B(n8437), .Z(n6907) );
  XNOR U8036 ( .A(n8427), .B(n8428), .Z(n8437) );
  AND U8037 ( .A(n8438), .B(n8439), .Z(n8428) );
  NANDN U8038 ( .A(n8440), .B(n8441), .Z(n8439) );
  NANDN U8039 ( .A(n8442), .B(n8443), .Z(n8438) );
  NANDN U8040 ( .A(n8441), .B(n8440), .Z(n8443) );
  ANDN U8041 ( .B(\stack[1][2] ), .A(n5374), .Z(n8427) );
  XNOR U8042 ( .A(n8444), .B(n8445), .Z(n8426) );
  XNOR U8043 ( .A(n8446), .B(n8447), .Z(n8445) );
  ANDN U8044 ( .B(\stack[1][1] ), .A(n5398), .Z(n6909) );
  AND U8045 ( .A(n8448), .B(n8449), .Z(n6910) );
  NANDN U8046 ( .A(n6849), .B(n6851), .Z(n8449) );
  NANDN U8047 ( .A(n6852), .B(n8450), .Z(n8448) );
  NANDN U8048 ( .A(n6851), .B(n6849), .Z(n8450) );
  XOR U8049 ( .A(n8440), .B(n8451), .Z(n6849) );
  XNOR U8050 ( .A(n8441), .B(n8442), .Z(n8451) );
  AND U8051 ( .A(n8452), .B(n8453), .Z(n8442) );
  NANDN U8052 ( .A(n8454), .B(n8455), .Z(n8453) );
  NANDN U8053 ( .A(n8456), .B(n8457), .Z(n8452) );
  OR U8054 ( .A(n8455), .B(n8458), .Z(n8457) );
  ANDN U8055 ( .B(\stack[0][8] ), .A(n5219), .Z(n8441) );
  XOR U8056 ( .A(n8459), .B(n8460), .Z(n8440) );
  XNOR U8057 ( .A(n8461), .B(n8462), .Z(n8460) );
  ANDN U8058 ( .B(\stack[1][1] ), .A(n5374), .Z(n6851) );
  AND U8059 ( .A(n8463), .B(n8464), .Z(n6852) );
  NANDN U8060 ( .A(n6856), .B(n6858), .Z(n8464) );
  IV U8061 ( .A(n8465), .Z(n6856) );
  NANDN U8062 ( .A(n6859), .B(n8466), .Z(n8463) );
  OR U8063 ( .A(n6858), .B(n8465), .Z(n8466) );
  XOR U8064 ( .A(n8455), .B(n8467), .Z(n8465) );
  XOR U8065 ( .A(n8454), .B(n8456), .Z(n8467) );
  AND U8066 ( .A(n8468), .B(n8469), .Z(n8456) );
  NANDN U8067 ( .A(n8472), .B(n8473), .Z(n8468) );
  NANDN U8068 ( .A(n8471), .B(n8470), .Z(n8473) );
  IV U8069 ( .A(n8458), .Z(n8454) );
  ANDN U8070 ( .B(\stack[0][7] ), .A(n5219), .Z(n8458) );
  XNOR U8071 ( .A(n8474), .B(n8475), .Z(n8455) );
  XNOR U8072 ( .A(n8476), .B(n8477), .Z(n8475) );
  AND U8073 ( .A(\stack[0][8] ), .B(\stack[1][1] ), .Z(n6858) );
  AND U8074 ( .A(n8478), .B(n8479), .Z(n6859) );
  NANDN U8075 ( .A(n6863), .B(n6865), .Z(n8479) );
  NANDN U8076 ( .A(n6866), .B(n8480), .Z(n8478) );
  NANDN U8077 ( .A(n6865), .B(n6863), .Z(n8480) );
  XOR U8078 ( .A(n8470), .B(n8481), .Z(n6863) );
  XNOR U8079 ( .A(n8471), .B(n8472), .Z(n8481) );
  AND U8080 ( .A(n8482), .B(n8483), .Z(n8472) );
  NANDN U8081 ( .A(n8484), .B(n8485), .Z(n8483) );
  NANDN U8082 ( .A(n8486), .B(n8487), .Z(n8482) );
  NANDN U8083 ( .A(n8485), .B(n8484), .Z(n8487) );
  ANDN U8084 ( .B(\stack[0][6] ), .A(n5219), .Z(n8471) );
  XOR U8085 ( .A(n8488), .B(n8489), .Z(n8470) );
  XNOR U8086 ( .A(n8490), .B(n8491), .Z(n8489) );
  ANDN U8087 ( .B(\stack[1][1] ), .A(n5326), .Z(n6865) );
  AND U8088 ( .A(n8492), .B(n8493), .Z(n6866) );
  NANDN U8089 ( .A(n6906), .B(n8494), .Z(n8492) );
  NANDN U8090 ( .A(n6905), .B(n6903), .Z(n8494) );
  XOR U8091 ( .A(n8484), .B(n8495), .Z(n6903) );
  XNOR U8092 ( .A(n8485), .B(n8486), .Z(n8495) );
  AND U8093 ( .A(n8496), .B(n8497), .Z(n8486) );
  NANDN U8094 ( .A(n8500), .B(n8501), .Z(n8496) );
  NANDN U8095 ( .A(n8499), .B(n8498), .Z(n8501) );
  ANDN U8096 ( .B(\stack[1][2] ), .A(n5278), .Z(n8485) );
  XOR U8097 ( .A(n8502), .B(n8503), .Z(n8484) );
  XNOR U8098 ( .A(n8504), .B(n8505), .Z(n8503) );
  ANDN U8099 ( .B(\stack[0][6] ), .A(n5195), .Z(n6905) );
  AND U8100 ( .A(n8506), .B(n8507), .Z(n6906) );
  NANDN U8101 ( .A(n6873), .B(n6875), .Z(n8507) );
  NANDN U8102 ( .A(n6876), .B(n8508), .Z(n8506) );
  NANDN U8103 ( .A(n6875), .B(n6873), .Z(n8508) );
  XOR U8104 ( .A(n8498), .B(n8509), .Z(n6873) );
  XNOR U8105 ( .A(n8499), .B(n8500), .Z(n8509) );
  AND U8106 ( .A(n8510), .B(n8511), .Z(n8500) );
  NANDN U8107 ( .A(n8512), .B(n8513), .Z(n8511) );
  NANDN U8108 ( .A(n8514), .B(n8515), .Z(n8510) );
  NANDN U8109 ( .A(n8513), .B(n8512), .Z(n8515) );
  ANDN U8110 ( .B(\stack[0][4] ), .A(n5219), .Z(n8499) );
  XOR U8111 ( .A(n8516), .B(n8517), .Z(n8498) );
  XNOR U8112 ( .A(n8518), .B(n8519), .Z(n8517) );
  ANDN U8113 ( .B(\stack[1][1] ), .A(n5278), .Z(n6875) );
  AND U8114 ( .A(n8520), .B(n8521), .Z(n6876) );
  NANDN U8115 ( .A(n6902), .B(n8522), .Z(n8520) );
  NANDN U8116 ( .A(n6901), .B(n6899), .Z(n8522) );
  XOR U8117 ( .A(n8512), .B(n8523), .Z(n6899) );
  XNOR U8118 ( .A(n8513), .B(n8514), .Z(n8523) );
  AND U8119 ( .A(n8524), .B(n8525), .Z(n8514) );
  NANDN U8120 ( .A(n8526), .B(n8527), .Z(n8525) );
  NAND U8121 ( .A(n8528), .B(n8529), .Z(n8524) );
  NANDN U8122 ( .A(n8527), .B(n8526), .Z(n8528) );
  ANDN U8123 ( .B(\stack[1][2] ), .A(n5230), .Z(n8513) );
  XNOR U8124 ( .A(n8530), .B(n8531), .Z(n8512) );
  XNOR U8125 ( .A(n8532), .B(n8533), .Z(n8531) );
  ANDN U8126 ( .B(\stack[0][4] ), .A(n5195), .Z(n6901) );
  AND U8127 ( .A(n8534), .B(n8535), .Z(n6902) );
  NANDN U8128 ( .A(n6883), .B(n6885), .Z(n8535) );
  NANDN U8129 ( .A(n6886), .B(n8536), .Z(n8534) );
  NANDN U8130 ( .A(n6885), .B(n6883), .Z(n8536) );
  XNOR U8131 ( .A(n8526), .B(n8537), .Z(n6883) );
  XNOR U8132 ( .A(n8527), .B(n8529), .Z(n8537) );
  ANDN U8133 ( .B(n8538), .A(n8539), .Z(n8529) );
  ANDN U8134 ( .B(\stack[0][0] ), .A(n5243), .Z(n8538) );
  ANDN U8135 ( .B(\stack[1][2] ), .A(n5206), .Z(n8527) );
  XNOR U8136 ( .A(n8540), .B(n8541), .Z(n8526) );
  NANDN U8137 ( .A(n5160), .B(\stack[1][4] ), .Z(n8541) );
  ANDN U8138 ( .B(\stack[1][1] ), .A(n5230), .Z(n6885) );
  AND U8139 ( .A(n8542), .B(n8543), .Z(n6886) );
  NANDN U8140 ( .A(n6890), .B(n6892), .Z(n8543) );
  NAND U8141 ( .A(n8544), .B(n6893), .Z(n8542) );
  ANDN U8142 ( .B(n8545), .A(n6897), .Z(n6893) );
  NANDN U8143 ( .A(n5195), .B(\stack[0][1] ), .Z(n6897) );
  ANDN U8144 ( .B(\stack[0][0] ), .A(n5219), .Z(n8545) );
  NANDN U8145 ( .A(n6892), .B(n6890), .Z(n8544) );
  XNOR U8146 ( .A(n8539), .B(n8546), .Z(n6890) );
  NANDN U8147 ( .A(n5160), .B(\stack[1][3] ), .Z(n8546) );
  NANDN U8148 ( .A(n5219), .B(\stack[0][1] ), .Z(n8539) );
  ANDN U8149 ( .B(\stack[1][1] ), .A(n5206), .Z(n6892) );
  XOR U8150 ( .A(n8547), .B(n8548), .Z(n7119) );
  AND U8151 ( .A(n8549), .B(n8550), .Z(n8548) );
  NANDN U8152 ( .A(n7730), .B(n7732), .Z(n8550) );
  NANDN U8153 ( .A(n7733), .B(n8551), .Z(n8549) );
  NANDN U8154 ( .A(n7732), .B(n7730), .Z(n8551) );
  XOR U8155 ( .A(n8552), .B(n8553), .Z(n7730) );
  XNOR U8156 ( .A(n8554), .B(n8555), .Z(n8553) );
  ANDN U8157 ( .B(\stack[0][59] ), .A(n5243), .Z(n7732) );
  AND U8158 ( .A(n8556), .B(n8557), .Z(n7733) );
  NANDN U8159 ( .A(n7747), .B(n8558), .Z(n8556) );
  NANDN U8160 ( .A(n7746), .B(n7744), .Z(n8558) );
  XOR U8161 ( .A(n8559), .B(n8560), .Z(n7744) );
  XNOR U8162 ( .A(n8561), .B(n8562), .Z(n8560) );
  ANDN U8163 ( .B(\stack[1][3] ), .A(n6550), .Z(n7746) );
  AND U8164 ( .A(n8563), .B(n8564), .Z(n7747) );
  NANDN U8165 ( .A(n7758), .B(n7760), .Z(n8564) );
  NANDN U8166 ( .A(n7761), .B(n8565), .Z(n8563) );
  NANDN U8167 ( .A(n7760), .B(n7758), .Z(n8565) );
  XOR U8168 ( .A(n8566), .B(n8567), .Z(n7758) );
  XNOR U8169 ( .A(n8568), .B(n8569), .Z(n8567) );
  ANDN U8170 ( .B(\stack[0][57] ), .A(n5243), .Z(n7760) );
  AND U8171 ( .A(n8570), .B(n8571), .Z(n7761) );
  NANDN U8172 ( .A(n7775), .B(n8572), .Z(n8570) );
  NANDN U8173 ( .A(n7774), .B(n7772), .Z(n8572) );
  XOR U8174 ( .A(n8573), .B(n8574), .Z(n7772) );
  XNOR U8175 ( .A(n8575), .B(n8576), .Z(n8574) );
  ANDN U8176 ( .B(\stack[1][3] ), .A(n6502), .Z(n7774) );
  AND U8177 ( .A(n8577), .B(n8578), .Z(n7775) );
  NANDN U8178 ( .A(n7786), .B(n7788), .Z(n8578) );
  NANDN U8179 ( .A(n7789), .B(n8579), .Z(n8577) );
  NANDN U8180 ( .A(n7788), .B(n7786), .Z(n8579) );
  XOR U8181 ( .A(n8580), .B(n8581), .Z(n7786) );
  XNOR U8182 ( .A(n8582), .B(n8583), .Z(n8581) );
  ANDN U8183 ( .B(\stack[0][55] ), .A(n5243), .Z(n7788) );
  AND U8184 ( .A(n8584), .B(n8585), .Z(n7789) );
  NANDN U8185 ( .A(n7803), .B(n8586), .Z(n8584) );
  NANDN U8186 ( .A(n7802), .B(n7800), .Z(n8586) );
  XOR U8187 ( .A(n8587), .B(n8588), .Z(n7800) );
  XNOR U8188 ( .A(n8589), .B(n8590), .Z(n8588) );
  ANDN U8189 ( .B(\stack[1][3] ), .A(n6454), .Z(n7802) );
  AND U8190 ( .A(n8591), .B(n8592), .Z(n7803) );
  NANDN U8191 ( .A(n7814), .B(n7816), .Z(n8592) );
  NANDN U8192 ( .A(n7817), .B(n8593), .Z(n8591) );
  NANDN U8193 ( .A(n7816), .B(n7814), .Z(n8593) );
  XOR U8194 ( .A(n8594), .B(n8595), .Z(n7814) );
  XNOR U8195 ( .A(n8596), .B(n8597), .Z(n8595) );
  ANDN U8196 ( .B(\stack[0][53] ), .A(n5243), .Z(n7816) );
  AND U8197 ( .A(n8598), .B(n8599), .Z(n7817) );
  NANDN U8198 ( .A(n7831), .B(n8600), .Z(n8598) );
  NANDN U8199 ( .A(n7830), .B(n7828), .Z(n8600) );
  XOR U8200 ( .A(n8601), .B(n8602), .Z(n7828) );
  XNOR U8201 ( .A(n8603), .B(n8604), .Z(n8602) );
  ANDN U8202 ( .B(\stack[1][3] ), .A(n6406), .Z(n7830) );
  AND U8203 ( .A(n8605), .B(n8606), .Z(n7831) );
  NANDN U8204 ( .A(n7842), .B(n7844), .Z(n8606) );
  NANDN U8205 ( .A(n7845), .B(n8607), .Z(n8605) );
  NANDN U8206 ( .A(n7844), .B(n7842), .Z(n8607) );
  XOR U8207 ( .A(n8608), .B(n8609), .Z(n7842) );
  XNOR U8208 ( .A(n8610), .B(n8611), .Z(n8609) );
  ANDN U8209 ( .B(\stack[0][51] ), .A(n5243), .Z(n7844) );
  AND U8210 ( .A(n8612), .B(n8613), .Z(n7845) );
  NANDN U8211 ( .A(n7859), .B(n8614), .Z(n8612) );
  NANDN U8212 ( .A(n7858), .B(n7856), .Z(n8614) );
  XOR U8213 ( .A(n8615), .B(n8616), .Z(n7856) );
  XNOR U8214 ( .A(n8617), .B(n8618), .Z(n8616) );
  ANDN U8215 ( .B(\stack[1][3] ), .A(n6358), .Z(n7858) );
  AND U8216 ( .A(n8619), .B(n8620), .Z(n7859) );
  NANDN U8217 ( .A(n7870), .B(n7872), .Z(n8620) );
  NANDN U8218 ( .A(n7873), .B(n8621), .Z(n8619) );
  NANDN U8219 ( .A(n7872), .B(n7870), .Z(n8621) );
  XOR U8220 ( .A(n8622), .B(n8623), .Z(n7870) );
  XNOR U8221 ( .A(n8624), .B(n8625), .Z(n8623) );
  ANDN U8222 ( .B(\stack[0][49] ), .A(n5243), .Z(n7872) );
  AND U8223 ( .A(n8626), .B(n8627), .Z(n7873) );
  NANDN U8224 ( .A(n7887), .B(n8628), .Z(n8626) );
  NANDN U8225 ( .A(n7886), .B(n7884), .Z(n8628) );
  XOR U8226 ( .A(n8629), .B(n8630), .Z(n7884) );
  XNOR U8227 ( .A(n8631), .B(n8632), .Z(n8630) );
  ANDN U8228 ( .B(\stack[1][3] ), .A(n6310), .Z(n7886) );
  AND U8229 ( .A(n8633), .B(n8634), .Z(n7887) );
  NANDN U8230 ( .A(n7898), .B(n7900), .Z(n8634) );
  NANDN U8231 ( .A(n7901), .B(n8635), .Z(n8633) );
  NANDN U8232 ( .A(n7900), .B(n7898), .Z(n8635) );
  XOR U8233 ( .A(n8636), .B(n8637), .Z(n7898) );
  XNOR U8234 ( .A(n8638), .B(n8639), .Z(n8637) );
  ANDN U8235 ( .B(\stack[0][47] ), .A(n5243), .Z(n7900) );
  AND U8236 ( .A(n8640), .B(n8641), .Z(n7901) );
  NANDN U8237 ( .A(n7915), .B(n8642), .Z(n8640) );
  NANDN U8238 ( .A(n7914), .B(n7912), .Z(n8642) );
  XOR U8239 ( .A(n8643), .B(n8644), .Z(n7912) );
  XNOR U8240 ( .A(n8645), .B(n8646), .Z(n8644) );
  ANDN U8241 ( .B(\stack[1][3] ), .A(n6262), .Z(n7914) );
  AND U8242 ( .A(n8647), .B(n8648), .Z(n7915) );
  NANDN U8243 ( .A(n7926), .B(n7928), .Z(n8648) );
  NANDN U8244 ( .A(n7929), .B(n8649), .Z(n8647) );
  NANDN U8245 ( .A(n7928), .B(n7926), .Z(n8649) );
  XOR U8246 ( .A(n8650), .B(n8651), .Z(n7926) );
  XNOR U8247 ( .A(n8652), .B(n8653), .Z(n8651) );
  ANDN U8248 ( .B(\stack[0][45] ), .A(n5243), .Z(n7928) );
  AND U8249 ( .A(n8654), .B(n8655), .Z(n7929) );
  NANDN U8250 ( .A(n7943), .B(n8656), .Z(n8654) );
  NANDN U8251 ( .A(n7942), .B(n7940), .Z(n8656) );
  XOR U8252 ( .A(n8657), .B(n8658), .Z(n7940) );
  XNOR U8253 ( .A(n8659), .B(n8660), .Z(n8658) );
  ANDN U8254 ( .B(\stack[1][3] ), .A(n6214), .Z(n7942) );
  AND U8255 ( .A(n8661), .B(n8662), .Z(n7943) );
  NANDN U8256 ( .A(n7954), .B(n7956), .Z(n8662) );
  NANDN U8257 ( .A(n7957), .B(n8663), .Z(n8661) );
  NANDN U8258 ( .A(n7956), .B(n7954), .Z(n8663) );
  XOR U8259 ( .A(n8664), .B(n8665), .Z(n7954) );
  XNOR U8260 ( .A(n8666), .B(n8667), .Z(n8665) );
  ANDN U8261 ( .B(\stack[0][43] ), .A(n5243), .Z(n7956) );
  AND U8262 ( .A(n8668), .B(n8669), .Z(n7957) );
  NANDN U8263 ( .A(n7971), .B(n8670), .Z(n8668) );
  NANDN U8264 ( .A(n7970), .B(n7968), .Z(n8670) );
  XOR U8265 ( .A(n8671), .B(n8672), .Z(n7968) );
  XNOR U8266 ( .A(n8673), .B(n8674), .Z(n8672) );
  ANDN U8267 ( .B(\stack[1][3] ), .A(n6166), .Z(n7970) );
  AND U8268 ( .A(n8675), .B(n8676), .Z(n7971) );
  NANDN U8269 ( .A(n7982), .B(n7984), .Z(n8676) );
  NANDN U8270 ( .A(n7985), .B(n8677), .Z(n8675) );
  NANDN U8271 ( .A(n7984), .B(n7982), .Z(n8677) );
  XOR U8272 ( .A(n8678), .B(n8679), .Z(n7982) );
  XNOR U8273 ( .A(n8680), .B(n8681), .Z(n8679) );
  ANDN U8274 ( .B(\stack[0][41] ), .A(n5243), .Z(n7984) );
  AND U8275 ( .A(n8682), .B(n8683), .Z(n7985) );
  NANDN U8276 ( .A(n7999), .B(n8684), .Z(n8682) );
  NANDN U8277 ( .A(n7998), .B(n7996), .Z(n8684) );
  XOR U8278 ( .A(n8685), .B(n8686), .Z(n7996) );
  XNOR U8279 ( .A(n8687), .B(n8688), .Z(n8686) );
  ANDN U8280 ( .B(\stack[1][3] ), .A(n6118), .Z(n7998) );
  AND U8281 ( .A(n8689), .B(n8690), .Z(n7999) );
  NANDN U8282 ( .A(n8010), .B(n8012), .Z(n8690) );
  NANDN U8283 ( .A(n8013), .B(n8691), .Z(n8689) );
  NANDN U8284 ( .A(n8012), .B(n8010), .Z(n8691) );
  XOR U8285 ( .A(n8692), .B(n8693), .Z(n8010) );
  XNOR U8286 ( .A(n8694), .B(n8695), .Z(n8693) );
  ANDN U8287 ( .B(\stack[0][39] ), .A(n5243), .Z(n8012) );
  AND U8288 ( .A(n8696), .B(n8697), .Z(n8013) );
  NANDN U8289 ( .A(n8027), .B(n8698), .Z(n8696) );
  NANDN U8290 ( .A(n8026), .B(n8024), .Z(n8698) );
  XOR U8291 ( .A(n8699), .B(n8700), .Z(n8024) );
  XNOR U8292 ( .A(n8701), .B(n8702), .Z(n8700) );
  ANDN U8293 ( .B(\stack[1][3] ), .A(n6070), .Z(n8026) );
  AND U8294 ( .A(n8703), .B(n8704), .Z(n8027) );
  NANDN U8295 ( .A(n8038), .B(n8040), .Z(n8704) );
  NANDN U8296 ( .A(n8041), .B(n8705), .Z(n8703) );
  NANDN U8297 ( .A(n8040), .B(n8038), .Z(n8705) );
  XOR U8298 ( .A(n8706), .B(n8707), .Z(n8038) );
  XNOR U8299 ( .A(n8708), .B(n8709), .Z(n8707) );
  ANDN U8300 ( .B(\stack[0][37] ), .A(n5243), .Z(n8040) );
  AND U8301 ( .A(n8710), .B(n8711), .Z(n8041) );
  NANDN U8302 ( .A(n8055), .B(n8712), .Z(n8710) );
  NANDN U8303 ( .A(n8054), .B(n8052), .Z(n8712) );
  XOR U8304 ( .A(n8713), .B(n8714), .Z(n8052) );
  XNOR U8305 ( .A(n8715), .B(n8716), .Z(n8714) );
  ANDN U8306 ( .B(\stack[1][3] ), .A(n6022), .Z(n8054) );
  AND U8307 ( .A(n8717), .B(n8718), .Z(n8055) );
  NANDN U8308 ( .A(n8066), .B(n8068), .Z(n8718) );
  NANDN U8309 ( .A(n8069), .B(n8719), .Z(n8717) );
  NANDN U8310 ( .A(n8068), .B(n8066), .Z(n8719) );
  XOR U8311 ( .A(n8720), .B(n8721), .Z(n8066) );
  XNOR U8312 ( .A(n8722), .B(n8723), .Z(n8721) );
  ANDN U8313 ( .B(\stack[0][35] ), .A(n5243), .Z(n8068) );
  AND U8314 ( .A(n8724), .B(n8725), .Z(n8069) );
  NANDN U8315 ( .A(n8083), .B(n8726), .Z(n8724) );
  NANDN U8316 ( .A(n8082), .B(n8080), .Z(n8726) );
  XOR U8317 ( .A(n8727), .B(n8728), .Z(n8080) );
  XNOR U8318 ( .A(n8729), .B(n8730), .Z(n8728) );
  ANDN U8319 ( .B(\stack[1][3] ), .A(n5974), .Z(n8082) );
  AND U8320 ( .A(n8731), .B(n8732), .Z(n8083) );
  NANDN U8321 ( .A(n8094), .B(n8096), .Z(n8732) );
  NANDN U8322 ( .A(n8097), .B(n8733), .Z(n8731) );
  NANDN U8323 ( .A(n8096), .B(n8094), .Z(n8733) );
  XOR U8324 ( .A(n8734), .B(n8735), .Z(n8094) );
  XNOR U8325 ( .A(n8736), .B(n8737), .Z(n8735) );
  ANDN U8326 ( .B(\stack[0][33] ), .A(n5243), .Z(n8096) );
  AND U8327 ( .A(n8738), .B(n8739), .Z(n8097) );
  NANDN U8328 ( .A(n8111), .B(n8740), .Z(n8738) );
  NANDN U8329 ( .A(n8110), .B(n8108), .Z(n8740) );
  XOR U8330 ( .A(n8741), .B(n8742), .Z(n8108) );
  XNOR U8331 ( .A(n8743), .B(n8744), .Z(n8742) );
  ANDN U8332 ( .B(\stack[1][3] ), .A(n5926), .Z(n8110) );
  AND U8333 ( .A(n8745), .B(n8746), .Z(n8111) );
  NANDN U8334 ( .A(n8122), .B(n8124), .Z(n8746) );
  NANDN U8335 ( .A(n8125), .B(n8747), .Z(n8745) );
  NANDN U8336 ( .A(n8124), .B(n8122), .Z(n8747) );
  XOR U8337 ( .A(n8748), .B(n8749), .Z(n8122) );
  XNOR U8338 ( .A(n8750), .B(n8751), .Z(n8749) );
  ANDN U8339 ( .B(\stack[0][31] ), .A(n5243), .Z(n8124) );
  AND U8340 ( .A(n8752), .B(n8753), .Z(n8125) );
  NANDN U8341 ( .A(n8139), .B(n8754), .Z(n8752) );
  NANDN U8342 ( .A(n8138), .B(n8136), .Z(n8754) );
  XOR U8343 ( .A(n8755), .B(n8756), .Z(n8136) );
  XNOR U8344 ( .A(n8757), .B(n8758), .Z(n8756) );
  ANDN U8345 ( .B(\stack[1][3] ), .A(n5878), .Z(n8138) );
  AND U8346 ( .A(n8759), .B(n8760), .Z(n8139) );
  NANDN U8347 ( .A(n8150), .B(n8152), .Z(n8760) );
  NANDN U8348 ( .A(n8153), .B(n8761), .Z(n8759) );
  NANDN U8349 ( .A(n8152), .B(n8150), .Z(n8761) );
  XOR U8350 ( .A(n8762), .B(n8763), .Z(n8150) );
  XNOR U8351 ( .A(n8764), .B(n8765), .Z(n8763) );
  ANDN U8352 ( .B(\stack[0][29] ), .A(n5243), .Z(n8152) );
  AND U8353 ( .A(n8766), .B(n8767), .Z(n8153) );
  NANDN U8354 ( .A(n8167), .B(n8768), .Z(n8766) );
  NANDN U8355 ( .A(n8166), .B(n8164), .Z(n8768) );
  XOR U8356 ( .A(n8769), .B(n8770), .Z(n8164) );
  XNOR U8357 ( .A(n8771), .B(n8772), .Z(n8770) );
  ANDN U8358 ( .B(\stack[1][3] ), .A(n5830), .Z(n8166) );
  AND U8359 ( .A(n8773), .B(n8774), .Z(n8167) );
  NANDN U8360 ( .A(n8178), .B(n8180), .Z(n8774) );
  NANDN U8361 ( .A(n8181), .B(n8775), .Z(n8773) );
  NANDN U8362 ( .A(n8180), .B(n8178), .Z(n8775) );
  XOR U8363 ( .A(n8776), .B(n8777), .Z(n8178) );
  XNOR U8364 ( .A(n8778), .B(n8779), .Z(n8777) );
  ANDN U8365 ( .B(\stack[0][27] ), .A(n5243), .Z(n8180) );
  AND U8366 ( .A(n8780), .B(n8781), .Z(n8181) );
  NANDN U8367 ( .A(n8195), .B(n8782), .Z(n8780) );
  NANDN U8368 ( .A(n8194), .B(n8192), .Z(n8782) );
  XOR U8369 ( .A(n8783), .B(n8784), .Z(n8192) );
  XNOR U8370 ( .A(n8785), .B(n8786), .Z(n8784) );
  ANDN U8371 ( .B(\stack[1][3] ), .A(n5782), .Z(n8194) );
  AND U8372 ( .A(n8787), .B(n8788), .Z(n8195) );
  NANDN U8373 ( .A(n8206), .B(n8208), .Z(n8788) );
  NANDN U8374 ( .A(n8209), .B(n8789), .Z(n8787) );
  NANDN U8375 ( .A(n8208), .B(n8206), .Z(n8789) );
  XOR U8376 ( .A(n8790), .B(n8791), .Z(n8206) );
  XNOR U8377 ( .A(n8792), .B(n8793), .Z(n8791) );
  ANDN U8378 ( .B(\stack[0][25] ), .A(n5243), .Z(n8208) );
  AND U8379 ( .A(n8794), .B(n8795), .Z(n8209) );
  NANDN U8380 ( .A(n8223), .B(n8796), .Z(n8794) );
  NANDN U8381 ( .A(n8222), .B(n8220), .Z(n8796) );
  XOR U8382 ( .A(n8797), .B(n8798), .Z(n8220) );
  XNOR U8383 ( .A(n8799), .B(n8800), .Z(n8798) );
  ANDN U8384 ( .B(\stack[1][3] ), .A(n5734), .Z(n8222) );
  AND U8385 ( .A(n8801), .B(n8802), .Z(n8223) );
  NANDN U8386 ( .A(n8234), .B(n8236), .Z(n8802) );
  NANDN U8387 ( .A(n8237), .B(n8803), .Z(n8801) );
  NANDN U8388 ( .A(n8236), .B(n8234), .Z(n8803) );
  XOR U8389 ( .A(n8804), .B(n8805), .Z(n8234) );
  XNOR U8390 ( .A(n8806), .B(n8807), .Z(n8805) );
  ANDN U8391 ( .B(\stack[0][23] ), .A(n5243), .Z(n8236) );
  AND U8392 ( .A(n8808), .B(n8809), .Z(n8237) );
  NANDN U8393 ( .A(n8251), .B(n8810), .Z(n8808) );
  NANDN U8394 ( .A(n8250), .B(n8248), .Z(n8810) );
  XOR U8395 ( .A(n8811), .B(n8812), .Z(n8248) );
  XNOR U8396 ( .A(n8813), .B(n8814), .Z(n8812) );
  ANDN U8397 ( .B(\stack[1][3] ), .A(n5686), .Z(n8250) );
  AND U8398 ( .A(n8815), .B(n8816), .Z(n8251) );
  NANDN U8399 ( .A(n8262), .B(n8264), .Z(n8816) );
  NANDN U8400 ( .A(n8265), .B(n8817), .Z(n8815) );
  NANDN U8401 ( .A(n8264), .B(n8262), .Z(n8817) );
  XOR U8402 ( .A(n8818), .B(n8819), .Z(n8262) );
  XNOR U8403 ( .A(n8820), .B(n8821), .Z(n8819) );
  ANDN U8404 ( .B(\stack[0][21] ), .A(n5243), .Z(n8264) );
  AND U8405 ( .A(n8822), .B(n8823), .Z(n8265) );
  NANDN U8406 ( .A(n8279), .B(n8824), .Z(n8822) );
  NANDN U8407 ( .A(n8278), .B(n8276), .Z(n8824) );
  XOR U8408 ( .A(n8825), .B(n8826), .Z(n8276) );
  XNOR U8409 ( .A(n8827), .B(n8828), .Z(n8826) );
  ANDN U8410 ( .B(\stack[1][3] ), .A(n5638), .Z(n8278) );
  AND U8411 ( .A(n8829), .B(n8830), .Z(n8279) );
  NANDN U8412 ( .A(n8290), .B(n8292), .Z(n8830) );
  NANDN U8413 ( .A(n8293), .B(n8831), .Z(n8829) );
  NANDN U8414 ( .A(n8292), .B(n8290), .Z(n8831) );
  XOR U8415 ( .A(n8832), .B(n8833), .Z(n8290) );
  XNOR U8416 ( .A(n8834), .B(n8835), .Z(n8833) );
  ANDN U8417 ( .B(\stack[0][19] ), .A(n5243), .Z(n8292) );
  AND U8418 ( .A(n8836), .B(n8837), .Z(n8293) );
  NANDN U8419 ( .A(n8307), .B(n8838), .Z(n8836) );
  NANDN U8420 ( .A(n8306), .B(n8304), .Z(n8838) );
  XOR U8421 ( .A(n8839), .B(n8840), .Z(n8304) );
  XNOR U8422 ( .A(n8841), .B(n8842), .Z(n8840) );
  ANDN U8423 ( .B(\stack[1][3] ), .A(n5590), .Z(n8306) );
  AND U8424 ( .A(n8843), .B(n8844), .Z(n8307) );
  NANDN U8425 ( .A(n8318), .B(n8320), .Z(n8844) );
  NANDN U8426 ( .A(n8321), .B(n8845), .Z(n8843) );
  NANDN U8427 ( .A(n8320), .B(n8318), .Z(n8845) );
  XOR U8428 ( .A(n8846), .B(n8847), .Z(n8318) );
  XNOR U8429 ( .A(n8848), .B(n8849), .Z(n8847) );
  ANDN U8430 ( .B(\stack[0][17] ), .A(n5243), .Z(n8320) );
  AND U8431 ( .A(n8850), .B(n8851), .Z(n8321) );
  NANDN U8432 ( .A(n8335), .B(n8852), .Z(n8850) );
  NANDN U8433 ( .A(n8334), .B(n8332), .Z(n8852) );
  XOR U8434 ( .A(n8853), .B(n8854), .Z(n8332) );
  XNOR U8435 ( .A(n8855), .B(n8856), .Z(n8854) );
  ANDN U8436 ( .B(\stack[1][3] ), .A(n5542), .Z(n8334) );
  AND U8437 ( .A(n8857), .B(n8858), .Z(n8335) );
  NANDN U8438 ( .A(n8346), .B(n8348), .Z(n8858) );
  NANDN U8439 ( .A(n8349), .B(n8859), .Z(n8857) );
  NANDN U8440 ( .A(n8348), .B(n8346), .Z(n8859) );
  XOR U8441 ( .A(n8860), .B(n8861), .Z(n8346) );
  XNOR U8442 ( .A(n8862), .B(n8863), .Z(n8861) );
  ANDN U8443 ( .B(\stack[0][15] ), .A(n5243), .Z(n8348) );
  AND U8444 ( .A(n8864), .B(n8865), .Z(n8349) );
  NANDN U8445 ( .A(n8363), .B(n8866), .Z(n8864) );
  NANDN U8446 ( .A(n8362), .B(n8360), .Z(n8866) );
  XOR U8447 ( .A(n8867), .B(n8868), .Z(n8360) );
  XNOR U8448 ( .A(n8869), .B(n8870), .Z(n8868) );
  ANDN U8449 ( .B(\stack[1][3] ), .A(n5494), .Z(n8362) );
  AND U8450 ( .A(n8871), .B(n8872), .Z(n8363) );
  NANDN U8451 ( .A(n8374), .B(n8376), .Z(n8872) );
  NANDN U8452 ( .A(n8377), .B(n8873), .Z(n8871) );
  NANDN U8453 ( .A(n8376), .B(n8374), .Z(n8873) );
  XOR U8454 ( .A(n8874), .B(n8875), .Z(n8374) );
  XNOR U8455 ( .A(n8876), .B(n8877), .Z(n8875) );
  ANDN U8456 ( .B(\stack[0][13] ), .A(n5243), .Z(n8376) );
  AND U8457 ( .A(n8878), .B(n8879), .Z(n8377) );
  NANDN U8458 ( .A(n8391), .B(n8880), .Z(n8878) );
  NANDN U8459 ( .A(n8390), .B(n8388), .Z(n8880) );
  XOR U8460 ( .A(n8881), .B(n8882), .Z(n8388) );
  XNOR U8461 ( .A(n8883), .B(n8884), .Z(n8882) );
  ANDN U8462 ( .B(\stack[1][3] ), .A(n5446), .Z(n8390) );
  AND U8463 ( .A(n8885), .B(n8886), .Z(n8391) );
  NANDN U8464 ( .A(n8402), .B(n8404), .Z(n8886) );
  NANDN U8465 ( .A(n8405), .B(n8887), .Z(n8885) );
  NANDN U8466 ( .A(n8404), .B(n8402), .Z(n8887) );
  XOR U8467 ( .A(n8888), .B(n8889), .Z(n8402) );
  XNOR U8468 ( .A(n8890), .B(n8891), .Z(n8889) );
  ANDN U8469 ( .B(\stack[0][11] ), .A(n5243), .Z(n8404) );
  AND U8470 ( .A(n8892), .B(n8893), .Z(n8405) );
  NANDN U8471 ( .A(n8419), .B(n8894), .Z(n8892) );
  NANDN U8472 ( .A(n8418), .B(n8416), .Z(n8894) );
  XOR U8473 ( .A(n8895), .B(n8896), .Z(n8416) );
  XNOR U8474 ( .A(n8897), .B(n8898), .Z(n8896) );
  ANDN U8475 ( .B(\stack[1][3] ), .A(n5398), .Z(n8418) );
  AND U8476 ( .A(n8899), .B(n8900), .Z(n8419) );
  NANDN U8477 ( .A(n8430), .B(n8432), .Z(n8900) );
  NANDN U8478 ( .A(n8433), .B(n8901), .Z(n8899) );
  NANDN U8479 ( .A(n8432), .B(n8430), .Z(n8901) );
  XOR U8480 ( .A(n8902), .B(n8903), .Z(n8430) );
  XNOR U8481 ( .A(n8904), .B(n8905), .Z(n8903) );
  ANDN U8482 ( .B(\stack[1][3] ), .A(n5374), .Z(n8432) );
  AND U8483 ( .A(n8906), .B(n8907), .Z(n8433) );
  NANDN U8484 ( .A(n8447), .B(n8908), .Z(n8906) );
  NANDN U8485 ( .A(n8446), .B(n8444), .Z(n8908) );
  XOR U8486 ( .A(n8909), .B(n8910), .Z(n8444) );
  XNOR U8487 ( .A(n8911), .B(n8912), .Z(n8910) );
  ANDN U8488 ( .B(\stack[1][3] ), .A(n5350), .Z(n8446) );
  AND U8489 ( .A(n8913), .B(n8914), .Z(n8447) );
  NANDN U8490 ( .A(n8459), .B(n8461), .Z(n8914) );
  NANDN U8491 ( .A(n8462), .B(n8915), .Z(n8913) );
  NANDN U8492 ( .A(n8461), .B(n8459), .Z(n8915) );
  XOR U8493 ( .A(n8916), .B(n8917), .Z(n8459) );
  XNOR U8494 ( .A(n8918), .B(n8919), .Z(n8917) );
  ANDN U8495 ( .B(\stack[0][7] ), .A(n5243), .Z(n8461) );
  AND U8496 ( .A(n8920), .B(n8921), .Z(n8462) );
  NANDN U8497 ( .A(n8474), .B(n8476), .Z(n8921) );
  NANDN U8498 ( .A(n8477), .B(n8922), .Z(n8920) );
  NANDN U8499 ( .A(n8476), .B(n8474), .Z(n8922) );
  XNOR U8500 ( .A(n8923), .B(n8924), .Z(n8474) );
  XOR U8501 ( .A(n8925), .B(n8926), .Z(n8924) );
  AND U8502 ( .A(\stack[0][6] ), .B(\stack[1][3] ), .Z(n8476) );
  AND U8503 ( .A(n8927), .B(n8928), .Z(n8477) );
  NANDN U8504 ( .A(n8488), .B(n8490), .Z(n8928) );
  NANDN U8505 ( .A(n8491), .B(n8929), .Z(n8927) );
  NANDN U8506 ( .A(n8490), .B(n8488), .Z(n8929) );
  XOR U8507 ( .A(n8930), .B(n8931), .Z(n8488) );
  XNOR U8508 ( .A(n8932), .B(n8933), .Z(n8931) );
  ANDN U8509 ( .B(\stack[1][3] ), .A(n5278), .Z(n8490) );
  AND U8510 ( .A(n8934), .B(n8935), .Z(n8491) );
  NANDN U8511 ( .A(n8505), .B(n8936), .Z(n8934) );
  NANDN U8512 ( .A(n8504), .B(n8502), .Z(n8936) );
  XOR U8513 ( .A(n8937), .B(n8938), .Z(n8502) );
  XNOR U8514 ( .A(n8939), .B(n8940), .Z(n8938) );
  ANDN U8515 ( .B(\stack[0][4] ), .A(n5243), .Z(n8504) );
  AND U8516 ( .A(n8941), .B(n8942), .Z(n8505) );
  NANDN U8517 ( .A(n8516), .B(n8518), .Z(n8942) );
  NANDN U8518 ( .A(n8519), .B(n8943), .Z(n8941) );
  NANDN U8519 ( .A(n8518), .B(n8516), .Z(n8943) );
  XNOR U8520 ( .A(n8944), .B(n8945), .Z(n8516) );
  XNOR U8521 ( .A(n8946), .B(n8947), .Z(n8945) );
  ANDN U8522 ( .B(\stack[1][3] ), .A(n5230), .Z(n8518) );
  AND U8523 ( .A(n8948), .B(n8949), .Z(n8519) );
  NANDN U8524 ( .A(n8530), .B(n8532), .Z(n8949) );
  NAND U8525 ( .A(n8950), .B(n8533), .Z(n8948) );
  ANDN U8526 ( .B(n8951), .A(n8540), .Z(n8533) );
  NANDN U8527 ( .A(n5243), .B(\stack[0][1] ), .Z(n8540) );
  ANDN U8528 ( .B(\stack[0][0] ), .A(n5267), .Z(n8951) );
  NANDN U8529 ( .A(n8532), .B(n8530), .Z(n8950) );
  XNOR U8530 ( .A(n8952), .B(n8953), .Z(n8530) );
  NANDN U8531 ( .A(n5160), .B(\stack[1][5] ), .Z(n8953) );
  ANDN U8532 ( .B(\stack[1][3] ), .A(n5206), .Z(n8532) );
  ANDN U8533 ( .B(\stack[1][3] ), .A(n6598), .Z(n8547) );
  XOR U8534 ( .A(n8954), .B(n8955), .Z(n7117) );
  XOR U8535 ( .A(n8956), .B(n8957), .Z(n8955) );
  AND U8536 ( .A(n8958), .B(n8959), .Z(n8957) );
  NANDN U8537 ( .A(n8555), .B(n8960), .Z(n8958) );
  NANDN U8538 ( .A(n8554), .B(n8552), .Z(n8960) );
  XOR U8539 ( .A(n8961), .B(n8962), .Z(n8552) );
  XNOR U8540 ( .A(n8963), .B(n8964), .Z(n8962) );
  ANDN U8541 ( .B(\stack[1][4] ), .A(n6550), .Z(n8554) );
  AND U8542 ( .A(n8965), .B(n8966), .Z(n8555) );
  NANDN U8543 ( .A(n8559), .B(n8561), .Z(n8966) );
  NANDN U8544 ( .A(n8562), .B(n8967), .Z(n8965) );
  NANDN U8545 ( .A(n8561), .B(n8559), .Z(n8967) );
  XOR U8546 ( .A(n8968), .B(n8969), .Z(n8559) );
  XNOR U8547 ( .A(n8970), .B(n8971), .Z(n8969) );
  ANDN U8548 ( .B(\stack[0][57] ), .A(n5267), .Z(n8561) );
  AND U8549 ( .A(n8972), .B(n8973), .Z(n8562) );
  NANDN U8550 ( .A(n8569), .B(n8974), .Z(n8972) );
  NANDN U8551 ( .A(n8568), .B(n8566), .Z(n8974) );
  XOR U8552 ( .A(n8975), .B(n8976), .Z(n8566) );
  XNOR U8553 ( .A(n8977), .B(n8978), .Z(n8976) );
  ANDN U8554 ( .B(\stack[1][4] ), .A(n6502), .Z(n8568) );
  AND U8555 ( .A(n8979), .B(n8980), .Z(n8569) );
  NANDN U8556 ( .A(n8573), .B(n8575), .Z(n8980) );
  NANDN U8557 ( .A(n8576), .B(n8981), .Z(n8979) );
  NANDN U8558 ( .A(n8575), .B(n8573), .Z(n8981) );
  XOR U8559 ( .A(n8982), .B(n8983), .Z(n8573) );
  XNOR U8560 ( .A(n8984), .B(n8985), .Z(n8983) );
  ANDN U8561 ( .B(\stack[0][55] ), .A(n5267), .Z(n8575) );
  AND U8562 ( .A(n8986), .B(n8987), .Z(n8576) );
  OR U8563 ( .A(n8580), .B(n8988), .Z(n8987) );
  IV U8564 ( .A(n8582), .Z(n8988) );
  NANDN U8565 ( .A(n8583), .B(n8989), .Z(n8986) );
  NANDN U8566 ( .A(n8582), .B(n8580), .Z(n8989) );
  XOR U8567 ( .A(n8990), .B(n8991), .Z(n8580) );
  XNOR U8568 ( .A(n8992), .B(n8993), .Z(n8991) );
  ANDN U8569 ( .B(\stack[1][4] ), .A(n6454), .Z(n8582) );
  AND U8570 ( .A(n8994), .B(n8995), .Z(n8583) );
  NANDN U8571 ( .A(n8587), .B(n8589), .Z(n8995) );
  NANDN U8572 ( .A(n8590), .B(n8996), .Z(n8994) );
  NANDN U8573 ( .A(n8589), .B(n8587), .Z(n8996) );
  XOR U8574 ( .A(n8997), .B(n8998), .Z(n8587) );
  XNOR U8575 ( .A(n8999), .B(n9000), .Z(n8998) );
  ANDN U8576 ( .B(\stack[0][53] ), .A(n5267), .Z(n8589) );
  AND U8577 ( .A(n9001), .B(n9002), .Z(n8590) );
  NANDN U8578 ( .A(n8597), .B(n9003), .Z(n9001) );
  NANDN U8579 ( .A(n8596), .B(n8594), .Z(n9003) );
  XOR U8580 ( .A(n9004), .B(n9005), .Z(n8594) );
  XNOR U8581 ( .A(n9006), .B(n9007), .Z(n9005) );
  ANDN U8582 ( .B(\stack[1][4] ), .A(n6406), .Z(n8596) );
  AND U8583 ( .A(n9008), .B(n9009), .Z(n8597) );
  NANDN U8584 ( .A(n8601), .B(n8603), .Z(n9009) );
  NANDN U8585 ( .A(n8604), .B(n9010), .Z(n9008) );
  NANDN U8586 ( .A(n8603), .B(n8601), .Z(n9010) );
  XOR U8587 ( .A(n9011), .B(n9012), .Z(n8601) );
  XNOR U8588 ( .A(n9013), .B(n9014), .Z(n9012) );
  ANDN U8589 ( .B(\stack[0][51] ), .A(n5267), .Z(n8603) );
  AND U8590 ( .A(n9015), .B(n9016), .Z(n8604) );
  NANDN U8591 ( .A(n8611), .B(n9017), .Z(n9015) );
  NANDN U8592 ( .A(n8610), .B(n8608), .Z(n9017) );
  XOR U8593 ( .A(n9018), .B(n9019), .Z(n8608) );
  XNOR U8594 ( .A(n9020), .B(n9021), .Z(n9019) );
  ANDN U8595 ( .B(\stack[1][4] ), .A(n6358), .Z(n8610) );
  AND U8596 ( .A(n9022), .B(n9023), .Z(n8611) );
  NANDN U8597 ( .A(n8615), .B(n8617), .Z(n9023) );
  NANDN U8598 ( .A(n8618), .B(n9024), .Z(n9022) );
  NANDN U8599 ( .A(n8617), .B(n8615), .Z(n9024) );
  XOR U8600 ( .A(n9025), .B(n9026), .Z(n8615) );
  XNOR U8601 ( .A(n9027), .B(n9028), .Z(n9026) );
  ANDN U8602 ( .B(\stack[0][49] ), .A(n5267), .Z(n8617) );
  AND U8603 ( .A(n9029), .B(n9030), .Z(n8618) );
  NANDN U8604 ( .A(n8625), .B(n9031), .Z(n9029) );
  NANDN U8605 ( .A(n8624), .B(n8622), .Z(n9031) );
  XOR U8606 ( .A(n9032), .B(n9033), .Z(n8622) );
  XNOR U8607 ( .A(n9034), .B(n9035), .Z(n9033) );
  ANDN U8608 ( .B(\stack[1][4] ), .A(n6310), .Z(n8624) );
  AND U8609 ( .A(n9036), .B(n9037), .Z(n8625) );
  NANDN U8610 ( .A(n8629), .B(n8631), .Z(n9037) );
  NANDN U8611 ( .A(n8632), .B(n9038), .Z(n9036) );
  NANDN U8612 ( .A(n8631), .B(n8629), .Z(n9038) );
  XOR U8613 ( .A(n9039), .B(n9040), .Z(n8629) );
  XNOR U8614 ( .A(n9041), .B(n9042), .Z(n9040) );
  ANDN U8615 ( .B(\stack[0][47] ), .A(n5267), .Z(n8631) );
  AND U8616 ( .A(n9043), .B(n9044), .Z(n8632) );
  NANDN U8617 ( .A(n8639), .B(n9045), .Z(n9043) );
  NANDN U8618 ( .A(n8638), .B(n8636), .Z(n9045) );
  XOR U8619 ( .A(n9046), .B(n9047), .Z(n8636) );
  XNOR U8620 ( .A(n9048), .B(n9049), .Z(n9047) );
  ANDN U8621 ( .B(\stack[1][4] ), .A(n6262), .Z(n8638) );
  AND U8622 ( .A(n9050), .B(n9051), .Z(n8639) );
  NANDN U8623 ( .A(n8643), .B(n8645), .Z(n9051) );
  NANDN U8624 ( .A(n8646), .B(n9052), .Z(n9050) );
  NANDN U8625 ( .A(n8645), .B(n8643), .Z(n9052) );
  XOR U8626 ( .A(n9053), .B(n9054), .Z(n8643) );
  XNOR U8627 ( .A(n9055), .B(n9056), .Z(n9054) );
  ANDN U8628 ( .B(\stack[0][45] ), .A(n5267), .Z(n8645) );
  AND U8629 ( .A(n9057), .B(n9058), .Z(n8646) );
  NANDN U8630 ( .A(n8653), .B(n9059), .Z(n9057) );
  NANDN U8631 ( .A(n8652), .B(n8650), .Z(n9059) );
  XOR U8632 ( .A(n9060), .B(n9061), .Z(n8650) );
  XNOR U8633 ( .A(n9062), .B(n9063), .Z(n9061) );
  ANDN U8634 ( .B(\stack[1][4] ), .A(n6214), .Z(n8652) );
  AND U8635 ( .A(n9064), .B(n9065), .Z(n8653) );
  NANDN U8636 ( .A(n8657), .B(n8659), .Z(n9065) );
  NANDN U8637 ( .A(n8660), .B(n9066), .Z(n9064) );
  NANDN U8638 ( .A(n8659), .B(n8657), .Z(n9066) );
  XOR U8639 ( .A(n9067), .B(n9068), .Z(n8657) );
  XNOR U8640 ( .A(n9069), .B(n9070), .Z(n9068) );
  ANDN U8641 ( .B(\stack[0][43] ), .A(n5267), .Z(n8659) );
  AND U8642 ( .A(n9071), .B(n9072), .Z(n8660) );
  NANDN U8643 ( .A(n8667), .B(n9073), .Z(n9071) );
  NANDN U8644 ( .A(n8666), .B(n8664), .Z(n9073) );
  XOR U8645 ( .A(n9074), .B(n9075), .Z(n8664) );
  XNOR U8646 ( .A(n9076), .B(n9077), .Z(n9075) );
  ANDN U8647 ( .B(\stack[1][4] ), .A(n6166), .Z(n8666) );
  AND U8648 ( .A(n9078), .B(n9079), .Z(n8667) );
  NANDN U8649 ( .A(n8671), .B(n8673), .Z(n9079) );
  NANDN U8650 ( .A(n8674), .B(n9080), .Z(n9078) );
  NANDN U8651 ( .A(n8673), .B(n8671), .Z(n9080) );
  XOR U8652 ( .A(n9081), .B(n9082), .Z(n8671) );
  XNOR U8653 ( .A(n9083), .B(n9084), .Z(n9082) );
  ANDN U8654 ( .B(\stack[0][41] ), .A(n5267), .Z(n8673) );
  AND U8655 ( .A(n9085), .B(n9086), .Z(n8674) );
  NANDN U8656 ( .A(n8681), .B(n9087), .Z(n9085) );
  NANDN U8657 ( .A(n8680), .B(n8678), .Z(n9087) );
  XOR U8658 ( .A(n9088), .B(n9089), .Z(n8678) );
  XNOR U8659 ( .A(n9090), .B(n9091), .Z(n9089) );
  ANDN U8660 ( .B(\stack[1][4] ), .A(n6118), .Z(n8680) );
  AND U8661 ( .A(n9092), .B(n9093), .Z(n8681) );
  NANDN U8662 ( .A(n8685), .B(n8687), .Z(n9093) );
  NANDN U8663 ( .A(n8688), .B(n9094), .Z(n9092) );
  NANDN U8664 ( .A(n8687), .B(n8685), .Z(n9094) );
  XOR U8665 ( .A(n9095), .B(n9096), .Z(n8685) );
  XNOR U8666 ( .A(n9097), .B(n9098), .Z(n9096) );
  ANDN U8667 ( .B(\stack[0][39] ), .A(n5267), .Z(n8687) );
  AND U8668 ( .A(n9099), .B(n9100), .Z(n8688) );
  NANDN U8669 ( .A(n8695), .B(n9101), .Z(n9099) );
  NANDN U8670 ( .A(n8694), .B(n8692), .Z(n9101) );
  XOR U8671 ( .A(n9102), .B(n9103), .Z(n8692) );
  XNOR U8672 ( .A(n9104), .B(n9105), .Z(n9103) );
  ANDN U8673 ( .B(\stack[1][4] ), .A(n6070), .Z(n8694) );
  AND U8674 ( .A(n9106), .B(n9107), .Z(n8695) );
  NANDN U8675 ( .A(n8699), .B(n8701), .Z(n9107) );
  NANDN U8676 ( .A(n8702), .B(n9108), .Z(n9106) );
  NANDN U8677 ( .A(n8701), .B(n8699), .Z(n9108) );
  XOR U8678 ( .A(n9109), .B(n9110), .Z(n8699) );
  XNOR U8679 ( .A(n9111), .B(n9112), .Z(n9110) );
  ANDN U8680 ( .B(\stack[0][37] ), .A(n5267), .Z(n8701) );
  AND U8681 ( .A(n9113), .B(n9114), .Z(n8702) );
  NANDN U8682 ( .A(n8709), .B(n9115), .Z(n9113) );
  NANDN U8683 ( .A(n8708), .B(n8706), .Z(n9115) );
  XOR U8684 ( .A(n9116), .B(n9117), .Z(n8706) );
  XNOR U8685 ( .A(n9118), .B(n9119), .Z(n9117) );
  ANDN U8686 ( .B(\stack[1][4] ), .A(n6022), .Z(n8708) );
  AND U8687 ( .A(n9120), .B(n9121), .Z(n8709) );
  NANDN U8688 ( .A(n8713), .B(n8715), .Z(n9121) );
  NANDN U8689 ( .A(n8716), .B(n9122), .Z(n9120) );
  NANDN U8690 ( .A(n8715), .B(n8713), .Z(n9122) );
  XOR U8691 ( .A(n9123), .B(n9124), .Z(n8713) );
  XNOR U8692 ( .A(n9125), .B(n9126), .Z(n9124) );
  ANDN U8693 ( .B(\stack[0][35] ), .A(n5267), .Z(n8715) );
  AND U8694 ( .A(n9127), .B(n9128), .Z(n8716) );
  NANDN U8695 ( .A(n8723), .B(n9129), .Z(n9127) );
  NANDN U8696 ( .A(n8722), .B(n8720), .Z(n9129) );
  XOR U8697 ( .A(n9130), .B(n9131), .Z(n8720) );
  XNOR U8698 ( .A(n9132), .B(n9133), .Z(n9131) );
  ANDN U8699 ( .B(\stack[1][4] ), .A(n5974), .Z(n8722) );
  AND U8700 ( .A(n9134), .B(n9135), .Z(n8723) );
  NANDN U8701 ( .A(n8727), .B(n8729), .Z(n9135) );
  NANDN U8702 ( .A(n8730), .B(n9136), .Z(n9134) );
  NANDN U8703 ( .A(n8729), .B(n8727), .Z(n9136) );
  XOR U8704 ( .A(n9137), .B(n9138), .Z(n8727) );
  XNOR U8705 ( .A(n9139), .B(n9140), .Z(n9138) );
  ANDN U8706 ( .B(\stack[0][33] ), .A(n5267), .Z(n8729) );
  AND U8707 ( .A(n9141), .B(n9142), .Z(n8730) );
  NANDN U8708 ( .A(n8737), .B(n9143), .Z(n9141) );
  NANDN U8709 ( .A(n8736), .B(n8734), .Z(n9143) );
  XOR U8710 ( .A(n9144), .B(n9145), .Z(n8734) );
  XNOR U8711 ( .A(n9146), .B(n9147), .Z(n9145) );
  ANDN U8712 ( .B(\stack[1][4] ), .A(n5926), .Z(n8736) );
  AND U8713 ( .A(n9148), .B(n9149), .Z(n8737) );
  NANDN U8714 ( .A(n8741), .B(n8743), .Z(n9149) );
  NANDN U8715 ( .A(n8744), .B(n9150), .Z(n9148) );
  NANDN U8716 ( .A(n8743), .B(n8741), .Z(n9150) );
  XOR U8717 ( .A(n9151), .B(n9152), .Z(n8741) );
  XNOR U8718 ( .A(n9153), .B(n9154), .Z(n9152) );
  ANDN U8719 ( .B(\stack[0][31] ), .A(n5267), .Z(n8743) );
  AND U8720 ( .A(n9155), .B(n9156), .Z(n8744) );
  NANDN U8721 ( .A(n8751), .B(n9157), .Z(n9155) );
  NANDN U8722 ( .A(n8750), .B(n8748), .Z(n9157) );
  XOR U8723 ( .A(n9158), .B(n9159), .Z(n8748) );
  XNOR U8724 ( .A(n9160), .B(n9161), .Z(n9159) );
  ANDN U8725 ( .B(\stack[1][4] ), .A(n5878), .Z(n8750) );
  AND U8726 ( .A(n9162), .B(n9163), .Z(n8751) );
  NANDN U8727 ( .A(n8755), .B(n8757), .Z(n9163) );
  NANDN U8728 ( .A(n8758), .B(n9164), .Z(n9162) );
  NANDN U8729 ( .A(n8757), .B(n8755), .Z(n9164) );
  XOR U8730 ( .A(n9165), .B(n9166), .Z(n8755) );
  XNOR U8731 ( .A(n9167), .B(n9168), .Z(n9166) );
  ANDN U8732 ( .B(\stack[0][29] ), .A(n5267), .Z(n8757) );
  AND U8733 ( .A(n9169), .B(n9170), .Z(n8758) );
  NANDN U8734 ( .A(n8765), .B(n9171), .Z(n9169) );
  NANDN U8735 ( .A(n8764), .B(n8762), .Z(n9171) );
  XOR U8736 ( .A(n9172), .B(n9173), .Z(n8762) );
  XNOR U8737 ( .A(n9174), .B(n9175), .Z(n9173) );
  ANDN U8738 ( .B(\stack[1][4] ), .A(n5830), .Z(n8764) );
  AND U8739 ( .A(n9176), .B(n9177), .Z(n8765) );
  NANDN U8740 ( .A(n8769), .B(n8771), .Z(n9177) );
  NANDN U8741 ( .A(n8772), .B(n9178), .Z(n9176) );
  NANDN U8742 ( .A(n8771), .B(n8769), .Z(n9178) );
  XOR U8743 ( .A(n9179), .B(n9180), .Z(n8769) );
  XNOR U8744 ( .A(n9181), .B(n9182), .Z(n9180) );
  ANDN U8745 ( .B(\stack[0][27] ), .A(n5267), .Z(n8771) );
  AND U8746 ( .A(n9183), .B(n9184), .Z(n8772) );
  NANDN U8747 ( .A(n8779), .B(n9185), .Z(n9183) );
  NANDN U8748 ( .A(n8778), .B(n8776), .Z(n9185) );
  XOR U8749 ( .A(n9186), .B(n9187), .Z(n8776) );
  XNOR U8750 ( .A(n9188), .B(n9189), .Z(n9187) );
  ANDN U8751 ( .B(\stack[1][4] ), .A(n5782), .Z(n8778) );
  AND U8752 ( .A(n9190), .B(n9191), .Z(n8779) );
  NANDN U8753 ( .A(n8783), .B(n8785), .Z(n9191) );
  NANDN U8754 ( .A(n8786), .B(n9192), .Z(n9190) );
  NANDN U8755 ( .A(n8785), .B(n8783), .Z(n9192) );
  XOR U8756 ( .A(n9193), .B(n9194), .Z(n8783) );
  XNOR U8757 ( .A(n9195), .B(n9196), .Z(n9194) );
  ANDN U8758 ( .B(\stack[0][25] ), .A(n5267), .Z(n8785) );
  AND U8759 ( .A(n9197), .B(n9198), .Z(n8786) );
  NANDN U8760 ( .A(n8793), .B(n9199), .Z(n9197) );
  NANDN U8761 ( .A(n8792), .B(n8790), .Z(n9199) );
  XOR U8762 ( .A(n9200), .B(n9201), .Z(n8790) );
  XNOR U8763 ( .A(n9202), .B(n9203), .Z(n9201) );
  ANDN U8764 ( .B(\stack[1][4] ), .A(n5734), .Z(n8792) );
  AND U8765 ( .A(n9204), .B(n9205), .Z(n8793) );
  NANDN U8766 ( .A(n8797), .B(n8799), .Z(n9205) );
  NANDN U8767 ( .A(n8800), .B(n9206), .Z(n9204) );
  NANDN U8768 ( .A(n8799), .B(n8797), .Z(n9206) );
  XOR U8769 ( .A(n9207), .B(n9208), .Z(n8797) );
  XNOR U8770 ( .A(n9209), .B(n9210), .Z(n9208) );
  ANDN U8771 ( .B(\stack[0][23] ), .A(n5267), .Z(n8799) );
  AND U8772 ( .A(n9211), .B(n9212), .Z(n8800) );
  NANDN U8773 ( .A(n8807), .B(n9213), .Z(n9211) );
  NANDN U8774 ( .A(n8806), .B(n8804), .Z(n9213) );
  XOR U8775 ( .A(n9214), .B(n9215), .Z(n8804) );
  XNOR U8776 ( .A(n9216), .B(n9217), .Z(n9215) );
  ANDN U8777 ( .B(\stack[1][4] ), .A(n5686), .Z(n8806) );
  AND U8778 ( .A(n9218), .B(n9219), .Z(n8807) );
  NANDN U8779 ( .A(n8811), .B(n8813), .Z(n9219) );
  NANDN U8780 ( .A(n8814), .B(n9220), .Z(n9218) );
  NANDN U8781 ( .A(n8813), .B(n8811), .Z(n9220) );
  XOR U8782 ( .A(n9221), .B(n9222), .Z(n8811) );
  XNOR U8783 ( .A(n9223), .B(n9224), .Z(n9222) );
  ANDN U8784 ( .B(\stack[0][21] ), .A(n5267), .Z(n8813) );
  AND U8785 ( .A(n9225), .B(n9226), .Z(n8814) );
  NANDN U8786 ( .A(n8821), .B(n9227), .Z(n9225) );
  NANDN U8787 ( .A(n8820), .B(n8818), .Z(n9227) );
  XOR U8788 ( .A(n9228), .B(n9229), .Z(n8818) );
  XNOR U8789 ( .A(n9230), .B(n9231), .Z(n9229) );
  ANDN U8790 ( .B(\stack[1][4] ), .A(n5638), .Z(n8820) );
  AND U8791 ( .A(n9232), .B(n9233), .Z(n8821) );
  NANDN U8792 ( .A(n8825), .B(n8827), .Z(n9233) );
  NANDN U8793 ( .A(n8828), .B(n9234), .Z(n9232) );
  NANDN U8794 ( .A(n8827), .B(n8825), .Z(n9234) );
  XOR U8795 ( .A(n9235), .B(n9236), .Z(n8825) );
  XNOR U8796 ( .A(n9237), .B(n9238), .Z(n9236) );
  ANDN U8797 ( .B(\stack[0][19] ), .A(n5267), .Z(n8827) );
  AND U8798 ( .A(n9239), .B(n9240), .Z(n8828) );
  NANDN U8799 ( .A(n8835), .B(n9241), .Z(n9239) );
  NANDN U8800 ( .A(n8834), .B(n8832), .Z(n9241) );
  XOR U8801 ( .A(n9242), .B(n9243), .Z(n8832) );
  XNOR U8802 ( .A(n9244), .B(n9245), .Z(n9243) );
  ANDN U8803 ( .B(\stack[1][4] ), .A(n5590), .Z(n8834) );
  AND U8804 ( .A(n9246), .B(n9247), .Z(n8835) );
  NANDN U8805 ( .A(n8839), .B(n8841), .Z(n9247) );
  NANDN U8806 ( .A(n8842), .B(n9248), .Z(n9246) );
  NANDN U8807 ( .A(n8841), .B(n8839), .Z(n9248) );
  XOR U8808 ( .A(n9249), .B(n9250), .Z(n8839) );
  XNOR U8809 ( .A(n9251), .B(n9252), .Z(n9250) );
  ANDN U8810 ( .B(\stack[0][17] ), .A(n5267), .Z(n8841) );
  AND U8811 ( .A(n9253), .B(n9254), .Z(n8842) );
  NANDN U8812 ( .A(n8849), .B(n9255), .Z(n9253) );
  NANDN U8813 ( .A(n8848), .B(n8846), .Z(n9255) );
  XOR U8814 ( .A(n9256), .B(n9257), .Z(n8846) );
  XNOR U8815 ( .A(n9258), .B(n9259), .Z(n9257) );
  ANDN U8816 ( .B(\stack[1][4] ), .A(n5542), .Z(n8848) );
  AND U8817 ( .A(n9260), .B(n9261), .Z(n8849) );
  NANDN U8818 ( .A(n8853), .B(n8855), .Z(n9261) );
  NANDN U8819 ( .A(n8856), .B(n9262), .Z(n9260) );
  NANDN U8820 ( .A(n8855), .B(n8853), .Z(n9262) );
  XOR U8821 ( .A(n9263), .B(n9264), .Z(n8853) );
  XNOR U8822 ( .A(n9265), .B(n9266), .Z(n9264) );
  ANDN U8823 ( .B(\stack[0][15] ), .A(n5267), .Z(n8855) );
  AND U8824 ( .A(n9267), .B(n9268), .Z(n8856) );
  NANDN U8825 ( .A(n8863), .B(n9269), .Z(n9267) );
  NANDN U8826 ( .A(n8862), .B(n8860), .Z(n9269) );
  XOR U8827 ( .A(n9270), .B(n9271), .Z(n8860) );
  XNOR U8828 ( .A(n9272), .B(n9273), .Z(n9271) );
  ANDN U8829 ( .B(\stack[1][4] ), .A(n5494), .Z(n8862) );
  AND U8830 ( .A(n9274), .B(n9275), .Z(n8863) );
  NANDN U8831 ( .A(n8867), .B(n8869), .Z(n9275) );
  NANDN U8832 ( .A(n8870), .B(n9276), .Z(n9274) );
  NANDN U8833 ( .A(n8869), .B(n8867), .Z(n9276) );
  XOR U8834 ( .A(n9277), .B(n9278), .Z(n8867) );
  XNOR U8835 ( .A(n9279), .B(n9280), .Z(n9278) );
  ANDN U8836 ( .B(\stack[0][13] ), .A(n5267), .Z(n8869) );
  AND U8837 ( .A(n9281), .B(n9282), .Z(n8870) );
  NANDN U8838 ( .A(n8877), .B(n9283), .Z(n9281) );
  NANDN U8839 ( .A(n8876), .B(n8874), .Z(n9283) );
  XOR U8840 ( .A(n9284), .B(n9285), .Z(n8874) );
  XNOR U8841 ( .A(n9286), .B(n9287), .Z(n9285) );
  ANDN U8842 ( .B(\stack[1][4] ), .A(n5446), .Z(n8876) );
  AND U8843 ( .A(n9288), .B(n9289), .Z(n8877) );
  NANDN U8844 ( .A(n8881), .B(n8883), .Z(n9289) );
  NANDN U8845 ( .A(n8884), .B(n9290), .Z(n9288) );
  NANDN U8846 ( .A(n8883), .B(n8881), .Z(n9290) );
  XOR U8847 ( .A(n9291), .B(n9292), .Z(n8881) );
  XNOR U8848 ( .A(n9293), .B(n9294), .Z(n9292) );
  ANDN U8849 ( .B(\stack[0][11] ), .A(n5267), .Z(n8883) );
  AND U8850 ( .A(n9295), .B(n9296), .Z(n8884) );
  NANDN U8851 ( .A(n8891), .B(n9297), .Z(n9295) );
  NANDN U8852 ( .A(n8890), .B(n8888), .Z(n9297) );
  XOR U8853 ( .A(n9298), .B(n9299), .Z(n8888) );
  XNOR U8854 ( .A(n9300), .B(n9301), .Z(n9299) );
  ANDN U8855 ( .B(\stack[1][4] ), .A(n5398), .Z(n8890) );
  AND U8856 ( .A(n9302), .B(n9303), .Z(n8891) );
  NANDN U8857 ( .A(n8895), .B(n8897), .Z(n9303) );
  NANDN U8858 ( .A(n8898), .B(n9304), .Z(n9302) );
  NANDN U8859 ( .A(n8897), .B(n8895), .Z(n9304) );
  XOR U8860 ( .A(n9305), .B(n9306), .Z(n8895) );
  XNOR U8861 ( .A(n9307), .B(n9308), .Z(n9306) );
  ANDN U8862 ( .B(\stack[1][4] ), .A(n5374), .Z(n8897) );
  AND U8863 ( .A(n9309), .B(n9310), .Z(n8898) );
  NANDN U8864 ( .A(n8905), .B(n9311), .Z(n9309) );
  NANDN U8865 ( .A(n8904), .B(n8902), .Z(n9311) );
  XOR U8866 ( .A(n9312), .B(n9313), .Z(n8902) );
  XNOR U8867 ( .A(n9314), .B(n9315), .Z(n9313) );
  ANDN U8868 ( .B(\stack[1][4] ), .A(n5350), .Z(n8904) );
  AND U8869 ( .A(n9316), .B(n9317), .Z(n8905) );
  NANDN U8870 ( .A(n8909), .B(n8911), .Z(n9317) );
  NANDN U8871 ( .A(n8912), .B(n9318), .Z(n9316) );
  NANDN U8872 ( .A(n8911), .B(n8909), .Z(n9318) );
  XOR U8873 ( .A(n9319), .B(n9320), .Z(n8909) );
  XNOR U8874 ( .A(n9321), .B(n9322), .Z(n9320) );
  ANDN U8875 ( .B(\stack[0][7] ), .A(n5267), .Z(n8911) );
  AND U8876 ( .A(n9323), .B(n9324), .Z(n8912) );
  NANDN U8877 ( .A(n8919), .B(n9325), .Z(n9323) );
  NANDN U8878 ( .A(n8918), .B(n8916), .Z(n9325) );
  XOR U8879 ( .A(n9326), .B(n9327), .Z(n8916) );
  XNOR U8880 ( .A(n9328), .B(n9329), .Z(n9327) );
  ANDN U8881 ( .B(\stack[1][4] ), .A(n5302), .Z(n8918) );
  AND U8882 ( .A(n9330), .B(n9331), .Z(n8919) );
  NANDN U8883 ( .A(n8925), .B(n8923), .Z(n9331) );
  IV U8884 ( .A(n9332), .Z(n8925) );
  NANDN U8885 ( .A(n8926), .B(n9333), .Z(n9330) );
  OR U8886 ( .A(n8923), .B(n9332), .Z(n9333) );
  ANDN U8887 ( .B(\stack[0][5] ), .A(n5267), .Z(n9332) );
  XNOR U8888 ( .A(n9334), .B(n9335), .Z(n8923) );
  XNOR U8889 ( .A(n9336), .B(n9337), .Z(n9335) );
  AND U8890 ( .A(n9338), .B(n9339), .Z(n8926) );
  NANDN U8891 ( .A(n8933), .B(n9340), .Z(n9338) );
  NANDN U8892 ( .A(n8932), .B(n8930), .Z(n9340) );
  XOR U8893 ( .A(n9341), .B(n9342), .Z(n8930) );
  XNOR U8894 ( .A(n9343), .B(n9344), .Z(n9342) );
  ANDN U8895 ( .B(\stack[0][4] ), .A(n5267), .Z(n8932) );
  AND U8896 ( .A(n9345), .B(n9346), .Z(n8933) );
  NANDN U8897 ( .A(n8937), .B(n8939), .Z(n9346) );
  NANDN U8898 ( .A(n8940), .B(n9347), .Z(n9345) );
  NANDN U8899 ( .A(n8939), .B(n8937), .Z(n9347) );
  XNOR U8900 ( .A(n9348), .B(n9349), .Z(n8937) );
  XNOR U8901 ( .A(n9350), .B(n9351), .Z(n9349) );
  ANDN U8902 ( .B(\stack[1][4] ), .A(n5230), .Z(n8939) );
  AND U8903 ( .A(n9352), .B(n9353), .Z(n8940) );
  NANDN U8904 ( .A(n8944), .B(n8946), .Z(n9353) );
  NAND U8905 ( .A(n9354), .B(n8947), .Z(n9352) );
  ANDN U8906 ( .B(n9355), .A(n8952), .Z(n8947) );
  NANDN U8907 ( .A(n5267), .B(\stack[0][1] ), .Z(n8952) );
  ANDN U8908 ( .B(\stack[0][0] ), .A(n5292), .Z(n9355) );
  NANDN U8909 ( .A(n8946), .B(n8944), .Z(n9354) );
  XNOR U8910 ( .A(n9356), .B(n9357), .Z(n8944) );
  NANDN U8911 ( .A(n5160), .B(\stack[1][6] ), .Z(n9357) );
  ANDN U8912 ( .B(\stack[1][4] ), .A(n5206), .Z(n8946) );
  ANDN U8913 ( .B(\stack[1][4] ), .A(n6574), .Z(n8956) );
  XOR U8914 ( .A(n9358), .B(n9359), .Z(n8954) );
  AND U8915 ( .A(n9360), .B(n9361), .Z(n9359) );
  NANDN U8916 ( .A(n8961), .B(n8963), .Z(n9361) );
  NANDN U8917 ( .A(n8964), .B(n9362), .Z(n9360) );
  NANDN U8918 ( .A(n8963), .B(n8961), .Z(n9362) );
  XOR U8919 ( .A(n7147), .B(n9363), .Z(n8961) );
  XNOR U8920 ( .A(n7148), .B(n7149), .Z(n9363) );
  AND U8921 ( .A(n9364), .B(n9365), .Z(n7149) );
  NAND U8922 ( .A(n9366), .B(n9367), .Z(n9365) );
  NANDN U8923 ( .A(n9368), .B(n9369), .Z(n9364) );
  OR U8924 ( .A(n9366), .B(n9367), .Z(n9369) );
  AND U8925 ( .A(\stack[1][6] ), .B(\stack[0][56] ), .Z(n7148) );
  IV U8926 ( .A(n7151), .Z(n7147) );
  XOR U8927 ( .A(n7697), .B(n9370), .Z(n7151) );
  XOR U8928 ( .A(n7696), .B(n7698), .Z(n9370) );
  AND U8929 ( .A(n9371), .B(n9372), .Z(n7698) );
  NANDN U8930 ( .A(n9373), .B(n9374), .Z(n9372) );
  NANDN U8931 ( .A(n9375), .B(n9376), .Z(n9371) );
  NANDN U8932 ( .A(n9374), .B(n9373), .Z(n9376) );
  IV U8933 ( .A(n7700), .Z(n7696) );
  ANDN U8934 ( .B(\stack[1][7] ), .A(n6478), .Z(n7700) );
  XNOR U8935 ( .A(n7707), .B(n9377), .Z(n7697) );
  XNOR U8936 ( .A(n7708), .B(n7709), .Z(n9377) );
  AND U8937 ( .A(n9378), .B(n9379), .Z(n7709) );
  NAND U8938 ( .A(n9380), .B(n9381), .Z(n9379) );
  NANDN U8939 ( .A(n9382), .B(n9383), .Z(n9378) );
  OR U8940 ( .A(n9380), .B(n9381), .Z(n9383) );
  AND U8941 ( .A(\stack[1][8] ), .B(\stack[0][54] ), .Z(n7708) );
  XNOR U8942 ( .A(n7716), .B(n9384), .Z(n7707) );
  XOR U8943 ( .A(n7715), .B(n7717), .Z(n9384) );
  AND U8944 ( .A(n9385), .B(n9386), .Z(n7717) );
  NANDN U8945 ( .A(n9387), .B(n9388), .Z(n9386) );
  NANDN U8946 ( .A(n9389), .B(n9390), .Z(n9385) );
  NANDN U8947 ( .A(n9388), .B(n9387), .Z(n9390) );
  IV U8948 ( .A(n7719), .Z(n7715) );
  ANDN U8949 ( .B(\stack[1][9] ), .A(n6430), .Z(n7719) );
  XNOR U8950 ( .A(n7162), .B(n9391), .Z(n7716) );
  XNOR U8951 ( .A(n7163), .B(n7164), .Z(n9391) );
  AND U8952 ( .A(n9392), .B(n9393), .Z(n7164) );
  NAND U8953 ( .A(n9394), .B(n9395), .Z(n9393) );
  NANDN U8954 ( .A(n9396), .B(n9397), .Z(n9392) );
  OR U8955 ( .A(n9394), .B(n9395), .Z(n9397) );
  AND U8956 ( .A(\stack[0][52] ), .B(\stack[1][10] ), .Z(n7163) );
  XNOR U8957 ( .A(n7669), .B(n9398), .Z(n7162) );
  XOR U8958 ( .A(n7668), .B(n7670), .Z(n9398) );
  AND U8959 ( .A(n9399), .B(n9400), .Z(n7670) );
  NANDN U8960 ( .A(n9401), .B(n9402), .Z(n9400) );
  NANDN U8961 ( .A(n9403), .B(n9404), .Z(n9399) );
  NANDN U8962 ( .A(n9402), .B(n9401), .Z(n9404) );
  IV U8963 ( .A(n7672), .Z(n7668) );
  ANDN U8964 ( .B(\stack[0][51] ), .A(n5435), .Z(n7672) );
  XNOR U8965 ( .A(n7679), .B(n9405), .Z(n7669) );
  XNOR U8966 ( .A(n7680), .B(n7681), .Z(n9405) );
  AND U8967 ( .A(n9406), .B(n9407), .Z(n7681) );
  NAND U8968 ( .A(n9408), .B(n9409), .Z(n9407) );
  NANDN U8969 ( .A(n9410), .B(n9411), .Z(n9406) );
  OR U8970 ( .A(n9408), .B(n9409), .Z(n9411) );
  AND U8971 ( .A(\stack[0][50] ), .B(\stack[1][12] ), .Z(n7680) );
  XNOR U8972 ( .A(n7688), .B(n9412), .Z(n7679) );
  XOR U8973 ( .A(n7687), .B(n7689), .Z(n9412) );
  AND U8974 ( .A(n9413), .B(n9414), .Z(n7689) );
  NANDN U8975 ( .A(n9415), .B(n9416), .Z(n9414) );
  NANDN U8976 ( .A(n9417), .B(n9418), .Z(n9413) );
  NANDN U8977 ( .A(n9416), .B(n9415), .Z(n9418) );
  IV U8978 ( .A(n7691), .Z(n7687) );
  ANDN U8979 ( .B(\stack[0][49] ), .A(n5483), .Z(n7691) );
  XNOR U8980 ( .A(n7176), .B(n9419), .Z(n7688) );
  XNOR U8981 ( .A(n7177), .B(n7178), .Z(n9419) );
  AND U8982 ( .A(n9420), .B(n9421), .Z(n7178) );
  NAND U8983 ( .A(n9422), .B(n9423), .Z(n9421) );
  NANDN U8984 ( .A(n9424), .B(n9425), .Z(n9420) );
  OR U8985 ( .A(n9422), .B(n9423), .Z(n9425) );
  AND U8986 ( .A(\stack[0][48] ), .B(\stack[1][14] ), .Z(n7177) );
  XNOR U8987 ( .A(n7641), .B(n9426), .Z(n7176) );
  XOR U8988 ( .A(n7640), .B(n7642), .Z(n9426) );
  AND U8989 ( .A(n9427), .B(n9428), .Z(n7642) );
  NANDN U8990 ( .A(n9429), .B(n9430), .Z(n9428) );
  NANDN U8991 ( .A(n9431), .B(n9432), .Z(n9427) );
  NANDN U8992 ( .A(n9430), .B(n9429), .Z(n9432) );
  IV U8993 ( .A(n7644), .Z(n7640) );
  ANDN U8994 ( .B(\stack[0][47] ), .A(n5531), .Z(n7644) );
  XNOR U8995 ( .A(n7651), .B(n9433), .Z(n7641) );
  XNOR U8996 ( .A(n7652), .B(n7653), .Z(n9433) );
  AND U8997 ( .A(n9434), .B(n9435), .Z(n7653) );
  NAND U8998 ( .A(n9436), .B(n9437), .Z(n9435) );
  NANDN U8999 ( .A(n9438), .B(n9439), .Z(n9434) );
  OR U9000 ( .A(n9436), .B(n9437), .Z(n9439) );
  AND U9001 ( .A(\stack[0][46] ), .B(\stack[1][16] ), .Z(n7652) );
  XNOR U9002 ( .A(n7660), .B(n9440), .Z(n7651) );
  XOR U9003 ( .A(n7659), .B(n7661), .Z(n9440) );
  AND U9004 ( .A(n9441), .B(n9442), .Z(n7661) );
  NANDN U9005 ( .A(n9443), .B(n9444), .Z(n9442) );
  NANDN U9006 ( .A(n9445), .B(n9446), .Z(n9441) );
  NANDN U9007 ( .A(n9444), .B(n9443), .Z(n9446) );
  IV U9008 ( .A(n7663), .Z(n7659) );
  ANDN U9009 ( .B(\stack[0][45] ), .A(n5579), .Z(n7663) );
  XNOR U9010 ( .A(n7190), .B(n9447), .Z(n7660) );
  XNOR U9011 ( .A(n7191), .B(n7192), .Z(n9447) );
  AND U9012 ( .A(n9448), .B(n9449), .Z(n7192) );
  NAND U9013 ( .A(n9450), .B(n9451), .Z(n9449) );
  NANDN U9014 ( .A(n9452), .B(n9453), .Z(n9448) );
  OR U9015 ( .A(n9450), .B(n9451), .Z(n9453) );
  AND U9016 ( .A(\stack[0][44] ), .B(\stack[1][18] ), .Z(n7191) );
  XNOR U9017 ( .A(n7613), .B(n9454), .Z(n7190) );
  XOR U9018 ( .A(n7612), .B(n7614), .Z(n9454) );
  AND U9019 ( .A(n9455), .B(n9456), .Z(n7614) );
  NANDN U9020 ( .A(n9457), .B(n9458), .Z(n9456) );
  NANDN U9021 ( .A(n9459), .B(n9460), .Z(n9455) );
  NANDN U9022 ( .A(n9458), .B(n9457), .Z(n9460) );
  IV U9023 ( .A(n7616), .Z(n7612) );
  ANDN U9024 ( .B(\stack[0][43] ), .A(n5627), .Z(n7616) );
  XNOR U9025 ( .A(n7623), .B(n9461), .Z(n7613) );
  XNOR U9026 ( .A(n7624), .B(n7625), .Z(n9461) );
  AND U9027 ( .A(n9462), .B(n9463), .Z(n7625) );
  NAND U9028 ( .A(n9464), .B(n9465), .Z(n9463) );
  NANDN U9029 ( .A(n9466), .B(n9467), .Z(n9462) );
  OR U9030 ( .A(n9464), .B(n9465), .Z(n9467) );
  AND U9031 ( .A(\stack[0][42] ), .B(\stack[1][20] ), .Z(n7624) );
  XNOR U9032 ( .A(n7632), .B(n9468), .Z(n7623) );
  XOR U9033 ( .A(n7631), .B(n7633), .Z(n9468) );
  AND U9034 ( .A(n9469), .B(n9470), .Z(n7633) );
  NANDN U9035 ( .A(n9471), .B(n9472), .Z(n9470) );
  NANDN U9036 ( .A(n9473), .B(n9474), .Z(n9469) );
  NANDN U9037 ( .A(n9472), .B(n9471), .Z(n9474) );
  IV U9038 ( .A(n7635), .Z(n7631) );
  ANDN U9039 ( .B(\stack[0][41] ), .A(n5675), .Z(n7635) );
  XNOR U9040 ( .A(n7204), .B(n9475), .Z(n7632) );
  XNOR U9041 ( .A(n7205), .B(n7206), .Z(n9475) );
  AND U9042 ( .A(n9476), .B(n9477), .Z(n7206) );
  NAND U9043 ( .A(n9478), .B(n9479), .Z(n9477) );
  NANDN U9044 ( .A(n9480), .B(n9481), .Z(n9476) );
  OR U9045 ( .A(n9478), .B(n9479), .Z(n9481) );
  AND U9046 ( .A(\stack[0][40] ), .B(\stack[1][22] ), .Z(n7205) );
  XNOR U9047 ( .A(n7585), .B(n9482), .Z(n7204) );
  XOR U9048 ( .A(n7584), .B(n7586), .Z(n9482) );
  AND U9049 ( .A(n9483), .B(n9484), .Z(n7586) );
  NANDN U9050 ( .A(n9485), .B(n9486), .Z(n9484) );
  NANDN U9051 ( .A(n9487), .B(n9488), .Z(n9483) );
  NANDN U9052 ( .A(n9486), .B(n9485), .Z(n9488) );
  IV U9053 ( .A(n7588), .Z(n7584) );
  ANDN U9054 ( .B(\stack[0][39] ), .A(n5723), .Z(n7588) );
  XNOR U9055 ( .A(n7595), .B(n9489), .Z(n7585) );
  XNOR U9056 ( .A(n7596), .B(n7597), .Z(n9489) );
  AND U9057 ( .A(n9490), .B(n9491), .Z(n7597) );
  NAND U9058 ( .A(n9492), .B(n9493), .Z(n9491) );
  NANDN U9059 ( .A(n9494), .B(n9495), .Z(n9490) );
  OR U9060 ( .A(n9492), .B(n9493), .Z(n9495) );
  AND U9061 ( .A(\stack[0][38] ), .B(\stack[1][24] ), .Z(n7596) );
  XNOR U9062 ( .A(n7604), .B(n9496), .Z(n7595) );
  XOR U9063 ( .A(n7603), .B(n7605), .Z(n9496) );
  AND U9064 ( .A(n9497), .B(n9498), .Z(n7605) );
  NANDN U9065 ( .A(n9499), .B(n9500), .Z(n9498) );
  NANDN U9066 ( .A(n9501), .B(n9502), .Z(n9497) );
  NANDN U9067 ( .A(n9500), .B(n9499), .Z(n9502) );
  IV U9068 ( .A(n7607), .Z(n7603) );
  ANDN U9069 ( .B(\stack[0][37] ), .A(n5771), .Z(n7607) );
  XNOR U9070 ( .A(n7218), .B(n9503), .Z(n7604) );
  XNOR U9071 ( .A(n7219), .B(n7220), .Z(n9503) );
  AND U9072 ( .A(n9504), .B(n9505), .Z(n7220) );
  NAND U9073 ( .A(n9506), .B(n9507), .Z(n9505) );
  NANDN U9074 ( .A(n9508), .B(n9509), .Z(n9504) );
  OR U9075 ( .A(n9506), .B(n9507), .Z(n9509) );
  AND U9076 ( .A(\stack[0][36] ), .B(\stack[1][26] ), .Z(n7219) );
  XNOR U9077 ( .A(n7557), .B(n9510), .Z(n7218) );
  XOR U9078 ( .A(n7556), .B(n7558), .Z(n9510) );
  AND U9079 ( .A(n9511), .B(n9512), .Z(n7558) );
  NANDN U9080 ( .A(n9513), .B(n9514), .Z(n9512) );
  NANDN U9081 ( .A(n9515), .B(n9516), .Z(n9511) );
  NANDN U9082 ( .A(n9514), .B(n9513), .Z(n9516) );
  IV U9083 ( .A(n7560), .Z(n7556) );
  ANDN U9084 ( .B(\stack[0][35] ), .A(n5819), .Z(n7560) );
  XNOR U9085 ( .A(n7567), .B(n9517), .Z(n7557) );
  XNOR U9086 ( .A(n7568), .B(n7569), .Z(n9517) );
  AND U9087 ( .A(n9518), .B(n9519), .Z(n7569) );
  NAND U9088 ( .A(n9520), .B(n9521), .Z(n9519) );
  NANDN U9089 ( .A(n9522), .B(n9523), .Z(n9518) );
  OR U9090 ( .A(n9520), .B(n9521), .Z(n9523) );
  AND U9091 ( .A(\stack[0][34] ), .B(\stack[1][28] ), .Z(n7568) );
  XNOR U9092 ( .A(n7576), .B(n9524), .Z(n7567) );
  XOR U9093 ( .A(n7575), .B(n7577), .Z(n9524) );
  AND U9094 ( .A(n9525), .B(n9526), .Z(n7577) );
  NANDN U9095 ( .A(n9527), .B(n9528), .Z(n9526) );
  NANDN U9096 ( .A(n9529), .B(n9530), .Z(n9525) );
  NANDN U9097 ( .A(n9528), .B(n9527), .Z(n9530) );
  IV U9098 ( .A(n7579), .Z(n7575) );
  ANDN U9099 ( .B(\stack[0][33] ), .A(n5867), .Z(n7579) );
  XNOR U9100 ( .A(n7232), .B(n9531), .Z(n7576) );
  XNOR U9101 ( .A(n7233), .B(n7234), .Z(n9531) );
  AND U9102 ( .A(n9532), .B(n9533), .Z(n7234) );
  NAND U9103 ( .A(n9534), .B(n9535), .Z(n9533) );
  NANDN U9104 ( .A(n9536), .B(n9537), .Z(n9532) );
  OR U9105 ( .A(n9534), .B(n9535), .Z(n9537) );
  AND U9106 ( .A(\stack[0][32] ), .B(\stack[1][30] ), .Z(n7233) );
  XNOR U9107 ( .A(n7529), .B(n9538), .Z(n7232) );
  XOR U9108 ( .A(n7528), .B(n7530), .Z(n9538) );
  AND U9109 ( .A(n9539), .B(n9540), .Z(n7530) );
  NANDN U9110 ( .A(n9541), .B(n9542), .Z(n9540) );
  NANDN U9111 ( .A(n9543), .B(n9544), .Z(n9539) );
  NANDN U9112 ( .A(n9542), .B(n9541), .Z(n9544) );
  IV U9113 ( .A(n7532), .Z(n7528) );
  ANDN U9114 ( .B(\stack[0][31] ), .A(n5915), .Z(n7532) );
  XNOR U9115 ( .A(n7539), .B(n9545), .Z(n7529) );
  XNOR U9116 ( .A(n7540), .B(n7541), .Z(n9545) );
  AND U9117 ( .A(n9546), .B(n9547), .Z(n7541) );
  NAND U9118 ( .A(n9548), .B(n9549), .Z(n9547) );
  NANDN U9119 ( .A(n9550), .B(n9551), .Z(n9546) );
  OR U9120 ( .A(n9548), .B(n9549), .Z(n9551) );
  AND U9121 ( .A(\stack[0][30] ), .B(\stack[1][32] ), .Z(n7540) );
  XNOR U9122 ( .A(n7548), .B(n9552), .Z(n7539) );
  XOR U9123 ( .A(n7547), .B(n7549), .Z(n9552) );
  AND U9124 ( .A(n9553), .B(n9554), .Z(n7549) );
  NANDN U9125 ( .A(n9555), .B(n9556), .Z(n9554) );
  NANDN U9126 ( .A(n9557), .B(n9558), .Z(n9553) );
  NANDN U9127 ( .A(n9556), .B(n9555), .Z(n9558) );
  IV U9128 ( .A(n7551), .Z(n7547) );
  ANDN U9129 ( .B(\stack[0][29] ), .A(n5964), .Z(n7551) );
  XNOR U9130 ( .A(n7244), .B(n9559), .Z(n7548) );
  XNOR U9131 ( .A(n7245), .B(n7246), .Z(n9559) );
  AND U9132 ( .A(n9560), .B(n9561), .Z(n7246) );
  NAND U9133 ( .A(n9562), .B(n9563), .Z(n9561) );
  NANDN U9134 ( .A(n9564), .B(n9565), .Z(n9560) );
  OR U9135 ( .A(n9562), .B(n9563), .Z(n9565) );
  AND U9136 ( .A(\stack[0][28] ), .B(\stack[1][34] ), .Z(n7245) );
  XNOR U9137 ( .A(n7508), .B(n9566), .Z(n7244) );
  XOR U9138 ( .A(n7507), .B(n7509), .Z(n9566) );
  AND U9139 ( .A(n9567), .B(n9568), .Z(n7509) );
  NANDN U9140 ( .A(n9569), .B(n9570), .Z(n9568) );
  NANDN U9141 ( .A(n9571), .B(n9572), .Z(n9567) );
  NANDN U9142 ( .A(n9570), .B(n9569), .Z(n9572) );
  IV U9143 ( .A(n7511), .Z(n7507) );
  ANDN U9144 ( .B(\stack[0][27] ), .A(n6012), .Z(n7511) );
  XNOR U9145 ( .A(n7518), .B(n9573), .Z(n7508) );
  XNOR U9146 ( .A(n7519), .B(n7520), .Z(n9573) );
  AND U9147 ( .A(n9574), .B(n9575), .Z(n7520) );
  NAND U9148 ( .A(n9576), .B(n9577), .Z(n9575) );
  NANDN U9149 ( .A(n9578), .B(n9579), .Z(n9574) );
  OR U9150 ( .A(n9576), .B(n9577), .Z(n9579) );
  AND U9151 ( .A(\stack[0][26] ), .B(\stack[1][36] ), .Z(n7519) );
  XOR U9152 ( .A(n7503), .B(n7504), .Z(n9580) );
  NAND U9153 ( .A(n9581), .B(n9582), .Z(n7504) );
  NANDN U9154 ( .A(n9583), .B(n9584), .Z(n9582) );
  OR U9155 ( .A(n9585), .B(n9586), .Z(n9584) );
  AND U9156 ( .A(\stack[0][25] ), .B(\stack[1][37] ), .Z(n7503) );
  XOR U9157 ( .A(n7256), .B(n9587), .Z(n7501) );
  XOR U9158 ( .A(n7258), .B(n7261), .Z(n9587) );
  IV U9159 ( .A(n7257), .Z(n7261) );
  NAND U9160 ( .A(n9588), .B(n9589), .Z(n7257) );
  NAND U9161 ( .A(n9590), .B(n9591), .Z(n9589) );
  OR U9162 ( .A(n9592), .B(n9593), .Z(n9590) );
  NANDN U9163 ( .A(n6084), .B(\stack[0][24] ), .Z(n7258) );
  IV U9164 ( .A(n7260), .Z(n7256) );
  XOR U9165 ( .A(n7485), .B(n9594), .Z(n7260) );
  XOR U9166 ( .A(n7484), .B(n7486), .Z(n9594) );
  AND U9167 ( .A(n9595), .B(n9596), .Z(n7486) );
  NANDN U9168 ( .A(n9597), .B(n9598), .Z(n9596) );
  NANDN U9169 ( .A(n9599), .B(n9600), .Z(n9595) );
  NANDN U9170 ( .A(n9598), .B(n9597), .Z(n9600) );
  IV U9171 ( .A(n7488), .Z(n7484) );
  ANDN U9172 ( .B(\stack[0][23] ), .A(n6108), .Z(n7488) );
  XNOR U9173 ( .A(n7493), .B(n9601), .Z(n7485) );
  XNOR U9174 ( .A(n7494), .B(n7495), .Z(n9601) );
  AND U9175 ( .A(n9602), .B(n9603), .Z(n7495) );
  NAND U9176 ( .A(n9604), .B(n9605), .Z(n9603) );
  NANDN U9177 ( .A(n9606), .B(n9607), .Z(n9602) );
  OR U9178 ( .A(n9604), .B(n9605), .Z(n9607) );
  AND U9179 ( .A(\stack[0][22] ), .B(\stack[1][40] ), .Z(n7494) );
  XNOR U9180 ( .A(n7271), .B(n9608), .Z(n7493) );
  XOR U9181 ( .A(n7270), .B(n7272), .Z(n9608) );
  AND U9182 ( .A(n9609), .B(n9610), .Z(n7272) );
  NANDN U9183 ( .A(n9611), .B(n9612), .Z(n9610) );
  NANDN U9184 ( .A(n9613), .B(n9614), .Z(n9609) );
  NANDN U9185 ( .A(n9612), .B(n9611), .Z(n9614) );
  IV U9186 ( .A(n7274), .Z(n7270) );
  ANDN U9187 ( .B(\stack[0][21] ), .A(n6156), .Z(n7274) );
  XNOR U9188 ( .A(n7465), .B(n9615), .Z(n7271) );
  XNOR U9189 ( .A(n7466), .B(n7467), .Z(n9615) );
  AND U9190 ( .A(n9616), .B(n9617), .Z(n7467) );
  NAND U9191 ( .A(n9618), .B(n9619), .Z(n9617) );
  NANDN U9192 ( .A(n9620), .B(n9621), .Z(n9616) );
  OR U9193 ( .A(n9618), .B(n9619), .Z(n9621) );
  AND U9194 ( .A(\stack[0][20] ), .B(\stack[1][42] ), .Z(n7466) );
  XNOR U9195 ( .A(n7474), .B(n9622), .Z(n7465) );
  XOR U9196 ( .A(n7473), .B(n7475), .Z(n9622) );
  AND U9197 ( .A(n9623), .B(n9624), .Z(n7475) );
  NANDN U9198 ( .A(n9625), .B(n9626), .Z(n9624) );
  NANDN U9199 ( .A(n9627), .B(n9628), .Z(n9623) );
  NANDN U9200 ( .A(n9626), .B(n9625), .Z(n9628) );
  IV U9201 ( .A(n7477), .Z(n7473) );
  ANDN U9202 ( .B(\stack[0][19] ), .A(n6204), .Z(n7477) );
  XNOR U9203 ( .A(n7283), .B(n9629), .Z(n7474) );
  XNOR U9204 ( .A(n7284), .B(n7285), .Z(n9629) );
  AND U9205 ( .A(n9630), .B(n9631), .Z(n7285) );
  NAND U9206 ( .A(n9632), .B(n9633), .Z(n9631) );
  NANDN U9207 ( .A(n9634), .B(n9635), .Z(n9630) );
  OR U9208 ( .A(n9632), .B(n9633), .Z(n9635) );
  AND U9209 ( .A(\stack[0][18] ), .B(\stack[1][44] ), .Z(n7284) );
  XNOR U9210 ( .A(n7447), .B(n9636), .Z(n7283) );
  XOR U9211 ( .A(n7446), .B(n7448), .Z(n9636) );
  AND U9212 ( .A(n9637), .B(n9638), .Z(n7448) );
  NANDN U9213 ( .A(n9639), .B(n9640), .Z(n9638) );
  NANDN U9214 ( .A(n9641), .B(n9642), .Z(n9637) );
  NANDN U9215 ( .A(n9640), .B(n9639), .Z(n9642) );
  IV U9216 ( .A(n7450), .Z(n7446) );
  ANDN U9217 ( .B(\stack[0][17] ), .A(n6252), .Z(n7450) );
  XNOR U9218 ( .A(n7455), .B(n9643), .Z(n7447) );
  XNOR U9219 ( .A(n7456), .B(n7457), .Z(n9643) );
  AND U9220 ( .A(n9644), .B(n9645), .Z(n7457) );
  NAND U9221 ( .A(n9646), .B(n9647), .Z(n9645) );
  NANDN U9222 ( .A(n9648), .B(n9649), .Z(n9644) );
  OR U9223 ( .A(n9646), .B(n9647), .Z(n9649) );
  AND U9224 ( .A(\stack[0][16] ), .B(\stack[1][46] ), .Z(n7456) );
  XNOR U9225 ( .A(n7296), .B(n9650), .Z(n7455) );
  XOR U9226 ( .A(n7295), .B(n7297), .Z(n9650) );
  AND U9227 ( .A(n9651), .B(n9652), .Z(n7297) );
  NANDN U9228 ( .A(n9653), .B(n9654), .Z(n9652) );
  NANDN U9229 ( .A(n9655), .B(n9656), .Z(n9651) );
  NANDN U9230 ( .A(n9654), .B(n9653), .Z(n9656) );
  IV U9231 ( .A(n7299), .Z(n7295) );
  ANDN U9232 ( .B(\stack[0][15] ), .A(n6300), .Z(n7299) );
  XNOR U9233 ( .A(n7427), .B(n9657), .Z(n7296) );
  XNOR U9234 ( .A(n7428), .B(n7429), .Z(n9657) );
  AND U9235 ( .A(n9658), .B(n9659), .Z(n7429) );
  NAND U9236 ( .A(n9660), .B(n9661), .Z(n9659) );
  NANDN U9237 ( .A(n9662), .B(n9663), .Z(n9658) );
  OR U9238 ( .A(n9660), .B(n9661), .Z(n9663) );
  AND U9239 ( .A(\stack[0][14] ), .B(\stack[1][48] ), .Z(n7428) );
  XNOR U9240 ( .A(n7436), .B(n9664), .Z(n7427) );
  XOR U9241 ( .A(n7435), .B(n7437), .Z(n9664) );
  AND U9242 ( .A(n9665), .B(n9666), .Z(n7437) );
  NANDN U9243 ( .A(n9667), .B(n9668), .Z(n9666) );
  NANDN U9244 ( .A(n9669), .B(n9670), .Z(n9665) );
  NANDN U9245 ( .A(n9668), .B(n9667), .Z(n9670) );
  IV U9246 ( .A(n7439), .Z(n7435) );
  ANDN U9247 ( .B(\stack[0][13] ), .A(n6348), .Z(n7439) );
  XNOR U9248 ( .A(n7308), .B(n9671), .Z(n7436) );
  XNOR U9249 ( .A(n7309), .B(n7310), .Z(n9671) );
  AND U9250 ( .A(n9672), .B(n9673), .Z(n7310) );
  NAND U9251 ( .A(n9674), .B(n9675), .Z(n9673) );
  NANDN U9252 ( .A(n9676), .B(n9677), .Z(n9672) );
  OR U9253 ( .A(n9674), .B(n9675), .Z(n9677) );
  AND U9254 ( .A(\stack[0][12] ), .B(\stack[1][50] ), .Z(n7309) );
  XNOR U9255 ( .A(n7409), .B(n9678), .Z(n7308) );
  XOR U9256 ( .A(n7408), .B(n7410), .Z(n9678) );
  AND U9257 ( .A(n9679), .B(n9680), .Z(n7410) );
  NANDN U9258 ( .A(n9681), .B(n9682), .Z(n9680) );
  NANDN U9259 ( .A(n9683), .B(n9684), .Z(n9679) );
  NANDN U9260 ( .A(n9682), .B(n9681), .Z(n9684) );
  IV U9261 ( .A(n7412), .Z(n7408) );
  ANDN U9262 ( .B(\stack[0][11] ), .A(n6396), .Z(n7412) );
  XNOR U9263 ( .A(n7417), .B(n9685), .Z(n7409) );
  XNOR U9264 ( .A(n7418), .B(n7419), .Z(n9685) );
  AND U9265 ( .A(n9686), .B(n9687), .Z(n7419) );
  NAND U9266 ( .A(n9688), .B(n9689), .Z(n9687) );
  NANDN U9267 ( .A(n9690), .B(n9691), .Z(n9686) );
  OR U9268 ( .A(n9688), .B(n9689), .Z(n9691) );
  AND U9269 ( .A(\stack[0][10] ), .B(\stack[1][52] ), .Z(n7418) );
  XNOR U9270 ( .A(n7321), .B(n9692), .Z(n7417) );
  XOR U9271 ( .A(n7320), .B(n7322), .Z(n9692) );
  AND U9272 ( .A(n9693), .B(n9694), .Z(n7322) );
  NANDN U9273 ( .A(n9695), .B(n9696), .Z(n9694) );
  NANDN U9274 ( .A(n9697), .B(n9698), .Z(n9693) );
  NANDN U9275 ( .A(n9696), .B(n9695), .Z(n9698) );
  IV U9276 ( .A(n7324), .Z(n7320) );
  ANDN U9277 ( .B(\stack[0][9] ), .A(n6444), .Z(n7324) );
  XNOR U9278 ( .A(n7389), .B(n9699), .Z(n7321) );
  XNOR U9279 ( .A(n7390), .B(n7391), .Z(n9699) );
  AND U9280 ( .A(n9700), .B(n9701), .Z(n7391) );
  NAND U9281 ( .A(n9702), .B(n9703), .Z(n9701) );
  NANDN U9282 ( .A(n9704), .B(n9705), .Z(n9700) );
  OR U9283 ( .A(n9702), .B(n9703), .Z(n9705) );
  AND U9284 ( .A(\stack[0][8] ), .B(\stack[1][54] ), .Z(n7390) );
  XNOR U9285 ( .A(n7398), .B(n9706), .Z(n7389) );
  XOR U9286 ( .A(n7397), .B(n7399), .Z(n9706) );
  AND U9287 ( .A(n9707), .B(n9708), .Z(n7399) );
  NANDN U9288 ( .A(n9709), .B(n9710), .Z(n9708) );
  NANDN U9289 ( .A(n9711), .B(n9712), .Z(n9707) );
  NANDN U9290 ( .A(n9710), .B(n9709), .Z(n9712) );
  IV U9291 ( .A(n7401), .Z(n7397) );
  ANDN U9292 ( .B(\stack[0][7] ), .A(n6492), .Z(n7401) );
  XNOR U9293 ( .A(n7339), .B(n9713), .Z(n7398) );
  XNOR U9294 ( .A(n7340), .B(n7341), .Z(n9713) );
  AND U9295 ( .A(n9714), .B(n9715), .Z(n7341) );
  NAND U9296 ( .A(n9716), .B(n9717), .Z(n9715) );
  NANDN U9297 ( .A(n9718), .B(n9719), .Z(n9714) );
  OR U9298 ( .A(n9716), .B(n9717), .Z(n9719) );
  AND U9299 ( .A(\stack[0][6] ), .B(\stack[1][56] ), .Z(n7340) );
  XNOR U9300 ( .A(n7371), .B(n9720), .Z(n7339) );
  XOR U9301 ( .A(n7370), .B(n7372), .Z(n9720) );
  AND U9302 ( .A(n9721), .B(n9722), .Z(n7372) );
  NANDN U9303 ( .A(n9723), .B(n9724), .Z(n9722) );
  NANDN U9304 ( .A(n9725), .B(n9726), .Z(n9721) );
  NANDN U9305 ( .A(n9724), .B(n9723), .Z(n9726) );
  IV U9306 ( .A(n7374), .Z(n7370) );
  ANDN U9307 ( .B(\stack[0][5] ), .A(n6540), .Z(n7374) );
  XNOR U9308 ( .A(n7379), .B(n9727), .Z(n7371) );
  XNOR U9309 ( .A(n7380), .B(n7381), .Z(n9727) );
  AND U9310 ( .A(n9728), .B(n9729), .Z(n7381) );
  NAND U9311 ( .A(n9730), .B(n9731), .Z(n9729) );
  NANDN U9312 ( .A(n9732), .B(n9733), .Z(n9728) );
  OR U9313 ( .A(n9730), .B(n9731), .Z(n9733) );
  AND U9314 ( .A(\stack[0][4] ), .B(\stack[1][58] ), .Z(n7380) );
  XNOR U9315 ( .A(n7348), .B(n9734), .Z(n7379) );
  XOR U9316 ( .A(n7347), .B(n7349), .Z(n9734) );
  AND U9317 ( .A(n9735), .B(n9736), .Z(n7349) );
  NAND U9318 ( .A(n9737), .B(n9738), .Z(n9736) );
  NAND U9319 ( .A(n9739), .B(n9740), .Z(n9735) );
  OR U9320 ( .A(n9737), .B(n9738), .Z(n9739) );
  IV U9321 ( .A(n7351), .Z(n7347) );
  ANDN U9322 ( .B(\stack[0][3] ), .A(n6588), .Z(n7351) );
  XNOR U9323 ( .A(n7358), .B(n9741), .Z(n7348) );
  XOR U9324 ( .A(n7360), .B(n7359), .Z(n9741) );
  ANDN U9325 ( .B(\stack[1][60] ), .A(n5206), .Z(n7359) );
  NANDN U9326 ( .A(n9742), .B(n9743), .Z(n7360) );
  ANDN U9327 ( .B(\stack[0][0] ), .A(n6636), .Z(n9743) );
  XOR U9328 ( .A(n7334), .B(n9744), .Z(n7358) );
  NANDN U9329 ( .A(n5160), .B(\stack[1][62] ), .Z(n9744) );
  NANDN U9330 ( .A(n6636), .B(\stack[0][1] ), .Z(n7334) );
  ANDN U9331 ( .B(\stack[0][57] ), .A(n5292), .Z(n8963) );
  AND U9332 ( .A(n9745), .B(n9746), .Z(n8964) );
  NANDN U9333 ( .A(n8971), .B(n9747), .Z(n9745) );
  NANDN U9334 ( .A(n8970), .B(n8968), .Z(n9747) );
  XNOR U9335 ( .A(n9366), .B(n9748), .Z(n8968) );
  XNOR U9336 ( .A(n9367), .B(n9368), .Z(n9748) );
  AND U9337 ( .A(n9749), .B(n9750), .Z(n9368) );
  NANDN U9338 ( .A(n9751), .B(n9752), .Z(n9750) );
  NANDN U9339 ( .A(n9753), .B(n9754), .Z(n9749) );
  NANDN U9340 ( .A(n9752), .B(n9751), .Z(n9754) );
  ANDN U9341 ( .B(\stack[0][55] ), .A(n5316), .Z(n9367) );
  XNOR U9342 ( .A(n9373), .B(n9755), .Z(n9366) );
  XNOR U9343 ( .A(n9374), .B(n9375), .Z(n9755) );
  AND U9344 ( .A(n9756), .B(n9757), .Z(n9375) );
  NAND U9345 ( .A(n9758), .B(n9759), .Z(n9757) );
  NANDN U9346 ( .A(n9760), .B(n9761), .Z(n9756) );
  OR U9347 ( .A(n9758), .B(n9759), .Z(n9761) );
  ANDN U9348 ( .B(\stack[0][54] ), .A(n5340), .Z(n9374) );
  XNOR U9349 ( .A(n9380), .B(n9762), .Z(n9373) );
  XNOR U9350 ( .A(n9381), .B(n9382), .Z(n9762) );
  AND U9351 ( .A(n9763), .B(n9764), .Z(n9382) );
  NANDN U9352 ( .A(n9765), .B(n9766), .Z(n9764) );
  NANDN U9353 ( .A(n9767), .B(n9768), .Z(n9763) );
  NANDN U9354 ( .A(n9766), .B(n9765), .Z(n9768) );
  ANDN U9355 ( .B(\stack[0][53] ), .A(n5364), .Z(n9381) );
  XNOR U9356 ( .A(n9387), .B(n9769), .Z(n9380) );
  XNOR U9357 ( .A(n9388), .B(n9389), .Z(n9769) );
  AND U9358 ( .A(n9770), .B(n9771), .Z(n9389) );
  NAND U9359 ( .A(n9772), .B(n9773), .Z(n9771) );
  NANDN U9360 ( .A(n9774), .B(n9775), .Z(n9770) );
  OR U9361 ( .A(n9772), .B(n9773), .Z(n9775) );
  ANDN U9362 ( .B(\stack[0][52] ), .A(n5387), .Z(n9388) );
  XNOR U9363 ( .A(n9394), .B(n9776), .Z(n9387) );
  XNOR U9364 ( .A(n9395), .B(n9396), .Z(n9776) );
  AND U9365 ( .A(n9777), .B(n9778), .Z(n9396) );
  NANDN U9366 ( .A(n9779), .B(n9780), .Z(n9778) );
  NANDN U9367 ( .A(n9781), .B(n9782), .Z(n9777) );
  NANDN U9368 ( .A(n9780), .B(n9779), .Z(n9782) );
  ANDN U9369 ( .B(\stack[1][10] ), .A(n6382), .Z(n9395) );
  XNOR U9370 ( .A(n9401), .B(n9783), .Z(n9394) );
  XNOR U9371 ( .A(n9402), .B(n9403), .Z(n9783) );
  AND U9372 ( .A(n9784), .B(n9785), .Z(n9403) );
  NAND U9373 ( .A(n9786), .B(n9787), .Z(n9785) );
  NANDN U9374 ( .A(n9788), .B(n9789), .Z(n9784) );
  OR U9375 ( .A(n9786), .B(n9787), .Z(n9789) );
  ANDN U9376 ( .B(\stack[1][11] ), .A(n6358), .Z(n9402) );
  XNOR U9377 ( .A(n9408), .B(n9790), .Z(n9401) );
  XNOR U9378 ( .A(n9409), .B(n9410), .Z(n9790) );
  AND U9379 ( .A(n9791), .B(n9792), .Z(n9410) );
  NANDN U9380 ( .A(n9793), .B(n9794), .Z(n9792) );
  NANDN U9381 ( .A(n9795), .B(n9796), .Z(n9791) );
  NANDN U9382 ( .A(n9794), .B(n9793), .Z(n9796) );
  ANDN U9383 ( .B(\stack[1][12] ), .A(n6334), .Z(n9409) );
  XNOR U9384 ( .A(n9415), .B(n9797), .Z(n9408) );
  XNOR U9385 ( .A(n9416), .B(n9417), .Z(n9797) );
  AND U9386 ( .A(n9798), .B(n9799), .Z(n9417) );
  NAND U9387 ( .A(n9800), .B(n9801), .Z(n9799) );
  NANDN U9388 ( .A(n9802), .B(n9803), .Z(n9798) );
  OR U9389 ( .A(n9800), .B(n9801), .Z(n9803) );
  ANDN U9390 ( .B(\stack[1][13] ), .A(n6310), .Z(n9416) );
  XNOR U9391 ( .A(n9422), .B(n9804), .Z(n9415) );
  XNOR U9392 ( .A(n9423), .B(n9424), .Z(n9804) );
  AND U9393 ( .A(n9805), .B(n9806), .Z(n9424) );
  NANDN U9394 ( .A(n9807), .B(n9808), .Z(n9806) );
  NANDN U9395 ( .A(n9809), .B(n9810), .Z(n9805) );
  NANDN U9396 ( .A(n9808), .B(n9807), .Z(n9810) );
  ANDN U9397 ( .B(\stack[1][14] ), .A(n6286), .Z(n9423) );
  XNOR U9398 ( .A(n9429), .B(n9811), .Z(n9422) );
  XNOR U9399 ( .A(n9430), .B(n9431), .Z(n9811) );
  AND U9400 ( .A(n9812), .B(n9813), .Z(n9431) );
  NAND U9401 ( .A(n9814), .B(n9815), .Z(n9813) );
  NANDN U9402 ( .A(n9816), .B(n9817), .Z(n9812) );
  OR U9403 ( .A(n9814), .B(n9815), .Z(n9817) );
  ANDN U9404 ( .B(\stack[1][15] ), .A(n6262), .Z(n9430) );
  XNOR U9405 ( .A(n9436), .B(n9818), .Z(n9429) );
  XNOR U9406 ( .A(n9437), .B(n9438), .Z(n9818) );
  AND U9407 ( .A(n9819), .B(n9820), .Z(n9438) );
  NANDN U9408 ( .A(n9821), .B(n9822), .Z(n9820) );
  NANDN U9409 ( .A(n9823), .B(n9824), .Z(n9819) );
  NANDN U9410 ( .A(n9822), .B(n9821), .Z(n9824) );
  ANDN U9411 ( .B(\stack[1][16] ), .A(n6238), .Z(n9437) );
  XNOR U9412 ( .A(n9443), .B(n9825), .Z(n9436) );
  XNOR U9413 ( .A(n9444), .B(n9445), .Z(n9825) );
  AND U9414 ( .A(n9826), .B(n9827), .Z(n9445) );
  NAND U9415 ( .A(n9828), .B(n9829), .Z(n9827) );
  NANDN U9416 ( .A(n9830), .B(n9831), .Z(n9826) );
  OR U9417 ( .A(n9828), .B(n9829), .Z(n9831) );
  ANDN U9418 ( .B(\stack[1][17] ), .A(n6214), .Z(n9444) );
  XNOR U9419 ( .A(n9450), .B(n9832), .Z(n9443) );
  XNOR U9420 ( .A(n9451), .B(n9452), .Z(n9832) );
  AND U9421 ( .A(n9833), .B(n9834), .Z(n9452) );
  NANDN U9422 ( .A(n9835), .B(n9836), .Z(n9834) );
  NANDN U9423 ( .A(n9837), .B(n9838), .Z(n9833) );
  NANDN U9424 ( .A(n9836), .B(n9835), .Z(n9838) );
  ANDN U9425 ( .B(\stack[1][18] ), .A(n6190), .Z(n9451) );
  XNOR U9426 ( .A(n9457), .B(n9839), .Z(n9450) );
  XNOR U9427 ( .A(n9458), .B(n9459), .Z(n9839) );
  AND U9428 ( .A(n9840), .B(n9841), .Z(n9459) );
  NAND U9429 ( .A(n9842), .B(n9843), .Z(n9841) );
  NANDN U9430 ( .A(n9844), .B(n9845), .Z(n9840) );
  OR U9431 ( .A(n9842), .B(n9843), .Z(n9845) );
  ANDN U9432 ( .B(\stack[1][19] ), .A(n6166), .Z(n9458) );
  XNOR U9433 ( .A(n9464), .B(n9846), .Z(n9457) );
  XNOR U9434 ( .A(n9465), .B(n9466), .Z(n9846) );
  AND U9435 ( .A(n9847), .B(n9848), .Z(n9466) );
  NANDN U9436 ( .A(n9849), .B(n9850), .Z(n9848) );
  NANDN U9437 ( .A(n9851), .B(n9852), .Z(n9847) );
  NANDN U9438 ( .A(n9850), .B(n9849), .Z(n9852) );
  ANDN U9439 ( .B(\stack[1][20] ), .A(n6142), .Z(n9465) );
  XNOR U9440 ( .A(n9471), .B(n9853), .Z(n9464) );
  XNOR U9441 ( .A(n9472), .B(n9473), .Z(n9853) );
  AND U9442 ( .A(n9854), .B(n9855), .Z(n9473) );
  NAND U9443 ( .A(n9856), .B(n9857), .Z(n9855) );
  NANDN U9444 ( .A(n9858), .B(n9859), .Z(n9854) );
  OR U9445 ( .A(n9856), .B(n9857), .Z(n9859) );
  ANDN U9446 ( .B(\stack[1][21] ), .A(n6118), .Z(n9472) );
  XNOR U9447 ( .A(n9478), .B(n9860), .Z(n9471) );
  XNOR U9448 ( .A(n9479), .B(n9480), .Z(n9860) );
  AND U9449 ( .A(n9861), .B(n9862), .Z(n9480) );
  NANDN U9450 ( .A(n9863), .B(n9864), .Z(n9862) );
  NANDN U9451 ( .A(n9865), .B(n9866), .Z(n9861) );
  NANDN U9452 ( .A(n9864), .B(n9863), .Z(n9866) );
  ANDN U9453 ( .B(\stack[1][22] ), .A(n6094), .Z(n9479) );
  XNOR U9454 ( .A(n9485), .B(n9867), .Z(n9478) );
  XNOR U9455 ( .A(n9486), .B(n9487), .Z(n9867) );
  AND U9456 ( .A(n9868), .B(n9869), .Z(n9487) );
  NAND U9457 ( .A(n9870), .B(n9871), .Z(n9869) );
  NANDN U9458 ( .A(n9872), .B(n9873), .Z(n9868) );
  OR U9459 ( .A(n9870), .B(n9871), .Z(n9873) );
  ANDN U9460 ( .B(\stack[1][23] ), .A(n6070), .Z(n9486) );
  XNOR U9461 ( .A(n9492), .B(n9874), .Z(n9485) );
  XNOR U9462 ( .A(n9493), .B(n9494), .Z(n9874) );
  AND U9463 ( .A(n9875), .B(n9876), .Z(n9494) );
  NANDN U9464 ( .A(n9877), .B(n9878), .Z(n9876) );
  NANDN U9465 ( .A(n9879), .B(n9880), .Z(n9875) );
  NANDN U9466 ( .A(n9878), .B(n9877), .Z(n9880) );
  ANDN U9467 ( .B(\stack[1][24] ), .A(n6046), .Z(n9493) );
  XNOR U9468 ( .A(n9499), .B(n9881), .Z(n9492) );
  XNOR U9469 ( .A(n9500), .B(n9501), .Z(n9881) );
  AND U9470 ( .A(n9882), .B(n9883), .Z(n9501) );
  NAND U9471 ( .A(n9884), .B(n9885), .Z(n9883) );
  NANDN U9472 ( .A(n9886), .B(n9887), .Z(n9882) );
  OR U9473 ( .A(n9884), .B(n9885), .Z(n9887) );
  ANDN U9474 ( .B(\stack[1][25] ), .A(n6022), .Z(n9500) );
  XNOR U9475 ( .A(n9506), .B(n9888), .Z(n9499) );
  XNOR U9476 ( .A(n9507), .B(n9508), .Z(n9888) );
  AND U9477 ( .A(n9889), .B(n9890), .Z(n9508) );
  NANDN U9478 ( .A(n9891), .B(n9892), .Z(n9890) );
  NANDN U9479 ( .A(n9893), .B(n9894), .Z(n9889) );
  NANDN U9480 ( .A(n9892), .B(n9891), .Z(n9894) );
  ANDN U9481 ( .B(\stack[1][26] ), .A(n5998), .Z(n9507) );
  XNOR U9482 ( .A(n9513), .B(n9895), .Z(n9506) );
  XNOR U9483 ( .A(n9514), .B(n9515), .Z(n9895) );
  AND U9484 ( .A(n9896), .B(n9897), .Z(n9515) );
  NAND U9485 ( .A(n9898), .B(n9899), .Z(n9897) );
  NANDN U9486 ( .A(n9900), .B(n9901), .Z(n9896) );
  OR U9487 ( .A(n9898), .B(n9899), .Z(n9901) );
  ANDN U9488 ( .B(\stack[1][27] ), .A(n5974), .Z(n9514) );
  XNOR U9489 ( .A(n9520), .B(n9902), .Z(n9513) );
  XNOR U9490 ( .A(n9521), .B(n9522), .Z(n9902) );
  AND U9491 ( .A(n9903), .B(n9904), .Z(n9522) );
  NANDN U9492 ( .A(n9905), .B(n9906), .Z(n9904) );
  NANDN U9493 ( .A(n9907), .B(n9908), .Z(n9903) );
  NANDN U9494 ( .A(n9906), .B(n9905), .Z(n9908) );
  ANDN U9495 ( .B(\stack[1][28] ), .A(n5950), .Z(n9521) );
  XNOR U9496 ( .A(n9527), .B(n9909), .Z(n9520) );
  XNOR U9497 ( .A(n9528), .B(n9529), .Z(n9909) );
  AND U9498 ( .A(n9910), .B(n9911), .Z(n9529) );
  NAND U9499 ( .A(n9912), .B(n9913), .Z(n9911) );
  NANDN U9500 ( .A(n9914), .B(n9915), .Z(n9910) );
  OR U9501 ( .A(n9912), .B(n9913), .Z(n9915) );
  ANDN U9502 ( .B(\stack[1][29] ), .A(n5926), .Z(n9528) );
  XNOR U9503 ( .A(n9534), .B(n9916), .Z(n9527) );
  XNOR U9504 ( .A(n9535), .B(n9536), .Z(n9916) );
  AND U9505 ( .A(n9917), .B(n9918), .Z(n9536) );
  NANDN U9506 ( .A(n9919), .B(n9920), .Z(n9918) );
  NANDN U9507 ( .A(n9921), .B(n9922), .Z(n9917) );
  NANDN U9508 ( .A(n9920), .B(n9919), .Z(n9922) );
  ANDN U9509 ( .B(\stack[1][30] ), .A(n5902), .Z(n9535) );
  XNOR U9510 ( .A(n9541), .B(n9923), .Z(n9534) );
  XNOR U9511 ( .A(n9542), .B(n9543), .Z(n9923) );
  AND U9512 ( .A(n9924), .B(n9925), .Z(n9543) );
  NAND U9513 ( .A(n9926), .B(n9927), .Z(n9925) );
  NANDN U9514 ( .A(n9928), .B(n9929), .Z(n9924) );
  OR U9515 ( .A(n9926), .B(n9927), .Z(n9929) );
  ANDN U9516 ( .B(\stack[1][31] ), .A(n5878), .Z(n9542) );
  XNOR U9517 ( .A(n9548), .B(n9930), .Z(n9541) );
  XNOR U9518 ( .A(n9549), .B(n9550), .Z(n9930) );
  AND U9519 ( .A(n9931), .B(n9932), .Z(n9550) );
  NANDN U9520 ( .A(n9933), .B(n9934), .Z(n9932) );
  NANDN U9521 ( .A(n9935), .B(n9936), .Z(n9931) );
  NANDN U9522 ( .A(n9934), .B(n9933), .Z(n9936) );
  ANDN U9523 ( .B(\stack[1][32] ), .A(n5854), .Z(n9549) );
  XNOR U9524 ( .A(n9555), .B(n9937), .Z(n9548) );
  XNOR U9525 ( .A(n9556), .B(n9557), .Z(n9937) );
  AND U9526 ( .A(n9938), .B(n9939), .Z(n9557) );
  NAND U9527 ( .A(n9940), .B(n9941), .Z(n9939) );
  NANDN U9528 ( .A(n9942), .B(n9943), .Z(n9938) );
  OR U9529 ( .A(n9940), .B(n9941), .Z(n9943) );
  ANDN U9530 ( .B(\stack[1][33] ), .A(n5830), .Z(n9556) );
  XNOR U9531 ( .A(n9562), .B(n9944), .Z(n9555) );
  XNOR U9532 ( .A(n9563), .B(n9564), .Z(n9944) );
  AND U9533 ( .A(n9945), .B(n9946), .Z(n9564) );
  NANDN U9534 ( .A(n9947), .B(n9948), .Z(n9946) );
  NANDN U9535 ( .A(n9949), .B(n9950), .Z(n9945) );
  NANDN U9536 ( .A(n9948), .B(n9947), .Z(n9950) );
  ANDN U9537 ( .B(\stack[1][34] ), .A(n5806), .Z(n9563) );
  XNOR U9538 ( .A(n9569), .B(n9951), .Z(n9562) );
  XNOR U9539 ( .A(n9570), .B(n9571), .Z(n9951) );
  AND U9540 ( .A(n9952), .B(n9953), .Z(n9571) );
  NAND U9541 ( .A(n9954), .B(n9955), .Z(n9953) );
  NANDN U9542 ( .A(n9956), .B(n9957), .Z(n9952) );
  OR U9543 ( .A(n9954), .B(n9955), .Z(n9957) );
  ANDN U9544 ( .B(\stack[1][35] ), .A(n5782), .Z(n9570) );
  XNOR U9545 ( .A(n9576), .B(n9958), .Z(n9569) );
  XNOR U9546 ( .A(n9577), .B(n9578), .Z(n9958) );
  AND U9547 ( .A(n9959), .B(n9960), .Z(n9578) );
  NANDN U9548 ( .A(n9961), .B(n9962), .Z(n9960) );
  NANDN U9549 ( .A(n9963), .B(n9964), .Z(n9959) );
  NANDN U9550 ( .A(n9962), .B(n9961), .Z(n9964) );
  ANDN U9551 ( .B(\stack[1][36] ), .A(n5758), .Z(n9577) );
  XNOR U9552 ( .A(n9583), .B(n9965), .Z(n9576) );
  XOR U9553 ( .A(n9585), .B(n9586), .Z(n9965) );
  NAND U9554 ( .A(n9966), .B(n9967), .Z(n9586) );
  NAND U9555 ( .A(n9968), .B(n9969), .Z(n9967) );
  OR U9556 ( .A(n9970), .B(n9971), .Z(n9968) );
  AND U9557 ( .A(\stack[0][24] ), .B(\stack[1][37] ), .Z(n9585) );
  XNOR U9558 ( .A(n9592), .B(n9972), .Z(n9583) );
  XOR U9559 ( .A(n9593), .B(n9591), .Z(n9972) );
  AND U9560 ( .A(\stack[0][23] ), .B(\stack[1][38] ), .Z(n9591) );
  NAND U9561 ( .A(n9973), .B(n9974), .Z(n9593) );
  OR U9562 ( .A(n9975), .B(n9976), .Z(n9974) );
  NAND U9563 ( .A(n9977), .B(n9978), .Z(n9973) );
  NAND U9564 ( .A(n9976), .B(n9975), .Z(n9977) );
  XNOR U9565 ( .A(n9597), .B(n9979), .Z(n9592) );
  XNOR U9566 ( .A(n9598), .B(n9599), .Z(n9979) );
  AND U9567 ( .A(n9980), .B(n9981), .Z(n9599) );
  NAND U9568 ( .A(n9982), .B(n9983), .Z(n9981) );
  NANDN U9569 ( .A(n9984), .B(n9985), .Z(n9980) );
  OR U9570 ( .A(n9982), .B(n9983), .Z(n9985) );
  ANDN U9571 ( .B(\stack[1][39] ), .A(n5686), .Z(n9598) );
  XNOR U9572 ( .A(n9604), .B(n9986), .Z(n9597) );
  XNOR U9573 ( .A(n9605), .B(n9606), .Z(n9986) );
  AND U9574 ( .A(n9987), .B(n9988), .Z(n9606) );
  NANDN U9575 ( .A(n9989), .B(n9990), .Z(n9988) );
  NANDN U9576 ( .A(n9991), .B(n9992), .Z(n9987) );
  NANDN U9577 ( .A(n9990), .B(n9989), .Z(n9992) );
  ANDN U9578 ( .B(\stack[1][40] ), .A(n5662), .Z(n9605) );
  XNOR U9579 ( .A(n9611), .B(n9993), .Z(n9604) );
  XNOR U9580 ( .A(n9612), .B(n9613), .Z(n9993) );
  AND U9581 ( .A(n9994), .B(n9995), .Z(n9613) );
  NAND U9582 ( .A(n9996), .B(n9997), .Z(n9995) );
  NANDN U9583 ( .A(n9998), .B(n9999), .Z(n9994) );
  OR U9584 ( .A(n9996), .B(n9997), .Z(n9999) );
  ANDN U9585 ( .B(\stack[1][41] ), .A(n5638), .Z(n9612) );
  XNOR U9586 ( .A(n9618), .B(n10000), .Z(n9611) );
  XNOR U9587 ( .A(n9619), .B(n9620), .Z(n10000) );
  AND U9588 ( .A(n10001), .B(n10002), .Z(n9620) );
  NANDN U9589 ( .A(n10003), .B(n10004), .Z(n10002) );
  NANDN U9590 ( .A(n10005), .B(n10006), .Z(n10001) );
  NANDN U9591 ( .A(n10004), .B(n10003), .Z(n10006) );
  ANDN U9592 ( .B(\stack[1][42] ), .A(n5614), .Z(n9619) );
  XNOR U9593 ( .A(n9625), .B(n10007), .Z(n9618) );
  XNOR U9594 ( .A(n9626), .B(n9627), .Z(n10007) );
  AND U9595 ( .A(n10008), .B(n10009), .Z(n9627) );
  NAND U9596 ( .A(n10010), .B(n10011), .Z(n10009) );
  NANDN U9597 ( .A(n10012), .B(n10013), .Z(n10008) );
  OR U9598 ( .A(n10010), .B(n10011), .Z(n10013) );
  ANDN U9599 ( .B(\stack[1][43] ), .A(n5590), .Z(n9626) );
  XNOR U9600 ( .A(n9632), .B(n10014), .Z(n9625) );
  XNOR U9601 ( .A(n9633), .B(n9634), .Z(n10014) );
  AND U9602 ( .A(n10015), .B(n10016), .Z(n9634) );
  NANDN U9603 ( .A(n10017), .B(n10018), .Z(n10016) );
  NANDN U9604 ( .A(n10019), .B(n10020), .Z(n10015) );
  NANDN U9605 ( .A(n10018), .B(n10017), .Z(n10020) );
  ANDN U9606 ( .B(\stack[1][44] ), .A(n5566), .Z(n9633) );
  XNOR U9607 ( .A(n9639), .B(n10021), .Z(n9632) );
  XNOR U9608 ( .A(n9640), .B(n9641), .Z(n10021) );
  AND U9609 ( .A(n10022), .B(n10023), .Z(n9641) );
  NAND U9610 ( .A(n10024), .B(n10025), .Z(n10023) );
  NANDN U9611 ( .A(n10026), .B(n10027), .Z(n10022) );
  OR U9612 ( .A(n10024), .B(n10025), .Z(n10027) );
  ANDN U9613 ( .B(\stack[1][45] ), .A(n5542), .Z(n9640) );
  XNOR U9614 ( .A(n9646), .B(n10028), .Z(n9639) );
  XNOR U9615 ( .A(n9647), .B(n9648), .Z(n10028) );
  AND U9616 ( .A(n10029), .B(n10030), .Z(n9648) );
  NANDN U9617 ( .A(n10031), .B(n10032), .Z(n10030) );
  NANDN U9618 ( .A(n10033), .B(n10034), .Z(n10029) );
  NANDN U9619 ( .A(n10032), .B(n10031), .Z(n10034) );
  ANDN U9620 ( .B(\stack[1][46] ), .A(n5518), .Z(n9647) );
  XNOR U9621 ( .A(n9653), .B(n10035), .Z(n9646) );
  XNOR U9622 ( .A(n9654), .B(n9655), .Z(n10035) );
  AND U9623 ( .A(n10036), .B(n10037), .Z(n9655) );
  NAND U9624 ( .A(n10038), .B(n10039), .Z(n10037) );
  NANDN U9625 ( .A(n10040), .B(n10041), .Z(n10036) );
  OR U9626 ( .A(n10038), .B(n10039), .Z(n10041) );
  ANDN U9627 ( .B(\stack[1][47] ), .A(n5494), .Z(n9654) );
  XNOR U9628 ( .A(n9660), .B(n10042), .Z(n9653) );
  XNOR U9629 ( .A(n9661), .B(n9662), .Z(n10042) );
  AND U9630 ( .A(n10043), .B(n10044), .Z(n9662) );
  NANDN U9631 ( .A(n10045), .B(n10046), .Z(n10044) );
  NANDN U9632 ( .A(n10047), .B(n10048), .Z(n10043) );
  NANDN U9633 ( .A(n10046), .B(n10045), .Z(n10048) );
  ANDN U9634 ( .B(\stack[1][48] ), .A(n5470), .Z(n9661) );
  XNOR U9635 ( .A(n9667), .B(n10049), .Z(n9660) );
  XNOR U9636 ( .A(n9668), .B(n9669), .Z(n10049) );
  AND U9637 ( .A(n10050), .B(n10051), .Z(n9669) );
  NAND U9638 ( .A(n10052), .B(n10053), .Z(n10051) );
  NANDN U9639 ( .A(n10054), .B(n10055), .Z(n10050) );
  OR U9640 ( .A(n10052), .B(n10053), .Z(n10055) );
  ANDN U9641 ( .B(\stack[1][49] ), .A(n5446), .Z(n9668) );
  XNOR U9642 ( .A(n9674), .B(n10056), .Z(n9667) );
  XNOR U9643 ( .A(n9675), .B(n9676), .Z(n10056) );
  AND U9644 ( .A(n10057), .B(n10058), .Z(n9676) );
  NANDN U9645 ( .A(n10059), .B(n10060), .Z(n10058) );
  NANDN U9646 ( .A(n10061), .B(n10062), .Z(n10057) );
  NANDN U9647 ( .A(n10060), .B(n10059), .Z(n10062) );
  ANDN U9648 ( .B(\stack[1][50] ), .A(n5422), .Z(n9675) );
  XNOR U9649 ( .A(n9681), .B(n10063), .Z(n9674) );
  XNOR U9650 ( .A(n9682), .B(n9683), .Z(n10063) );
  AND U9651 ( .A(n10064), .B(n10065), .Z(n9683) );
  NAND U9652 ( .A(n10066), .B(n10067), .Z(n10065) );
  NANDN U9653 ( .A(n10068), .B(n10069), .Z(n10064) );
  OR U9654 ( .A(n10066), .B(n10067), .Z(n10069) );
  ANDN U9655 ( .B(\stack[1][51] ), .A(n5398), .Z(n9682) );
  XNOR U9656 ( .A(n9688), .B(n10070), .Z(n9681) );
  XNOR U9657 ( .A(n9689), .B(n9690), .Z(n10070) );
  AND U9658 ( .A(n10071), .B(n10072), .Z(n9690) );
  NANDN U9659 ( .A(n10073), .B(n10074), .Z(n10072) );
  NANDN U9660 ( .A(n10075), .B(n10076), .Z(n10071) );
  NANDN U9661 ( .A(n10074), .B(n10073), .Z(n10076) );
  ANDN U9662 ( .B(\stack[1][52] ), .A(n5374), .Z(n9689) );
  XNOR U9663 ( .A(n9695), .B(n10077), .Z(n9688) );
  XNOR U9664 ( .A(n9696), .B(n9697), .Z(n10077) );
  AND U9665 ( .A(n10078), .B(n10079), .Z(n9697) );
  NAND U9666 ( .A(n10080), .B(n10081), .Z(n10079) );
  NANDN U9667 ( .A(n10082), .B(n10083), .Z(n10078) );
  OR U9668 ( .A(n10080), .B(n10081), .Z(n10083) );
  ANDN U9669 ( .B(\stack[1][53] ), .A(n5350), .Z(n9696) );
  XNOR U9670 ( .A(n9702), .B(n10084), .Z(n9695) );
  XNOR U9671 ( .A(n9703), .B(n9704), .Z(n10084) );
  AND U9672 ( .A(n10085), .B(n10086), .Z(n9704) );
  NANDN U9673 ( .A(n10087), .B(n10088), .Z(n10086) );
  NANDN U9674 ( .A(n10089), .B(n10090), .Z(n10085) );
  NANDN U9675 ( .A(n10088), .B(n10087), .Z(n10090) );
  ANDN U9676 ( .B(\stack[1][54] ), .A(n5326), .Z(n9703) );
  XNOR U9677 ( .A(n9709), .B(n10091), .Z(n9702) );
  XNOR U9678 ( .A(n9710), .B(n9711), .Z(n10091) );
  AND U9679 ( .A(n10092), .B(n10093), .Z(n9711) );
  NAND U9680 ( .A(n10094), .B(n10095), .Z(n10093) );
  NANDN U9681 ( .A(n10096), .B(n10097), .Z(n10092) );
  OR U9682 ( .A(n10094), .B(n10095), .Z(n10097) );
  ANDN U9683 ( .B(\stack[1][55] ), .A(n5302), .Z(n9710) );
  XNOR U9684 ( .A(n9716), .B(n10098), .Z(n9709) );
  XNOR U9685 ( .A(n9717), .B(n9718), .Z(n10098) );
  AND U9686 ( .A(n10099), .B(n10100), .Z(n9718) );
  NANDN U9687 ( .A(n10101), .B(n10102), .Z(n10100) );
  NANDN U9688 ( .A(n10103), .B(n10104), .Z(n10099) );
  NANDN U9689 ( .A(n10102), .B(n10101), .Z(n10104) );
  ANDN U9690 ( .B(\stack[1][56] ), .A(n5278), .Z(n9717) );
  XNOR U9691 ( .A(n9723), .B(n10105), .Z(n9716) );
  XNOR U9692 ( .A(n9724), .B(n9725), .Z(n10105) );
  AND U9693 ( .A(n10106), .B(n10107), .Z(n9725) );
  NAND U9694 ( .A(n10108), .B(n10109), .Z(n10107) );
  NANDN U9695 ( .A(n10110), .B(n10111), .Z(n10106) );
  OR U9696 ( .A(n10108), .B(n10109), .Z(n10111) );
  ANDN U9697 ( .B(\stack[1][57] ), .A(n5254), .Z(n9724) );
  XNOR U9698 ( .A(n9730), .B(n10112), .Z(n9723) );
  XNOR U9699 ( .A(n9731), .B(n9732), .Z(n10112) );
  AND U9700 ( .A(n10113), .B(n10114), .Z(n9732) );
  NAND U9701 ( .A(n10115), .B(n10116), .Z(n10114) );
  NAND U9702 ( .A(n10117), .B(n10118), .Z(n10113) );
  OR U9703 ( .A(n10115), .B(n10116), .Z(n10117) );
  ANDN U9704 ( .B(\stack[1][58] ), .A(n5230), .Z(n9731) );
  XNOR U9705 ( .A(n9737), .B(n10119), .Z(n9730) );
  XNOR U9706 ( .A(n9738), .B(n9740), .Z(n10119) );
  ANDN U9707 ( .B(n10120), .A(n10121), .Z(n9740) );
  ANDN U9708 ( .B(\stack[0][0] ), .A(n6612), .Z(n10120) );
  ANDN U9709 ( .B(\stack[1][59] ), .A(n5206), .Z(n9738) );
  XOR U9710 ( .A(n9742), .B(n10122), .Z(n9737) );
  NANDN U9711 ( .A(n5160), .B(\stack[1][61] ), .Z(n10122) );
  NANDN U9712 ( .A(n6612), .B(\stack[0][1] ), .Z(n9742) );
  ANDN U9713 ( .B(\stack[1][5] ), .A(n6502), .Z(n8970) );
  AND U9714 ( .A(n10123), .B(n10124), .Z(n8971) );
  NANDN U9715 ( .A(n8975), .B(n8977), .Z(n10124) );
  NANDN U9716 ( .A(n8978), .B(n10125), .Z(n10123) );
  NANDN U9717 ( .A(n8977), .B(n8975), .Z(n10125) );
  XOR U9718 ( .A(n9751), .B(n10126), .Z(n8975) );
  XNOR U9719 ( .A(n9752), .B(n9753), .Z(n10126) );
  AND U9720 ( .A(n10127), .B(n10128), .Z(n9753) );
  NAND U9721 ( .A(n10129), .B(n10130), .Z(n10128) );
  NANDN U9722 ( .A(n10131), .B(n10132), .Z(n10127) );
  OR U9723 ( .A(n10129), .B(n10130), .Z(n10132) );
  ANDN U9724 ( .B(\stack[0][54] ), .A(n5316), .Z(n9752) );
  XNOR U9725 ( .A(n9758), .B(n10133), .Z(n9751) );
  XNOR U9726 ( .A(n9759), .B(n9760), .Z(n10133) );
  AND U9727 ( .A(n10134), .B(n10135), .Z(n9760) );
  NANDN U9728 ( .A(n10136), .B(n10137), .Z(n10135) );
  NANDN U9729 ( .A(n10138), .B(n10139), .Z(n10134) );
  NANDN U9730 ( .A(n10137), .B(n10136), .Z(n10139) );
  ANDN U9731 ( .B(\stack[0][53] ), .A(n5340), .Z(n9759) );
  XNOR U9732 ( .A(n9765), .B(n10140), .Z(n9758) );
  XNOR U9733 ( .A(n9766), .B(n9767), .Z(n10140) );
  AND U9734 ( .A(n10141), .B(n10142), .Z(n9767) );
  NAND U9735 ( .A(n10143), .B(n10144), .Z(n10142) );
  NANDN U9736 ( .A(n10145), .B(n10146), .Z(n10141) );
  OR U9737 ( .A(n10143), .B(n10144), .Z(n10146) );
  ANDN U9738 ( .B(\stack[0][52] ), .A(n5364), .Z(n9766) );
  XNOR U9739 ( .A(n9772), .B(n10147), .Z(n9765) );
  XNOR U9740 ( .A(n9773), .B(n9774), .Z(n10147) );
  AND U9741 ( .A(n10148), .B(n10149), .Z(n9774) );
  NANDN U9742 ( .A(n10150), .B(n10151), .Z(n10149) );
  NANDN U9743 ( .A(n10152), .B(n10153), .Z(n10148) );
  NANDN U9744 ( .A(n10151), .B(n10150), .Z(n10153) );
  ANDN U9745 ( .B(\stack[0][51] ), .A(n5387), .Z(n9773) );
  XNOR U9746 ( .A(n9779), .B(n10154), .Z(n9772) );
  XNOR U9747 ( .A(n9780), .B(n9781), .Z(n10154) );
  AND U9748 ( .A(n10155), .B(n10156), .Z(n9781) );
  NAND U9749 ( .A(n10157), .B(n10158), .Z(n10156) );
  NANDN U9750 ( .A(n10159), .B(n10160), .Z(n10155) );
  OR U9751 ( .A(n10157), .B(n10158), .Z(n10160) );
  ANDN U9752 ( .B(\stack[1][10] ), .A(n6358), .Z(n9780) );
  XNOR U9753 ( .A(n9786), .B(n10161), .Z(n9779) );
  XNOR U9754 ( .A(n9787), .B(n9788), .Z(n10161) );
  AND U9755 ( .A(n10162), .B(n10163), .Z(n9788) );
  NANDN U9756 ( .A(n10164), .B(n10165), .Z(n10163) );
  NANDN U9757 ( .A(n10166), .B(n10167), .Z(n10162) );
  NANDN U9758 ( .A(n10165), .B(n10164), .Z(n10167) );
  ANDN U9759 ( .B(\stack[1][11] ), .A(n6334), .Z(n9787) );
  XNOR U9760 ( .A(n9793), .B(n10168), .Z(n9786) );
  XNOR U9761 ( .A(n9794), .B(n9795), .Z(n10168) );
  AND U9762 ( .A(n10169), .B(n10170), .Z(n9795) );
  NAND U9763 ( .A(n10171), .B(n10172), .Z(n10170) );
  NANDN U9764 ( .A(n10173), .B(n10174), .Z(n10169) );
  OR U9765 ( .A(n10171), .B(n10172), .Z(n10174) );
  ANDN U9766 ( .B(\stack[1][12] ), .A(n6310), .Z(n9794) );
  XNOR U9767 ( .A(n9800), .B(n10175), .Z(n9793) );
  XNOR U9768 ( .A(n9801), .B(n9802), .Z(n10175) );
  AND U9769 ( .A(n10176), .B(n10177), .Z(n9802) );
  NANDN U9770 ( .A(n10178), .B(n10179), .Z(n10177) );
  NANDN U9771 ( .A(n10180), .B(n10181), .Z(n10176) );
  NANDN U9772 ( .A(n10179), .B(n10178), .Z(n10181) );
  ANDN U9773 ( .B(\stack[1][13] ), .A(n6286), .Z(n9801) );
  XNOR U9774 ( .A(n9807), .B(n10182), .Z(n9800) );
  XNOR U9775 ( .A(n9808), .B(n9809), .Z(n10182) );
  AND U9776 ( .A(n10183), .B(n10184), .Z(n9809) );
  NAND U9777 ( .A(n10185), .B(n10186), .Z(n10184) );
  NANDN U9778 ( .A(n10187), .B(n10188), .Z(n10183) );
  OR U9779 ( .A(n10185), .B(n10186), .Z(n10188) );
  ANDN U9780 ( .B(\stack[1][14] ), .A(n6262), .Z(n9808) );
  XNOR U9781 ( .A(n9814), .B(n10189), .Z(n9807) );
  XNOR U9782 ( .A(n9815), .B(n9816), .Z(n10189) );
  AND U9783 ( .A(n10190), .B(n10191), .Z(n9816) );
  NANDN U9784 ( .A(n10192), .B(n10193), .Z(n10191) );
  NANDN U9785 ( .A(n10194), .B(n10195), .Z(n10190) );
  NANDN U9786 ( .A(n10193), .B(n10192), .Z(n10195) );
  ANDN U9787 ( .B(\stack[1][15] ), .A(n6238), .Z(n9815) );
  XNOR U9788 ( .A(n9821), .B(n10196), .Z(n9814) );
  XNOR U9789 ( .A(n9822), .B(n9823), .Z(n10196) );
  AND U9790 ( .A(n10197), .B(n10198), .Z(n9823) );
  NAND U9791 ( .A(n10199), .B(n10200), .Z(n10198) );
  NANDN U9792 ( .A(n10201), .B(n10202), .Z(n10197) );
  OR U9793 ( .A(n10199), .B(n10200), .Z(n10202) );
  ANDN U9794 ( .B(\stack[1][16] ), .A(n6214), .Z(n9822) );
  XNOR U9795 ( .A(n9828), .B(n10203), .Z(n9821) );
  XNOR U9796 ( .A(n9829), .B(n9830), .Z(n10203) );
  AND U9797 ( .A(n10204), .B(n10205), .Z(n9830) );
  NANDN U9798 ( .A(n10206), .B(n10207), .Z(n10205) );
  NANDN U9799 ( .A(n10208), .B(n10209), .Z(n10204) );
  NANDN U9800 ( .A(n10207), .B(n10206), .Z(n10209) );
  ANDN U9801 ( .B(\stack[1][17] ), .A(n6190), .Z(n9829) );
  XNOR U9802 ( .A(n9835), .B(n10210), .Z(n9828) );
  XNOR U9803 ( .A(n9836), .B(n9837), .Z(n10210) );
  AND U9804 ( .A(n10211), .B(n10212), .Z(n9837) );
  NAND U9805 ( .A(n10213), .B(n10214), .Z(n10212) );
  NANDN U9806 ( .A(n10215), .B(n10216), .Z(n10211) );
  OR U9807 ( .A(n10213), .B(n10214), .Z(n10216) );
  ANDN U9808 ( .B(\stack[1][18] ), .A(n6166), .Z(n9836) );
  XNOR U9809 ( .A(n9842), .B(n10217), .Z(n9835) );
  XNOR U9810 ( .A(n9843), .B(n9844), .Z(n10217) );
  AND U9811 ( .A(n10218), .B(n10219), .Z(n9844) );
  NANDN U9812 ( .A(n10220), .B(n10221), .Z(n10219) );
  NANDN U9813 ( .A(n10222), .B(n10223), .Z(n10218) );
  NANDN U9814 ( .A(n10221), .B(n10220), .Z(n10223) );
  ANDN U9815 ( .B(\stack[1][19] ), .A(n6142), .Z(n9843) );
  XNOR U9816 ( .A(n9849), .B(n10224), .Z(n9842) );
  XNOR U9817 ( .A(n9850), .B(n9851), .Z(n10224) );
  AND U9818 ( .A(n10225), .B(n10226), .Z(n9851) );
  NAND U9819 ( .A(n10227), .B(n10228), .Z(n10226) );
  NANDN U9820 ( .A(n10229), .B(n10230), .Z(n10225) );
  OR U9821 ( .A(n10227), .B(n10228), .Z(n10230) );
  ANDN U9822 ( .B(\stack[1][20] ), .A(n6118), .Z(n9850) );
  XNOR U9823 ( .A(n9856), .B(n10231), .Z(n9849) );
  XNOR U9824 ( .A(n9857), .B(n9858), .Z(n10231) );
  AND U9825 ( .A(n10232), .B(n10233), .Z(n9858) );
  NANDN U9826 ( .A(n10234), .B(n10235), .Z(n10233) );
  NANDN U9827 ( .A(n10236), .B(n10237), .Z(n10232) );
  NANDN U9828 ( .A(n10235), .B(n10234), .Z(n10237) );
  ANDN U9829 ( .B(\stack[1][21] ), .A(n6094), .Z(n9857) );
  XNOR U9830 ( .A(n9863), .B(n10238), .Z(n9856) );
  XNOR U9831 ( .A(n9864), .B(n9865), .Z(n10238) );
  AND U9832 ( .A(n10239), .B(n10240), .Z(n9865) );
  NAND U9833 ( .A(n10241), .B(n10242), .Z(n10240) );
  NANDN U9834 ( .A(n10243), .B(n10244), .Z(n10239) );
  OR U9835 ( .A(n10241), .B(n10242), .Z(n10244) );
  ANDN U9836 ( .B(\stack[1][22] ), .A(n6070), .Z(n9864) );
  XNOR U9837 ( .A(n9870), .B(n10245), .Z(n9863) );
  XNOR U9838 ( .A(n9871), .B(n9872), .Z(n10245) );
  AND U9839 ( .A(n10246), .B(n10247), .Z(n9872) );
  NANDN U9840 ( .A(n10248), .B(n10249), .Z(n10247) );
  NANDN U9841 ( .A(n10250), .B(n10251), .Z(n10246) );
  NANDN U9842 ( .A(n10249), .B(n10248), .Z(n10251) );
  ANDN U9843 ( .B(\stack[1][23] ), .A(n6046), .Z(n9871) );
  XNOR U9844 ( .A(n9877), .B(n10252), .Z(n9870) );
  XNOR U9845 ( .A(n9878), .B(n9879), .Z(n10252) );
  AND U9846 ( .A(n10253), .B(n10254), .Z(n9879) );
  NAND U9847 ( .A(n10255), .B(n10256), .Z(n10254) );
  NANDN U9848 ( .A(n10257), .B(n10258), .Z(n10253) );
  OR U9849 ( .A(n10255), .B(n10256), .Z(n10258) );
  ANDN U9850 ( .B(\stack[1][24] ), .A(n6022), .Z(n9878) );
  XNOR U9851 ( .A(n9884), .B(n10259), .Z(n9877) );
  XNOR U9852 ( .A(n9885), .B(n9886), .Z(n10259) );
  AND U9853 ( .A(n10260), .B(n10261), .Z(n9886) );
  NANDN U9854 ( .A(n10262), .B(n10263), .Z(n10261) );
  NANDN U9855 ( .A(n10264), .B(n10265), .Z(n10260) );
  NANDN U9856 ( .A(n10263), .B(n10262), .Z(n10265) );
  ANDN U9857 ( .B(\stack[1][25] ), .A(n5998), .Z(n9885) );
  XNOR U9858 ( .A(n9891), .B(n10266), .Z(n9884) );
  XNOR U9859 ( .A(n9892), .B(n9893), .Z(n10266) );
  AND U9860 ( .A(n10267), .B(n10268), .Z(n9893) );
  NAND U9861 ( .A(n10269), .B(n10270), .Z(n10268) );
  NANDN U9862 ( .A(n10271), .B(n10272), .Z(n10267) );
  OR U9863 ( .A(n10269), .B(n10270), .Z(n10272) );
  ANDN U9864 ( .B(\stack[1][26] ), .A(n5974), .Z(n9892) );
  XNOR U9865 ( .A(n9898), .B(n10273), .Z(n9891) );
  XNOR U9866 ( .A(n9899), .B(n9900), .Z(n10273) );
  AND U9867 ( .A(n10274), .B(n10275), .Z(n9900) );
  NANDN U9868 ( .A(n10276), .B(n10277), .Z(n10275) );
  NANDN U9869 ( .A(n10278), .B(n10279), .Z(n10274) );
  NANDN U9870 ( .A(n10277), .B(n10276), .Z(n10279) );
  ANDN U9871 ( .B(\stack[1][27] ), .A(n5950), .Z(n9899) );
  XNOR U9872 ( .A(n9905), .B(n10280), .Z(n9898) );
  XNOR U9873 ( .A(n9906), .B(n9907), .Z(n10280) );
  AND U9874 ( .A(n10281), .B(n10282), .Z(n9907) );
  NAND U9875 ( .A(n10283), .B(n10284), .Z(n10282) );
  NANDN U9876 ( .A(n10285), .B(n10286), .Z(n10281) );
  OR U9877 ( .A(n10283), .B(n10284), .Z(n10286) );
  ANDN U9878 ( .B(\stack[1][28] ), .A(n5926), .Z(n9906) );
  XNOR U9879 ( .A(n9912), .B(n10287), .Z(n9905) );
  XNOR U9880 ( .A(n9913), .B(n9914), .Z(n10287) );
  AND U9881 ( .A(n10288), .B(n10289), .Z(n9914) );
  NANDN U9882 ( .A(n10290), .B(n10291), .Z(n10289) );
  NANDN U9883 ( .A(n10292), .B(n10293), .Z(n10288) );
  NANDN U9884 ( .A(n10291), .B(n10290), .Z(n10293) );
  ANDN U9885 ( .B(\stack[1][29] ), .A(n5902), .Z(n9913) );
  XNOR U9886 ( .A(n9919), .B(n10294), .Z(n9912) );
  XNOR U9887 ( .A(n9920), .B(n9921), .Z(n10294) );
  AND U9888 ( .A(n10295), .B(n10296), .Z(n9921) );
  NAND U9889 ( .A(n10297), .B(n10298), .Z(n10296) );
  NANDN U9890 ( .A(n10299), .B(n10300), .Z(n10295) );
  OR U9891 ( .A(n10297), .B(n10298), .Z(n10300) );
  ANDN U9892 ( .B(\stack[1][30] ), .A(n5878), .Z(n9920) );
  XNOR U9893 ( .A(n9926), .B(n10301), .Z(n9919) );
  XNOR U9894 ( .A(n9927), .B(n9928), .Z(n10301) );
  AND U9895 ( .A(n10302), .B(n10303), .Z(n9928) );
  NANDN U9896 ( .A(n10304), .B(n10305), .Z(n10303) );
  NANDN U9897 ( .A(n10306), .B(n10307), .Z(n10302) );
  NANDN U9898 ( .A(n10305), .B(n10304), .Z(n10307) );
  ANDN U9899 ( .B(\stack[1][31] ), .A(n5854), .Z(n9927) );
  XNOR U9900 ( .A(n9933), .B(n10308), .Z(n9926) );
  XNOR U9901 ( .A(n9934), .B(n9935), .Z(n10308) );
  AND U9902 ( .A(n10309), .B(n10310), .Z(n9935) );
  NAND U9903 ( .A(n10311), .B(n10312), .Z(n10310) );
  NANDN U9904 ( .A(n10313), .B(n10314), .Z(n10309) );
  OR U9905 ( .A(n10311), .B(n10312), .Z(n10314) );
  ANDN U9906 ( .B(\stack[1][32] ), .A(n5830), .Z(n9934) );
  XNOR U9907 ( .A(n9940), .B(n10315), .Z(n9933) );
  XNOR U9908 ( .A(n9941), .B(n9942), .Z(n10315) );
  AND U9909 ( .A(n10316), .B(n10317), .Z(n9942) );
  NANDN U9910 ( .A(n10318), .B(n10319), .Z(n10317) );
  NANDN U9911 ( .A(n10320), .B(n10321), .Z(n10316) );
  NANDN U9912 ( .A(n10319), .B(n10318), .Z(n10321) );
  ANDN U9913 ( .B(\stack[1][33] ), .A(n5806), .Z(n9941) );
  XNOR U9914 ( .A(n9947), .B(n10322), .Z(n9940) );
  XNOR U9915 ( .A(n9948), .B(n9949), .Z(n10322) );
  AND U9916 ( .A(n10323), .B(n10324), .Z(n9949) );
  NAND U9917 ( .A(n10325), .B(n10326), .Z(n10324) );
  NANDN U9918 ( .A(n10327), .B(n10328), .Z(n10323) );
  OR U9919 ( .A(n10325), .B(n10326), .Z(n10328) );
  ANDN U9920 ( .B(\stack[1][34] ), .A(n5782), .Z(n9948) );
  XNOR U9921 ( .A(n9954), .B(n10329), .Z(n9947) );
  XNOR U9922 ( .A(n9955), .B(n9956), .Z(n10329) );
  AND U9923 ( .A(n10330), .B(n10331), .Z(n9956) );
  NANDN U9924 ( .A(n10332), .B(n10333), .Z(n10331) );
  NANDN U9925 ( .A(n10334), .B(n10335), .Z(n10330) );
  NANDN U9926 ( .A(n10333), .B(n10332), .Z(n10335) );
  ANDN U9927 ( .B(\stack[1][35] ), .A(n5758), .Z(n9955) );
  XNOR U9928 ( .A(n9961), .B(n10336), .Z(n9954) );
  XNOR U9929 ( .A(n9962), .B(n9963), .Z(n10336) );
  AND U9930 ( .A(n10337), .B(n10338), .Z(n9963) );
  NAND U9931 ( .A(n10339), .B(n10340), .Z(n10338) );
  NANDN U9932 ( .A(n10341), .B(n10342), .Z(n10337) );
  OR U9933 ( .A(n10339), .B(n10340), .Z(n10342) );
  ANDN U9934 ( .B(\stack[1][36] ), .A(n5734), .Z(n9962) );
  XNOR U9935 ( .A(n9969), .B(n10343), .Z(n9961) );
  XOR U9936 ( .A(n9970), .B(n9971), .Z(n10343) );
  NAND U9937 ( .A(n10344), .B(n10345), .Z(n9971) );
  NANDN U9938 ( .A(n10346), .B(n10347), .Z(n10345) );
  OR U9939 ( .A(n10348), .B(n10349), .Z(n10347) );
  AND U9940 ( .A(\stack[0][23] ), .B(\stack[1][37] ), .Z(n9970) );
  XNOR U9941 ( .A(n9976), .B(n10350), .Z(n9969) );
  XNOR U9942 ( .A(n9975), .B(n9978), .Z(n10350) );
  AND U9943 ( .A(\stack[0][22] ), .B(\stack[1][38] ), .Z(n9978) );
  AND U9944 ( .A(n10351), .B(n10352), .Z(n9975) );
  NAND U9945 ( .A(n10353), .B(n10354), .Z(n10352) );
  OR U9946 ( .A(n10355), .B(n10356), .Z(n10353) );
  XNOR U9947 ( .A(n9982), .B(n10357), .Z(n9976) );
  XNOR U9948 ( .A(n9983), .B(n9984), .Z(n10357) );
  AND U9949 ( .A(n10358), .B(n10359), .Z(n9984) );
  NANDN U9950 ( .A(n10360), .B(n10361), .Z(n10359) );
  NANDN U9951 ( .A(n10362), .B(n10363), .Z(n10358) );
  NANDN U9952 ( .A(n10361), .B(n10360), .Z(n10363) );
  ANDN U9953 ( .B(\stack[1][39] ), .A(n5662), .Z(n9983) );
  XNOR U9954 ( .A(n9989), .B(n10364), .Z(n9982) );
  XNOR U9955 ( .A(n9990), .B(n9991), .Z(n10364) );
  AND U9956 ( .A(n10365), .B(n10366), .Z(n9991) );
  NAND U9957 ( .A(n10367), .B(n10368), .Z(n10366) );
  NANDN U9958 ( .A(n10369), .B(n10370), .Z(n10365) );
  OR U9959 ( .A(n10367), .B(n10368), .Z(n10370) );
  ANDN U9960 ( .B(\stack[1][40] ), .A(n5638), .Z(n9990) );
  XNOR U9961 ( .A(n9996), .B(n10371), .Z(n9989) );
  XNOR U9962 ( .A(n9997), .B(n9998), .Z(n10371) );
  AND U9963 ( .A(n10372), .B(n10373), .Z(n9998) );
  NANDN U9964 ( .A(n10374), .B(n10375), .Z(n10373) );
  NANDN U9965 ( .A(n10376), .B(n10377), .Z(n10372) );
  NANDN U9966 ( .A(n10375), .B(n10374), .Z(n10377) );
  ANDN U9967 ( .B(\stack[1][41] ), .A(n5614), .Z(n9997) );
  XNOR U9968 ( .A(n10003), .B(n10378), .Z(n9996) );
  XNOR U9969 ( .A(n10004), .B(n10005), .Z(n10378) );
  AND U9970 ( .A(n10379), .B(n10380), .Z(n10005) );
  NAND U9971 ( .A(n10381), .B(n10382), .Z(n10380) );
  NANDN U9972 ( .A(n10383), .B(n10384), .Z(n10379) );
  OR U9973 ( .A(n10381), .B(n10382), .Z(n10384) );
  ANDN U9974 ( .B(\stack[1][42] ), .A(n5590), .Z(n10004) );
  XNOR U9975 ( .A(n10010), .B(n10385), .Z(n10003) );
  XNOR U9976 ( .A(n10011), .B(n10012), .Z(n10385) );
  AND U9977 ( .A(n10386), .B(n10387), .Z(n10012) );
  NANDN U9978 ( .A(n10388), .B(n10389), .Z(n10387) );
  NANDN U9979 ( .A(n10390), .B(n10391), .Z(n10386) );
  NANDN U9980 ( .A(n10389), .B(n10388), .Z(n10391) );
  ANDN U9981 ( .B(\stack[1][43] ), .A(n5566), .Z(n10011) );
  XNOR U9982 ( .A(n10017), .B(n10392), .Z(n10010) );
  XNOR U9983 ( .A(n10018), .B(n10019), .Z(n10392) );
  AND U9984 ( .A(n10393), .B(n10394), .Z(n10019) );
  NAND U9985 ( .A(n10395), .B(n10396), .Z(n10394) );
  NANDN U9986 ( .A(n10397), .B(n10398), .Z(n10393) );
  OR U9987 ( .A(n10395), .B(n10396), .Z(n10398) );
  ANDN U9988 ( .B(\stack[1][44] ), .A(n5542), .Z(n10018) );
  XNOR U9989 ( .A(n10024), .B(n10399), .Z(n10017) );
  XNOR U9990 ( .A(n10025), .B(n10026), .Z(n10399) );
  AND U9991 ( .A(n10400), .B(n10401), .Z(n10026) );
  NANDN U9992 ( .A(n10402), .B(n10403), .Z(n10401) );
  NANDN U9993 ( .A(n10404), .B(n10405), .Z(n10400) );
  NANDN U9994 ( .A(n10403), .B(n10402), .Z(n10405) );
  ANDN U9995 ( .B(\stack[1][45] ), .A(n5518), .Z(n10025) );
  XNOR U9996 ( .A(n10031), .B(n10406), .Z(n10024) );
  XNOR U9997 ( .A(n10032), .B(n10033), .Z(n10406) );
  AND U9998 ( .A(n10407), .B(n10408), .Z(n10033) );
  NAND U9999 ( .A(n10409), .B(n10410), .Z(n10408) );
  NANDN U10000 ( .A(n10411), .B(n10412), .Z(n10407) );
  OR U10001 ( .A(n10409), .B(n10410), .Z(n10412) );
  ANDN U10002 ( .B(\stack[1][46] ), .A(n5494), .Z(n10032) );
  XNOR U10003 ( .A(n10038), .B(n10413), .Z(n10031) );
  XNOR U10004 ( .A(n10039), .B(n10040), .Z(n10413) );
  AND U10005 ( .A(n10414), .B(n10415), .Z(n10040) );
  NANDN U10006 ( .A(n10416), .B(n10417), .Z(n10415) );
  NANDN U10007 ( .A(n10418), .B(n10419), .Z(n10414) );
  NANDN U10008 ( .A(n10417), .B(n10416), .Z(n10419) );
  ANDN U10009 ( .B(\stack[1][47] ), .A(n5470), .Z(n10039) );
  XNOR U10010 ( .A(n10045), .B(n10420), .Z(n10038) );
  XNOR U10011 ( .A(n10046), .B(n10047), .Z(n10420) );
  AND U10012 ( .A(n10421), .B(n10422), .Z(n10047) );
  NAND U10013 ( .A(n10423), .B(n10424), .Z(n10422) );
  NANDN U10014 ( .A(n10425), .B(n10426), .Z(n10421) );
  OR U10015 ( .A(n10423), .B(n10424), .Z(n10426) );
  ANDN U10016 ( .B(\stack[1][48] ), .A(n5446), .Z(n10046) );
  XNOR U10017 ( .A(n10052), .B(n10427), .Z(n10045) );
  XNOR U10018 ( .A(n10053), .B(n10054), .Z(n10427) );
  AND U10019 ( .A(n10428), .B(n10429), .Z(n10054) );
  NANDN U10020 ( .A(n10430), .B(n10431), .Z(n10429) );
  NANDN U10021 ( .A(n10432), .B(n10433), .Z(n10428) );
  NANDN U10022 ( .A(n10431), .B(n10430), .Z(n10433) );
  ANDN U10023 ( .B(\stack[1][49] ), .A(n5422), .Z(n10053) );
  XNOR U10024 ( .A(n10059), .B(n10434), .Z(n10052) );
  XNOR U10025 ( .A(n10060), .B(n10061), .Z(n10434) );
  AND U10026 ( .A(n10435), .B(n10436), .Z(n10061) );
  NAND U10027 ( .A(n10437), .B(n10438), .Z(n10436) );
  NANDN U10028 ( .A(n10439), .B(n10440), .Z(n10435) );
  OR U10029 ( .A(n10437), .B(n10438), .Z(n10440) );
  ANDN U10030 ( .B(\stack[1][50] ), .A(n5398), .Z(n10060) );
  XNOR U10031 ( .A(n10066), .B(n10441), .Z(n10059) );
  XNOR U10032 ( .A(n10067), .B(n10068), .Z(n10441) );
  AND U10033 ( .A(n10442), .B(n10443), .Z(n10068) );
  NANDN U10034 ( .A(n10444), .B(n10445), .Z(n10443) );
  NANDN U10035 ( .A(n10446), .B(n10447), .Z(n10442) );
  NANDN U10036 ( .A(n10445), .B(n10444), .Z(n10447) );
  ANDN U10037 ( .B(\stack[1][51] ), .A(n5374), .Z(n10067) );
  XNOR U10038 ( .A(n10073), .B(n10448), .Z(n10066) );
  XNOR U10039 ( .A(n10074), .B(n10075), .Z(n10448) );
  AND U10040 ( .A(n10449), .B(n10450), .Z(n10075) );
  NAND U10041 ( .A(n10451), .B(n10452), .Z(n10450) );
  NANDN U10042 ( .A(n10453), .B(n10454), .Z(n10449) );
  OR U10043 ( .A(n10451), .B(n10452), .Z(n10454) );
  ANDN U10044 ( .B(\stack[1][52] ), .A(n5350), .Z(n10074) );
  XNOR U10045 ( .A(n10080), .B(n10455), .Z(n10073) );
  XNOR U10046 ( .A(n10081), .B(n10082), .Z(n10455) );
  AND U10047 ( .A(n10456), .B(n10457), .Z(n10082) );
  NANDN U10048 ( .A(n10458), .B(n10459), .Z(n10457) );
  NANDN U10049 ( .A(n10460), .B(n10461), .Z(n10456) );
  NANDN U10050 ( .A(n10459), .B(n10458), .Z(n10461) );
  ANDN U10051 ( .B(\stack[1][53] ), .A(n5326), .Z(n10081) );
  XNOR U10052 ( .A(n10087), .B(n10462), .Z(n10080) );
  XNOR U10053 ( .A(n10088), .B(n10089), .Z(n10462) );
  AND U10054 ( .A(n10463), .B(n10464), .Z(n10089) );
  NAND U10055 ( .A(n10465), .B(n10466), .Z(n10464) );
  NANDN U10056 ( .A(n10467), .B(n10468), .Z(n10463) );
  OR U10057 ( .A(n10465), .B(n10466), .Z(n10468) );
  ANDN U10058 ( .B(\stack[1][54] ), .A(n5302), .Z(n10088) );
  XNOR U10059 ( .A(n10094), .B(n10469), .Z(n10087) );
  XNOR U10060 ( .A(n10095), .B(n10096), .Z(n10469) );
  AND U10061 ( .A(n10470), .B(n10471), .Z(n10096) );
  NANDN U10062 ( .A(n10472), .B(n10473), .Z(n10471) );
  NANDN U10063 ( .A(n10474), .B(n10475), .Z(n10470) );
  NANDN U10064 ( .A(n10473), .B(n10472), .Z(n10475) );
  ANDN U10065 ( .B(\stack[1][55] ), .A(n5278), .Z(n10095) );
  XNOR U10066 ( .A(n10101), .B(n10476), .Z(n10094) );
  XNOR U10067 ( .A(n10102), .B(n10103), .Z(n10476) );
  AND U10068 ( .A(n10477), .B(n10478), .Z(n10103) );
  NAND U10069 ( .A(n10479), .B(n10480), .Z(n10478) );
  NANDN U10070 ( .A(n10481), .B(n10482), .Z(n10477) );
  OR U10071 ( .A(n10479), .B(n10480), .Z(n10482) );
  ANDN U10072 ( .B(\stack[1][56] ), .A(n5254), .Z(n10102) );
  XNOR U10073 ( .A(n10108), .B(n10483), .Z(n10101) );
  XNOR U10074 ( .A(n10109), .B(n10110), .Z(n10483) );
  AND U10075 ( .A(n10484), .B(n10485), .Z(n10110) );
  NAND U10076 ( .A(n10486), .B(n10487), .Z(n10485) );
  NAND U10077 ( .A(n10488), .B(n10489), .Z(n10484) );
  OR U10078 ( .A(n10486), .B(n10487), .Z(n10488) );
  ANDN U10079 ( .B(\stack[1][57] ), .A(n5230), .Z(n10109) );
  XNOR U10080 ( .A(n10115), .B(n10490), .Z(n10108) );
  XNOR U10081 ( .A(n10116), .B(n10118), .Z(n10490) );
  ANDN U10082 ( .B(n10491), .A(n10492), .Z(n10118) );
  ANDN U10083 ( .B(\stack[0][0] ), .A(n6588), .Z(n10491) );
  ANDN U10084 ( .B(\stack[1][58] ), .A(n5206), .Z(n10116) );
  XOR U10085 ( .A(n10121), .B(n10493), .Z(n10115) );
  NANDN U10086 ( .A(n5160), .B(\stack[1][60] ), .Z(n10493) );
  NANDN U10087 ( .A(n6588), .B(\stack[0][1] ), .Z(n10121) );
  ANDN U10088 ( .B(\stack[0][55] ), .A(n5292), .Z(n8977) );
  AND U10089 ( .A(n10494), .B(n10495), .Z(n8978) );
  NANDN U10090 ( .A(n8985), .B(n10496), .Z(n10494) );
  NANDN U10091 ( .A(n8984), .B(n8982), .Z(n10496) );
  XNOR U10092 ( .A(n10129), .B(n10497), .Z(n8982) );
  XNOR U10093 ( .A(n10130), .B(n10131), .Z(n10497) );
  AND U10094 ( .A(n10498), .B(n10499), .Z(n10131) );
  NANDN U10095 ( .A(n10500), .B(n10501), .Z(n10499) );
  NANDN U10096 ( .A(n10502), .B(n10503), .Z(n10498) );
  NANDN U10097 ( .A(n10501), .B(n10500), .Z(n10503) );
  ANDN U10098 ( .B(\stack[0][53] ), .A(n5316), .Z(n10130) );
  XNOR U10099 ( .A(n10136), .B(n10504), .Z(n10129) );
  XNOR U10100 ( .A(n10137), .B(n10138), .Z(n10504) );
  AND U10101 ( .A(n10505), .B(n10506), .Z(n10138) );
  NAND U10102 ( .A(n10507), .B(n10508), .Z(n10506) );
  NANDN U10103 ( .A(n10509), .B(n10510), .Z(n10505) );
  OR U10104 ( .A(n10507), .B(n10508), .Z(n10510) );
  ANDN U10105 ( .B(\stack[0][52] ), .A(n5340), .Z(n10137) );
  XNOR U10106 ( .A(n10143), .B(n10511), .Z(n10136) );
  XNOR U10107 ( .A(n10144), .B(n10145), .Z(n10511) );
  AND U10108 ( .A(n10512), .B(n10513), .Z(n10145) );
  NANDN U10109 ( .A(n10514), .B(n10515), .Z(n10513) );
  NANDN U10110 ( .A(n10516), .B(n10517), .Z(n10512) );
  NANDN U10111 ( .A(n10515), .B(n10514), .Z(n10517) );
  ANDN U10112 ( .B(\stack[0][51] ), .A(n5364), .Z(n10144) );
  XNOR U10113 ( .A(n10150), .B(n10518), .Z(n10143) );
  XNOR U10114 ( .A(n10151), .B(n10152), .Z(n10518) );
  AND U10115 ( .A(n10519), .B(n10520), .Z(n10152) );
  NAND U10116 ( .A(n10521), .B(n10522), .Z(n10520) );
  NANDN U10117 ( .A(n10523), .B(n10524), .Z(n10519) );
  OR U10118 ( .A(n10521), .B(n10522), .Z(n10524) );
  ANDN U10119 ( .B(\stack[0][50] ), .A(n5387), .Z(n10151) );
  XNOR U10120 ( .A(n10157), .B(n10525), .Z(n10150) );
  XNOR U10121 ( .A(n10158), .B(n10159), .Z(n10525) );
  AND U10122 ( .A(n10526), .B(n10527), .Z(n10159) );
  NANDN U10123 ( .A(n10528), .B(n10529), .Z(n10527) );
  NANDN U10124 ( .A(n10530), .B(n10531), .Z(n10526) );
  NANDN U10125 ( .A(n10529), .B(n10528), .Z(n10531) );
  ANDN U10126 ( .B(\stack[1][10] ), .A(n6334), .Z(n10158) );
  XNOR U10127 ( .A(n10164), .B(n10532), .Z(n10157) );
  XNOR U10128 ( .A(n10165), .B(n10166), .Z(n10532) );
  AND U10129 ( .A(n10533), .B(n10534), .Z(n10166) );
  NAND U10130 ( .A(n10535), .B(n10536), .Z(n10534) );
  NANDN U10131 ( .A(n10537), .B(n10538), .Z(n10533) );
  OR U10132 ( .A(n10535), .B(n10536), .Z(n10538) );
  ANDN U10133 ( .B(\stack[1][11] ), .A(n6310), .Z(n10165) );
  XNOR U10134 ( .A(n10171), .B(n10539), .Z(n10164) );
  XNOR U10135 ( .A(n10172), .B(n10173), .Z(n10539) );
  AND U10136 ( .A(n10540), .B(n10541), .Z(n10173) );
  NANDN U10137 ( .A(n10542), .B(n10543), .Z(n10541) );
  NANDN U10138 ( .A(n10544), .B(n10545), .Z(n10540) );
  NANDN U10139 ( .A(n10543), .B(n10542), .Z(n10545) );
  ANDN U10140 ( .B(\stack[1][12] ), .A(n6286), .Z(n10172) );
  XNOR U10141 ( .A(n10178), .B(n10546), .Z(n10171) );
  XNOR U10142 ( .A(n10179), .B(n10180), .Z(n10546) );
  AND U10143 ( .A(n10547), .B(n10548), .Z(n10180) );
  NAND U10144 ( .A(n10549), .B(n10550), .Z(n10548) );
  NANDN U10145 ( .A(n10551), .B(n10552), .Z(n10547) );
  OR U10146 ( .A(n10549), .B(n10550), .Z(n10552) );
  ANDN U10147 ( .B(\stack[1][13] ), .A(n6262), .Z(n10179) );
  XNOR U10148 ( .A(n10185), .B(n10553), .Z(n10178) );
  XNOR U10149 ( .A(n10186), .B(n10187), .Z(n10553) );
  AND U10150 ( .A(n10554), .B(n10555), .Z(n10187) );
  NANDN U10151 ( .A(n10556), .B(n10557), .Z(n10555) );
  NANDN U10152 ( .A(n10558), .B(n10559), .Z(n10554) );
  NANDN U10153 ( .A(n10557), .B(n10556), .Z(n10559) );
  ANDN U10154 ( .B(\stack[1][14] ), .A(n6238), .Z(n10186) );
  XNOR U10155 ( .A(n10192), .B(n10560), .Z(n10185) );
  XNOR U10156 ( .A(n10193), .B(n10194), .Z(n10560) );
  AND U10157 ( .A(n10561), .B(n10562), .Z(n10194) );
  NAND U10158 ( .A(n10563), .B(n10564), .Z(n10562) );
  NANDN U10159 ( .A(n10565), .B(n10566), .Z(n10561) );
  OR U10160 ( .A(n10563), .B(n10564), .Z(n10566) );
  ANDN U10161 ( .B(\stack[1][15] ), .A(n6214), .Z(n10193) );
  XNOR U10162 ( .A(n10199), .B(n10567), .Z(n10192) );
  XNOR U10163 ( .A(n10200), .B(n10201), .Z(n10567) );
  AND U10164 ( .A(n10568), .B(n10569), .Z(n10201) );
  NANDN U10165 ( .A(n10570), .B(n10571), .Z(n10569) );
  NANDN U10166 ( .A(n10572), .B(n10573), .Z(n10568) );
  NANDN U10167 ( .A(n10571), .B(n10570), .Z(n10573) );
  ANDN U10168 ( .B(\stack[1][16] ), .A(n6190), .Z(n10200) );
  XNOR U10169 ( .A(n10206), .B(n10574), .Z(n10199) );
  XNOR U10170 ( .A(n10207), .B(n10208), .Z(n10574) );
  AND U10171 ( .A(n10575), .B(n10576), .Z(n10208) );
  NAND U10172 ( .A(n10577), .B(n10578), .Z(n10576) );
  NANDN U10173 ( .A(n10579), .B(n10580), .Z(n10575) );
  OR U10174 ( .A(n10577), .B(n10578), .Z(n10580) );
  ANDN U10175 ( .B(\stack[1][17] ), .A(n6166), .Z(n10207) );
  XNOR U10176 ( .A(n10213), .B(n10581), .Z(n10206) );
  XNOR U10177 ( .A(n10214), .B(n10215), .Z(n10581) );
  AND U10178 ( .A(n10582), .B(n10583), .Z(n10215) );
  NANDN U10179 ( .A(n10584), .B(n10585), .Z(n10583) );
  NANDN U10180 ( .A(n10586), .B(n10587), .Z(n10582) );
  NANDN U10181 ( .A(n10585), .B(n10584), .Z(n10587) );
  ANDN U10182 ( .B(\stack[1][18] ), .A(n6142), .Z(n10214) );
  XNOR U10183 ( .A(n10220), .B(n10588), .Z(n10213) );
  XNOR U10184 ( .A(n10221), .B(n10222), .Z(n10588) );
  AND U10185 ( .A(n10589), .B(n10590), .Z(n10222) );
  NAND U10186 ( .A(n10591), .B(n10592), .Z(n10590) );
  NANDN U10187 ( .A(n10593), .B(n10594), .Z(n10589) );
  OR U10188 ( .A(n10591), .B(n10592), .Z(n10594) );
  ANDN U10189 ( .B(\stack[1][19] ), .A(n6118), .Z(n10221) );
  XNOR U10190 ( .A(n10227), .B(n10595), .Z(n10220) );
  XNOR U10191 ( .A(n10228), .B(n10229), .Z(n10595) );
  AND U10192 ( .A(n10596), .B(n10597), .Z(n10229) );
  NANDN U10193 ( .A(n10598), .B(n10599), .Z(n10597) );
  NANDN U10194 ( .A(n10600), .B(n10601), .Z(n10596) );
  NANDN U10195 ( .A(n10599), .B(n10598), .Z(n10601) );
  ANDN U10196 ( .B(\stack[1][20] ), .A(n6094), .Z(n10228) );
  XNOR U10197 ( .A(n10234), .B(n10602), .Z(n10227) );
  XNOR U10198 ( .A(n10235), .B(n10236), .Z(n10602) );
  AND U10199 ( .A(n10603), .B(n10604), .Z(n10236) );
  NAND U10200 ( .A(n10605), .B(n10606), .Z(n10604) );
  NANDN U10201 ( .A(n10607), .B(n10608), .Z(n10603) );
  OR U10202 ( .A(n10605), .B(n10606), .Z(n10608) );
  ANDN U10203 ( .B(\stack[1][21] ), .A(n6070), .Z(n10235) );
  XNOR U10204 ( .A(n10241), .B(n10609), .Z(n10234) );
  XNOR U10205 ( .A(n10242), .B(n10243), .Z(n10609) );
  AND U10206 ( .A(n10610), .B(n10611), .Z(n10243) );
  NANDN U10207 ( .A(n10612), .B(n10613), .Z(n10611) );
  NANDN U10208 ( .A(n10614), .B(n10615), .Z(n10610) );
  NANDN U10209 ( .A(n10613), .B(n10612), .Z(n10615) );
  ANDN U10210 ( .B(\stack[1][22] ), .A(n6046), .Z(n10242) );
  XNOR U10211 ( .A(n10248), .B(n10616), .Z(n10241) );
  XNOR U10212 ( .A(n10249), .B(n10250), .Z(n10616) );
  AND U10213 ( .A(n10617), .B(n10618), .Z(n10250) );
  NAND U10214 ( .A(n10619), .B(n10620), .Z(n10618) );
  NANDN U10215 ( .A(n10621), .B(n10622), .Z(n10617) );
  OR U10216 ( .A(n10619), .B(n10620), .Z(n10622) );
  ANDN U10217 ( .B(\stack[1][23] ), .A(n6022), .Z(n10249) );
  XNOR U10218 ( .A(n10255), .B(n10623), .Z(n10248) );
  XNOR U10219 ( .A(n10256), .B(n10257), .Z(n10623) );
  AND U10220 ( .A(n10624), .B(n10625), .Z(n10257) );
  NANDN U10221 ( .A(n10626), .B(n10627), .Z(n10625) );
  NANDN U10222 ( .A(n10628), .B(n10629), .Z(n10624) );
  NANDN U10223 ( .A(n10627), .B(n10626), .Z(n10629) );
  ANDN U10224 ( .B(\stack[1][24] ), .A(n5998), .Z(n10256) );
  XNOR U10225 ( .A(n10262), .B(n10630), .Z(n10255) );
  XNOR U10226 ( .A(n10263), .B(n10264), .Z(n10630) );
  AND U10227 ( .A(n10631), .B(n10632), .Z(n10264) );
  NAND U10228 ( .A(n10633), .B(n10634), .Z(n10632) );
  NANDN U10229 ( .A(n10635), .B(n10636), .Z(n10631) );
  OR U10230 ( .A(n10633), .B(n10634), .Z(n10636) );
  ANDN U10231 ( .B(\stack[1][25] ), .A(n5974), .Z(n10263) );
  XNOR U10232 ( .A(n10269), .B(n10637), .Z(n10262) );
  XNOR U10233 ( .A(n10270), .B(n10271), .Z(n10637) );
  AND U10234 ( .A(n10638), .B(n10639), .Z(n10271) );
  NANDN U10235 ( .A(n10640), .B(n10641), .Z(n10639) );
  NANDN U10236 ( .A(n10642), .B(n10643), .Z(n10638) );
  NANDN U10237 ( .A(n10641), .B(n10640), .Z(n10643) );
  ANDN U10238 ( .B(\stack[1][26] ), .A(n5950), .Z(n10270) );
  XNOR U10239 ( .A(n10276), .B(n10644), .Z(n10269) );
  XNOR U10240 ( .A(n10277), .B(n10278), .Z(n10644) );
  AND U10241 ( .A(n10645), .B(n10646), .Z(n10278) );
  NAND U10242 ( .A(n10647), .B(n10648), .Z(n10646) );
  NANDN U10243 ( .A(n10649), .B(n10650), .Z(n10645) );
  OR U10244 ( .A(n10647), .B(n10648), .Z(n10650) );
  ANDN U10245 ( .B(\stack[1][27] ), .A(n5926), .Z(n10277) );
  XNOR U10246 ( .A(n10283), .B(n10651), .Z(n10276) );
  XNOR U10247 ( .A(n10284), .B(n10285), .Z(n10651) );
  AND U10248 ( .A(n10652), .B(n10653), .Z(n10285) );
  NANDN U10249 ( .A(n10654), .B(n10655), .Z(n10653) );
  NANDN U10250 ( .A(n10656), .B(n10657), .Z(n10652) );
  NANDN U10251 ( .A(n10655), .B(n10654), .Z(n10657) );
  ANDN U10252 ( .B(\stack[1][28] ), .A(n5902), .Z(n10284) );
  XNOR U10253 ( .A(n10290), .B(n10658), .Z(n10283) );
  XNOR U10254 ( .A(n10291), .B(n10292), .Z(n10658) );
  AND U10255 ( .A(n10659), .B(n10660), .Z(n10292) );
  NAND U10256 ( .A(n10661), .B(n10662), .Z(n10660) );
  NANDN U10257 ( .A(n10663), .B(n10664), .Z(n10659) );
  OR U10258 ( .A(n10661), .B(n10662), .Z(n10664) );
  ANDN U10259 ( .B(\stack[1][29] ), .A(n5878), .Z(n10291) );
  XNOR U10260 ( .A(n10297), .B(n10665), .Z(n10290) );
  XNOR U10261 ( .A(n10298), .B(n10299), .Z(n10665) );
  AND U10262 ( .A(n10666), .B(n10667), .Z(n10299) );
  NANDN U10263 ( .A(n10668), .B(n10669), .Z(n10667) );
  NANDN U10264 ( .A(n10670), .B(n10671), .Z(n10666) );
  NANDN U10265 ( .A(n10669), .B(n10668), .Z(n10671) );
  ANDN U10266 ( .B(\stack[1][30] ), .A(n5854), .Z(n10298) );
  XNOR U10267 ( .A(n10304), .B(n10672), .Z(n10297) );
  XNOR U10268 ( .A(n10305), .B(n10306), .Z(n10672) );
  AND U10269 ( .A(n10673), .B(n10674), .Z(n10306) );
  NAND U10270 ( .A(n10675), .B(n10676), .Z(n10674) );
  NANDN U10271 ( .A(n10677), .B(n10678), .Z(n10673) );
  OR U10272 ( .A(n10675), .B(n10676), .Z(n10678) );
  ANDN U10273 ( .B(\stack[1][31] ), .A(n5830), .Z(n10305) );
  XNOR U10274 ( .A(n10311), .B(n10679), .Z(n10304) );
  XNOR U10275 ( .A(n10312), .B(n10313), .Z(n10679) );
  AND U10276 ( .A(n10680), .B(n10681), .Z(n10313) );
  NANDN U10277 ( .A(n10682), .B(n10683), .Z(n10681) );
  NANDN U10278 ( .A(n10684), .B(n10685), .Z(n10680) );
  NANDN U10279 ( .A(n10683), .B(n10682), .Z(n10685) );
  ANDN U10280 ( .B(\stack[1][32] ), .A(n5806), .Z(n10312) );
  XNOR U10281 ( .A(n10318), .B(n10686), .Z(n10311) );
  XNOR U10282 ( .A(n10319), .B(n10320), .Z(n10686) );
  AND U10283 ( .A(n10687), .B(n10688), .Z(n10320) );
  NAND U10284 ( .A(n10689), .B(n10690), .Z(n10688) );
  NANDN U10285 ( .A(n10691), .B(n10692), .Z(n10687) );
  OR U10286 ( .A(n10689), .B(n10690), .Z(n10692) );
  ANDN U10287 ( .B(\stack[1][33] ), .A(n5782), .Z(n10319) );
  XNOR U10288 ( .A(n10325), .B(n10693), .Z(n10318) );
  XNOR U10289 ( .A(n10326), .B(n10327), .Z(n10693) );
  AND U10290 ( .A(n10694), .B(n10695), .Z(n10327) );
  NANDN U10291 ( .A(n10696), .B(n10697), .Z(n10695) );
  NANDN U10292 ( .A(n10698), .B(n10699), .Z(n10694) );
  NANDN U10293 ( .A(n10697), .B(n10696), .Z(n10699) );
  ANDN U10294 ( .B(\stack[1][34] ), .A(n5758), .Z(n10326) );
  XNOR U10295 ( .A(n10332), .B(n10700), .Z(n10325) );
  XNOR U10296 ( .A(n10333), .B(n10334), .Z(n10700) );
  AND U10297 ( .A(n10701), .B(n10702), .Z(n10334) );
  NAND U10298 ( .A(n10703), .B(n10704), .Z(n10702) );
  NANDN U10299 ( .A(n10705), .B(n10706), .Z(n10701) );
  OR U10300 ( .A(n10703), .B(n10704), .Z(n10706) );
  ANDN U10301 ( .B(\stack[1][35] ), .A(n5734), .Z(n10333) );
  XNOR U10302 ( .A(n10339), .B(n10707), .Z(n10332) );
  XNOR U10303 ( .A(n10340), .B(n10341), .Z(n10707) );
  AND U10304 ( .A(n10708), .B(n10709), .Z(n10341) );
  NANDN U10305 ( .A(n10710), .B(n10711), .Z(n10709) );
  NANDN U10306 ( .A(n10712), .B(n10713), .Z(n10708) );
  NANDN U10307 ( .A(n10711), .B(n10710), .Z(n10713) );
  ANDN U10308 ( .B(\stack[1][36] ), .A(n5710), .Z(n10340) );
  XNOR U10309 ( .A(n10346), .B(n10714), .Z(n10339) );
  XOR U10310 ( .A(n10348), .B(n10349), .Z(n10714) );
  NAND U10311 ( .A(n10715), .B(n10716), .Z(n10349) );
  NAND U10312 ( .A(n10717), .B(n10718), .Z(n10716) );
  OR U10313 ( .A(n10719), .B(n10720), .Z(n10717) );
  AND U10314 ( .A(\stack[0][22] ), .B(\stack[1][37] ), .Z(n10348) );
  XNOR U10315 ( .A(n10355), .B(n10721), .Z(n10346) );
  XOR U10316 ( .A(n10356), .B(n10354), .Z(n10721) );
  AND U10317 ( .A(\stack[0][21] ), .B(\stack[1][38] ), .Z(n10354) );
  NAND U10318 ( .A(n10722), .B(n10723), .Z(n10356) );
  OR U10319 ( .A(n10724), .B(n10725), .Z(n10723) );
  NAND U10320 ( .A(n10726), .B(n10727), .Z(n10722) );
  NAND U10321 ( .A(n10725), .B(n10724), .Z(n10726) );
  XNOR U10322 ( .A(n10360), .B(n10728), .Z(n10355) );
  XNOR U10323 ( .A(n10361), .B(n10362), .Z(n10728) );
  AND U10324 ( .A(n10729), .B(n10730), .Z(n10362) );
  NAND U10325 ( .A(n10731), .B(n10732), .Z(n10730) );
  NANDN U10326 ( .A(n10733), .B(n10734), .Z(n10729) );
  OR U10327 ( .A(n10731), .B(n10732), .Z(n10734) );
  ANDN U10328 ( .B(\stack[1][39] ), .A(n5638), .Z(n10361) );
  XNOR U10329 ( .A(n10367), .B(n10735), .Z(n10360) );
  XNOR U10330 ( .A(n10368), .B(n10369), .Z(n10735) );
  AND U10331 ( .A(n10736), .B(n10737), .Z(n10369) );
  NANDN U10332 ( .A(n10738), .B(n10739), .Z(n10737) );
  NANDN U10333 ( .A(n10740), .B(n10741), .Z(n10736) );
  NANDN U10334 ( .A(n10739), .B(n10738), .Z(n10741) );
  ANDN U10335 ( .B(\stack[1][40] ), .A(n5614), .Z(n10368) );
  XNOR U10336 ( .A(n10374), .B(n10742), .Z(n10367) );
  XNOR U10337 ( .A(n10375), .B(n10376), .Z(n10742) );
  AND U10338 ( .A(n10743), .B(n10744), .Z(n10376) );
  NAND U10339 ( .A(n10745), .B(n10746), .Z(n10744) );
  NANDN U10340 ( .A(n10747), .B(n10748), .Z(n10743) );
  OR U10341 ( .A(n10745), .B(n10746), .Z(n10748) );
  ANDN U10342 ( .B(\stack[1][41] ), .A(n5590), .Z(n10375) );
  XNOR U10343 ( .A(n10381), .B(n10749), .Z(n10374) );
  XNOR U10344 ( .A(n10382), .B(n10383), .Z(n10749) );
  AND U10345 ( .A(n10750), .B(n10751), .Z(n10383) );
  NANDN U10346 ( .A(n10752), .B(n10753), .Z(n10751) );
  NANDN U10347 ( .A(n10754), .B(n10755), .Z(n10750) );
  NANDN U10348 ( .A(n10753), .B(n10752), .Z(n10755) );
  ANDN U10349 ( .B(\stack[1][42] ), .A(n5566), .Z(n10382) );
  XNOR U10350 ( .A(n10388), .B(n10756), .Z(n10381) );
  XNOR U10351 ( .A(n10389), .B(n10390), .Z(n10756) );
  AND U10352 ( .A(n10757), .B(n10758), .Z(n10390) );
  NAND U10353 ( .A(n10759), .B(n10760), .Z(n10758) );
  NANDN U10354 ( .A(n10761), .B(n10762), .Z(n10757) );
  OR U10355 ( .A(n10759), .B(n10760), .Z(n10762) );
  ANDN U10356 ( .B(\stack[1][43] ), .A(n5542), .Z(n10389) );
  XNOR U10357 ( .A(n10395), .B(n10763), .Z(n10388) );
  XNOR U10358 ( .A(n10396), .B(n10397), .Z(n10763) );
  AND U10359 ( .A(n10764), .B(n10765), .Z(n10397) );
  NANDN U10360 ( .A(n10766), .B(n10767), .Z(n10765) );
  NANDN U10361 ( .A(n10768), .B(n10769), .Z(n10764) );
  NANDN U10362 ( .A(n10767), .B(n10766), .Z(n10769) );
  ANDN U10363 ( .B(\stack[1][44] ), .A(n5518), .Z(n10396) );
  XNOR U10364 ( .A(n10402), .B(n10770), .Z(n10395) );
  XNOR U10365 ( .A(n10403), .B(n10404), .Z(n10770) );
  AND U10366 ( .A(n10771), .B(n10772), .Z(n10404) );
  NAND U10367 ( .A(n10773), .B(n10774), .Z(n10772) );
  NANDN U10368 ( .A(n10775), .B(n10776), .Z(n10771) );
  OR U10369 ( .A(n10773), .B(n10774), .Z(n10776) );
  ANDN U10370 ( .B(\stack[1][45] ), .A(n5494), .Z(n10403) );
  XNOR U10371 ( .A(n10409), .B(n10777), .Z(n10402) );
  XNOR U10372 ( .A(n10410), .B(n10411), .Z(n10777) );
  AND U10373 ( .A(n10778), .B(n10779), .Z(n10411) );
  NANDN U10374 ( .A(n10780), .B(n10781), .Z(n10779) );
  NANDN U10375 ( .A(n10782), .B(n10783), .Z(n10778) );
  NANDN U10376 ( .A(n10781), .B(n10780), .Z(n10783) );
  ANDN U10377 ( .B(\stack[1][46] ), .A(n5470), .Z(n10410) );
  XNOR U10378 ( .A(n10416), .B(n10784), .Z(n10409) );
  XNOR U10379 ( .A(n10417), .B(n10418), .Z(n10784) );
  AND U10380 ( .A(n10785), .B(n10786), .Z(n10418) );
  NAND U10381 ( .A(n10787), .B(n10788), .Z(n10786) );
  NANDN U10382 ( .A(n10789), .B(n10790), .Z(n10785) );
  OR U10383 ( .A(n10787), .B(n10788), .Z(n10790) );
  ANDN U10384 ( .B(\stack[1][47] ), .A(n5446), .Z(n10417) );
  XNOR U10385 ( .A(n10423), .B(n10791), .Z(n10416) );
  XNOR U10386 ( .A(n10424), .B(n10425), .Z(n10791) );
  AND U10387 ( .A(n10792), .B(n10793), .Z(n10425) );
  NANDN U10388 ( .A(n10794), .B(n10795), .Z(n10793) );
  NANDN U10389 ( .A(n10796), .B(n10797), .Z(n10792) );
  NANDN U10390 ( .A(n10795), .B(n10794), .Z(n10797) );
  ANDN U10391 ( .B(\stack[1][48] ), .A(n5422), .Z(n10424) );
  XNOR U10392 ( .A(n10430), .B(n10798), .Z(n10423) );
  XNOR U10393 ( .A(n10431), .B(n10432), .Z(n10798) );
  AND U10394 ( .A(n10799), .B(n10800), .Z(n10432) );
  NAND U10395 ( .A(n10801), .B(n10802), .Z(n10800) );
  NANDN U10396 ( .A(n10803), .B(n10804), .Z(n10799) );
  OR U10397 ( .A(n10801), .B(n10802), .Z(n10804) );
  ANDN U10398 ( .B(\stack[1][49] ), .A(n5398), .Z(n10431) );
  XNOR U10399 ( .A(n10437), .B(n10805), .Z(n10430) );
  XNOR U10400 ( .A(n10438), .B(n10439), .Z(n10805) );
  AND U10401 ( .A(n10806), .B(n10807), .Z(n10439) );
  NANDN U10402 ( .A(n10808), .B(n10809), .Z(n10807) );
  NANDN U10403 ( .A(n10810), .B(n10811), .Z(n10806) );
  NANDN U10404 ( .A(n10809), .B(n10808), .Z(n10811) );
  ANDN U10405 ( .B(\stack[1][50] ), .A(n5374), .Z(n10438) );
  XNOR U10406 ( .A(n10444), .B(n10812), .Z(n10437) );
  XNOR U10407 ( .A(n10445), .B(n10446), .Z(n10812) );
  AND U10408 ( .A(n10813), .B(n10814), .Z(n10446) );
  NAND U10409 ( .A(n10815), .B(n10816), .Z(n10814) );
  NANDN U10410 ( .A(n10817), .B(n10818), .Z(n10813) );
  OR U10411 ( .A(n10815), .B(n10816), .Z(n10818) );
  ANDN U10412 ( .B(\stack[1][51] ), .A(n5350), .Z(n10445) );
  XNOR U10413 ( .A(n10451), .B(n10819), .Z(n10444) );
  XNOR U10414 ( .A(n10452), .B(n10453), .Z(n10819) );
  AND U10415 ( .A(n10820), .B(n10821), .Z(n10453) );
  NANDN U10416 ( .A(n10822), .B(n10823), .Z(n10821) );
  NANDN U10417 ( .A(n10824), .B(n10825), .Z(n10820) );
  NANDN U10418 ( .A(n10823), .B(n10822), .Z(n10825) );
  ANDN U10419 ( .B(\stack[1][52] ), .A(n5326), .Z(n10452) );
  XNOR U10420 ( .A(n10458), .B(n10826), .Z(n10451) );
  XNOR U10421 ( .A(n10459), .B(n10460), .Z(n10826) );
  AND U10422 ( .A(n10827), .B(n10828), .Z(n10460) );
  NAND U10423 ( .A(n10829), .B(n10830), .Z(n10828) );
  NANDN U10424 ( .A(n10831), .B(n10832), .Z(n10827) );
  OR U10425 ( .A(n10829), .B(n10830), .Z(n10832) );
  ANDN U10426 ( .B(\stack[1][53] ), .A(n5302), .Z(n10459) );
  XNOR U10427 ( .A(n10465), .B(n10833), .Z(n10458) );
  XNOR U10428 ( .A(n10466), .B(n10467), .Z(n10833) );
  AND U10429 ( .A(n10834), .B(n10835), .Z(n10467) );
  NANDN U10430 ( .A(n10836), .B(n10837), .Z(n10835) );
  NANDN U10431 ( .A(n10838), .B(n10839), .Z(n10834) );
  NANDN U10432 ( .A(n10837), .B(n10836), .Z(n10839) );
  ANDN U10433 ( .B(\stack[1][54] ), .A(n5278), .Z(n10466) );
  XNOR U10434 ( .A(n10472), .B(n10840), .Z(n10465) );
  XNOR U10435 ( .A(n10473), .B(n10474), .Z(n10840) );
  AND U10436 ( .A(n10841), .B(n10842), .Z(n10474) );
  NAND U10437 ( .A(n10843), .B(n10844), .Z(n10842) );
  NANDN U10438 ( .A(n10845), .B(n10846), .Z(n10841) );
  OR U10439 ( .A(n10843), .B(n10844), .Z(n10846) );
  ANDN U10440 ( .B(\stack[1][55] ), .A(n5254), .Z(n10473) );
  XNOR U10441 ( .A(n10479), .B(n10847), .Z(n10472) );
  XNOR U10442 ( .A(n10480), .B(n10481), .Z(n10847) );
  AND U10443 ( .A(n10848), .B(n10849), .Z(n10481) );
  NAND U10444 ( .A(n10850), .B(n10851), .Z(n10849) );
  NAND U10445 ( .A(n10852), .B(n10853), .Z(n10848) );
  OR U10446 ( .A(n10850), .B(n10851), .Z(n10852) );
  ANDN U10447 ( .B(\stack[1][56] ), .A(n5230), .Z(n10480) );
  XNOR U10448 ( .A(n10486), .B(n10854), .Z(n10479) );
  XNOR U10449 ( .A(n10487), .B(n10489), .Z(n10854) );
  ANDN U10450 ( .B(n10855), .A(n10856), .Z(n10489) );
  ANDN U10451 ( .B(\stack[0][0] ), .A(n6564), .Z(n10855) );
  ANDN U10452 ( .B(\stack[1][57] ), .A(n5206), .Z(n10487) );
  XOR U10453 ( .A(n10492), .B(n10857), .Z(n10486) );
  NANDN U10454 ( .A(n5160), .B(\stack[1][59] ), .Z(n10857) );
  NANDN U10455 ( .A(n6564), .B(\stack[0][1] ), .Z(n10492) );
  ANDN U10456 ( .B(\stack[1][5] ), .A(n6454), .Z(n8984) );
  AND U10457 ( .A(n10858), .B(n10859), .Z(n8985) );
  NANDN U10458 ( .A(n8990), .B(n8992), .Z(n10859) );
  NANDN U10459 ( .A(n8993), .B(n10860), .Z(n10858) );
  NANDN U10460 ( .A(n8992), .B(n8990), .Z(n10860) );
  XOR U10461 ( .A(n10500), .B(n10861), .Z(n8990) );
  XNOR U10462 ( .A(n10501), .B(n10502), .Z(n10861) );
  AND U10463 ( .A(n10862), .B(n10863), .Z(n10502) );
  NAND U10464 ( .A(n10864), .B(n10865), .Z(n10863) );
  NANDN U10465 ( .A(n10866), .B(n10867), .Z(n10862) );
  OR U10466 ( .A(n10864), .B(n10865), .Z(n10867) );
  ANDN U10467 ( .B(\stack[0][52] ), .A(n5316), .Z(n10501) );
  XNOR U10468 ( .A(n10507), .B(n10868), .Z(n10500) );
  XNOR U10469 ( .A(n10508), .B(n10509), .Z(n10868) );
  AND U10470 ( .A(n10869), .B(n10870), .Z(n10509) );
  NANDN U10471 ( .A(n10871), .B(n10872), .Z(n10870) );
  NANDN U10472 ( .A(n10873), .B(n10874), .Z(n10869) );
  NANDN U10473 ( .A(n10872), .B(n10871), .Z(n10874) );
  ANDN U10474 ( .B(\stack[0][51] ), .A(n5340), .Z(n10508) );
  XNOR U10475 ( .A(n10514), .B(n10875), .Z(n10507) );
  XNOR U10476 ( .A(n10515), .B(n10516), .Z(n10875) );
  AND U10477 ( .A(n10876), .B(n10877), .Z(n10516) );
  NAND U10478 ( .A(n10878), .B(n10879), .Z(n10877) );
  NANDN U10479 ( .A(n10880), .B(n10881), .Z(n10876) );
  OR U10480 ( .A(n10878), .B(n10879), .Z(n10881) );
  ANDN U10481 ( .B(\stack[0][50] ), .A(n5364), .Z(n10515) );
  XNOR U10482 ( .A(n10521), .B(n10882), .Z(n10514) );
  XNOR U10483 ( .A(n10522), .B(n10523), .Z(n10882) );
  AND U10484 ( .A(n10883), .B(n10884), .Z(n10523) );
  NANDN U10485 ( .A(n10885), .B(n10886), .Z(n10884) );
  NANDN U10486 ( .A(n10887), .B(n10888), .Z(n10883) );
  NANDN U10487 ( .A(n10886), .B(n10885), .Z(n10888) );
  ANDN U10488 ( .B(\stack[0][49] ), .A(n5387), .Z(n10522) );
  XNOR U10489 ( .A(n10528), .B(n10889), .Z(n10521) );
  XNOR U10490 ( .A(n10529), .B(n10530), .Z(n10889) );
  AND U10491 ( .A(n10890), .B(n10891), .Z(n10530) );
  NAND U10492 ( .A(n10892), .B(n10893), .Z(n10891) );
  NANDN U10493 ( .A(n10894), .B(n10895), .Z(n10890) );
  OR U10494 ( .A(n10892), .B(n10893), .Z(n10895) );
  ANDN U10495 ( .B(\stack[1][10] ), .A(n6310), .Z(n10529) );
  XNOR U10496 ( .A(n10535), .B(n10896), .Z(n10528) );
  XNOR U10497 ( .A(n10536), .B(n10537), .Z(n10896) );
  AND U10498 ( .A(n10897), .B(n10898), .Z(n10537) );
  NANDN U10499 ( .A(n10899), .B(n10900), .Z(n10898) );
  NANDN U10500 ( .A(n10901), .B(n10902), .Z(n10897) );
  NANDN U10501 ( .A(n10900), .B(n10899), .Z(n10902) );
  ANDN U10502 ( .B(\stack[1][11] ), .A(n6286), .Z(n10536) );
  XNOR U10503 ( .A(n10542), .B(n10903), .Z(n10535) );
  XNOR U10504 ( .A(n10543), .B(n10544), .Z(n10903) );
  AND U10505 ( .A(n10904), .B(n10905), .Z(n10544) );
  NAND U10506 ( .A(n10906), .B(n10907), .Z(n10905) );
  NANDN U10507 ( .A(n10908), .B(n10909), .Z(n10904) );
  OR U10508 ( .A(n10906), .B(n10907), .Z(n10909) );
  ANDN U10509 ( .B(\stack[1][12] ), .A(n6262), .Z(n10543) );
  XNOR U10510 ( .A(n10549), .B(n10910), .Z(n10542) );
  XNOR U10511 ( .A(n10550), .B(n10551), .Z(n10910) );
  AND U10512 ( .A(n10911), .B(n10912), .Z(n10551) );
  NANDN U10513 ( .A(n10913), .B(n10914), .Z(n10912) );
  NANDN U10514 ( .A(n10915), .B(n10916), .Z(n10911) );
  NANDN U10515 ( .A(n10914), .B(n10913), .Z(n10916) );
  ANDN U10516 ( .B(\stack[1][13] ), .A(n6238), .Z(n10550) );
  XNOR U10517 ( .A(n10556), .B(n10917), .Z(n10549) );
  XNOR U10518 ( .A(n10557), .B(n10558), .Z(n10917) );
  AND U10519 ( .A(n10918), .B(n10919), .Z(n10558) );
  NAND U10520 ( .A(n10920), .B(n10921), .Z(n10919) );
  NANDN U10521 ( .A(n10922), .B(n10923), .Z(n10918) );
  OR U10522 ( .A(n10920), .B(n10921), .Z(n10923) );
  ANDN U10523 ( .B(\stack[1][14] ), .A(n6214), .Z(n10557) );
  XNOR U10524 ( .A(n10563), .B(n10924), .Z(n10556) );
  XNOR U10525 ( .A(n10564), .B(n10565), .Z(n10924) );
  AND U10526 ( .A(n10925), .B(n10926), .Z(n10565) );
  NANDN U10527 ( .A(n10927), .B(n10928), .Z(n10926) );
  NANDN U10528 ( .A(n10929), .B(n10930), .Z(n10925) );
  NANDN U10529 ( .A(n10928), .B(n10927), .Z(n10930) );
  ANDN U10530 ( .B(\stack[1][15] ), .A(n6190), .Z(n10564) );
  XNOR U10531 ( .A(n10570), .B(n10931), .Z(n10563) );
  XNOR U10532 ( .A(n10571), .B(n10572), .Z(n10931) );
  AND U10533 ( .A(n10932), .B(n10933), .Z(n10572) );
  NAND U10534 ( .A(n10934), .B(n10935), .Z(n10933) );
  NANDN U10535 ( .A(n10936), .B(n10937), .Z(n10932) );
  OR U10536 ( .A(n10934), .B(n10935), .Z(n10937) );
  ANDN U10537 ( .B(\stack[1][16] ), .A(n6166), .Z(n10571) );
  XNOR U10538 ( .A(n10577), .B(n10938), .Z(n10570) );
  XNOR U10539 ( .A(n10578), .B(n10579), .Z(n10938) );
  AND U10540 ( .A(n10939), .B(n10940), .Z(n10579) );
  NANDN U10541 ( .A(n10941), .B(n10942), .Z(n10940) );
  NANDN U10542 ( .A(n10943), .B(n10944), .Z(n10939) );
  NANDN U10543 ( .A(n10942), .B(n10941), .Z(n10944) );
  ANDN U10544 ( .B(\stack[1][17] ), .A(n6142), .Z(n10578) );
  XNOR U10545 ( .A(n10584), .B(n10945), .Z(n10577) );
  XNOR U10546 ( .A(n10585), .B(n10586), .Z(n10945) );
  AND U10547 ( .A(n10946), .B(n10947), .Z(n10586) );
  NAND U10548 ( .A(n10948), .B(n10949), .Z(n10947) );
  NANDN U10549 ( .A(n10950), .B(n10951), .Z(n10946) );
  OR U10550 ( .A(n10948), .B(n10949), .Z(n10951) );
  ANDN U10551 ( .B(\stack[1][18] ), .A(n6118), .Z(n10585) );
  XNOR U10552 ( .A(n10591), .B(n10952), .Z(n10584) );
  XNOR U10553 ( .A(n10592), .B(n10593), .Z(n10952) );
  AND U10554 ( .A(n10953), .B(n10954), .Z(n10593) );
  NANDN U10555 ( .A(n10955), .B(n10956), .Z(n10954) );
  NANDN U10556 ( .A(n10957), .B(n10958), .Z(n10953) );
  NANDN U10557 ( .A(n10956), .B(n10955), .Z(n10958) );
  ANDN U10558 ( .B(\stack[1][19] ), .A(n6094), .Z(n10592) );
  XNOR U10559 ( .A(n10598), .B(n10959), .Z(n10591) );
  XNOR U10560 ( .A(n10599), .B(n10600), .Z(n10959) );
  AND U10561 ( .A(n10960), .B(n10961), .Z(n10600) );
  NAND U10562 ( .A(n10962), .B(n10963), .Z(n10961) );
  NANDN U10563 ( .A(n10964), .B(n10965), .Z(n10960) );
  OR U10564 ( .A(n10962), .B(n10963), .Z(n10965) );
  ANDN U10565 ( .B(\stack[1][20] ), .A(n6070), .Z(n10599) );
  XNOR U10566 ( .A(n10605), .B(n10966), .Z(n10598) );
  XNOR U10567 ( .A(n10606), .B(n10607), .Z(n10966) );
  AND U10568 ( .A(n10967), .B(n10968), .Z(n10607) );
  NANDN U10569 ( .A(n10969), .B(n10970), .Z(n10968) );
  NANDN U10570 ( .A(n10971), .B(n10972), .Z(n10967) );
  NANDN U10571 ( .A(n10970), .B(n10969), .Z(n10972) );
  ANDN U10572 ( .B(\stack[1][21] ), .A(n6046), .Z(n10606) );
  XNOR U10573 ( .A(n10612), .B(n10973), .Z(n10605) );
  XNOR U10574 ( .A(n10613), .B(n10614), .Z(n10973) );
  AND U10575 ( .A(n10974), .B(n10975), .Z(n10614) );
  NAND U10576 ( .A(n10976), .B(n10977), .Z(n10975) );
  NANDN U10577 ( .A(n10978), .B(n10979), .Z(n10974) );
  OR U10578 ( .A(n10976), .B(n10977), .Z(n10979) );
  ANDN U10579 ( .B(\stack[1][22] ), .A(n6022), .Z(n10613) );
  XNOR U10580 ( .A(n10619), .B(n10980), .Z(n10612) );
  XNOR U10581 ( .A(n10620), .B(n10621), .Z(n10980) );
  AND U10582 ( .A(n10981), .B(n10982), .Z(n10621) );
  NANDN U10583 ( .A(n10983), .B(n10984), .Z(n10982) );
  NANDN U10584 ( .A(n10985), .B(n10986), .Z(n10981) );
  NANDN U10585 ( .A(n10984), .B(n10983), .Z(n10986) );
  ANDN U10586 ( .B(\stack[1][23] ), .A(n5998), .Z(n10620) );
  XNOR U10587 ( .A(n10626), .B(n10987), .Z(n10619) );
  XNOR U10588 ( .A(n10627), .B(n10628), .Z(n10987) );
  AND U10589 ( .A(n10988), .B(n10989), .Z(n10628) );
  NAND U10590 ( .A(n10990), .B(n10991), .Z(n10989) );
  NANDN U10591 ( .A(n10992), .B(n10993), .Z(n10988) );
  OR U10592 ( .A(n10990), .B(n10991), .Z(n10993) );
  ANDN U10593 ( .B(\stack[1][24] ), .A(n5974), .Z(n10627) );
  XNOR U10594 ( .A(n10633), .B(n10994), .Z(n10626) );
  XNOR U10595 ( .A(n10634), .B(n10635), .Z(n10994) );
  AND U10596 ( .A(n10995), .B(n10996), .Z(n10635) );
  NANDN U10597 ( .A(n10997), .B(n10998), .Z(n10996) );
  NANDN U10598 ( .A(n10999), .B(n11000), .Z(n10995) );
  NANDN U10599 ( .A(n10998), .B(n10997), .Z(n11000) );
  ANDN U10600 ( .B(\stack[1][25] ), .A(n5950), .Z(n10634) );
  XNOR U10601 ( .A(n10640), .B(n11001), .Z(n10633) );
  XNOR U10602 ( .A(n10641), .B(n10642), .Z(n11001) );
  AND U10603 ( .A(n11002), .B(n11003), .Z(n10642) );
  NAND U10604 ( .A(n11004), .B(n11005), .Z(n11003) );
  NANDN U10605 ( .A(n11006), .B(n11007), .Z(n11002) );
  OR U10606 ( .A(n11004), .B(n11005), .Z(n11007) );
  ANDN U10607 ( .B(\stack[1][26] ), .A(n5926), .Z(n10641) );
  XNOR U10608 ( .A(n10647), .B(n11008), .Z(n10640) );
  XNOR U10609 ( .A(n10648), .B(n10649), .Z(n11008) );
  AND U10610 ( .A(n11009), .B(n11010), .Z(n10649) );
  NANDN U10611 ( .A(n11011), .B(n11012), .Z(n11010) );
  NANDN U10612 ( .A(n11013), .B(n11014), .Z(n11009) );
  NANDN U10613 ( .A(n11012), .B(n11011), .Z(n11014) );
  ANDN U10614 ( .B(\stack[1][27] ), .A(n5902), .Z(n10648) );
  XNOR U10615 ( .A(n10654), .B(n11015), .Z(n10647) );
  XNOR U10616 ( .A(n10655), .B(n10656), .Z(n11015) );
  AND U10617 ( .A(n11016), .B(n11017), .Z(n10656) );
  NAND U10618 ( .A(n11018), .B(n11019), .Z(n11017) );
  NANDN U10619 ( .A(n11020), .B(n11021), .Z(n11016) );
  OR U10620 ( .A(n11018), .B(n11019), .Z(n11021) );
  ANDN U10621 ( .B(\stack[1][28] ), .A(n5878), .Z(n10655) );
  XNOR U10622 ( .A(n10661), .B(n11022), .Z(n10654) );
  XNOR U10623 ( .A(n10662), .B(n10663), .Z(n11022) );
  AND U10624 ( .A(n11023), .B(n11024), .Z(n10663) );
  NANDN U10625 ( .A(n11025), .B(n11026), .Z(n11024) );
  NANDN U10626 ( .A(n11027), .B(n11028), .Z(n11023) );
  NANDN U10627 ( .A(n11026), .B(n11025), .Z(n11028) );
  ANDN U10628 ( .B(\stack[1][29] ), .A(n5854), .Z(n10662) );
  XNOR U10629 ( .A(n10668), .B(n11029), .Z(n10661) );
  XNOR U10630 ( .A(n10669), .B(n10670), .Z(n11029) );
  AND U10631 ( .A(n11030), .B(n11031), .Z(n10670) );
  NAND U10632 ( .A(n11032), .B(n11033), .Z(n11031) );
  NANDN U10633 ( .A(n11034), .B(n11035), .Z(n11030) );
  OR U10634 ( .A(n11032), .B(n11033), .Z(n11035) );
  ANDN U10635 ( .B(\stack[1][30] ), .A(n5830), .Z(n10669) );
  XNOR U10636 ( .A(n10675), .B(n11036), .Z(n10668) );
  XNOR U10637 ( .A(n10676), .B(n10677), .Z(n11036) );
  AND U10638 ( .A(n11037), .B(n11038), .Z(n10677) );
  NANDN U10639 ( .A(n11039), .B(n11040), .Z(n11038) );
  NANDN U10640 ( .A(n11041), .B(n11042), .Z(n11037) );
  NANDN U10641 ( .A(n11040), .B(n11039), .Z(n11042) );
  ANDN U10642 ( .B(\stack[1][31] ), .A(n5806), .Z(n10676) );
  XNOR U10643 ( .A(n10682), .B(n11043), .Z(n10675) );
  XNOR U10644 ( .A(n10683), .B(n10684), .Z(n11043) );
  AND U10645 ( .A(n11044), .B(n11045), .Z(n10684) );
  NAND U10646 ( .A(n11046), .B(n11047), .Z(n11045) );
  NANDN U10647 ( .A(n11048), .B(n11049), .Z(n11044) );
  OR U10648 ( .A(n11046), .B(n11047), .Z(n11049) );
  ANDN U10649 ( .B(\stack[1][32] ), .A(n5782), .Z(n10683) );
  XNOR U10650 ( .A(n10689), .B(n11050), .Z(n10682) );
  XNOR U10651 ( .A(n10690), .B(n10691), .Z(n11050) );
  AND U10652 ( .A(n11051), .B(n11052), .Z(n10691) );
  NANDN U10653 ( .A(n11053), .B(n11054), .Z(n11052) );
  NANDN U10654 ( .A(n11055), .B(n11056), .Z(n11051) );
  NANDN U10655 ( .A(n11054), .B(n11053), .Z(n11056) );
  ANDN U10656 ( .B(\stack[1][33] ), .A(n5758), .Z(n10690) );
  XNOR U10657 ( .A(n10696), .B(n11057), .Z(n10689) );
  XNOR U10658 ( .A(n10697), .B(n10698), .Z(n11057) );
  AND U10659 ( .A(n11058), .B(n11059), .Z(n10698) );
  NAND U10660 ( .A(n11060), .B(n11061), .Z(n11059) );
  NANDN U10661 ( .A(n11062), .B(n11063), .Z(n11058) );
  OR U10662 ( .A(n11060), .B(n11061), .Z(n11063) );
  ANDN U10663 ( .B(\stack[1][34] ), .A(n5734), .Z(n10697) );
  XNOR U10664 ( .A(n10703), .B(n11064), .Z(n10696) );
  XNOR U10665 ( .A(n10704), .B(n10705), .Z(n11064) );
  AND U10666 ( .A(n11065), .B(n11066), .Z(n10705) );
  NANDN U10667 ( .A(n11067), .B(n11068), .Z(n11066) );
  NANDN U10668 ( .A(n11069), .B(n11070), .Z(n11065) );
  NANDN U10669 ( .A(n11068), .B(n11067), .Z(n11070) );
  ANDN U10670 ( .B(\stack[1][35] ), .A(n5710), .Z(n10704) );
  XNOR U10671 ( .A(n10710), .B(n11071), .Z(n10703) );
  XNOR U10672 ( .A(n10711), .B(n10712), .Z(n11071) );
  AND U10673 ( .A(n11072), .B(n11073), .Z(n10712) );
  NAND U10674 ( .A(n11074), .B(n11075), .Z(n11073) );
  NANDN U10675 ( .A(n11076), .B(n11077), .Z(n11072) );
  OR U10676 ( .A(n11074), .B(n11075), .Z(n11077) );
  ANDN U10677 ( .B(\stack[1][36] ), .A(n5686), .Z(n10711) );
  XNOR U10678 ( .A(n10718), .B(n11078), .Z(n10710) );
  XOR U10679 ( .A(n10719), .B(n10720), .Z(n11078) );
  NAND U10680 ( .A(n11079), .B(n11080), .Z(n10720) );
  NANDN U10681 ( .A(n11081), .B(n11082), .Z(n11080) );
  OR U10682 ( .A(n11083), .B(n11084), .Z(n11082) );
  AND U10683 ( .A(\stack[0][21] ), .B(\stack[1][37] ), .Z(n10719) );
  XNOR U10684 ( .A(n10725), .B(n11085), .Z(n10718) );
  XNOR U10685 ( .A(n10724), .B(n10727), .Z(n11085) );
  AND U10686 ( .A(\stack[0][20] ), .B(\stack[1][38] ), .Z(n10727) );
  AND U10687 ( .A(n11086), .B(n11087), .Z(n10724) );
  NAND U10688 ( .A(n11088), .B(n11089), .Z(n11087) );
  OR U10689 ( .A(n11090), .B(n11091), .Z(n11088) );
  XNOR U10690 ( .A(n10731), .B(n11092), .Z(n10725) );
  XNOR U10691 ( .A(n10732), .B(n10733), .Z(n11092) );
  AND U10692 ( .A(n11093), .B(n11094), .Z(n10733) );
  NANDN U10693 ( .A(n11095), .B(n11096), .Z(n11094) );
  NANDN U10694 ( .A(n11097), .B(n11098), .Z(n11093) );
  NANDN U10695 ( .A(n11096), .B(n11095), .Z(n11098) );
  ANDN U10696 ( .B(\stack[1][39] ), .A(n5614), .Z(n10732) );
  XNOR U10697 ( .A(n10738), .B(n11099), .Z(n10731) );
  XNOR U10698 ( .A(n10739), .B(n10740), .Z(n11099) );
  AND U10699 ( .A(n11100), .B(n11101), .Z(n10740) );
  NAND U10700 ( .A(n11102), .B(n11103), .Z(n11101) );
  NANDN U10701 ( .A(n11104), .B(n11105), .Z(n11100) );
  OR U10702 ( .A(n11102), .B(n11103), .Z(n11105) );
  ANDN U10703 ( .B(\stack[1][40] ), .A(n5590), .Z(n10739) );
  XNOR U10704 ( .A(n10745), .B(n11106), .Z(n10738) );
  XNOR U10705 ( .A(n10746), .B(n10747), .Z(n11106) );
  AND U10706 ( .A(n11107), .B(n11108), .Z(n10747) );
  NANDN U10707 ( .A(n11109), .B(n11110), .Z(n11108) );
  NANDN U10708 ( .A(n11111), .B(n11112), .Z(n11107) );
  NANDN U10709 ( .A(n11110), .B(n11109), .Z(n11112) );
  ANDN U10710 ( .B(\stack[1][41] ), .A(n5566), .Z(n10746) );
  XNOR U10711 ( .A(n10752), .B(n11113), .Z(n10745) );
  XNOR U10712 ( .A(n10753), .B(n10754), .Z(n11113) );
  AND U10713 ( .A(n11114), .B(n11115), .Z(n10754) );
  NAND U10714 ( .A(n11116), .B(n11117), .Z(n11115) );
  NANDN U10715 ( .A(n11118), .B(n11119), .Z(n11114) );
  OR U10716 ( .A(n11116), .B(n11117), .Z(n11119) );
  ANDN U10717 ( .B(\stack[1][42] ), .A(n5542), .Z(n10753) );
  XNOR U10718 ( .A(n10759), .B(n11120), .Z(n10752) );
  XNOR U10719 ( .A(n10760), .B(n10761), .Z(n11120) );
  AND U10720 ( .A(n11121), .B(n11122), .Z(n10761) );
  NANDN U10721 ( .A(n11123), .B(n11124), .Z(n11122) );
  NANDN U10722 ( .A(n11125), .B(n11126), .Z(n11121) );
  NANDN U10723 ( .A(n11124), .B(n11123), .Z(n11126) );
  ANDN U10724 ( .B(\stack[1][43] ), .A(n5518), .Z(n10760) );
  XNOR U10725 ( .A(n10766), .B(n11127), .Z(n10759) );
  XNOR U10726 ( .A(n10767), .B(n10768), .Z(n11127) );
  AND U10727 ( .A(n11128), .B(n11129), .Z(n10768) );
  NAND U10728 ( .A(n11130), .B(n11131), .Z(n11129) );
  NANDN U10729 ( .A(n11132), .B(n11133), .Z(n11128) );
  OR U10730 ( .A(n11130), .B(n11131), .Z(n11133) );
  ANDN U10731 ( .B(\stack[1][44] ), .A(n5494), .Z(n10767) );
  XNOR U10732 ( .A(n10773), .B(n11134), .Z(n10766) );
  XNOR U10733 ( .A(n10774), .B(n10775), .Z(n11134) );
  AND U10734 ( .A(n11135), .B(n11136), .Z(n10775) );
  NANDN U10735 ( .A(n11137), .B(n11138), .Z(n11136) );
  NANDN U10736 ( .A(n11139), .B(n11140), .Z(n11135) );
  NANDN U10737 ( .A(n11138), .B(n11137), .Z(n11140) );
  ANDN U10738 ( .B(\stack[1][45] ), .A(n5470), .Z(n10774) );
  XNOR U10739 ( .A(n10780), .B(n11141), .Z(n10773) );
  XNOR U10740 ( .A(n10781), .B(n10782), .Z(n11141) );
  AND U10741 ( .A(n11142), .B(n11143), .Z(n10782) );
  NAND U10742 ( .A(n11144), .B(n11145), .Z(n11143) );
  NANDN U10743 ( .A(n11146), .B(n11147), .Z(n11142) );
  OR U10744 ( .A(n11144), .B(n11145), .Z(n11147) );
  ANDN U10745 ( .B(\stack[1][46] ), .A(n5446), .Z(n10781) );
  XNOR U10746 ( .A(n10787), .B(n11148), .Z(n10780) );
  XNOR U10747 ( .A(n10788), .B(n10789), .Z(n11148) );
  AND U10748 ( .A(n11149), .B(n11150), .Z(n10789) );
  NANDN U10749 ( .A(n11151), .B(n11152), .Z(n11150) );
  NANDN U10750 ( .A(n11153), .B(n11154), .Z(n11149) );
  NANDN U10751 ( .A(n11152), .B(n11151), .Z(n11154) );
  ANDN U10752 ( .B(\stack[1][47] ), .A(n5422), .Z(n10788) );
  XNOR U10753 ( .A(n10794), .B(n11155), .Z(n10787) );
  XNOR U10754 ( .A(n10795), .B(n10796), .Z(n11155) );
  AND U10755 ( .A(n11156), .B(n11157), .Z(n10796) );
  NAND U10756 ( .A(n11158), .B(n11159), .Z(n11157) );
  NANDN U10757 ( .A(n11160), .B(n11161), .Z(n11156) );
  OR U10758 ( .A(n11158), .B(n11159), .Z(n11161) );
  ANDN U10759 ( .B(\stack[1][48] ), .A(n5398), .Z(n10795) );
  XNOR U10760 ( .A(n10801), .B(n11162), .Z(n10794) );
  XNOR U10761 ( .A(n10802), .B(n10803), .Z(n11162) );
  AND U10762 ( .A(n11163), .B(n11164), .Z(n10803) );
  NANDN U10763 ( .A(n11165), .B(n11166), .Z(n11164) );
  NANDN U10764 ( .A(n11167), .B(n11168), .Z(n11163) );
  NANDN U10765 ( .A(n11166), .B(n11165), .Z(n11168) );
  ANDN U10766 ( .B(\stack[1][49] ), .A(n5374), .Z(n10802) );
  XNOR U10767 ( .A(n10808), .B(n11169), .Z(n10801) );
  XNOR U10768 ( .A(n10809), .B(n10810), .Z(n11169) );
  AND U10769 ( .A(n11170), .B(n11171), .Z(n10810) );
  NAND U10770 ( .A(n11172), .B(n11173), .Z(n11171) );
  NANDN U10771 ( .A(n11174), .B(n11175), .Z(n11170) );
  OR U10772 ( .A(n11172), .B(n11173), .Z(n11175) );
  ANDN U10773 ( .B(\stack[1][50] ), .A(n5350), .Z(n10809) );
  XNOR U10774 ( .A(n10815), .B(n11176), .Z(n10808) );
  XNOR U10775 ( .A(n10816), .B(n10817), .Z(n11176) );
  AND U10776 ( .A(n11177), .B(n11178), .Z(n10817) );
  NANDN U10777 ( .A(n11179), .B(n11180), .Z(n11178) );
  NANDN U10778 ( .A(n11181), .B(n11182), .Z(n11177) );
  NANDN U10779 ( .A(n11180), .B(n11179), .Z(n11182) );
  ANDN U10780 ( .B(\stack[1][51] ), .A(n5326), .Z(n10816) );
  XNOR U10781 ( .A(n10822), .B(n11183), .Z(n10815) );
  XNOR U10782 ( .A(n10823), .B(n10824), .Z(n11183) );
  AND U10783 ( .A(n11184), .B(n11185), .Z(n10824) );
  NAND U10784 ( .A(n11186), .B(n11187), .Z(n11185) );
  NANDN U10785 ( .A(n11188), .B(n11189), .Z(n11184) );
  OR U10786 ( .A(n11186), .B(n11187), .Z(n11189) );
  ANDN U10787 ( .B(\stack[1][52] ), .A(n5302), .Z(n10823) );
  XNOR U10788 ( .A(n10829), .B(n11190), .Z(n10822) );
  XNOR U10789 ( .A(n10830), .B(n10831), .Z(n11190) );
  AND U10790 ( .A(n11191), .B(n11192), .Z(n10831) );
  NANDN U10791 ( .A(n11193), .B(n11194), .Z(n11192) );
  NANDN U10792 ( .A(n11195), .B(n11196), .Z(n11191) );
  NANDN U10793 ( .A(n11194), .B(n11193), .Z(n11196) );
  ANDN U10794 ( .B(\stack[1][53] ), .A(n5278), .Z(n10830) );
  XNOR U10795 ( .A(n10836), .B(n11197), .Z(n10829) );
  XNOR U10796 ( .A(n10837), .B(n10838), .Z(n11197) );
  AND U10797 ( .A(n11198), .B(n11199), .Z(n10838) );
  NAND U10798 ( .A(n11200), .B(n11201), .Z(n11199) );
  NANDN U10799 ( .A(n11202), .B(n11203), .Z(n11198) );
  OR U10800 ( .A(n11200), .B(n11201), .Z(n11203) );
  ANDN U10801 ( .B(\stack[1][54] ), .A(n5254), .Z(n10837) );
  XNOR U10802 ( .A(n10843), .B(n11204), .Z(n10836) );
  XNOR U10803 ( .A(n10844), .B(n10845), .Z(n11204) );
  AND U10804 ( .A(n11205), .B(n11206), .Z(n10845) );
  NAND U10805 ( .A(n11207), .B(n11208), .Z(n11206) );
  NAND U10806 ( .A(n11209), .B(n11210), .Z(n11205) );
  OR U10807 ( .A(n11207), .B(n11208), .Z(n11209) );
  ANDN U10808 ( .B(\stack[1][55] ), .A(n5230), .Z(n10844) );
  XNOR U10809 ( .A(n10850), .B(n11211), .Z(n10843) );
  XNOR U10810 ( .A(n10851), .B(n10853), .Z(n11211) );
  ANDN U10811 ( .B(n11212), .A(n11213), .Z(n10853) );
  ANDN U10812 ( .B(\stack[0][0] ), .A(n6540), .Z(n11212) );
  ANDN U10813 ( .B(\stack[1][56] ), .A(n5206), .Z(n10851) );
  XOR U10814 ( .A(n10856), .B(n11214), .Z(n10850) );
  NANDN U10815 ( .A(n5160), .B(\stack[1][58] ), .Z(n11214) );
  NANDN U10816 ( .A(n6540), .B(\stack[0][1] ), .Z(n10856) );
  ANDN U10817 ( .B(\stack[0][53] ), .A(n5292), .Z(n8992) );
  AND U10818 ( .A(n11215), .B(n11216), .Z(n8993) );
  NANDN U10819 ( .A(n9000), .B(n11217), .Z(n11215) );
  NANDN U10820 ( .A(n8999), .B(n8997), .Z(n11217) );
  XNOR U10821 ( .A(n10864), .B(n11218), .Z(n8997) );
  XNOR U10822 ( .A(n10865), .B(n10866), .Z(n11218) );
  AND U10823 ( .A(n11219), .B(n11220), .Z(n10866) );
  NANDN U10824 ( .A(n11221), .B(n11222), .Z(n11220) );
  NANDN U10825 ( .A(n11223), .B(n11224), .Z(n11219) );
  NANDN U10826 ( .A(n11222), .B(n11221), .Z(n11224) );
  ANDN U10827 ( .B(\stack[0][51] ), .A(n5316), .Z(n10865) );
  XNOR U10828 ( .A(n10871), .B(n11225), .Z(n10864) );
  XNOR U10829 ( .A(n10872), .B(n10873), .Z(n11225) );
  AND U10830 ( .A(n11226), .B(n11227), .Z(n10873) );
  NAND U10831 ( .A(n11228), .B(n11229), .Z(n11227) );
  NANDN U10832 ( .A(n11230), .B(n11231), .Z(n11226) );
  OR U10833 ( .A(n11228), .B(n11229), .Z(n11231) );
  ANDN U10834 ( .B(\stack[0][50] ), .A(n5340), .Z(n10872) );
  XNOR U10835 ( .A(n10878), .B(n11232), .Z(n10871) );
  XNOR U10836 ( .A(n10879), .B(n10880), .Z(n11232) );
  AND U10837 ( .A(n11233), .B(n11234), .Z(n10880) );
  NANDN U10838 ( .A(n11235), .B(n11236), .Z(n11234) );
  NANDN U10839 ( .A(n11237), .B(n11238), .Z(n11233) );
  NANDN U10840 ( .A(n11236), .B(n11235), .Z(n11238) );
  ANDN U10841 ( .B(\stack[0][49] ), .A(n5364), .Z(n10879) );
  XNOR U10842 ( .A(n10885), .B(n11239), .Z(n10878) );
  XNOR U10843 ( .A(n10886), .B(n10887), .Z(n11239) );
  AND U10844 ( .A(n11240), .B(n11241), .Z(n10887) );
  NAND U10845 ( .A(n11242), .B(n11243), .Z(n11241) );
  NANDN U10846 ( .A(n11244), .B(n11245), .Z(n11240) );
  OR U10847 ( .A(n11242), .B(n11243), .Z(n11245) );
  ANDN U10848 ( .B(\stack[0][48] ), .A(n5387), .Z(n10886) );
  XNOR U10849 ( .A(n10892), .B(n11246), .Z(n10885) );
  XNOR U10850 ( .A(n10893), .B(n10894), .Z(n11246) );
  AND U10851 ( .A(n11247), .B(n11248), .Z(n10894) );
  NANDN U10852 ( .A(n11249), .B(n11250), .Z(n11248) );
  NANDN U10853 ( .A(n11251), .B(n11252), .Z(n11247) );
  NANDN U10854 ( .A(n11250), .B(n11249), .Z(n11252) );
  ANDN U10855 ( .B(\stack[1][10] ), .A(n6286), .Z(n10893) );
  XNOR U10856 ( .A(n10899), .B(n11253), .Z(n10892) );
  XNOR U10857 ( .A(n10900), .B(n10901), .Z(n11253) );
  AND U10858 ( .A(n11254), .B(n11255), .Z(n10901) );
  NAND U10859 ( .A(n11256), .B(n11257), .Z(n11255) );
  NANDN U10860 ( .A(n11258), .B(n11259), .Z(n11254) );
  OR U10861 ( .A(n11256), .B(n11257), .Z(n11259) );
  ANDN U10862 ( .B(\stack[1][11] ), .A(n6262), .Z(n10900) );
  XNOR U10863 ( .A(n10906), .B(n11260), .Z(n10899) );
  XNOR U10864 ( .A(n10907), .B(n10908), .Z(n11260) );
  AND U10865 ( .A(n11261), .B(n11262), .Z(n10908) );
  NANDN U10866 ( .A(n11263), .B(n11264), .Z(n11262) );
  NANDN U10867 ( .A(n11265), .B(n11266), .Z(n11261) );
  NANDN U10868 ( .A(n11264), .B(n11263), .Z(n11266) );
  ANDN U10869 ( .B(\stack[1][12] ), .A(n6238), .Z(n10907) );
  XNOR U10870 ( .A(n10913), .B(n11267), .Z(n10906) );
  XNOR U10871 ( .A(n10914), .B(n10915), .Z(n11267) );
  AND U10872 ( .A(n11268), .B(n11269), .Z(n10915) );
  NAND U10873 ( .A(n11270), .B(n11271), .Z(n11269) );
  NANDN U10874 ( .A(n11272), .B(n11273), .Z(n11268) );
  OR U10875 ( .A(n11270), .B(n11271), .Z(n11273) );
  ANDN U10876 ( .B(\stack[1][13] ), .A(n6214), .Z(n10914) );
  XNOR U10877 ( .A(n10920), .B(n11274), .Z(n10913) );
  XNOR U10878 ( .A(n10921), .B(n10922), .Z(n11274) );
  AND U10879 ( .A(n11275), .B(n11276), .Z(n10922) );
  NANDN U10880 ( .A(n11277), .B(n11278), .Z(n11276) );
  NANDN U10881 ( .A(n11279), .B(n11280), .Z(n11275) );
  NANDN U10882 ( .A(n11278), .B(n11277), .Z(n11280) );
  ANDN U10883 ( .B(\stack[1][14] ), .A(n6190), .Z(n10921) );
  XNOR U10884 ( .A(n10927), .B(n11281), .Z(n10920) );
  XNOR U10885 ( .A(n10928), .B(n10929), .Z(n11281) );
  AND U10886 ( .A(n11282), .B(n11283), .Z(n10929) );
  NAND U10887 ( .A(n11284), .B(n11285), .Z(n11283) );
  NANDN U10888 ( .A(n11286), .B(n11287), .Z(n11282) );
  OR U10889 ( .A(n11284), .B(n11285), .Z(n11287) );
  ANDN U10890 ( .B(\stack[1][15] ), .A(n6166), .Z(n10928) );
  XNOR U10891 ( .A(n10934), .B(n11288), .Z(n10927) );
  XNOR U10892 ( .A(n10935), .B(n10936), .Z(n11288) );
  AND U10893 ( .A(n11289), .B(n11290), .Z(n10936) );
  NANDN U10894 ( .A(n11291), .B(n11292), .Z(n11290) );
  NANDN U10895 ( .A(n11293), .B(n11294), .Z(n11289) );
  NANDN U10896 ( .A(n11292), .B(n11291), .Z(n11294) );
  ANDN U10897 ( .B(\stack[1][16] ), .A(n6142), .Z(n10935) );
  XNOR U10898 ( .A(n10941), .B(n11295), .Z(n10934) );
  XNOR U10899 ( .A(n10942), .B(n10943), .Z(n11295) );
  AND U10900 ( .A(n11296), .B(n11297), .Z(n10943) );
  NAND U10901 ( .A(n11298), .B(n11299), .Z(n11297) );
  NANDN U10902 ( .A(n11300), .B(n11301), .Z(n11296) );
  OR U10903 ( .A(n11298), .B(n11299), .Z(n11301) );
  ANDN U10904 ( .B(\stack[1][17] ), .A(n6118), .Z(n10942) );
  XNOR U10905 ( .A(n10948), .B(n11302), .Z(n10941) );
  XNOR U10906 ( .A(n10949), .B(n10950), .Z(n11302) );
  AND U10907 ( .A(n11303), .B(n11304), .Z(n10950) );
  NANDN U10908 ( .A(n11305), .B(n11306), .Z(n11304) );
  NANDN U10909 ( .A(n11307), .B(n11308), .Z(n11303) );
  NANDN U10910 ( .A(n11306), .B(n11305), .Z(n11308) );
  ANDN U10911 ( .B(\stack[1][18] ), .A(n6094), .Z(n10949) );
  XNOR U10912 ( .A(n10955), .B(n11309), .Z(n10948) );
  XNOR U10913 ( .A(n10956), .B(n10957), .Z(n11309) );
  AND U10914 ( .A(n11310), .B(n11311), .Z(n10957) );
  NAND U10915 ( .A(n11312), .B(n11313), .Z(n11311) );
  NANDN U10916 ( .A(n11314), .B(n11315), .Z(n11310) );
  OR U10917 ( .A(n11312), .B(n11313), .Z(n11315) );
  ANDN U10918 ( .B(\stack[1][19] ), .A(n6070), .Z(n10956) );
  XNOR U10919 ( .A(n10962), .B(n11316), .Z(n10955) );
  XNOR U10920 ( .A(n10963), .B(n10964), .Z(n11316) );
  AND U10921 ( .A(n11317), .B(n11318), .Z(n10964) );
  NANDN U10922 ( .A(n11319), .B(n11320), .Z(n11318) );
  NANDN U10923 ( .A(n11321), .B(n11322), .Z(n11317) );
  NANDN U10924 ( .A(n11320), .B(n11319), .Z(n11322) );
  ANDN U10925 ( .B(\stack[1][20] ), .A(n6046), .Z(n10963) );
  XNOR U10926 ( .A(n10969), .B(n11323), .Z(n10962) );
  XNOR U10927 ( .A(n10970), .B(n10971), .Z(n11323) );
  AND U10928 ( .A(n11324), .B(n11325), .Z(n10971) );
  NAND U10929 ( .A(n11326), .B(n11327), .Z(n11325) );
  NANDN U10930 ( .A(n11328), .B(n11329), .Z(n11324) );
  OR U10931 ( .A(n11326), .B(n11327), .Z(n11329) );
  ANDN U10932 ( .B(\stack[1][21] ), .A(n6022), .Z(n10970) );
  XNOR U10933 ( .A(n10976), .B(n11330), .Z(n10969) );
  XNOR U10934 ( .A(n10977), .B(n10978), .Z(n11330) );
  AND U10935 ( .A(n11331), .B(n11332), .Z(n10978) );
  NANDN U10936 ( .A(n11333), .B(n11334), .Z(n11332) );
  NANDN U10937 ( .A(n11335), .B(n11336), .Z(n11331) );
  NANDN U10938 ( .A(n11334), .B(n11333), .Z(n11336) );
  ANDN U10939 ( .B(\stack[1][22] ), .A(n5998), .Z(n10977) );
  XNOR U10940 ( .A(n10983), .B(n11337), .Z(n10976) );
  XNOR U10941 ( .A(n10984), .B(n10985), .Z(n11337) );
  AND U10942 ( .A(n11338), .B(n11339), .Z(n10985) );
  NAND U10943 ( .A(n11340), .B(n11341), .Z(n11339) );
  NANDN U10944 ( .A(n11342), .B(n11343), .Z(n11338) );
  OR U10945 ( .A(n11340), .B(n11341), .Z(n11343) );
  ANDN U10946 ( .B(\stack[1][23] ), .A(n5974), .Z(n10984) );
  XNOR U10947 ( .A(n10990), .B(n11344), .Z(n10983) );
  XNOR U10948 ( .A(n10991), .B(n10992), .Z(n11344) );
  AND U10949 ( .A(n11345), .B(n11346), .Z(n10992) );
  NANDN U10950 ( .A(n11347), .B(n11348), .Z(n11346) );
  NANDN U10951 ( .A(n11349), .B(n11350), .Z(n11345) );
  NANDN U10952 ( .A(n11348), .B(n11347), .Z(n11350) );
  ANDN U10953 ( .B(\stack[1][24] ), .A(n5950), .Z(n10991) );
  XNOR U10954 ( .A(n10997), .B(n11351), .Z(n10990) );
  XNOR U10955 ( .A(n10998), .B(n10999), .Z(n11351) );
  AND U10956 ( .A(n11352), .B(n11353), .Z(n10999) );
  NAND U10957 ( .A(n11354), .B(n11355), .Z(n11353) );
  NANDN U10958 ( .A(n11356), .B(n11357), .Z(n11352) );
  OR U10959 ( .A(n11354), .B(n11355), .Z(n11357) );
  ANDN U10960 ( .B(\stack[1][25] ), .A(n5926), .Z(n10998) );
  XNOR U10961 ( .A(n11004), .B(n11358), .Z(n10997) );
  XNOR U10962 ( .A(n11005), .B(n11006), .Z(n11358) );
  AND U10963 ( .A(n11359), .B(n11360), .Z(n11006) );
  NANDN U10964 ( .A(n11361), .B(n11362), .Z(n11360) );
  NANDN U10965 ( .A(n11363), .B(n11364), .Z(n11359) );
  NANDN U10966 ( .A(n11362), .B(n11361), .Z(n11364) );
  ANDN U10967 ( .B(\stack[1][26] ), .A(n5902), .Z(n11005) );
  XNOR U10968 ( .A(n11011), .B(n11365), .Z(n11004) );
  XNOR U10969 ( .A(n11012), .B(n11013), .Z(n11365) );
  AND U10970 ( .A(n11366), .B(n11367), .Z(n11013) );
  NAND U10971 ( .A(n11368), .B(n11369), .Z(n11367) );
  NANDN U10972 ( .A(n11370), .B(n11371), .Z(n11366) );
  OR U10973 ( .A(n11368), .B(n11369), .Z(n11371) );
  ANDN U10974 ( .B(\stack[1][27] ), .A(n5878), .Z(n11012) );
  XNOR U10975 ( .A(n11018), .B(n11372), .Z(n11011) );
  XNOR U10976 ( .A(n11019), .B(n11020), .Z(n11372) );
  AND U10977 ( .A(n11373), .B(n11374), .Z(n11020) );
  NANDN U10978 ( .A(n11375), .B(n11376), .Z(n11374) );
  NANDN U10979 ( .A(n11377), .B(n11378), .Z(n11373) );
  NANDN U10980 ( .A(n11376), .B(n11375), .Z(n11378) );
  ANDN U10981 ( .B(\stack[1][28] ), .A(n5854), .Z(n11019) );
  XNOR U10982 ( .A(n11025), .B(n11379), .Z(n11018) );
  XNOR U10983 ( .A(n11026), .B(n11027), .Z(n11379) );
  AND U10984 ( .A(n11380), .B(n11381), .Z(n11027) );
  NAND U10985 ( .A(n11382), .B(n11383), .Z(n11381) );
  NANDN U10986 ( .A(n11384), .B(n11385), .Z(n11380) );
  OR U10987 ( .A(n11382), .B(n11383), .Z(n11385) );
  ANDN U10988 ( .B(\stack[1][29] ), .A(n5830), .Z(n11026) );
  XNOR U10989 ( .A(n11032), .B(n11386), .Z(n11025) );
  XNOR U10990 ( .A(n11033), .B(n11034), .Z(n11386) );
  AND U10991 ( .A(n11387), .B(n11388), .Z(n11034) );
  NANDN U10992 ( .A(n11389), .B(n11390), .Z(n11388) );
  NANDN U10993 ( .A(n11391), .B(n11392), .Z(n11387) );
  NANDN U10994 ( .A(n11390), .B(n11389), .Z(n11392) );
  ANDN U10995 ( .B(\stack[1][30] ), .A(n5806), .Z(n11033) );
  XNOR U10996 ( .A(n11039), .B(n11393), .Z(n11032) );
  XNOR U10997 ( .A(n11040), .B(n11041), .Z(n11393) );
  AND U10998 ( .A(n11394), .B(n11395), .Z(n11041) );
  NAND U10999 ( .A(n11396), .B(n11397), .Z(n11395) );
  NANDN U11000 ( .A(n11398), .B(n11399), .Z(n11394) );
  OR U11001 ( .A(n11396), .B(n11397), .Z(n11399) );
  ANDN U11002 ( .B(\stack[1][31] ), .A(n5782), .Z(n11040) );
  XNOR U11003 ( .A(n11046), .B(n11400), .Z(n11039) );
  XNOR U11004 ( .A(n11047), .B(n11048), .Z(n11400) );
  AND U11005 ( .A(n11401), .B(n11402), .Z(n11048) );
  NANDN U11006 ( .A(n11403), .B(n11404), .Z(n11402) );
  NANDN U11007 ( .A(n11405), .B(n11406), .Z(n11401) );
  NANDN U11008 ( .A(n11404), .B(n11403), .Z(n11406) );
  ANDN U11009 ( .B(\stack[1][32] ), .A(n5758), .Z(n11047) );
  XNOR U11010 ( .A(n11053), .B(n11407), .Z(n11046) );
  XNOR U11011 ( .A(n11054), .B(n11055), .Z(n11407) );
  AND U11012 ( .A(n11408), .B(n11409), .Z(n11055) );
  NAND U11013 ( .A(n11410), .B(n11411), .Z(n11409) );
  NANDN U11014 ( .A(n11412), .B(n11413), .Z(n11408) );
  OR U11015 ( .A(n11410), .B(n11411), .Z(n11413) );
  ANDN U11016 ( .B(\stack[1][33] ), .A(n5734), .Z(n11054) );
  XNOR U11017 ( .A(n11060), .B(n11414), .Z(n11053) );
  XNOR U11018 ( .A(n11061), .B(n11062), .Z(n11414) );
  AND U11019 ( .A(n11415), .B(n11416), .Z(n11062) );
  NANDN U11020 ( .A(n11417), .B(n11418), .Z(n11416) );
  NANDN U11021 ( .A(n11419), .B(n11420), .Z(n11415) );
  NANDN U11022 ( .A(n11418), .B(n11417), .Z(n11420) );
  ANDN U11023 ( .B(\stack[1][34] ), .A(n5710), .Z(n11061) );
  XNOR U11024 ( .A(n11067), .B(n11421), .Z(n11060) );
  XNOR U11025 ( .A(n11068), .B(n11069), .Z(n11421) );
  AND U11026 ( .A(n11422), .B(n11423), .Z(n11069) );
  NAND U11027 ( .A(n11424), .B(n11425), .Z(n11423) );
  NANDN U11028 ( .A(n11426), .B(n11427), .Z(n11422) );
  OR U11029 ( .A(n11424), .B(n11425), .Z(n11427) );
  ANDN U11030 ( .B(\stack[1][35] ), .A(n5686), .Z(n11068) );
  XNOR U11031 ( .A(n11074), .B(n11428), .Z(n11067) );
  XNOR U11032 ( .A(n11075), .B(n11076), .Z(n11428) );
  AND U11033 ( .A(n11429), .B(n11430), .Z(n11076) );
  NANDN U11034 ( .A(n11431), .B(n11432), .Z(n11430) );
  NANDN U11035 ( .A(n11433), .B(n11434), .Z(n11429) );
  NANDN U11036 ( .A(n11432), .B(n11431), .Z(n11434) );
  ANDN U11037 ( .B(\stack[1][36] ), .A(n5662), .Z(n11075) );
  XNOR U11038 ( .A(n11081), .B(n11435), .Z(n11074) );
  XOR U11039 ( .A(n11083), .B(n11084), .Z(n11435) );
  NAND U11040 ( .A(n11436), .B(n11437), .Z(n11084) );
  NAND U11041 ( .A(n11438), .B(n11439), .Z(n11437) );
  OR U11042 ( .A(n11440), .B(n11441), .Z(n11438) );
  AND U11043 ( .A(\stack[0][20] ), .B(\stack[1][37] ), .Z(n11083) );
  XNOR U11044 ( .A(n11090), .B(n11442), .Z(n11081) );
  XOR U11045 ( .A(n11091), .B(n11089), .Z(n11442) );
  AND U11046 ( .A(\stack[0][19] ), .B(\stack[1][38] ), .Z(n11089) );
  NAND U11047 ( .A(n11443), .B(n11444), .Z(n11091) );
  OR U11048 ( .A(n11445), .B(n11446), .Z(n11444) );
  NAND U11049 ( .A(n11447), .B(n11448), .Z(n11443) );
  NAND U11050 ( .A(n11446), .B(n11445), .Z(n11447) );
  XNOR U11051 ( .A(n11095), .B(n11449), .Z(n11090) );
  XNOR U11052 ( .A(n11096), .B(n11097), .Z(n11449) );
  AND U11053 ( .A(n11450), .B(n11451), .Z(n11097) );
  NAND U11054 ( .A(n11452), .B(n11453), .Z(n11451) );
  NANDN U11055 ( .A(n11454), .B(n11455), .Z(n11450) );
  OR U11056 ( .A(n11452), .B(n11453), .Z(n11455) );
  ANDN U11057 ( .B(\stack[1][39] ), .A(n5590), .Z(n11096) );
  XNOR U11058 ( .A(n11102), .B(n11456), .Z(n11095) );
  XNOR U11059 ( .A(n11103), .B(n11104), .Z(n11456) );
  AND U11060 ( .A(n11457), .B(n11458), .Z(n11104) );
  NANDN U11061 ( .A(n11459), .B(n11460), .Z(n11458) );
  NANDN U11062 ( .A(n11461), .B(n11462), .Z(n11457) );
  NANDN U11063 ( .A(n11460), .B(n11459), .Z(n11462) );
  ANDN U11064 ( .B(\stack[1][40] ), .A(n5566), .Z(n11103) );
  XNOR U11065 ( .A(n11109), .B(n11463), .Z(n11102) );
  XNOR U11066 ( .A(n11110), .B(n11111), .Z(n11463) );
  AND U11067 ( .A(n11464), .B(n11465), .Z(n11111) );
  NAND U11068 ( .A(n11466), .B(n11467), .Z(n11465) );
  NANDN U11069 ( .A(n11468), .B(n11469), .Z(n11464) );
  OR U11070 ( .A(n11466), .B(n11467), .Z(n11469) );
  ANDN U11071 ( .B(\stack[1][41] ), .A(n5542), .Z(n11110) );
  XNOR U11072 ( .A(n11116), .B(n11470), .Z(n11109) );
  XNOR U11073 ( .A(n11117), .B(n11118), .Z(n11470) );
  AND U11074 ( .A(n11471), .B(n11472), .Z(n11118) );
  NANDN U11075 ( .A(n11473), .B(n11474), .Z(n11472) );
  NANDN U11076 ( .A(n11475), .B(n11476), .Z(n11471) );
  NANDN U11077 ( .A(n11474), .B(n11473), .Z(n11476) );
  ANDN U11078 ( .B(\stack[1][42] ), .A(n5518), .Z(n11117) );
  XNOR U11079 ( .A(n11123), .B(n11477), .Z(n11116) );
  XNOR U11080 ( .A(n11124), .B(n11125), .Z(n11477) );
  AND U11081 ( .A(n11478), .B(n11479), .Z(n11125) );
  NAND U11082 ( .A(n11480), .B(n11481), .Z(n11479) );
  NANDN U11083 ( .A(n11482), .B(n11483), .Z(n11478) );
  OR U11084 ( .A(n11480), .B(n11481), .Z(n11483) );
  ANDN U11085 ( .B(\stack[1][43] ), .A(n5494), .Z(n11124) );
  XNOR U11086 ( .A(n11130), .B(n11484), .Z(n11123) );
  XNOR U11087 ( .A(n11131), .B(n11132), .Z(n11484) );
  AND U11088 ( .A(n11485), .B(n11486), .Z(n11132) );
  NANDN U11089 ( .A(n11487), .B(n11488), .Z(n11486) );
  NANDN U11090 ( .A(n11489), .B(n11490), .Z(n11485) );
  NANDN U11091 ( .A(n11488), .B(n11487), .Z(n11490) );
  ANDN U11092 ( .B(\stack[1][44] ), .A(n5470), .Z(n11131) );
  XNOR U11093 ( .A(n11137), .B(n11491), .Z(n11130) );
  XNOR U11094 ( .A(n11138), .B(n11139), .Z(n11491) );
  AND U11095 ( .A(n11492), .B(n11493), .Z(n11139) );
  NAND U11096 ( .A(n11494), .B(n11495), .Z(n11493) );
  NANDN U11097 ( .A(n11496), .B(n11497), .Z(n11492) );
  OR U11098 ( .A(n11494), .B(n11495), .Z(n11497) );
  ANDN U11099 ( .B(\stack[1][45] ), .A(n5446), .Z(n11138) );
  XNOR U11100 ( .A(n11144), .B(n11498), .Z(n11137) );
  XNOR U11101 ( .A(n11145), .B(n11146), .Z(n11498) );
  AND U11102 ( .A(n11499), .B(n11500), .Z(n11146) );
  NANDN U11103 ( .A(n11501), .B(n11502), .Z(n11500) );
  NANDN U11104 ( .A(n11503), .B(n11504), .Z(n11499) );
  NANDN U11105 ( .A(n11502), .B(n11501), .Z(n11504) );
  ANDN U11106 ( .B(\stack[1][46] ), .A(n5422), .Z(n11145) );
  XNOR U11107 ( .A(n11151), .B(n11505), .Z(n11144) );
  XNOR U11108 ( .A(n11152), .B(n11153), .Z(n11505) );
  AND U11109 ( .A(n11506), .B(n11507), .Z(n11153) );
  NAND U11110 ( .A(n11508), .B(n11509), .Z(n11507) );
  NANDN U11111 ( .A(n11510), .B(n11511), .Z(n11506) );
  OR U11112 ( .A(n11508), .B(n11509), .Z(n11511) );
  ANDN U11113 ( .B(\stack[1][47] ), .A(n5398), .Z(n11152) );
  XNOR U11114 ( .A(n11158), .B(n11512), .Z(n11151) );
  XNOR U11115 ( .A(n11159), .B(n11160), .Z(n11512) );
  AND U11116 ( .A(n11513), .B(n11514), .Z(n11160) );
  NANDN U11117 ( .A(n11515), .B(n11516), .Z(n11514) );
  NANDN U11118 ( .A(n11517), .B(n11518), .Z(n11513) );
  NANDN U11119 ( .A(n11516), .B(n11515), .Z(n11518) );
  ANDN U11120 ( .B(\stack[1][48] ), .A(n5374), .Z(n11159) );
  XNOR U11121 ( .A(n11165), .B(n11519), .Z(n11158) );
  XNOR U11122 ( .A(n11166), .B(n11167), .Z(n11519) );
  AND U11123 ( .A(n11520), .B(n11521), .Z(n11167) );
  NAND U11124 ( .A(n11522), .B(n11523), .Z(n11521) );
  NANDN U11125 ( .A(n11524), .B(n11525), .Z(n11520) );
  OR U11126 ( .A(n11522), .B(n11523), .Z(n11525) );
  ANDN U11127 ( .B(\stack[1][49] ), .A(n5350), .Z(n11166) );
  XNOR U11128 ( .A(n11172), .B(n11526), .Z(n11165) );
  XNOR U11129 ( .A(n11173), .B(n11174), .Z(n11526) );
  AND U11130 ( .A(n11527), .B(n11528), .Z(n11174) );
  NANDN U11131 ( .A(n11529), .B(n11530), .Z(n11528) );
  NANDN U11132 ( .A(n11531), .B(n11532), .Z(n11527) );
  NANDN U11133 ( .A(n11530), .B(n11529), .Z(n11532) );
  ANDN U11134 ( .B(\stack[1][50] ), .A(n5326), .Z(n11173) );
  XNOR U11135 ( .A(n11179), .B(n11533), .Z(n11172) );
  XNOR U11136 ( .A(n11180), .B(n11181), .Z(n11533) );
  AND U11137 ( .A(n11534), .B(n11535), .Z(n11181) );
  NAND U11138 ( .A(n11536), .B(n11537), .Z(n11535) );
  NANDN U11139 ( .A(n11538), .B(n11539), .Z(n11534) );
  OR U11140 ( .A(n11536), .B(n11537), .Z(n11539) );
  ANDN U11141 ( .B(\stack[1][51] ), .A(n5302), .Z(n11180) );
  XNOR U11142 ( .A(n11186), .B(n11540), .Z(n11179) );
  XNOR U11143 ( .A(n11187), .B(n11188), .Z(n11540) );
  AND U11144 ( .A(n11541), .B(n11542), .Z(n11188) );
  NANDN U11145 ( .A(n11543), .B(n11544), .Z(n11542) );
  NANDN U11146 ( .A(n11545), .B(n11546), .Z(n11541) );
  NANDN U11147 ( .A(n11544), .B(n11543), .Z(n11546) );
  ANDN U11148 ( .B(\stack[1][52] ), .A(n5278), .Z(n11187) );
  XNOR U11149 ( .A(n11193), .B(n11547), .Z(n11186) );
  XNOR U11150 ( .A(n11194), .B(n11195), .Z(n11547) );
  AND U11151 ( .A(n11548), .B(n11549), .Z(n11195) );
  NAND U11152 ( .A(n11550), .B(n11551), .Z(n11549) );
  NANDN U11153 ( .A(n11552), .B(n11553), .Z(n11548) );
  OR U11154 ( .A(n11550), .B(n11551), .Z(n11553) );
  ANDN U11155 ( .B(\stack[1][53] ), .A(n5254), .Z(n11194) );
  XNOR U11156 ( .A(n11200), .B(n11554), .Z(n11193) );
  XNOR U11157 ( .A(n11201), .B(n11202), .Z(n11554) );
  AND U11158 ( .A(n11555), .B(n11556), .Z(n11202) );
  NAND U11159 ( .A(n11557), .B(n11558), .Z(n11556) );
  NAND U11160 ( .A(n11559), .B(n11560), .Z(n11555) );
  OR U11161 ( .A(n11557), .B(n11558), .Z(n11559) );
  ANDN U11162 ( .B(\stack[1][54] ), .A(n5230), .Z(n11201) );
  XNOR U11163 ( .A(n11207), .B(n11561), .Z(n11200) );
  XNOR U11164 ( .A(n11208), .B(n11210), .Z(n11561) );
  ANDN U11165 ( .B(n11562), .A(n11563), .Z(n11210) );
  ANDN U11166 ( .B(\stack[0][0] ), .A(n6516), .Z(n11562) );
  ANDN U11167 ( .B(\stack[1][55] ), .A(n5206), .Z(n11208) );
  XOR U11168 ( .A(n11213), .B(n11564), .Z(n11207) );
  NANDN U11169 ( .A(n5160), .B(\stack[1][57] ), .Z(n11564) );
  NANDN U11170 ( .A(n6516), .B(\stack[0][1] ), .Z(n11213) );
  ANDN U11171 ( .B(\stack[1][5] ), .A(n6406), .Z(n8999) );
  AND U11172 ( .A(n11565), .B(n11566), .Z(n9000) );
  NANDN U11173 ( .A(n9004), .B(n9006), .Z(n11566) );
  NANDN U11174 ( .A(n9007), .B(n11567), .Z(n11565) );
  NANDN U11175 ( .A(n9006), .B(n9004), .Z(n11567) );
  XOR U11176 ( .A(n11221), .B(n11568), .Z(n9004) );
  XNOR U11177 ( .A(n11222), .B(n11223), .Z(n11568) );
  AND U11178 ( .A(n11569), .B(n11570), .Z(n11223) );
  NAND U11179 ( .A(n11571), .B(n11572), .Z(n11570) );
  NANDN U11180 ( .A(n11573), .B(n11574), .Z(n11569) );
  OR U11181 ( .A(n11571), .B(n11572), .Z(n11574) );
  ANDN U11182 ( .B(\stack[0][50] ), .A(n5316), .Z(n11222) );
  XNOR U11183 ( .A(n11228), .B(n11575), .Z(n11221) );
  XNOR U11184 ( .A(n11229), .B(n11230), .Z(n11575) );
  AND U11185 ( .A(n11576), .B(n11577), .Z(n11230) );
  NANDN U11186 ( .A(n11578), .B(n11579), .Z(n11577) );
  NANDN U11187 ( .A(n11580), .B(n11581), .Z(n11576) );
  NANDN U11188 ( .A(n11579), .B(n11578), .Z(n11581) );
  ANDN U11189 ( .B(\stack[0][49] ), .A(n5340), .Z(n11229) );
  XNOR U11190 ( .A(n11235), .B(n11582), .Z(n11228) );
  XNOR U11191 ( .A(n11236), .B(n11237), .Z(n11582) );
  AND U11192 ( .A(n11583), .B(n11584), .Z(n11237) );
  NAND U11193 ( .A(n11585), .B(n11586), .Z(n11584) );
  NANDN U11194 ( .A(n11587), .B(n11588), .Z(n11583) );
  OR U11195 ( .A(n11585), .B(n11586), .Z(n11588) );
  ANDN U11196 ( .B(\stack[0][48] ), .A(n5364), .Z(n11236) );
  XNOR U11197 ( .A(n11242), .B(n11589), .Z(n11235) );
  XNOR U11198 ( .A(n11243), .B(n11244), .Z(n11589) );
  AND U11199 ( .A(n11590), .B(n11591), .Z(n11244) );
  NANDN U11200 ( .A(n11592), .B(n11593), .Z(n11591) );
  NANDN U11201 ( .A(n11594), .B(n11595), .Z(n11590) );
  NANDN U11202 ( .A(n11593), .B(n11592), .Z(n11595) );
  ANDN U11203 ( .B(\stack[0][47] ), .A(n5387), .Z(n11243) );
  XNOR U11204 ( .A(n11249), .B(n11596), .Z(n11242) );
  XNOR U11205 ( .A(n11250), .B(n11251), .Z(n11596) );
  AND U11206 ( .A(n11597), .B(n11598), .Z(n11251) );
  NAND U11207 ( .A(n11599), .B(n11600), .Z(n11598) );
  NANDN U11208 ( .A(n11601), .B(n11602), .Z(n11597) );
  OR U11209 ( .A(n11599), .B(n11600), .Z(n11602) );
  ANDN U11210 ( .B(\stack[1][10] ), .A(n6262), .Z(n11250) );
  XNOR U11211 ( .A(n11256), .B(n11603), .Z(n11249) );
  XNOR U11212 ( .A(n11257), .B(n11258), .Z(n11603) );
  AND U11213 ( .A(n11604), .B(n11605), .Z(n11258) );
  NANDN U11214 ( .A(n11606), .B(n11607), .Z(n11605) );
  NANDN U11215 ( .A(n11608), .B(n11609), .Z(n11604) );
  NANDN U11216 ( .A(n11607), .B(n11606), .Z(n11609) );
  ANDN U11217 ( .B(\stack[1][11] ), .A(n6238), .Z(n11257) );
  XNOR U11218 ( .A(n11263), .B(n11610), .Z(n11256) );
  XNOR U11219 ( .A(n11264), .B(n11265), .Z(n11610) );
  AND U11220 ( .A(n11611), .B(n11612), .Z(n11265) );
  NAND U11221 ( .A(n11613), .B(n11614), .Z(n11612) );
  NANDN U11222 ( .A(n11615), .B(n11616), .Z(n11611) );
  OR U11223 ( .A(n11613), .B(n11614), .Z(n11616) );
  ANDN U11224 ( .B(\stack[1][12] ), .A(n6214), .Z(n11264) );
  XNOR U11225 ( .A(n11270), .B(n11617), .Z(n11263) );
  XNOR U11226 ( .A(n11271), .B(n11272), .Z(n11617) );
  AND U11227 ( .A(n11618), .B(n11619), .Z(n11272) );
  NANDN U11228 ( .A(n11620), .B(n11621), .Z(n11619) );
  NANDN U11229 ( .A(n11622), .B(n11623), .Z(n11618) );
  NANDN U11230 ( .A(n11621), .B(n11620), .Z(n11623) );
  ANDN U11231 ( .B(\stack[1][13] ), .A(n6190), .Z(n11271) );
  XNOR U11232 ( .A(n11277), .B(n11624), .Z(n11270) );
  XNOR U11233 ( .A(n11278), .B(n11279), .Z(n11624) );
  AND U11234 ( .A(n11625), .B(n11626), .Z(n11279) );
  NAND U11235 ( .A(n11627), .B(n11628), .Z(n11626) );
  NANDN U11236 ( .A(n11629), .B(n11630), .Z(n11625) );
  OR U11237 ( .A(n11627), .B(n11628), .Z(n11630) );
  ANDN U11238 ( .B(\stack[1][14] ), .A(n6166), .Z(n11278) );
  XNOR U11239 ( .A(n11284), .B(n11631), .Z(n11277) );
  XNOR U11240 ( .A(n11285), .B(n11286), .Z(n11631) );
  AND U11241 ( .A(n11632), .B(n11633), .Z(n11286) );
  NANDN U11242 ( .A(n11634), .B(n11635), .Z(n11633) );
  NANDN U11243 ( .A(n11636), .B(n11637), .Z(n11632) );
  NANDN U11244 ( .A(n11635), .B(n11634), .Z(n11637) );
  ANDN U11245 ( .B(\stack[1][15] ), .A(n6142), .Z(n11285) );
  XNOR U11246 ( .A(n11291), .B(n11638), .Z(n11284) );
  XNOR U11247 ( .A(n11292), .B(n11293), .Z(n11638) );
  AND U11248 ( .A(n11639), .B(n11640), .Z(n11293) );
  NAND U11249 ( .A(n11641), .B(n11642), .Z(n11640) );
  NANDN U11250 ( .A(n11643), .B(n11644), .Z(n11639) );
  OR U11251 ( .A(n11641), .B(n11642), .Z(n11644) );
  ANDN U11252 ( .B(\stack[1][16] ), .A(n6118), .Z(n11292) );
  XNOR U11253 ( .A(n11298), .B(n11645), .Z(n11291) );
  XNOR U11254 ( .A(n11299), .B(n11300), .Z(n11645) );
  AND U11255 ( .A(n11646), .B(n11647), .Z(n11300) );
  NANDN U11256 ( .A(n11648), .B(n11649), .Z(n11647) );
  NANDN U11257 ( .A(n11650), .B(n11651), .Z(n11646) );
  NANDN U11258 ( .A(n11649), .B(n11648), .Z(n11651) );
  ANDN U11259 ( .B(\stack[1][17] ), .A(n6094), .Z(n11299) );
  XNOR U11260 ( .A(n11305), .B(n11652), .Z(n11298) );
  XNOR U11261 ( .A(n11306), .B(n11307), .Z(n11652) );
  AND U11262 ( .A(n11653), .B(n11654), .Z(n11307) );
  NAND U11263 ( .A(n11655), .B(n11656), .Z(n11654) );
  NANDN U11264 ( .A(n11657), .B(n11658), .Z(n11653) );
  OR U11265 ( .A(n11655), .B(n11656), .Z(n11658) );
  ANDN U11266 ( .B(\stack[1][18] ), .A(n6070), .Z(n11306) );
  XNOR U11267 ( .A(n11312), .B(n11659), .Z(n11305) );
  XNOR U11268 ( .A(n11313), .B(n11314), .Z(n11659) );
  AND U11269 ( .A(n11660), .B(n11661), .Z(n11314) );
  NANDN U11270 ( .A(n11662), .B(n11663), .Z(n11661) );
  NANDN U11271 ( .A(n11664), .B(n11665), .Z(n11660) );
  NANDN U11272 ( .A(n11663), .B(n11662), .Z(n11665) );
  ANDN U11273 ( .B(\stack[1][19] ), .A(n6046), .Z(n11313) );
  XNOR U11274 ( .A(n11319), .B(n11666), .Z(n11312) );
  XNOR U11275 ( .A(n11320), .B(n11321), .Z(n11666) );
  AND U11276 ( .A(n11667), .B(n11668), .Z(n11321) );
  NAND U11277 ( .A(n11669), .B(n11670), .Z(n11668) );
  NANDN U11278 ( .A(n11671), .B(n11672), .Z(n11667) );
  OR U11279 ( .A(n11669), .B(n11670), .Z(n11672) );
  ANDN U11280 ( .B(\stack[1][20] ), .A(n6022), .Z(n11320) );
  XNOR U11281 ( .A(n11326), .B(n11673), .Z(n11319) );
  XNOR U11282 ( .A(n11327), .B(n11328), .Z(n11673) );
  AND U11283 ( .A(n11674), .B(n11675), .Z(n11328) );
  NANDN U11284 ( .A(n11676), .B(n11677), .Z(n11675) );
  NANDN U11285 ( .A(n11678), .B(n11679), .Z(n11674) );
  NANDN U11286 ( .A(n11677), .B(n11676), .Z(n11679) );
  ANDN U11287 ( .B(\stack[1][21] ), .A(n5998), .Z(n11327) );
  XNOR U11288 ( .A(n11333), .B(n11680), .Z(n11326) );
  XNOR U11289 ( .A(n11334), .B(n11335), .Z(n11680) );
  AND U11290 ( .A(n11681), .B(n11682), .Z(n11335) );
  NAND U11291 ( .A(n11683), .B(n11684), .Z(n11682) );
  NANDN U11292 ( .A(n11685), .B(n11686), .Z(n11681) );
  OR U11293 ( .A(n11683), .B(n11684), .Z(n11686) );
  ANDN U11294 ( .B(\stack[1][22] ), .A(n5974), .Z(n11334) );
  XNOR U11295 ( .A(n11340), .B(n11687), .Z(n11333) );
  XNOR U11296 ( .A(n11341), .B(n11342), .Z(n11687) );
  AND U11297 ( .A(n11688), .B(n11689), .Z(n11342) );
  NANDN U11298 ( .A(n11690), .B(n11691), .Z(n11689) );
  NANDN U11299 ( .A(n11692), .B(n11693), .Z(n11688) );
  NANDN U11300 ( .A(n11691), .B(n11690), .Z(n11693) );
  ANDN U11301 ( .B(\stack[1][23] ), .A(n5950), .Z(n11341) );
  XNOR U11302 ( .A(n11347), .B(n11694), .Z(n11340) );
  XNOR U11303 ( .A(n11348), .B(n11349), .Z(n11694) );
  AND U11304 ( .A(n11695), .B(n11696), .Z(n11349) );
  NAND U11305 ( .A(n11697), .B(n11698), .Z(n11696) );
  NANDN U11306 ( .A(n11699), .B(n11700), .Z(n11695) );
  OR U11307 ( .A(n11697), .B(n11698), .Z(n11700) );
  ANDN U11308 ( .B(\stack[1][24] ), .A(n5926), .Z(n11348) );
  XNOR U11309 ( .A(n11354), .B(n11701), .Z(n11347) );
  XNOR U11310 ( .A(n11355), .B(n11356), .Z(n11701) );
  AND U11311 ( .A(n11702), .B(n11703), .Z(n11356) );
  NANDN U11312 ( .A(n11704), .B(n11705), .Z(n11703) );
  NANDN U11313 ( .A(n11706), .B(n11707), .Z(n11702) );
  NANDN U11314 ( .A(n11705), .B(n11704), .Z(n11707) );
  ANDN U11315 ( .B(\stack[1][25] ), .A(n5902), .Z(n11355) );
  XNOR U11316 ( .A(n11361), .B(n11708), .Z(n11354) );
  XNOR U11317 ( .A(n11362), .B(n11363), .Z(n11708) );
  AND U11318 ( .A(n11709), .B(n11710), .Z(n11363) );
  NAND U11319 ( .A(n11711), .B(n11712), .Z(n11710) );
  NANDN U11320 ( .A(n11713), .B(n11714), .Z(n11709) );
  OR U11321 ( .A(n11711), .B(n11712), .Z(n11714) );
  ANDN U11322 ( .B(\stack[1][26] ), .A(n5878), .Z(n11362) );
  XNOR U11323 ( .A(n11368), .B(n11715), .Z(n11361) );
  XNOR U11324 ( .A(n11369), .B(n11370), .Z(n11715) );
  AND U11325 ( .A(n11716), .B(n11717), .Z(n11370) );
  NANDN U11326 ( .A(n11718), .B(n11719), .Z(n11717) );
  NANDN U11327 ( .A(n11720), .B(n11721), .Z(n11716) );
  NANDN U11328 ( .A(n11719), .B(n11718), .Z(n11721) );
  ANDN U11329 ( .B(\stack[1][27] ), .A(n5854), .Z(n11369) );
  XNOR U11330 ( .A(n11375), .B(n11722), .Z(n11368) );
  XNOR U11331 ( .A(n11376), .B(n11377), .Z(n11722) );
  AND U11332 ( .A(n11723), .B(n11724), .Z(n11377) );
  NAND U11333 ( .A(n11725), .B(n11726), .Z(n11724) );
  NANDN U11334 ( .A(n11727), .B(n11728), .Z(n11723) );
  OR U11335 ( .A(n11725), .B(n11726), .Z(n11728) );
  ANDN U11336 ( .B(\stack[1][28] ), .A(n5830), .Z(n11376) );
  XNOR U11337 ( .A(n11382), .B(n11729), .Z(n11375) );
  XNOR U11338 ( .A(n11383), .B(n11384), .Z(n11729) );
  AND U11339 ( .A(n11730), .B(n11731), .Z(n11384) );
  NANDN U11340 ( .A(n11732), .B(n11733), .Z(n11731) );
  NANDN U11341 ( .A(n11734), .B(n11735), .Z(n11730) );
  NANDN U11342 ( .A(n11733), .B(n11732), .Z(n11735) );
  ANDN U11343 ( .B(\stack[1][29] ), .A(n5806), .Z(n11383) );
  XNOR U11344 ( .A(n11389), .B(n11736), .Z(n11382) );
  XNOR U11345 ( .A(n11390), .B(n11391), .Z(n11736) );
  AND U11346 ( .A(n11737), .B(n11738), .Z(n11391) );
  NAND U11347 ( .A(n11739), .B(n11740), .Z(n11738) );
  NANDN U11348 ( .A(n11741), .B(n11742), .Z(n11737) );
  OR U11349 ( .A(n11739), .B(n11740), .Z(n11742) );
  ANDN U11350 ( .B(\stack[1][30] ), .A(n5782), .Z(n11390) );
  XNOR U11351 ( .A(n11396), .B(n11743), .Z(n11389) );
  XNOR U11352 ( .A(n11397), .B(n11398), .Z(n11743) );
  AND U11353 ( .A(n11744), .B(n11745), .Z(n11398) );
  NANDN U11354 ( .A(n11746), .B(n11747), .Z(n11745) );
  NANDN U11355 ( .A(n11748), .B(n11749), .Z(n11744) );
  NANDN U11356 ( .A(n11747), .B(n11746), .Z(n11749) );
  ANDN U11357 ( .B(\stack[1][31] ), .A(n5758), .Z(n11397) );
  XNOR U11358 ( .A(n11403), .B(n11750), .Z(n11396) );
  XNOR U11359 ( .A(n11404), .B(n11405), .Z(n11750) );
  AND U11360 ( .A(n11751), .B(n11752), .Z(n11405) );
  NAND U11361 ( .A(n11753), .B(n11754), .Z(n11752) );
  NANDN U11362 ( .A(n11755), .B(n11756), .Z(n11751) );
  OR U11363 ( .A(n11753), .B(n11754), .Z(n11756) );
  ANDN U11364 ( .B(\stack[1][32] ), .A(n5734), .Z(n11404) );
  XNOR U11365 ( .A(n11410), .B(n11757), .Z(n11403) );
  XNOR U11366 ( .A(n11411), .B(n11412), .Z(n11757) );
  AND U11367 ( .A(n11758), .B(n11759), .Z(n11412) );
  NANDN U11368 ( .A(n11760), .B(n11761), .Z(n11759) );
  NANDN U11369 ( .A(n11762), .B(n11763), .Z(n11758) );
  NANDN U11370 ( .A(n11761), .B(n11760), .Z(n11763) );
  ANDN U11371 ( .B(\stack[1][33] ), .A(n5710), .Z(n11411) );
  XNOR U11372 ( .A(n11417), .B(n11764), .Z(n11410) );
  XNOR U11373 ( .A(n11418), .B(n11419), .Z(n11764) );
  AND U11374 ( .A(n11765), .B(n11766), .Z(n11419) );
  NAND U11375 ( .A(n11767), .B(n11768), .Z(n11766) );
  NANDN U11376 ( .A(n11769), .B(n11770), .Z(n11765) );
  OR U11377 ( .A(n11767), .B(n11768), .Z(n11770) );
  ANDN U11378 ( .B(\stack[1][34] ), .A(n5686), .Z(n11418) );
  XNOR U11379 ( .A(n11424), .B(n11771), .Z(n11417) );
  XNOR U11380 ( .A(n11425), .B(n11426), .Z(n11771) );
  AND U11381 ( .A(n11772), .B(n11773), .Z(n11426) );
  NANDN U11382 ( .A(n11774), .B(n11775), .Z(n11773) );
  NANDN U11383 ( .A(n11776), .B(n11777), .Z(n11772) );
  NANDN U11384 ( .A(n11775), .B(n11774), .Z(n11777) );
  ANDN U11385 ( .B(\stack[1][35] ), .A(n5662), .Z(n11425) );
  XNOR U11386 ( .A(n11431), .B(n11778), .Z(n11424) );
  XNOR U11387 ( .A(n11432), .B(n11433), .Z(n11778) );
  AND U11388 ( .A(n11779), .B(n11780), .Z(n11433) );
  NAND U11389 ( .A(n11781), .B(n11782), .Z(n11780) );
  NANDN U11390 ( .A(n11783), .B(n11784), .Z(n11779) );
  OR U11391 ( .A(n11781), .B(n11782), .Z(n11784) );
  ANDN U11392 ( .B(\stack[1][36] ), .A(n5638), .Z(n11432) );
  XNOR U11393 ( .A(n11439), .B(n11785), .Z(n11431) );
  XOR U11394 ( .A(n11440), .B(n11441), .Z(n11785) );
  NAND U11395 ( .A(n11786), .B(n11787), .Z(n11441) );
  NANDN U11396 ( .A(n11788), .B(n11789), .Z(n11787) );
  OR U11397 ( .A(n11790), .B(n11791), .Z(n11789) );
  AND U11398 ( .A(\stack[0][19] ), .B(\stack[1][37] ), .Z(n11440) );
  XNOR U11399 ( .A(n11446), .B(n11792), .Z(n11439) );
  XNOR U11400 ( .A(n11445), .B(n11448), .Z(n11792) );
  AND U11401 ( .A(\stack[0][18] ), .B(\stack[1][38] ), .Z(n11448) );
  AND U11402 ( .A(n11793), .B(n11794), .Z(n11445) );
  NAND U11403 ( .A(n11795), .B(n11796), .Z(n11794) );
  OR U11404 ( .A(n11797), .B(n11798), .Z(n11795) );
  XNOR U11405 ( .A(n11452), .B(n11799), .Z(n11446) );
  XNOR U11406 ( .A(n11453), .B(n11454), .Z(n11799) );
  AND U11407 ( .A(n11800), .B(n11801), .Z(n11454) );
  NANDN U11408 ( .A(n11802), .B(n11803), .Z(n11801) );
  NANDN U11409 ( .A(n11804), .B(n11805), .Z(n11800) );
  NANDN U11410 ( .A(n11803), .B(n11802), .Z(n11805) );
  ANDN U11411 ( .B(\stack[1][39] ), .A(n5566), .Z(n11453) );
  XNOR U11412 ( .A(n11459), .B(n11806), .Z(n11452) );
  XNOR U11413 ( .A(n11460), .B(n11461), .Z(n11806) );
  AND U11414 ( .A(n11807), .B(n11808), .Z(n11461) );
  NAND U11415 ( .A(n11809), .B(n11810), .Z(n11808) );
  NANDN U11416 ( .A(n11811), .B(n11812), .Z(n11807) );
  OR U11417 ( .A(n11809), .B(n11810), .Z(n11812) );
  ANDN U11418 ( .B(\stack[1][40] ), .A(n5542), .Z(n11460) );
  XNOR U11419 ( .A(n11466), .B(n11813), .Z(n11459) );
  XNOR U11420 ( .A(n11467), .B(n11468), .Z(n11813) );
  AND U11421 ( .A(n11814), .B(n11815), .Z(n11468) );
  NANDN U11422 ( .A(n11816), .B(n11817), .Z(n11815) );
  NANDN U11423 ( .A(n11818), .B(n11819), .Z(n11814) );
  NANDN U11424 ( .A(n11817), .B(n11816), .Z(n11819) );
  ANDN U11425 ( .B(\stack[1][41] ), .A(n5518), .Z(n11467) );
  XNOR U11426 ( .A(n11473), .B(n11820), .Z(n11466) );
  XNOR U11427 ( .A(n11474), .B(n11475), .Z(n11820) );
  AND U11428 ( .A(n11821), .B(n11822), .Z(n11475) );
  NAND U11429 ( .A(n11823), .B(n11824), .Z(n11822) );
  NANDN U11430 ( .A(n11825), .B(n11826), .Z(n11821) );
  OR U11431 ( .A(n11823), .B(n11824), .Z(n11826) );
  ANDN U11432 ( .B(\stack[1][42] ), .A(n5494), .Z(n11474) );
  XNOR U11433 ( .A(n11480), .B(n11827), .Z(n11473) );
  XNOR U11434 ( .A(n11481), .B(n11482), .Z(n11827) );
  AND U11435 ( .A(n11828), .B(n11829), .Z(n11482) );
  NANDN U11436 ( .A(n11830), .B(n11831), .Z(n11829) );
  NANDN U11437 ( .A(n11832), .B(n11833), .Z(n11828) );
  NANDN U11438 ( .A(n11831), .B(n11830), .Z(n11833) );
  ANDN U11439 ( .B(\stack[1][43] ), .A(n5470), .Z(n11481) );
  XNOR U11440 ( .A(n11487), .B(n11834), .Z(n11480) );
  XNOR U11441 ( .A(n11488), .B(n11489), .Z(n11834) );
  AND U11442 ( .A(n11835), .B(n11836), .Z(n11489) );
  NAND U11443 ( .A(n11837), .B(n11838), .Z(n11836) );
  NANDN U11444 ( .A(n11839), .B(n11840), .Z(n11835) );
  OR U11445 ( .A(n11837), .B(n11838), .Z(n11840) );
  ANDN U11446 ( .B(\stack[1][44] ), .A(n5446), .Z(n11488) );
  XNOR U11447 ( .A(n11494), .B(n11841), .Z(n11487) );
  XNOR U11448 ( .A(n11495), .B(n11496), .Z(n11841) );
  AND U11449 ( .A(n11842), .B(n11843), .Z(n11496) );
  NANDN U11450 ( .A(n11844), .B(n11845), .Z(n11843) );
  NANDN U11451 ( .A(n11846), .B(n11847), .Z(n11842) );
  NANDN U11452 ( .A(n11845), .B(n11844), .Z(n11847) );
  ANDN U11453 ( .B(\stack[1][45] ), .A(n5422), .Z(n11495) );
  XNOR U11454 ( .A(n11501), .B(n11848), .Z(n11494) );
  XNOR U11455 ( .A(n11502), .B(n11503), .Z(n11848) );
  AND U11456 ( .A(n11849), .B(n11850), .Z(n11503) );
  NAND U11457 ( .A(n11851), .B(n11852), .Z(n11850) );
  NANDN U11458 ( .A(n11853), .B(n11854), .Z(n11849) );
  OR U11459 ( .A(n11851), .B(n11852), .Z(n11854) );
  ANDN U11460 ( .B(\stack[1][46] ), .A(n5398), .Z(n11502) );
  XNOR U11461 ( .A(n11508), .B(n11855), .Z(n11501) );
  XNOR U11462 ( .A(n11509), .B(n11510), .Z(n11855) );
  AND U11463 ( .A(n11856), .B(n11857), .Z(n11510) );
  NANDN U11464 ( .A(n11858), .B(n11859), .Z(n11857) );
  NANDN U11465 ( .A(n11860), .B(n11861), .Z(n11856) );
  NANDN U11466 ( .A(n11859), .B(n11858), .Z(n11861) );
  ANDN U11467 ( .B(\stack[1][47] ), .A(n5374), .Z(n11509) );
  XNOR U11468 ( .A(n11515), .B(n11862), .Z(n11508) );
  XNOR U11469 ( .A(n11516), .B(n11517), .Z(n11862) );
  AND U11470 ( .A(n11863), .B(n11864), .Z(n11517) );
  NAND U11471 ( .A(n11865), .B(n11866), .Z(n11864) );
  NANDN U11472 ( .A(n11867), .B(n11868), .Z(n11863) );
  OR U11473 ( .A(n11865), .B(n11866), .Z(n11868) );
  ANDN U11474 ( .B(\stack[1][48] ), .A(n5350), .Z(n11516) );
  XNOR U11475 ( .A(n11522), .B(n11869), .Z(n11515) );
  XNOR U11476 ( .A(n11523), .B(n11524), .Z(n11869) );
  AND U11477 ( .A(n11870), .B(n11871), .Z(n11524) );
  NANDN U11478 ( .A(n11872), .B(n11873), .Z(n11871) );
  NANDN U11479 ( .A(n11874), .B(n11875), .Z(n11870) );
  NANDN U11480 ( .A(n11873), .B(n11872), .Z(n11875) );
  ANDN U11481 ( .B(\stack[1][49] ), .A(n5326), .Z(n11523) );
  XNOR U11482 ( .A(n11529), .B(n11876), .Z(n11522) );
  XNOR U11483 ( .A(n11530), .B(n11531), .Z(n11876) );
  AND U11484 ( .A(n11877), .B(n11878), .Z(n11531) );
  NAND U11485 ( .A(n11879), .B(n11880), .Z(n11878) );
  NANDN U11486 ( .A(n11881), .B(n11882), .Z(n11877) );
  OR U11487 ( .A(n11879), .B(n11880), .Z(n11882) );
  ANDN U11488 ( .B(\stack[1][50] ), .A(n5302), .Z(n11530) );
  XNOR U11489 ( .A(n11536), .B(n11883), .Z(n11529) );
  XNOR U11490 ( .A(n11537), .B(n11538), .Z(n11883) );
  AND U11491 ( .A(n11884), .B(n11885), .Z(n11538) );
  NANDN U11492 ( .A(n11886), .B(n11887), .Z(n11885) );
  NANDN U11493 ( .A(n11888), .B(n11889), .Z(n11884) );
  NANDN U11494 ( .A(n11887), .B(n11886), .Z(n11889) );
  ANDN U11495 ( .B(\stack[1][51] ), .A(n5278), .Z(n11537) );
  XNOR U11496 ( .A(n11543), .B(n11890), .Z(n11536) );
  XNOR U11497 ( .A(n11544), .B(n11545), .Z(n11890) );
  AND U11498 ( .A(n11891), .B(n11892), .Z(n11545) );
  NAND U11499 ( .A(n11893), .B(n11894), .Z(n11892) );
  NANDN U11500 ( .A(n11895), .B(n11896), .Z(n11891) );
  OR U11501 ( .A(n11893), .B(n11894), .Z(n11896) );
  ANDN U11502 ( .B(\stack[1][52] ), .A(n5254), .Z(n11544) );
  XNOR U11503 ( .A(n11550), .B(n11897), .Z(n11543) );
  XNOR U11504 ( .A(n11551), .B(n11552), .Z(n11897) );
  AND U11505 ( .A(n11898), .B(n11899), .Z(n11552) );
  NAND U11506 ( .A(n11900), .B(n11901), .Z(n11899) );
  NAND U11507 ( .A(n11902), .B(n11903), .Z(n11898) );
  OR U11508 ( .A(n11900), .B(n11901), .Z(n11902) );
  ANDN U11509 ( .B(\stack[1][53] ), .A(n5230), .Z(n11551) );
  XNOR U11510 ( .A(n11557), .B(n11904), .Z(n11550) );
  XNOR U11511 ( .A(n11558), .B(n11560), .Z(n11904) );
  ANDN U11512 ( .B(n11905), .A(n11906), .Z(n11560) );
  ANDN U11513 ( .B(\stack[0][0] ), .A(n6492), .Z(n11905) );
  ANDN U11514 ( .B(\stack[1][54] ), .A(n5206), .Z(n11558) );
  XOR U11515 ( .A(n11563), .B(n11907), .Z(n11557) );
  NANDN U11516 ( .A(n5160), .B(\stack[1][56] ), .Z(n11907) );
  NANDN U11517 ( .A(n6492), .B(\stack[0][1] ), .Z(n11563) );
  ANDN U11518 ( .B(\stack[0][51] ), .A(n5292), .Z(n9006) );
  AND U11519 ( .A(n11908), .B(n11909), .Z(n9007) );
  OR U11520 ( .A(n9011), .B(n11910), .Z(n11909) );
  IV U11521 ( .A(n9013), .Z(n11910) );
  NANDN U11522 ( .A(n9014), .B(n11911), .Z(n11908) );
  NANDN U11523 ( .A(n9013), .B(n9011), .Z(n11911) );
  XNOR U11524 ( .A(n11571), .B(n11912), .Z(n9011) );
  XNOR U11525 ( .A(n11572), .B(n11573), .Z(n11912) );
  AND U11526 ( .A(n11913), .B(n11914), .Z(n11573) );
  NANDN U11527 ( .A(n11915), .B(n11916), .Z(n11914) );
  NANDN U11528 ( .A(n11917), .B(n11918), .Z(n11913) );
  NANDN U11529 ( .A(n11916), .B(n11915), .Z(n11918) );
  ANDN U11530 ( .B(\stack[0][49] ), .A(n5316), .Z(n11572) );
  XNOR U11531 ( .A(n11578), .B(n11919), .Z(n11571) );
  XNOR U11532 ( .A(n11579), .B(n11580), .Z(n11919) );
  AND U11533 ( .A(n11920), .B(n11921), .Z(n11580) );
  NAND U11534 ( .A(n11922), .B(n11923), .Z(n11921) );
  NANDN U11535 ( .A(n11924), .B(n11925), .Z(n11920) );
  OR U11536 ( .A(n11922), .B(n11923), .Z(n11925) );
  ANDN U11537 ( .B(\stack[0][48] ), .A(n5340), .Z(n11579) );
  XNOR U11538 ( .A(n11585), .B(n11926), .Z(n11578) );
  XNOR U11539 ( .A(n11586), .B(n11587), .Z(n11926) );
  AND U11540 ( .A(n11927), .B(n11928), .Z(n11587) );
  NANDN U11541 ( .A(n11929), .B(n11930), .Z(n11928) );
  NANDN U11542 ( .A(n11931), .B(n11932), .Z(n11927) );
  NANDN U11543 ( .A(n11930), .B(n11929), .Z(n11932) );
  ANDN U11544 ( .B(\stack[0][47] ), .A(n5364), .Z(n11586) );
  XNOR U11545 ( .A(n11592), .B(n11933), .Z(n11585) );
  XNOR U11546 ( .A(n11593), .B(n11594), .Z(n11933) );
  AND U11547 ( .A(n11934), .B(n11935), .Z(n11594) );
  NAND U11548 ( .A(n11936), .B(n11937), .Z(n11935) );
  NANDN U11549 ( .A(n11938), .B(n11939), .Z(n11934) );
  OR U11550 ( .A(n11936), .B(n11937), .Z(n11939) );
  ANDN U11551 ( .B(\stack[0][46] ), .A(n5387), .Z(n11593) );
  XNOR U11552 ( .A(n11599), .B(n11940), .Z(n11592) );
  XNOR U11553 ( .A(n11600), .B(n11601), .Z(n11940) );
  AND U11554 ( .A(n11941), .B(n11942), .Z(n11601) );
  NANDN U11555 ( .A(n11943), .B(n11944), .Z(n11942) );
  NANDN U11556 ( .A(n11945), .B(n11946), .Z(n11941) );
  NANDN U11557 ( .A(n11944), .B(n11943), .Z(n11946) );
  ANDN U11558 ( .B(\stack[1][10] ), .A(n6238), .Z(n11600) );
  XNOR U11559 ( .A(n11606), .B(n11947), .Z(n11599) );
  XNOR U11560 ( .A(n11607), .B(n11608), .Z(n11947) );
  AND U11561 ( .A(n11948), .B(n11949), .Z(n11608) );
  NAND U11562 ( .A(n11950), .B(n11951), .Z(n11949) );
  NANDN U11563 ( .A(n11952), .B(n11953), .Z(n11948) );
  OR U11564 ( .A(n11950), .B(n11951), .Z(n11953) );
  ANDN U11565 ( .B(\stack[1][11] ), .A(n6214), .Z(n11607) );
  XNOR U11566 ( .A(n11613), .B(n11954), .Z(n11606) );
  XNOR U11567 ( .A(n11614), .B(n11615), .Z(n11954) );
  AND U11568 ( .A(n11955), .B(n11956), .Z(n11615) );
  NANDN U11569 ( .A(n11957), .B(n11958), .Z(n11956) );
  NANDN U11570 ( .A(n11959), .B(n11960), .Z(n11955) );
  NANDN U11571 ( .A(n11958), .B(n11957), .Z(n11960) );
  ANDN U11572 ( .B(\stack[1][12] ), .A(n6190), .Z(n11614) );
  XNOR U11573 ( .A(n11620), .B(n11961), .Z(n11613) );
  XNOR U11574 ( .A(n11621), .B(n11622), .Z(n11961) );
  AND U11575 ( .A(n11962), .B(n11963), .Z(n11622) );
  NAND U11576 ( .A(n11964), .B(n11965), .Z(n11963) );
  NANDN U11577 ( .A(n11966), .B(n11967), .Z(n11962) );
  OR U11578 ( .A(n11964), .B(n11965), .Z(n11967) );
  ANDN U11579 ( .B(\stack[1][13] ), .A(n6166), .Z(n11621) );
  XNOR U11580 ( .A(n11627), .B(n11968), .Z(n11620) );
  XNOR U11581 ( .A(n11628), .B(n11629), .Z(n11968) );
  AND U11582 ( .A(n11969), .B(n11970), .Z(n11629) );
  NANDN U11583 ( .A(n11971), .B(n11972), .Z(n11970) );
  NANDN U11584 ( .A(n11973), .B(n11974), .Z(n11969) );
  NANDN U11585 ( .A(n11972), .B(n11971), .Z(n11974) );
  ANDN U11586 ( .B(\stack[1][14] ), .A(n6142), .Z(n11628) );
  XNOR U11587 ( .A(n11634), .B(n11975), .Z(n11627) );
  XNOR U11588 ( .A(n11635), .B(n11636), .Z(n11975) );
  AND U11589 ( .A(n11976), .B(n11977), .Z(n11636) );
  NAND U11590 ( .A(n11978), .B(n11979), .Z(n11977) );
  NANDN U11591 ( .A(n11980), .B(n11981), .Z(n11976) );
  OR U11592 ( .A(n11978), .B(n11979), .Z(n11981) );
  ANDN U11593 ( .B(\stack[1][15] ), .A(n6118), .Z(n11635) );
  XNOR U11594 ( .A(n11641), .B(n11982), .Z(n11634) );
  XNOR U11595 ( .A(n11642), .B(n11643), .Z(n11982) );
  AND U11596 ( .A(n11983), .B(n11984), .Z(n11643) );
  NANDN U11597 ( .A(n11985), .B(n11986), .Z(n11984) );
  NANDN U11598 ( .A(n11987), .B(n11988), .Z(n11983) );
  NANDN U11599 ( .A(n11986), .B(n11985), .Z(n11988) );
  ANDN U11600 ( .B(\stack[1][16] ), .A(n6094), .Z(n11642) );
  XNOR U11601 ( .A(n11648), .B(n11989), .Z(n11641) );
  XNOR U11602 ( .A(n11649), .B(n11650), .Z(n11989) );
  AND U11603 ( .A(n11990), .B(n11991), .Z(n11650) );
  NAND U11604 ( .A(n11992), .B(n11993), .Z(n11991) );
  NANDN U11605 ( .A(n11994), .B(n11995), .Z(n11990) );
  OR U11606 ( .A(n11992), .B(n11993), .Z(n11995) );
  ANDN U11607 ( .B(\stack[1][17] ), .A(n6070), .Z(n11649) );
  XNOR U11608 ( .A(n11655), .B(n11996), .Z(n11648) );
  XNOR U11609 ( .A(n11656), .B(n11657), .Z(n11996) );
  AND U11610 ( .A(n11997), .B(n11998), .Z(n11657) );
  NANDN U11611 ( .A(n11999), .B(n12000), .Z(n11998) );
  NANDN U11612 ( .A(n12001), .B(n12002), .Z(n11997) );
  NANDN U11613 ( .A(n12000), .B(n11999), .Z(n12002) );
  ANDN U11614 ( .B(\stack[1][18] ), .A(n6046), .Z(n11656) );
  XNOR U11615 ( .A(n11662), .B(n12003), .Z(n11655) );
  XNOR U11616 ( .A(n11663), .B(n11664), .Z(n12003) );
  AND U11617 ( .A(n12004), .B(n12005), .Z(n11664) );
  NAND U11618 ( .A(n12006), .B(n12007), .Z(n12005) );
  NANDN U11619 ( .A(n12008), .B(n12009), .Z(n12004) );
  OR U11620 ( .A(n12006), .B(n12007), .Z(n12009) );
  ANDN U11621 ( .B(\stack[1][19] ), .A(n6022), .Z(n11663) );
  XNOR U11622 ( .A(n11669), .B(n12010), .Z(n11662) );
  XNOR U11623 ( .A(n11670), .B(n11671), .Z(n12010) );
  AND U11624 ( .A(n12011), .B(n12012), .Z(n11671) );
  NANDN U11625 ( .A(n12013), .B(n12014), .Z(n12012) );
  NANDN U11626 ( .A(n12015), .B(n12016), .Z(n12011) );
  NANDN U11627 ( .A(n12014), .B(n12013), .Z(n12016) );
  ANDN U11628 ( .B(\stack[1][20] ), .A(n5998), .Z(n11670) );
  XNOR U11629 ( .A(n11676), .B(n12017), .Z(n11669) );
  XNOR U11630 ( .A(n11677), .B(n11678), .Z(n12017) );
  AND U11631 ( .A(n12018), .B(n12019), .Z(n11678) );
  NAND U11632 ( .A(n12020), .B(n12021), .Z(n12019) );
  NANDN U11633 ( .A(n12022), .B(n12023), .Z(n12018) );
  OR U11634 ( .A(n12020), .B(n12021), .Z(n12023) );
  ANDN U11635 ( .B(\stack[1][21] ), .A(n5974), .Z(n11677) );
  XNOR U11636 ( .A(n11683), .B(n12024), .Z(n11676) );
  XNOR U11637 ( .A(n11684), .B(n11685), .Z(n12024) );
  AND U11638 ( .A(n12025), .B(n12026), .Z(n11685) );
  NANDN U11639 ( .A(n12027), .B(n12028), .Z(n12026) );
  NANDN U11640 ( .A(n12029), .B(n12030), .Z(n12025) );
  NANDN U11641 ( .A(n12028), .B(n12027), .Z(n12030) );
  ANDN U11642 ( .B(\stack[1][22] ), .A(n5950), .Z(n11684) );
  XNOR U11643 ( .A(n11690), .B(n12031), .Z(n11683) );
  XNOR U11644 ( .A(n11691), .B(n11692), .Z(n12031) );
  AND U11645 ( .A(n12032), .B(n12033), .Z(n11692) );
  NAND U11646 ( .A(n12034), .B(n12035), .Z(n12033) );
  NANDN U11647 ( .A(n12036), .B(n12037), .Z(n12032) );
  OR U11648 ( .A(n12034), .B(n12035), .Z(n12037) );
  ANDN U11649 ( .B(\stack[1][23] ), .A(n5926), .Z(n11691) );
  XNOR U11650 ( .A(n11697), .B(n12038), .Z(n11690) );
  XNOR U11651 ( .A(n11698), .B(n11699), .Z(n12038) );
  AND U11652 ( .A(n12039), .B(n12040), .Z(n11699) );
  NANDN U11653 ( .A(n12041), .B(n12042), .Z(n12040) );
  NANDN U11654 ( .A(n12043), .B(n12044), .Z(n12039) );
  NANDN U11655 ( .A(n12042), .B(n12041), .Z(n12044) );
  ANDN U11656 ( .B(\stack[1][24] ), .A(n5902), .Z(n11698) );
  XNOR U11657 ( .A(n11704), .B(n12045), .Z(n11697) );
  XNOR U11658 ( .A(n11705), .B(n11706), .Z(n12045) );
  AND U11659 ( .A(n12046), .B(n12047), .Z(n11706) );
  NAND U11660 ( .A(n12048), .B(n12049), .Z(n12047) );
  NANDN U11661 ( .A(n12050), .B(n12051), .Z(n12046) );
  OR U11662 ( .A(n12048), .B(n12049), .Z(n12051) );
  ANDN U11663 ( .B(\stack[1][25] ), .A(n5878), .Z(n11705) );
  XNOR U11664 ( .A(n11711), .B(n12052), .Z(n11704) );
  XNOR U11665 ( .A(n11712), .B(n11713), .Z(n12052) );
  AND U11666 ( .A(n12053), .B(n12054), .Z(n11713) );
  NANDN U11667 ( .A(n12055), .B(n12056), .Z(n12054) );
  NANDN U11668 ( .A(n12057), .B(n12058), .Z(n12053) );
  NANDN U11669 ( .A(n12056), .B(n12055), .Z(n12058) );
  ANDN U11670 ( .B(\stack[1][26] ), .A(n5854), .Z(n11712) );
  XNOR U11671 ( .A(n11718), .B(n12059), .Z(n11711) );
  XNOR U11672 ( .A(n11719), .B(n11720), .Z(n12059) );
  AND U11673 ( .A(n12060), .B(n12061), .Z(n11720) );
  NAND U11674 ( .A(n12062), .B(n12063), .Z(n12061) );
  NANDN U11675 ( .A(n12064), .B(n12065), .Z(n12060) );
  OR U11676 ( .A(n12062), .B(n12063), .Z(n12065) );
  ANDN U11677 ( .B(\stack[1][27] ), .A(n5830), .Z(n11719) );
  XNOR U11678 ( .A(n11725), .B(n12066), .Z(n11718) );
  XNOR U11679 ( .A(n11726), .B(n11727), .Z(n12066) );
  AND U11680 ( .A(n12067), .B(n12068), .Z(n11727) );
  NANDN U11681 ( .A(n12069), .B(n12070), .Z(n12068) );
  NANDN U11682 ( .A(n12071), .B(n12072), .Z(n12067) );
  NANDN U11683 ( .A(n12070), .B(n12069), .Z(n12072) );
  ANDN U11684 ( .B(\stack[1][28] ), .A(n5806), .Z(n11726) );
  XNOR U11685 ( .A(n11732), .B(n12073), .Z(n11725) );
  XNOR U11686 ( .A(n11733), .B(n11734), .Z(n12073) );
  AND U11687 ( .A(n12074), .B(n12075), .Z(n11734) );
  NAND U11688 ( .A(n12076), .B(n12077), .Z(n12075) );
  NANDN U11689 ( .A(n12078), .B(n12079), .Z(n12074) );
  OR U11690 ( .A(n12076), .B(n12077), .Z(n12079) );
  ANDN U11691 ( .B(\stack[1][29] ), .A(n5782), .Z(n11733) );
  XNOR U11692 ( .A(n11739), .B(n12080), .Z(n11732) );
  XNOR U11693 ( .A(n11740), .B(n11741), .Z(n12080) );
  AND U11694 ( .A(n12081), .B(n12082), .Z(n11741) );
  NANDN U11695 ( .A(n12083), .B(n12084), .Z(n12082) );
  NANDN U11696 ( .A(n12085), .B(n12086), .Z(n12081) );
  NANDN U11697 ( .A(n12084), .B(n12083), .Z(n12086) );
  ANDN U11698 ( .B(\stack[1][30] ), .A(n5758), .Z(n11740) );
  XNOR U11699 ( .A(n11746), .B(n12087), .Z(n11739) );
  XNOR U11700 ( .A(n11747), .B(n11748), .Z(n12087) );
  AND U11701 ( .A(n12088), .B(n12089), .Z(n11748) );
  NAND U11702 ( .A(n12090), .B(n12091), .Z(n12089) );
  NANDN U11703 ( .A(n12092), .B(n12093), .Z(n12088) );
  OR U11704 ( .A(n12090), .B(n12091), .Z(n12093) );
  ANDN U11705 ( .B(\stack[1][31] ), .A(n5734), .Z(n11747) );
  XNOR U11706 ( .A(n11753), .B(n12094), .Z(n11746) );
  XNOR U11707 ( .A(n11754), .B(n11755), .Z(n12094) );
  AND U11708 ( .A(n12095), .B(n12096), .Z(n11755) );
  NANDN U11709 ( .A(n12097), .B(n12098), .Z(n12096) );
  NANDN U11710 ( .A(n12099), .B(n12100), .Z(n12095) );
  NANDN U11711 ( .A(n12098), .B(n12097), .Z(n12100) );
  ANDN U11712 ( .B(\stack[1][32] ), .A(n5710), .Z(n11754) );
  XNOR U11713 ( .A(n11760), .B(n12101), .Z(n11753) );
  XNOR U11714 ( .A(n11761), .B(n11762), .Z(n12101) );
  AND U11715 ( .A(n12102), .B(n12103), .Z(n11762) );
  NAND U11716 ( .A(n12104), .B(n12105), .Z(n12103) );
  NANDN U11717 ( .A(n12106), .B(n12107), .Z(n12102) );
  OR U11718 ( .A(n12104), .B(n12105), .Z(n12107) );
  ANDN U11719 ( .B(\stack[1][33] ), .A(n5686), .Z(n11761) );
  XNOR U11720 ( .A(n11767), .B(n12108), .Z(n11760) );
  XNOR U11721 ( .A(n11768), .B(n11769), .Z(n12108) );
  AND U11722 ( .A(n12109), .B(n12110), .Z(n11769) );
  NANDN U11723 ( .A(n12111), .B(n12112), .Z(n12110) );
  NANDN U11724 ( .A(n12113), .B(n12114), .Z(n12109) );
  NANDN U11725 ( .A(n12112), .B(n12111), .Z(n12114) );
  ANDN U11726 ( .B(\stack[1][34] ), .A(n5662), .Z(n11768) );
  XNOR U11727 ( .A(n11774), .B(n12115), .Z(n11767) );
  XNOR U11728 ( .A(n11775), .B(n11776), .Z(n12115) );
  AND U11729 ( .A(n12116), .B(n12117), .Z(n11776) );
  NAND U11730 ( .A(n12118), .B(n12119), .Z(n12117) );
  NANDN U11731 ( .A(n12120), .B(n12121), .Z(n12116) );
  OR U11732 ( .A(n12118), .B(n12119), .Z(n12121) );
  ANDN U11733 ( .B(\stack[1][35] ), .A(n5638), .Z(n11775) );
  XNOR U11734 ( .A(n11781), .B(n12122), .Z(n11774) );
  XNOR U11735 ( .A(n11782), .B(n11783), .Z(n12122) );
  AND U11736 ( .A(n12123), .B(n12124), .Z(n11783) );
  NANDN U11737 ( .A(n12125), .B(n12126), .Z(n12124) );
  NANDN U11738 ( .A(n12127), .B(n12128), .Z(n12123) );
  NANDN U11739 ( .A(n12126), .B(n12125), .Z(n12128) );
  ANDN U11740 ( .B(\stack[1][36] ), .A(n5614), .Z(n11782) );
  XNOR U11741 ( .A(n11788), .B(n12129), .Z(n11781) );
  XOR U11742 ( .A(n11790), .B(n11791), .Z(n12129) );
  NAND U11743 ( .A(n12130), .B(n12131), .Z(n11791) );
  NAND U11744 ( .A(n12132), .B(n12133), .Z(n12131) );
  OR U11745 ( .A(n12134), .B(n12135), .Z(n12132) );
  AND U11746 ( .A(\stack[0][18] ), .B(\stack[1][37] ), .Z(n11790) );
  XNOR U11747 ( .A(n11797), .B(n12136), .Z(n11788) );
  XOR U11748 ( .A(n11798), .B(n11796), .Z(n12136) );
  AND U11749 ( .A(\stack[0][17] ), .B(\stack[1][38] ), .Z(n11796) );
  NAND U11750 ( .A(n12137), .B(n12138), .Z(n11798) );
  OR U11751 ( .A(n12139), .B(n12140), .Z(n12138) );
  NAND U11752 ( .A(n12141), .B(n12142), .Z(n12137) );
  NAND U11753 ( .A(n12140), .B(n12139), .Z(n12141) );
  XNOR U11754 ( .A(n11802), .B(n12143), .Z(n11797) );
  XNOR U11755 ( .A(n11803), .B(n11804), .Z(n12143) );
  AND U11756 ( .A(n12144), .B(n12145), .Z(n11804) );
  NAND U11757 ( .A(n12146), .B(n12147), .Z(n12145) );
  NANDN U11758 ( .A(n12148), .B(n12149), .Z(n12144) );
  OR U11759 ( .A(n12146), .B(n12147), .Z(n12149) );
  ANDN U11760 ( .B(\stack[1][39] ), .A(n5542), .Z(n11803) );
  XNOR U11761 ( .A(n11809), .B(n12150), .Z(n11802) );
  XNOR U11762 ( .A(n11810), .B(n11811), .Z(n12150) );
  AND U11763 ( .A(n12151), .B(n12152), .Z(n11811) );
  NANDN U11764 ( .A(n12153), .B(n12154), .Z(n12152) );
  NANDN U11765 ( .A(n12155), .B(n12156), .Z(n12151) );
  NANDN U11766 ( .A(n12154), .B(n12153), .Z(n12156) );
  ANDN U11767 ( .B(\stack[1][40] ), .A(n5518), .Z(n11810) );
  XNOR U11768 ( .A(n11816), .B(n12157), .Z(n11809) );
  XNOR U11769 ( .A(n11817), .B(n11818), .Z(n12157) );
  AND U11770 ( .A(n12158), .B(n12159), .Z(n11818) );
  NAND U11771 ( .A(n12160), .B(n12161), .Z(n12159) );
  NANDN U11772 ( .A(n12162), .B(n12163), .Z(n12158) );
  OR U11773 ( .A(n12160), .B(n12161), .Z(n12163) );
  ANDN U11774 ( .B(\stack[1][41] ), .A(n5494), .Z(n11817) );
  XNOR U11775 ( .A(n11823), .B(n12164), .Z(n11816) );
  XNOR U11776 ( .A(n11824), .B(n11825), .Z(n12164) );
  AND U11777 ( .A(n12165), .B(n12166), .Z(n11825) );
  NANDN U11778 ( .A(n12167), .B(n12168), .Z(n12166) );
  NANDN U11779 ( .A(n12169), .B(n12170), .Z(n12165) );
  NANDN U11780 ( .A(n12168), .B(n12167), .Z(n12170) );
  ANDN U11781 ( .B(\stack[1][42] ), .A(n5470), .Z(n11824) );
  XNOR U11782 ( .A(n11830), .B(n12171), .Z(n11823) );
  XNOR U11783 ( .A(n11831), .B(n11832), .Z(n12171) );
  AND U11784 ( .A(n12172), .B(n12173), .Z(n11832) );
  NAND U11785 ( .A(n12174), .B(n12175), .Z(n12173) );
  NANDN U11786 ( .A(n12176), .B(n12177), .Z(n12172) );
  OR U11787 ( .A(n12174), .B(n12175), .Z(n12177) );
  ANDN U11788 ( .B(\stack[1][43] ), .A(n5446), .Z(n11831) );
  XNOR U11789 ( .A(n11837), .B(n12178), .Z(n11830) );
  XNOR U11790 ( .A(n11838), .B(n11839), .Z(n12178) );
  AND U11791 ( .A(n12179), .B(n12180), .Z(n11839) );
  NANDN U11792 ( .A(n12181), .B(n12182), .Z(n12180) );
  NANDN U11793 ( .A(n12183), .B(n12184), .Z(n12179) );
  NANDN U11794 ( .A(n12182), .B(n12181), .Z(n12184) );
  ANDN U11795 ( .B(\stack[1][44] ), .A(n5422), .Z(n11838) );
  XNOR U11796 ( .A(n11844), .B(n12185), .Z(n11837) );
  XNOR U11797 ( .A(n11845), .B(n11846), .Z(n12185) );
  AND U11798 ( .A(n12186), .B(n12187), .Z(n11846) );
  NAND U11799 ( .A(n12188), .B(n12189), .Z(n12187) );
  NANDN U11800 ( .A(n12190), .B(n12191), .Z(n12186) );
  OR U11801 ( .A(n12188), .B(n12189), .Z(n12191) );
  ANDN U11802 ( .B(\stack[1][45] ), .A(n5398), .Z(n11845) );
  XNOR U11803 ( .A(n11851), .B(n12192), .Z(n11844) );
  XNOR U11804 ( .A(n11852), .B(n11853), .Z(n12192) );
  AND U11805 ( .A(n12193), .B(n12194), .Z(n11853) );
  NANDN U11806 ( .A(n12195), .B(n12196), .Z(n12194) );
  NANDN U11807 ( .A(n12197), .B(n12198), .Z(n12193) );
  NANDN U11808 ( .A(n12196), .B(n12195), .Z(n12198) );
  ANDN U11809 ( .B(\stack[1][46] ), .A(n5374), .Z(n11852) );
  XNOR U11810 ( .A(n11858), .B(n12199), .Z(n11851) );
  XNOR U11811 ( .A(n11859), .B(n11860), .Z(n12199) );
  AND U11812 ( .A(n12200), .B(n12201), .Z(n11860) );
  NAND U11813 ( .A(n12202), .B(n12203), .Z(n12201) );
  NANDN U11814 ( .A(n12204), .B(n12205), .Z(n12200) );
  OR U11815 ( .A(n12202), .B(n12203), .Z(n12205) );
  ANDN U11816 ( .B(\stack[1][47] ), .A(n5350), .Z(n11859) );
  XNOR U11817 ( .A(n11865), .B(n12206), .Z(n11858) );
  XNOR U11818 ( .A(n11866), .B(n11867), .Z(n12206) );
  AND U11819 ( .A(n12207), .B(n12208), .Z(n11867) );
  NANDN U11820 ( .A(n12209), .B(n12210), .Z(n12208) );
  NANDN U11821 ( .A(n12211), .B(n12212), .Z(n12207) );
  NANDN U11822 ( .A(n12210), .B(n12209), .Z(n12212) );
  ANDN U11823 ( .B(\stack[1][48] ), .A(n5326), .Z(n11866) );
  XNOR U11824 ( .A(n11872), .B(n12213), .Z(n11865) );
  XNOR U11825 ( .A(n11873), .B(n11874), .Z(n12213) );
  AND U11826 ( .A(n12214), .B(n12215), .Z(n11874) );
  NAND U11827 ( .A(n12216), .B(n12217), .Z(n12215) );
  NANDN U11828 ( .A(n12218), .B(n12219), .Z(n12214) );
  OR U11829 ( .A(n12216), .B(n12217), .Z(n12219) );
  ANDN U11830 ( .B(\stack[1][49] ), .A(n5302), .Z(n11873) );
  XNOR U11831 ( .A(n11879), .B(n12220), .Z(n11872) );
  XNOR U11832 ( .A(n11880), .B(n11881), .Z(n12220) );
  AND U11833 ( .A(n12221), .B(n12222), .Z(n11881) );
  NANDN U11834 ( .A(n12223), .B(n12224), .Z(n12222) );
  NANDN U11835 ( .A(n12225), .B(n12226), .Z(n12221) );
  NANDN U11836 ( .A(n12224), .B(n12223), .Z(n12226) );
  ANDN U11837 ( .B(\stack[1][50] ), .A(n5278), .Z(n11880) );
  XNOR U11838 ( .A(n11886), .B(n12227), .Z(n11879) );
  XNOR U11839 ( .A(n11887), .B(n11888), .Z(n12227) );
  AND U11840 ( .A(n12228), .B(n12229), .Z(n11888) );
  NAND U11841 ( .A(n12230), .B(n12231), .Z(n12229) );
  NANDN U11842 ( .A(n12232), .B(n12233), .Z(n12228) );
  OR U11843 ( .A(n12230), .B(n12231), .Z(n12233) );
  ANDN U11844 ( .B(\stack[1][51] ), .A(n5254), .Z(n11887) );
  XNOR U11845 ( .A(n11893), .B(n12234), .Z(n11886) );
  XNOR U11846 ( .A(n11894), .B(n11895), .Z(n12234) );
  AND U11847 ( .A(n12235), .B(n12236), .Z(n11895) );
  NAND U11848 ( .A(n12237), .B(n12238), .Z(n12236) );
  NAND U11849 ( .A(n12239), .B(n12240), .Z(n12235) );
  OR U11850 ( .A(n12237), .B(n12238), .Z(n12239) );
  ANDN U11851 ( .B(\stack[1][52] ), .A(n5230), .Z(n11894) );
  XNOR U11852 ( .A(n11900), .B(n12241), .Z(n11893) );
  XNOR U11853 ( .A(n11901), .B(n11903), .Z(n12241) );
  ANDN U11854 ( .B(n12242), .A(n12243), .Z(n11903) );
  ANDN U11855 ( .B(\stack[0][0] ), .A(n6468), .Z(n12242) );
  ANDN U11856 ( .B(\stack[1][53] ), .A(n5206), .Z(n11901) );
  XOR U11857 ( .A(n11906), .B(n12244), .Z(n11900) );
  NANDN U11858 ( .A(n5160), .B(\stack[1][55] ), .Z(n12244) );
  NANDN U11859 ( .A(n6468), .B(\stack[0][1] ), .Z(n11906) );
  ANDN U11860 ( .B(\stack[1][5] ), .A(n6358), .Z(n9013) );
  AND U11861 ( .A(n12245), .B(n12246), .Z(n9014) );
  NANDN U11862 ( .A(n9018), .B(n9020), .Z(n12246) );
  NANDN U11863 ( .A(n9021), .B(n12247), .Z(n12245) );
  NANDN U11864 ( .A(n9020), .B(n9018), .Z(n12247) );
  XOR U11865 ( .A(n11915), .B(n12248), .Z(n9018) );
  XNOR U11866 ( .A(n11916), .B(n11917), .Z(n12248) );
  AND U11867 ( .A(n12249), .B(n12250), .Z(n11917) );
  NAND U11868 ( .A(n12251), .B(n12252), .Z(n12250) );
  NANDN U11869 ( .A(n12253), .B(n12254), .Z(n12249) );
  OR U11870 ( .A(n12251), .B(n12252), .Z(n12254) );
  ANDN U11871 ( .B(\stack[0][48] ), .A(n5316), .Z(n11916) );
  XNOR U11872 ( .A(n11922), .B(n12255), .Z(n11915) );
  XNOR U11873 ( .A(n11923), .B(n11924), .Z(n12255) );
  AND U11874 ( .A(n12256), .B(n12257), .Z(n11924) );
  NANDN U11875 ( .A(n12258), .B(n12259), .Z(n12257) );
  NANDN U11876 ( .A(n12260), .B(n12261), .Z(n12256) );
  NANDN U11877 ( .A(n12259), .B(n12258), .Z(n12261) );
  ANDN U11878 ( .B(\stack[0][47] ), .A(n5340), .Z(n11923) );
  XNOR U11879 ( .A(n11929), .B(n12262), .Z(n11922) );
  XNOR U11880 ( .A(n11930), .B(n11931), .Z(n12262) );
  AND U11881 ( .A(n12263), .B(n12264), .Z(n11931) );
  NAND U11882 ( .A(n12265), .B(n12266), .Z(n12264) );
  NANDN U11883 ( .A(n12267), .B(n12268), .Z(n12263) );
  OR U11884 ( .A(n12265), .B(n12266), .Z(n12268) );
  ANDN U11885 ( .B(\stack[0][46] ), .A(n5364), .Z(n11930) );
  XNOR U11886 ( .A(n11936), .B(n12269), .Z(n11929) );
  XNOR U11887 ( .A(n11937), .B(n11938), .Z(n12269) );
  AND U11888 ( .A(n12270), .B(n12271), .Z(n11938) );
  NANDN U11889 ( .A(n12272), .B(n12273), .Z(n12271) );
  NANDN U11890 ( .A(n12274), .B(n12275), .Z(n12270) );
  NANDN U11891 ( .A(n12273), .B(n12272), .Z(n12275) );
  ANDN U11892 ( .B(\stack[0][45] ), .A(n5387), .Z(n11937) );
  XNOR U11893 ( .A(n11943), .B(n12276), .Z(n11936) );
  XNOR U11894 ( .A(n11944), .B(n11945), .Z(n12276) );
  AND U11895 ( .A(n12277), .B(n12278), .Z(n11945) );
  NAND U11896 ( .A(n12279), .B(n12280), .Z(n12278) );
  NANDN U11897 ( .A(n12281), .B(n12282), .Z(n12277) );
  OR U11898 ( .A(n12279), .B(n12280), .Z(n12282) );
  ANDN U11899 ( .B(\stack[1][10] ), .A(n6214), .Z(n11944) );
  XNOR U11900 ( .A(n11950), .B(n12283), .Z(n11943) );
  XNOR U11901 ( .A(n11951), .B(n11952), .Z(n12283) );
  AND U11902 ( .A(n12284), .B(n12285), .Z(n11952) );
  NANDN U11903 ( .A(n12286), .B(n12287), .Z(n12285) );
  NANDN U11904 ( .A(n12288), .B(n12289), .Z(n12284) );
  NANDN U11905 ( .A(n12287), .B(n12286), .Z(n12289) );
  ANDN U11906 ( .B(\stack[1][11] ), .A(n6190), .Z(n11951) );
  XNOR U11907 ( .A(n11957), .B(n12290), .Z(n11950) );
  XNOR U11908 ( .A(n11958), .B(n11959), .Z(n12290) );
  AND U11909 ( .A(n12291), .B(n12292), .Z(n11959) );
  NAND U11910 ( .A(n12293), .B(n12294), .Z(n12292) );
  NANDN U11911 ( .A(n12295), .B(n12296), .Z(n12291) );
  OR U11912 ( .A(n12293), .B(n12294), .Z(n12296) );
  ANDN U11913 ( .B(\stack[1][12] ), .A(n6166), .Z(n11958) );
  XNOR U11914 ( .A(n11964), .B(n12297), .Z(n11957) );
  XNOR U11915 ( .A(n11965), .B(n11966), .Z(n12297) );
  AND U11916 ( .A(n12298), .B(n12299), .Z(n11966) );
  NANDN U11917 ( .A(n12300), .B(n12301), .Z(n12299) );
  NANDN U11918 ( .A(n12302), .B(n12303), .Z(n12298) );
  NANDN U11919 ( .A(n12301), .B(n12300), .Z(n12303) );
  ANDN U11920 ( .B(\stack[1][13] ), .A(n6142), .Z(n11965) );
  XNOR U11921 ( .A(n11971), .B(n12304), .Z(n11964) );
  XNOR U11922 ( .A(n11972), .B(n11973), .Z(n12304) );
  AND U11923 ( .A(n12305), .B(n12306), .Z(n11973) );
  NAND U11924 ( .A(n12307), .B(n12308), .Z(n12306) );
  NANDN U11925 ( .A(n12309), .B(n12310), .Z(n12305) );
  OR U11926 ( .A(n12307), .B(n12308), .Z(n12310) );
  ANDN U11927 ( .B(\stack[1][14] ), .A(n6118), .Z(n11972) );
  XNOR U11928 ( .A(n11978), .B(n12311), .Z(n11971) );
  XNOR U11929 ( .A(n11979), .B(n11980), .Z(n12311) );
  AND U11930 ( .A(n12312), .B(n12313), .Z(n11980) );
  NANDN U11931 ( .A(n12314), .B(n12315), .Z(n12313) );
  NANDN U11932 ( .A(n12316), .B(n12317), .Z(n12312) );
  NANDN U11933 ( .A(n12315), .B(n12314), .Z(n12317) );
  ANDN U11934 ( .B(\stack[1][15] ), .A(n6094), .Z(n11979) );
  XNOR U11935 ( .A(n11985), .B(n12318), .Z(n11978) );
  XNOR U11936 ( .A(n11986), .B(n11987), .Z(n12318) );
  AND U11937 ( .A(n12319), .B(n12320), .Z(n11987) );
  NAND U11938 ( .A(n12321), .B(n12322), .Z(n12320) );
  NANDN U11939 ( .A(n12323), .B(n12324), .Z(n12319) );
  OR U11940 ( .A(n12321), .B(n12322), .Z(n12324) );
  ANDN U11941 ( .B(\stack[1][16] ), .A(n6070), .Z(n11986) );
  XNOR U11942 ( .A(n11992), .B(n12325), .Z(n11985) );
  XNOR U11943 ( .A(n11993), .B(n11994), .Z(n12325) );
  AND U11944 ( .A(n12326), .B(n12327), .Z(n11994) );
  NANDN U11945 ( .A(n12328), .B(n12329), .Z(n12327) );
  NANDN U11946 ( .A(n12330), .B(n12331), .Z(n12326) );
  NANDN U11947 ( .A(n12329), .B(n12328), .Z(n12331) );
  ANDN U11948 ( .B(\stack[1][17] ), .A(n6046), .Z(n11993) );
  XNOR U11949 ( .A(n11999), .B(n12332), .Z(n11992) );
  XNOR U11950 ( .A(n12000), .B(n12001), .Z(n12332) );
  AND U11951 ( .A(n12333), .B(n12334), .Z(n12001) );
  NAND U11952 ( .A(n12335), .B(n12336), .Z(n12334) );
  NANDN U11953 ( .A(n12337), .B(n12338), .Z(n12333) );
  OR U11954 ( .A(n12335), .B(n12336), .Z(n12338) );
  ANDN U11955 ( .B(\stack[1][18] ), .A(n6022), .Z(n12000) );
  XNOR U11956 ( .A(n12006), .B(n12339), .Z(n11999) );
  XNOR U11957 ( .A(n12007), .B(n12008), .Z(n12339) );
  AND U11958 ( .A(n12340), .B(n12341), .Z(n12008) );
  NANDN U11959 ( .A(n12342), .B(n12343), .Z(n12341) );
  NANDN U11960 ( .A(n12344), .B(n12345), .Z(n12340) );
  NANDN U11961 ( .A(n12343), .B(n12342), .Z(n12345) );
  ANDN U11962 ( .B(\stack[1][19] ), .A(n5998), .Z(n12007) );
  XNOR U11963 ( .A(n12013), .B(n12346), .Z(n12006) );
  XNOR U11964 ( .A(n12014), .B(n12015), .Z(n12346) );
  AND U11965 ( .A(n12347), .B(n12348), .Z(n12015) );
  NAND U11966 ( .A(n12349), .B(n12350), .Z(n12348) );
  NANDN U11967 ( .A(n12351), .B(n12352), .Z(n12347) );
  OR U11968 ( .A(n12349), .B(n12350), .Z(n12352) );
  ANDN U11969 ( .B(\stack[1][20] ), .A(n5974), .Z(n12014) );
  XNOR U11970 ( .A(n12020), .B(n12353), .Z(n12013) );
  XNOR U11971 ( .A(n12021), .B(n12022), .Z(n12353) );
  AND U11972 ( .A(n12354), .B(n12355), .Z(n12022) );
  NANDN U11973 ( .A(n12356), .B(n12357), .Z(n12355) );
  NANDN U11974 ( .A(n12358), .B(n12359), .Z(n12354) );
  NANDN U11975 ( .A(n12357), .B(n12356), .Z(n12359) );
  ANDN U11976 ( .B(\stack[1][21] ), .A(n5950), .Z(n12021) );
  XNOR U11977 ( .A(n12027), .B(n12360), .Z(n12020) );
  XNOR U11978 ( .A(n12028), .B(n12029), .Z(n12360) );
  AND U11979 ( .A(n12361), .B(n12362), .Z(n12029) );
  NAND U11980 ( .A(n12363), .B(n12364), .Z(n12362) );
  NANDN U11981 ( .A(n12365), .B(n12366), .Z(n12361) );
  OR U11982 ( .A(n12363), .B(n12364), .Z(n12366) );
  ANDN U11983 ( .B(\stack[1][22] ), .A(n5926), .Z(n12028) );
  XNOR U11984 ( .A(n12034), .B(n12367), .Z(n12027) );
  XNOR U11985 ( .A(n12035), .B(n12036), .Z(n12367) );
  AND U11986 ( .A(n12368), .B(n12369), .Z(n12036) );
  NANDN U11987 ( .A(n12370), .B(n12371), .Z(n12369) );
  NANDN U11988 ( .A(n12372), .B(n12373), .Z(n12368) );
  NANDN U11989 ( .A(n12371), .B(n12370), .Z(n12373) );
  ANDN U11990 ( .B(\stack[1][23] ), .A(n5902), .Z(n12035) );
  XNOR U11991 ( .A(n12041), .B(n12374), .Z(n12034) );
  XNOR U11992 ( .A(n12042), .B(n12043), .Z(n12374) );
  AND U11993 ( .A(n12375), .B(n12376), .Z(n12043) );
  NAND U11994 ( .A(n12377), .B(n12378), .Z(n12376) );
  NANDN U11995 ( .A(n12379), .B(n12380), .Z(n12375) );
  OR U11996 ( .A(n12377), .B(n12378), .Z(n12380) );
  ANDN U11997 ( .B(\stack[1][24] ), .A(n5878), .Z(n12042) );
  XNOR U11998 ( .A(n12048), .B(n12381), .Z(n12041) );
  XNOR U11999 ( .A(n12049), .B(n12050), .Z(n12381) );
  AND U12000 ( .A(n12382), .B(n12383), .Z(n12050) );
  NANDN U12001 ( .A(n12384), .B(n12385), .Z(n12383) );
  NANDN U12002 ( .A(n12386), .B(n12387), .Z(n12382) );
  NANDN U12003 ( .A(n12385), .B(n12384), .Z(n12387) );
  ANDN U12004 ( .B(\stack[1][25] ), .A(n5854), .Z(n12049) );
  XNOR U12005 ( .A(n12055), .B(n12388), .Z(n12048) );
  XNOR U12006 ( .A(n12056), .B(n12057), .Z(n12388) );
  AND U12007 ( .A(n12389), .B(n12390), .Z(n12057) );
  NAND U12008 ( .A(n12391), .B(n12392), .Z(n12390) );
  NANDN U12009 ( .A(n12393), .B(n12394), .Z(n12389) );
  OR U12010 ( .A(n12391), .B(n12392), .Z(n12394) );
  ANDN U12011 ( .B(\stack[1][26] ), .A(n5830), .Z(n12056) );
  XNOR U12012 ( .A(n12062), .B(n12395), .Z(n12055) );
  XNOR U12013 ( .A(n12063), .B(n12064), .Z(n12395) );
  AND U12014 ( .A(n12396), .B(n12397), .Z(n12064) );
  NANDN U12015 ( .A(n12398), .B(n12399), .Z(n12397) );
  NANDN U12016 ( .A(n12400), .B(n12401), .Z(n12396) );
  NANDN U12017 ( .A(n12399), .B(n12398), .Z(n12401) );
  ANDN U12018 ( .B(\stack[1][27] ), .A(n5806), .Z(n12063) );
  XNOR U12019 ( .A(n12069), .B(n12402), .Z(n12062) );
  XNOR U12020 ( .A(n12070), .B(n12071), .Z(n12402) );
  AND U12021 ( .A(n12403), .B(n12404), .Z(n12071) );
  NAND U12022 ( .A(n12405), .B(n12406), .Z(n12404) );
  NANDN U12023 ( .A(n12407), .B(n12408), .Z(n12403) );
  OR U12024 ( .A(n12405), .B(n12406), .Z(n12408) );
  ANDN U12025 ( .B(\stack[1][28] ), .A(n5782), .Z(n12070) );
  XNOR U12026 ( .A(n12076), .B(n12409), .Z(n12069) );
  XNOR U12027 ( .A(n12077), .B(n12078), .Z(n12409) );
  AND U12028 ( .A(n12410), .B(n12411), .Z(n12078) );
  NANDN U12029 ( .A(n12412), .B(n12413), .Z(n12411) );
  NANDN U12030 ( .A(n12414), .B(n12415), .Z(n12410) );
  NANDN U12031 ( .A(n12413), .B(n12412), .Z(n12415) );
  ANDN U12032 ( .B(\stack[1][29] ), .A(n5758), .Z(n12077) );
  XNOR U12033 ( .A(n12083), .B(n12416), .Z(n12076) );
  XNOR U12034 ( .A(n12084), .B(n12085), .Z(n12416) );
  AND U12035 ( .A(n12417), .B(n12418), .Z(n12085) );
  NAND U12036 ( .A(n12419), .B(n12420), .Z(n12418) );
  NANDN U12037 ( .A(n12421), .B(n12422), .Z(n12417) );
  OR U12038 ( .A(n12419), .B(n12420), .Z(n12422) );
  ANDN U12039 ( .B(\stack[1][30] ), .A(n5734), .Z(n12084) );
  XNOR U12040 ( .A(n12090), .B(n12423), .Z(n12083) );
  XNOR U12041 ( .A(n12091), .B(n12092), .Z(n12423) );
  AND U12042 ( .A(n12424), .B(n12425), .Z(n12092) );
  NANDN U12043 ( .A(n12426), .B(n12427), .Z(n12425) );
  NANDN U12044 ( .A(n12428), .B(n12429), .Z(n12424) );
  NANDN U12045 ( .A(n12427), .B(n12426), .Z(n12429) );
  ANDN U12046 ( .B(\stack[1][31] ), .A(n5710), .Z(n12091) );
  XNOR U12047 ( .A(n12097), .B(n12430), .Z(n12090) );
  XNOR U12048 ( .A(n12098), .B(n12099), .Z(n12430) );
  AND U12049 ( .A(n12431), .B(n12432), .Z(n12099) );
  NAND U12050 ( .A(n12433), .B(n12434), .Z(n12432) );
  NANDN U12051 ( .A(n12435), .B(n12436), .Z(n12431) );
  OR U12052 ( .A(n12433), .B(n12434), .Z(n12436) );
  ANDN U12053 ( .B(\stack[1][32] ), .A(n5686), .Z(n12098) );
  XNOR U12054 ( .A(n12104), .B(n12437), .Z(n12097) );
  XNOR U12055 ( .A(n12105), .B(n12106), .Z(n12437) );
  AND U12056 ( .A(n12438), .B(n12439), .Z(n12106) );
  NANDN U12057 ( .A(n12440), .B(n12441), .Z(n12439) );
  NANDN U12058 ( .A(n12442), .B(n12443), .Z(n12438) );
  NANDN U12059 ( .A(n12441), .B(n12440), .Z(n12443) );
  ANDN U12060 ( .B(\stack[1][33] ), .A(n5662), .Z(n12105) );
  XNOR U12061 ( .A(n12111), .B(n12444), .Z(n12104) );
  XNOR U12062 ( .A(n12112), .B(n12113), .Z(n12444) );
  AND U12063 ( .A(n12445), .B(n12446), .Z(n12113) );
  NAND U12064 ( .A(n12447), .B(n12448), .Z(n12446) );
  NANDN U12065 ( .A(n12449), .B(n12450), .Z(n12445) );
  OR U12066 ( .A(n12447), .B(n12448), .Z(n12450) );
  ANDN U12067 ( .B(\stack[1][34] ), .A(n5638), .Z(n12112) );
  XNOR U12068 ( .A(n12118), .B(n12451), .Z(n12111) );
  XNOR U12069 ( .A(n12119), .B(n12120), .Z(n12451) );
  AND U12070 ( .A(n12452), .B(n12453), .Z(n12120) );
  NANDN U12071 ( .A(n12454), .B(n12455), .Z(n12453) );
  NANDN U12072 ( .A(n12456), .B(n12457), .Z(n12452) );
  NANDN U12073 ( .A(n12455), .B(n12454), .Z(n12457) );
  ANDN U12074 ( .B(\stack[1][35] ), .A(n5614), .Z(n12119) );
  XNOR U12075 ( .A(n12125), .B(n12458), .Z(n12118) );
  XNOR U12076 ( .A(n12126), .B(n12127), .Z(n12458) );
  AND U12077 ( .A(n12459), .B(n12460), .Z(n12127) );
  NAND U12078 ( .A(n12461), .B(n12462), .Z(n12460) );
  NANDN U12079 ( .A(n12463), .B(n12464), .Z(n12459) );
  OR U12080 ( .A(n12461), .B(n12462), .Z(n12464) );
  ANDN U12081 ( .B(\stack[1][36] ), .A(n5590), .Z(n12126) );
  XNOR U12082 ( .A(n12133), .B(n12465), .Z(n12125) );
  XOR U12083 ( .A(n12134), .B(n12135), .Z(n12465) );
  NAND U12084 ( .A(n12466), .B(n12467), .Z(n12135) );
  NANDN U12085 ( .A(n12468), .B(n12469), .Z(n12467) );
  OR U12086 ( .A(n12470), .B(n12471), .Z(n12469) );
  AND U12087 ( .A(\stack[0][17] ), .B(\stack[1][37] ), .Z(n12134) );
  XNOR U12088 ( .A(n12140), .B(n12472), .Z(n12133) );
  XNOR U12089 ( .A(n12139), .B(n12142), .Z(n12472) );
  AND U12090 ( .A(\stack[0][16] ), .B(\stack[1][38] ), .Z(n12142) );
  AND U12091 ( .A(n12473), .B(n12474), .Z(n12139) );
  NAND U12092 ( .A(n12475), .B(n12476), .Z(n12474) );
  OR U12093 ( .A(n12477), .B(n12478), .Z(n12475) );
  XNOR U12094 ( .A(n12146), .B(n12479), .Z(n12140) );
  XNOR U12095 ( .A(n12147), .B(n12148), .Z(n12479) );
  AND U12096 ( .A(n12480), .B(n12481), .Z(n12148) );
  NANDN U12097 ( .A(n12482), .B(n12483), .Z(n12481) );
  NANDN U12098 ( .A(n12484), .B(n12485), .Z(n12480) );
  NANDN U12099 ( .A(n12483), .B(n12482), .Z(n12485) );
  ANDN U12100 ( .B(\stack[1][39] ), .A(n5518), .Z(n12147) );
  XNOR U12101 ( .A(n12153), .B(n12486), .Z(n12146) );
  XNOR U12102 ( .A(n12154), .B(n12155), .Z(n12486) );
  AND U12103 ( .A(n12487), .B(n12488), .Z(n12155) );
  NAND U12104 ( .A(n12489), .B(n12490), .Z(n12488) );
  NANDN U12105 ( .A(n12491), .B(n12492), .Z(n12487) );
  OR U12106 ( .A(n12489), .B(n12490), .Z(n12492) );
  ANDN U12107 ( .B(\stack[1][40] ), .A(n5494), .Z(n12154) );
  XNOR U12108 ( .A(n12160), .B(n12493), .Z(n12153) );
  XNOR U12109 ( .A(n12161), .B(n12162), .Z(n12493) );
  AND U12110 ( .A(n12494), .B(n12495), .Z(n12162) );
  NANDN U12111 ( .A(n12496), .B(n12497), .Z(n12495) );
  NANDN U12112 ( .A(n12498), .B(n12499), .Z(n12494) );
  NANDN U12113 ( .A(n12497), .B(n12496), .Z(n12499) );
  ANDN U12114 ( .B(\stack[1][41] ), .A(n5470), .Z(n12161) );
  XNOR U12115 ( .A(n12167), .B(n12500), .Z(n12160) );
  XNOR U12116 ( .A(n12168), .B(n12169), .Z(n12500) );
  AND U12117 ( .A(n12501), .B(n12502), .Z(n12169) );
  NAND U12118 ( .A(n12503), .B(n12504), .Z(n12502) );
  NANDN U12119 ( .A(n12505), .B(n12506), .Z(n12501) );
  OR U12120 ( .A(n12503), .B(n12504), .Z(n12506) );
  ANDN U12121 ( .B(\stack[1][42] ), .A(n5446), .Z(n12168) );
  XNOR U12122 ( .A(n12174), .B(n12507), .Z(n12167) );
  XNOR U12123 ( .A(n12175), .B(n12176), .Z(n12507) );
  AND U12124 ( .A(n12508), .B(n12509), .Z(n12176) );
  NANDN U12125 ( .A(n12510), .B(n12511), .Z(n12509) );
  NANDN U12126 ( .A(n12512), .B(n12513), .Z(n12508) );
  NANDN U12127 ( .A(n12511), .B(n12510), .Z(n12513) );
  ANDN U12128 ( .B(\stack[1][43] ), .A(n5422), .Z(n12175) );
  XNOR U12129 ( .A(n12181), .B(n12514), .Z(n12174) );
  XNOR U12130 ( .A(n12182), .B(n12183), .Z(n12514) );
  AND U12131 ( .A(n12515), .B(n12516), .Z(n12183) );
  NAND U12132 ( .A(n12517), .B(n12518), .Z(n12516) );
  NANDN U12133 ( .A(n12519), .B(n12520), .Z(n12515) );
  OR U12134 ( .A(n12517), .B(n12518), .Z(n12520) );
  ANDN U12135 ( .B(\stack[1][44] ), .A(n5398), .Z(n12182) );
  XNOR U12136 ( .A(n12188), .B(n12521), .Z(n12181) );
  XNOR U12137 ( .A(n12189), .B(n12190), .Z(n12521) );
  AND U12138 ( .A(n12522), .B(n12523), .Z(n12190) );
  NANDN U12139 ( .A(n12524), .B(n12525), .Z(n12523) );
  NANDN U12140 ( .A(n12526), .B(n12527), .Z(n12522) );
  NANDN U12141 ( .A(n12525), .B(n12524), .Z(n12527) );
  ANDN U12142 ( .B(\stack[1][45] ), .A(n5374), .Z(n12189) );
  XNOR U12143 ( .A(n12195), .B(n12528), .Z(n12188) );
  XNOR U12144 ( .A(n12196), .B(n12197), .Z(n12528) );
  AND U12145 ( .A(n12529), .B(n12530), .Z(n12197) );
  NAND U12146 ( .A(n12531), .B(n12532), .Z(n12530) );
  NANDN U12147 ( .A(n12533), .B(n12534), .Z(n12529) );
  OR U12148 ( .A(n12531), .B(n12532), .Z(n12534) );
  ANDN U12149 ( .B(\stack[1][46] ), .A(n5350), .Z(n12196) );
  XNOR U12150 ( .A(n12202), .B(n12535), .Z(n12195) );
  XNOR U12151 ( .A(n12203), .B(n12204), .Z(n12535) );
  AND U12152 ( .A(n12536), .B(n12537), .Z(n12204) );
  NANDN U12153 ( .A(n12538), .B(n12539), .Z(n12537) );
  NANDN U12154 ( .A(n12540), .B(n12541), .Z(n12536) );
  NANDN U12155 ( .A(n12539), .B(n12538), .Z(n12541) );
  ANDN U12156 ( .B(\stack[1][47] ), .A(n5326), .Z(n12203) );
  XNOR U12157 ( .A(n12209), .B(n12542), .Z(n12202) );
  XNOR U12158 ( .A(n12210), .B(n12211), .Z(n12542) );
  AND U12159 ( .A(n12543), .B(n12544), .Z(n12211) );
  NAND U12160 ( .A(n12545), .B(n12546), .Z(n12544) );
  NANDN U12161 ( .A(n12547), .B(n12548), .Z(n12543) );
  OR U12162 ( .A(n12545), .B(n12546), .Z(n12548) );
  ANDN U12163 ( .B(\stack[1][48] ), .A(n5302), .Z(n12210) );
  XNOR U12164 ( .A(n12216), .B(n12549), .Z(n12209) );
  XNOR U12165 ( .A(n12217), .B(n12218), .Z(n12549) );
  AND U12166 ( .A(n12550), .B(n12551), .Z(n12218) );
  NANDN U12167 ( .A(n12552), .B(n12553), .Z(n12551) );
  NANDN U12168 ( .A(n12554), .B(n12555), .Z(n12550) );
  NANDN U12169 ( .A(n12553), .B(n12552), .Z(n12555) );
  ANDN U12170 ( .B(\stack[1][49] ), .A(n5278), .Z(n12217) );
  XNOR U12171 ( .A(n12223), .B(n12556), .Z(n12216) );
  XNOR U12172 ( .A(n12224), .B(n12225), .Z(n12556) );
  AND U12173 ( .A(n12557), .B(n12558), .Z(n12225) );
  NAND U12174 ( .A(n12559), .B(n12560), .Z(n12558) );
  NANDN U12175 ( .A(n12561), .B(n12562), .Z(n12557) );
  OR U12176 ( .A(n12559), .B(n12560), .Z(n12562) );
  ANDN U12177 ( .B(\stack[1][50] ), .A(n5254), .Z(n12224) );
  XNOR U12178 ( .A(n12230), .B(n12563), .Z(n12223) );
  XNOR U12179 ( .A(n12231), .B(n12232), .Z(n12563) );
  AND U12180 ( .A(n12564), .B(n12565), .Z(n12232) );
  NAND U12181 ( .A(n12566), .B(n12567), .Z(n12565) );
  NAND U12182 ( .A(n12568), .B(n12569), .Z(n12564) );
  OR U12183 ( .A(n12566), .B(n12567), .Z(n12568) );
  ANDN U12184 ( .B(\stack[1][51] ), .A(n5230), .Z(n12231) );
  XNOR U12185 ( .A(n12237), .B(n12570), .Z(n12230) );
  XNOR U12186 ( .A(n12238), .B(n12240), .Z(n12570) );
  ANDN U12187 ( .B(n12571), .A(n12572), .Z(n12240) );
  ANDN U12188 ( .B(\stack[0][0] ), .A(n6444), .Z(n12571) );
  ANDN U12189 ( .B(\stack[1][52] ), .A(n5206), .Z(n12238) );
  XOR U12190 ( .A(n12243), .B(n12573), .Z(n12237) );
  NANDN U12191 ( .A(n5160), .B(\stack[1][54] ), .Z(n12573) );
  NANDN U12192 ( .A(n6444), .B(\stack[0][1] ), .Z(n12243) );
  ANDN U12193 ( .B(\stack[0][49] ), .A(n5292), .Z(n9020) );
  AND U12194 ( .A(n12574), .B(n12575), .Z(n9021) );
  NANDN U12195 ( .A(n9028), .B(n12576), .Z(n12574) );
  NANDN U12196 ( .A(n9027), .B(n9025), .Z(n12576) );
  XNOR U12197 ( .A(n12251), .B(n12577), .Z(n9025) );
  XNOR U12198 ( .A(n12252), .B(n12253), .Z(n12577) );
  AND U12199 ( .A(n12578), .B(n12579), .Z(n12253) );
  NANDN U12200 ( .A(n12580), .B(n12581), .Z(n12579) );
  NANDN U12201 ( .A(n12582), .B(n12583), .Z(n12578) );
  NANDN U12202 ( .A(n12581), .B(n12580), .Z(n12583) );
  ANDN U12203 ( .B(\stack[0][47] ), .A(n5316), .Z(n12252) );
  XNOR U12204 ( .A(n12258), .B(n12584), .Z(n12251) );
  XNOR U12205 ( .A(n12259), .B(n12260), .Z(n12584) );
  AND U12206 ( .A(n12585), .B(n12586), .Z(n12260) );
  NAND U12207 ( .A(n12587), .B(n12588), .Z(n12586) );
  NANDN U12208 ( .A(n12589), .B(n12590), .Z(n12585) );
  OR U12209 ( .A(n12587), .B(n12588), .Z(n12590) );
  ANDN U12210 ( .B(\stack[0][46] ), .A(n5340), .Z(n12259) );
  XNOR U12211 ( .A(n12265), .B(n12591), .Z(n12258) );
  XNOR U12212 ( .A(n12266), .B(n12267), .Z(n12591) );
  AND U12213 ( .A(n12592), .B(n12593), .Z(n12267) );
  NANDN U12214 ( .A(n12594), .B(n12595), .Z(n12593) );
  NANDN U12215 ( .A(n12596), .B(n12597), .Z(n12592) );
  NANDN U12216 ( .A(n12595), .B(n12594), .Z(n12597) );
  ANDN U12217 ( .B(\stack[0][45] ), .A(n5364), .Z(n12266) );
  XNOR U12218 ( .A(n12272), .B(n12598), .Z(n12265) );
  XNOR U12219 ( .A(n12273), .B(n12274), .Z(n12598) );
  AND U12220 ( .A(n12599), .B(n12600), .Z(n12274) );
  NAND U12221 ( .A(n12601), .B(n12602), .Z(n12600) );
  NANDN U12222 ( .A(n12603), .B(n12604), .Z(n12599) );
  OR U12223 ( .A(n12601), .B(n12602), .Z(n12604) );
  ANDN U12224 ( .B(\stack[0][44] ), .A(n5387), .Z(n12273) );
  XNOR U12225 ( .A(n12279), .B(n12605), .Z(n12272) );
  XNOR U12226 ( .A(n12280), .B(n12281), .Z(n12605) );
  AND U12227 ( .A(n12606), .B(n12607), .Z(n12281) );
  NANDN U12228 ( .A(n12608), .B(n12609), .Z(n12607) );
  NANDN U12229 ( .A(n12610), .B(n12611), .Z(n12606) );
  NANDN U12230 ( .A(n12609), .B(n12608), .Z(n12611) );
  ANDN U12231 ( .B(\stack[1][10] ), .A(n6190), .Z(n12280) );
  XNOR U12232 ( .A(n12286), .B(n12612), .Z(n12279) );
  XNOR U12233 ( .A(n12287), .B(n12288), .Z(n12612) );
  AND U12234 ( .A(n12613), .B(n12614), .Z(n12288) );
  NAND U12235 ( .A(n12615), .B(n12616), .Z(n12614) );
  NANDN U12236 ( .A(n12617), .B(n12618), .Z(n12613) );
  OR U12237 ( .A(n12615), .B(n12616), .Z(n12618) );
  ANDN U12238 ( .B(\stack[1][11] ), .A(n6166), .Z(n12287) );
  XNOR U12239 ( .A(n12293), .B(n12619), .Z(n12286) );
  XNOR U12240 ( .A(n12294), .B(n12295), .Z(n12619) );
  AND U12241 ( .A(n12620), .B(n12621), .Z(n12295) );
  NANDN U12242 ( .A(n12622), .B(n12623), .Z(n12621) );
  NANDN U12243 ( .A(n12624), .B(n12625), .Z(n12620) );
  NANDN U12244 ( .A(n12623), .B(n12622), .Z(n12625) );
  ANDN U12245 ( .B(\stack[1][12] ), .A(n6142), .Z(n12294) );
  XNOR U12246 ( .A(n12300), .B(n12626), .Z(n12293) );
  XNOR U12247 ( .A(n12301), .B(n12302), .Z(n12626) );
  AND U12248 ( .A(n12627), .B(n12628), .Z(n12302) );
  NAND U12249 ( .A(n12629), .B(n12630), .Z(n12628) );
  NANDN U12250 ( .A(n12631), .B(n12632), .Z(n12627) );
  OR U12251 ( .A(n12629), .B(n12630), .Z(n12632) );
  ANDN U12252 ( .B(\stack[1][13] ), .A(n6118), .Z(n12301) );
  XNOR U12253 ( .A(n12307), .B(n12633), .Z(n12300) );
  XNOR U12254 ( .A(n12308), .B(n12309), .Z(n12633) );
  AND U12255 ( .A(n12634), .B(n12635), .Z(n12309) );
  NANDN U12256 ( .A(n12636), .B(n12637), .Z(n12635) );
  NANDN U12257 ( .A(n12638), .B(n12639), .Z(n12634) );
  NANDN U12258 ( .A(n12637), .B(n12636), .Z(n12639) );
  ANDN U12259 ( .B(\stack[1][14] ), .A(n6094), .Z(n12308) );
  XNOR U12260 ( .A(n12314), .B(n12640), .Z(n12307) );
  XNOR U12261 ( .A(n12315), .B(n12316), .Z(n12640) );
  AND U12262 ( .A(n12641), .B(n12642), .Z(n12316) );
  NAND U12263 ( .A(n12643), .B(n12644), .Z(n12642) );
  NANDN U12264 ( .A(n12645), .B(n12646), .Z(n12641) );
  OR U12265 ( .A(n12643), .B(n12644), .Z(n12646) );
  ANDN U12266 ( .B(\stack[1][15] ), .A(n6070), .Z(n12315) );
  XNOR U12267 ( .A(n12321), .B(n12647), .Z(n12314) );
  XNOR U12268 ( .A(n12322), .B(n12323), .Z(n12647) );
  AND U12269 ( .A(n12648), .B(n12649), .Z(n12323) );
  NANDN U12270 ( .A(n12650), .B(n12651), .Z(n12649) );
  NANDN U12271 ( .A(n12652), .B(n12653), .Z(n12648) );
  NANDN U12272 ( .A(n12651), .B(n12650), .Z(n12653) );
  ANDN U12273 ( .B(\stack[1][16] ), .A(n6046), .Z(n12322) );
  XNOR U12274 ( .A(n12328), .B(n12654), .Z(n12321) );
  XNOR U12275 ( .A(n12329), .B(n12330), .Z(n12654) );
  AND U12276 ( .A(n12655), .B(n12656), .Z(n12330) );
  NAND U12277 ( .A(n12657), .B(n12658), .Z(n12656) );
  NANDN U12278 ( .A(n12659), .B(n12660), .Z(n12655) );
  OR U12279 ( .A(n12657), .B(n12658), .Z(n12660) );
  ANDN U12280 ( .B(\stack[1][17] ), .A(n6022), .Z(n12329) );
  XNOR U12281 ( .A(n12335), .B(n12661), .Z(n12328) );
  XNOR U12282 ( .A(n12336), .B(n12337), .Z(n12661) );
  AND U12283 ( .A(n12662), .B(n12663), .Z(n12337) );
  NANDN U12284 ( .A(n12664), .B(n12665), .Z(n12663) );
  NANDN U12285 ( .A(n12666), .B(n12667), .Z(n12662) );
  NANDN U12286 ( .A(n12665), .B(n12664), .Z(n12667) );
  ANDN U12287 ( .B(\stack[1][18] ), .A(n5998), .Z(n12336) );
  XNOR U12288 ( .A(n12342), .B(n12668), .Z(n12335) );
  XNOR U12289 ( .A(n12343), .B(n12344), .Z(n12668) );
  AND U12290 ( .A(n12669), .B(n12670), .Z(n12344) );
  NAND U12291 ( .A(n12671), .B(n12672), .Z(n12670) );
  NANDN U12292 ( .A(n12673), .B(n12674), .Z(n12669) );
  OR U12293 ( .A(n12671), .B(n12672), .Z(n12674) );
  ANDN U12294 ( .B(\stack[1][19] ), .A(n5974), .Z(n12343) );
  XNOR U12295 ( .A(n12349), .B(n12675), .Z(n12342) );
  XNOR U12296 ( .A(n12350), .B(n12351), .Z(n12675) );
  AND U12297 ( .A(n12676), .B(n12677), .Z(n12351) );
  NANDN U12298 ( .A(n12678), .B(n12679), .Z(n12677) );
  NANDN U12299 ( .A(n12680), .B(n12681), .Z(n12676) );
  NANDN U12300 ( .A(n12679), .B(n12678), .Z(n12681) );
  ANDN U12301 ( .B(\stack[1][20] ), .A(n5950), .Z(n12350) );
  XNOR U12302 ( .A(n12356), .B(n12682), .Z(n12349) );
  XNOR U12303 ( .A(n12357), .B(n12358), .Z(n12682) );
  AND U12304 ( .A(n12683), .B(n12684), .Z(n12358) );
  NAND U12305 ( .A(n12685), .B(n12686), .Z(n12684) );
  NANDN U12306 ( .A(n12687), .B(n12688), .Z(n12683) );
  OR U12307 ( .A(n12685), .B(n12686), .Z(n12688) );
  ANDN U12308 ( .B(\stack[1][21] ), .A(n5926), .Z(n12357) );
  XNOR U12309 ( .A(n12363), .B(n12689), .Z(n12356) );
  XNOR U12310 ( .A(n12364), .B(n12365), .Z(n12689) );
  AND U12311 ( .A(n12690), .B(n12691), .Z(n12365) );
  NANDN U12312 ( .A(n12692), .B(n12693), .Z(n12691) );
  NANDN U12313 ( .A(n12694), .B(n12695), .Z(n12690) );
  NANDN U12314 ( .A(n12693), .B(n12692), .Z(n12695) );
  ANDN U12315 ( .B(\stack[1][22] ), .A(n5902), .Z(n12364) );
  XNOR U12316 ( .A(n12370), .B(n12696), .Z(n12363) );
  XNOR U12317 ( .A(n12371), .B(n12372), .Z(n12696) );
  AND U12318 ( .A(n12697), .B(n12698), .Z(n12372) );
  NAND U12319 ( .A(n12699), .B(n12700), .Z(n12698) );
  NANDN U12320 ( .A(n12701), .B(n12702), .Z(n12697) );
  OR U12321 ( .A(n12699), .B(n12700), .Z(n12702) );
  ANDN U12322 ( .B(\stack[1][23] ), .A(n5878), .Z(n12371) );
  XNOR U12323 ( .A(n12377), .B(n12703), .Z(n12370) );
  XNOR U12324 ( .A(n12378), .B(n12379), .Z(n12703) );
  AND U12325 ( .A(n12704), .B(n12705), .Z(n12379) );
  NANDN U12326 ( .A(n12706), .B(n12707), .Z(n12705) );
  NANDN U12327 ( .A(n12708), .B(n12709), .Z(n12704) );
  NANDN U12328 ( .A(n12707), .B(n12706), .Z(n12709) );
  ANDN U12329 ( .B(\stack[1][24] ), .A(n5854), .Z(n12378) );
  XNOR U12330 ( .A(n12384), .B(n12710), .Z(n12377) );
  XNOR U12331 ( .A(n12385), .B(n12386), .Z(n12710) );
  AND U12332 ( .A(n12711), .B(n12712), .Z(n12386) );
  NAND U12333 ( .A(n12713), .B(n12714), .Z(n12712) );
  NANDN U12334 ( .A(n12715), .B(n12716), .Z(n12711) );
  OR U12335 ( .A(n12713), .B(n12714), .Z(n12716) );
  ANDN U12336 ( .B(\stack[1][25] ), .A(n5830), .Z(n12385) );
  XNOR U12337 ( .A(n12391), .B(n12717), .Z(n12384) );
  XNOR U12338 ( .A(n12392), .B(n12393), .Z(n12717) );
  AND U12339 ( .A(n12718), .B(n12719), .Z(n12393) );
  NANDN U12340 ( .A(n12720), .B(n12721), .Z(n12719) );
  NANDN U12341 ( .A(n12722), .B(n12723), .Z(n12718) );
  NANDN U12342 ( .A(n12721), .B(n12720), .Z(n12723) );
  ANDN U12343 ( .B(\stack[1][26] ), .A(n5806), .Z(n12392) );
  XNOR U12344 ( .A(n12398), .B(n12724), .Z(n12391) );
  XNOR U12345 ( .A(n12399), .B(n12400), .Z(n12724) );
  AND U12346 ( .A(n12725), .B(n12726), .Z(n12400) );
  NAND U12347 ( .A(n12727), .B(n12728), .Z(n12726) );
  NANDN U12348 ( .A(n12729), .B(n12730), .Z(n12725) );
  OR U12349 ( .A(n12727), .B(n12728), .Z(n12730) );
  ANDN U12350 ( .B(\stack[1][27] ), .A(n5782), .Z(n12399) );
  XNOR U12351 ( .A(n12405), .B(n12731), .Z(n12398) );
  XNOR U12352 ( .A(n12406), .B(n12407), .Z(n12731) );
  AND U12353 ( .A(n12732), .B(n12733), .Z(n12407) );
  NANDN U12354 ( .A(n12734), .B(n12735), .Z(n12733) );
  NANDN U12355 ( .A(n12736), .B(n12737), .Z(n12732) );
  NANDN U12356 ( .A(n12735), .B(n12734), .Z(n12737) );
  ANDN U12357 ( .B(\stack[1][28] ), .A(n5758), .Z(n12406) );
  XNOR U12358 ( .A(n12412), .B(n12738), .Z(n12405) );
  XNOR U12359 ( .A(n12413), .B(n12414), .Z(n12738) );
  AND U12360 ( .A(n12739), .B(n12740), .Z(n12414) );
  NAND U12361 ( .A(n12741), .B(n12742), .Z(n12740) );
  NANDN U12362 ( .A(n12743), .B(n12744), .Z(n12739) );
  OR U12363 ( .A(n12741), .B(n12742), .Z(n12744) );
  ANDN U12364 ( .B(\stack[1][29] ), .A(n5734), .Z(n12413) );
  XNOR U12365 ( .A(n12419), .B(n12745), .Z(n12412) );
  XNOR U12366 ( .A(n12420), .B(n12421), .Z(n12745) );
  AND U12367 ( .A(n12746), .B(n12747), .Z(n12421) );
  NANDN U12368 ( .A(n12748), .B(n12749), .Z(n12747) );
  NANDN U12369 ( .A(n12750), .B(n12751), .Z(n12746) );
  NANDN U12370 ( .A(n12749), .B(n12748), .Z(n12751) );
  ANDN U12371 ( .B(\stack[1][30] ), .A(n5710), .Z(n12420) );
  XNOR U12372 ( .A(n12426), .B(n12752), .Z(n12419) );
  XNOR U12373 ( .A(n12427), .B(n12428), .Z(n12752) );
  AND U12374 ( .A(n12753), .B(n12754), .Z(n12428) );
  NAND U12375 ( .A(n12755), .B(n12756), .Z(n12754) );
  NANDN U12376 ( .A(n12757), .B(n12758), .Z(n12753) );
  OR U12377 ( .A(n12755), .B(n12756), .Z(n12758) );
  ANDN U12378 ( .B(\stack[1][31] ), .A(n5686), .Z(n12427) );
  XNOR U12379 ( .A(n12433), .B(n12759), .Z(n12426) );
  XNOR U12380 ( .A(n12434), .B(n12435), .Z(n12759) );
  AND U12381 ( .A(n12760), .B(n12761), .Z(n12435) );
  NANDN U12382 ( .A(n12762), .B(n12763), .Z(n12761) );
  NANDN U12383 ( .A(n12764), .B(n12765), .Z(n12760) );
  NANDN U12384 ( .A(n12763), .B(n12762), .Z(n12765) );
  ANDN U12385 ( .B(\stack[1][32] ), .A(n5662), .Z(n12434) );
  XNOR U12386 ( .A(n12440), .B(n12766), .Z(n12433) );
  XNOR U12387 ( .A(n12441), .B(n12442), .Z(n12766) );
  AND U12388 ( .A(n12767), .B(n12768), .Z(n12442) );
  NAND U12389 ( .A(n12769), .B(n12770), .Z(n12768) );
  NANDN U12390 ( .A(n12771), .B(n12772), .Z(n12767) );
  OR U12391 ( .A(n12769), .B(n12770), .Z(n12772) );
  ANDN U12392 ( .B(\stack[1][33] ), .A(n5638), .Z(n12441) );
  XNOR U12393 ( .A(n12447), .B(n12773), .Z(n12440) );
  XNOR U12394 ( .A(n12448), .B(n12449), .Z(n12773) );
  AND U12395 ( .A(n12774), .B(n12775), .Z(n12449) );
  NANDN U12396 ( .A(n12776), .B(n12777), .Z(n12775) );
  NANDN U12397 ( .A(n12778), .B(n12779), .Z(n12774) );
  NANDN U12398 ( .A(n12777), .B(n12776), .Z(n12779) );
  ANDN U12399 ( .B(\stack[1][34] ), .A(n5614), .Z(n12448) );
  XNOR U12400 ( .A(n12454), .B(n12780), .Z(n12447) );
  XNOR U12401 ( .A(n12455), .B(n12456), .Z(n12780) );
  AND U12402 ( .A(n12781), .B(n12782), .Z(n12456) );
  NAND U12403 ( .A(n12783), .B(n12784), .Z(n12782) );
  NANDN U12404 ( .A(n12785), .B(n12786), .Z(n12781) );
  OR U12405 ( .A(n12783), .B(n12784), .Z(n12786) );
  ANDN U12406 ( .B(\stack[1][35] ), .A(n5590), .Z(n12455) );
  XNOR U12407 ( .A(n12461), .B(n12787), .Z(n12454) );
  XNOR U12408 ( .A(n12462), .B(n12463), .Z(n12787) );
  AND U12409 ( .A(n12788), .B(n12789), .Z(n12463) );
  NANDN U12410 ( .A(n12790), .B(n12791), .Z(n12789) );
  NANDN U12411 ( .A(n12792), .B(n12793), .Z(n12788) );
  NANDN U12412 ( .A(n12791), .B(n12790), .Z(n12793) );
  ANDN U12413 ( .B(\stack[1][36] ), .A(n5566), .Z(n12462) );
  XNOR U12414 ( .A(n12468), .B(n12794), .Z(n12461) );
  XOR U12415 ( .A(n12470), .B(n12471), .Z(n12794) );
  NAND U12416 ( .A(n12795), .B(n12796), .Z(n12471) );
  NAND U12417 ( .A(n12797), .B(n12798), .Z(n12796) );
  OR U12418 ( .A(n12799), .B(n12800), .Z(n12797) );
  AND U12419 ( .A(\stack[0][16] ), .B(\stack[1][37] ), .Z(n12470) );
  XNOR U12420 ( .A(n12477), .B(n12801), .Z(n12468) );
  XOR U12421 ( .A(n12478), .B(n12476), .Z(n12801) );
  AND U12422 ( .A(\stack[0][15] ), .B(\stack[1][38] ), .Z(n12476) );
  NAND U12423 ( .A(n12802), .B(n12803), .Z(n12478) );
  OR U12424 ( .A(n12804), .B(n12805), .Z(n12803) );
  NAND U12425 ( .A(n12806), .B(n12807), .Z(n12802) );
  NAND U12426 ( .A(n12805), .B(n12804), .Z(n12806) );
  XNOR U12427 ( .A(n12482), .B(n12808), .Z(n12477) );
  XNOR U12428 ( .A(n12483), .B(n12484), .Z(n12808) );
  AND U12429 ( .A(n12809), .B(n12810), .Z(n12484) );
  NAND U12430 ( .A(n12811), .B(n12812), .Z(n12810) );
  NANDN U12431 ( .A(n12813), .B(n12814), .Z(n12809) );
  OR U12432 ( .A(n12811), .B(n12812), .Z(n12814) );
  ANDN U12433 ( .B(\stack[1][39] ), .A(n5494), .Z(n12483) );
  XNOR U12434 ( .A(n12489), .B(n12815), .Z(n12482) );
  XNOR U12435 ( .A(n12490), .B(n12491), .Z(n12815) );
  AND U12436 ( .A(n12816), .B(n12817), .Z(n12491) );
  NANDN U12437 ( .A(n12818), .B(n12819), .Z(n12817) );
  NANDN U12438 ( .A(n12820), .B(n12821), .Z(n12816) );
  NANDN U12439 ( .A(n12819), .B(n12818), .Z(n12821) );
  ANDN U12440 ( .B(\stack[1][40] ), .A(n5470), .Z(n12490) );
  XNOR U12441 ( .A(n12496), .B(n12822), .Z(n12489) );
  XNOR U12442 ( .A(n12497), .B(n12498), .Z(n12822) );
  AND U12443 ( .A(n12823), .B(n12824), .Z(n12498) );
  NAND U12444 ( .A(n12825), .B(n12826), .Z(n12824) );
  NANDN U12445 ( .A(n12827), .B(n12828), .Z(n12823) );
  OR U12446 ( .A(n12825), .B(n12826), .Z(n12828) );
  ANDN U12447 ( .B(\stack[1][41] ), .A(n5446), .Z(n12497) );
  XNOR U12448 ( .A(n12503), .B(n12829), .Z(n12496) );
  XNOR U12449 ( .A(n12504), .B(n12505), .Z(n12829) );
  AND U12450 ( .A(n12830), .B(n12831), .Z(n12505) );
  NANDN U12451 ( .A(n12832), .B(n12833), .Z(n12831) );
  NANDN U12452 ( .A(n12834), .B(n12835), .Z(n12830) );
  NANDN U12453 ( .A(n12833), .B(n12832), .Z(n12835) );
  ANDN U12454 ( .B(\stack[1][42] ), .A(n5422), .Z(n12504) );
  XNOR U12455 ( .A(n12510), .B(n12836), .Z(n12503) );
  XNOR U12456 ( .A(n12511), .B(n12512), .Z(n12836) );
  AND U12457 ( .A(n12837), .B(n12838), .Z(n12512) );
  NAND U12458 ( .A(n12839), .B(n12840), .Z(n12838) );
  NANDN U12459 ( .A(n12841), .B(n12842), .Z(n12837) );
  OR U12460 ( .A(n12839), .B(n12840), .Z(n12842) );
  ANDN U12461 ( .B(\stack[1][43] ), .A(n5398), .Z(n12511) );
  XNOR U12462 ( .A(n12517), .B(n12843), .Z(n12510) );
  XNOR U12463 ( .A(n12518), .B(n12519), .Z(n12843) );
  AND U12464 ( .A(n12844), .B(n12845), .Z(n12519) );
  NANDN U12465 ( .A(n12846), .B(n12847), .Z(n12845) );
  NANDN U12466 ( .A(n12848), .B(n12849), .Z(n12844) );
  NANDN U12467 ( .A(n12847), .B(n12846), .Z(n12849) );
  ANDN U12468 ( .B(\stack[1][44] ), .A(n5374), .Z(n12518) );
  XNOR U12469 ( .A(n12524), .B(n12850), .Z(n12517) );
  XNOR U12470 ( .A(n12525), .B(n12526), .Z(n12850) );
  AND U12471 ( .A(n12851), .B(n12852), .Z(n12526) );
  NAND U12472 ( .A(n12853), .B(n12854), .Z(n12852) );
  NANDN U12473 ( .A(n12855), .B(n12856), .Z(n12851) );
  OR U12474 ( .A(n12853), .B(n12854), .Z(n12856) );
  ANDN U12475 ( .B(\stack[1][45] ), .A(n5350), .Z(n12525) );
  XNOR U12476 ( .A(n12531), .B(n12857), .Z(n12524) );
  XNOR U12477 ( .A(n12532), .B(n12533), .Z(n12857) );
  AND U12478 ( .A(n12858), .B(n12859), .Z(n12533) );
  NANDN U12479 ( .A(n12860), .B(n12861), .Z(n12859) );
  NANDN U12480 ( .A(n12862), .B(n12863), .Z(n12858) );
  NANDN U12481 ( .A(n12861), .B(n12860), .Z(n12863) );
  ANDN U12482 ( .B(\stack[1][46] ), .A(n5326), .Z(n12532) );
  XNOR U12483 ( .A(n12538), .B(n12864), .Z(n12531) );
  XNOR U12484 ( .A(n12539), .B(n12540), .Z(n12864) );
  AND U12485 ( .A(n12865), .B(n12866), .Z(n12540) );
  NAND U12486 ( .A(n12867), .B(n12868), .Z(n12866) );
  NANDN U12487 ( .A(n12869), .B(n12870), .Z(n12865) );
  OR U12488 ( .A(n12867), .B(n12868), .Z(n12870) );
  ANDN U12489 ( .B(\stack[1][47] ), .A(n5302), .Z(n12539) );
  XNOR U12490 ( .A(n12545), .B(n12871), .Z(n12538) );
  XNOR U12491 ( .A(n12546), .B(n12547), .Z(n12871) );
  AND U12492 ( .A(n12872), .B(n12873), .Z(n12547) );
  NANDN U12493 ( .A(n12874), .B(n12875), .Z(n12873) );
  NANDN U12494 ( .A(n12876), .B(n12877), .Z(n12872) );
  NANDN U12495 ( .A(n12875), .B(n12874), .Z(n12877) );
  ANDN U12496 ( .B(\stack[1][48] ), .A(n5278), .Z(n12546) );
  XNOR U12497 ( .A(n12552), .B(n12878), .Z(n12545) );
  XNOR U12498 ( .A(n12553), .B(n12554), .Z(n12878) );
  AND U12499 ( .A(n12879), .B(n12880), .Z(n12554) );
  NAND U12500 ( .A(n12881), .B(n12882), .Z(n12880) );
  NANDN U12501 ( .A(n12883), .B(n12884), .Z(n12879) );
  OR U12502 ( .A(n12881), .B(n12882), .Z(n12884) );
  ANDN U12503 ( .B(\stack[1][49] ), .A(n5254), .Z(n12553) );
  XNOR U12504 ( .A(n12559), .B(n12885), .Z(n12552) );
  XNOR U12505 ( .A(n12560), .B(n12561), .Z(n12885) );
  AND U12506 ( .A(n12886), .B(n12887), .Z(n12561) );
  NAND U12507 ( .A(n12888), .B(n12889), .Z(n12887) );
  NAND U12508 ( .A(n12890), .B(n12891), .Z(n12886) );
  OR U12509 ( .A(n12888), .B(n12889), .Z(n12890) );
  ANDN U12510 ( .B(\stack[1][50] ), .A(n5230), .Z(n12560) );
  XNOR U12511 ( .A(n12566), .B(n12892), .Z(n12559) );
  XNOR U12512 ( .A(n12567), .B(n12569), .Z(n12892) );
  ANDN U12513 ( .B(n12893), .A(n12894), .Z(n12569) );
  ANDN U12514 ( .B(\stack[0][0] ), .A(n6420), .Z(n12893) );
  ANDN U12515 ( .B(\stack[1][51] ), .A(n5206), .Z(n12567) );
  XOR U12516 ( .A(n12572), .B(n12895), .Z(n12566) );
  NANDN U12517 ( .A(n5160), .B(\stack[1][53] ), .Z(n12895) );
  NANDN U12518 ( .A(n6420), .B(\stack[0][1] ), .Z(n12572) );
  ANDN U12519 ( .B(\stack[1][5] ), .A(n6310), .Z(n9027) );
  AND U12520 ( .A(n12896), .B(n12897), .Z(n9028) );
  NANDN U12521 ( .A(n9032), .B(n9034), .Z(n12897) );
  NANDN U12522 ( .A(n9035), .B(n12898), .Z(n12896) );
  NANDN U12523 ( .A(n9034), .B(n9032), .Z(n12898) );
  XOR U12524 ( .A(n12580), .B(n12899), .Z(n9032) );
  XNOR U12525 ( .A(n12581), .B(n12582), .Z(n12899) );
  AND U12526 ( .A(n12900), .B(n12901), .Z(n12582) );
  NAND U12527 ( .A(n12902), .B(n12903), .Z(n12901) );
  NANDN U12528 ( .A(n12904), .B(n12905), .Z(n12900) );
  OR U12529 ( .A(n12902), .B(n12903), .Z(n12905) );
  ANDN U12530 ( .B(\stack[0][46] ), .A(n5316), .Z(n12581) );
  XNOR U12531 ( .A(n12587), .B(n12906), .Z(n12580) );
  XNOR U12532 ( .A(n12588), .B(n12589), .Z(n12906) );
  AND U12533 ( .A(n12907), .B(n12908), .Z(n12589) );
  NANDN U12534 ( .A(n12909), .B(n12910), .Z(n12908) );
  NANDN U12535 ( .A(n12911), .B(n12912), .Z(n12907) );
  NANDN U12536 ( .A(n12910), .B(n12909), .Z(n12912) );
  ANDN U12537 ( .B(\stack[0][45] ), .A(n5340), .Z(n12588) );
  XNOR U12538 ( .A(n12594), .B(n12913), .Z(n12587) );
  XNOR U12539 ( .A(n12595), .B(n12596), .Z(n12913) );
  AND U12540 ( .A(n12914), .B(n12915), .Z(n12596) );
  NAND U12541 ( .A(n12916), .B(n12917), .Z(n12915) );
  NANDN U12542 ( .A(n12918), .B(n12919), .Z(n12914) );
  OR U12543 ( .A(n12916), .B(n12917), .Z(n12919) );
  ANDN U12544 ( .B(\stack[0][44] ), .A(n5364), .Z(n12595) );
  XNOR U12545 ( .A(n12601), .B(n12920), .Z(n12594) );
  XNOR U12546 ( .A(n12602), .B(n12603), .Z(n12920) );
  AND U12547 ( .A(n12921), .B(n12922), .Z(n12603) );
  NANDN U12548 ( .A(n12923), .B(n12924), .Z(n12922) );
  NANDN U12549 ( .A(n12925), .B(n12926), .Z(n12921) );
  NANDN U12550 ( .A(n12924), .B(n12923), .Z(n12926) );
  ANDN U12551 ( .B(\stack[0][43] ), .A(n5387), .Z(n12602) );
  XNOR U12552 ( .A(n12608), .B(n12927), .Z(n12601) );
  XNOR U12553 ( .A(n12609), .B(n12610), .Z(n12927) );
  AND U12554 ( .A(n12928), .B(n12929), .Z(n12610) );
  NAND U12555 ( .A(n12930), .B(n12931), .Z(n12929) );
  NANDN U12556 ( .A(n12932), .B(n12933), .Z(n12928) );
  OR U12557 ( .A(n12930), .B(n12931), .Z(n12933) );
  ANDN U12558 ( .B(\stack[1][10] ), .A(n6166), .Z(n12609) );
  XNOR U12559 ( .A(n12615), .B(n12934), .Z(n12608) );
  XNOR U12560 ( .A(n12616), .B(n12617), .Z(n12934) );
  AND U12561 ( .A(n12935), .B(n12936), .Z(n12617) );
  NANDN U12562 ( .A(n12937), .B(n12938), .Z(n12936) );
  NANDN U12563 ( .A(n12939), .B(n12940), .Z(n12935) );
  NANDN U12564 ( .A(n12938), .B(n12937), .Z(n12940) );
  ANDN U12565 ( .B(\stack[1][11] ), .A(n6142), .Z(n12616) );
  XNOR U12566 ( .A(n12622), .B(n12941), .Z(n12615) );
  XNOR U12567 ( .A(n12623), .B(n12624), .Z(n12941) );
  AND U12568 ( .A(n12942), .B(n12943), .Z(n12624) );
  NAND U12569 ( .A(n12944), .B(n12945), .Z(n12943) );
  NANDN U12570 ( .A(n12946), .B(n12947), .Z(n12942) );
  OR U12571 ( .A(n12944), .B(n12945), .Z(n12947) );
  ANDN U12572 ( .B(\stack[1][12] ), .A(n6118), .Z(n12623) );
  XNOR U12573 ( .A(n12629), .B(n12948), .Z(n12622) );
  XNOR U12574 ( .A(n12630), .B(n12631), .Z(n12948) );
  AND U12575 ( .A(n12949), .B(n12950), .Z(n12631) );
  NANDN U12576 ( .A(n12951), .B(n12952), .Z(n12950) );
  NANDN U12577 ( .A(n12953), .B(n12954), .Z(n12949) );
  NANDN U12578 ( .A(n12952), .B(n12951), .Z(n12954) );
  ANDN U12579 ( .B(\stack[1][13] ), .A(n6094), .Z(n12630) );
  XNOR U12580 ( .A(n12636), .B(n12955), .Z(n12629) );
  XNOR U12581 ( .A(n12637), .B(n12638), .Z(n12955) );
  AND U12582 ( .A(n12956), .B(n12957), .Z(n12638) );
  NAND U12583 ( .A(n12958), .B(n12959), .Z(n12957) );
  NANDN U12584 ( .A(n12960), .B(n12961), .Z(n12956) );
  OR U12585 ( .A(n12958), .B(n12959), .Z(n12961) );
  ANDN U12586 ( .B(\stack[1][14] ), .A(n6070), .Z(n12637) );
  XNOR U12587 ( .A(n12643), .B(n12962), .Z(n12636) );
  XNOR U12588 ( .A(n12644), .B(n12645), .Z(n12962) );
  AND U12589 ( .A(n12963), .B(n12964), .Z(n12645) );
  NANDN U12590 ( .A(n12965), .B(n12966), .Z(n12964) );
  NANDN U12591 ( .A(n12967), .B(n12968), .Z(n12963) );
  NANDN U12592 ( .A(n12966), .B(n12965), .Z(n12968) );
  ANDN U12593 ( .B(\stack[1][15] ), .A(n6046), .Z(n12644) );
  XNOR U12594 ( .A(n12650), .B(n12969), .Z(n12643) );
  XNOR U12595 ( .A(n12651), .B(n12652), .Z(n12969) );
  AND U12596 ( .A(n12970), .B(n12971), .Z(n12652) );
  NAND U12597 ( .A(n12972), .B(n12973), .Z(n12971) );
  NANDN U12598 ( .A(n12974), .B(n12975), .Z(n12970) );
  OR U12599 ( .A(n12972), .B(n12973), .Z(n12975) );
  ANDN U12600 ( .B(\stack[1][16] ), .A(n6022), .Z(n12651) );
  XNOR U12601 ( .A(n12657), .B(n12976), .Z(n12650) );
  XNOR U12602 ( .A(n12658), .B(n12659), .Z(n12976) );
  AND U12603 ( .A(n12977), .B(n12978), .Z(n12659) );
  NANDN U12604 ( .A(n12979), .B(n12980), .Z(n12978) );
  NANDN U12605 ( .A(n12981), .B(n12982), .Z(n12977) );
  NANDN U12606 ( .A(n12980), .B(n12979), .Z(n12982) );
  ANDN U12607 ( .B(\stack[1][17] ), .A(n5998), .Z(n12658) );
  XNOR U12608 ( .A(n12664), .B(n12983), .Z(n12657) );
  XNOR U12609 ( .A(n12665), .B(n12666), .Z(n12983) );
  AND U12610 ( .A(n12984), .B(n12985), .Z(n12666) );
  NAND U12611 ( .A(n12986), .B(n12987), .Z(n12985) );
  NANDN U12612 ( .A(n12988), .B(n12989), .Z(n12984) );
  OR U12613 ( .A(n12986), .B(n12987), .Z(n12989) );
  ANDN U12614 ( .B(\stack[1][18] ), .A(n5974), .Z(n12665) );
  XNOR U12615 ( .A(n12671), .B(n12990), .Z(n12664) );
  XNOR U12616 ( .A(n12672), .B(n12673), .Z(n12990) );
  AND U12617 ( .A(n12991), .B(n12992), .Z(n12673) );
  NANDN U12618 ( .A(n12993), .B(n12994), .Z(n12992) );
  NANDN U12619 ( .A(n12995), .B(n12996), .Z(n12991) );
  NANDN U12620 ( .A(n12994), .B(n12993), .Z(n12996) );
  ANDN U12621 ( .B(\stack[1][19] ), .A(n5950), .Z(n12672) );
  XNOR U12622 ( .A(n12678), .B(n12997), .Z(n12671) );
  XNOR U12623 ( .A(n12679), .B(n12680), .Z(n12997) );
  AND U12624 ( .A(n12998), .B(n12999), .Z(n12680) );
  NAND U12625 ( .A(n13000), .B(n13001), .Z(n12999) );
  NANDN U12626 ( .A(n13002), .B(n13003), .Z(n12998) );
  OR U12627 ( .A(n13000), .B(n13001), .Z(n13003) );
  ANDN U12628 ( .B(\stack[1][20] ), .A(n5926), .Z(n12679) );
  XNOR U12629 ( .A(n12685), .B(n13004), .Z(n12678) );
  XNOR U12630 ( .A(n12686), .B(n12687), .Z(n13004) );
  AND U12631 ( .A(n13005), .B(n13006), .Z(n12687) );
  NANDN U12632 ( .A(n13007), .B(n13008), .Z(n13006) );
  NANDN U12633 ( .A(n13009), .B(n13010), .Z(n13005) );
  NANDN U12634 ( .A(n13008), .B(n13007), .Z(n13010) );
  ANDN U12635 ( .B(\stack[1][21] ), .A(n5902), .Z(n12686) );
  XNOR U12636 ( .A(n12692), .B(n13011), .Z(n12685) );
  XNOR U12637 ( .A(n12693), .B(n12694), .Z(n13011) );
  AND U12638 ( .A(n13012), .B(n13013), .Z(n12694) );
  NAND U12639 ( .A(n13014), .B(n13015), .Z(n13013) );
  NANDN U12640 ( .A(n13016), .B(n13017), .Z(n13012) );
  OR U12641 ( .A(n13014), .B(n13015), .Z(n13017) );
  ANDN U12642 ( .B(\stack[1][22] ), .A(n5878), .Z(n12693) );
  XNOR U12643 ( .A(n12699), .B(n13018), .Z(n12692) );
  XNOR U12644 ( .A(n12700), .B(n12701), .Z(n13018) );
  AND U12645 ( .A(n13019), .B(n13020), .Z(n12701) );
  NANDN U12646 ( .A(n13021), .B(n13022), .Z(n13020) );
  NANDN U12647 ( .A(n13023), .B(n13024), .Z(n13019) );
  NANDN U12648 ( .A(n13022), .B(n13021), .Z(n13024) );
  ANDN U12649 ( .B(\stack[1][23] ), .A(n5854), .Z(n12700) );
  XNOR U12650 ( .A(n12706), .B(n13025), .Z(n12699) );
  XNOR U12651 ( .A(n12707), .B(n12708), .Z(n13025) );
  AND U12652 ( .A(n13026), .B(n13027), .Z(n12708) );
  NAND U12653 ( .A(n13028), .B(n13029), .Z(n13027) );
  NANDN U12654 ( .A(n13030), .B(n13031), .Z(n13026) );
  OR U12655 ( .A(n13028), .B(n13029), .Z(n13031) );
  ANDN U12656 ( .B(\stack[1][24] ), .A(n5830), .Z(n12707) );
  XNOR U12657 ( .A(n12713), .B(n13032), .Z(n12706) );
  XNOR U12658 ( .A(n12714), .B(n12715), .Z(n13032) );
  AND U12659 ( .A(n13033), .B(n13034), .Z(n12715) );
  NANDN U12660 ( .A(n13035), .B(n13036), .Z(n13034) );
  NANDN U12661 ( .A(n13037), .B(n13038), .Z(n13033) );
  NANDN U12662 ( .A(n13036), .B(n13035), .Z(n13038) );
  ANDN U12663 ( .B(\stack[1][25] ), .A(n5806), .Z(n12714) );
  XNOR U12664 ( .A(n12720), .B(n13039), .Z(n12713) );
  XNOR U12665 ( .A(n12721), .B(n12722), .Z(n13039) );
  AND U12666 ( .A(n13040), .B(n13041), .Z(n12722) );
  NAND U12667 ( .A(n13042), .B(n13043), .Z(n13041) );
  NANDN U12668 ( .A(n13044), .B(n13045), .Z(n13040) );
  OR U12669 ( .A(n13042), .B(n13043), .Z(n13045) );
  ANDN U12670 ( .B(\stack[1][26] ), .A(n5782), .Z(n12721) );
  XNOR U12671 ( .A(n12727), .B(n13046), .Z(n12720) );
  XNOR U12672 ( .A(n12728), .B(n12729), .Z(n13046) );
  AND U12673 ( .A(n13047), .B(n13048), .Z(n12729) );
  NANDN U12674 ( .A(n13049), .B(n13050), .Z(n13048) );
  NANDN U12675 ( .A(n13051), .B(n13052), .Z(n13047) );
  NANDN U12676 ( .A(n13050), .B(n13049), .Z(n13052) );
  ANDN U12677 ( .B(\stack[1][27] ), .A(n5758), .Z(n12728) );
  XNOR U12678 ( .A(n12734), .B(n13053), .Z(n12727) );
  XNOR U12679 ( .A(n12735), .B(n12736), .Z(n13053) );
  AND U12680 ( .A(n13054), .B(n13055), .Z(n12736) );
  NAND U12681 ( .A(n13056), .B(n13057), .Z(n13055) );
  NANDN U12682 ( .A(n13058), .B(n13059), .Z(n13054) );
  OR U12683 ( .A(n13056), .B(n13057), .Z(n13059) );
  ANDN U12684 ( .B(\stack[1][28] ), .A(n5734), .Z(n12735) );
  XNOR U12685 ( .A(n12741), .B(n13060), .Z(n12734) );
  XNOR U12686 ( .A(n12742), .B(n12743), .Z(n13060) );
  AND U12687 ( .A(n13061), .B(n13062), .Z(n12743) );
  NANDN U12688 ( .A(n13063), .B(n13064), .Z(n13062) );
  NANDN U12689 ( .A(n13065), .B(n13066), .Z(n13061) );
  NANDN U12690 ( .A(n13064), .B(n13063), .Z(n13066) );
  ANDN U12691 ( .B(\stack[1][29] ), .A(n5710), .Z(n12742) );
  XNOR U12692 ( .A(n12748), .B(n13067), .Z(n12741) );
  XNOR U12693 ( .A(n12749), .B(n12750), .Z(n13067) );
  AND U12694 ( .A(n13068), .B(n13069), .Z(n12750) );
  NAND U12695 ( .A(n13070), .B(n13071), .Z(n13069) );
  NANDN U12696 ( .A(n13072), .B(n13073), .Z(n13068) );
  OR U12697 ( .A(n13070), .B(n13071), .Z(n13073) );
  ANDN U12698 ( .B(\stack[1][30] ), .A(n5686), .Z(n12749) );
  XNOR U12699 ( .A(n12755), .B(n13074), .Z(n12748) );
  XNOR U12700 ( .A(n12756), .B(n12757), .Z(n13074) );
  AND U12701 ( .A(n13075), .B(n13076), .Z(n12757) );
  NANDN U12702 ( .A(n13077), .B(n13078), .Z(n13076) );
  NANDN U12703 ( .A(n13079), .B(n13080), .Z(n13075) );
  NANDN U12704 ( .A(n13078), .B(n13077), .Z(n13080) );
  ANDN U12705 ( .B(\stack[1][31] ), .A(n5662), .Z(n12756) );
  XNOR U12706 ( .A(n12762), .B(n13081), .Z(n12755) );
  XNOR U12707 ( .A(n12763), .B(n12764), .Z(n13081) );
  AND U12708 ( .A(n13082), .B(n13083), .Z(n12764) );
  NAND U12709 ( .A(n13084), .B(n13085), .Z(n13083) );
  NANDN U12710 ( .A(n13086), .B(n13087), .Z(n13082) );
  OR U12711 ( .A(n13084), .B(n13085), .Z(n13087) );
  ANDN U12712 ( .B(\stack[1][32] ), .A(n5638), .Z(n12763) );
  XNOR U12713 ( .A(n12769), .B(n13088), .Z(n12762) );
  XNOR U12714 ( .A(n12770), .B(n12771), .Z(n13088) );
  AND U12715 ( .A(n13089), .B(n13090), .Z(n12771) );
  NANDN U12716 ( .A(n13091), .B(n13092), .Z(n13090) );
  NANDN U12717 ( .A(n13093), .B(n13094), .Z(n13089) );
  NANDN U12718 ( .A(n13092), .B(n13091), .Z(n13094) );
  ANDN U12719 ( .B(\stack[1][33] ), .A(n5614), .Z(n12770) );
  XNOR U12720 ( .A(n12776), .B(n13095), .Z(n12769) );
  XNOR U12721 ( .A(n12777), .B(n12778), .Z(n13095) );
  AND U12722 ( .A(n13096), .B(n13097), .Z(n12778) );
  NAND U12723 ( .A(n13098), .B(n13099), .Z(n13097) );
  NANDN U12724 ( .A(n13100), .B(n13101), .Z(n13096) );
  OR U12725 ( .A(n13098), .B(n13099), .Z(n13101) );
  ANDN U12726 ( .B(\stack[1][34] ), .A(n5590), .Z(n12777) );
  XNOR U12727 ( .A(n12783), .B(n13102), .Z(n12776) );
  XNOR U12728 ( .A(n12784), .B(n12785), .Z(n13102) );
  AND U12729 ( .A(n13103), .B(n13104), .Z(n12785) );
  NANDN U12730 ( .A(n13105), .B(n13106), .Z(n13104) );
  NANDN U12731 ( .A(n13107), .B(n13108), .Z(n13103) );
  NANDN U12732 ( .A(n13106), .B(n13105), .Z(n13108) );
  ANDN U12733 ( .B(\stack[1][35] ), .A(n5566), .Z(n12784) );
  XNOR U12734 ( .A(n12790), .B(n13109), .Z(n12783) );
  XNOR U12735 ( .A(n12791), .B(n12792), .Z(n13109) );
  AND U12736 ( .A(n13110), .B(n13111), .Z(n12792) );
  NAND U12737 ( .A(n13112), .B(n13113), .Z(n13111) );
  NANDN U12738 ( .A(n13114), .B(n13115), .Z(n13110) );
  OR U12739 ( .A(n13112), .B(n13113), .Z(n13115) );
  ANDN U12740 ( .B(\stack[1][36] ), .A(n5542), .Z(n12791) );
  XNOR U12741 ( .A(n12798), .B(n13116), .Z(n12790) );
  XOR U12742 ( .A(n12799), .B(n12800), .Z(n13116) );
  NAND U12743 ( .A(n13117), .B(n13118), .Z(n12800) );
  NANDN U12744 ( .A(n13119), .B(n13120), .Z(n13118) );
  OR U12745 ( .A(n13121), .B(n13122), .Z(n13120) );
  AND U12746 ( .A(\stack[0][15] ), .B(\stack[1][37] ), .Z(n12799) );
  XNOR U12747 ( .A(n12805), .B(n13123), .Z(n12798) );
  XNOR U12748 ( .A(n12804), .B(n12807), .Z(n13123) );
  AND U12749 ( .A(\stack[0][14] ), .B(\stack[1][38] ), .Z(n12807) );
  AND U12750 ( .A(n13124), .B(n13125), .Z(n12804) );
  NAND U12751 ( .A(n13126), .B(n13127), .Z(n13125) );
  OR U12752 ( .A(n13128), .B(n13129), .Z(n13126) );
  XNOR U12753 ( .A(n12811), .B(n13130), .Z(n12805) );
  XNOR U12754 ( .A(n12812), .B(n12813), .Z(n13130) );
  AND U12755 ( .A(n13131), .B(n13132), .Z(n12813) );
  NANDN U12756 ( .A(n13133), .B(n13134), .Z(n13132) );
  NANDN U12757 ( .A(n13135), .B(n13136), .Z(n13131) );
  NANDN U12758 ( .A(n13134), .B(n13133), .Z(n13136) );
  ANDN U12759 ( .B(\stack[1][39] ), .A(n5470), .Z(n12812) );
  XNOR U12760 ( .A(n12818), .B(n13137), .Z(n12811) );
  XNOR U12761 ( .A(n12819), .B(n12820), .Z(n13137) );
  AND U12762 ( .A(n13138), .B(n13139), .Z(n12820) );
  NAND U12763 ( .A(n13140), .B(n13141), .Z(n13139) );
  NANDN U12764 ( .A(n13142), .B(n13143), .Z(n13138) );
  OR U12765 ( .A(n13140), .B(n13141), .Z(n13143) );
  ANDN U12766 ( .B(\stack[1][40] ), .A(n5446), .Z(n12819) );
  XNOR U12767 ( .A(n12825), .B(n13144), .Z(n12818) );
  XNOR U12768 ( .A(n12826), .B(n12827), .Z(n13144) );
  AND U12769 ( .A(n13145), .B(n13146), .Z(n12827) );
  NANDN U12770 ( .A(n13147), .B(n13148), .Z(n13146) );
  NANDN U12771 ( .A(n13149), .B(n13150), .Z(n13145) );
  NANDN U12772 ( .A(n13148), .B(n13147), .Z(n13150) );
  ANDN U12773 ( .B(\stack[1][41] ), .A(n5422), .Z(n12826) );
  XNOR U12774 ( .A(n12832), .B(n13151), .Z(n12825) );
  XNOR U12775 ( .A(n12833), .B(n12834), .Z(n13151) );
  AND U12776 ( .A(n13152), .B(n13153), .Z(n12834) );
  NAND U12777 ( .A(n13154), .B(n13155), .Z(n13153) );
  NANDN U12778 ( .A(n13156), .B(n13157), .Z(n13152) );
  OR U12779 ( .A(n13154), .B(n13155), .Z(n13157) );
  ANDN U12780 ( .B(\stack[1][42] ), .A(n5398), .Z(n12833) );
  XNOR U12781 ( .A(n12839), .B(n13158), .Z(n12832) );
  XNOR U12782 ( .A(n12840), .B(n12841), .Z(n13158) );
  AND U12783 ( .A(n13159), .B(n13160), .Z(n12841) );
  NANDN U12784 ( .A(n13161), .B(n13162), .Z(n13160) );
  NANDN U12785 ( .A(n13163), .B(n13164), .Z(n13159) );
  NANDN U12786 ( .A(n13162), .B(n13161), .Z(n13164) );
  ANDN U12787 ( .B(\stack[1][43] ), .A(n5374), .Z(n12840) );
  XNOR U12788 ( .A(n12846), .B(n13165), .Z(n12839) );
  XNOR U12789 ( .A(n12847), .B(n12848), .Z(n13165) );
  AND U12790 ( .A(n13166), .B(n13167), .Z(n12848) );
  NAND U12791 ( .A(n13168), .B(n13169), .Z(n13167) );
  NANDN U12792 ( .A(n13170), .B(n13171), .Z(n13166) );
  OR U12793 ( .A(n13168), .B(n13169), .Z(n13171) );
  ANDN U12794 ( .B(\stack[1][44] ), .A(n5350), .Z(n12847) );
  XNOR U12795 ( .A(n12853), .B(n13172), .Z(n12846) );
  XNOR U12796 ( .A(n12854), .B(n12855), .Z(n13172) );
  AND U12797 ( .A(n13173), .B(n13174), .Z(n12855) );
  NANDN U12798 ( .A(n13175), .B(n13176), .Z(n13174) );
  NANDN U12799 ( .A(n13177), .B(n13178), .Z(n13173) );
  NANDN U12800 ( .A(n13176), .B(n13175), .Z(n13178) );
  ANDN U12801 ( .B(\stack[1][45] ), .A(n5326), .Z(n12854) );
  XNOR U12802 ( .A(n12860), .B(n13179), .Z(n12853) );
  XNOR U12803 ( .A(n12861), .B(n12862), .Z(n13179) );
  AND U12804 ( .A(n13180), .B(n13181), .Z(n12862) );
  NAND U12805 ( .A(n13182), .B(n13183), .Z(n13181) );
  NANDN U12806 ( .A(n13184), .B(n13185), .Z(n13180) );
  OR U12807 ( .A(n13182), .B(n13183), .Z(n13185) );
  ANDN U12808 ( .B(\stack[1][46] ), .A(n5302), .Z(n12861) );
  XNOR U12809 ( .A(n12867), .B(n13186), .Z(n12860) );
  XNOR U12810 ( .A(n12868), .B(n12869), .Z(n13186) );
  AND U12811 ( .A(n13187), .B(n13188), .Z(n12869) );
  NANDN U12812 ( .A(n13189), .B(n13190), .Z(n13188) );
  NANDN U12813 ( .A(n13191), .B(n13192), .Z(n13187) );
  NANDN U12814 ( .A(n13190), .B(n13189), .Z(n13192) );
  ANDN U12815 ( .B(\stack[1][47] ), .A(n5278), .Z(n12868) );
  XNOR U12816 ( .A(n12874), .B(n13193), .Z(n12867) );
  XNOR U12817 ( .A(n12875), .B(n12876), .Z(n13193) );
  AND U12818 ( .A(n13194), .B(n13195), .Z(n12876) );
  NAND U12819 ( .A(n13196), .B(n13197), .Z(n13195) );
  NANDN U12820 ( .A(n13198), .B(n13199), .Z(n13194) );
  OR U12821 ( .A(n13196), .B(n13197), .Z(n13199) );
  ANDN U12822 ( .B(\stack[1][48] ), .A(n5254), .Z(n12875) );
  XNOR U12823 ( .A(n12881), .B(n13200), .Z(n12874) );
  XNOR U12824 ( .A(n12882), .B(n12883), .Z(n13200) );
  AND U12825 ( .A(n13201), .B(n13202), .Z(n12883) );
  NAND U12826 ( .A(n13203), .B(n13204), .Z(n13202) );
  NAND U12827 ( .A(n13205), .B(n13206), .Z(n13201) );
  OR U12828 ( .A(n13203), .B(n13204), .Z(n13205) );
  ANDN U12829 ( .B(\stack[1][49] ), .A(n5230), .Z(n12882) );
  XNOR U12830 ( .A(n12888), .B(n13207), .Z(n12881) );
  XNOR U12831 ( .A(n12889), .B(n12891), .Z(n13207) );
  ANDN U12832 ( .B(n13208), .A(n13209), .Z(n12891) );
  ANDN U12833 ( .B(\stack[0][0] ), .A(n6396), .Z(n13208) );
  ANDN U12834 ( .B(\stack[1][50] ), .A(n5206), .Z(n12889) );
  XOR U12835 ( .A(n12894), .B(n13210), .Z(n12888) );
  NANDN U12836 ( .A(n5160), .B(\stack[1][52] ), .Z(n13210) );
  NANDN U12837 ( .A(n6396), .B(\stack[0][1] ), .Z(n12894) );
  ANDN U12838 ( .B(\stack[0][47] ), .A(n5292), .Z(n9034) );
  AND U12839 ( .A(n13211), .B(n13212), .Z(n9035) );
  OR U12840 ( .A(n9039), .B(n13213), .Z(n13212) );
  IV U12841 ( .A(n9041), .Z(n13213) );
  NANDN U12842 ( .A(n9042), .B(n13214), .Z(n13211) );
  NANDN U12843 ( .A(n9041), .B(n9039), .Z(n13214) );
  XNOR U12844 ( .A(n12902), .B(n13215), .Z(n9039) );
  XNOR U12845 ( .A(n12903), .B(n12904), .Z(n13215) );
  AND U12846 ( .A(n13216), .B(n13217), .Z(n12904) );
  NANDN U12847 ( .A(n13218), .B(n13219), .Z(n13217) );
  NANDN U12848 ( .A(n13220), .B(n13221), .Z(n13216) );
  NANDN U12849 ( .A(n13219), .B(n13218), .Z(n13221) );
  ANDN U12850 ( .B(\stack[0][45] ), .A(n5316), .Z(n12903) );
  XNOR U12851 ( .A(n12909), .B(n13222), .Z(n12902) );
  XNOR U12852 ( .A(n12910), .B(n12911), .Z(n13222) );
  AND U12853 ( .A(n13223), .B(n13224), .Z(n12911) );
  NAND U12854 ( .A(n13225), .B(n13226), .Z(n13224) );
  NANDN U12855 ( .A(n13227), .B(n13228), .Z(n13223) );
  OR U12856 ( .A(n13225), .B(n13226), .Z(n13228) );
  ANDN U12857 ( .B(\stack[0][44] ), .A(n5340), .Z(n12910) );
  XNOR U12858 ( .A(n12916), .B(n13229), .Z(n12909) );
  XNOR U12859 ( .A(n12917), .B(n12918), .Z(n13229) );
  AND U12860 ( .A(n13230), .B(n13231), .Z(n12918) );
  NANDN U12861 ( .A(n13232), .B(n13233), .Z(n13231) );
  NANDN U12862 ( .A(n13234), .B(n13235), .Z(n13230) );
  NANDN U12863 ( .A(n13233), .B(n13232), .Z(n13235) );
  ANDN U12864 ( .B(\stack[0][43] ), .A(n5364), .Z(n12917) );
  XNOR U12865 ( .A(n12923), .B(n13236), .Z(n12916) );
  XNOR U12866 ( .A(n12924), .B(n12925), .Z(n13236) );
  AND U12867 ( .A(n13237), .B(n13238), .Z(n12925) );
  NAND U12868 ( .A(n13239), .B(n13240), .Z(n13238) );
  NANDN U12869 ( .A(n13241), .B(n13242), .Z(n13237) );
  OR U12870 ( .A(n13239), .B(n13240), .Z(n13242) );
  ANDN U12871 ( .B(\stack[0][42] ), .A(n5387), .Z(n12924) );
  XNOR U12872 ( .A(n12930), .B(n13243), .Z(n12923) );
  XNOR U12873 ( .A(n12931), .B(n12932), .Z(n13243) );
  AND U12874 ( .A(n13244), .B(n13245), .Z(n12932) );
  NANDN U12875 ( .A(n13246), .B(n13247), .Z(n13245) );
  NANDN U12876 ( .A(n13248), .B(n13249), .Z(n13244) );
  NANDN U12877 ( .A(n13247), .B(n13246), .Z(n13249) );
  ANDN U12878 ( .B(\stack[1][10] ), .A(n6142), .Z(n12931) );
  XNOR U12879 ( .A(n12937), .B(n13250), .Z(n12930) );
  XNOR U12880 ( .A(n12938), .B(n12939), .Z(n13250) );
  AND U12881 ( .A(n13251), .B(n13252), .Z(n12939) );
  NAND U12882 ( .A(n13253), .B(n13254), .Z(n13252) );
  NANDN U12883 ( .A(n13255), .B(n13256), .Z(n13251) );
  OR U12884 ( .A(n13253), .B(n13254), .Z(n13256) );
  ANDN U12885 ( .B(\stack[1][11] ), .A(n6118), .Z(n12938) );
  XNOR U12886 ( .A(n12944), .B(n13257), .Z(n12937) );
  XNOR U12887 ( .A(n12945), .B(n12946), .Z(n13257) );
  AND U12888 ( .A(n13258), .B(n13259), .Z(n12946) );
  NANDN U12889 ( .A(n13260), .B(n13261), .Z(n13259) );
  NANDN U12890 ( .A(n13262), .B(n13263), .Z(n13258) );
  NANDN U12891 ( .A(n13261), .B(n13260), .Z(n13263) );
  ANDN U12892 ( .B(\stack[1][12] ), .A(n6094), .Z(n12945) );
  XNOR U12893 ( .A(n12951), .B(n13264), .Z(n12944) );
  XNOR U12894 ( .A(n12952), .B(n12953), .Z(n13264) );
  AND U12895 ( .A(n13265), .B(n13266), .Z(n12953) );
  NAND U12896 ( .A(n13267), .B(n13268), .Z(n13266) );
  NANDN U12897 ( .A(n13269), .B(n13270), .Z(n13265) );
  OR U12898 ( .A(n13267), .B(n13268), .Z(n13270) );
  ANDN U12899 ( .B(\stack[1][13] ), .A(n6070), .Z(n12952) );
  XNOR U12900 ( .A(n12958), .B(n13271), .Z(n12951) );
  XNOR U12901 ( .A(n12959), .B(n12960), .Z(n13271) );
  AND U12902 ( .A(n13272), .B(n13273), .Z(n12960) );
  NANDN U12903 ( .A(n13274), .B(n13275), .Z(n13273) );
  NANDN U12904 ( .A(n13276), .B(n13277), .Z(n13272) );
  NANDN U12905 ( .A(n13275), .B(n13274), .Z(n13277) );
  ANDN U12906 ( .B(\stack[1][14] ), .A(n6046), .Z(n12959) );
  XNOR U12907 ( .A(n12965), .B(n13278), .Z(n12958) );
  XNOR U12908 ( .A(n12966), .B(n12967), .Z(n13278) );
  AND U12909 ( .A(n13279), .B(n13280), .Z(n12967) );
  NAND U12910 ( .A(n13281), .B(n13282), .Z(n13280) );
  NANDN U12911 ( .A(n13283), .B(n13284), .Z(n13279) );
  OR U12912 ( .A(n13281), .B(n13282), .Z(n13284) );
  ANDN U12913 ( .B(\stack[1][15] ), .A(n6022), .Z(n12966) );
  XNOR U12914 ( .A(n12972), .B(n13285), .Z(n12965) );
  XNOR U12915 ( .A(n12973), .B(n12974), .Z(n13285) );
  AND U12916 ( .A(n13286), .B(n13287), .Z(n12974) );
  NANDN U12917 ( .A(n13288), .B(n13289), .Z(n13287) );
  NANDN U12918 ( .A(n13290), .B(n13291), .Z(n13286) );
  NANDN U12919 ( .A(n13289), .B(n13288), .Z(n13291) );
  ANDN U12920 ( .B(\stack[1][16] ), .A(n5998), .Z(n12973) );
  XNOR U12921 ( .A(n12979), .B(n13292), .Z(n12972) );
  XNOR U12922 ( .A(n12980), .B(n12981), .Z(n13292) );
  AND U12923 ( .A(n13293), .B(n13294), .Z(n12981) );
  NAND U12924 ( .A(n13295), .B(n13296), .Z(n13294) );
  NANDN U12925 ( .A(n13297), .B(n13298), .Z(n13293) );
  OR U12926 ( .A(n13295), .B(n13296), .Z(n13298) );
  ANDN U12927 ( .B(\stack[1][17] ), .A(n5974), .Z(n12980) );
  XNOR U12928 ( .A(n12986), .B(n13299), .Z(n12979) );
  XNOR U12929 ( .A(n12987), .B(n12988), .Z(n13299) );
  AND U12930 ( .A(n13300), .B(n13301), .Z(n12988) );
  NANDN U12931 ( .A(n13302), .B(n13303), .Z(n13301) );
  NANDN U12932 ( .A(n13304), .B(n13305), .Z(n13300) );
  NANDN U12933 ( .A(n13303), .B(n13302), .Z(n13305) );
  ANDN U12934 ( .B(\stack[1][18] ), .A(n5950), .Z(n12987) );
  XNOR U12935 ( .A(n12993), .B(n13306), .Z(n12986) );
  XNOR U12936 ( .A(n12994), .B(n12995), .Z(n13306) );
  AND U12937 ( .A(n13307), .B(n13308), .Z(n12995) );
  NAND U12938 ( .A(n13309), .B(n13310), .Z(n13308) );
  NANDN U12939 ( .A(n13311), .B(n13312), .Z(n13307) );
  OR U12940 ( .A(n13309), .B(n13310), .Z(n13312) );
  ANDN U12941 ( .B(\stack[1][19] ), .A(n5926), .Z(n12994) );
  XNOR U12942 ( .A(n13000), .B(n13313), .Z(n12993) );
  XNOR U12943 ( .A(n13001), .B(n13002), .Z(n13313) );
  AND U12944 ( .A(n13314), .B(n13315), .Z(n13002) );
  NANDN U12945 ( .A(n13316), .B(n13317), .Z(n13315) );
  NANDN U12946 ( .A(n13318), .B(n13319), .Z(n13314) );
  NANDN U12947 ( .A(n13317), .B(n13316), .Z(n13319) );
  ANDN U12948 ( .B(\stack[1][20] ), .A(n5902), .Z(n13001) );
  XNOR U12949 ( .A(n13007), .B(n13320), .Z(n13000) );
  XNOR U12950 ( .A(n13008), .B(n13009), .Z(n13320) );
  AND U12951 ( .A(n13321), .B(n13322), .Z(n13009) );
  NAND U12952 ( .A(n13323), .B(n13324), .Z(n13322) );
  NANDN U12953 ( .A(n13325), .B(n13326), .Z(n13321) );
  OR U12954 ( .A(n13323), .B(n13324), .Z(n13326) );
  ANDN U12955 ( .B(\stack[1][21] ), .A(n5878), .Z(n13008) );
  XNOR U12956 ( .A(n13014), .B(n13327), .Z(n13007) );
  XNOR U12957 ( .A(n13015), .B(n13016), .Z(n13327) );
  AND U12958 ( .A(n13328), .B(n13329), .Z(n13016) );
  NANDN U12959 ( .A(n13330), .B(n13331), .Z(n13329) );
  NANDN U12960 ( .A(n13332), .B(n13333), .Z(n13328) );
  NANDN U12961 ( .A(n13331), .B(n13330), .Z(n13333) );
  ANDN U12962 ( .B(\stack[1][22] ), .A(n5854), .Z(n13015) );
  XNOR U12963 ( .A(n13021), .B(n13334), .Z(n13014) );
  XNOR U12964 ( .A(n13022), .B(n13023), .Z(n13334) );
  AND U12965 ( .A(n13335), .B(n13336), .Z(n13023) );
  NAND U12966 ( .A(n13337), .B(n13338), .Z(n13336) );
  NANDN U12967 ( .A(n13339), .B(n13340), .Z(n13335) );
  OR U12968 ( .A(n13337), .B(n13338), .Z(n13340) );
  ANDN U12969 ( .B(\stack[1][23] ), .A(n5830), .Z(n13022) );
  XNOR U12970 ( .A(n13028), .B(n13341), .Z(n13021) );
  XNOR U12971 ( .A(n13029), .B(n13030), .Z(n13341) );
  AND U12972 ( .A(n13342), .B(n13343), .Z(n13030) );
  NANDN U12973 ( .A(n13344), .B(n13345), .Z(n13343) );
  NANDN U12974 ( .A(n13346), .B(n13347), .Z(n13342) );
  NANDN U12975 ( .A(n13345), .B(n13344), .Z(n13347) );
  ANDN U12976 ( .B(\stack[1][24] ), .A(n5806), .Z(n13029) );
  XNOR U12977 ( .A(n13035), .B(n13348), .Z(n13028) );
  XNOR U12978 ( .A(n13036), .B(n13037), .Z(n13348) );
  AND U12979 ( .A(n13349), .B(n13350), .Z(n13037) );
  NAND U12980 ( .A(n13351), .B(n13352), .Z(n13350) );
  NANDN U12981 ( .A(n13353), .B(n13354), .Z(n13349) );
  OR U12982 ( .A(n13351), .B(n13352), .Z(n13354) );
  ANDN U12983 ( .B(\stack[1][25] ), .A(n5782), .Z(n13036) );
  XNOR U12984 ( .A(n13042), .B(n13355), .Z(n13035) );
  XNOR U12985 ( .A(n13043), .B(n13044), .Z(n13355) );
  AND U12986 ( .A(n13356), .B(n13357), .Z(n13044) );
  NANDN U12987 ( .A(n13358), .B(n13359), .Z(n13357) );
  NANDN U12988 ( .A(n13360), .B(n13361), .Z(n13356) );
  NANDN U12989 ( .A(n13359), .B(n13358), .Z(n13361) );
  ANDN U12990 ( .B(\stack[1][26] ), .A(n5758), .Z(n13043) );
  XNOR U12991 ( .A(n13049), .B(n13362), .Z(n13042) );
  XNOR U12992 ( .A(n13050), .B(n13051), .Z(n13362) );
  AND U12993 ( .A(n13363), .B(n13364), .Z(n13051) );
  NAND U12994 ( .A(n13365), .B(n13366), .Z(n13364) );
  NANDN U12995 ( .A(n13367), .B(n13368), .Z(n13363) );
  OR U12996 ( .A(n13365), .B(n13366), .Z(n13368) );
  ANDN U12997 ( .B(\stack[1][27] ), .A(n5734), .Z(n13050) );
  XNOR U12998 ( .A(n13056), .B(n13369), .Z(n13049) );
  XNOR U12999 ( .A(n13057), .B(n13058), .Z(n13369) );
  AND U13000 ( .A(n13370), .B(n13371), .Z(n13058) );
  NANDN U13001 ( .A(n13372), .B(n13373), .Z(n13371) );
  NANDN U13002 ( .A(n13374), .B(n13375), .Z(n13370) );
  NANDN U13003 ( .A(n13373), .B(n13372), .Z(n13375) );
  ANDN U13004 ( .B(\stack[1][28] ), .A(n5710), .Z(n13057) );
  XNOR U13005 ( .A(n13063), .B(n13376), .Z(n13056) );
  XNOR U13006 ( .A(n13064), .B(n13065), .Z(n13376) );
  AND U13007 ( .A(n13377), .B(n13378), .Z(n13065) );
  NAND U13008 ( .A(n13379), .B(n13380), .Z(n13378) );
  NANDN U13009 ( .A(n13381), .B(n13382), .Z(n13377) );
  OR U13010 ( .A(n13379), .B(n13380), .Z(n13382) );
  ANDN U13011 ( .B(\stack[1][29] ), .A(n5686), .Z(n13064) );
  XNOR U13012 ( .A(n13070), .B(n13383), .Z(n13063) );
  XNOR U13013 ( .A(n13071), .B(n13072), .Z(n13383) );
  AND U13014 ( .A(n13384), .B(n13385), .Z(n13072) );
  NANDN U13015 ( .A(n13386), .B(n13387), .Z(n13385) );
  NANDN U13016 ( .A(n13388), .B(n13389), .Z(n13384) );
  NANDN U13017 ( .A(n13387), .B(n13386), .Z(n13389) );
  ANDN U13018 ( .B(\stack[1][30] ), .A(n5662), .Z(n13071) );
  XNOR U13019 ( .A(n13077), .B(n13390), .Z(n13070) );
  XNOR U13020 ( .A(n13078), .B(n13079), .Z(n13390) );
  AND U13021 ( .A(n13391), .B(n13392), .Z(n13079) );
  NAND U13022 ( .A(n13393), .B(n13394), .Z(n13392) );
  NANDN U13023 ( .A(n13395), .B(n13396), .Z(n13391) );
  OR U13024 ( .A(n13393), .B(n13394), .Z(n13396) );
  ANDN U13025 ( .B(\stack[1][31] ), .A(n5638), .Z(n13078) );
  XNOR U13026 ( .A(n13084), .B(n13397), .Z(n13077) );
  XNOR U13027 ( .A(n13085), .B(n13086), .Z(n13397) );
  AND U13028 ( .A(n13398), .B(n13399), .Z(n13086) );
  NANDN U13029 ( .A(n13400), .B(n13401), .Z(n13399) );
  NANDN U13030 ( .A(n13402), .B(n13403), .Z(n13398) );
  NANDN U13031 ( .A(n13401), .B(n13400), .Z(n13403) );
  ANDN U13032 ( .B(\stack[1][32] ), .A(n5614), .Z(n13085) );
  XNOR U13033 ( .A(n13091), .B(n13404), .Z(n13084) );
  XNOR U13034 ( .A(n13092), .B(n13093), .Z(n13404) );
  AND U13035 ( .A(n13405), .B(n13406), .Z(n13093) );
  NAND U13036 ( .A(n13407), .B(n13408), .Z(n13406) );
  NANDN U13037 ( .A(n13409), .B(n13410), .Z(n13405) );
  OR U13038 ( .A(n13407), .B(n13408), .Z(n13410) );
  ANDN U13039 ( .B(\stack[1][33] ), .A(n5590), .Z(n13092) );
  XNOR U13040 ( .A(n13098), .B(n13411), .Z(n13091) );
  XNOR U13041 ( .A(n13099), .B(n13100), .Z(n13411) );
  AND U13042 ( .A(n13412), .B(n13413), .Z(n13100) );
  NANDN U13043 ( .A(n13414), .B(n13415), .Z(n13413) );
  NANDN U13044 ( .A(n13416), .B(n13417), .Z(n13412) );
  NANDN U13045 ( .A(n13415), .B(n13414), .Z(n13417) );
  ANDN U13046 ( .B(\stack[1][34] ), .A(n5566), .Z(n13099) );
  XNOR U13047 ( .A(n13105), .B(n13418), .Z(n13098) );
  XNOR U13048 ( .A(n13106), .B(n13107), .Z(n13418) );
  AND U13049 ( .A(n13419), .B(n13420), .Z(n13107) );
  NAND U13050 ( .A(n13421), .B(n13422), .Z(n13420) );
  NANDN U13051 ( .A(n13423), .B(n13424), .Z(n13419) );
  OR U13052 ( .A(n13421), .B(n13422), .Z(n13424) );
  ANDN U13053 ( .B(\stack[1][35] ), .A(n5542), .Z(n13106) );
  XNOR U13054 ( .A(n13112), .B(n13425), .Z(n13105) );
  XNOR U13055 ( .A(n13113), .B(n13114), .Z(n13425) );
  AND U13056 ( .A(n13426), .B(n13427), .Z(n13114) );
  NANDN U13057 ( .A(n13428), .B(n13429), .Z(n13427) );
  NANDN U13058 ( .A(n13430), .B(n13431), .Z(n13426) );
  NANDN U13059 ( .A(n13429), .B(n13428), .Z(n13431) );
  ANDN U13060 ( .B(\stack[1][36] ), .A(n5518), .Z(n13113) );
  XNOR U13061 ( .A(n13119), .B(n13432), .Z(n13112) );
  XOR U13062 ( .A(n13121), .B(n13122), .Z(n13432) );
  NAND U13063 ( .A(n13433), .B(n13434), .Z(n13122) );
  NAND U13064 ( .A(n13435), .B(n13436), .Z(n13434) );
  OR U13065 ( .A(n13437), .B(n13438), .Z(n13435) );
  AND U13066 ( .A(\stack[0][14] ), .B(\stack[1][37] ), .Z(n13121) );
  XNOR U13067 ( .A(n13128), .B(n13439), .Z(n13119) );
  XOR U13068 ( .A(n13129), .B(n13127), .Z(n13439) );
  AND U13069 ( .A(\stack[0][13] ), .B(\stack[1][38] ), .Z(n13127) );
  NAND U13070 ( .A(n13440), .B(n13441), .Z(n13129) );
  OR U13071 ( .A(n13442), .B(n13443), .Z(n13441) );
  NAND U13072 ( .A(n13444), .B(n13445), .Z(n13440) );
  NAND U13073 ( .A(n13443), .B(n13442), .Z(n13444) );
  XNOR U13074 ( .A(n13133), .B(n13446), .Z(n13128) );
  XNOR U13075 ( .A(n13134), .B(n13135), .Z(n13446) );
  AND U13076 ( .A(n13447), .B(n13448), .Z(n13135) );
  NAND U13077 ( .A(n13449), .B(n13450), .Z(n13448) );
  NANDN U13078 ( .A(n13451), .B(n13452), .Z(n13447) );
  OR U13079 ( .A(n13449), .B(n13450), .Z(n13452) );
  ANDN U13080 ( .B(\stack[1][39] ), .A(n5446), .Z(n13134) );
  XNOR U13081 ( .A(n13140), .B(n13453), .Z(n13133) );
  XNOR U13082 ( .A(n13141), .B(n13142), .Z(n13453) );
  AND U13083 ( .A(n13454), .B(n13455), .Z(n13142) );
  NANDN U13084 ( .A(n13456), .B(n13457), .Z(n13455) );
  NANDN U13085 ( .A(n13458), .B(n13459), .Z(n13454) );
  NANDN U13086 ( .A(n13457), .B(n13456), .Z(n13459) );
  ANDN U13087 ( .B(\stack[1][40] ), .A(n5422), .Z(n13141) );
  XNOR U13088 ( .A(n13147), .B(n13460), .Z(n13140) );
  XNOR U13089 ( .A(n13148), .B(n13149), .Z(n13460) );
  AND U13090 ( .A(n13461), .B(n13462), .Z(n13149) );
  NAND U13091 ( .A(n13463), .B(n13464), .Z(n13462) );
  NANDN U13092 ( .A(n13465), .B(n13466), .Z(n13461) );
  OR U13093 ( .A(n13463), .B(n13464), .Z(n13466) );
  ANDN U13094 ( .B(\stack[1][41] ), .A(n5398), .Z(n13148) );
  XNOR U13095 ( .A(n13154), .B(n13467), .Z(n13147) );
  XNOR U13096 ( .A(n13155), .B(n13156), .Z(n13467) );
  AND U13097 ( .A(n13468), .B(n13469), .Z(n13156) );
  NANDN U13098 ( .A(n13470), .B(n13471), .Z(n13469) );
  NANDN U13099 ( .A(n13472), .B(n13473), .Z(n13468) );
  NANDN U13100 ( .A(n13471), .B(n13470), .Z(n13473) );
  ANDN U13101 ( .B(\stack[1][42] ), .A(n5374), .Z(n13155) );
  XNOR U13102 ( .A(n13161), .B(n13474), .Z(n13154) );
  XNOR U13103 ( .A(n13162), .B(n13163), .Z(n13474) );
  AND U13104 ( .A(n13475), .B(n13476), .Z(n13163) );
  NAND U13105 ( .A(n13477), .B(n13478), .Z(n13476) );
  NANDN U13106 ( .A(n13479), .B(n13480), .Z(n13475) );
  OR U13107 ( .A(n13477), .B(n13478), .Z(n13480) );
  ANDN U13108 ( .B(\stack[1][43] ), .A(n5350), .Z(n13162) );
  XNOR U13109 ( .A(n13168), .B(n13481), .Z(n13161) );
  XNOR U13110 ( .A(n13169), .B(n13170), .Z(n13481) );
  AND U13111 ( .A(n13482), .B(n13483), .Z(n13170) );
  NANDN U13112 ( .A(n13484), .B(n13485), .Z(n13483) );
  NANDN U13113 ( .A(n13486), .B(n13487), .Z(n13482) );
  NANDN U13114 ( .A(n13485), .B(n13484), .Z(n13487) );
  ANDN U13115 ( .B(\stack[1][44] ), .A(n5326), .Z(n13169) );
  XNOR U13116 ( .A(n13175), .B(n13488), .Z(n13168) );
  XNOR U13117 ( .A(n13176), .B(n13177), .Z(n13488) );
  AND U13118 ( .A(n13489), .B(n13490), .Z(n13177) );
  NAND U13119 ( .A(n13491), .B(n13492), .Z(n13490) );
  NANDN U13120 ( .A(n13493), .B(n13494), .Z(n13489) );
  OR U13121 ( .A(n13491), .B(n13492), .Z(n13494) );
  ANDN U13122 ( .B(\stack[1][45] ), .A(n5302), .Z(n13176) );
  XNOR U13123 ( .A(n13182), .B(n13495), .Z(n13175) );
  XNOR U13124 ( .A(n13183), .B(n13184), .Z(n13495) );
  AND U13125 ( .A(n13496), .B(n13497), .Z(n13184) );
  NANDN U13126 ( .A(n13498), .B(n13499), .Z(n13497) );
  NANDN U13127 ( .A(n13500), .B(n13501), .Z(n13496) );
  NANDN U13128 ( .A(n13499), .B(n13498), .Z(n13501) );
  ANDN U13129 ( .B(\stack[1][46] ), .A(n5278), .Z(n13183) );
  XNOR U13130 ( .A(n13189), .B(n13502), .Z(n13182) );
  XNOR U13131 ( .A(n13190), .B(n13191), .Z(n13502) );
  AND U13132 ( .A(n13503), .B(n13504), .Z(n13191) );
  NAND U13133 ( .A(n13505), .B(n13506), .Z(n13504) );
  NANDN U13134 ( .A(n13507), .B(n13508), .Z(n13503) );
  OR U13135 ( .A(n13505), .B(n13506), .Z(n13508) );
  ANDN U13136 ( .B(\stack[1][47] ), .A(n5254), .Z(n13190) );
  XNOR U13137 ( .A(n13196), .B(n13509), .Z(n13189) );
  XNOR U13138 ( .A(n13197), .B(n13198), .Z(n13509) );
  AND U13139 ( .A(n13510), .B(n13511), .Z(n13198) );
  NAND U13140 ( .A(n13512), .B(n13513), .Z(n13511) );
  NAND U13141 ( .A(n13514), .B(n13515), .Z(n13510) );
  OR U13142 ( .A(n13512), .B(n13513), .Z(n13514) );
  ANDN U13143 ( .B(\stack[1][48] ), .A(n5230), .Z(n13197) );
  XNOR U13144 ( .A(n13203), .B(n13516), .Z(n13196) );
  XNOR U13145 ( .A(n13204), .B(n13206), .Z(n13516) );
  ANDN U13146 ( .B(n13517), .A(n13518), .Z(n13206) );
  ANDN U13147 ( .B(\stack[0][0] ), .A(n6372), .Z(n13517) );
  ANDN U13148 ( .B(\stack[1][49] ), .A(n5206), .Z(n13204) );
  XOR U13149 ( .A(n13209), .B(n13519), .Z(n13203) );
  NANDN U13150 ( .A(n5160), .B(\stack[1][51] ), .Z(n13519) );
  NANDN U13151 ( .A(n6372), .B(\stack[0][1] ), .Z(n13209) );
  ANDN U13152 ( .B(\stack[1][5] ), .A(n6262), .Z(n9041) );
  AND U13153 ( .A(n13520), .B(n13521), .Z(n9042) );
  NANDN U13154 ( .A(n9046), .B(n9048), .Z(n13521) );
  NANDN U13155 ( .A(n9049), .B(n13522), .Z(n13520) );
  NANDN U13156 ( .A(n9048), .B(n9046), .Z(n13522) );
  XOR U13157 ( .A(n13218), .B(n13523), .Z(n9046) );
  XNOR U13158 ( .A(n13219), .B(n13220), .Z(n13523) );
  AND U13159 ( .A(n13524), .B(n13525), .Z(n13220) );
  NAND U13160 ( .A(n13526), .B(n13527), .Z(n13525) );
  NANDN U13161 ( .A(n13528), .B(n13529), .Z(n13524) );
  OR U13162 ( .A(n13526), .B(n13527), .Z(n13529) );
  ANDN U13163 ( .B(\stack[0][44] ), .A(n5316), .Z(n13219) );
  XNOR U13164 ( .A(n13225), .B(n13530), .Z(n13218) );
  XNOR U13165 ( .A(n13226), .B(n13227), .Z(n13530) );
  AND U13166 ( .A(n13531), .B(n13532), .Z(n13227) );
  NANDN U13167 ( .A(n13533), .B(n13534), .Z(n13532) );
  NANDN U13168 ( .A(n13535), .B(n13536), .Z(n13531) );
  NANDN U13169 ( .A(n13534), .B(n13533), .Z(n13536) );
  ANDN U13170 ( .B(\stack[0][43] ), .A(n5340), .Z(n13226) );
  XNOR U13171 ( .A(n13232), .B(n13537), .Z(n13225) );
  XNOR U13172 ( .A(n13233), .B(n13234), .Z(n13537) );
  AND U13173 ( .A(n13538), .B(n13539), .Z(n13234) );
  NAND U13174 ( .A(n13540), .B(n13541), .Z(n13539) );
  NANDN U13175 ( .A(n13542), .B(n13543), .Z(n13538) );
  OR U13176 ( .A(n13540), .B(n13541), .Z(n13543) );
  ANDN U13177 ( .B(\stack[0][42] ), .A(n5364), .Z(n13233) );
  XNOR U13178 ( .A(n13239), .B(n13544), .Z(n13232) );
  XNOR U13179 ( .A(n13240), .B(n13241), .Z(n13544) );
  AND U13180 ( .A(n13545), .B(n13546), .Z(n13241) );
  NANDN U13181 ( .A(n13547), .B(n13548), .Z(n13546) );
  NANDN U13182 ( .A(n13549), .B(n13550), .Z(n13545) );
  NANDN U13183 ( .A(n13548), .B(n13547), .Z(n13550) );
  ANDN U13184 ( .B(\stack[0][41] ), .A(n5387), .Z(n13240) );
  XNOR U13185 ( .A(n13246), .B(n13551), .Z(n13239) );
  XNOR U13186 ( .A(n13247), .B(n13248), .Z(n13551) );
  AND U13187 ( .A(n13552), .B(n13553), .Z(n13248) );
  NAND U13188 ( .A(n13554), .B(n13555), .Z(n13553) );
  NANDN U13189 ( .A(n13556), .B(n13557), .Z(n13552) );
  OR U13190 ( .A(n13554), .B(n13555), .Z(n13557) );
  ANDN U13191 ( .B(\stack[1][10] ), .A(n6118), .Z(n13247) );
  XNOR U13192 ( .A(n13253), .B(n13558), .Z(n13246) );
  XNOR U13193 ( .A(n13254), .B(n13255), .Z(n13558) );
  AND U13194 ( .A(n13559), .B(n13560), .Z(n13255) );
  NANDN U13195 ( .A(n13561), .B(n13562), .Z(n13560) );
  NANDN U13196 ( .A(n13563), .B(n13564), .Z(n13559) );
  NANDN U13197 ( .A(n13562), .B(n13561), .Z(n13564) );
  ANDN U13198 ( .B(\stack[1][11] ), .A(n6094), .Z(n13254) );
  XNOR U13199 ( .A(n13260), .B(n13565), .Z(n13253) );
  XNOR U13200 ( .A(n13261), .B(n13262), .Z(n13565) );
  AND U13201 ( .A(n13566), .B(n13567), .Z(n13262) );
  NAND U13202 ( .A(n13568), .B(n13569), .Z(n13567) );
  NANDN U13203 ( .A(n13570), .B(n13571), .Z(n13566) );
  OR U13204 ( .A(n13568), .B(n13569), .Z(n13571) );
  ANDN U13205 ( .B(\stack[1][12] ), .A(n6070), .Z(n13261) );
  XNOR U13206 ( .A(n13267), .B(n13572), .Z(n13260) );
  XNOR U13207 ( .A(n13268), .B(n13269), .Z(n13572) );
  AND U13208 ( .A(n13573), .B(n13574), .Z(n13269) );
  NANDN U13209 ( .A(n13575), .B(n13576), .Z(n13574) );
  NANDN U13210 ( .A(n13577), .B(n13578), .Z(n13573) );
  NANDN U13211 ( .A(n13576), .B(n13575), .Z(n13578) );
  ANDN U13212 ( .B(\stack[1][13] ), .A(n6046), .Z(n13268) );
  XNOR U13213 ( .A(n13274), .B(n13579), .Z(n13267) );
  XNOR U13214 ( .A(n13275), .B(n13276), .Z(n13579) );
  AND U13215 ( .A(n13580), .B(n13581), .Z(n13276) );
  NAND U13216 ( .A(n13582), .B(n13583), .Z(n13581) );
  NANDN U13217 ( .A(n13584), .B(n13585), .Z(n13580) );
  OR U13218 ( .A(n13582), .B(n13583), .Z(n13585) );
  ANDN U13219 ( .B(\stack[1][14] ), .A(n6022), .Z(n13275) );
  XNOR U13220 ( .A(n13281), .B(n13586), .Z(n13274) );
  XNOR U13221 ( .A(n13282), .B(n13283), .Z(n13586) );
  AND U13222 ( .A(n13587), .B(n13588), .Z(n13283) );
  NANDN U13223 ( .A(n13589), .B(n13590), .Z(n13588) );
  NANDN U13224 ( .A(n13591), .B(n13592), .Z(n13587) );
  NANDN U13225 ( .A(n13590), .B(n13589), .Z(n13592) );
  ANDN U13226 ( .B(\stack[1][15] ), .A(n5998), .Z(n13282) );
  XNOR U13227 ( .A(n13288), .B(n13593), .Z(n13281) );
  XNOR U13228 ( .A(n13289), .B(n13290), .Z(n13593) );
  AND U13229 ( .A(n13594), .B(n13595), .Z(n13290) );
  NAND U13230 ( .A(n13596), .B(n13597), .Z(n13595) );
  NANDN U13231 ( .A(n13598), .B(n13599), .Z(n13594) );
  OR U13232 ( .A(n13596), .B(n13597), .Z(n13599) );
  ANDN U13233 ( .B(\stack[1][16] ), .A(n5974), .Z(n13289) );
  XNOR U13234 ( .A(n13295), .B(n13600), .Z(n13288) );
  XNOR U13235 ( .A(n13296), .B(n13297), .Z(n13600) );
  AND U13236 ( .A(n13601), .B(n13602), .Z(n13297) );
  NANDN U13237 ( .A(n13603), .B(n13604), .Z(n13602) );
  NANDN U13238 ( .A(n13605), .B(n13606), .Z(n13601) );
  NANDN U13239 ( .A(n13604), .B(n13603), .Z(n13606) );
  ANDN U13240 ( .B(\stack[1][17] ), .A(n5950), .Z(n13296) );
  XNOR U13241 ( .A(n13302), .B(n13607), .Z(n13295) );
  XNOR U13242 ( .A(n13303), .B(n13304), .Z(n13607) );
  AND U13243 ( .A(n13608), .B(n13609), .Z(n13304) );
  NAND U13244 ( .A(n13610), .B(n13611), .Z(n13609) );
  NANDN U13245 ( .A(n13612), .B(n13613), .Z(n13608) );
  OR U13246 ( .A(n13610), .B(n13611), .Z(n13613) );
  ANDN U13247 ( .B(\stack[1][18] ), .A(n5926), .Z(n13303) );
  XNOR U13248 ( .A(n13309), .B(n13614), .Z(n13302) );
  XNOR U13249 ( .A(n13310), .B(n13311), .Z(n13614) );
  AND U13250 ( .A(n13615), .B(n13616), .Z(n13311) );
  NANDN U13251 ( .A(n13617), .B(n13618), .Z(n13616) );
  NANDN U13252 ( .A(n13619), .B(n13620), .Z(n13615) );
  NANDN U13253 ( .A(n13618), .B(n13617), .Z(n13620) );
  ANDN U13254 ( .B(\stack[1][19] ), .A(n5902), .Z(n13310) );
  XNOR U13255 ( .A(n13316), .B(n13621), .Z(n13309) );
  XNOR U13256 ( .A(n13317), .B(n13318), .Z(n13621) );
  AND U13257 ( .A(n13622), .B(n13623), .Z(n13318) );
  NAND U13258 ( .A(n13624), .B(n13625), .Z(n13623) );
  NANDN U13259 ( .A(n13626), .B(n13627), .Z(n13622) );
  OR U13260 ( .A(n13624), .B(n13625), .Z(n13627) );
  ANDN U13261 ( .B(\stack[1][20] ), .A(n5878), .Z(n13317) );
  XNOR U13262 ( .A(n13323), .B(n13628), .Z(n13316) );
  XNOR U13263 ( .A(n13324), .B(n13325), .Z(n13628) );
  AND U13264 ( .A(n13629), .B(n13630), .Z(n13325) );
  NANDN U13265 ( .A(n13631), .B(n13632), .Z(n13630) );
  NANDN U13266 ( .A(n13633), .B(n13634), .Z(n13629) );
  NANDN U13267 ( .A(n13632), .B(n13631), .Z(n13634) );
  ANDN U13268 ( .B(\stack[1][21] ), .A(n5854), .Z(n13324) );
  XNOR U13269 ( .A(n13330), .B(n13635), .Z(n13323) );
  XNOR U13270 ( .A(n13331), .B(n13332), .Z(n13635) );
  AND U13271 ( .A(n13636), .B(n13637), .Z(n13332) );
  NAND U13272 ( .A(n13638), .B(n13639), .Z(n13637) );
  NANDN U13273 ( .A(n13640), .B(n13641), .Z(n13636) );
  OR U13274 ( .A(n13638), .B(n13639), .Z(n13641) );
  ANDN U13275 ( .B(\stack[1][22] ), .A(n5830), .Z(n13331) );
  XNOR U13276 ( .A(n13337), .B(n13642), .Z(n13330) );
  XNOR U13277 ( .A(n13338), .B(n13339), .Z(n13642) );
  AND U13278 ( .A(n13643), .B(n13644), .Z(n13339) );
  NANDN U13279 ( .A(n13645), .B(n13646), .Z(n13644) );
  NANDN U13280 ( .A(n13647), .B(n13648), .Z(n13643) );
  NANDN U13281 ( .A(n13646), .B(n13645), .Z(n13648) );
  ANDN U13282 ( .B(\stack[1][23] ), .A(n5806), .Z(n13338) );
  XNOR U13283 ( .A(n13344), .B(n13649), .Z(n13337) );
  XNOR U13284 ( .A(n13345), .B(n13346), .Z(n13649) );
  AND U13285 ( .A(n13650), .B(n13651), .Z(n13346) );
  NAND U13286 ( .A(n13652), .B(n13653), .Z(n13651) );
  NANDN U13287 ( .A(n13654), .B(n13655), .Z(n13650) );
  OR U13288 ( .A(n13652), .B(n13653), .Z(n13655) );
  ANDN U13289 ( .B(\stack[1][24] ), .A(n5782), .Z(n13345) );
  XNOR U13290 ( .A(n13351), .B(n13656), .Z(n13344) );
  XNOR U13291 ( .A(n13352), .B(n13353), .Z(n13656) );
  AND U13292 ( .A(n13657), .B(n13658), .Z(n13353) );
  NANDN U13293 ( .A(n13659), .B(n13660), .Z(n13658) );
  NANDN U13294 ( .A(n13661), .B(n13662), .Z(n13657) );
  NANDN U13295 ( .A(n13660), .B(n13659), .Z(n13662) );
  ANDN U13296 ( .B(\stack[1][25] ), .A(n5758), .Z(n13352) );
  XNOR U13297 ( .A(n13358), .B(n13663), .Z(n13351) );
  XNOR U13298 ( .A(n13359), .B(n13360), .Z(n13663) );
  AND U13299 ( .A(n13664), .B(n13665), .Z(n13360) );
  NAND U13300 ( .A(n13666), .B(n13667), .Z(n13665) );
  NANDN U13301 ( .A(n13668), .B(n13669), .Z(n13664) );
  OR U13302 ( .A(n13666), .B(n13667), .Z(n13669) );
  ANDN U13303 ( .B(\stack[1][26] ), .A(n5734), .Z(n13359) );
  XNOR U13304 ( .A(n13365), .B(n13670), .Z(n13358) );
  XNOR U13305 ( .A(n13366), .B(n13367), .Z(n13670) );
  AND U13306 ( .A(n13671), .B(n13672), .Z(n13367) );
  NANDN U13307 ( .A(n13673), .B(n13674), .Z(n13672) );
  NANDN U13308 ( .A(n13675), .B(n13676), .Z(n13671) );
  NANDN U13309 ( .A(n13674), .B(n13673), .Z(n13676) );
  ANDN U13310 ( .B(\stack[1][27] ), .A(n5710), .Z(n13366) );
  XNOR U13311 ( .A(n13372), .B(n13677), .Z(n13365) );
  XNOR U13312 ( .A(n13373), .B(n13374), .Z(n13677) );
  AND U13313 ( .A(n13678), .B(n13679), .Z(n13374) );
  NAND U13314 ( .A(n13680), .B(n13681), .Z(n13679) );
  NANDN U13315 ( .A(n13682), .B(n13683), .Z(n13678) );
  OR U13316 ( .A(n13680), .B(n13681), .Z(n13683) );
  ANDN U13317 ( .B(\stack[1][28] ), .A(n5686), .Z(n13373) );
  XNOR U13318 ( .A(n13379), .B(n13684), .Z(n13372) );
  XNOR U13319 ( .A(n13380), .B(n13381), .Z(n13684) );
  AND U13320 ( .A(n13685), .B(n13686), .Z(n13381) );
  NANDN U13321 ( .A(n13687), .B(n13688), .Z(n13686) );
  NANDN U13322 ( .A(n13689), .B(n13690), .Z(n13685) );
  NANDN U13323 ( .A(n13688), .B(n13687), .Z(n13690) );
  ANDN U13324 ( .B(\stack[1][29] ), .A(n5662), .Z(n13380) );
  XNOR U13325 ( .A(n13386), .B(n13691), .Z(n13379) );
  XNOR U13326 ( .A(n13387), .B(n13388), .Z(n13691) );
  AND U13327 ( .A(n13692), .B(n13693), .Z(n13388) );
  NAND U13328 ( .A(n13694), .B(n13695), .Z(n13693) );
  NANDN U13329 ( .A(n13696), .B(n13697), .Z(n13692) );
  OR U13330 ( .A(n13694), .B(n13695), .Z(n13697) );
  ANDN U13331 ( .B(\stack[1][30] ), .A(n5638), .Z(n13387) );
  XNOR U13332 ( .A(n13393), .B(n13698), .Z(n13386) );
  XNOR U13333 ( .A(n13394), .B(n13395), .Z(n13698) );
  AND U13334 ( .A(n13699), .B(n13700), .Z(n13395) );
  NANDN U13335 ( .A(n13701), .B(n13702), .Z(n13700) );
  NANDN U13336 ( .A(n13703), .B(n13704), .Z(n13699) );
  NANDN U13337 ( .A(n13702), .B(n13701), .Z(n13704) );
  ANDN U13338 ( .B(\stack[1][31] ), .A(n5614), .Z(n13394) );
  XNOR U13339 ( .A(n13400), .B(n13705), .Z(n13393) );
  XNOR U13340 ( .A(n13401), .B(n13402), .Z(n13705) );
  AND U13341 ( .A(n13706), .B(n13707), .Z(n13402) );
  NAND U13342 ( .A(n13708), .B(n13709), .Z(n13707) );
  NANDN U13343 ( .A(n13710), .B(n13711), .Z(n13706) );
  OR U13344 ( .A(n13708), .B(n13709), .Z(n13711) );
  ANDN U13345 ( .B(\stack[1][32] ), .A(n5590), .Z(n13401) );
  XNOR U13346 ( .A(n13407), .B(n13712), .Z(n13400) );
  XNOR U13347 ( .A(n13408), .B(n13409), .Z(n13712) );
  AND U13348 ( .A(n13713), .B(n13714), .Z(n13409) );
  NANDN U13349 ( .A(n13715), .B(n13716), .Z(n13714) );
  NANDN U13350 ( .A(n13717), .B(n13718), .Z(n13713) );
  NANDN U13351 ( .A(n13716), .B(n13715), .Z(n13718) );
  ANDN U13352 ( .B(\stack[1][33] ), .A(n5566), .Z(n13408) );
  XNOR U13353 ( .A(n13414), .B(n13719), .Z(n13407) );
  XNOR U13354 ( .A(n13415), .B(n13416), .Z(n13719) );
  AND U13355 ( .A(n13720), .B(n13721), .Z(n13416) );
  NAND U13356 ( .A(n13722), .B(n13723), .Z(n13721) );
  NANDN U13357 ( .A(n13724), .B(n13725), .Z(n13720) );
  OR U13358 ( .A(n13722), .B(n13723), .Z(n13725) );
  ANDN U13359 ( .B(\stack[1][34] ), .A(n5542), .Z(n13415) );
  XNOR U13360 ( .A(n13421), .B(n13726), .Z(n13414) );
  XNOR U13361 ( .A(n13422), .B(n13423), .Z(n13726) );
  AND U13362 ( .A(n13727), .B(n13728), .Z(n13423) );
  NANDN U13363 ( .A(n13729), .B(n13730), .Z(n13728) );
  NANDN U13364 ( .A(n13731), .B(n13732), .Z(n13727) );
  NANDN U13365 ( .A(n13730), .B(n13729), .Z(n13732) );
  ANDN U13366 ( .B(\stack[1][35] ), .A(n5518), .Z(n13422) );
  XNOR U13367 ( .A(n13428), .B(n13733), .Z(n13421) );
  XNOR U13368 ( .A(n13429), .B(n13430), .Z(n13733) );
  AND U13369 ( .A(n13734), .B(n13735), .Z(n13430) );
  NAND U13370 ( .A(n13736), .B(n13737), .Z(n13735) );
  NANDN U13371 ( .A(n13738), .B(n13739), .Z(n13734) );
  OR U13372 ( .A(n13736), .B(n13737), .Z(n13739) );
  ANDN U13373 ( .B(\stack[1][36] ), .A(n5494), .Z(n13429) );
  XNOR U13374 ( .A(n13436), .B(n13740), .Z(n13428) );
  XOR U13375 ( .A(n13437), .B(n13438), .Z(n13740) );
  NAND U13376 ( .A(n13741), .B(n13742), .Z(n13438) );
  NANDN U13377 ( .A(n13743), .B(n13744), .Z(n13742) );
  OR U13378 ( .A(n13745), .B(n13746), .Z(n13744) );
  AND U13379 ( .A(\stack[0][13] ), .B(\stack[1][37] ), .Z(n13437) );
  XNOR U13380 ( .A(n13443), .B(n13747), .Z(n13436) );
  XNOR U13381 ( .A(n13442), .B(n13445), .Z(n13747) );
  AND U13382 ( .A(\stack[0][12] ), .B(\stack[1][38] ), .Z(n13445) );
  AND U13383 ( .A(n13748), .B(n13749), .Z(n13442) );
  NAND U13384 ( .A(n13750), .B(n13751), .Z(n13749) );
  OR U13385 ( .A(n13752), .B(n13753), .Z(n13750) );
  XNOR U13386 ( .A(n13449), .B(n13754), .Z(n13443) );
  XNOR U13387 ( .A(n13450), .B(n13451), .Z(n13754) );
  AND U13388 ( .A(n13755), .B(n13756), .Z(n13451) );
  NANDN U13389 ( .A(n13757), .B(n13758), .Z(n13756) );
  NANDN U13390 ( .A(n13759), .B(n13760), .Z(n13755) );
  NANDN U13391 ( .A(n13758), .B(n13757), .Z(n13760) );
  ANDN U13392 ( .B(\stack[1][39] ), .A(n5422), .Z(n13450) );
  XNOR U13393 ( .A(n13456), .B(n13761), .Z(n13449) );
  XNOR U13394 ( .A(n13457), .B(n13458), .Z(n13761) );
  AND U13395 ( .A(n13762), .B(n13763), .Z(n13458) );
  NAND U13396 ( .A(n13764), .B(n13765), .Z(n13763) );
  NANDN U13397 ( .A(n13766), .B(n13767), .Z(n13762) );
  OR U13398 ( .A(n13764), .B(n13765), .Z(n13767) );
  ANDN U13399 ( .B(\stack[1][40] ), .A(n5398), .Z(n13457) );
  XNOR U13400 ( .A(n13463), .B(n13768), .Z(n13456) );
  XNOR U13401 ( .A(n13464), .B(n13465), .Z(n13768) );
  AND U13402 ( .A(n13769), .B(n13770), .Z(n13465) );
  NANDN U13403 ( .A(n13771), .B(n13772), .Z(n13770) );
  NANDN U13404 ( .A(n13773), .B(n13774), .Z(n13769) );
  NANDN U13405 ( .A(n13772), .B(n13771), .Z(n13774) );
  ANDN U13406 ( .B(\stack[1][41] ), .A(n5374), .Z(n13464) );
  XNOR U13407 ( .A(n13470), .B(n13775), .Z(n13463) );
  XNOR U13408 ( .A(n13471), .B(n13472), .Z(n13775) );
  AND U13409 ( .A(n13776), .B(n13777), .Z(n13472) );
  NAND U13410 ( .A(n13778), .B(n13779), .Z(n13777) );
  NANDN U13411 ( .A(n13780), .B(n13781), .Z(n13776) );
  OR U13412 ( .A(n13778), .B(n13779), .Z(n13781) );
  ANDN U13413 ( .B(\stack[1][42] ), .A(n5350), .Z(n13471) );
  XNOR U13414 ( .A(n13477), .B(n13782), .Z(n13470) );
  XNOR U13415 ( .A(n13478), .B(n13479), .Z(n13782) );
  AND U13416 ( .A(n13783), .B(n13784), .Z(n13479) );
  NANDN U13417 ( .A(n13785), .B(n13786), .Z(n13784) );
  NANDN U13418 ( .A(n13787), .B(n13788), .Z(n13783) );
  NANDN U13419 ( .A(n13786), .B(n13785), .Z(n13788) );
  ANDN U13420 ( .B(\stack[1][43] ), .A(n5326), .Z(n13478) );
  XNOR U13421 ( .A(n13484), .B(n13789), .Z(n13477) );
  XNOR U13422 ( .A(n13485), .B(n13486), .Z(n13789) );
  AND U13423 ( .A(n13790), .B(n13791), .Z(n13486) );
  NAND U13424 ( .A(n13792), .B(n13793), .Z(n13791) );
  NANDN U13425 ( .A(n13794), .B(n13795), .Z(n13790) );
  OR U13426 ( .A(n13792), .B(n13793), .Z(n13795) );
  ANDN U13427 ( .B(\stack[1][44] ), .A(n5302), .Z(n13485) );
  XNOR U13428 ( .A(n13491), .B(n13796), .Z(n13484) );
  XNOR U13429 ( .A(n13492), .B(n13493), .Z(n13796) );
  AND U13430 ( .A(n13797), .B(n13798), .Z(n13493) );
  NANDN U13431 ( .A(n13799), .B(n13800), .Z(n13798) );
  NANDN U13432 ( .A(n13801), .B(n13802), .Z(n13797) );
  NANDN U13433 ( .A(n13800), .B(n13799), .Z(n13802) );
  ANDN U13434 ( .B(\stack[1][45] ), .A(n5278), .Z(n13492) );
  XNOR U13435 ( .A(n13498), .B(n13803), .Z(n13491) );
  XNOR U13436 ( .A(n13499), .B(n13500), .Z(n13803) );
  AND U13437 ( .A(n13804), .B(n13805), .Z(n13500) );
  NAND U13438 ( .A(n13806), .B(n13807), .Z(n13805) );
  NANDN U13439 ( .A(n13808), .B(n13809), .Z(n13804) );
  OR U13440 ( .A(n13806), .B(n13807), .Z(n13809) );
  ANDN U13441 ( .B(\stack[1][46] ), .A(n5254), .Z(n13499) );
  XNOR U13442 ( .A(n13505), .B(n13810), .Z(n13498) );
  XNOR U13443 ( .A(n13506), .B(n13507), .Z(n13810) );
  AND U13444 ( .A(n13811), .B(n13812), .Z(n13507) );
  NAND U13445 ( .A(n13813), .B(n13814), .Z(n13812) );
  NAND U13446 ( .A(n13815), .B(n13816), .Z(n13811) );
  OR U13447 ( .A(n13813), .B(n13814), .Z(n13815) );
  ANDN U13448 ( .B(\stack[1][47] ), .A(n5230), .Z(n13506) );
  XNOR U13449 ( .A(n13512), .B(n13817), .Z(n13505) );
  XNOR U13450 ( .A(n13513), .B(n13515), .Z(n13817) );
  ANDN U13451 ( .B(n13818), .A(n13819), .Z(n13515) );
  ANDN U13452 ( .B(\stack[0][0] ), .A(n6348), .Z(n13818) );
  ANDN U13453 ( .B(\stack[1][48] ), .A(n5206), .Z(n13513) );
  XOR U13454 ( .A(n13518), .B(n13820), .Z(n13512) );
  NANDN U13455 ( .A(n5160), .B(\stack[1][50] ), .Z(n13820) );
  NANDN U13456 ( .A(n6348), .B(\stack[0][1] ), .Z(n13518) );
  ANDN U13457 ( .B(\stack[0][45] ), .A(n5292), .Z(n9048) );
  AND U13458 ( .A(n13821), .B(n13822), .Z(n9049) );
  NANDN U13459 ( .A(n9056), .B(n13823), .Z(n13821) );
  NANDN U13460 ( .A(n9055), .B(n9053), .Z(n13823) );
  XNOR U13461 ( .A(n13526), .B(n13824), .Z(n9053) );
  XNOR U13462 ( .A(n13527), .B(n13528), .Z(n13824) );
  AND U13463 ( .A(n13825), .B(n13826), .Z(n13528) );
  NANDN U13464 ( .A(n13827), .B(n13828), .Z(n13826) );
  NANDN U13465 ( .A(n13829), .B(n13830), .Z(n13825) );
  NANDN U13466 ( .A(n13828), .B(n13827), .Z(n13830) );
  ANDN U13467 ( .B(\stack[0][43] ), .A(n5316), .Z(n13527) );
  XNOR U13468 ( .A(n13533), .B(n13831), .Z(n13526) );
  XNOR U13469 ( .A(n13534), .B(n13535), .Z(n13831) );
  AND U13470 ( .A(n13832), .B(n13833), .Z(n13535) );
  NAND U13471 ( .A(n13834), .B(n13835), .Z(n13833) );
  NANDN U13472 ( .A(n13836), .B(n13837), .Z(n13832) );
  OR U13473 ( .A(n13834), .B(n13835), .Z(n13837) );
  ANDN U13474 ( .B(\stack[0][42] ), .A(n5340), .Z(n13534) );
  XNOR U13475 ( .A(n13540), .B(n13838), .Z(n13533) );
  XNOR U13476 ( .A(n13541), .B(n13542), .Z(n13838) );
  AND U13477 ( .A(n13839), .B(n13840), .Z(n13542) );
  NANDN U13478 ( .A(n13841), .B(n13842), .Z(n13840) );
  NANDN U13479 ( .A(n13843), .B(n13844), .Z(n13839) );
  NANDN U13480 ( .A(n13842), .B(n13841), .Z(n13844) );
  ANDN U13481 ( .B(\stack[0][41] ), .A(n5364), .Z(n13541) );
  XNOR U13482 ( .A(n13547), .B(n13845), .Z(n13540) );
  XNOR U13483 ( .A(n13548), .B(n13549), .Z(n13845) );
  AND U13484 ( .A(n13846), .B(n13847), .Z(n13549) );
  NAND U13485 ( .A(n13848), .B(n13849), .Z(n13847) );
  NANDN U13486 ( .A(n13850), .B(n13851), .Z(n13846) );
  OR U13487 ( .A(n13848), .B(n13849), .Z(n13851) );
  ANDN U13488 ( .B(\stack[0][40] ), .A(n5387), .Z(n13548) );
  XNOR U13489 ( .A(n13554), .B(n13852), .Z(n13547) );
  XNOR U13490 ( .A(n13555), .B(n13556), .Z(n13852) );
  AND U13491 ( .A(n13853), .B(n13854), .Z(n13556) );
  NANDN U13492 ( .A(n13855), .B(n13856), .Z(n13854) );
  NANDN U13493 ( .A(n13857), .B(n13858), .Z(n13853) );
  NANDN U13494 ( .A(n13856), .B(n13855), .Z(n13858) );
  ANDN U13495 ( .B(\stack[1][10] ), .A(n6094), .Z(n13555) );
  XNOR U13496 ( .A(n13561), .B(n13859), .Z(n13554) );
  XNOR U13497 ( .A(n13562), .B(n13563), .Z(n13859) );
  AND U13498 ( .A(n13860), .B(n13861), .Z(n13563) );
  NAND U13499 ( .A(n13862), .B(n13863), .Z(n13861) );
  NANDN U13500 ( .A(n13864), .B(n13865), .Z(n13860) );
  OR U13501 ( .A(n13862), .B(n13863), .Z(n13865) );
  ANDN U13502 ( .B(\stack[1][11] ), .A(n6070), .Z(n13562) );
  XNOR U13503 ( .A(n13568), .B(n13866), .Z(n13561) );
  XNOR U13504 ( .A(n13569), .B(n13570), .Z(n13866) );
  AND U13505 ( .A(n13867), .B(n13868), .Z(n13570) );
  NANDN U13506 ( .A(n13869), .B(n13870), .Z(n13868) );
  NANDN U13507 ( .A(n13871), .B(n13872), .Z(n13867) );
  NANDN U13508 ( .A(n13870), .B(n13869), .Z(n13872) );
  ANDN U13509 ( .B(\stack[1][12] ), .A(n6046), .Z(n13569) );
  XNOR U13510 ( .A(n13575), .B(n13873), .Z(n13568) );
  XNOR U13511 ( .A(n13576), .B(n13577), .Z(n13873) );
  AND U13512 ( .A(n13874), .B(n13875), .Z(n13577) );
  NAND U13513 ( .A(n13876), .B(n13877), .Z(n13875) );
  NANDN U13514 ( .A(n13878), .B(n13879), .Z(n13874) );
  OR U13515 ( .A(n13876), .B(n13877), .Z(n13879) );
  ANDN U13516 ( .B(\stack[1][13] ), .A(n6022), .Z(n13576) );
  XNOR U13517 ( .A(n13582), .B(n13880), .Z(n13575) );
  XNOR U13518 ( .A(n13583), .B(n13584), .Z(n13880) );
  AND U13519 ( .A(n13881), .B(n13882), .Z(n13584) );
  NANDN U13520 ( .A(n13883), .B(n13884), .Z(n13882) );
  NANDN U13521 ( .A(n13885), .B(n13886), .Z(n13881) );
  NANDN U13522 ( .A(n13884), .B(n13883), .Z(n13886) );
  ANDN U13523 ( .B(\stack[1][14] ), .A(n5998), .Z(n13583) );
  XNOR U13524 ( .A(n13589), .B(n13887), .Z(n13582) );
  XNOR U13525 ( .A(n13590), .B(n13591), .Z(n13887) );
  AND U13526 ( .A(n13888), .B(n13889), .Z(n13591) );
  NAND U13527 ( .A(n13890), .B(n13891), .Z(n13889) );
  NANDN U13528 ( .A(n13892), .B(n13893), .Z(n13888) );
  OR U13529 ( .A(n13890), .B(n13891), .Z(n13893) );
  ANDN U13530 ( .B(\stack[1][15] ), .A(n5974), .Z(n13590) );
  XNOR U13531 ( .A(n13596), .B(n13894), .Z(n13589) );
  XNOR U13532 ( .A(n13597), .B(n13598), .Z(n13894) );
  AND U13533 ( .A(n13895), .B(n13896), .Z(n13598) );
  NANDN U13534 ( .A(n13897), .B(n13898), .Z(n13896) );
  NANDN U13535 ( .A(n13899), .B(n13900), .Z(n13895) );
  NANDN U13536 ( .A(n13898), .B(n13897), .Z(n13900) );
  ANDN U13537 ( .B(\stack[1][16] ), .A(n5950), .Z(n13597) );
  XNOR U13538 ( .A(n13603), .B(n13901), .Z(n13596) );
  XNOR U13539 ( .A(n13604), .B(n13605), .Z(n13901) );
  AND U13540 ( .A(n13902), .B(n13903), .Z(n13605) );
  NAND U13541 ( .A(n13904), .B(n13905), .Z(n13903) );
  NANDN U13542 ( .A(n13906), .B(n13907), .Z(n13902) );
  OR U13543 ( .A(n13904), .B(n13905), .Z(n13907) );
  ANDN U13544 ( .B(\stack[1][17] ), .A(n5926), .Z(n13604) );
  XNOR U13545 ( .A(n13610), .B(n13908), .Z(n13603) );
  XNOR U13546 ( .A(n13611), .B(n13612), .Z(n13908) );
  AND U13547 ( .A(n13909), .B(n13910), .Z(n13612) );
  NANDN U13548 ( .A(n13911), .B(n13912), .Z(n13910) );
  NANDN U13549 ( .A(n13913), .B(n13914), .Z(n13909) );
  NANDN U13550 ( .A(n13912), .B(n13911), .Z(n13914) );
  ANDN U13551 ( .B(\stack[1][18] ), .A(n5902), .Z(n13611) );
  XNOR U13552 ( .A(n13617), .B(n13915), .Z(n13610) );
  XNOR U13553 ( .A(n13618), .B(n13619), .Z(n13915) );
  AND U13554 ( .A(n13916), .B(n13917), .Z(n13619) );
  NAND U13555 ( .A(n13918), .B(n13919), .Z(n13917) );
  NANDN U13556 ( .A(n13920), .B(n13921), .Z(n13916) );
  OR U13557 ( .A(n13918), .B(n13919), .Z(n13921) );
  ANDN U13558 ( .B(\stack[1][19] ), .A(n5878), .Z(n13618) );
  XNOR U13559 ( .A(n13624), .B(n13922), .Z(n13617) );
  XNOR U13560 ( .A(n13625), .B(n13626), .Z(n13922) );
  AND U13561 ( .A(n13923), .B(n13924), .Z(n13626) );
  NANDN U13562 ( .A(n13925), .B(n13926), .Z(n13924) );
  NANDN U13563 ( .A(n13927), .B(n13928), .Z(n13923) );
  NANDN U13564 ( .A(n13926), .B(n13925), .Z(n13928) );
  ANDN U13565 ( .B(\stack[1][20] ), .A(n5854), .Z(n13625) );
  XNOR U13566 ( .A(n13631), .B(n13929), .Z(n13624) );
  XNOR U13567 ( .A(n13632), .B(n13633), .Z(n13929) );
  AND U13568 ( .A(n13930), .B(n13931), .Z(n13633) );
  NAND U13569 ( .A(n13932), .B(n13933), .Z(n13931) );
  NANDN U13570 ( .A(n13934), .B(n13935), .Z(n13930) );
  OR U13571 ( .A(n13932), .B(n13933), .Z(n13935) );
  ANDN U13572 ( .B(\stack[1][21] ), .A(n5830), .Z(n13632) );
  XNOR U13573 ( .A(n13638), .B(n13936), .Z(n13631) );
  XNOR U13574 ( .A(n13639), .B(n13640), .Z(n13936) );
  AND U13575 ( .A(n13937), .B(n13938), .Z(n13640) );
  NANDN U13576 ( .A(n13939), .B(n13940), .Z(n13938) );
  NANDN U13577 ( .A(n13941), .B(n13942), .Z(n13937) );
  NANDN U13578 ( .A(n13940), .B(n13939), .Z(n13942) );
  ANDN U13579 ( .B(\stack[1][22] ), .A(n5806), .Z(n13639) );
  XNOR U13580 ( .A(n13645), .B(n13943), .Z(n13638) );
  XNOR U13581 ( .A(n13646), .B(n13647), .Z(n13943) );
  AND U13582 ( .A(n13944), .B(n13945), .Z(n13647) );
  NAND U13583 ( .A(n13946), .B(n13947), .Z(n13945) );
  NANDN U13584 ( .A(n13948), .B(n13949), .Z(n13944) );
  OR U13585 ( .A(n13946), .B(n13947), .Z(n13949) );
  ANDN U13586 ( .B(\stack[1][23] ), .A(n5782), .Z(n13646) );
  XNOR U13587 ( .A(n13652), .B(n13950), .Z(n13645) );
  XNOR U13588 ( .A(n13653), .B(n13654), .Z(n13950) );
  AND U13589 ( .A(n13951), .B(n13952), .Z(n13654) );
  NANDN U13590 ( .A(n13953), .B(n13954), .Z(n13952) );
  NANDN U13591 ( .A(n13955), .B(n13956), .Z(n13951) );
  NANDN U13592 ( .A(n13954), .B(n13953), .Z(n13956) );
  ANDN U13593 ( .B(\stack[1][24] ), .A(n5758), .Z(n13653) );
  XNOR U13594 ( .A(n13659), .B(n13957), .Z(n13652) );
  XNOR U13595 ( .A(n13660), .B(n13661), .Z(n13957) );
  AND U13596 ( .A(n13958), .B(n13959), .Z(n13661) );
  NAND U13597 ( .A(n13960), .B(n13961), .Z(n13959) );
  NANDN U13598 ( .A(n13962), .B(n13963), .Z(n13958) );
  OR U13599 ( .A(n13960), .B(n13961), .Z(n13963) );
  ANDN U13600 ( .B(\stack[1][25] ), .A(n5734), .Z(n13660) );
  XNOR U13601 ( .A(n13666), .B(n13964), .Z(n13659) );
  XNOR U13602 ( .A(n13667), .B(n13668), .Z(n13964) );
  AND U13603 ( .A(n13965), .B(n13966), .Z(n13668) );
  NANDN U13604 ( .A(n13967), .B(n13968), .Z(n13966) );
  NANDN U13605 ( .A(n13969), .B(n13970), .Z(n13965) );
  NANDN U13606 ( .A(n13968), .B(n13967), .Z(n13970) );
  ANDN U13607 ( .B(\stack[1][26] ), .A(n5710), .Z(n13667) );
  XNOR U13608 ( .A(n13673), .B(n13971), .Z(n13666) );
  XNOR U13609 ( .A(n13674), .B(n13675), .Z(n13971) );
  AND U13610 ( .A(n13972), .B(n13973), .Z(n13675) );
  NAND U13611 ( .A(n13974), .B(n13975), .Z(n13973) );
  NANDN U13612 ( .A(n13976), .B(n13977), .Z(n13972) );
  OR U13613 ( .A(n13974), .B(n13975), .Z(n13977) );
  ANDN U13614 ( .B(\stack[1][27] ), .A(n5686), .Z(n13674) );
  XNOR U13615 ( .A(n13680), .B(n13978), .Z(n13673) );
  XNOR U13616 ( .A(n13681), .B(n13682), .Z(n13978) );
  AND U13617 ( .A(n13979), .B(n13980), .Z(n13682) );
  NANDN U13618 ( .A(n13981), .B(n13982), .Z(n13980) );
  NANDN U13619 ( .A(n13983), .B(n13984), .Z(n13979) );
  NANDN U13620 ( .A(n13982), .B(n13981), .Z(n13984) );
  ANDN U13621 ( .B(\stack[1][28] ), .A(n5662), .Z(n13681) );
  XNOR U13622 ( .A(n13687), .B(n13985), .Z(n13680) );
  XNOR U13623 ( .A(n13688), .B(n13689), .Z(n13985) );
  AND U13624 ( .A(n13986), .B(n13987), .Z(n13689) );
  NAND U13625 ( .A(n13988), .B(n13989), .Z(n13987) );
  NANDN U13626 ( .A(n13990), .B(n13991), .Z(n13986) );
  OR U13627 ( .A(n13988), .B(n13989), .Z(n13991) );
  ANDN U13628 ( .B(\stack[1][29] ), .A(n5638), .Z(n13688) );
  XNOR U13629 ( .A(n13694), .B(n13992), .Z(n13687) );
  XNOR U13630 ( .A(n13695), .B(n13696), .Z(n13992) );
  AND U13631 ( .A(n13993), .B(n13994), .Z(n13696) );
  NANDN U13632 ( .A(n13995), .B(n13996), .Z(n13994) );
  NANDN U13633 ( .A(n13997), .B(n13998), .Z(n13993) );
  NANDN U13634 ( .A(n13996), .B(n13995), .Z(n13998) );
  ANDN U13635 ( .B(\stack[1][30] ), .A(n5614), .Z(n13695) );
  XNOR U13636 ( .A(n13701), .B(n13999), .Z(n13694) );
  XNOR U13637 ( .A(n13702), .B(n13703), .Z(n13999) );
  AND U13638 ( .A(n14000), .B(n14001), .Z(n13703) );
  NAND U13639 ( .A(n14002), .B(n14003), .Z(n14001) );
  NANDN U13640 ( .A(n14004), .B(n14005), .Z(n14000) );
  OR U13641 ( .A(n14002), .B(n14003), .Z(n14005) );
  ANDN U13642 ( .B(\stack[1][31] ), .A(n5590), .Z(n13702) );
  XNOR U13643 ( .A(n13708), .B(n14006), .Z(n13701) );
  XNOR U13644 ( .A(n13709), .B(n13710), .Z(n14006) );
  AND U13645 ( .A(n14007), .B(n14008), .Z(n13710) );
  NANDN U13646 ( .A(n14009), .B(n14010), .Z(n14008) );
  NANDN U13647 ( .A(n14011), .B(n14012), .Z(n14007) );
  NANDN U13648 ( .A(n14010), .B(n14009), .Z(n14012) );
  ANDN U13649 ( .B(\stack[1][32] ), .A(n5566), .Z(n13709) );
  XNOR U13650 ( .A(n13715), .B(n14013), .Z(n13708) );
  XNOR U13651 ( .A(n13716), .B(n13717), .Z(n14013) );
  AND U13652 ( .A(n14014), .B(n14015), .Z(n13717) );
  NAND U13653 ( .A(n14016), .B(n14017), .Z(n14015) );
  NANDN U13654 ( .A(n14018), .B(n14019), .Z(n14014) );
  OR U13655 ( .A(n14016), .B(n14017), .Z(n14019) );
  ANDN U13656 ( .B(\stack[1][33] ), .A(n5542), .Z(n13716) );
  XNOR U13657 ( .A(n13722), .B(n14020), .Z(n13715) );
  XNOR U13658 ( .A(n13723), .B(n13724), .Z(n14020) );
  AND U13659 ( .A(n14021), .B(n14022), .Z(n13724) );
  NANDN U13660 ( .A(n14023), .B(n14024), .Z(n14022) );
  NANDN U13661 ( .A(n14025), .B(n14026), .Z(n14021) );
  NANDN U13662 ( .A(n14024), .B(n14023), .Z(n14026) );
  ANDN U13663 ( .B(\stack[1][34] ), .A(n5518), .Z(n13723) );
  XNOR U13664 ( .A(n13729), .B(n14027), .Z(n13722) );
  XNOR U13665 ( .A(n13730), .B(n13731), .Z(n14027) );
  AND U13666 ( .A(n14028), .B(n14029), .Z(n13731) );
  NAND U13667 ( .A(n14030), .B(n14031), .Z(n14029) );
  NANDN U13668 ( .A(n14032), .B(n14033), .Z(n14028) );
  OR U13669 ( .A(n14030), .B(n14031), .Z(n14033) );
  ANDN U13670 ( .B(\stack[1][35] ), .A(n5494), .Z(n13730) );
  XNOR U13671 ( .A(n13736), .B(n14034), .Z(n13729) );
  XNOR U13672 ( .A(n13737), .B(n13738), .Z(n14034) );
  AND U13673 ( .A(n14035), .B(n14036), .Z(n13738) );
  NANDN U13674 ( .A(n14037), .B(n14038), .Z(n14036) );
  NANDN U13675 ( .A(n14039), .B(n14040), .Z(n14035) );
  NANDN U13676 ( .A(n14038), .B(n14037), .Z(n14040) );
  ANDN U13677 ( .B(\stack[1][36] ), .A(n5470), .Z(n13737) );
  XNOR U13678 ( .A(n13743), .B(n14041), .Z(n13736) );
  XOR U13679 ( .A(n13745), .B(n13746), .Z(n14041) );
  NAND U13680 ( .A(n14042), .B(n14043), .Z(n13746) );
  NAND U13681 ( .A(n14044), .B(n14045), .Z(n14043) );
  OR U13682 ( .A(n14046), .B(n14047), .Z(n14044) );
  AND U13683 ( .A(\stack[0][12] ), .B(\stack[1][37] ), .Z(n13745) );
  XNOR U13684 ( .A(n13752), .B(n14048), .Z(n13743) );
  XOR U13685 ( .A(n13753), .B(n13751), .Z(n14048) );
  AND U13686 ( .A(\stack[0][11] ), .B(\stack[1][38] ), .Z(n13751) );
  NAND U13687 ( .A(n14049), .B(n14050), .Z(n13753) );
  OR U13688 ( .A(n14051), .B(n14052), .Z(n14050) );
  NAND U13689 ( .A(n14053), .B(n14054), .Z(n14049) );
  NAND U13690 ( .A(n14052), .B(n14051), .Z(n14053) );
  XNOR U13691 ( .A(n13757), .B(n14055), .Z(n13752) );
  XNOR U13692 ( .A(n13758), .B(n13759), .Z(n14055) );
  AND U13693 ( .A(n14056), .B(n14057), .Z(n13759) );
  NAND U13694 ( .A(n14058), .B(n14059), .Z(n14057) );
  NANDN U13695 ( .A(n14060), .B(n14061), .Z(n14056) );
  OR U13696 ( .A(n14058), .B(n14059), .Z(n14061) );
  ANDN U13697 ( .B(\stack[1][39] ), .A(n5398), .Z(n13758) );
  XNOR U13698 ( .A(n13764), .B(n14062), .Z(n13757) );
  XNOR U13699 ( .A(n13765), .B(n13766), .Z(n14062) );
  AND U13700 ( .A(n14063), .B(n14064), .Z(n13766) );
  NANDN U13701 ( .A(n14065), .B(n14066), .Z(n14064) );
  NANDN U13702 ( .A(n14067), .B(n14068), .Z(n14063) );
  NANDN U13703 ( .A(n14066), .B(n14065), .Z(n14068) );
  ANDN U13704 ( .B(\stack[1][40] ), .A(n5374), .Z(n13765) );
  XNOR U13705 ( .A(n13771), .B(n14069), .Z(n13764) );
  XNOR U13706 ( .A(n13772), .B(n13773), .Z(n14069) );
  AND U13707 ( .A(n14070), .B(n14071), .Z(n13773) );
  NAND U13708 ( .A(n14072), .B(n14073), .Z(n14071) );
  NANDN U13709 ( .A(n14074), .B(n14075), .Z(n14070) );
  OR U13710 ( .A(n14072), .B(n14073), .Z(n14075) );
  ANDN U13711 ( .B(\stack[1][41] ), .A(n5350), .Z(n13772) );
  XNOR U13712 ( .A(n13778), .B(n14076), .Z(n13771) );
  XNOR U13713 ( .A(n13779), .B(n13780), .Z(n14076) );
  AND U13714 ( .A(n14077), .B(n14078), .Z(n13780) );
  NANDN U13715 ( .A(n14079), .B(n14080), .Z(n14078) );
  NANDN U13716 ( .A(n14081), .B(n14082), .Z(n14077) );
  NANDN U13717 ( .A(n14080), .B(n14079), .Z(n14082) );
  ANDN U13718 ( .B(\stack[1][42] ), .A(n5326), .Z(n13779) );
  XNOR U13719 ( .A(n13785), .B(n14083), .Z(n13778) );
  XNOR U13720 ( .A(n13786), .B(n13787), .Z(n14083) );
  AND U13721 ( .A(n14084), .B(n14085), .Z(n13787) );
  NAND U13722 ( .A(n14086), .B(n14087), .Z(n14085) );
  NANDN U13723 ( .A(n14088), .B(n14089), .Z(n14084) );
  OR U13724 ( .A(n14086), .B(n14087), .Z(n14089) );
  ANDN U13725 ( .B(\stack[1][43] ), .A(n5302), .Z(n13786) );
  XNOR U13726 ( .A(n13792), .B(n14090), .Z(n13785) );
  XNOR U13727 ( .A(n13793), .B(n13794), .Z(n14090) );
  AND U13728 ( .A(n14091), .B(n14092), .Z(n13794) );
  NANDN U13729 ( .A(n14093), .B(n14094), .Z(n14092) );
  NANDN U13730 ( .A(n14095), .B(n14096), .Z(n14091) );
  NANDN U13731 ( .A(n14094), .B(n14093), .Z(n14096) );
  ANDN U13732 ( .B(\stack[1][44] ), .A(n5278), .Z(n13793) );
  XNOR U13733 ( .A(n13799), .B(n14097), .Z(n13792) );
  XNOR U13734 ( .A(n13800), .B(n13801), .Z(n14097) );
  AND U13735 ( .A(n14098), .B(n14099), .Z(n13801) );
  NAND U13736 ( .A(n14100), .B(n14101), .Z(n14099) );
  NANDN U13737 ( .A(n14102), .B(n14103), .Z(n14098) );
  OR U13738 ( .A(n14100), .B(n14101), .Z(n14103) );
  ANDN U13739 ( .B(\stack[1][45] ), .A(n5254), .Z(n13800) );
  XNOR U13740 ( .A(n13806), .B(n14104), .Z(n13799) );
  XNOR U13741 ( .A(n13807), .B(n13808), .Z(n14104) );
  AND U13742 ( .A(n14105), .B(n14106), .Z(n13808) );
  NAND U13743 ( .A(n14107), .B(n14108), .Z(n14106) );
  NAND U13744 ( .A(n14109), .B(n14110), .Z(n14105) );
  OR U13745 ( .A(n14107), .B(n14108), .Z(n14109) );
  ANDN U13746 ( .B(\stack[1][46] ), .A(n5230), .Z(n13807) );
  XNOR U13747 ( .A(n13813), .B(n14111), .Z(n13806) );
  XNOR U13748 ( .A(n13814), .B(n13816), .Z(n14111) );
  ANDN U13749 ( .B(n14112), .A(n14113), .Z(n13816) );
  ANDN U13750 ( .B(\stack[0][0] ), .A(n6324), .Z(n14112) );
  ANDN U13751 ( .B(\stack[1][47] ), .A(n5206), .Z(n13814) );
  XOR U13752 ( .A(n13819), .B(n14114), .Z(n13813) );
  NANDN U13753 ( .A(n5160), .B(\stack[1][49] ), .Z(n14114) );
  NANDN U13754 ( .A(n6324), .B(\stack[0][1] ), .Z(n13819) );
  ANDN U13755 ( .B(\stack[1][5] ), .A(n6214), .Z(n9055) );
  AND U13756 ( .A(n14115), .B(n14116), .Z(n9056) );
  NANDN U13757 ( .A(n9060), .B(n9062), .Z(n14116) );
  NANDN U13758 ( .A(n9063), .B(n14117), .Z(n14115) );
  NANDN U13759 ( .A(n9062), .B(n9060), .Z(n14117) );
  XOR U13760 ( .A(n13827), .B(n14118), .Z(n9060) );
  XNOR U13761 ( .A(n13828), .B(n13829), .Z(n14118) );
  AND U13762 ( .A(n14119), .B(n14120), .Z(n13829) );
  NAND U13763 ( .A(n14121), .B(n14122), .Z(n14120) );
  NANDN U13764 ( .A(n14123), .B(n14124), .Z(n14119) );
  OR U13765 ( .A(n14121), .B(n14122), .Z(n14124) );
  ANDN U13766 ( .B(\stack[0][42] ), .A(n5316), .Z(n13828) );
  XNOR U13767 ( .A(n13834), .B(n14125), .Z(n13827) );
  XNOR U13768 ( .A(n13835), .B(n13836), .Z(n14125) );
  AND U13769 ( .A(n14126), .B(n14127), .Z(n13836) );
  NANDN U13770 ( .A(n14128), .B(n14129), .Z(n14127) );
  NANDN U13771 ( .A(n14130), .B(n14131), .Z(n14126) );
  NANDN U13772 ( .A(n14129), .B(n14128), .Z(n14131) );
  ANDN U13773 ( .B(\stack[0][41] ), .A(n5340), .Z(n13835) );
  XNOR U13774 ( .A(n13841), .B(n14132), .Z(n13834) );
  XNOR U13775 ( .A(n13842), .B(n13843), .Z(n14132) );
  AND U13776 ( .A(n14133), .B(n14134), .Z(n13843) );
  NAND U13777 ( .A(n14135), .B(n14136), .Z(n14134) );
  NANDN U13778 ( .A(n14137), .B(n14138), .Z(n14133) );
  OR U13779 ( .A(n14135), .B(n14136), .Z(n14138) );
  ANDN U13780 ( .B(\stack[0][40] ), .A(n5364), .Z(n13842) );
  XNOR U13781 ( .A(n13848), .B(n14139), .Z(n13841) );
  XNOR U13782 ( .A(n13849), .B(n13850), .Z(n14139) );
  AND U13783 ( .A(n14140), .B(n14141), .Z(n13850) );
  NANDN U13784 ( .A(n14142), .B(n14143), .Z(n14141) );
  NANDN U13785 ( .A(n14144), .B(n14145), .Z(n14140) );
  NANDN U13786 ( .A(n14143), .B(n14142), .Z(n14145) );
  ANDN U13787 ( .B(\stack[0][39] ), .A(n5387), .Z(n13849) );
  XNOR U13788 ( .A(n13855), .B(n14146), .Z(n13848) );
  XNOR U13789 ( .A(n13856), .B(n13857), .Z(n14146) );
  AND U13790 ( .A(n14147), .B(n14148), .Z(n13857) );
  NAND U13791 ( .A(n14149), .B(n14150), .Z(n14148) );
  NANDN U13792 ( .A(n14151), .B(n14152), .Z(n14147) );
  OR U13793 ( .A(n14149), .B(n14150), .Z(n14152) );
  ANDN U13794 ( .B(\stack[1][10] ), .A(n6070), .Z(n13856) );
  XNOR U13795 ( .A(n13862), .B(n14153), .Z(n13855) );
  XNOR U13796 ( .A(n13863), .B(n13864), .Z(n14153) );
  AND U13797 ( .A(n14154), .B(n14155), .Z(n13864) );
  NANDN U13798 ( .A(n14156), .B(n14157), .Z(n14155) );
  NANDN U13799 ( .A(n14158), .B(n14159), .Z(n14154) );
  NANDN U13800 ( .A(n14157), .B(n14156), .Z(n14159) );
  ANDN U13801 ( .B(\stack[1][11] ), .A(n6046), .Z(n13863) );
  XNOR U13802 ( .A(n13869), .B(n14160), .Z(n13862) );
  XNOR U13803 ( .A(n13870), .B(n13871), .Z(n14160) );
  AND U13804 ( .A(n14161), .B(n14162), .Z(n13871) );
  NAND U13805 ( .A(n14163), .B(n14164), .Z(n14162) );
  NANDN U13806 ( .A(n14165), .B(n14166), .Z(n14161) );
  OR U13807 ( .A(n14163), .B(n14164), .Z(n14166) );
  ANDN U13808 ( .B(\stack[1][12] ), .A(n6022), .Z(n13870) );
  XNOR U13809 ( .A(n13876), .B(n14167), .Z(n13869) );
  XNOR U13810 ( .A(n13877), .B(n13878), .Z(n14167) );
  AND U13811 ( .A(n14168), .B(n14169), .Z(n13878) );
  NANDN U13812 ( .A(n14170), .B(n14171), .Z(n14169) );
  NANDN U13813 ( .A(n14172), .B(n14173), .Z(n14168) );
  NANDN U13814 ( .A(n14171), .B(n14170), .Z(n14173) );
  ANDN U13815 ( .B(\stack[1][13] ), .A(n5998), .Z(n13877) );
  XNOR U13816 ( .A(n13883), .B(n14174), .Z(n13876) );
  XNOR U13817 ( .A(n13884), .B(n13885), .Z(n14174) );
  AND U13818 ( .A(n14175), .B(n14176), .Z(n13885) );
  NAND U13819 ( .A(n14177), .B(n14178), .Z(n14176) );
  NANDN U13820 ( .A(n14179), .B(n14180), .Z(n14175) );
  OR U13821 ( .A(n14177), .B(n14178), .Z(n14180) );
  ANDN U13822 ( .B(\stack[1][14] ), .A(n5974), .Z(n13884) );
  XNOR U13823 ( .A(n13890), .B(n14181), .Z(n13883) );
  XNOR U13824 ( .A(n13891), .B(n13892), .Z(n14181) );
  AND U13825 ( .A(n14182), .B(n14183), .Z(n13892) );
  NANDN U13826 ( .A(n14184), .B(n14185), .Z(n14183) );
  NANDN U13827 ( .A(n14186), .B(n14187), .Z(n14182) );
  NANDN U13828 ( .A(n14185), .B(n14184), .Z(n14187) );
  ANDN U13829 ( .B(\stack[1][15] ), .A(n5950), .Z(n13891) );
  XNOR U13830 ( .A(n13897), .B(n14188), .Z(n13890) );
  XNOR U13831 ( .A(n13898), .B(n13899), .Z(n14188) );
  AND U13832 ( .A(n14189), .B(n14190), .Z(n13899) );
  NAND U13833 ( .A(n14191), .B(n14192), .Z(n14190) );
  NANDN U13834 ( .A(n14193), .B(n14194), .Z(n14189) );
  OR U13835 ( .A(n14191), .B(n14192), .Z(n14194) );
  ANDN U13836 ( .B(\stack[1][16] ), .A(n5926), .Z(n13898) );
  XNOR U13837 ( .A(n13904), .B(n14195), .Z(n13897) );
  XNOR U13838 ( .A(n13905), .B(n13906), .Z(n14195) );
  AND U13839 ( .A(n14196), .B(n14197), .Z(n13906) );
  NANDN U13840 ( .A(n14198), .B(n14199), .Z(n14197) );
  NANDN U13841 ( .A(n14200), .B(n14201), .Z(n14196) );
  NANDN U13842 ( .A(n14199), .B(n14198), .Z(n14201) );
  ANDN U13843 ( .B(\stack[1][17] ), .A(n5902), .Z(n13905) );
  XNOR U13844 ( .A(n13911), .B(n14202), .Z(n13904) );
  XNOR U13845 ( .A(n13912), .B(n13913), .Z(n14202) );
  AND U13846 ( .A(n14203), .B(n14204), .Z(n13913) );
  NAND U13847 ( .A(n14205), .B(n14206), .Z(n14204) );
  NANDN U13848 ( .A(n14207), .B(n14208), .Z(n14203) );
  OR U13849 ( .A(n14205), .B(n14206), .Z(n14208) );
  ANDN U13850 ( .B(\stack[1][18] ), .A(n5878), .Z(n13912) );
  XNOR U13851 ( .A(n13918), .B(n14209), .Z(n13911) );
  XNOR U13852 ( .A(n13919), .B(n13920), .Z(n14209) );
  AND U13853 ( .A(n14210), .B(n14211), .Z(n13920) );
  NANDN U13854 ( .A(n14212), .B(n14213), .Z(n14211) );
  NANDN U13855 ( .A(n14214), .B(n14215), .Z(n14210) );
  NANDN U13856 ( .A(n14213), .B(n14212), .Z(n14215) );
  ANDN U13857 ( .B(\stack[1][19] ), .A(n5854), .Z(n13919) );
  XNOR U13858 ( .A(n13925), .B(n14216), .Z(n13918) );
  XNOR U13859 ( .A(n13926), .B(n13927), .Z(n14216) );
  AND U13860 ( .A(n14217), .B(n14218), .Z(n13927) );
  NAND U13861 ( .A(n14219), .B(n14220), .Z(n14218) );
  NANDN U13862 ( .A(n14221), .B(n14222), .Z(n14217) );
  OR U13863 ( .A(n14219), .B(n14220), .Z(n14222) );
  ANDN U13864 ( .B(\stack[1][20] ), .A(n5830), .Z(n13926) );
  XNOR U13865 ( .A(n13932), .B(n14223), .Z(n13925) );
  XNOR U13866 ( .A(n13933), .B(n13934), .Z(n14223) );
  AND U13867 ( .A(n14224), .B(n14225), .Z(n13934) );
  NANDN U13868 ( .A(n14226), .B(n14227), .Z(n14225) );
  NANDN U13869 ( .A(n14228), .B(n14229), .Z(n14224) );
  NANDN U13870 ( .A(n14227), .B(n14226), .Z(n14229) );
  ANDN U13871 ( .B(\stack[1][21] ), .A(n5806), .Z(n13933) );
  XNOR U13872 ( .A(n13939), .B(n14230), .Z(n13932) );
  XNOR U13873 ( .A(n13940), .B(n13941), .Z(n14230) );
  AND U13874 ( .A(n14231), .B(n14232), .Z(n13941) );
  NAND U13875 ( .A(n14233), .B(n14234), .Z(n14232) );
  NANDN U13876 ( .A(n14235), .B(n14236), .Z(n14231) );
  OR U13877 ( .A(n14233), .B(n14234), .Z(n14236) );
  ANDN U13878 ( .B(\stack[1][22] ), .A(n5782), .Z(n13940) );
  XNOR U13879 ( .A(n13946), .B(n14237), .Z(n13939) );
  XNOR U13880 ( .A(n13947), .B(n13948), .Z(n14237) );
  AND U13881 ( .A(n14238), .B(n14239), .Z(n13948) );
  NANDN U13882 ( .A(n14240), .B(n14241), .Z(n14239) );
  NANDN U13883 ( .A(n14242), .B(n14243), .Z(n14238) );
  NANDN U13884 ( .A(n14241), .B(n14240), .Z(n14243) );
  ANDN U13885 ( .B(\stack[1][23] ), .A(n5758), .Z(n13947) );
  XNOR U13886 ( .A(n13953), .B(n14244), .Z(n13946) );
  XNOR U13887 ( .A(n13954), .B(n13955), .Z(n14244) );
  AND U13888 ( .A(n14245), .B(n14246), .Z(n13955) );
  NAND U13889 ( .A(n14247), .B(n14248), .Z(n14246) );
  NANDN U13890 ( .A(n14249), .B(n14250), .Z(n14245) );
  OR U13891 ( .A(n14247), .B(n14248), .Z(n14250) );
  ANDN U13892 ( .B(\stack[1][24] ), .A(n5734), .Z(n13954) );
  XNOR U13893 ( .A(n13960), .B(n14251), .Z(n13953) );
  XNOR U13894 ( .A(n13961), .B(n13962), .Z(n14251) );
  AND U13895 ( .A(n14252), .B(n14253), .Z(n13962) );
  NANDN U13896 ( .A(n14254), .B(n14255), .Z(n14253) );
  NANDN U13897 ( .A(n14256), .B(n14257), .Z(n14252) );
  NANDN U13898 ( .A(n14255), .B(n14254), .Z(n14257) );
  ANDN U13899 ( .B(\stack[1][25] ), .A(n5710), .Z(n13961) );
  XNOR U13900 ( .A(n13967), .B(n14258), .Z(n13960) );
  XNOR U13901 ( .A(n13968), .B(n13969), .Z(n14258) );
  AND U13902 ( .A(n14259), .B(n14260), .Z(n13969) );
  NAND U13903 ( .A(n14261), .B(n14262), .Z(n14260) );
  NANDN U13904 ( .A(n14263), .B(n14264), .Z(n14259) );
  OR U13905 ( .A(n14261), .B(n14262), .Z(n14264) );
  ANDN U13906 ( .B(\stack[1][26] ), .A(n5686), .Z(n13968) );
  XNOR U13907 ( .A(n13974), .B(n14265), .Z(n13967) );
  XNOR U13908 ( .A(n13975), .B(n13976), .Z(n14265) );
  AND U13909 ( .A(n14266), .B(n14267), .Z(n13976) );
  NANDN U13910 ( .A(n14268), .B(n14269), .Z(n14267) );
  NANDN U13911 ( .A(n14270), .B(n14271), .Z(n14266) );
  NANDN U13912 ( .A(n14269), .B(n14268), .Z(n14271) );
  ANDN U13913 ( .B(\stack[1][27] ), .A(n5662), .Z(n13975) );
  XNOR U13914 ( .A(n13981), .B(n14272), .Z(n13974) );
  XNOR U13915 ( .A(n13982), .B(n13983), .Z(n14272) );
  AND U13916 ( .A(n14273), .B(n14274), .Z(n13983) );
  NAND U13917 ( .A(n14275), .B(n14276), .Z(n14274) );
  NANDN U13918 ( .A(n14277), .B(n14278), .Z(n14273) );
  OR U13919 ( .A(n14275), .B(n14276), .Z(n14278) );
  ANDN U13920 ( .B(\stack[1][28] ), .A(n5638), .Z(n13982) );
  XNOR U13921 ( .A(n13988), .B(n14279), .Z(n13981) );
  XNOR U13922 ( .A(n13989), .B(n13990), .Z(n14279) );
  AND U13923 ( .A(n14280), .B(n14281), .Z(n13990) );
  NANDN U13924 ( .A(n14282), .B(n14283), .Z(n14281) );
  NANDN U13925 ( .A(n14284), .B(n14285), .Z(n14280) );
  NANDN U13926 ( .A(n14283), .B(n14282), .Z(n14285) );
  ANDN U13927 ( .B(\stack[1][29] ), .A(n5614), .Z(n13989) );
  XNOR U13928 ( .A(n13995), .B(n14286), .Z(n13988) );
  XNOR U13929 ( .A(n13996), .B(n13997), .Z(n14286) );
  AND U13930 ( .A(n14287), .B(n14288), .Z(n13997) );
  NAND U13931 ( .A(n14289), .B(n14290), .Z(n14288) );
  NANDN U13932 ( .A(n14291), .B(n14292), .Z(n14287) );
  OR U13933 ( .A(n14289), .B(n14290), .Z(n14292) );
  ANDN U13934 ( .B(\stack[1][30] ), .A(n5590), .Z(n13996) );
  XNOR U13935 ( .A(n14002), .B(n14293), .Z(n13995) );
  XNOR U13936 ( .A(n14003), .B(n14004), .Z(n14293) );
  AND U13937 ( .A(n14294), .B(n14295), .Z(n14004) );
  NANDN U13938 ( .A(n14296), .B(n14297), .Z(n14295) );
  NANDN U13939 ( .A(n14298), .B(n14299), .Z(n14294) );
  NANDN U13940 ( .A(n14297), .B(n14296), .Z(n14299) );
  ANDN U13941 ( .B(\stack[1][31] ), .A(n5566), .Z(n14003) );
  XNOR U13942 ( .A(n14009), .B(n14300), .Z(n14002) );
  XNOR U13943 ( .A(n14010), .B(n14011), .Z(n14300) );
  AND U13944 ( .A(n14301), .B(n14302), .Z(n14011) );
  NAND U13945 ( .A(n14303), .B(n14304), .Z(n14302) );
  NANDN U13946 ( .A(n14305), .B(n14306), .Z(n14301) );
  OR U13947 ( .A(n14303), .B(n14304), .Z(n14306) );
  ANDN U13948 ( .B(\stack[1][32] ), .A(n5542), .Z(n14010) );
  XNOR U13949 ( .A(n14016), .B(n14307), .Z(n14009) );
  XNOR U13950 ( .A(n14017), .B(n14018), .Z(n14307) );
  AND U13951 ( .A(n14308), .B(n14309), .Z(n14018) );
  NANDN U13952 ( .A(n14310), .B(n14311), .Z(n14309) );
  NANDN U13953 ( .A(n14312), .B(n14313), .Z(n14308) );
  NANDN U13954 ( .A(n14311), .B(n14310), .Z(n14313) );
  ANDN U13955 ( .B(\stack[1][33] ), .A(n5518), .Z(n14017) );
  XNOR U13956 ( .A(n14023), .B(n14314), .Z(n14016) );
  XNOR U13957 ( .A(n14024), .B(n14025), .Z(n14314) );
  AND U13958 ( .A(n14315), .B(n14316), .Z(n14025) );
  NAND U13959 ( .A(n14317), .B(n14318), .Z(n14316) );
  NANDN U13960 ( .A(n14319), .B(n14320), .Z(n14315) );
  OR U13961 ( .A(n14317), .B(n14318), .Z(n14320) );
  ANDN U13962 ( .B(\stack[1][34] ), .A(n5494), .Z(n14024) );
  XNOR U13963 ( .A(n14030), .B(n14321), .Z(n14023) );
  XNOR U13964 ( .A(n14031), .B(n14032), .Z(n14321) );
  AND U13965 ( .A(n14322), .B(n14323), .Z(n14032) );
  NANDN U13966 ( .A(n14324), .B(n14325), .Z(n14323) );
  NANDN U13967 ( .A(n14326), .B(n14327), .Z(n14322) );
  NANDN U13968 ( .A(n14325), .B(n14324), .Z(n14327) );
  ANDN U13969 ( .B(\stack[1][35] ), .A(n5470), .Z(n14031) );
  XNOR U13970 ( .A(n14037), .B(n14328), .Z(n14030) );
  XNOR U13971 ( .A(n14038), .B(n14039), .Z(n14328) );
  AND U13972 ( .A(n14329), .B(n14330), .Z(n14039) );
  NAND U13973 ( .A(n14331), .B(n14332), .Z(n14330) );
  NANDN U13974 ( .A(n14333), .B(n14334), .Z(n14329) );
  OR U13975 ( .A(n14331), .B(n14332), .Z(n14334) );
  ANDN U13976 ( .B(\stack[1][36] ), .A(n5446), .Z(n14038) );
  XNOR U13977 ( .A(n14045), .B(n14335), .Z(n14037) );
  XOR U13978 ( .A(n14046), .B(n14047), .Z(n14335) );
  NAND U13979 ( .A(n14336), .B(n14337), .Z(n14047) );
  NANDN U13980 ( .A(n14338), .B(n14339), .Z(n14337) );
  OR U13981 ( .A(n14340), .B(n14341), .Z(n14339) );
  AND U13982 ( .A(\stack[0][11] ), .B(\stack[1][37] ), .Z(n14046) );
  XNOR U13983 ( .A(n14052), .B(n14342), .Z(n14045) );
  XNOR U13984 ( .A(n14051), .B(n14054), .Z(n14342) );
  AND U13985 ( .A(\stack[0][10] ), .B(\stack[1][38] ), .Z(n14054) );
  AND U13986 ( .A(n14343), .B(n14344), .Z(n14051) );
  NAND U13987 ( .A(n14345), .B(n14346), .Z(n14344) );
  OR U13988 ( .A(n14347), .B(n14348), .Z(n14345) );
  XNOR U13989 ( .A(n14058), .B(n14349), .Z(n14052) );
  XNOR U13990 ( .A(n14059), .B(n14060), .Z(n14349) );
  AND U13991 ( .A(n14350), .B(n14351), .Z(n14060) );
  NANDN U13992 ( .A(n14352), .B(n14353), .Z(n14351) );
  NANDN U13993 ( .A(n14354), .B(n14355), .Z(n14350) );
  NANDN U13994 ( .A(n14353), .B(n14352), .Z(n14355) );
  ANDN U13995 ( .B(\stack[1][39] ), .A(n5374), .Z(n14059) );
  XNOR U13996 ( .A(n14065), .B(n14356), .Z(n14058) );
  XNOR U13997 ( .A(n14066), .B(n14067), .Z(n14356) );
  AND U13998 ( .A(n14357), .B(n14358), .Z(n14067) );
  NAND U13999 ( .A(n14359), .B(n14360), .Z(n14358) );
  NANDN U14000 ( .A(n14361), .B(n14362), .Z(n14357) );
  OR U14001 ( .A(n14359), .B(n14360), .Z(n14362) );
  ANDN U14002 ( .B(\stack[1][40] ), .A(n5350), .Z(n14066) );
  XNOR U14003 ( .A(n14072), .B(n14363), .Z(n14065) );
  XNOR U14004 ( .A(n14073), .B(n14074), .Z(n14363) );
  AND U14005 ( .A(n14364), .B(n14365), .Z(n14074) );
  NANDN U14006 ( .A(n14366), .B(n14367), .Z(n14365) );
  NANDN U14007 ( .A(n14368), .B(n14369), .Z(n14364) );
  NANDN U14008 ( .A(n14367), .B(n14366), .Z(n14369) );
  ANDN U14009 ( .B(\stack[1][41] ), .A(n5326), .Z(n14073) );
  XNOR U14010 ( .A(n14079), .B(n14370), .Z(n14072) );
  XNOR U14011 ( .A(n14080), .B(n14081), .Z(n14370) );
  AND U14012 ( .A(n14371), .B(n14372), .Z(n14081) );
  NAND U14013 ( .A(n14373), .B(n14374), .Z(n14372) );
  NANDN U14014 ( .A(n14375), .B(n14376), .Z(n14371) );
  OR U14015 ( .A(n14373), .B(n14374), .Z(n14376) );
  ANDN U14016 ( .B(\stack[1][42] ), .A(n5302), .Z(n14080) );
  XNOR U14017 ( .A(n14086), .B(n14377), .Z(n14079) );
  XNOR U14018 ( .A(n14087), .B(n14088), .Z(n14377) );
  AND U14019 ( .A(n14378), .B(n14379), .Z(n14088) );
  NANDN U14020 ( .A(n14380), .B(n14381), .Z(n14379) );
  NANDN U14021 ( .A(n14382), .B(n14383), .Z(n14378) );
  NANDN U14022 ( .A(n14381), .B(n14380), .Z(n14383) );
  ANDN U14023 ( .B(\stack[1][43] ), .A(n5278), .Z(n14087) );
  XNOR U14024 ( .A(n14093), .B(n14384), .Z(n14086) );
  XNOR U14025 ( .A(n14094), .B(n14095), .Z(n14384) );
  AND U14026 ( .A(n14385), .B(n14386), .Z(n14095) );
  NAND U14027 ( .A(n14387), .B(n14388), .Z(n14386) );
  NANDN U14028 ( .A(n14389), .B(n14390), .Z(n14385) );
  OR U14029 ( .A(n14387), .B(n14388), .Z(n14390) );
  ANDN U14030 ( .B(\stack[1][44] ), .A(n5254), .Z(n14094) );
  XNOR U14031 ( .A(n14100), .B(n14391), .Z(n14093) );
  XNOR U14032 ( .A(n14101), .B(n14102), .Z(n14391) );
  AND U14033 ( .A(n14392), .B(n14393), .Z(n14102) );
  NAND U14034 ( .A(n14394), .B(n14395), .Z(n14393) );
  NAND U14035 ( .A(n14396), .B(n14397), .Z(n14392) );
  OR U14036 ( .A(n14394), .B(n14395), .Z(n14396) );
  ANDN U14037 ( .B(\stack[1][45] ), .A(n5230), .Z(n14101) );
  XNOR U14038 ( .A(n14107), .B(n14398), .Z(n14100) );
  XNOR U14039 ( .A(n14108), .B(n14110), .Z(n14398) );
  ANDN U14040 ( .B(n14399), .A(n14400), .Z(n14110) );
  ANDN U14041 ( .B(\stack[0][0] ), .A(n6300), .Z(n14399) );
  ANDN U14042 ( .B(\stack[1][46] ), .A(n5206), .Z(n14108) );
  XOR U14043 ( .A(n14113), .B(n14401), .Z(n14107) );
  NANDN U14044 ( .A(n5160), .B(\stack[1][48] ), .Z(n14401) );
  NANDN U14045 ( .A(n6300), .B(\stack[0][1] ), .Z(n14113) );
  ANDN U14046 ( .B(\stack[0][43] ), .A(n5292), .Z(n9062) );
  AND U14047 ( .A(n14402), .B(n14403), .Z(n9063) );
  NANDN U14048 ( .A(n9070), .B(n14404), .Z(n14402) );
  NANDN U14049 ( .A(n9069), .B(n9067), .Z(n14404) );
  XNOR U14050 ( .A(n14121), .B(n14405), .Z(n9067) );
  XNOR U14051 ( .A(n14122), .B(n14123), .Z(n14405) );
  AND U14052 ( .A(n14406), .B(n14407), .Z(n14123) );
  NANDN U14053 ( .A(n14408), .B(n14409), .Z(n14407) );
  NANDN U14054 ( .A(n14410), .B(n14411), .Z(n14406) );
  NANDN U14055 ( .A(n14409), .B(n14408), .Z(n14411) );
  ANDN U14056 ( .B(\stack[0][41] ), .A(n5316), .Z(n14122) );
  XNOR U14057 ( .A(n14128), .B(n14412), .Z(n14121) );
  XNOR U14058 ( .A(n14129), .B(n14130), .Z(n14412) );
  AND U14059 ( .A(n14413), .B(n14414), .Z(n14130) );
  NAND U14060 ( .A(n14415), .B(n14416), .Z(n14414) );
  NANDN U14061 ( .A(n14417), .B(n14418), .Z(n14413) );
  OR U14062 ( .A(n14415), .B(n14416), .Z(n14418) );
  ANDN U14063 ( .B(\stack[0][40] ), .A(n5340), .Z(n14129) );
  XNOR U14064 ( .A(n14135), .B(n14419), .Z(n14128) );
  XNOR U14065 ( .A(n14136), .B(n14137), .Z(n14419) );
  AND U14066 ( .A(n14420), .B(n14421), .Z(n14137) );
  NANDN U14067 ( .A(n14422), .B(n14423), .Z(n14421) );
  NANDN U14068 ( .A(n14424), .B(n14425), .Z(n14420) );
  NANDN U14069 ( .A(n14423), .B(n14422), .Z(n14425) );
  ANDN U14070 ( .B(\stack[0][39] ), .A(n5364), .Z(n14136) );
  XNOR U14071 ( .A(n14142), .B(n14426), .Z(n14135) );
  XNOR U14072 ( .A(n14143), .B(n14144), .Z(n14426) );
  AND U14073 ( .A(n14427), .B(n14428), .Z(n14144) );
  NAND U14074 ( .A(n14429), .B(n14430), .Z(n14428) );
  NANDN U14075 ( .A(n14431), .B(n14432), .Z(n14427) );
  OR U14076 ( .A(n14429), .B(n14430), .Z(n14432) );
  ANDN U14077 ( .B(\stack[0][38] ), .A(n5387), .Z(n14143) );
  XNOR U14078 ( .A(n14149), .B(n14433), .Z(n14142) );
  XNOR U14079 ( .A(n14150), .B(n14151), .Z(n14433) );
  AND U14080 ( .A(n14434), .B(n14435), .Z(n14151) );
  NANDN U14081 ( .A(n14436), .B(n14437), .Z(n14435) );
  NANDN U14082 ( .A(n14438), .B(n14439), .Z(n14434) );
  NANDN U14083 ( .A(n14437), .B(n14436), .Z(n14439) );
  ANDN U14084 ( .B(\stack[1][10] ), .A(n6046), .Z(n14150) );
  XNOR U14085 ( .A(n14156), .B(n14440), .Z(n14149) );
  XNOR U14086 ( .A(n14157), .B(n14158), .Z(n14440) );
  AND U14087 ( .A(n14441), .B(n14442), .Z(n14158) );
  NAND U14088 ( .A(n14443), .B(n14444), .Z(n14442) );
  NANDN U14089 ( .A(n14445), .B(n14446), .Z(n14441) );
  OR U14090 ( .A(n14443), .B(n14444), .Z(n14446) );
  ANDN U14091 ( .B(\stack[1][11] ), .A(n6022), .Z(n14157) );
  XNOR U14092 ( .A(n14163), .B(n14447), .Z(n14156) );
  XNOR U14093 ( .A(n14164), .B(n14165), .Z(n14447) );
  AND U14094 ( .A(n14448), .B(n14449), .Z(n14165) );
  NANDN U14095 ( .A(n14450), .B(n14451), .Z(n14449) );
  NANDN U14096 ( .A(n14452), .B(n14453), .Z(n14448) );
  NANDN U14097 ( .A(n14451), .B(n14450), .Z(n14453) );
  ANDN U14098 ( .B(\stack[1][12] ), .A(n5998), .Z(n14164) );
  XNOR U14099 ( .A(n14170), .B(n14454), .Z(n14163) );
  XNOR U14100 ( .A(n14171), .B(n14172), .Z(n14454) );
  AND U14101 ( .A(n14455), .B(n14456), .Z(n14172) );
  NAND U14102 ( .A(n14457), .B(n14458), .Z(n14456) );
  NANDN U14103 ( .A(n14459), .B(n14460), .Z(n14455) );
  OR U14104 ( .A(n14457), .B(n14458), .Z(n14460) );
  ANDN U14105 ( .B(\stack[1][13] ), .A(n5974), .Z(n14171) );
  XNOR U14106 ( .A(n14177), .B(n14461), .Z(n14170) );
  XNOR U14107 ( .A(n14178), .B(n14179), .Z(n14461) );
  AND U14108 ( .A(n14462), .B(n14463), .Z(n14179) );
  NANDN U14109 ( .A(n14464), .B(n14465), .Z(n14463) );
  NANDN U14110 ( .A(n14466), .B(n14467), .Z(n14462) );
  NANDN U14111 ( .A(n14465), .B(n14464), .Z(n14467) );
  ANDN U14112 ( .B(\stack[1][14] ), .A(n5950), .Z(n14178) );
  XNOR U14113 ( .A(n14184), .B(n14468), .Z(n14177) );
  XNOR U14114 ( .A(n14185), .B(n14186), .Z(n14468) );
  AND U14115 ( .A(n14469), .B(n14470), .Z(n14186) );
  NAND U14116 ( .A(n14471), .B(n14472), .Z(n14470) );
  NANDN U14117 ( .A(n14473), .B(n14474), .Z(n14469) );
  OR U14118 ( .A(n14471), .B(n14472), .Z(n14474) );
  ANDN U14119 ( .B(\stack[1][15] ), .A(n5926), .Z(n14185) );
  XNOR U14120 ( .A(n14191), .B(n14475), .Z(n14184) );
  XNOR U14121 ( .A(n14192), .B(n14193), .Z(n14475) );
  AND U14122 ( .A(n14476), .B(n14477), .Z(n14193) );
  NANDN U14123 ( .A(n14478), .B(n14479), .Z(n14477) );
  NANDN U14124 ( .A(n14480), .B(n14481), .Z(n14476) );
  NANDN U14125 ( .A(n14479), .B(n14478), .Z(n14481) );
  ANDN U14126 ( .B(\stack[1][16] ), .A(n5902), .Z(n14192) );
  XNOR U14127 ( .A(n14198), .B(n14482), .Z(n14191) );
  XNOR U14128 ( .A(n14199), .B(n14200), .Z(n14482) );
  AND U14129 ( .A(n14483), .B(n14484), .Z(n14200) );
  NAND U14130 ( .A(n14485), .B(n14486), .Z(n14484) );
  NANDN U14131 ( .A(n14487), .B(n14488), .Z(n14483) );
  OR U14132 ( .A(n14485), .B(n14486), .Z(n14488) );
  ANDN U14133 ( .B(\stack[1][17] ), .A(n5878), .Z(n14199) );
  XNOR U14134 ( .A(n14205), .B(n14489), .Z(n14198) );
  XNOR U14135 ( .A(n14206), .B(n14207), .Z(n14489) );
  AND U14136 ( .A(n14490), .B(n14491), .Z(n14207) );
  NANDN U14137 ( .A(n14492), .B(n14493), .Z(n14491) );
  NANDN U14138 ( .A(n14494), .B(n14495), .Z(n14490) );
  NANDN U14139 ( .A(n14493), .B(n14492), .Z(n14495) );
  ANDN U14140 ( .B(\stack[1][18] ), .A(n5854), .Z(n14206) );
  XNOR U14141 ( .A(n14212), .B(n14496), .Z(n14205) );
  XNOR U14142 ( .A(n14213), .B(n14214), .Z(n14496) );
  AND U14143 ( .A(n14497), .B(n14498), .Z(n14214) );
  NAND U14144 ( .A(n14499), .B(n14500), .Z(n14498) );
  NANDN U14145 ( .A(n14501), .B(n14502), .Z(n14497) );
  OR U14146 ( .A(n14499), .B(n14500), .Z(n14502) );
  ANDN U14147 ( .B(\stack[1][19] ), .A(n5830), .Z(n14213) );
  XNOR U14148 ( .A(n14219), .B(n14503), .Z(n14212) );
  XNOR U14149 ( .A(n14220), .B(n14221), .Z(n14503) );
  AND U14150 ( .A(n14504), .B(n14505), .Z(n14221) );
  NANDN U14151 ( .A(n14506), .B(n14507), .Z(n14505) );
  NANDN U14152 ( .A(n14508), .B(n14509), .Z(n14504) );
  NANDN U14153 ( .A(n14507), .B(n14506), .Z(n14509) );
  ANDN U14154 ( .B(\stack[1][20] ), .A(n5806), .Z(n14220) );
  XNOR U14155 ( .A(n14226), .B(n14510), .Z(n14219) );
  XNOR U14156 ( .A(n14227), .B(n14228), .Z(n14510) );
  AND U14157 ( .A(n14511), .B(n14512), .Z(n14228) );
  NAND U14158 ( .A(n14513), .B(n14514), .Z(n14512) );
  NANDN U14159 ( .A(n14515), .B(n14516), .Z(n14511) );
  OR U14160 ( .A(n14513), .B(n14514), .Z(n14516) );
  ANDN U14161 ( .B(\stack[1][21] ), .A(n5782), .Z(n14227) );
  XNOR U14162 ( .A(n14233), .B(n14517), .Z(n14226) );
  XNOR U14163 ( .A(n14234), .B(n14235), .Z(n14517) );
  AND U14164 ( .A(n14518), .B(n14519), .Z(n14235) );
  NANDN U14165 ( .A(n14520), .B(n14521), .Z(n14519) );
  NANDN U14166 ( .A(n14522), .B(n14523), .Z(n14518) );
  NANDN U14167 ( .A(n14521), .B(n14520), .Z(n14523) );
  ANDN U14168 ( .B(\stack[1][22] ), .A(n5758), .Z(n14234) );
  XNOR U14169 ( .A(n14240), .B(n14524), .Z(n14233) );
  XNOR U14170 ( .A(n14241), .B(n14242), .Z(n14524) );
  AND U14171 ( .A(n14525), .B(n14526), .Z(n14242) );
  NAND U14172 ( .A(n14527), .B(n14528), .Z(n14526) );
  NANDN U14173 ( .A(n14529), .B(n14530), .Z(n14525) );
  OR U14174 ( .A(n14527), .B(n14528), .Z(n14530) );
  ANDN U14175 ( .B(\stack[1][23] ), .A(n5734), .Z(n14241) );
  XNOR U14176 ( .A(n14247), .B(n14531), .Z(n14240) );
  XNOR U14177 ( .A(n14248), .B(n14249), .Z(n14531) );
  AND U14178 ( .A(n14532), .B(n14533), .Z(n14249) );
  NANDN U14179 ( .A(n14534), .B(n14535), .Z(n14533) );
  NANDN U14180 ( .A(n14536), .B(n14537), .Z(n14532) );
  NANDN U14181 ( .A(n14535), .B(n14534), .Z(n14537) );
  ANDN U14182 ( .B(\stack[1][24] ), .A(n5710), .Z(n14248) );
  XNOR U14183 ( .A(n14254), .B(n14538), .Z(n14247) );
  XNOR U14184 ( .A(n14255), .B(n14256), .Z(n14538) );
  AND U14185 ( .A(n14539), .B(n14540), .Z(n14256) );
  NAND U14186 ( .A(n14541), .B(n14542), .Z(n14540) );
  NANDN U14187 ( .A(n14543), .B(n14544), .Z(n14539) );
  OR U14188 ( .A(n14541), .B(n14542), .Z(n14544) );
  ANDN U14189 ( .B(\stack[1][25] ), .A(n5686), .Z(n14255) );
  XNOR U14190 ( .A(n14261), .B(n14545), .Z(n14254) );
  XNOR U14191 ( .A(n14262), .B(n14263), .Z(n14545) );
  AND U14192 ( .A(n14546), .B(n14547), .Z(n14263) );
  NANDN U14193 ( .A(n14548), .B(n14549), .Z(n14547) );
  NANDN U14194 ( .A(n14550), .B(n14551), .Z(n14546) );
  NANDN U14195 ( .A(n14549), .B(n14548), .Z(n14551) );
  ANDN U14196 ( .B(\stack[1][26] ), .A(n5662), .Z(n14262) );
  XNOR U14197 ( .A(n14268), .B(n14552), .Z(n14261) );
  XNOR U14198 ( .A(n14269), .B(n14270), .Z(n14552) );
  AND U14199 ( .A(n14553), .B(n14554), .Z(n14270) );
  NAND U14200 ( .A(n14555), .B(n14556), .Z(n14554) );
  NANDN U14201 ( .A(n14557), .B(n14558), .Z(n14553) );
  OR U14202 ( .A(n14555), .B(n14556), .Z(n14558) );
  ANDN U14203 ( .B(\stack[1][27] ), .A(n5638), .Z(n14269) );
  XNOR U14204 ( .A(n14275), .B(n14559), .Z(n14268) );
  XNOR U14205 ( .A(n14276), .B(n14277), .Z(n14559) );
  AND U14206 ( .A(n14560), .B(n14561), .Z(n14277) );
  NANDN U14207 ( .A(n14562), .B(n14563), .Z(n14561) );
  NANDN U14208 ( .A(n14564), .B(n14565), .Z(n14560) );
  NANDN U14209 ( .A(n14563), .B(n14562), .Z(n14565) );
  ANDN U14210 ( .B(\stack[1][28] ), .A(n5614), .Z(n14276) );
  XNOR U14211 ( .A(n14282), .B(n14566), .Z(n14275) );
  XNOR U14212 ( .A(n14283), .B(n14284), .Z(n14566) );
  AND U14213 ( .A(n14567), .B(n14568), .Z(n14284) );
  NAND U14214 ( .A(n14569), .B(n14570), .Z(n14568) );
  NANDN U14215 ( .A(n14571), .B(n14572), .Z(n14567) );
  OR U14216 ( .A(n14569), .B(n14570), .Z(n14572) );
  ANDN U14217 ( .B(\stack[1][29] ), .A(n5590), .Z(n14283) );
  XNOR U14218 ( .A(n14289), .B(n14573), .Z(n14282) );
  XNOR U14219 ( .A(n14290), .B(n14291), .Z(n14573) );
  AND U14220 ( .A(n14574), .B(n14575), .Z(n14291) );
  NANDN U14221 ( .A(n14576), .B(n14577), .Z(n14575) );
  NANDN U14222 ( .A(n14578), .B(n14579), .Z(n14574) );
  NANDN U14223 ( .A(n14577), .B(n14576), .Z(n14579) );
  ANDN U14224 ( .B(\stack[1][30] ), .A(n5566), .Z(n14290) );
  XNOR U14225 ( .A(n14296), .B(n14580), .Z(n14289) );
  XNOR U14226 ( .A(n14297), .B(n14298), .Z(n14580) );
  AND U14227 ( .A(n14581), .B(n14582), .Z(n14298) );
  NAND U14228 ( .A(n14583), .B(n14584), .Z(n14582) );
  NANDN U14229 ( .A(n14585), .B(n14586), .Z(n14581) );
  OR U14230 ( .A(n14583), .B(n14584), .Z(n14586) );
  ANDN U14231 ( .B(\stack[1][31] ), .A(n5542), .Z(n14297) );
  XNOR U14232 ( .A(n14303), .B(n14587), .Z(n14296) );
  XNOR U14233 ( .A(n14304), .B(n14305), .Z(n14587) );
  AND U14234 ( .A(n14588), .B(n14589), .Z(n14305) );
  NANDN U14235 ( .A(n14590), .B(n14591), .Z(n14589) );
  NANDN U14236 ( .A(n14592), .B(n14593), .Z(n14588) );
  NANDN U14237 ( .A(n14591), .B(n14590), .Z(n14593) );
  ANDN U14238 ( .B(\stack[1][32] ), .A(n5518), .Z(n14304) );
  XNOR U14239 ( .A(n14310), .B(n14594), .Z(n14303) );
  XNOR U14240 ( .A(n14311), .B(n14312), .Z(n14594) );
  AND U14241 ( .A(n14595), .B(n14596), .Z(n14312) );
  NAND U14242 ( .A(n14597), .B(n14598), .Z(n14596) );
  NANDN U14243 ( .A(n14599), .B(n14600), .Z(n14595) );
  OR U14244 ( .A(n14597), .B(n14598), .Z(n14600) );
  ANDN U14245 ( .B(\stack[1][33] ), .A(n5494), .Z(n14311) );
  XNOR U14246 ( .A(n14317), .B(n14601), .Z(n14310) );
  XNOR U14247 ( .A(n14318), .B(n14319), .Z(n14601) );
  AND U14248 ( .A(n14602), .B(n14603), .Z(n14319) );
  NANDN U14249 ( .A(n14604), .B(n14605), .Z(n14603) );
  NANDN U14250 ( .A(n14606), .B(n14607), .Z(n14602) );
  NANDN U14251 ( .A(n14605), .B(n14604), .Z(n14607) );
  ANDN U14252 ( .B(\stack[1][34] ), .A(n5470), .Z(n14318) );
  XNOR U14253 ( .A(n14324), .B(n14608), .Z(n14317) );
  XNOR U14254 ( .A(n14325), .B(n14326), .Z(n14608) );
  AND U14255 ( .A(n14609), .B(n14610), .Z(n14326) );
  NAND U14256 ( .A(n14611), .B(n14612), .Z(n14610) );
  NANDN U14257 ( .A(n14613), .B(n14614), .Z(n14609) );
  OR U14258 ( .A(n14611), .B(n14612), .Z(n14614) );
  ANDN U14259 ( .B(\stack[1][35] ), .A(n5446), .Z(n14325) );
  XNOR U14260 ( .A(n14331), .B(n14615), .Z(n14324) );
  XNOR U14261 ( .A(n14332), .B(n14333), .Z(n14615) );
  AND U14262 ( .A(n14616), .B(n14617), .Z(n14333) );
  NANDN U14263 ( .A(n14618), .B(n14619), .Z(n14617) );
  NANDN U14264 ( .A(n14620), .B(n14621), .Z(n14616) );
  NANDN U14265 ( .A(n14619), .B(n14618), .Z(n14621) );
  ANDN U14266 ( .B(\stack[1][36] ), .A(n5422), .Z(n14332) );
  XNOR U14267 ( .A(n14338), .B(n14622), .Z(n14331) );
  XOR U14268 ( .A(n14340), .B(n14341), .Z(n14622) );
  NAND U14269 ( .A(n14623), .B(n14624), .Z(n14341) );
  NAND U14270 ( .A(n14625), .B(n14626), .Z(n14624) );
  OR U14271 ( .A(n14627), .B(n14628), .Z(n14625) );
  AND U14272 ( .A(\stack[0][10] ), .B(\stack[1][37] ), .Z(n14340) );
  XNOR U14273 ( .A(n14347), .B(n14629), .Z(n14338) );
  XOR U14274 ( .A(n14348), .B(n14346), .Z(n14629) );
  AND U14275 ( .A(\stack[0][9] ), .B(\stack[1][38] ), .Z(n14346) );
  NAND U14276 ( .A(n14630), .B(n14631), .Z(n14348) );
  OR U14277 ( .A(n14632), .B(n14633), .Z(n14631) );
  NAND U14278 ( .A(n14634), .B(n14635), .Z(n14630) );
  NAND U14279 ( .A(n14633), .B(n14632), .Z(n14634) );
  XNOR U14280 ( .A(n14352), .B(n14636), .Z(n14347) );
  XNOR U14281 ( .A(n14353), .B(n14354), .Z(n14636) );
  AND U14282 ( .A(n14637), .B(n14638), .Z(n14354) );
  NAND U14283 ( .A(n14639), .B(n14640), .Z(n14638) );
  NANDN U14284 ( .A(n14641), .B(n14642), .Z(n14637) );
  OR U14285 ( .A(n14639), .B(n14640), .Z(n14642) );
  ANDN U14286 ( .B(\stack[1][39] ), .A(n5350), .Z(n14353) );
  XNOR U14287 ( .A(n14359), .B(n14643), .Z(n14352) );
  XNOR U14288 ( .A(n14360), .B(n14361), .Z(n14643) );
  AND U14289 ( .A(n14644), .B(n14645), .Z(n14361) );
  NANDN U14290 ( .A(n14646), .B(n14647), .Z(n14645) );
  NANDN U14291 ( .A(n14648), .B(n14649), .Z(n14644) );
  NANDN U14292 ( .A(n14647), .B(n14646), .Z(n14649) );
  ANDN U14293 ( .B(\stack[1][40] ), .A(n5326), .Z(n14360) );
  XNOR U14294 ( .A(n14366), .B(n14650), .Z(n14359) );
  XNOR U14295 ( .A(n14367), .B(n14368), .Z(n14650) );
  AND U14296 ( .A(n14651), .B(n14652), .Z(n14368) );
  NAND U14297 ( .A(n14653), .B(n14654), .Z(n14652) );
  NANDN U14298 ( .A(n14655), .B(n14656), .Z(n14651) );
  OR U14299 ( .A(n14653), .B(n14654), .Z(n14656) );
  ANDN U14300 ( .B(\stack[1][41] ), .A(n5302), .Z(n14367) );
  XNOR U14301 ( .A(n14373), .B(n14657), .Z(n14366) );
  XNOR U14302 ( .A(n14374), .B(n14375), .Z(n14657) );
  AND U14303 ( .A(n14658), .B(n14659), .Z(n14375) );
  NANDN U14304 ( .A(n14660), .B(n14661), .Z(n14659) );
  NANDN U14305 ( .A(n14662), .B(n14663), .Z(n14658) );
  NANDN U14306 ( .A(n14661), .B(n14660), .Z(n14663) );
  ANDN U14307 ( .B(\stack[1][42] ), .A(n5278), .Z(n14374) );
  XNOR U14308 ( .A(n14380), .B(n14664), .Z(n14373) );
  XNOR U14309 ( .A(n14381), .B(n14382), .Z(n14664) );
  AND U14310 ( .A(n14665), .B(n14666), .Z(n14382) );
  NAND U14311 ( .A(n14667), .B(n14668), .Z(n14666) );
  NANDN U14312 ( .A(n14669), .B(n14670), .Z(n14665) );
  OR U14313 ( .A(n14667), .B(n14668), .Z(n14670) );
  ANDN U14314 ( .B(\stack[1][43] ), .A(n5254), .Z(n14381) );
  XNOR U14315 ( .A(n14387), .B(n14671), .Z(n14380) );
  XNOR U14316 ( .A(n14388), .B(n14389), .Z(n14671) );
  AND U14317 ( .A(n14672), .B(n14673), .Z(n14389) );
  NAND U14318 ( .A(n14674), .B(n14675), .Z(n14673) );
  NAND U14319 ( .A(n14676), .B(n14677), .Z(n14672) );
  OR U14320 ( .A(n14674), .B(n14675), .Z(n14676) );
  ANDN U14321 ( .B(\stack[1][44] ), .A(n5230), .Z(n14388) );
  XNOR U14322 ( .A(n14394), .B(n14678), .Z(n14387) );
  XNOR U14323 ( .A(n14395), .B(n14397), .Z(n14678) );
  ANDN U14324 ( .B(n14679), .A(n14680), .Z(n14397) );
  ANDN U14325 ( .B(\stack[0][0] ), .A(n6276), .Z(n14679) );
  ANDN U14326 ( .B(\stack[1][45] ), .A(n5206), .Z(n14395) );
  XOR U14327 ( .A(n14400), .B(n14681), .Z(n14394) );
  NANDN U14328 ( .A(n5160), .B(\stack[1][47] ), .Z(n14681) );
  NANDN U14329 ( .A(n6276), .B(\stack[0][1] ), .Z(n14400) );
  ANDN U14330 ( .B(\stack[1][5] ), .A(n6166), .Z(n9069) );
  AND U14331 ( .A(n14682), .B(n14683), .Z(n9070) );
  NANDN U14332 ( .A(n9074), .B(n9076), .Z(n14683) );
  NANDN U14333 ( .A(n9077), .B(n14684), .Z(n14682) );
  NANDN U14334 ( .A(n9076), .B(n9074), .Z(n14684) );
  XOR U14335 ( .A(n14408), .B(n14685), .Z(n9074) );
  XNOR U14336 ( .A(n14409), .B(n14410), .Z(n14685) );
  AND U14337 ( .A(n14686), .B(n14687), .Z(n14410) );
  NAND U14338 ( .A(n14688), .B(n14689), .Z(n14687) );
  NANDN U14339 ( .A(n14690), .B(n14691), .Z(n14686) );
  OR U14340 ( .A(n14688), .B(n14689), .Z(n14691) );
  ANDN U14341 ( .B(\stack[0][40] ), .A(n5316), .Z(n14409) );
  XNOR U14342 ( .A(n14415), .B(n14692), .Z(n14408) );
  XNOR U14343 ( .A(n14416), .B(n14417), .Z(n14692) );
  AND U14344 ( .A(n14693), .B(n14694), .Z(n14417) );
  NANDN U14345 ( .A(n14695), .B(n14696), .Z(n14694) );
  NANDN U14346 ( .A(n14697), .B(n14698), .Z(n14693) );
  NANDN U14347 ( .A(n14696), .B(n14695), .Z(n14698) );
  ANDN U14348 ( .B(\stack[0][39] ), .A(n5340), .Z(n14416) );
  XNOR U14349 ( .A(n14422), .B(n14699), .Z(n14415) );
  XNOR U14350 ( .A(n14423), .B(n14424), .Z(n14699) );
  AND U14351 ( .A(n14700), .B(n14701), .Z(n14424) );
  NAND U14352 ( .A(n14702), .B(n14703), .Z(n14701) );
  NANDN U14353 ( .A(n14704), .B(n14705), .Z(n14700) );
  OR U14354 ( .A(n14702), .B(n14703), .Z(n14705) );
  ANDN U14355 ( .B(\stack[0][38] ), .A(n5364), .Z(n14423) );
  XNOR U14356 ( .A(n14429), .B(n14706), .Z(n14422) );
  XNOR U14357 ( .A(n14430), .B(n14431), .Z(n14706) );
  AND U14358 ( .A(n14707), .B(n14708), .Z(n14431) );
  NANDN U14359 ( .A(n14709), .B(n14710), .Z(n14708) );
  NANDN U14360 ( .A(n14711), .B(n14712), .Z(n14707) );
  NANDN U14361 ( .A(n14710), .B(n14709), .Z(n14712) );
  ANDN U14362 ( .B(\stack[0][37] ), .A(n5387), .Z(n14430) );
  XNOR U14363 ( .A(n14436), .B(n14713), .Z(n14429) );
  XNOR U14364 ( .A(n14437), .B(n14438), .Z(n14713) );
  AND U14365 ( .A(n14714), .B(n14715), .Z(n14438) );
  NAND U14366 ( .A(n14716), .B(n14717), .Z(n14715) );
  NANDN U14367 ( .A(n14718), .B(n14719), .Z(n14714) );
  OR U14368 ( .A(n14716), .B(n14717), .Z(n14719) );
  ANDN U14369 ( .B(\stack[1][10] ), .A(n6022), .Z(n14437) );
  XNOR U14370 ( .A(n14443), .B(n14720), .Z(n14436) );
  XNOR U14371 ( .A(n14444), .B(n14445), .Z(n14720) );
  AND U14372 ( .A(n14721), .B(n14722), .Z(n14445) );
  NANDN U14373 ( .A(n14723), .B(n14724), .Z(n14722) );
  NANDN U14374 ( .A(n14725), .B(n14726), .Z(n14721) );
  NANDN U14375 ( .A(n14724), .B(n14723), .Z(n14726) );
  ANDN U14376 ( .B(\stack[1][11] ), .A(n5998), .Z(n14444) );
  XNOR U14377 ( .A(n14450), .B(n14727), .Z(n14443) );
  XNOR U14378 ( .A(n14451), .B(n14452), .Z(n14727) );
  AND U14379 ( .A(n14728), .B(n14729), .Z(n14452) );
  NAND U14380 ( .A(n14730), .B(n14731), .Z(n14729) );
  NANDN U14381 ( .A(n14732), .B(n14733), .Z(n14728) );
  OR U14382 ( .A(n14730), .B(n14731), .Z(n14733) );
  ANDN U14383 ( .B(\stack[1][12] ), .A(n5974), .Z(n14451) );
  XNOR U14384 ( .A(n14457), .B(n14734), .Z(n14450) );
  XNOR U14385 ( .A(n14458), .B(n14459), .Z(n14734) );
  AND U14386 ( .A(n14735), .B(n14736), .Z(n14459) );
  NANDN U14387 ( .A(n14737), .B(n14738), .Z(n14736) );
  NANDN U14388 ( .A(n14739), .B(n14740), .Z(n14735) );
  NANDN U14389 ( .A(n14738), .B(n14737), .Z(n14740) );
  ANDN U14390 ( .B(\stack[1][13] ), .A(n5950), .Z(n14458) );
  XNOR U14391 ( .A(n14464), .B(n14741), .Z(n14457) );
  XNOR U14392 ( .A(n14465), .B(n14466), .Z(n14741) );
  AND U14393 ( .A(n14742), .B(n14743), .Z(n14466) );
  NAND U14394 ( .A(n14744), .B(n14745), .Z(n14743) );
  NANDN U14395 ( .A(n14746), .B(n14747), .Z(n14742) );
  OR U14396 ( .A(n14744), .B(n14745), .Z(n14747) );
  ANDN U14397 ( .B(\stack[1][14] ), .A(n5926), .Z(n14465) );
  XNOR U14398 ( .A(n14471), .B(n14748), .Z(n14464) );
  XNOR U14399 ( .A(n14472), .B(n14473), .Z(n14748) );
  AND U14400 ( .A(n14749), .B(n14750), .Z(n14473) );
  NANDN U14401 ( .A(n14751), .B(n14752), .Z(n14750) );
  NANDN U14402 ( .A(n14753), .B(n14754), .Z(n14749) );
  NANDN U14403 ( .A(n14752), .B(n14751), .Z(n14754) );
  ANDN U14404 ( .B(\stack[1][15] ), .A(n5902), .Z(n14472) );
  XNOR U14405 ( .A(n14478), .B(n14755), .Z(n14471) );
  XNOR U14406 ( .A(n14479), .B(n14480), .Z(n14755) );
  AND U14407 ( .A(n14756), .B(n14757), .Z(n14480) );
  NAND U14408 ( .A(n14758), .B(n14759), .Z(n14757) );
  NANDN U14409 ( .A(n14760), .B(n14761), .Z(n14756) );
  OR U14410 ( .A(n14758), .B(n14759), .Z(n14761) );
  ANDN U14411 ( .B(\stack[1][16] ), .A(n5878), .Z(n14479) );
  XNOR U14412 ( .A(n14485), .B(n14762), .Z(n14478) );
  XNOR U14413 ( .A(n14486), .B(n14487), .Z(n14762) );
  AND U14414 ( .A(n14763), .B(n14764), .Z(n14487) );
  NANDN U14415 ( .A(n14765), .B(n14766), .Z(n14764) );
  NANDN U14416 ( .A(n14767), .B(n14768), .Z(n14763) );
  NANDN U14417 ( .A(n14766), .B(n14765), .Z(n14768) );
  ANDN U14418 ( .B(\stack[1][17] ), .A(n5854), .Z(n14486) );
  XNOR U14419 ( .A(n14492), .B(n14769), .Z(n14485) );
  XNOR U14420 ( .A(n14493), .B(n14494), .Z(n14769) );
  AND U14421 ( .A(n14770), .B(n14771), .Z(n14494) );
  NAND U14422 ( .A(n14772), .B(n14773), .Z(n14771) );
  NANDN U14423 ( .A(n14774), .B(n14775), .Z(n14770) );
  OR U14424 ( .A(n14772), .B(n14773), .Z(n14775) );
  ANDN U14425 ( .B(\stack[1][18] ), .A(n5830), .Z(n14493) );
  XNOR U14426 ( .A(n14499), .B(n14776), .Z(n14492) );
  XNOR U14427 ( .A(n14500), .B(n14501), .Z(n14776) );
  AND U14428 ( .A(n14777), .B(n14778), .Z(n14501) );
  NANDN U14429 ( .A(n14779), .B(n14780), .Z(n14778) );
  NANDN U14430 ( .A(n14781), .B(n14782), .Z(n14777) );
  NANDN U14431 ( .A(n14780), .B(n14779), .Z(n14782) );
  ANDN U14432 ( .B(\stack[1][19] ), .A(n5806), .Z(n14500) );
  XNOR U14433 ( .A(n14506), .B(n14783), .Z(n14499) );
  XNOR U14434 ( .A(n14507), .B(n14508), .Z(n14783) );
  AND U14435 ( .A(n14784), .B(n14785), .Z(n14508) );
  NAND U14436 ( .A(n14786), .B(n14787), .Z(n14785) );
  NANDN U14437 ( .A(n14788), .B(n14789), .Z(n14784) );
  OR U14438 ( .A(n14786), .B(n14787), .Z(n14789) );
  ANDN U14439 ( .B(\stack[1][20] ), .A(n5782), .Z(n14507) );
  XNOR U14440 ( .A(n14513), .B(n14790), .Z(n14506) );
  XNOR U14441 ( .A(n14514), .B(n14515), .Z(n14790) );
  AND U14442 ( .A(n14791), .B(n14792), .Z(n14515) );
  NANDN U14443 ( .A(n14793), .B(n14794), .Z(n14792) );
  NANDN U14444 ( .A(n14795), .B(n14796), .Z(n14791) );
  NANDN U14445 ( .A(n14794), .B(n14793), .Z(n14796) );
  ANDN U14446 ( .B(\stack[1][21] ), .A(n5758), .Z(n14514) );
  XNOR U14447 ( .A(n14520), .B(n14797), .Z(n14513) );
  XNOR U14448 ( .A(n14521), .B(n14522), .Z(n14797) );
  AND U14449 ( .A(n14798), .B(n14799), .Z(n14522) );
  NAND U14450 ( .A(n14800), .B(n14801), .Z(n14799) );
  NANDN U14451 ( .A(n14802), .B(n14803), .Z(n14798) );
  OR U14452 ( .A(n14800), .B(n14801), .Z(n14803) );
  ANDN U14453 ( .B(\stack[1][22] ), .A(n5734), .Z(n14521) );
  XNOR U14454 ( .A(n14527), .B(n14804), .Z(n14520) );
  XNOR U14455 ( .A(n14528), .B(n14529), .Z(n14804) );
  AND U14456 ( .A(n14805), .B(n14806), .Z(n14529) );
  NANDN U14457 ( .A(n14807), .B(n14808), .Z(n14806) );
  NANDN U14458 ( .A(n14809), .B(n14810), .Z(n14805) );
  NANDN U14459 ( .A(n14808), .B(n14807), .Z(n14810) );
  ANDN U14460 ( .B(\stack[1][23] ), .A(n5710), .Z(n14528) );
  XNOR U14461 ( .A(n14534), .B(n14811), .Z(n14527) );
  XNOR U14462 ( .A(n14535), .B(n14536), .Z(n14811) );
  AND U14463 ( .A(n14812), .B(n14813), .Z(n14536) );
  NAND U14464 ( .A(n14814), .B(n14815), .Z(n14813) );
  NANDN U14465 ( .A(n14816), .B(n14817), .Z(n14812) );
  OR U14466 ( .A(n14814), .B(n14815), .Z(n14817) );
  ANDN U14467 ( .B(\stack[1][24] ), .A(n5686), .Z(n14535) );
  XNOR U14468 ( .A(n14541), .B(n14818), .Z(n14534) );
  XNOR U14469 ( .A(n14542), .B(n14543), .Z(n14818) );
  AND U14470 ( .A(n14819), .B(n14820), .Z(n14543) );
  NANDN U14471 ( .A(n14821), .B(n14822), .Z(n14820) );
  NANDN U14472 ( .A(n14823), .B(n14824), .Z(n14819) );
  NANDN U14473 ( .A(n14822), .B(n14821), .Z(n14824) );
  ANDN U14474 ( .B(\stack[1][25] ), .A(n5662), .Z(n14542) );
  XNOR U14475 ( .A(n14548), .B(n14825), .Z(n14541) );
  XNOR U14476 ( .A(n14549), .B(n14550), .Z(n14825) );
  AND U14477 ( .A(n14826), .B(n14827), .Z(n14550) );
  NAND U14478 ( .A(n14828), .B(n14829), .Z(n14827) );
  NANDN U14479 ( .A(n14830), .B(n14831), .Z(n14826) );
  OR U14480 ( .A(n14828), .B(n14829), .Z(n14831) );
  ANDN U14481 ( .B(\stack[1][26] ), .A(n5638), .Z(n14549) );
  XNOR U14482 ( .A(n14555), .B(n14832), .Z(n14548) );
  XNOR U14483 ( .A(n14556), .B(n14557), .Z(n14832) );
  AND U14484 ( .A(n14833), .B(n14834), .Z(n14557) );
  NANDN U14485 ( .A(n14835), .B(n14836), .Z(n14834) );
  NANDN U14486 ( .A(n14837), .B(n14838), .Z(n14833) );
  NANDN U14487 ( .A(n14836), .B(n14835), .Z(n14838) );
  ANDN U14488 ( .B(\stack[1][27] ), .A(n5614), .Z(n14556) );
  XNOR U14489 ( .A(n14562), .B(n14839), .Z(n14555) );
  XNOR U14490 ( .A(n14563), .B(n14564), .Z(n14839) );
  AND U14491 ( .A(n14840), .B(n14841), .Z(n14564) );
  NAND U14492 ( .A(n14842), .B(n14843), .Z(n14841) );
  NANDN U14493 ( .A(n14844), .B(n14845), .Z(n14840) );
  OR U14494 ( .A(n14842), .B(n14843), .Z(n14845) );
  ANDN U14495 ( .B(\stack[1][28] ), .A(n5590), .Z(n14563) );
  XNOR U14496 ( .A(n14569), .B(n14846), .Z(n14562) );
  XNOR U14497 ( .A(n14570), .B(n14571), .Z(n14846) );
  AND U14498 ( .A(n14847), .B(n14848), .Z(n14571) );
  NANDN U14499 ( .A(n14849), .B(n14850), .Z(n14848) );
  NANDN U14500 ( .A(n14851), .B(n14852), .Z(n14847) );
  NANDN U14501 ( .A(n14850), .B(n14849), .Z(n14852) );
  ANDN U14502 ( .B(\stack[1][29] ), .A(n5566), .Z(n14570) );
  XNOR U14503 ( .A(n14576), .B(n14853), .Z(n14569) );
  XNOR U14504 ( .A(n14577), .B(n14578), .Z(n14853) );
  AND U14505 ( .A(n14854), .B(n14855), .Z(n14578) );
  NAND U14506 ( .A(n14856), .B(n14857), .Z(n14855) );
  NANDN U14507 ( .A(n14858), .B(n14859), .Z(n14854) );
  OR U14508 ( .A(n14856), .B(n14857), .Z(n14859) );
  ANDN U14509 ( .B(\stack[1][30] ), .A(n5542), .Z(n14577) );
  XNOR U14510 ( .A(n14583), .B(n14860), .Z(n14576) );
  XNOR U14511 ( .A(n14584), .B(n14585), .Z(n14860) );
  AND U14512 ( .A(n14861), .B(n14862), .Z(n14585) );
  NANDN U14513 ( .A(n14863), .B(n14864), .Z(n14862) );
  NANDN U14514 ( .A(n14865), .B(n14866), .Z(n14861) );
  NANDN U14515 ( .A(n14864), .B(n14863), .Z(n14866) );
  ANDN U14516 ( .B(\stack[1][31] ), .A(n5518), .Z(n14584) );
  XNOR U14517 ( .A(n14590), .B(n14867), .Z(n14583) );
  XNOR U14518 ( .A(n14591), .B(n14592), .Z(n14867) );
  AND U14519 ( .A(n14868), .B(n14869), .Z(n14592) );
  NAND U14520 ( .A(n14870), .B(n14871), .Z(n14869) );
  NANDN U14521 ( .A(n14872), .B(n14873), .Z(n14868) );
  OR U14522 ( .A(n14870), .B(n14871), .Z(n14873) );
  ANDN U14523 ( .B(\stack[1][32] ), .A(n5494), .Z(n14591) );
  XNOR U14524 ( .A(n14597), .B(n14874), .Z(n14590) );
  XNOR U14525 ( .A(n14598), .B(n14599), .Z(n14874) );
  AND U14526 ( .A(n14875), .B(n14876), .Z(n14599) );
  NANDN U14527 ( .A(n14877), .B(n14878), .Z(n14876) );
  NANDN U14528 ( .A(n14879), .B(n14880), .Z(n14875) );
  NANDN U14529 ( .A(n14878), .B(n14877), .Z(n14880) );
  ANDN U14530 ( .B(\stack[1][33] ), .A(n5470), .Z(n14598) );
  XNOR U14531 ( .A(n14604), .B(n14881), .Z(n14597) );
  XNOR U14532 ( .A(n14605), .B(n14606), .Z(n14881) );
  AND U14533 ( .A(n14882), .B(n14883), .Z(n14606) );
  NAND U14534 ( .A(n14884), .B(n14885), .Z(n14883) );
  NANDN U14535 ( .A(n14886), .B(n14887), .Z(n14882) );
  OR U14536 ( .A(n14884), .B(n14885), .Z(n14887) );
  ANDN U14537 ( .B(\stack[1][34] ), .A(n5446), .Z(n14605) );
  XNOR U14538 ( .A(n14611), .B(n14888), .Z(n14604) );
  XNOR U14539 ( .A(n14612), .B(n14613), .Z(n14888) );
  AND U14540 ( .A(n14889), .B(n14890), .Z(n14613) );
  NANDN U14541 ( .A(n14891), .B(n14892), .Z(n14890) );
  NANDN U14542 ( .A(n14893), .B(n14894), .Z(n14889) );
  NANDN U14543 ( .A(n14892), .B(n14891), .Z(n14894) );
  ANDN U14544 ( .B(\stack[1][35] ), .A(n5422), .Z(n14612) );
  XNOR U14545 ( .A(n14618), .B(n14895), .Z(n14611) );
  XNOR U14546 ( .A(n14619), .B(n14620), .Z(n14895) );
  AND U14547 ( .A(n14896), .B(n14897), .Z(n14620) );
  NAND U14548 ( .A(n14898), .B(n14899), .Z(n14897) );
  NANDN U14549 ( .A(n14900), .B(n14901), .Z(n14896) );
  OR U14550 ( .A(n14898), .B(n14899), .Z(n14901) );
  ANDN U14551 ( .B(\stack[1][36] ), .A(n5398), .Z(n14619) );
  XNOR U14552 ( .A(n14626), .B(n14902), .Z(n14618) );
  XOR U14553 ( .A(n14627), .B(n14628), .Z(n14902) );
  NAND U14554 ( .A(n14903), .B(n14904), .Z(n14628) );
  NANDN U14555 ( .A(n14905), .B(n14906), .Z(n14904) );
  OR U14556 ( .A(n14907), .B(n14908), .Z(n14906) );
  AND U14557 ( .A(\stack[0][9] ), .B(\stack[1][37] ), .Z(n14627) );
  XNOR U14558 ( .A(n14633), .B(n14909), .Z(n14626) );
  XNOR U14559 ( .A(n14632), .B(n14635), .Z(n14909) );
  AND U14560 ( .A(\stack[0][8] ), .B(\stack[1][38] ), .Z(n14635) );
  AND U14561 ( .A(n14910), .B(n14911), .Z(n14632) );
  NAND U14562 ( .A(n14912), .B(n14913), .Z(n14911) );
  OR U14563 ( .A(n14914), .B(n14915), .Z(n14912) );
  XNOR U14564 ( .A(n14639), .B(n14916), .Z(n14633) );
  XNOR U14565 ( .A(n14640), .B(n14641), .Z(n14916) );
  AND U14566 ( .A(n14917), .B(n14918), .Z(n14641) );
  NANDN U14567 ( .A(n14919), .B(n14920), .Z(n14918) );
  NANDN U14568 ( .A(n14921), .B(n14922), .Z(n14917) );
  NANDN U14569 ( .A(n14920), .B(n14919), .Z(n14922) );
  ANDN U14570 ( .B(\stack[1][39] ), .A(n5326), .Z(n14640) );
  XNOR U14571 ( .A(n14646), .B(n14923), .Z(n14639) );
  XNOR U14572 ( .A(n14647), .B(n14648), .Z(n14923) );
  AND U14573 ( .A(n14924), .B(n14925), .Z(n14648) );
  NAND U14574 ( .A(n14926), .B(n14927), .Z(n14925) );
  NANDN U14575 ( .A(n14928), .B(n14929), .Z(n14924) );
  OR U14576 ( .A(n14926), .B(n14927), .Z(n14929) );
  ANDN U14577 ( .B(\stack[1][40] ), .A(n5302), .Z(n14647) );
  XNOR U14578 ( .A(n14653), .B(n14930), .Z(n14646) );
  XNOR U14579 ( .A(n14654), .B(n14655), .Z(n14930) );
  AND U14580 ( .A(n14931), .B(n14932), .Z(n14655) );
  NANDN U14581 ( .A(n14933), .B(n14934), .Z(n14932) );
  NANDN U14582 ( .A(n14935), .B(n14936), .Z(n14931) );
  NANDN U14583 ( .A(n14934), .B(n14933), .Z(n14936) );
  ANDN U14584 ( .B(\stack[1][41] ), .A(n5278), .Z(n14654) );
  XNOR U14585 ( .A(n14660), .B(n14937), .Z(n14653) );
  XNOR U14586 ( .A(n14661), .B(n14662), .Z(n14937) );
  AND U14587 ( .A(n14938), .B(n14939), .Z(n14662) );
  NAND U14588 ( .A(n14940), .B(n14941), .Z(n14939) );
  NANDN U14589 ( .A(n14942), .B(n14943), .Z(n14938) );
  OR U14590 ( .A(n14940), .B(n14941), .Z(n14943) );
  ANDN U14591 ( .B(\stack[1][42] ), .A(n5254), .Z(n14661) );
  XNOR U14592 ( .A(n14667), .B(n14944), .Z(n14660) );
  XNOR U14593 ( .A(n14668), .B(n14669), .Z(n14944) );
  AND U14594 ( .A(n14945), .B(n14946), .Z(n14669) );
  NAND U14595 ( .A(n14947), .B(n14948), .Z(n14946) );
  NAND U14596 ( .A(n14949), .B(n14950), .Z(n14945) );
  OR U14597 ( .A(n14947), .B(n14948), .Z(n14949) );
  ANDN U14598 ( .B(\stack[1][43] ), .A(n5230), .Z(n14668) );
  XNOR U14599 ( .A(n14674), .B(n14951), .Z(n14667) );
  XNOR U14600 ( .A(n14675), .B(n14677), .Z(n14951) );
  ANDN U14601 ( .B(n14952), .A(n14953), .Z(n14677) );
  ANDN U14602 ( .B(\stack[0][0] ), .A(n6252), .Z(n14952) );
  ANDN U14603 ( .B(\stack[1][44] ), .A(n5206), .Z(n14675) );
  XOR U14604 ( .A(n14680), .B(n14954), .Z(n14674) );
  NANDN U14605 ( .A(n5160), .B(\stack[1][46] ), .Z(n14954) );
  NANDN U14606 ( .A(n6252), .B(\stack[0][1] ), .Z(n14680) );
  ANDN U14607 ( .B(\stack[0][41] ), .A(n5292), .Z(n9076) );
  AND U14608 ( .A(n14955), .B(n14956), .Z(n9077) );
  NANDN U14609 ( .A(n9084), .B(n14957), .Z(n14955) );
  NANDN U14610 ( .A(n9083), .B(n9081), .Z(n14957) );
  XNOR U14611 ( .A(n14688), .B(n14958), .Z(n9081) );
  XNOR U14612 ( .A(n14689), .B(n14690), .Z(n14958) );
  AND U14613 ( .A(n14959), .B(n14960), .Z(n14690) );
  NANDN U14614 ( .A(n14961), .B(n14962), .Z(n14960) );
  NANDN U14615 ( .A(n14963), .B(n14964), .Z(n14959) );
  NANDN U14616 ( .A(n14962), .B(n14961), .Z(n14964) );
  ANDN U14617 ( .B(\stack[0][39] ), .A(n5316), .Z(n14689) );
  XNOR U14618 ( .A(n14695), .B(n14965), .Z(n14688) );
  XNOR U14619 ( .A(n14696), .B(n14697), .Z(n14965) );
  AND U14620 ( .A(n14966), .B(n14967), .Z(n14697) );
  NAND U14621 ( .A(n14968), .B(n14969), .Z(n14967) );
  NANDN U14622 ( .A(n14970), .B(n14971), .Z(n14966) );
  OR U14623 ( .A(n14968), .B(n14969), .Z(n14971) );
  ANDN U14624 ( .B(\stack[0][38] ), .A(n5340), .Z(n14696) );
  XNOR U14625 ( .A(n14702), .B(n14972), .Z(n14695) );
  XNOR U14626 ( .A(n14703), .B(n14704), .Z(n14972) );
  AND U14627 ( .A(n14973), .B(n14974), .Z(n14704) );
  NANDN U14628 ( .A(n14975), .B(n14976), .Z(n14974) );
  NANDN U14629 ( .A(n14977), .B(n14978), .Z(n14973) );
  NANDN U14630 ( .A(n14976), .B(n14975), .Z(n14978) );
  ANDN U14631 ( .B(\stack[0][37] ), .A(n5364), .Z(n14703) );
  XNOR U14632 ( .A(n14709), .B(n14979), .Z(n14702) );
  XNOR U14633 ( .A(n14710), .B(n14711), .Z(n14979) );
  AND U14634 ( .A(n14980), .B(n14981), .Z(n14711) );
  NAND U14635 ( .A(n14982), .B(n14983), .Z(n14981) );
  NANDN U14636 ( .A(n14984), .B(n14985), .Z(n14980) );
  OR U14637 ( .A(n14982), .B(n14983), .Z(n14985) );
  ANDN U14638 ( .B(\stack[0][36] ), .A(n5387), .Z(n14710) );
  XNOR U14639 ( .A(n14716), .B(n14986), .Z(n14709) );
  XNOR U14640 ( .A(n14717), .B(n14718), .Z(n14986) );
  AND U14641 ( .A(n14987), .B(n14988), .Z(n14718) );
  NANDN U14642 ( .A(n14989), .B(n14990), .Z(n14988) );
  NANDN U14643 ( .A(n14991), .B(n14992), .Z(n14987) );
  NANDN U14644 ( .A(n14990), .B(n14989), .Z(n14992) );
  ANDN U14645 ( .B(\stack[1][10] ), .A(n5998), .Z(n14717) );
  XNOR U14646 ( .A(n14723), .B(n14993), .Z(n14716) );
  XNOR U14647 ( .A(n14724), .B(n14725), .Z(n14993) );
  AND U14648 ( .A(n14994), .B(n14995), .Z(n14725) );
  NAND U14649 ( .A(n14996), .B(n14997), .Z(n14995) );
  NANDN U14650 ( .A(n14998), .B(n14999), .Z(n14994) );
  OR U14651 ( .A(n14996), .B(n14997), .Z(n14999) );
  ANDN U14652 ( .B(\stack[1][11] ), .A(n5974), .Z(n14724) );
  XNOR U14653 ( .A(n14730), .B(n15000), .Z(n14723) );
  XNOR U14654 ( .A(n14731), .B(n14732), .Z(n15000) );
  AND U14655 ( .A(n15001), .B(n15002), .Z(n14732) );
  NANDN U14656 ( .A(n15003), .B(n15004), .Z(n15002) );
  NANDN U14657 ( .A(n15005), .B(n15006), .Z(n15001) );
  NANDN U14658 ( .A(n15004), .B(n15003), .Z(n15006) );
  ANDN U14659 ( .B(\stack[1][12] ), .A(n5950), .Z(n14731) );
  XNOR U14660 ( .A(n14737), .B(n15007), .Z(n14730) );
  XNOR U14661 ( .A(n14738), .B(n14739), .Z(n15007) );
  AND U14662 ( .A(n15008), .B(n15009), .Z(n14739) );
  NAND U14663 ( .A(n15010), .B(n15011), .Z(n15009) );
  NANDN U14664 ( .A(n15012), .B(n15013), .Z(n15008) );
  OR U14665 ( .A(n15010), .B(n15011), .Z(n15013) );
  ANDN U14666 ( .B(\stack[1][13] ), .A(n5926), .Z(n14738) );
  XNOR U14667 ( .A(n14744), .B(n15014), .Z(n14737) );
  XNOR U14668 ( .A(n14745), .B(n14746), .Z(n15014) );
  AND U14669 ( .A(n15015), .B(n15016), .Z(n14746) );
  NANDN U14670 ( .A(n15017), .B(n15018), .Z(n15016) );
  NANDN U14671 ( .A(n15019), .B(n15020), .Z(n15015) );
  NANDN U14672 ( .A(n15018), .B(n15017), .Z(n15020) );
  ANDN U14673 ( .B(\stack[1][14] ), .A(n5902), .Z(n14745) );
  XNOR U14674 ( .A(n14751), .B(n15021), .Z(n14744) );
  XNOR U14675 ( .A(n14752), .B(n14753), .Z(n15021) );
  AND U14676 ( .A(n15022), .B(n15023), .Z(n14753) );
  NAND U14677 ( .A(n15024), .B(n15025), .Z(n15023) );
  NANDN U14678 ( .A(n15026), .B(n15027), .Z(n15022) );
  OR U14679 ( .A(n15024), .B(n15025), .Z(n15027) );
  ANDN U14680 ( .B(\stack[1][15] ), .A(n5878), .Z(n14752) );
  XNOR U14681 ( .A(n14758), .B(n15028), .Z(n14751) );
  XNOR U14682 ( .A(n14759), .B(n14760), .Z(n15028) );
  AND U14683 ( .A(n15029), .B(n15030), .Z(n14760) );
  NANDN U14684 ( .A(n15031), .B(n15032), .Z(n15030) );
  NANDN U14685 ( .A(n15033), .B(n15034), .Z(n15029) );
  NANDN U14686 ( .A(n15032), .B(n15031), .Z(n15034) );
  ANDN U14687 ( .B(\stack[1][16] ), .A(n5854), .Z(n14759) );
  XNOR U14688 ( .A(n14765), .B(n15035), .Z(n14758) );
  XNOR U14689 ( .A(n14766), .B(n14767), .Z(n15035) );
  AND U14690 ( .A(n15036), .B(n15037), .Z(n14767) );
  NAND U14691 ( .A(n15038), .B(n15039), .Z(n15037) );
  NANDN U14692 ( .A(n15040), .B(n15041), .Z(n15036) );
  OR U14693 ( .A(n15038), .B(n15039), .Z(n15041) );
  ANDN U14694 ( .B(\stack[1][17] ), .A(n5830), .Z(n14766) );
  XNOR U14695 ( .A(n14772), .B(n15042), .Z(n14765) );
  XNOR U14696 ( .A(n14773), .B(n14774), .Z(n15042) );
  AND U14697 ( .A(n15043), .B(n15044), .Z(n14774) );
  NANDN U14698 ( .A(n15045), .B(n15046), .Z(n15044) );
  NANDN U14699 ( .A(n15047), .B(n15048), .Z(n15043) );
  NANDN U14700 ( .A(n15046), .B(n15045), .Z(n15048) );
  ANDN U14701 ( .B(\stack[1][18] ), .A(n5806), .Z(n14773) );
  XNOR U14702 ( .A(n14779), .B(n15049), .Z(n14772) );
  XNOR U14703 ( .A(n14780), .B(n14781), .Z(n15049) );
  AND U14704 ( .A(n15050), .B(n15051), .Z(n14781) );
  NAND U14705 ( .A(n15052), .B(n15053), .Z(n15051) );
  NANDN U14706 ( .A(n15054), .B(n15055), .Z(n15050) );
  OR U14707 ( .A(n15052), .B(n15053), .Z(n15055) );
  ANDN U14708 ( .B(\stack[1][19] ), .A(n5782), .Z(n14780) );
  XNOR U14709 ( .A(n14786), .B(n15056), .Z(n14779) );
  XNOR U14710 ( .A(n14787), .B(n14788), .Z(n15056) );
  AND U14711 ( .A(n15057), .B(n15058), .Z(n14788) );
  NANDN U14712 ( .A(n15059), .B(n15060), .Z(n15058) );
  NANDN U14713 ( .A(n15061), .B(n15062), .Z(n15057) );
  NANDN U14714 ( .A(n15060), .B(n15059), .Z(n15062) );
  ANDN U14715 ( .B(\stack[1][20] ), .A(n5758), .Z(n14787) );
  XNOR U14716 ( .A(n14793), .B(n15063), .Z(n14786) );
  XNOR U14717 ( .A(n14794), .B(n14795), .Z(n15063) );
  AND U14718 ( .A(n15064), .B(n15065), .Z(n14795) );
  NAND U14719 ( .A(n15066), .B(n15067), .Z(n15065) );
  NANDN U14720 ( .A(n15068), .B(n15069), .Z(n15064) );
  OR U14721 ( .A(n15066), .B(n15067), .Z(n15069) );
  ANDN U14722 ( .B(\stack[1][21] ), .A(n5734), .Z(n14794) );
  XNOR U14723 ( .A(n14800), .B(n15070), .Z(n14793) );
  XNOR U14724 ( .A(n14801), .B(n14802), .Z(n15070) );
  AND U14725 ( .A(n15071), .B(n15072), .Z(n14802) );
  NANDN U14726 ( .A(n15073), .B(n15074), .Z(n15072) );
  NANDN U14727 ( .A(n15075), .B(n15076), .Z(n15071) );
  NANDN U14728 ( .A(n15074), .B(n15073), .Z(n15076) );
  ANDN U14729 ( .B(\stack[1][22] ), .A(n5710), .Z(n14801) );
  XNOR U14730 ( .A(n14807), .B(n15077), .Z(n14800) );
  XNOR U14731 ( .A(n14808), .B(n14809), .Z(n15077) );
  AND U14732 ( .A(n15078), .B(n15079), .Z(n14809) );
  NAND U14733 ( .A(n15080), .B(n15081), .Z(n15079) );
  NANDN U14734 ( .A(n15082), .B(n15083), .Z(n15078) );
  OR U14735 ( .A(n15080), .B(n15081), .Z(n15083) );
  ANDN U14736 ( .B(\stack[1][23] ), .A(n5686), .Z(n14808) );
  XNOR U14737 ( .A(n14814), .B(n15084), .Z(n14807) );
  XNOR U14738 ( .A(n14815), .B(n14816), .Z(n15084) );
  AND U14739 ( .A(n15085), .B(n15086), .Z(n14816) );
  NANDN U14740 ( .A(n15087), .B(n15088), .Z(n15086) );
  NANDN U14741 ( .A(n15089), .B(n15090), .Z(n15085) );
  NANDN U14742 ( .A(n15088), .B(n15087), .Z(n15090) );
  ANDN U14743 ( .B(\stack[1][24] ), .A(n5662), .Z(n14815) );
  XNOR U14744 ( .A(n14821), .B(n15091), .Z(n14814) );
  XNOR U14745 ( .A(n14822), .B(n14823), .Z(n15091) );
  AND U14746 ( .A(n15092), .B(n15093), .Z(n14823) );
  NAND U14747 ( .A(n15094), .B(n15095), .Z(n15093) );
  NANDN U14748 ( .A(n15096), .B(n15097), .Z(n15092) );
  OR U14749 ( .A(n15094), .B(n15095), .Z(n15097) );
  ANDN U14750 ( .B(\stack[1][25] ), .A(n5638), .Z(n14822) );
  XNOR U14751 ( .A(n14828), .B(n15098), .Z(n14821) );
  XNOR U14752 ( .A(n14829), .B(n14830), .Z(n15098) );
  AND U14753 ( .A(n15099), .B(n15100), .Z(n14830) );
  NANDN U14754 ( .A(n15101), .B(n15102), .Z(n15100) );
  NANDN U14755 ( .A(n15103), .B(n15104), .Z(n15099) );
  NANDN U14756 ( .A(n15102), .B(n15101), .Z(n15104) );
  ANDN U14757 ( .B(\stack[1][26] ), .A(n5614), .Z(n14829) );
  XNOR U14758 ( .A(n14835), .B(n15105), .Z(n14828) );
  XNOR U14759 ( .A(n14836), .B(n14837), .Z(n15105) );
  AND U14760 ( .A(n15106), .B(n15107), .Z(n14837) );
  NAND U14761 ( .A(n15108), .B(n15109), .Z(n15107) );
  NANDN U14762 ( .A(n15110), .B(n15111), .Z(n15106) );
  OR U14763 ( .A(n15108), .B(n15109), .Z(n15111) );
  ANDN U14764 ( .B(\stack[1][27] ), .A(n5590), .Z(n14836) );
  XNOR U14765 ( .A(n14842), .B(n15112), .Z(n14835) );
  XNOR U14766 ( .A(n14843), .B(n14844), .Z(n15112) );
  AND U14767 ( .A(n15113), .B(n15114), .Z(n14844) );
  NANDN U14768 ( .A(n15115), .B(n15116), .Z(n15114) );
  NANDN U14769 ( .A(n15117), .B(n15118), .Z(n15113) );
  NANDN U14770 ( .A(n15116), .B(n15115), .Z(n15118) );
  ANDN U14771 ( .B(\stack[1][28] ), .A(n5566), .Z(n14843) );
  XNOR U14772 ( .A(n14849), .B(n15119), .Z(n14842) );
  XNOR U14773 ( .A(n14850), .B(n14851), .Z(n15119) );
  AND U14774 ( .A(n15120), .B(n15121), .Z(n14851) );
  NAND U14775 ( .A(n15122), .B(n15123), .Z(n15121) );
  NANDN U14776 ( .A(n15124), .B(n15125), .Z(n15120) );
  OR U14777 ( .A(n15122), .B(n15123), .Z(n15125) );
  ANDN U14778 ( .B(\stack[1][29] ), .A(n5542), .Z(n14850) );
  XNOR U14779 ( .A(n14856), .B(n15126), .Z(n14849) );
  XNOR U14780 ( .A(n14857), .B(n14858), .Z(n15126) );
  AND U14781 ( .A(n15127), .B(n15128), .Z(n14858) );
  NANDN U14782 ( .A(n15129), .B(n15130), .Z(n15128) );
  NANDN U14783 ( .A(n15131), .B(n15132), .Z(n15127) );
  NANDN U14784 ( .A(n15130), .B(n15129), .Z(n15132) );
  ANDN U14785 ( .B(\stack[1][30] ), .A(n5518), .Z(n14857) );
  XNOR U14786 ( .A(n14863), .B(n15133), .Z(n14856) );
  XNOR U14787 ( .A(n14864), .B(n14865), .Z(n15133) );
  AND U14788 ( .A(n15134), .B(n15135), .Z(n14865) );
  NAND U14789 ( .A(n15136), .B(n15137), .Z(n15135) );
  NANDN U14790 ( .A(n15138), .B(n15139), .Z(n15134) );
  OR U14791 ( .A(n15136), .B(n15137), .Z(n15139) );
  ANDN U14792 ( .B(\stack[1][31] ), .A(n5494), .Z(n14864) );
  XNOR U14793 ( .A(n14870), .B(n15140), .Z(n14863) );
  XNOR U14794 ( .A(n14871), .B(n14872), .Z(n15140) );
  AND U14795 ( .A(n15141), .B(n15142), .Z(n14872) );
  NANDN U14796 ( .A(n15143), .B(n15144), .Z(n15142) );
  NANDN U14797 ( .A(n15145), .B(n15146), .Z(n15141) );
  NANDN U14798 ( .A(n15144), .B(n15143), .Z(n15146) );
  ANDN U14799 ( .B(\stack[1][32] ), .A(n5470), .Z(n14871) );
  XNOR U14800 ( .A(n14877), .B(n15147), .Z(n14870) );
  XNOR U14801 ( .A(n14878), .B(n14879), .Z(n15147) );
  AND U14802 ( .A(n15148), .B(n15149), .Z(n14879) );
  NAND U14803 ( .A(n15150), .B(n15151), .Z(n15149) );
  NANDN U14804 ( .A(n15152), .B(n15153), .Z(n15148) );
  OR U14805 ( .A(n15150), .B(n15151), .Z(n15153) );
  ANDN U14806 ( .B(\stack[1][33] ), .A(n5446), .Z(n14878) );
  XNOR U14807 ( .A(n14884), .B(n15154), .Z(n14877) );
  XNOR U14808 ( .A(n14885), .B(n14886), .Z(n15154) );
  AND U14809 ( .A(n15155), .B(n15156), .Z(n14886) );
  NANDN U14810 ( .A(n15157), .B(n15158), .Z(n15156) );
  NANDN U14811 ( .A(n15159), .B(n15160), .Z(n15155) );
  NANDN U14812 ( .A(n15158), .B(n15157), .Z(n15160) );
  ANDN U14813 ( .B(\stack[1][34] ), .A(n5422), .Z(n14885) );
  XNOR U14814 ( .A(n14891), .B(n15161), .Z(n14884) );
  XNOR U14815 ( .A(n14892), .B(n14893), .Z(n15161) );
  AND U14816 ( .A(n15162), .B(n15163), .Z(n14893) );
  NAND U14817 ( .A(n15164), .B(n15165), .Z(n15163) );
  NANDN U14818 ( .A(n15166), .B(n15167), .Z(n15162) );
  OR U14819 ( .A(n15164), .B(n15165), .Z(n15167) );
  ANDN U14820 ( .B(\stack[1][35] ), .A(n5398), .Z(n14892) );
  XNOR U14821 ( .A(n14898), .B(n15168), .Z(n14891) );
  XNOR U14822 ( .A(n14899), .B(n14900), .Z(n15168) );
  AND U14823 ( .A(n15169), .B(n15170), .Z(n14900) );
  NANDN U14824 ( .A(n15171), .B(n15172), .Z(n15170) );
  NANDN U14825 ( .A(n15173), .B(n15174), .Z(n15169) );
  NANDN U14826 ( .A(n15172), .B(n15171), .Z(n15174) );
  ANDN U14827 ( .B(\stack[1][36] ), .A(n5374), .Z(n14899) );
  XNOR U14828 ( .A(n14905), .B(n15175), .Z(n14898) );
  XOR U14829 ( .A(n14907), .B(n14908), .Z(n15175) );
  NAND U14830 ( .A(n15176), .B(n15177), .Z(n14908) );
  NAND U14831 ( .A(n15178), .B(n15179), .Z(n15177) );
  OR U14832 ( .A(n15180), .B(n15181), .Z(n15178) );
  AND U14833 ( .A(\stack[0][8] ), .B(\stack[1][37] ), .Z(n14907) );
  XNOR U14834 ( .A(n14914), .B(n15182), .Z(n14905) );
  XOR U14835 ( .A(n14915), .B(n14913), .Z(n15182) );
  AND U14836 ( .A(\stack[0][7] ), .B(\stack[1][38] ), .Z(n14913) );
  NAND U14837 ( .A(n15183), .B(n15184), .Z(n14915) );
  OR U14838 ( .A(n15185), .B(n15186), .Z(n15184) );
  NAND U14839 ( .A(n15187), .B(n15188), .Z(n15183) );
  NAND U14840 ( .A(n15186), .B(n15185), .Z(n15187) );
  XNOR U14841 ( .A(n14919), .B(n15189), .Z(n14914) );
  XNOR U14842 ( .A(n14920), .B(n14921), .Z(n15189) );
  AND U14843 ( .A(n15190), .B(n15191), .Z(n14921) );
  NAND U14844 ( .A(n15192), .B(n15193), .Z(n15191) );
  NANDN U14845 ( .A(n15194), .B(n15195), .Z(n15190) );
  OR U14846 ( .A(n15192), .B(n15193), .Z(n15195) );
  ANDN U14847 ( .B(\stack[1][39] ), .A(n5302), .Z(n14920) );
  XNOR U14848 ( .A(n14926), .B(n15196), .Z(n14919) );
  XNOR U14849 ( .A(n14927), .B(n14928), .Z(n15196) );
  AND U14850 ( .A(n15197), .B(n15198), .Z(n14928) );
  NANDN U14851 ( .A(n15199), .B(n15200), .Z(n15198) );
  NANDN U14852 ( .A(n15201), .B(n15202), .Z(n15197) );
  NANDN U14853 ( .A(n15200), .B(n15199), .Z(n15202) );
  ANDN U14854 ( .B(\stack[1][40] ), .A(n5278), .Z(n14927) );
  XNOR U14855 ( .A(n14933), .B(n15203), .Z(n14926) );
  XNOR U14856 ( .A(n14934), .B(n14935), .Z(n15203) );
  AND U14857 ( .A(n15204), .B(n15205), .Z(n14935) );
  NAND U14858 ( .A(n15206), .B(n15207), .Z(n15205) );
  NANDN U14859 ( .A(n15208), .B(n15209), .Z(n15204) );
  OR U14860 ( .A(n15206), .B(n15207), .Z(n15209) );
  ANDN U14861 ( .B(\stack[1][41] ), .A(n5254), .Z(n14934) );
  XNOR U14862 ( .A(n14940), .B(n15210), .Z(n14933) );
  XNOR U14863 ( .A(n14941), .B(n14942), .Z(n15210) );
  AND U14864 ( .A(n15211), .B(n15212), .Z(n14942) );
  NAND U14865 ( .A(n15213), .B(n15214), .Z(n15212) );
  NAND U14866 ( .A(n15215), .B(n15216), .Z(n15211) );
  OR U14867 ( .A(n15213), .B(n15214), .Z(n15215) );
  ANDN U14868 ( .B(\stack[1][42] ), .A(n5230), .Z(n14941) );
  XNOR U14869 ( .A(n14947), .B(n15217), .Z(n14940) );
  XNOR U14870 ( .A(n14948), .B(n14950), .Z(n15217) );
  ANDN U14871 ( .B(n15218), .A(n15219), .Z(n14950) );
  ANDN U14872 ( .B(\stack[0][0] ), .A(n6228), .Z(n15218) );
  ANDN U14873 ( .B(\stack[1][43] ), .A(n5206), .Z(n14948) );
  XOR U14874 ( .A(n14953), .B(n15220), .Z(n14947) );
  NANDN U14875 ( .A(n5160), .B(\stack[1][45] ), .Z(n15220) );
  NANDN U14876 ( .A(n6228), .B(\stack[0][1] ), .Z(n14953) );
  ANDN U14877 ( .B(\stack[1][5] ), .A(n6118), .Z(n9083) );
  AND U14878 ( .A(n15221), .B(n15222), .Z(n9084) );
  NANDN U14879 ( .A(n9088), .B(n9090), .Z(n15222) );
  NANDN U14880 ( .A(n9091), .B(n15223), .Z(n15221) );
  NANDN U14881 ( .A(n9090), .B(n9088), .Z(n15223) );
  XOR U14882 ( .A(n14961), .B(n15224), .Z(n9088) );
  XNOR U14883 ( .A(n14962), .B(n14963), .Z(n15224) );
  AND U14884 ( .A(n15225), .B(n15226), .Z(n14963) );
  NAND U14885 ( .A(n15227), .B(n15228), .Z(n15226) );
  NANDN U14886 ( .A(n15229), .B(n15230), .Z(n15225) );
  OR U14887 ( .A(n15227), .B(n15228), .Z(n15230) );
  ANDN U14888 ( .B(\stack[0][38] ), .A(n5316), .Z(n14962) );
  XNOR U14889 ( .A(n14968), .B(n15231), .Z(n14961) );
  XNOR U14890 ( .A(n14969), .B(n14970), .Z(n15231) );
  AND U14891 ( .A(n15232), .B(n15233), .Z(n14970) );
  NANDN U14892 ( .A(n15234), .B(n15235), .Z(n15233) );
  NANDN U14893 ( .A(n15236), .B(n15237), .Z(n15232) );
  NANDN U14894 ( .A(n15235), .B(n15234), .Z(n15237) );
  ANDN U14895 ( .B(\stack[0][37] ), .A(n5340), .Z(n14969) );
  XNOR U14896 ( .A(n14975), .B(n15238), .Z(n14968) );
  XNOR U14897 ( .A(n14976), .B(n14977), .Z(n15238) );
  AND U14898 ( .A(n15239), .B(n15240), .Z(n14977) );
  NAND U14899 ( .A(n15241), .B(n15242), .Z(n15240) );
  NANDN U14900 ( .A(n15243), .B(n15244), .Z(n15239) );
  OR U14901 ( .A(n15241), .B(n15242), .Z(n15244) );
  ANDN U14902 ( .B(\stack[0][36] ), .A(n5364), .Z(n14976) );
  XNOR U14903 ( .A(n14982), .B(n15245), .Z(n14975) );
  XNOR U14904 ( .A(n14983), .B(n14984), .Z(n15245) );
  AND U14905 ( .A(n15246), .B(n15247), .Z(n14984) );
  NANDN U14906 ( .A(n15248), .B(n15249), .Z(n15247) );
  NANDN U14907 ( .A(n15250), .B(n15251), .Z(n15246) );
  NANDN U14908 ( .A(n15249), .B(n15248), .Z(n15251) );
  ANDN U14909 ( .B(\stack[0][35] ), .A(n5387), .Z(n14983) );
  XNOR U14910 ( .A(n14989), .B(n15252), .Z(n14982) );
  XNOR U14911 ( .A(n14990), .B(n14991), .Z(n15252) );
  AND U14912 ( .A(n15253), .B(n15254), .Z(n14991) );
  NAND U14913 ( .A(n15255), .B(n15256), .Z(n15254) );
  NANDN U14914 ( .A(n15257), .B(n15258), .Z(n15253) );
  OR U14915 ( .A(n15255), .B(n15256), .Z(n15258) );
  ANDN U14916 ( .B(\stack[1][10] ), .A(n5974), .Z(n14990) );
  XNOR U14917 ( .A(n14996), .B(n15259), .Z(n14989) );
  XNOR U14918 ( .A(n14997), .B(n14998), .Z(n15259) );
  AND U14919 ( .A(n15260), .B(n15261), .Z(n14998) );
  NANDN U14920 ( .A(n15262), .B(n15263), .Z(n15261) );
  NANDN U14921 ( .A(n15264), .B(n15265), .Z(n15260) );
  NANDN U14922 ( .A(n15263), .B(n15262), .Z(n15265) );
  ANDN U14923 ( .B(\stack[1][11] ), .A(n5950), .Z(n14997) );
  XNOR U14924 ( .A(n15003), .B(n15266), .Z(n14996) );
  XNOR U14925 ( .A(n15004), .B(n15005), .Z(n15266) );
  AND U14926 ( .A(n15267), .B(n15268), .Z(n15005) );
  NAND U14927 ( .A(n15269), .B(n15270), .Z(n15268) );
  NANDN U14928 ( .A(n15271), .B(n15272), .Z(n15267) );
  OR U14929 ( .A(n15269), .B(n15270), .Z(n15272) );
  ANDN U14930 ( .B(\stack[1][12] ), .A(n5926), .Z(n15004) );
  XNOR U14931 ( .A(n15010), .B(n15273), .Z(n15003) );
  XNOR U14932 ( .A(n15011), .B(n15012), .Z(n15273) );
  AND U14933 ( .A(n15274), .B(n15275), .Z(n15012) );
  NANDN U14934 ( .A(n15276), .B(n15277), .Z(n15275) );
  NANDN U14935 ( .A(n15278), .B(n15279), .Z(n15274) );
  NANDN U14936 ( .A(n15277), .B(n15276), .Z(n15279) );
  ANDN U14937 ( .B(\stack[1][13] ), .A(n5902), .Z(n15011) );
  XNOR U14938 ( .A(n15017), .B(n15280), .Z(n15010) );
  XNOR U14939 ( .A(n15018), .B(n15019), .Z(n15280) );
  AND U14940 ( .A(n15281), .B(n15282), .Z(n15019) );
  NAND U14941 ( .A(n15283), .B(n15284), .Z(n15282) );
  NANDN U14942 ( .A(n15285), .B(n15286), .Z(n15281) );
  OR U14943 ( .A(n15283), .B(n15284), .Z(n15286) );
  ANDN U14944 ( .B(\stack[1][14] ), .A(n5878), .Z(n15018) );
  XNOR U14945 ( .A(n15024), .B(n15287), .Z(n15017) );
  XNOR U14946 ( .A(n15025), .B(n15026), .Z(n15287) );
  AND U14947 ( .A(n15288), .B(n15289), .Z(n15026) );
  NANDN U14948 ( .A(n15290), .B(n15291), .Z(n15289) );
  NANDN U14949 ( .A(n15292), .B(n15293), .Z(n15288) );
  NANDN U14950 ( .A(n15291), .B(n15290), .Z(n15293) );
  ANDN U14951 ( .B(\stack[1][15] ), .A(n5854), .Z(n15025) );
  XNOR U14952 ( .A(n15031), .B(n15294), .Z(n15024) );
  XNOR U14953 ( .A(n15032), .B(n15033), .Z(n15294) );
  AND U14954 ( .A(n15295), .B(n15296), .Z(n15033) );
  NAND U14955 ( .A(n15297), .B(n15298), .Z(n15296) );
  NANDN U14956 ( .A(n15299), .B(n15300), .Z(n15295) );
  OR U14957 ( .A(n15297), .B(n15298), .Z(n15300) );
  ANDN U14958 ( .B(\stack[1][16] ), .A(n5830), .Z(n15032) );
  XNOR U14959 ( .A(n15038), .B(n15301), .Z(n15031) );
  XNOR U14960 ( .A(n15039), .B(n15040), .Z(n15301) );
  AND U14961 ( .A(n15302), .B(n15303), .Z(n15040) );
  NANDN U14962 ( .A(n15304), .B(n15305), .Z(n15303) );
  NANDN U14963 ( .A(n15306), .B(n15307), .Z(n15302) );
  NANDN U14964 ( .A(n15305), .B(n15304), .Z(n15307) );
  ANDN U14965 ( .B(\stack[1][17] ), .A(n5806), .Z(n15039) );
  XNOR U14966 ( .A(n15045), .B(n15308), .Z(n15038) );
  XNOR U14967 ( .A(n15046), .B(n15047), .Z(n15308) );
  AND U14968 ( .A(n15309), .B(n15310), .Z(n15047) );
  NAND U14969 ( .A(n15311), .B(n15312), .Z(n15310) );
  NANDN U14970 ( .A(n15313), .B(n15314), .Z(n15309) );
  OR U14971 ( .A(n15311), .B(n15312), .Z(n15314) );
  ANDN U14972 ( .B(\stack[1][18] ), .A(n5782), .Z(n15046) );
  XNOR U14973 ( .A(n15052), .B(n15315), .Z(n15045) );
  XNOR U14974 ( .A(n15053), .B(n15054), .Z(n15315) );
  AND U14975 ( .A(n15316), .B(n15317), .Z(n15054) );
  NANDN U14976 ( .A(n15318), .B(n15319), .Z(n15317) );
  NANDN U14977 ( .A(n15320), .B(n15321), .Z(n15316) );
  NANDN U14978 ( .A(n15319), .B(n15318), .Z(n15321) );
  ANDN U14979 ( .B(\stack[1][19] ), .A(n5758), .Z(n15053) );
  XNOR U14980 ( .A(n15059), .B(n15322), .Z(n15052) );
  XNOR U14981 ( .A(n15060), .B(n15061), .Z(n15322) );
  AND U14982 ( .A(n15323), .B(n15324), .Z(n15061) );
  NAND U14983 ( .A(n15325), .B(n15326), .Z(n15324) );
  NANDN U14984 ( .A(n15327), .B(n15328), .Z(n15323) );
  OR U14985 ( .A(n15325), .B(n15326), .Z(n15328) );
  ANDN U14986 ( .B(\stack[1][20] ), .A(n5734), .Z(n15060) );
  XNOR U14987 ( .A(n15066), .B(n15329), .Z(n15059) );
  XNOR U14988 ( .A(n15067), .B(n15068), .Z(n15329) );
  AND U14989 ( .A(n15330), .B(n15331), .Z(n15068) );
  NANDN U14990 ( .A(n15332), .B(n15333), .Z(n15331) );
  NANDN U14991 ( .A(n15334), .B(n15335), .Z(n15330) );
  NANDN U14992 ( .A(n15333), .B(n15332), .Z(n15335) );
  ANDN U14993 ( .B(\stack[1][21] ), .A(n5710), .Z(n15067) );
  XNOR U14994 ( .A(n15073), .B(n15336), .Z(n15066) );
  XNOR U14995 ( .A(n15074), .B(n15075), .Z(n15336) );
  AND U14996 ( .A(n15337), .B(n15338), .Z(n15075) );
  NAND U14997 ( .A(n15339), .B(n15340), .Z(n15338) );
  NANDN U14998 ( .A(n15341), .B(n15342), .Z(n15337) );
  OR U14999 ( .A(n15339), .B(n15340), .Z(n15342) );
  ANDN U15000 ( .B(\stack[1][22] ), .A(n5686), .Z(n15074) );
  XNOR U15001 ( .A(n15080), .B(n15343), .Z(n15073) );
  XNOR U15002 ( .A(n15081), .B(n15082), .Z(n15343) );
  AND U15003 ( .A(n15344), .B(n15345), .Z(n15082) );
  NANDN U15004 ( .A(n15346), .B(n15347), .Z(n15345) );
  NANDN U15005 ( .A(n15348), .B(n15349), .Z(n15344) );
  NANDN U15006 ( .A(n15347), .B(n15346), .Z(n15349) );
  ANDN U15007 ( .B(\stack[1][23] ), .A(n5662), .Z(n15081) );
  XNOR U15008 ( .A(n15087), .B(n15350), .Z(n15080) );
  XNOR U15009 ( .A(n15088), .B(n15089), .Z(n15350) );
  AND U15010 ( .A(n15351), .B(n15352), .Z(n15089) );
  NAND U15011 ( .A(n15353), .B(n15354), .Z(n15352) );
  NANDN U15012 ( .A(n15355), .B(n15356), .Z(n15351) );
  OR U15013 ( .A(n15353), .B(n15354), .Z(n15356) );
  ANDN U15014 ( .B(\stack[1][24] ), .A(n5638), .Z(n15088) );
  XNOR U15015 ( .A(n15094), .B(n15357), .Z(n15087) );
  XNOR U15016 ( .A(n15095), .B(n15096), .Z(n15357) );
  AND U15017 ( .A(n15358), .B(n15359), .Z(n15096) );
  NANDN U15018 ( .A(n15360), .B(n15361), .Z(n15359) );
  NANDN U15019 ( .A(n15362), .B(n15363), .Z(n15358) );
  NANDN U15020 ( .A(n15361), .B(n15360), .Z(n15363) );
  ANDN U15021 ( .B(\stack[1][25] ), .A(n5614), .Z(n15095) );
  XNOR U15022 ( .A(n15101), .B(n15364), .Z(n15094) );
  XNOR U15023 ( .A(n15102), .B(n15103), .Z(n15364) );
  AND U15024 ( .A(n15365), .B(n15366), .Z(n15103) );
  NAND U15025 ( .A(n15367), .B(n15368), .Z(n15366) );
  NANDN U15026 ( .A(n15369), .B(n15370), .Z(n15365) );
  OR U15027 ( .A(n15367), .B(n15368), .Z(n15370) );
  ANDN U15028 ( .B(\stack[1][26] ), .A(n5590), .Z(n15102) );
  XNOR U15029 ( .A(n15108), .B(n15371), .Z(n15101) );
  XNOR U15030 ( .A(n15109), .B(n15110), .Z(n15371) );
  AND U15031 ( .A(n15372), .B(n15373), .Z(n15110) );
  NANDN U15032 ( .A(n15374), .B(n15375), .Z(n15373) );
  NANDN U15033 ( .A(n15376), .B(n15377), .Z(n15372) );
  NANDN U15034 ( .A(n15375), .B(n15374), .Z(n15377) );
  ANDN U15035 ( .B(\stack[1][27] ), .A(n5566), .Z(n15109) );
  XNOR U15036 ( .A(n15115), .B(n15378), .Z(n15108) );
  XNOR U15037 ( .A(n15116), .B(n15117), .Z(n15378) );
  AND U15038 ( .A(n15379), .B(n15380), .Z(n15117) );
  NAND U15039 ( .A(n15381), .B(n15382), .Z(n15380) );
  NANDN U15040 ( .A(n15383), .B(n15384), .Z(n15379) );
  OR U15041 ( .A(n15381), .B(n15382), .Z(n15384) );
  ANDN U15042 ( .B(\stack[1][28] ), .A(n5542), .Z(n15116) );
  XNOR U15043 ( .A(n15122), .B(n15385), .Z(n15115) );
  XNOR U15044 ( .A(n15123), .B(n15124), .Z(n15385) );
  AND U15045 ( .A(n15386), .B(n15387), .Z(n15124) );
  NANDN U15046 ( .A(n15388), .B(n15389), .Z(n15387) );
  NANDN U15047 ( .A(n15390), .B(n15391), .Z(n15386) );
  NANDN U15048 ( .A(n15389), .B(n15388), .Z(n15391) );
  ANDN U15049 ( .B(\stack[1][29] ), .A(n5518), .Z(n15123) );
  XNOR U15050 ( .A(n15129), .B(n15392), .Z(n15122) );
  XNOR U15051 ( .A(n15130), .B(n15131), .Z(n15392) );
  AND U15052 ( .A(n15393), .B(n15394), .Z(n15131) );
  NAND U15053 ( .A(n15395), .B(n15396), .Z(n15394) );
  NANDN U15054 ( .A(n15397), .B(n15398), .Z(n15393) );
  OR U15055 ( .A(n15395), .B(n15396), .Z(n15398) );
  ANDN U15056 ( .B(\stack[1][30] ), .A(n5494), .Z(n15130) );
  XNOR U15057 ( .A(n15136), .B(n15399), .Z(n15129) );
  XNOR U15058 ( .A(n15137), .B(n15138), .Z(n15399) );
  AND U15059 ( .A(n15400), .B(n15401), .Z(n15138) );
  NANDN U15060 ( .A(n15402), .B(n15403), .Z(n15401) );
  NANDN U15061 ( .A(n15404), .B(n15405), .Z(n15400) );
  NANDN U15062 ( .A(n15403), .B(n15402), .Z(n15405) );
  ANDN U15063 ( .B(\stack[1][31] ), .A(n5470), .Z(n15137) );
  XNOR U15064 ( .A(n15143), .B(n15406), .Z(n15136) );
  XNOR U15065 ( .A(n15144), .B(n15145), .Z(n15406) );
  AND U15066 ( .A(n15407), .B(n15408), .Z(n15145) );
  NAND U15067 ( .A(n15409), .B(n15410), .Z(n15408) );
  NANDN U15068 ( .A(n15411), .B(n15412), .Z(n15407) );
  OR U15069 ( .A(n15409), .B(n15410), .Z(n15412) );
  ANDN U15070 ( .B(\stack[1][32] ), .A(n5446), .Z(n15144) );
  XNOR U15071 ( .A(n15150), .B(n15413), .Z(n15143) );
  XNOR U15072 ( .A(n15151), .B(n15152), .Z(n15413) );
  AND U15073 ( .A(n15414), .B(n15415), .Z(n15152) );
  NANDN U15074 ( .A(n15416), .B(n15417), .Z(n15415) );
  NANDN U15075 ( .A(n15418), .B(n15419), .Z(n15414) );
  NANDN U15076 ( .A(n15417), .B(n15416), .Z(n15419) );
  ANDN U15077 ( .B(\stack[1][33] ), .A(n5422), .Z(n15151) );
  XNOR U15078 ( .A(n15157), .B(n15420), .Z(n15150) );
  XNOR U15079 ( .A(n15158), .B(n15159), .Z(n15420) );
  AND U15080 ( .A(n15421), .B(n15422), .Z(n15159) );
  NAND U15081 ( .A(n15423), .B(n15424), .Z(n15422) );
  NANDN U15082 ( .A(n15425), .B(n15426), .Z(n15421) );
  OR U15083 ( .A(n15423), .B(n15424), .Z(n15426) );
  ANDN U15084 ( .B(\stack[1][34] ), .A(n5398), .Z(n15158) );
  XNOR U15085 ( .A(n15164), .B(n15427), .Z(n15157) );
  XNOR U15086 ( .A(n15165), .B(n15166), .Z(n15427) );
  AND U15087 ( .A(n15428), .B(n15429), .Z(n15166) );
  NANDN U15088 ( .A(n15430), .B(n15431), .Z(n15429) );
  NANDN U15089 ( .A(n15432), .B(n15433), .Z(n15428) );
  NANDN U15090 ( .A(n15431), .B(n15430), .Z(n15433) );
  ANDN U15091 ( .B(\stack[1][35] ), .A(n5374), .Z(n15165) );
  XNOR U15092 ( .A(n15171), .B(n15434), .Z(n15164) );
  XNOR U15093 ( .A(n15172), .B(n15173), .Z(n15434) );
  AND U15094 ( .A(n15435), .B(n15436), .Z(n15173) );
  NAND U15095 ( .A(n15437), .B(n15438), .Z(n15436) );
  NANDN U15096 ( .A(n15439), .B(n15440), .Z(n15435) );
  OR U15097 ( .A(n15437), .B(n15438), .Z(n15440) );
  ANDN U15098 ( .B(\stack[1][36] ), .A(n5350), .Z(n15172) );
  XNOR U15099 ( .A(n15179), .B(n15441), .Z(n15171) );
  XOR U15100 ( .A(n15180), .B(n15181), .Z(n15441) );
  NAND U15101 ( .A(n15442), .B(n15443), .Z(n15181) );
  NANDN U15102 ( .A(n15444), .B(n15445), .Z(n15443) );
  OR U15103 ( .A(n15446), .B(n15447), .Z(n15445) );
  AND U15104 ( .A(\stack[0][7] ), .B(\stack[1][37] ), .Z(n15180) );
  XNOR U15105 ( .A(n15186), .B(n15448), .Z(n15179) );
  XNOR U15106 ( .A(n15185), .B(n15188), .Z(n15448) );
  AND U15107 ( .A(\stack[0][6] ), .B(\stack[1][38] ), .Z(n15188) );
  AND U15108 ( .A(n15449), .B(n15450), .Z(n15185) );
  NAND U15109 ( .A(n15451), .B(n15452), .Z(n15450) );
  OR U15110 ( .A(n15453), .B(n15454), .Z(n15451) );
  XNOR U15111 ( .A(n15192), .B(n15455), .Z(n15186) );
  XNOR U15112 ( .A(n15193), .B(n15194), .Z(n15455) );
  AND U15113 ( .A(n15456), .B(n15457), .Z(n15194) );
  NANDN U15114 ( .A(n15458), .B(n15459), .Z(n15457) );
  NANDN U15115 ( .A(n15460), .B(n15461), .Z(n15456) );
  NANDN U15116 ( .A(n15459), .B(n15458), .Z(n15461) );
  ANDN U15117 ( .B(\stack[1][39] ), .A(n5278), .Z(n15193) );
  XNOR U15118 ( .A(n15199), .B(n15462), .Z(n15192) );
  XNOR U15119 ( .A(n15200), .B(n15201), .Z(n15462) );
  AND U15120 ( .A(n15463), .B(n15464), .Z(n15201) );
  NAND U15121 ( .A(n15465), .B(n15466), .Z(n15464) );
  NANDN U15122 ( .A(n15467), .B(n15468), .Z(n15463) );
  OR U15123 ( .A(n15465), .B(n15466), .Z(n15468) );
  ANDN U15124 ( .B(\stack[1][40] ), .A(n5254), .Z(n15200) );
  XNOR U15125 ( .A(n15206), .B(n15469), .Z(n15199) );
  XNOR U15126 ( .A(n15207), .B(n15208), .Z(n15469) );
  AND U15127 ( .A(n15470), .B(n15471), .Z(n15208) );
  NAND U15128 ( .A(n15472), .B(n15473), .Z(n15471) );
  NAND U15129 ( .A(n15474), .B(n15475), .Z(n15470) );
  OR U15130 ( .A(n15472), .B(n15473), .Z(n15474) );
  ANDN U15131 ( .B(\stack[1][41] ), .A(n5230), .Z(n15207) );
  XNOR U15132 ( .A(n15213), .B(n15476), .Z(n15206) );
  XNOR U15133 ( .A(n15214), .B(n15216), .Z(n15476) );
  ANDN U15134 ( .B(n15477), .A(n15478), .Z(n15216) );
  ANDN U15135 ( .B(\stack[0][0] ), .A(n6204), .Z(n15477) );
  ANDN U15136 ( .B(\stack[1][42] ), .A(n5206), .Z(n15214) );
  XOR U15137 ( .A(n15219), .B(n15479), .Z(n15213) );
  NANDN U15138 ( .A(n5160), .B(\stack[1][44] ), .Z(n15479) );
  NANDN U15139 ( .A(n6204), .B(\stack[0][1] ), .Z(n15219) );
  ANDN U15140 ( .B(\stack[0][39] ), .A(n5292), .Z(n9090) );
  AND U15141 ( .A(n15480), .B(n15481), .Z(n9091) );
  NANDN U15142 ( .A(n9098), .B(n15482), .Z(n15480) );
  NANDN U15143 ( .A(n9097), .B(n9095), .Z(n15482) );
  XNOR U15144 ( .A(n15227), .B(n15483), .Z(n9095) );
  XNOR U15145 ( .A(n15228), .B(n15229), .Z(n15483) );
  AND U15146 ( .A(n15484), .B(n15485), .Z(n15229) );
  NANDN U15147 ( .A(n15486), .B(n15487), .Z(n15485) );
  NANDN U15148 ( .A(n15488), .B(n15489), .Z(n15484) );
  NANDN U15149 ( .A(n15487), .B(n15486), .Z(n15489) );
  ANDN U15150 ( .B(\stack[0][37] ), .A(n5316), .Z(n15228) );
  XNOR U15151 ( .A(n15234), .B(n15490), .Z(n15227) );
  XNOR U15152 ( .A(n15235), .B(n15236), .Z(n15490) );
  AND U15153 ( .A(n15491), .B(n15492), .Z(n15236) );
  NAND U15154 ( .A(n15493), .B(n15494), .Z(n15492) );
  NANDN U15155 ( .A(n15495), .B(n15496), .Z(n15491) );
  OR U15156 ( .A(n15493), .B(n15494), .Z(n15496) );
  ANDN U15157 ( .B(\stack[0][36] ), .A(n5340), .Z(n15235) );
  XNOR U15158 ( .A(n15241), .B(n15497), .Z(n15234) );
  XNOR U15159 ( .A(n15242), .B(n15243), .Z(n15497) );
  AND U15160 ( .A(n15498), .B(n15499), .Z(n15243) );
  NANDN U15161 ( .A(n15500), .B(n15501), .Z(n15499) );
  NANDN U15162 ( .A(n15502), .B(n15503), .Z(n15498) );
  NANDN U15163 ( .A(n15501), .B(n15500), .Z(n15503) );
  ANDN U15164 ( .B(\stack[0][35] ), .A(n5364), .Z(n15242) );
  XNOR U15165 ( .A(n15248), .B(n15504), .Z(n15241) );
  XNOR U15166 ( .A(n15249), .B(n15250), .Z(n15504) );
  AND U15167 ( .A(n15505), .B(n15506), .Z(n15250) );
  NAND U15168 ( .A(n15507), .B(n15508), .Z(n15506) );
  NANDN U15169 ( .A(n15509), .B(n15510), .Z(n15505) );
  OR U15170 ( .A(n15507), .B(n15508), .Z(n15510) );
  ANDN U15171 ( .B(\stack[0][34] ), .A(n5387), .Z(n15249) );
  XNOR U15172 ( .A(n15255), .B(n15511), .Z(n15248) );
  XNOR U15173 ( .A(n15256), .B(n15257), .Z(n15511) );
  AND U15174 ( .A(n15512), .B(n15513), .Z(n15257) );
  NANDN U15175 ( .A(n15514), .B(n15515), .Z(n15513) );
  NANDN U15176 ( .A(n15516), .B(n15517), .Z(n15512) );
  NANDN U15177 ( .A(n15515), .B(n15514), .Z(n15517) );
  ANDN U15178 ( .B(\stack[1][10] ), .A(n5950), .Z(n15256) );
  XNOR U15179 ( .A(n15262), .B(n15518), .Z(n15255) );
  XNOR U15180 ( .A(n15263), .B(n15264), .Z(n15518) );
  AND U15181 ( .A(n15519), .B(n15520), .Z(n15264) );
  NAND U15182 ( .A(n15521), .B(n15522), .Z(n15520) );
  NANDN U15183 ( .A(n15523), .B(n15524), .Z(n15519) );
  OR U15184 ( .A(n15521), .B(n15522), .Z(n15524) );
  ANDN U15185 ( .B(\stack[1][11] ), .A(n5926), .Z(n15263) );
  XNOR U15186 ( .A(n15269), .B(n15525), .Z(n15262) );
  XNOR U15187 ( .A(n15270), .B(n15271), .Z(n15525) );
  AND U15188 ( .A(n15526), .B(n15527), .Z(n15271) );
  NANDN U15189 ( .A(n15528), .B(n15529), .Z(n15527) );
  NANDN U15190 ( .A(n15530), .B(n15531), .Z(n15526) );
  NANDN U15191 ( .A(n15529), .B(n15528), .Z(n15531) );
  ANDN U15192 ( .B(\stack[1][12] ), .A(n5902), .Z(n15270) );
  XNOR U15193 ( .A(n15276), .B(n15532), .Z(n15269) );
  XNOR U15194 ( .A(n15277), .B(n15278), .Z(n15532) );
  AND U15195 ( .A(n15533), .B(n15534), .Z(n15278) );
  NAND U15196 ( .A(n15535), .B(n15536), .Z(n15534) );
  NANDN U15197 ( .A(n15537), .B(n15538), .Z(n15533) );
  OR U15198 ( .A(n15535), .B(n15536), .Z(n15538) );
  ANDN U15199 ( .B(\stack[1][13] ), .A(n5878), .Z(n15277) );
  XNOR U15200 ( .A(n15283), .B(n15539), .Z(n15276) );
  XNOR U15201 ( .A(n15284), .B(n15285), .Z(n15539) );
  AND U15202 ( .A(n15540), .B(n15541), .Z(n15285) );
  NANDN U15203 ( .A(n15542), .B(n15543), .Z(n15541) );
  NANDN U15204 ( .A(n15544), .B(n15545), .Z(n15540) );
  NANDN U15205 ( .A(n15543), .B(n15542), .Z(n15545) );
  ANDN U15206 ( .B(\stack[1][14] ), .A(n5854), .Z(n15284) );
  XNOR U15207 ( .A(n15290), .B(n15546), .Z(n15283) );
  XNOR U15208 ( .A(n15291), .B(n15292), .Z(n15546) );
  AND U15209 ( .A(n15547), .B(n15548), .Z(n15292) );
  NAND U15210 ( .A(n15549), .B(n15550), .Z(n15548) );
  NANDN U15211 ( .A(n15551), .B(n15552), .Z(n15547) );
  OR U15212 ( .A(n15549), .B(n15550), .Z(n15552) );
  ANDN U15213 ( .B(\stack[1][15] ), .A(n5830), .Z(n15291) );
  XNOR U15214 ( .A(n15297), .B(n15553), .Z(n15290) );
  XNOR U15215 ( .A(n15298), .B(n15299), .Z(n15553) );
  AND U15216 ( .A(n15554), .B(n15555), .Z(n15299) );
  NANDN U15217 ( .A(n15556), .B(n15557), .Z(n15555) );
  NANDN U15218 ( .A(n15558), .B(n15559), .Z(n15554) );
  NANDN U15219 ( .A(n15557), .B(n15556), .Z(n15559) );
  ANDN U15220 ( .B(\stack[1][16] ), .A(n5806), .Z(n15298) );
  XNOR U15221 ( .A(n15304), .B(n15560), .Z(n15297) );
  XNOR U15222 ( .A(n15305), .B(n15306), .Z(n15560) );
  AND U15223 ( .A(n15561), .B(n15562), .Z(n15306) );
  NAND U15224 ( .A(n15563), .B(n15564), .Z(n15562) );
  NANDN U15225 ( .A(n15565), .B(n15566), .Z(n15561) );
  OR U15226 ( .A(n15563), .B(n15564), .Z(n15566) );
  ANDN U15227 ( .B(\stack[1][17] ), .A(n5782), .Z(n15305) );
  XNOR U15228 ( .A(n15311), .B(n15567), .Z(n15304) );
  XNOR U15229 ( .A(n15312), .B(n15313), .Z(n15567) );
  AND U15230 ( .A(n15568), .B(n15569), .Z(n15313) );
  NANDN U15231 ( .A(n15570), .B(n15571), .Z(n15569) );
  NANDN U15232 ( .A(n15572), .B(n15573), .Z(n15568) );
  NANDN U15233 ( .A(n15571), .B(n15570), .Z(n15573) );
  ANDN U15234 ( .B(\stack[1][18] ), .A(n5758), .Z(n15312) );
  XNOR U15235 ( .A(n15318), .B(n15574), .Z(n15311) );
  XNOR U15236 ( .A(n15319), .B(n15320), .Z(n15574) );
  AND U15237 ( .A(n15575), .B(n15576), .Z(n15320) );
  NAND U15238 ( .A(n15577), .B(n15578), .Z(n15576) );
  NANDN U15239 ( .A(n15579), .B(n15580), .Z(n15575) );
  OR U15240 ( .A(n15577), .B(n15578), .Z(n15580) );
  ANDN U15241 ( .B(\stack[1][19] ), .A(n5734), .Z(n15319) );
  XNOR U15242 ( .A(n15325), .B(n15581), .Z(n15318) );
  XNOR U15243 ( .A(n15326), .B(n15327), .Z(n15581) );
  AND U15244 ( .A(n15582), .B(n15583), .Z(n15327) );
  NANDN U15245 ( .A(n15584), .B(n15585), .Z(n15583) );
  NANDN U15246 ( .A(n15586), .B(n15587), .Z(n15582) );
  NANDN U15247 ( .A(n15585), .B(n15584), .Z(n15587) );
  ANDN U15248 ( .B(\stack[1][20] ), .A(n5710), .Z(n15326) );
  XNOR U15249 ( .A(n15332), .B(n15588), .Z(n15325) );
  XNOR U15250 ( .A(n15333), .B(n15334), .Z(n15588) );
  AND U15251 ( .A(n15589), .B(n15590), .Z(n15334) );
  NAND U15252 ( .A(n15591), .B(n15592), .Z(n15590) );
  NANDN U15253 ( .A(n15593), .B(n15594), .Z(n15589) );
  OR U15254 ( .A(n15591), .B(n15592), .Z(n15594) );
  ANDN U15255 ( .B(\stack[1][21] ), .A(n5686), .Z(n15333) );
  XNOR U15256 ( .A(n15339), .B(n15595), .Z(n15332) );
  XNOR U15257 ( .A(n15340), .B(n15341), .Z(n15595) );
  AND U15258 ( .A(n15596), .B(n15597), .Z(n15341) );
  NANDN U15259 ( .A(n15598), .B(n15599), .Z(n15597) );
  NANDN U15260 ( .A(n15600), .B(n15601), .Z(n15596) );
  NANDN U15261 ( .A(n15599), .B(n15598), .Z(n15601) );
  ANDN U15262 ( .B(\stack[1][22] ), .A(n5662), .Z(n15340) );
  XNOR U15263 ( .A(n15346), .B(n15602), .Z(n15339) );
  XNOR U15264 ( .A(n15347), .B(n15348), .Z(n15602) );
  AND U15265 ( .A(n15603), .B(n15604), .Z(n15348) );
  NAND U15266 ( .A(n15605), .B(n15606), .Z(n15604) );
  NANDN U15267 ( .A(n15607), .B(n15608), .Z(n15603) );
  OR U15268 ( .A(n15605), .B(n15606), .Z(n15608) );
  ANDN U15269 ( .B(\stack[1][23] ), .A(n5638), .Z(n15347) );
  XNOR U15270 ( .A(n15353), .B(n15609), .Z(n15346) );
  XNOR U15271 ( .A(n15354), .B(n15355), .Z(n15609) );
  AND U15272 ( .A(n15610), .B(n15611), .Z(n15355) );
  NANDN U15273 ( .A(n15612), .B(n15613), .Z(n15611) );
  NANDN U15274 ( .A(n15614), .B(n15615), .Z(n15610) );
  NANDN U15275 ( .A(n15613), .B(n15612), .Z(n15615) );
  ANDN U15276 ( .B(\stack[1][24] ), .A(n5614), .Z(n15354) );
  XNOR U15277 ( .A(n15360), .B(n15616), .Z(n15353) );
  XNOR U15278 ( .A(n15361), .B(n15362), .Z(n15616) );
  AND U15279 ( .A(n15617), .B(n15618), .Z(n15362) );
  NAND U15280 ( .A(n15619), .B(n15620), .Z(n15618) );
  NANDN U15281 ( .A(n15621), .B(n15622), .Z(n15617) );
  OR U15282 ( .A(n15619), .B(n15620), .Z(n15622) );
  ANDN U15283 ( .B(\stack[1][25] ), .A(n5590), .Z(n15361) );
  XNOR U15284 ( .A(n15367), .B(n15623), .Z(n15360) );
  XNOR U15285 ( .A(n15368), .B(n15369), .Z(n15623) );
  AND U15286 ( .A(n15624), .B(n15625), .Z(n15369) );
  NANDN U15287 ( .A(n15626), .B(n15627), .Z(n15625) );
  NANDN U15288 ( .A(n15628), .B(n15629), .Z(n15624) );
  NANDN U15289 ( .A(n15627), .B(n15626), .Z(n15629) );
  ANDN U15290 ( .B(\stack[1][26] ), .A(n5566), .Z(n15368) );
  XNOR U15291 ( .A(n15374), .B(n15630), .Z(n15367) );
  XNOR U15292 ( .A(n15375), .B(n15376), .Z(n15630) );
  AND U15293 ( .A(n15631), .B(n15632), .Z(n15376) );
  NAND U15294 ( .A(n15633), .B(n15634), .Z(n15632) );
  NANDN U15295 ( .A(n15635), .B(n15636), .Z(n15631) );
  OR U15296 ( .A(n15633), .B(n15634), .Z(n15636) );
  ANDN U15297 ( .B(\stack[1][27] ), .A(n5542), .Z(n15375) );
  XNOR U15298 ( .A(n15381), .B(n15637), .Z(n15374) );
  XNOR U15299 ( .A(n15382), .B(n15383), .Z(n15637) );
  AND U15300 ( .A(n15638), .B(n15639), .Z(n15383) );
  NANDN U15301 ( .A(n15640), .B(n15641), .Z(n15639) );
  NANDN U15302 ( .A(n15642), .B(n15643), .Z(n15638) );
  NANDN U15303 ( .A(n15641), .B(n15640), .Z(n15643) );
  ANDN U15304 ( .B(\stack[1][28] ), .A(n5518), .Z(n15382) );
  XNOR U15305 ( .A(n15388), .B(n15644), .Z(n15381) );
  XNOR U15306 ( .A(n15389), .B(n15390), .Z(n15644) );
  AND U15307 ( .A(n15645), .B(n15646), .Z(n15390) );
  NAND U15308 ( .A(n15647), .B(n15648), .Z(n15646) );
  NANDN U15309 ( .A(n15649), .B(n15650), .Z(n15645) );
  OR U15310 ( .A(n15647), .B(n15648), .Z(n15650) );
  ANDN U15311 ( .B(\stack[1][29] ), .A(n5494), .Z(n15389) );
  XNOR U15312 ( .A(n15395), .B(n15651), .Z(n15388) );
  XNOR U15313 ( .A(n15396), .B(n15397), .Z(n15651) );
  AND U15314 ( .A(n15652), .B(n15653), .Z(n15397) );
  NANDN U15315 ( .A(n15654), .B(n15655), .Z(n15653) );
  NANDN U15316 ( .A(n15656), .B(n15657), .Z(n15652) );
  NANDN U15317 ( .A(n15655), .B(n15654), .Z(n15657) );
  ANDN U15318 ( .B(\stack[1][30] ), .A(n5470), .Z(n15396) );
  XNOR U15319 ( .A(n15402), .B(n15658), .Z(n15395) );
  XNOR U15320 ( .A(n15403), .B(n15404), .Z(n15658) );
  AND U15321 ( .A(n15659), .B(n15660), .Z(n15404) );
  NAND U15322 ( .A(n15661), .B(n15662), .Z(n15660) );
  NANDN U15323 ( .A(n15663), .B(n15664), .Z(n15659) );
  OR U15324 ( .A(n15661), .B(n15662), .Z(n15664) );
  ANDN U15325 ( .B(\stack[1][31] ), .A(n5446), .Z(n15403) );
  XNOR U15326 ( .A(n15409), .B(n15665), .Z(n15402) );
  XNOR U15327 ( .A(n15410), .B(n15411), .Z(n15665) );
  AND U15328 ( .A(n15666), .B(n15667), .Z(n15411) );
  NANDN U15329 ( .A(n15668), .B(n15669), .Z(n15667) );
  NANDN U15330 ( .A(n15670), .B(n15671), .Z(n15666) );
  NANDN U15331 ( .A(n15669), .B(n15668), .Z(n15671) );
  ANDN U15332 ( .B(\stack[1][32] ), .A(n5422), .Z(n15410) );
  XNOR U15333 ( .A(n15416), .B(n15672), .Z(n15409) );
  XNOR U15334 ( .A(n15417), .B(n15418), .Z(n15672) );
  AND U15335 ( .A(n15673), .B(n15674), .Z(n15418) );
  NAND U15336 ( .A(n15675), .B(n15676), .Z(n15674) );
  NANDN U15337 ( .A(n15677), .B(n15678), .Z(n15673) );
  OR U15338 ( .A(n15675), .B(n15676), .Z(n15678) );
  ANDN U15339 ( .B(\stack[1][33] ), .A(n5398), .Z(n15417) );
  XNOR U15340 ( .A(n15423), .B(n15679), .Z(n15416) );
  XNOR U15341 ( .A(n15424), .B(n15425), .Z(n15679) );
  AND U15342 ( .A(n15680), .B(n15681), .Z(n15425) );
  NANDN U15343 ( .A(n15682), .B(n15683), .Z(n15681) );
  NANDN U15344 ( .A(n15684), .B(n15685), .Z(n15680) );
  NANDN U15345 ( .A(n15683), .B(n15682), .Z(n15685) );
  ANDN U15346 ( .B(\stack[1][34] ), .A(n5374), .Z(n15424) );
  XNOR U15347 ( .A(n15430), .B(n15686), .Z(n15423) );
  XNOR U15348 ( .A(n15431), .B(n15432), .Z(n15686) );
  AND U15349 ( .A(n15687), .B(n15688), .Z(n15432) );
  NAND U15350 ( .A(n15689), .B(n15690), .Z(n15688) );
  NANDN U15351 ( .A(n15691), .B(n15692), .Z(n15687) );
  OR U15352 ( .A(n15689), .B(n15690), .Z(n15692) );
  ANDN U15353 ( .B(\stack[1][35] ), .A(n5350), .Z(n15431) );
  XNOR U15354 ( .A(n15437), .B(n15693), .Z(n15430) );
  XNOR U15355 ( .A(n15438), .B(n15439), .Z(n15693) );
  AND U15356 ( .A(n15694), .B(n15695), .Z(n15439) );
  NANDN U15357 ( .A(n15696), .B(n15697), .Z(n15695) );
  NANDN U15358 ( .A(n15698), .B(n15699), .Z(n15694) );
  NANDN U15359 ( .A(n15697), .B(n15696), .Z(n15699) );
  ANDN U15360 ( .B(\stack[1][36] ), .A(n5326), .Z(n15438) );
  XNOR U15361 ( .A(n15444), .B(n15700), .Z(n15437) );
  XOR U15362 ( .A(n15446), .B(n15447), .Z(n15700) );
  NAND U15363 ( .A(n15701), .B(n15702), .Z(n15447) );
  NAND U15364 ( .A(n15703), .B(n15704), .Z(n15702) );
  OR U15365 ( .A(n15705), .B(n15706), .Z(n15703) );
  AND U15366 ( .A(\stack[0][6] ), .B(\stack[1][37] ), .Z(n15446) );
  XNOR U15367 ( .A(n15453), .B(n15707), .Z(n15444) );
  XOR U15368 ( .A(n15454), .B(n15452), .Z(n15707) );
  AND U15369 ( .A(\stack[0][5] ), .B(\stack[1][38] ), .Z(n15452) );
  NAND U15370 ( .A(n15708), .B(n15709), .Z(n15454) );
  OR U15371 ( .A(n15710), .B(n15711), .Z(n15709) );
  NAND U15372 ( .A(n15712), .B(n15713), .Z(n15708) );
  NAND U15373 ( .A(n15711), .B(n15710), .Z(n15712) );
  XNOR U15374 ( .A(n15458), .B(n15714), .Z(n15453) );
  XNOR U15375 ( .A(n15459), .B(n15460), .Z(n15714) );
  AND U15376 ( .A(n15715), .B(n15716), .Z(n15460) );
  NAND U15377 ( .A(n15717), .B(n15718), .Z(n15716) );
  NANDN U15378 ( .A(n15719), .B(n15720), .Z(n15715) );
  OR U15379 ( .A(n15717), .B(n15718), .Z(n15720) );
  ANDN U15380 ( .B(\stack[1][39] ), .A(n5254), .Z(n15459) );
  XNOR U15381 ( .A(n15465), .B(n15721), .Z(n15458) );
  XNOR U15382 ( .A(n15466), .B(n15467), .Z(n15721) );
  AND U15383 ( .A(n15722), .B(n15723), .Z(n15467) );
  NAND U15384 ( .A(n15724), .B(n15725), .Z(n15723) );
  NAND U15385 ( .A(n15726), .B(n15727), .Z(n15722) );
  OR U15386 ( .A(n15724), .B(n15725), .Z(n15726) );
  ANDN U15387 ( .B(\stack[1][40] ), .A(n5230), .Z(n15466) );
  XNOR U15388 ( .A(n15472), .B(n15728), .Z(n15465) );
  XNOR U15389 ( .A(n15473), .B(n15475), .Z(n15728) );
  ANDN U15390 ( .B(n15729), .A(n15730), .Z(n15475) );
  ANDN U15391 ( .B(\stack[0][0] ), .A(n6180), .Z(n15729) );
  ANDN U15392 ( .B(\stack[1][41] ), .A(n5206), .Z(n15473) );
  XOR U15393 ( .A(n15478), .B(n15731), .Z(n15472) );
  NANDN U15394 ( .A(n5160), .B(\stack[1][43] ), .Z(n15731) );
  NANDN U15395 ( .A(n6180), .B(\stack[0][1] ), .Z(n15478) );
  ANDN U15396 ( .B(\stack[1][5] ), .A(n6070), .Z(n9097) );
  AND U15397 ( .A(n15732), .B(n15733), .Z(n9098) );
  NANDN U15398 ( .A(n9102), .B(n9104), .Z(n15733) );
  NANDN U15399 ( .A(n9105), .B(n15734), .Z(n15732) );
  NANDN U15400 ( .A(n9104), .B(n9102), .Z(n15734) );
  XOR U15401 ( .A(n15486), .B(n15735), .Z(n9102) );
  XNOR U15402 ( .A(n15487), .B(n15488), .Z(n15735) );
  AND U15403 ( .A(n15736), .B(n15737), .Z(n15488) );
  NAND U15404 ( .A(n15738), .B(n15739), .Z(n15737) );
  NANDN U15405 ( .A(n15740), .B(n15741), .Z(n15736) );
  OR U15406 ( .A(n15738), .B(n15739), .Z(n15741) );
  ANDN U15407 ( .B(\stack[0][36] ), .A(n5316), .Z(n15487) );
  XNOR U15408 ( .A(n15493), .B(n15742), .Z(n15486) );
  XNOR U15409 ( .A(n15494), .B(n15495), .Z(n15742) );
  AND U15410 ( .A(n15743), .B(n15744), .Z(n15495) );
  NANDN U15411 ( .A(n15745), .B(n15746), .Z(n15744) );
  NANDN U15412 ( .A(n15747), .B(n15748), .Z(n15743) );
  NANDN U15413 ( .A(n15746), .B(n15745), .Z(n15748) );
  ANDN U15414 ( .B(\stack[0][35] ), .A(n5340), .Z(n15494) );
  XNOR U15415 ( .A(n15500), .B(n15749), .Z(n15493) );
  XNOR U15416 ( .A(n15501), .B(n15502), .Z(n15749) );
  AND U15417 ( .A(n15750), .B(n15751), .Z(n15502) );
  NAND U15418 ( .A(n15752), .B(n15753), .Z(n15751) );
  NANDN U15419 ( .A(n15754), .B(n15755), .Z(n15750) );
  OR U15420 ( .A(n15752), .B(n15753), .Z(n15755) );
  ANDN U15421 ( .B(\stack[0][34] ), .A(n5364), .Z(n15501) );
  XNOR U15422 ( .A(n15507), .B(n15756), .Z(n15500) );
  XNOR U15423 ( .A(n15508), .B(n15509), .Z(n15756) );
  AND U15424 ( .A(n15757), .B(n15758), .Z(n15509) );
  NANDN U15425 ( .A(n15759), .B(n15760), .Z(n15758) );
  NANDN U15426 ( .A(n15761), .B(n15762), .Z(n15757) );
  NANDN U15427 ( .A(n15760), .B(n15759), .Z(n15762) );
  ANDN U15428 ( .B(\stack[0][33] ), .A(n5387), .Z(n15508) );
  XNOR U15429 ( .A(n15514), .B(n15763), .Z(n15507) );
  XNOR U15430 ( .A(n15515), .B(n15516), .Z(n15763) );
  AND U15431 ( .A(n15764), .B(n15765), .Z(n15516) );
  NAND U15432 ( .A(n15766), .B(n15767), .Z(n15765) );
  NANDN U15433 ( .A(n15768), .B(n15769), .Z(n15764) );
  OR U15434 ( .A(n15766), .B(n15767), .Z(n15769) );
  ANDN U15435 ( .B(\stack[1][10] ), .A(n5926), .Z(n15515) );
  XNOR U15436 ( .A(n15521), .B(n15770), .Z(n15514) );
  XNOR U15437 ( .A(n15522), .B(n15523), .Z(n15770) );
  AND U15438 ( .A(n15771), .B(n15772), .Z(n15523) );
  NANDN U15439 ( .A(n15773), .B(n15774), .Z(n15772) );
  NANDN U15440 ( .A(n15775), .B(n15776), .Z(n15771) );
  NANDN U15441 ( .A(n15774), .B(n15773), .Z(n15776) );
  ANDN U15442 ( .B(\stack[1][11] ), .A(n5902), .Z(n15522) );
  XNOR U15443 ( .A(n15528), .B(n15777), .Z(n15521) );
  XNOR U15444 ( .A(n15529), .B(n15530), .Z(n15777) );
  AND U15445 ( .A(n15778), .B(n15779), .Z(n15530) );
  NAND U15446 ( .A(n15780), .B(n15781), .Z(n15779) );
  NANDN U15447 ( .A(n15782), .B(n15783), .Z(n15778) );
  OR U15448 ( .A(n15780), .B(n15781), .Z(n15783) );
  ANDN U15449 ( .B(\stack[1][12] ), .A(n5878), .Z(n15529) );
  XNOR U15450 ( .A(n15535), .B(n15784), .Z(n15528) );
  XNOR U15451 ( .A(n15536), .B(n15537), .Z(n15784) );
  AND U15452 ( .A(n15785), .B(n15786), .Z(n15537) );
  NANDN U15453 ( .A(n15787), .B(n15788), .Z(n15786) );
  NANDN U15454 ( .A(n15789), .B(n15790), .Z(n15785) );
  NANDN U15455 ( .A(n15788), .B(n15787), .Z(n15790) );
  ANDN U15456 ( .B(\stack[1][13] ), .A(n5854), .Z(n15536) );
  XNOR U15457 ( .A(n15542), .B(n15791), .Z(n15535) );
  XNOR U15458 ( .A(n15543), .B(n15544), .Z(n15791) );
  AND U15459 ( .A(n15792), .B(n15793), .Z(n15544) );
  NAND U15460 ( .A(n15794), .B(n15795), .Z(n15793) );
  NANDN U15461 ( .A(n15796), .B(n15797), .Z(n15792) );
  OR U15462 ( .A(n15794), .B(n15795), .Z(n15797) );
  ANDN U15463 ( .B(\stack[1][14] ), .A(n5830), .Z(n15543) );
  XNOR U15464 ( .A(n15549), .B(n15798), .Z(n15542) );
  XNOR U15465 ( .A(n15550), .B(n15551), .Z(n15798) );
  AND U15466 ( .A(n15799), .B(n15800), .Z(n15551) );
  NANDN U15467 ( .A(n15801), .B(n15802), .Z(n15800) );
  NANDN U15468 ( .A(n15803), .B(n15804), .Z(n15799) );
  NANDN U15469 ( .A(n15802), .B(n15801), .Z(n15804) );
  ANDN U15470 ( .B(\stack[1][15] ), .A(n5806), .Z(n15550) );
  XNOR U15471 ( .A(n15556), .B(n15805), .Z(n15549) );
  XNOR U15472 ( .A(n15557), .B(n15558), .Z(n15805) );
  AND U15473 ( .A(n15806), .B(n15807), .Z(n15558) );
  NAND U15474 ( .A(n15808), .B(n15809), .Z(n15807) );
  NANDN U15475 ( .A(n15810), .B(n15811), .Z(n15806) );
  OR U15476 ( .A(n15808), .B(n15809), .Z(n15811) );
  ANDN U15477 ( .B(\stack[1][16] ), .A(n5782), .Z(n15557) );
  XNOR U15478 ( .A(n15563), .B(n15812), .Z(n15556) );
  XNOR U15479 ( .A(n15564), .B(n15565), .Z(n15812) );
  AND U15480 ( .A(n15813), .B(n15814), .Z(n15565) );
  NANDN U15481 ( .A(n15815), .B(n15816), .Z(n15814) );
  NANDN U15482 ( .A(n15817), .B(n15818), .Z(n15813) );
  NANDN U15483 ( .A(n15816), .B(n15815), .Z(n15818) );
  ANDN U15484 ( .B(\stack[1][17] ), .A(n5758), .Z(n15564) );
  XNOR U15485 ( .A(n15570), .B(n15819), .Z(n15563) );
  XNOR U15486 ( .A(n15571), .B(n15572), .Z(n15819) );
  AND U15487 ( .A(n15820), .B(n15821), .Z(n15572) );
  NAND U15488 ( .A(n15822), .B(n15823), .Z(n15821) );
  NANDN U15489 ( .A(n15824), .B(n15825), .Z(n15820) );
  OR U15490 ( .A(n15822), .B(n15823), .Z(n15825) );
  ANDN U15491 ( .B(\stack[1][18] ), .A(n5734), .Z(n15571) );
  XNOR U15492 ( .A(n15577), .B(n15826), .Z(n15570) );
  XNOR U15493 ( .A(n15578), .B(n15579), .Z(n15826) );
  AND U15494 ( .A(n15827), .B(n15828), .Z(n15579) );
  NANDN U15495 ( .A(n15829), .B(n15830), .Z(n15828) );
  NANDN U15496 ( .A(n15831), .B(n15832), .Z(n15827) );
  NANDN U15497 ( .A(n15830), .B(n15829), .Z(n15832) );
  ANDN U15498 ( .B(\stack[1][19] ), .A(n5710), .Z(n15578) );
  XNOR U15499 ( .A(n15584), .B(n15833), .Z(n15577) );
  XNOR U15500 ( .A(n15585), .B(n15586), .Z(n15833) );
  AND U15501 ( .A(n15834), .B(n15835), .Z(n15586) );
  NAND U15502 ( .A(n15836), .B(n15837), .Z(n15835) );
  NANDN U15503 ( .A(n15838), .B(n15839), .Z(n15834) );
  OR U15504 ( .A(n15836), .B(n15837), .Z(n15839) );
  ANDN U15505 ( .B(\stack[1][20] ), .A(n5686), .Z(n15585) );
  XNOR U15506 ( .A(n15591), .B(n15840), .Z(n15584) );
  XNOR U15507 ( .A(n15592), .B(n15593), .Z(n15840) );
  AND U15508 ( .A(n15841), .B(n15842), .Z(n15593) );
  NANDN U15509 ( .A(n15843), .B(n15844), .Z(n15842) );
  NANDN U15510 ( .A(n15845), .B(n15846), .Z(n15841) );
  NANDN U15511 ( .A(n15844), .B(n15843), .Z(n15846) );
  ANDN U15512 ( .B(\stack[1][21] ), .A(n5662), .Z(n15592) );
  XNOR U15513 ( .A(n15598), .B(n15847), .Z(n15591) );
  XNOR U15514 ( .A(n15599), .B(n15600), .Z(n15847) );
  AND U15515 ( .A(n15848), .B(n15849), .Z(n15600) );
  NAND U15516 ( .A(n15850), .B(n15851), .Z(n15849) );
  NANDN U15517 ( .A(n15852), .B(n15853), .Z(n15848) );
  OR U15518 ( .A(n15850), .B(n15851), .Z(n15853) );
  ANDN U15519 ( .B(\stack[1][22] ), .A(n5638), .Z(n15599) );
  XNOR U15520 ( .A(n15605), .B(n15854), .Z(n15598) );
  XNOR U15521 ( .A(n15606), .B(n15607), .Z(n15854) );
  AND U15522 ( .A(n15855), .B(n15856), .Z(n15607) );
  NANDN U15523 ( .A(n15857), .B(n15858), .Z(n15856) );
  NANDN U15524 ( .A(n15859), .B(n15860), .Z(n15855) );
  NANDN U15525 ( .A(n15858), .B(n15857), .Z(n15860) );
  ANDN U15526 ( .B(\stack[1][23] ), .A(n5614), .Z(n15606) );
  XNOR U15527 ( .A(n15612), .B(n15861), .Z(n15605) );
  XNOR U15528 ( .A(n15613), .B(n15614), .Z(n15861) );
  AND U15529 ( .A(n15862), .B(n15863), .Z(n15614) );
  NAND U15530 ( .A(n15864), .B(n15865), .Z(n15863) );
  NANDN U15531 ( .A(n15866), .B(n15867), .Z(n15862) );
  OR U15532 ( .A(n15864), .B(n15865), .Z(n15867) );
  ANDN U15533 ( .B(\stack[1][24] ), .A(n5590), .Z(n15613) );
  XNOR U15534 ( .A(n15619), .B(n15868), .Z(n15612) );
  XNOR U15535 ( .A(n15620), .B(n15621), .Z(n15868) );
  AND U15536 ( .A(n15869), .B(n15870), .Z(n15621) );
  NANDN U15537 ( .A(n15871), .B(n15872), .Z(n15870) );
  NANDN U15538 ( .A(n15873), .B(n15874), .Z(n15869) );
  NANDN U15539 ( .A(n15872), .B(n15871), .Z(n15874) );
  ANDN U15540 ( .B(\stack[1][25] ), .A(n5566), .Z(n15620) );
  XNOR U15541 ( .A(n15626), .B(n15875), .Z(n15619) );
  XNOR U15542 ( .A(n15627), .B(n15628), .Z(n15875) );
  AND U15543 ( .A(n15876), .B(n15877), .Z(n15628) );
  NAND U15544 ( .A(n15878), .B(n15879), .Z(n15877) );
  NANDN U15545 ( .A(n15880), .B(n15881), .Z(n15876) );
  OR U15546 ( .A(n15878), .B(n15879), .Z(n15881) );
  ANDN U15547 ( .B(\stack[1][26] ), .A(n5542), .Z(n15627) );
  XNOR U15548 ( .A(n15633), .B(n15882), .Z(n15626) );
  XNOR U15549 ( .A(n15634), .B(n15635), .Z(n15882) );
  AND U15550 ( .A(n15883), .B(n15884), .Z(n15635) );
  NANDN U15551 ( .A(n15885), .B(n15886), .Z(n15884) );
  NANDN U15552 ( .A(n15887), .B(n15888), .Z(n15883) );
  NANDN U15553 ( .A(n15886), .B(n15885), .Z(n15888) );
  ANDN U15554 ( .B(\stack[1][27] ), .A(n5518), .Z(n15634) );
  XNOR U15555 ( .A(n15640), .B(n15889), .Z(n15633) );
  XNOR U15556 ( .A(n15641), .B(n15642), .Z(n15889) );
  AND U15557 ( .A(n15890), .B(n15891), .Z(n15642) );
  NAND U15558 ( .A(n15892), .B(n15893), .Z(n15891) );
  NANDN U15559 ( .A(n15894), .B(n15895), .Z(n15890) );
  OR U15560 ( .A(n15892), .B(n15893), .Z(n15895) );
  ANDN U15561 ( .B(\stack[1][28] ), .A(n5494), .Z(n15641) );
  XNOR U15562 ( .A(n15647), .B(n15896), .Z(n15640) );
  XNOR U15563 ( .A(n15648), .B(n15649), .Z(n15896) );
  AND U15564 ( .A(n15897), .B(n15898), .Z(n15649) );
  NANDN U15565 ( .A(n15899), .B(n15900), .Z(n15898) );
  NANDN U15566 ( .A(n15901), .B(n15902), .Z(n15897) );
  NANDN U15567 ( .A(n15900), .B(n15899), .Z(n15902) );
  ANDN U15568 ( .B(\stack[1][29] ), .A(n5470), .Z(n15648) );
  XNOR U15569 ( .A(n15654), .B(n15903), .Z(n15647) );
  XNOR U15570 ( .A(n15655), .B(n15656), .Z(n15903) );
  AND U15571 ( .A(n15904), .B(n15905), .Z(n15656) );
  NAND U15572 ( .A(n15906), .B(n15907), .Z(n15905) );
  NANDN U15573 ( .A(n15908), .B(n15909), .Z(n15904) );
  OR U15574 ( .A(n15906), .B(n15907), .Z(n15909) );
  ANDN U15575 ( .B(\stack[1][30] ), .A(n5446), .Z(n15655) );
  XNOR U15576 ( .A(n15661), .B(n15910), .Z(n15654) );
  XNOR U15577 ( .A(n15662), .B(n15663), .Z(n15910) );
  AND U15578 ( .A(n15911), .B(n15912), .Z(n15663) );
  NANDN U15579 ( .A(n15913), .B(n15914), .Z(n15912) );
  NANDN U15580 ( .A(n15915), .B(n15916), .Z(n15911) );
  NANDN U15581 ( .A(n15914), .B(n15913), .Z(n15916) );
  ANDN U15582 ( .B(\stack[1][31] ), .A(n5422), .Z(n15662) );
  XNOR U15583 ( .A(n15668), .B(n15917), .Z(n15661) );
  XNOR U15584 ( .A(n15669), .B(n15670), .Z(n15917) );
  AND U15585 ( .A(n15918), .B(n15919), .Z(n15670) );
  NAND U15586 ( .A(n15920), .B(n15921), .Z(n15919) );
  NANDN U15587 ( .A(n15922), .B(n15923), .Z(n15918) );
  OR U15588 ( .A(n15920), .B(n15921), .Z(n15923) );
  ANDN U15589 ( .B(\stack[1][32] ), .A(n5398), .Z(n15669) );
  XNOR U15590 ( .A(n15675), .B(n15924), .Z(n15668) );
  XNOR U15591 ( .A(n15676), .B(n15677), .Z(n15924) );
  AND U15592 ( .A(n15925), .B(n15926), .Z(n15677) );
  NANDN U15593 ( .A(n15927), .B(n15928), .Z(n15926) );
  NANDN U15594 ( .A(n15929), .B(n15930), .Z(n15925) );
  NANDN U15595 ( .A(n15928), .B(n15927), .Z(n15930) );
  ANDN U15596 ( .B(\stack[1][33] ), .A(n5374), .Z(n15676) );
  XNOR U15597 ( .A(n15682), .B(n15931), .Z(n15675) );
  XNOR U15598 ( .A(n15683), .B(n15684), .Z(n15931) );
  AND U15599 ( .A(n15932), .B(n15933), .Z(n15684) );
  NAND U15600 ( .A(n15934), .B(n15935), .Z(n15933) );
  NANDN U15601 ( .A(n15936), .B(n15937), .Z(n15932) );
  OR U15602 ( .A(n15934), .B(n15935), .Z(n15937) );
  ANDN U15603 ( .B(\stack[1][34] ), .A(n5350), .Z(n15683) );
  XNOR U15604 ( .A(n15689), .B(n15938), .Z(n15682) );
  XNOR U15605 ( .A(n15690), .B(n15691), .Z(n15938) );
  AND U15606 ( .A(n15939), .B(n15940), .Z(n15691) );
  NANDN U15607 ( .A(n15941), .B(n15942), .Z(n15940) );
  NANDN U15608 ( .A(n15943), .B(n15944), .Z(n15939) );
  NANDN U15609 ( .A(n15942), .B(n15941), .Z(n15944) );
  ANDN U15610 ( .B(\stack[1][35] ), .A(n5326), .Z(n15690) );
  XNOR U15611 ( .A(n15696), .B(n15945), .Z(n15689) );
  XNOR U15612 ( .A(n15697), .B(n15698), .Z(n15945) );
  AND U15613 ( .A(n15946), .B(n15947), .Z(n15698) );
  NAND U15614 ( .A(n15948), .B(n15949), .Z(n15947) );
  NANDN U15615 ( .A(n15950), .B(n15951), .Z(n15946) );
  OR U15616 ( .A(n15948), .B(n15949), .Z(n15951) );
  ANDN U15617 ( .B(\stack[1][36] ), .A(n5302), .Z(n15697) );
  XNOR U15618 ( .A(n15704), .B(n15952), .Z(n15696) );
  XOR U15619 ( .A(n15705), .B(n15706), .Z(n15952) );
  NAND U15620 ( .A(n15953), .B(n15954), .Z(n15706) );
  NANDN U15621 ( .A(n15955), .B(n15956), .Z(n15954) );
  OR U15622 ( .A(n15957), .B(n15958), .Z(n15956) );
  AND U15623 ( .A(\stack[0][5] ), .B(\stack[1][37] ), .Z(n15705) );
  XNOR U15624 ( .A(n15711), .B(n15959), .Z(n15704) );
  XNOR U15625 ( .A(n15710), .B(n15713), .Z(n15959) );
  AND U15626 ( .A(\stack[0][4] ), .B(\stack[1][38] ), .Z(n15713) );
  AND U15627 ( .A(n15960), .B(n15961), .Z(n15710) );
  NAND U15628 ( .A(n15962), .B(n15963), .Z(n15961) );
  OR U15629 ( .A(n15964), .B(n15965), .Z(n15962) );
  XNOR U15630 ( .A(n15717), .B(n15966), .Z(n15711) );
  XNOR U15631 ( .A(n15718), .B(n15719), .Z(n15966) );
  AND U15632 ( .A(n15967), .B(n15968), .Z(n15719) );
  NAND U15633 ( .A(n15969), .B(n15970), .Z(n15968) );
  NAND U15634 ( .A(n15971), .B(n15972), .Z(n15967) );
  OR U15635 ( .A(n15969), .B(n15970), .Z(n15971) );
  ANDN U15636 ( .B(\stack[1][39] ), .A(n5230), .Z(n15718) );
  XNOR U15637 ( .A(n15724), .B(n15973), .Z(n15717) );
  XNOR U15638 ( .A(n15725), .B(n15727), .Z(n15973) );
  ANDN U15639 ( .B(n15974), .A(n15975), .Z(n15727) );
  ANDN U15640 ( .B(\stack[0][0] ), .A(n6156), .Z(n15974) );
  ANDN U15641 ( .B(\stack[1][40] ), .A(n5206), .Z(n15725) );
  XOR U15642 ( .A(n15730), .B(n15976), .Z(n15724) );
  NANDN U15643 ( .A(n5160), .B(\stack[1][42] ), .Z(n15976) );
  NANDN U15644 ( .A(n6156), .B(\stack[0][1] ), .Z(n15730) );
  ANDN U15645 ( .B(\stack[0][37] ), .A(n5292), .Z(n9104) );
  AND U15646 ( .A(n15977), .B(n15978), .Z(n9105) );
  NANDN U15647 ( .A(n9112), .B(n15979), .Z(n15977) );
  NANDN U15648 ( .A(n9111), .B(n9109), .Z(n15979) );
  XNOR U15649 ( .A(n15738), .B(n15980), .Z(n9109) );
  XNOR U15650 ( .A(n15739), .B(n15740), .Z(n15980) );
  AND U15651 ( .A(n15981), .B(n15982), .Z(n15740) );
  NANDN U15652 ( .A(n15983), .B(n15984), .Z(n15982) );
  NANDN U15653 ( .A(n15985), .B(n15986), .Z(n15981) );
  NANDN U15654 ( .A(n15984), .B(n15983), .Z(n15986) );
  ANDN U15655 ( .B(\stack[0][35] ), .A(n5316), .Z(n15739) );
  XNOR U15656 ( .A(n15745), .B(n15987), .Z(n15738) );
  XNOR U15657 ( .A(n15746), .B(n15747), .Z(n15987) );
  AND U15658 ( .A(n15988), .B(n15989), .Z(n15747) );
  NAND U15659 ( .A(n15990), .B(n15991), .Z(n15989) );
  NANDN U15660 ( .A(n15992), .B(n15993), .Z(n15988) );
  OR U15661 ( .A(n15990), .B(n15991), .Z(n15993) );
  ANDN U15662 ( .B(\stack[0][34] ), .A(n5340), .Z(n15746) );
  XNOR U15663 ( .A(n15752), .B(n15994), .Z(n15745) );
  XNOR U15664 ( .A(n15753), .B(n15754), .Z(n15994) );
  AND U15665 ( .A(n15995), .B(n15996), .Z(n15754) );
  NANDN U15666 ( .A(n15997), .B(n15998), .Z(n15996) );
  NANDN U15667 ( .A(n15999), .B(n16000), .Z(n15995) );
  NANDN U15668 ( .A(n15998), .B(n15997), .Z(n16000) );
  ANDN U15669 ( .B(\stack[0][33] ), .A(n5364), .Z(n15753) );
  XNOR U15670 ( .A(n15759), .B(n16001), .Z(n15752) );
  XNOR U15671 ( .A(n15760), .B(n15761), .Z(n16001) );
  AND U15672 ( .A(n16002), .B(n16003), .Z(n15761) );
  NAND U15673 ( .A(n16004), .B(n16005), .Z(n16003) );
  NANDN U15674 ( .A(n16006), .B(n16007), .Z(n16002) );
  OR U15675 ( .A(n16004), .B(n16005), .Z(n16007) );
  ANDN U15676 ( .B(\stack[0][32] ), .A(n5387), .Z(n15760) );
  XNOR U15677 ( .A(n15766), .B(n16008), .Z(n15759) );
  XNOR U15678 ( .A(n15767), .B(n15768), .Z(n16008) );
  AND U15679 ( .A(n16009), .B(n16010), .Z(n15768) );
  NANDN U15680 ( .A(n16011), .B(n16012), .Z(n16010) );
  NANDN U15681 ( .A(n16013), .B(n16014), .Z(n16009) );
  NANDN U15682 ( .A(n16012), .B(n16011), .Z(n16014) );
  ANDN U15683 ( .B(\stack[1][10] ), .A(n5902), .Z(n15767) );
  XNOR U15684 ( .A(n15773), .B(n16015), .Z(n15766) );
  XNOR U15685 ( .A(n15774), .B(n15775), .Z(n16015) );
  AND U15686 ( .A(n16016), .B(n16017), .Z(n15775) );
  NAND U15687 ( .A(n16018), .B(n16019), .Z(n16017) );
  NANDN U15688 ( .A(n16020), .B(n16021), .Z(n16016) );
  OR U15689 ( .A(n16018), .B(n16019), .Z(n16021) );
  ANDN U15690 ( .B(\stack[1][11] ), .A(n5878), .Z(n15774) );
  XNOR U15691 ( .A(n15780), .B(n16022), .Z(n15773) );
  XNOR U15692 ( .A(n15781), .B(n15782), .Z(n16022) );
  AND U15693 ( .A(n16023), .B(n16024), .Z(n15782) );
  NANDN U15694 ( .A(n16025), .B(n16026), .Z(n16024) );
  NANDN U15695 ( .A(n16027), .B(n16028), .Z(n16023) );
  NANDN U15696 ( .A(n16026), .B(n16025), .Z(n16028) );
  ANDN U15697 ( .B(\stack[1][12] ), .A(n5854), .Z(n15781) );
  XNOR U15698 ( .A(n15787), .B(n16029), .Z(n15780) );
  XNOR U15699 ( .A(n15788), .B(n15789), .Z(n16029) );
  AND U15700 ( .A(n16030), .B(n16031), .Z(n15789) );
  NAND U15701 ( .A(n16032), .B(n16033), .Z(n16031) );
  NANDN U15702 ( .A(n16034), .B(n16035), .Z(n16030) );
  OR U15703 ( .A(n16032), .B(n16033), .Z(n16035) );
  ANDN U15704 ( .B(\stack[1][13] ), .A(n5830), .Z(n15788) );
  XNOR U15705 ( .A(n15794), .B(n16036), .Z(n15787) );
  XNOR U15706 ( .A(n15795), .B(n15796), .Z(n16036) );
  AND U15707 ( .A(n16037), .B(n16038), .Z(n15796) );
  NANDN U15708 ( .A(n16039), .B(n16040), .Z(n16038) );
  NANDN U15709 ( .A(n16041), .B(n16042), .Z(n16037) );
  NANDN U15710 ( .A(n16040), .B(n16039), .Z(n16042) );
  ANDN U15711 ( .B(\stack[1][14] ), .A(n5806), .Z(n15795) );
  XNOR U15712 ( .A(n15801), .B(n16043), .Z(n15794) );
  XNOR U15713 ( .A(n15802), .B(n15803), .Z(n16043) );
  AND U15714 ( .A(n16044), .B(n16045), .Z(n15803) );
  NAND U15715 ( .A(n16046), .B(n16047), .Z(n16045) );
  NANDN U15716 ( .A(n16048), .B(n16049), .Z(n16044) );
  OR U15717 ( .A(n16046), .B(n16047), .Z(n16049) );
  ANDN U15718 ( .B(\stack[1][15] ), .A(n5782), .Z(n15802) );
  XNOR U15719 ( .A(n15808), .B(n16050), .Z(n15801) );
  XNOR U15720 ( .A(n15809), .B(n15810), .Z(n16050) );
  AND U15721 ( .A(n16051), .B(n16052), .Z(n15810) );
  NANDN U15722 ( .A(n16053), .B(n16054), .Z(n16052) );
  NANDN U15723 ( .A(n16055), .B(n16056), .Z(n16051) );
  NANDN U15724 ( .A(n16054), .B(n16053), .Z(n16056) );
  ANDN U15725 ( .B(\stack[1][16] ), .A(n5758), .Z(n15809) );
  XNOR U15726 ( .A(n15815), .B(n16057), .Z(n15808) );
  XNOR U15727 ( .A(n15816), .B(n15817), .Z(n16057) );
  AND U15728 ( .A(n16058), .B(n16059), .Z(n15817) );
  NAND U15729 ( .A(n16060), .B(n16061), .Z(n16059) );
  NANDN U15730 ( .A(n16062), .B(n16063), .Z(n16058) );
  OR U15731 ( .A(n16060), .B(n16061), .Z(n16063) );
  ANDN U15732 ( .B(\stack[1][17] ), .A(n5734), .Z(n15816) );
  XNOR U15733 ( .A(n15822), .B(n16064), .Z(n15815) );
  XNOR U15734 ( .A(n15823), .B(n15824), .Z(n16064) );
  AND U15735 ( .A(n16065), .B(n16066), .Z(n15824) );
  NANDN U15736 ( .A(n16067), .B(n16068), .Z(n16066) );
  NANDN U15737 ( .A(n16069), .B(n16070), .Z(n16065) );
  NANDN U15738 ( .A(n16068), .B(n16067), .Z(n16070) );
  ANDN U15739 ( .B(\stack[1][18] ), .A(n5710), .Z(n15823) );
  XNOR U15740 ( .A(n15829), .B(n16071), .Z(n15822) );
  XNOR U15741 ( .A(n15830), .B(n15831), .Z(n16071) );
  AND U15742 ( .A(n16072), .B(n16073), .Z(n15831) );
  NAND U15743 ( .A(n16074), .B(n16075), .Z(n16073) );
  NANDN U15744 ( .A(n16076), .B(n16077), .Z(n16072) );
  OR U15745 ( .A(n16074), .B(n16075), .Z(n16077) );
  ANDN U15746 ( .B(\stack[1][19] ), .A(n5686), .Z(n15830) );
  XNOR U15747 ( .A(n15836), .B(n16078), .Z(n15829) );
  XNOR U15748 ( .A(n15837), .B(n15838), .Z(n16078) );
  AND U15749 ( .A(n16079), .B(n16080), .Z(n15838) );
  NANDN U15750 ( .A(n16081), .B(n16082), .Z(n16080) );
  NANDN U15751 ( .A(n16083), .B(n16084), .Z(n16079) );
  NANDN U15752 ( .A(n16082), .B(n16081), .Z(n16084) );
  ANDN U15753 ( .B(\stack[1][20] ), .A(n5662), .Z(n15837) );
  XNOR U15754 ( .A(n15843), .B(n16085), .Z(n15836) );
  XNOR U15755 ( .A(n15844), .B(n15845), .Z(n16085) );
  AND U15756 ( .A(n16086), .B(n16087), .Z(n15845) );
  NAND U15757 ( .A(n16088), .B(n16089), .Z(n16087) );
  NANDN U15758 ( .A(n16090), .B(n16091), .Z(n16086) );
  OR U15759 ( .A(n16088), .B(n16089), .Z(n16091) );
  ANDN U15760 ( .B(\stack[1][21] ), .A(n5638), .Z(n15844) );
  XNOR U15761 ( .A(n15850), .B(n16092), .Z(n15843) );
  XNOR U15762 ( .A(n15851), .B(n15852), .Z(n16092) );
  AND U15763 ( .A(n16093), .B(n16094), .Z(n15852) );
  NANDN U15764 ( .A(n16095), .B(n16096), .Z(n16094) );
  NANDN U15765 ( .A(n16097), .B(n16098), .Z(n16093) );
  NANDN U15766 ( .A(n16096), .B(n16095), .Z(n16098) );
  ANDN U15767 ( .B(\stack[1][22] ), .A(n5614), .Z(n15851) );
  XNOR U15768 ( .A(n15857), .B(n16099), .Z(n15850) );
  XNOR U15769 ( .A(n15858), .B(n15859), .Z(n16099) );
  AND U15770 ( .A(n16100), .B(n16101), .Z(n15859) );
  NAND U15771 ( .A(n16102), .B(n16103), .Z(n16101) );
  NANDN U15772 ( .A(n16104), .B(n16105), .Z(n16100) );
  OR U15773 ( .A(n16102), .B(n16103), .Z(n16105) );
  ANDN U15774 ( .B(\stack[1][23] ), .A(n5590), .Z(n15858) );
  XNOR U15775 ( .A(n15864), .B(n16106), .Z(n15857) );
  XNOR U15776 ( .A(n15865), .B(n15866), .Z(n16106) );
  AND U15777 ( .A(n16107), .B(n16108), .Z(n15866) );
  NANDN U15778 ( .A(n16109), .B(n16110), .Z(n16108) );
  NANDN U15779 ( .A(n16111), .B(n16112), .Z(n16107) );
  NANDN U15780 ( .A(n16110), .B(n16109), .Z(n16112) );
  ANDN U15781 ( .B(\stack[1][24] ), .A(n5566), .Z(n15865) );
  XNOR U15782 ( .A(n15871), .B(n16113), .Z(n15864) );
  XNOR U15783 ( .A(n15872), .B(n15873), .Z(n16113) );
  AND U15784 ( .A(n16114), .B(n16115), .Z(n15873) );
  NAND U15785 ( .A(n16116), .B(n16117), .Z(n16115) );
  NANDN U15786 ( .A(n16118), .B(n16119), .Z(n16114) );
  OR U15787 ( .A(n16116), .B(n16117), .Z(n16119) );
  ANDN U15788 ( .B(\stack[1][25] ), .A(n5542), .Z(n15872) );
  XNOR U15789 ( .A(n15878), .B(n16120), .Z(n15871) );
  XNOR U15790 ( .A(n15879), .B(n15880), .Z(n16120) );
  AND U15791 ( .A(n16121), .B(n16122), .Z(n15880) );
  NANDN U15792 ( .A(n16123), .B(n16124), .Z(n16122) );
  NANDN U15793 ( .A(n16125), .B(n16126), .Z(n16121) );
  NANDN U15794 ( .A(n16124), .B(n16123), .Z(n16126) );
  ANDN U15795 ( .B(\stack[1][26] ), .A(n5518), .Z(n15879) );
  XNOR U15796 ( .A(n15885), .B(n16127), .Z(n15878) );
  XNOR U15797 ( .A(n15886), .B(n15887), .Z(n16127) );
  AND U15798 ( .A(n16128), .B(n16129), .Z(n15887) );
  NAND U15799 ( .A(n16130), .B(n16131), .Z(n16129) );
  NANDN U15800 ( .A(n16132), .B(n16133), .Z(n16128) );
  OR U15801 ( .A(n16130), .B(n16131), .Z(n16133) );
  ANDN U15802 ( .B(\stack[1][27] ), .A(n5494), .Z(n15886) );
  XNOR U15803 ( .A(n15892), .B(n16134), .Z(n15885) );
  XNOR U15804 ( .A(n15893), .B(n15894), .Z(n16134) );
  AND U15805 ( .A(n16135), .B(n16136), .Z(n15894) );
  NANDN U15806 ( .A(n16137), .B(n16138), .Z(n16136) );
  NANDN U15807 ( .A(n16139), .B(n16140), .Z(n16135) );
  NANDN U15808 ( .A(n16138), .B(n16137), .Z(n16140) );
  ANDN U15809 ( .B(\stack[1][28] ), .A(n5470), .Z(n15893) );
  XNOR U15810 ( .A(n15899), .B(n16141), .Z(n15892) );
  XNOR U15811 ( .A(n15900), .B(n15901), .Z(n16141) );
  AND U15812 ( .A(n16142), .B(n16143), .Z(n15901) );
  NAND U15813 ( .A(n16144), .B(n16145), .Z(n16143) );
  NANDN U15814 ( .A(n16146), .B(n16147), .Z(n16142) );
  OR U15815 ( .A(n16144), .B(n16145), .Z(n16147) );
  ANDN U15816 ( .B(\stack[1][29] ), .A(n5446), .Z(n15900) );
  XNOR U15817 ( .A(n15906), .B(n16148), .Z(n15899) );
  XNOR U15818 ( .A(n15907), .B(n15908), .Z(n16148) );
  AND U15819 ( .A(n16149), .B(n16150), .Z(n15908) );
  NANDN U15820 ( .A(n16151), .B(n16152), .Z(n16150) );
  NANDN U15821 ( .A(n16153), .B(n16154), .Z(n16149) );
  NANDN U15822 ( .A(n16152), .B(n16151), .Z(n16154) );
  ANDN U15823 ( .B(\stack[1][30] ), .A(n5422), .Z(n15907) );
  XNOR U15824 ( .A(n15913), .B(n16155), .Z(n15906) );
  XNOR U15825 ( .A(n15914), .B(n15915), .Z(n16155) );
  AND U15826 ( .A(n16156), .B(n16157), .Z(n15915) );
  NAND U15827 ( .A(n16158), .B(n16159), .Z(n16157) );
  NANDN U15828 ( .A(n16160), .B(n16161), .Z(n16156) );
  OR U15829 ( .A(n16158), .B(n16159), .Z(n16161) );
  ANDN U15830 ( .B(\stack[1][31] ), .A(n5398), .Z(n15914) );
  XNOR U15831 ( .A(n15920), .B(n16162), .Z(n15913) );
  XNOR U15832 ( .A(n15921), .B(n15922), .Z(n16162) );
  AND U15833 ( .A(n16163), .B(n16164), .Z(n15922) );
  NANDN U15834 ( .A(n16165), .B(n16166), .Z(n16164) );
  NANDN U15835 ( .A(n16167), .B(n16168), .Z(n16163) );
  NANDN U15836 ( .A(n16166), .B(n16165), .Z(n16168) );
  ANDN U15837 ( .B(\stack[1][32] ), .A(n5374), .Z(n15921) );
  XNOR U15838 ( .A(n15927), .B(n16169), .Z(n15920) );
  XNOR U15839 ( .A(n15928), .B(n15929), .Z(n16169) );
  AND U15840 ( .A(n16170), .B(n16171), .Z(n15929) );
  NAND U15841 ( .A(n16172), .B(n16173), .Z(n16171) );
  NANDN U15842 ( .A(n16174), .B(n16175), .Z(n16170) );
  OR U15843 ( .A(n16172), .B(n16173), .Z(n16175) );
  ANDN U15844 ( .B(\stack[1][33] ), .A(n5350), .Z(n15928) );
  XNOR U15845 ( .A(n15934), .B(n16176), .Z(n15927) );
  XNOR U15846 ( .A(n15935), .B(n15936), .Z(n16176) );
  AND U15847 ( .A(n16177), .B(n16178), .Z(n15936) );
  NANDN U15848 ( .A(n16179), .B(n16180), .Z(n16178) );
  NANDN U15849 ( .A(n16181), .B(n16182), .Z(n16177) );
  NANDN U15850 ( .A(n16180), .B(n16179), .Z(n16182) );
  ANDN U15851 ( .B(\stack[1][34] ), .A(n5326), .Z(n15935) );
  XNOR U15852 ( .A(n15941), .B(n16183), .Z(n15934) );
  XNOR U15853 ( .A(n15942), .B(n15943), .Z(n16183) );
  AND U15854 ( .A(n16184), .B(n16185), .Z(n15943) );
  NAND U15855 ( .A(n16186), .B(n16187), .Z(n16185) );
  NANDN U15856 ( .A(n16188), .B(n16189), .Z(n16184) );
  OR U15857 ( .A(n16186), .B(n16187), .Z(n16189) );
  ANDN U15858 ( .B(\stack[1][35] ), .A(n5302), .Z(n15942) );
  XNOR U15859 ( .A(n15948), .B(n16190), .Z(n15941) );
  XNOR U15860 ( .A(n15949), .B(n15950), .Z(n16190) );
  AND U15861 ( .A(n16191), .B(n16192), .Z(n15950) );
  NANDN U15862 ( .A(n16193), .B(n16194), .Z(n16192) );
  NANDN U15863 ( .A(n16195), .B(n16196), .Z(n16191) );
  NANDN U15864 ( .A(n16194), .B(n16193), .Z(n16196) );
  ANDN U15865 ( .B(\stack[1][36] ), .A(n5278), .Z(n15949) );
  XNOR U15866 ( .A(n15955), .B(n16197), .Z(n15948) );
  XOR U15867 ( .A(n15957), .B(n15958), .Z(n16197) );
  NAND U15868 ( .A(n16198), .B(n16199), .Z(n15958) );
  NAND U15869 ( .A(n16200), .B(n16201), .Z(n16199) );
  OR U15870 ( .A(n16202), .B(n16203), .Z(n16200) );
  AND U15871 ( .A(\stack[0][4] ), .B(\stack[1][37] ), .Z(n15957) );
  XNOR U15872 ( .A(n15964), .B(n16204), .Z(n15955) );
  XOR U15873 ( .A(n15965), .B(n15963), .Z(n16204) );
  AND U15874 ( .A(\stack[0][3] ), .B(\stack[1][38] ), .Z(n15963) );
  NAND U15875 ( .A(n16205), .B(n16206), .Z(n15965) );
  NAND U15876 ( .A(n16207), .B(n16208), .Z(n16206) );
  NAND U15877 ( .A(n16209), .B(n16210), .Z(n16205) );
  OR U15878 ( .A(n16207), .B(n16208), .Z(n16209) );
  XNOR U15879 ( .A(n15969), .B(n16211), .Z(n15964) );
  XNOR U15880 ( .A(n15970), .B(n15972), .Z(n16211) );
  ANDN U15881 ( .B(n16212), .A(n16213), .Z(n15972) );
  ANDN U15882 ( .B(\stack[0][0] ), .A(n6132), .Z(n16212) );
  ANDN U15883 ( .B(\stack[1][39] ), .A(n5206), .Z(n15970) );
  XOR U15884 ( .A(n15975), .B(n16214), .Z(n15969) );
  NANDN U15885 ( .A(n5160), .B(\stack[1][41] ), .Z(n16214) );
  NANDN U15886 ( .A(n6132), .B(\stack[0][1] ), .Z(n15975) );
  ANDN U15887 ( .B(\stack[1][5] ), .A(n6022), .Z(n9111) );
  AND U15888 ( .A(n16215), .B(n16216), .Z(n9112) );
  NANDN U15889 ( .A(n9116), .B(n9118), .Z(n16216) );
  NANDN U15890 ( .A(n9119), .B(n16217), .Z(n16215) );
  NANDN U15891 ( .A(n9118), .B(n9116), .Z(n16217) );
  XOR U15892 ( .A(n15983), .B(n16218), .Z(n9116) );
  XNOR U15893 ( .A(n15984), .B(n15985), .Z(n16218) );
  AND U15894 ( .A(n16219), .B(n16220), .Z(n15985) );
  NAND U15895 ( .A(n16221), .B(n16222), .Z(n16220) );
  NANDN U15896 ( .A(n16223), .B(n16224), .Z(n16219) );
  OR U15897 ( .A(n16221), .B(n16222), .Z(n16224) );
  ANDN U15898 ( .B(\stack[0][34] ), .A(n5316), .Z(n15984) );
  XNOR U15899 ( .A(n15990), .B(n16225), .Z(n15983) );
  XNOR U15900 ( .A(n15991), .B(n15992), .Z(n16225) );
  AND U15901 ( .A(n16226), .B(n16227), .Z(n15992) );
  NANDN U15902 ( .A(n16228), .B(n16229), .Z(n16227) );
  NANDN U15903 ( .A(n16230), .B(n16231), .Z(n16226) );
  NANDN U15904 ( .A(n16229), .B(n16228), .Z(n16231) );
  ANDN U15905 ( .B(\stack[0][33] ), .A(n5340), .Z(n15991) );
  XNOR U15906 ( .A(n15997), .B(n16232), .Z(n15990) );
  XNOR U15907 ( .A(n15998), .B(n15999), .Z(n16232) );
  AND U15908 ( .A(n16233), .B(n16234), .Z(n15999) );
  NAND U15909 ( .A(n16235), .B(n16236), .Z(n16234) );
  NANDN U15910 ( .A(n16237), .B(n16238), .Z(n16233) );
  OR U15911 ( .A(n16235), .B(n16236), .Z(n16238) );
  ANDN U15912 ( .B(\stack[0][32] ), .A(n5364), .Z(n15998) );
  XNOR U15913 ( .A(n16004), .B(n16239), .Z(n15997) );
  XNOR U15914 ( .A(n16005), .B(n16006), .Z(n16239) );
  AND U15915 ( .A(n16240), .B(n16241), .Z(n16006) );
  NANDN U15916 ( .A(n16242), .B(n16243), .Z(n16241) );
  NANDN U15917 ( .A(n16244), .B(n16245), .Z(n16240) );
  NANDN U15918 ( .A(n16243), .B(n16242), .Z(n16245) );
  ANDN U15919 ( .B(\stack[0][31] ), .A(n5387), .Z(n16005) );
  XNOR U15920 ( .A(n16011), .B(n16246), .Z(n16004) );
  XNOR U15921 ( .A(n16012), .B(n16013), .Z(n16246) );
  AND U15922 ( .A(n16247), .B(n16248), .Z(n16013) );
  NAND U15923 ( .A(n16249), .B(n16250), .Z(n16248) );
  NANDN U15924 ( .A(n16251), .B(n16252), .Z(n16247) );
  OR U15925 ( .A(n16249), .B(n16250), .Z(n16252) );
  ANDN U15926 ( .B(\stack[1][10] ), .A(n5878), .Z(n16012) );
  XNOR U15927 ( .A(n16018), .B(n16253), .Z(n16011) );
  XNOR U15928 ( .A(n16019), .B(n16020), .Z(n16253) );
  AND U15929 ( .A(n16254), .B(n16255), .Z(n16020) );
  NANDN U15930 ( .A(n16256), .B(n16257), .Z(n16255) );
  NANDN U15931 ( .A(n16258), .B(n16259), .Z(n16254) );
  NANDN U15932 ( .A(n16257), .B(n16256), .Z(n16259) );
  ANDN U15933 ( .B(\stack[1][11] ), .A(n5854), .Z(n16019) );
  XNOR U15934 ( .A(n16025), .B(n16260), .Z(n16018) );
  XNOR U15935 ( .A(n16026), .B(n16027), .Z(n16260) );
  AND U15936 ( .A(n16261), .B(n16262), .Z(n16027) );
  NAND U15937 ( .A(n16263), .B(n16264), .Z(n16262) );
  NANDN U15938 ( .A(n16265), .B(n16266), .Z(n16261) );
  OR U15939 ( .A(n16263), .B(n16264), .Z(n16266) );
  ANDN U15940 ( .B(\stack[1][12] ), .A(n5830), .Z(n16026) );
  XNOR U15941 ( .A(n16032), .B(n16267), .Z(n16025) );
  XNOR U15942 ( .A(n16033), .B(n16034), .Z(n16267) );
  AND U15943 ( .A(n16268), .B(n16269), .Z(n16034) );
  NANDN U15944 ( .A(n16270), .B(n16271), .Z(n16269) );
  NANDN U15945 ( .A(n16272), .B(n16273), .Z(n16268) );
  NANDN U15946 ( .A(n16271), .B(n16270), .Z(n16273) );
  ANDN U15947 ( .B(\stack[1][13] ), .A(n5806), .Z(n16033) );
  XNOR U15948 ( .A(n16039), .B(n16274), .Z(n16032) );
  XNOR U15949 ( .A(n16040), .B(n16041), .Z(n16274) );
  AND U15950 ( .A(n16275), .B(n16276), .Z(n16041) );
  NAND U15951 ( .A(n16277), .B(n16278), .Z(n16276) );
  NANDN U15952 ( .A(n16279), .B(n16280), .Z(n16275) );
  OR U15953 ( .A(n16277), .B(n16278), .Z(n16280) );
  ANDN U15954 ( .B(\stack[1][14] ), .A(n5782), .Z(n16040) );
  XNOR U15955 ( .A(n16046), .B(n16281), .Z(n16039) );
  XNOR U15956 ( .A(n16047), .B(n16048), .Z(n16281) );
  AND U15957 ( .A(n16282), .B(n16283), .Z(n16048) );
  NANDN U15958 ( .A(n16284), .B(n16285), .Z(n16283) );
  NANDN U15959 ( .A(n16286), .B(n16287), .Z(n16282) );
  NANDN U15960 ( .A(n16285), .B(n16284), .Z(n16287) );
  ANDN U15961 ( .B(\stack[1][15] ), .A(n5758), .Z(n16047) );
  XNOR U15962 ( .A(n16053), .B(n16288), .Z(n16046) );
  XNOR U15963 ( .A(n16054), .B(n16055), .Z(n16288) );
  AND U15964 ( .A(n16289), .B(n16290), .Z(n16055) );
  NAND U15965 ( .A(n16291), .B(n16292), .Z(n16290) );
  NANDN U15966 ( .A(n16293), .B(n16294), .Z(n16289) );
  OR U15967 ( .A(n16291), .B(n16292), .Z(n16294) );
  ANDN U15968 ( .B(\stack[1][16] ), .A(n5734), .Z(n16054) );
  XNOR U15969 ( .A(n16060), .B(n16295), .Z(n16053) );
  XNOR U15970 ( .A(n16061), .B(n16062), .Z(n16295) );
  AND U15971 ( .A(n16296), .B(n16297), .Z(n16062) );
  NANDN U15972 ( .A(n16298), .B(n16299), .Z(n16297) );
  NANDN U15973 ( .A(n16300), .B(n16301), .Z(n16296) );
  NANDN U15974 ( .A(n16299), .B(n16298), .Z(n16301) );
  ANDN U15975 ( .B(\stack[1][17] ), .A(n5710), .Z(n16061) );
  XNOR U15976 ( .A(n16067), .B(n16302), .Z(n16060) );
  XNOR U15977 ( .A(n16068), .B(n16069), .Z(n16302) );
  AND U15978 ( .A(n16303), .B(n16304), .Z(n16069) );
  NAND U15979 ( .A(n16305), .B(n16306), .Z(n16304) );
  NANDN U15980 ( .A(n16307), .B(n16308), .Z(n16303) );
  OR U15981 ( .A(n16305), .B(n16306), .Z(n16308) );
  ANDN U15982 ( .B(\stack[1][18] ), .A(n5686), .Z(n16068) );
  XNOR U15983 ( .A(n16074), .B(n16309), .Z(n16067) );
  XNOR U15984 ( .A(n16075), .B(n16076), .Z(n16309) );
  AND U15985 ( .A(n16310), .B(n16311), .Z(n16076) );
  NANDN U15986 ( .A(n16312), .B(n16313), .Z(n16311) );
  NANDN U15987 ( .A(n16314), .B(n16315), .Z(n16310) );
  NANDN U15988 ( .A(n16313), .B(n16312), .Z(n16315) );
  ANDN U15989 ( .B(\stack[1][19] ), .A(n5662), .Z(n16075) );
  XNOR U15990 ( .A(n16081), .B(n16316), .Z(n16074) );
  XNOR U15991 ( .A(n16082), .B(n16083), .Z(n16316) );
  AND U15992 ( .A(n16317), .B(n16318), .Z(n16083) );
  NAND U15993 ( .A(n16319), .B(n16320), .Z(n16318) );
  NANDN U15994 ( .A(n16321), .B(n16322), .Z(n16317) );
  OR U15995 ( .A(n16319), .B(n16320), .Z(n16322) );
  ANDN U15996 ( .B(\stack[1][20] ), .A(n5638), .Z(n16082) );
  XNOR U15997 ( .A(n16088), .B(n16323), .Z(n16081) );
  XNOR U15998 ( .A(n16089), .B(n16090), .Z(n16323) );
  AND U15999 ( .A(n16324), .B(n16325), .Z(n16090) );
  NANDN U16000 ( .A(n16326), .B(n16327), .Z(n16325) );
  NANDN U16001 ( .A(n16328), .B(n16329), .Z(n16324) );
  NANDN U16002 ( .A(n16327), .B(n16326), .Z(n16329) );
  ANDN U16003 ( .B(\stack[1][21] ), .A(n5614), .Z(n16089) );
  XNOR U16004 ( .A(n16095), .B(n16330), .Z(n16088) );
  XNOR U16005 ( .A(n16096), .B(n16097), .Z(n16330) );
  AND U16006 ( .A(n16331), .B(n16332), .Z(n16097) );
  NAND U16007 ( .A(n16333), .B(n16334), .Z(n16332) );
  NANDN U16008 ( .A(n16335), .B(n16336), .Z(n16331) );
  OR U16009 ( .A(n16333), .B(n16334), .Z(n16336) );
  ANDN U16010 ( .B(\stack[1][22] ), .A(n5590), .Z(n16096) );
  XNOR U16011 ( .A(n16102), .B(n16337), .Z(n16095) );
  XNOR U16012 ( .A(n16103), .B(n16104), .Z(n16337) );
  AND U16013 ( .A(n16338), .B(n16339), .Z(n16104) );
  NANDN U16014 ( .A(n16340), .B(n16341), .Z(n16339) );
  NANDN U16015 ( .A(n16342), .B(n16343), .Z(n16338) );
  NANDN U16016 ( .A(n16341), .B(n16340), .Z(n16343) );
  ANDN U16017 ( .B(\stack[1][23] ), .A(n5566), .Z(n16103) );
  XNOR U16018 ( .A(n16109), .B(n16344), .Z(n16102) );
  XNOR U16019 ( .A(n16110), .B(n16111), .Z(n16344) );
  AND U16020 ( .A(n16345), .B(n16346), .Z(n16111) );
  NAND U16021 ( .A(n16347), .B(n16348), .Z(n16346) );
  NANDN U16022 ( .A(n16349), .B(n16350), .Z(n16345) );
  OR U16023 ( .A(n16347), .B(n16348), .Z(n16350) );
  ANDN U16024 ( .B(\stack[1][24] ), .A(n5542), .Z(n16110) );
  XNOR U16025 ( .A(n16116), .B(n16351), .Z(n16109) );
  XNOR U16026 ( .A(n16117), .B(n16118), .Z(n16351) );
  AND U16027 ( .A(n16352), .B(n16353), .Z(n16118) );
  NANDN U16028 ( .A(n16354), .B(n16355), .Z(n16353) );
  NANDN U16029 ( .A(n16356), .B(n16357), .Z(n16352) );
  NANDN U16030 ( .A(n16355), .B(n16354), .Z(n16357) );
  ANDN U16031 ( .B(\stack[1][25] ), .A(n5518), .Z(n16117) );
  XNOR U16032 ( .A(n16123), .B(n16358), .Z(n16116) );
  XNOR U16033 ( .A(n16124), .B(n16125), .Z(n16358) );
  AND U16034 ( .A(n16359), .B(n16360), .Z(n16125) );
  NAND U16035 ( .A(n16361), .B(n16362), .Z(n16360) );
  NANDN U16036 ( .A(n16363), .B(n16364), .Z(n16359) );
  OR U16037 ( .A(n16361), .B(n16362), .Z(n16364) );
  ANDN U16038 ( .B(\stack[1][26] ), .A(n5494), .Z(n16124) );
  XNOR U16039 ( .A(n16130), .B(n16365), .Z(n16123) );
  XNOR U16040 ( .A(n16131), .B(n16132), .Z(n16365) );
  AND U16041 ( .A(n16366), .B(n16367), .Z(n16132) );
  NANDN U16042 ( .A(n16368), .B(n16369), .Z(n16367) );
  NANDN U16043 ( .A(n16370), .B(n16371), .Z(n16366) );
  NANDN U16044 ( .A(n16369), .B(n16368), .Z(n16371) );
  ANDN U16045 ( .B(\stack[1][27] ), .A(n5470), .Z(n16131) );
  XNOR U16046 ( .A(n16137), .B(n16372), .Z(n16130) );
  XNOR U16047 ( .A(n16138), .B(n16139), .Z(n16372) );
  AND U16048 ( .A(n16373), .B(n16374), .Z(n16139) );
  NAND U16049 ( .A(n16375), .B(n16376), .Z(n16374) );
  NANDN U16050 ( .A(n16377), .B(n16378), .Z(n16373) );
  OR U16051 ( .A(n16375), .B(n16376), .Z(n16378) );
  ANDN U16052 ( .B(\stack[1][28] ), .A(n5446), .Z(n16138) );
  XNOR U16053 ( .A(n16144), .B(n16379), .Z(n16137) );
  XNOR U16054 ( .A(n16145), .B(n16146), .Z(n16379) );
  AND U16055 ( .A(n16380), .B(n16381), .Z(n16146) );
  NANDN U16056 ( .A(n16382), .B(n16383), .Z(n16381) );
  NANDN U16057 ( .A(n16384), .B(n16385), .Z(n16380) );
  NANDN U16058 ( .A(n16383), .B(n16382), .Z(n16385) );
  ANDN U16059 ( .B(\stack[1][29] ), .A(n5422), .Z(n16145) );
  XNOR U16060 ( .A(n16151), .B(n16386), .Z(n16144) );
  XNOR U16061 ( .A(n16152), .B(n16153), .Z(n16386) );
  AND U16062 ( .A(n16387), .B(n16388), .Z(n16153) );
  NAND U16063 ( .A(n16389), .B(n16390), .Z(n16388) );
  NANDN U16064 ( .A(n16391), .B(n16392), .Z(n16387) );
  OR U16065 ( .A(n16389), .B(n16390), .Z(n16392) );
  ANDN U16066 ( .B(\stack[1][30] ), .A(n5398), .Z(n16152) );
  XNOR U16067 ( .A(n16158), .B(n16393), .Z(n16151) );
  XNOR U16068 ( .A(n16159), .B(n16160), .Z(n16393) );
  AND U16069 ( .A(n16394), .B(n16395), .Z(n16160) );
  NANDN U16070 ( .A(n16396), .B(n16397), .Z(n16395) );
  NANDN U16071 ( .A(n16398), .B(n16399), .Z(n16394) );
  NANDN U16072 ( .A(n16397), .B(n16396), .Z(n16399) );
  ANDN U16073 ( .B(\stack[1][31] ), .A(n5374), .Z(n16159) );
  XNOR U16074 ( .A(n16165), .B(n16400), .Z(n16158) );
  XNOR U16075 ( .A(n16166), .B(n16167), .Z(n16400) );
  AND U16076 ( .A(n16401), .B(n16402), .Z(n16167) );
  NAND U16077 ( .A(n16403), .B(n16404), .Z(n16402) );
  NANDN U16078 ( .A(n16405), .B(n16406), .Z(n16401) );
  OR U16079 ( .A(n16403), .B(n16404), .Z(n16406) );
  ANDN U16080 ( .B(\stack[1][32] ), .A(n5350), .Z(n16166) );
  XNOR U16081 ( .A(n16172), .B(n16407), .Z(n16165) );
  XNOR U16082 ( .A(n16173), .B(n16174), .Z(n16407) );
  AND U16083 ( .A(n16408), .B(n16409), .Z(n16174) );
  NANDN U16084 ( .A(n16410), .B(n16411), .Z(n16409) );
  NANDN U16085 ( .A(n16412), .B(n16413), .Z(n16408) );
  NANDN U16086 ( .A(n16411), .B(n16410), .Z(n16413) );
  ANDN U16087 ( .B(\stack[1][33] ), .A(n5326), .Z(n16173) );
  XNOR U16088 ( .A(n16179), .B(n16414), .Z(n16172) );
  XNOR U16089 ( .A(n16180), .B(n16181), .Z(n16414) );
  AND U16090 ( .A(n16415), .B(n16416), .Z(n16181) );
  NAND U16091 ( .A(n16417), .B(n16418), .Z(n16416) );
  NANDN U16092 ( .A(n16419), .B(n16420), .Z(n16415) );
  OR U16093 ( .A(n16417), .B(n16418), .Z(n16420) );
  ANDN U16094 ( .B(\stack[1][34] ), .A(n5302), .Z(n16180) );
  XNOR U16095 ( .A(n16186), .B(n16421), .Z(n16179) );
  XNOR U16096 ( .A(n16187), .B(n16188), .Z(n16421) );
  AND U16097 ( .A(n16422), .B(n16423), .Z(n16188) );
  NANDN U16098 ( .A(n16424), .B(n16425), .Z(n16423) );
  NANDN U16099 ( .A(n16426), .B(n16427), .Z(n16422) );
  NANDN U16100 ( .A(n16425), .B(n16424), .Z(n16427) );
  ANDN U16101 ( .B(\stack[1][35] ), .A(n5278), .Z(n16187) );
  XNOR U16102 ( .A(n16193), .B(n16428), .Z(n16186) );
  XNOR U16103 ( .A(n16194), .B(n16195), .Z(n16428) );
  AND U16104 ( .A(n16429), .B(n16430), .Z(n16195) );
  NAND U16105 ( .A(n16431), .B(n16432), .Z(n16430) );
  NANDN U16106 ( .A(n16433), .B(n16434), .Z(n16429) );
  OR U16107 ( .A(n16431), .B(n16432), .Z(n16434) );
  ANDN U16108 ( .B(\stack[1][36] ), .A(n5254), .Z(n16194) );
  XNOR U16109 ( .A(n16201), .B(n16435), .Z(n16193) );
  XOR U16110 ( .A(n16202), .B(n16203), .Z(n16435) );
  NAND U16111 ( .A(n16436), .B(n16437), .Z(n16203) );
  NANDN U16112 ( .A(n16438), .B(n16439), .Z(n16437) );
  OR U16113 ( .A(n16440), .B(n16441), .Z(n16439) );
  NAND U16114 ( .A(n16441), .B(n16440), .Z(n16436) );
  AND U16115 ( .A(\stack[0][3] ), .B(\stack[1][37] ), .Z(n16202) );
  XNOR U16116 ( .A(n16207), .B(n16442), .Z(n16201) );
  XNOR U16117 ( .A(n16208), .B(n16210), .Z(n16442) );
  AND U16118 ( .A(\stack[0][2] ), .B(\stack[1][38] ), .Z(n16210) );
  ANDN U16119 ( .B(n16443), .A(n16444), .Z(n16208) );
  ANDN U16120 ( .B(\stack[0][0] ), .A(n6108), .Z(n16443) );
  XOR U16121 ( .A(n16213), .B(n16445), .Z(n16207) );
  NANDN U16122 ( .A(n5160), .B(\stack[1][40] ), .Z(n16445) );
  NANDN U16123 ( .A(n6108), .B(\stack[0][1] ), .Z(n16213) );
  ANDN U16124 ( .B(\stack[0][35] ), .A(n5292), .Z(n9118) );
  AND U16125 ( .A(n16446), .B(n16447), .Z(n9119) );
  NANDN U16126 ( .A(n9126), .B(n16448), .Z(n16446) );
  NANDN U16127 ( .A(n9125), .B(n9123), .Z(n16448) );
  XNOR U16128 ( .A(n16221), .B(n16449), .Z(n9123) );
  XNOR U16129 ( .A(n16222), .B(n16223), .Z(n16449) );
  AND U16130 ( .A(n16450), .B(n16451), .Z(n16223) );
  NANDN U16131 ( .A(n16452), .B(n16453), .Z(n16451) );
  NANDN U16132 ( .A(n16454), .B(n16455), .Z(n16450) );
  NANDN U16133 ( .A(n16453), .B(n16452), .Z(n16455) );
  ANDN U16134 ( .B(\stack[0][33] ), .A(n5316), .Z(n16222) );
  XNOR U16135 ( .A(n16228), .B(n16456), .Z(n16221) );
  XNOR U16136 ( .A(n16229), .B(n16230), .Z(n16456) );
  AND U16137 ( .A(n16457), .B(n16458), .Z(n16230) );
  NAND U16138 ( .A(n16459), .B(n16460), .Z(n16458) );
  NANDN U16139 ( .A(n16461), .B(n16462), .Z(n16457) );
  OR U16140 ( .A(n16459), .B(n16460), .Z(n16462) );
  ANDN U16141 ( .B(\stack[0][32] ), .A(n5340), .Z(n16229) );
  XNOR U16142 ( .A(n16235), .B(n16463), .Z(n16228) );
  XNOR U16143 ( .A(n16236), .B(n16237), .Z(n16463) );
  AND U16144 ( .A(n16464), .B(n16465), .Z(n16237) );
  NANDN U16145 ( .A(n16466), .B(n16467), .Z(n16465) );
  NANDN U16146 ( .A(n16468), .B(n16469), .Z(n16464) );
  NANDN U16147 ( .A(n16467), .B(n16466), .Z(n16469) );
  ANDN U16148 ( .B(\stack[0][31] ), .A(n5364), .Z(n16236) );
  XNOR U16149 ( .A(n16242), .B(n16470), .Z(n16235) );
  XNOR U16150 ( .A(n16243), .B(n16244), .Z(n16470) );
  AND U16151 ( .A(n16471), .B(n16472), .Z(n16244) );
  NAND U16152 ( .A(n16473), .B(n16474), .Z(n16472) );
  NANDN U16153 ( .A(n16475), .B(n16476), .Z(n16471) );
  OR U16154 ( .A(n16473), .B(n16474), .Z(n16476) );
  ANDN U16155 ( .B(\stack[0][30] ), .A(n5387), .Z(n16243) );
  XNOR U16156 ( .A(n16249), .B(n16477), .Z(n16242) );
  XNOR U16157 ( .A(n16250), .B(n16251), .Z(n16477) );
  AND U16158 ( .A(n16478), .B(n16479), .Z(n16251) );
  NANDN U16159 ( .A(n16480), .B(n16481), .Z(n16479) );
  NANDN U16160 ( .A(n16482), .B(n16483), .Z(n16478) );
  NANDN U16161 ( .A(n16481), .B(n16480), .Z(n16483) );
  ANDN U16162 ( .B(\stack[1][10] ), .A(n5854), .Z(n16250) );
  XNOR U16163 ( .A(n16256), .B(n16484), .Z(n16249) );
  XNOR U16164 ( .A(n16257), .B(n16258), .Z(n16484) );
  AND U16165 ( .A(n16485), .B(n16486), .Z(n16258) );
  NAND U16166 ( .A(n16487), .B(n16488), .Z(n16486) );
  NANDN U16167 ( .A(n16489), .B(n16490), .Z(n16485) );
  OR U16168 ( .A(n16487), .B(n16488), .Z(n16490) );
  ANDN U16169 ( .B(\stack[1][11] ), .A(n5830), .Z(n16257) );
  XNOR U16170 ( .A(n16263), .B(n16491), .Z(n16256) );
  XNOR U16171 ( .A(n16264), .B(n16265), .Z(n16491) );
  AND U16172 ( .A(n16492), .B(n16493), .Z(n16265) );
  NANDN U16173 ( .A(n16494), .B(n16495), .Z(n16493) );
  NANDN U16174 ( .A(n16496), .B(n16497), .Z(n16492) );
  NANDN U16175 ( .A(n16495), .B(n16494), .Z(n16497) );
  ANDN U16176 ( .B(\stack[1][12] ), .A(n5806), .Z(n16264) );
  XNOR U16177 ( .A(n16270), .B(n16498), .Z(n16263) );
  XNOR U16178 ( .A(n16271), .B(n16272), .Z(n16498) );
  AND U16179 ( .A(n16499), .B(n16500), .Z(n16272) );
  NAND U16180 ( .A(n16501), .B(n16502), .Z(n16500) );
  NANDN U16181 ( .A(n16503), .B(n16504), .Z(n16499) );
  OR U16182 ( .A(n16501), .B(n16502), .Z(n16504) );
  ANDN U16183 ( .B(\stack[1][13] ), .A(n5782), .Z(n16271) );
  XNOR U16184 ( .A(n16277), .B(n16505), .Z(n16270) );
  XNOR U16185 ( .A(n16278), .B(n16279), .Z(n16505) );
  AND U16186 ( .A(n16506), .B(n16507), .Z(n16279) );
  NANDN U16187 ( .A(n16508), .B(n16509), .Z(n16507) );
  NANDN U16188 ( .A(n16510), .B(n16511), .Z(n16506) );
  NANDN U16189 ( .A(n16509), .B(n16508), .Z(n16511) );
  ANDN U16190 ( .B(\stack[1][14] ), .A(n5758), .Z(n16278) );
  XNOR U16191 ( .A(n16284), .B(n16512), .Z(n16277) );
  XNOR U16192 ( .A(n16285), .B(n16286), .Z(n16512) );
  AND U16193 ( .A(n16513), .B(n16514), .Z(n16286) );
  NAND U16194 ( .A(n16515), .B(n16516), .Z(n16514) );
  NANDN U16195 ( .A(n16517), .B(n16518), .Z(n16513) );
  OR U16196 ( .A(n16515), .B(n16516), .Z(n16518) );
  ANDN U16197 ( .B(\stack[1][15] ), .A(n5734), .Z(n16285) );
  XNOR U16198 ( .A(n16291), .B(n16519), .Z(n16284) );
  XNOR U16199 ( .A(n16292), .B(n16293), .Z(n16519) );
  AND U16200 ( .A(n16520), .B(n16521), .Z(n16293) );
  NANDN U16201 ( .A(n16522), .B(n16523), .Z(n16521) );
  NANDN U16202 ( .A(n16524), .B(n16525), .Z(n16520) );
  NANDN U16203 ( .A(n16523), .B(n16522), .Z(n16525) );
  ANDN U16204 ( .B(\stack[1][16] ), .A(n5710), .Z(n16292) );
  XNOR U16205 ( .A(n16298), .B(n16526), .Z(n16291) );
  XNOR U16206 ( .A(n16299), .B(n16300), .Z(n16526) );
  AND U16207 ( .A(n16527), .B(n16528), .Z(n16300) );
  NAND U16208 ( .A(n16529), .B(n16530), .Z(n16528) );
  NANDN U16209 ( .A(n16531), .B(n16532), .Z(n16527) );
  OR U16210 ( .A(n16529), .B(n16530), .Z(n16532) );
  ANDN U16211 ( .B(\stack[1][17] ), .A(n5686), .Z(n16299) );
  XNOR U16212 ( .A(n16305), .B(n16533), .Z(n16298) );
  XNOR U16213 ( .A(n16306), .B(n16307), .Z(n16533) );
  AND U16214 ( .A(n16534), .B(n16535), .Z(n16307) );
  NANDN U16215 ( .A(n16536), .B(n16537), .Z(n16535) );
  NANDN U16216 ( .A(n16538), .B(n16539), .Z(n16534) );
  NANDN U16217 ( .A(n16537), .B(n16536), .Z(n16539) );
  ANDN U16218 ( .B(\stack[1][18] ), .A(n5662), .Z(n16306) );
  XNOR U16219 ( .A(n16312), .B(n16540), .Z(n16305) );
  XNOR U16220 ( .A(n16313), .B(n16314), .Z(n16540) );
  AND U16221 ( .A(n16541), .B(n16542), .Z(n16314) );
  NAND U16222 ( .A(n16543), .B(n16544), .Z(n16542) );
  NANDN U16223 ( .A(n16545), .B(n16546), .Z(n16541) );
  OR U16224 ( .A(n16543), .B(n16544), .Z(n16546) );
  ANDN U16225 ( .B(\stack[1][19] ), .A(n5638), .Z(n16313) );
  XNOR U16226 ( .A(n16319), .B(n16547), .Z(n16312) );
  XNOR U16227 ( .A(n16320), .B(n16321), .Z(n16547) );
  AND U16228 ( .A(n16548), .B(n16549), .Z(n16321) );
  NANDN U16229 ( .A(n16550), .B(n16551), .Z(n16549) );
  NANDN U16230 ( .A(n16552), .B(n16553), .Z(n16548) );
  NANDN U16231 ( .A(n16551), .B(n16550), .Z(n16553) );
  ANDN U16232 ( .B(\stack[1][20] ), .A(n5614), .Z(n16320) );
  XNOR U16233 ( .A(n16326), .B(n16554), .Z(n16319) );
  XNOR U16234 ( .A(n16327), .B(n16328), .Z(n16554) );
  AND U16235 ( .A(n16555), .B(n16556), .Z(n16328) );
  NAND U16236 ( .A(n16557), .B(n16558), .Z(n16556) );
  NANDN U16237 ( .A(n16559), .B(n16560), .Z(n16555) );
  OR U16238 ( .A(n16557), .B(n16558), .Z(n16560) );
  ANDN U16239 ( .B(\stack[1][21] ), .A(n5590), .Z(n16327) );
  XNOR U16240 ( .A(n16333), .B(n16561), .Z(n16326) );
  XNOR U16241 ( .A(n16334), .B(n16335), .Z(n16561) );
  AND U16242 ( .A(n16562), .B(n16563), .Z(n16335) );
  NANDN U16243 ( .A(n16564), .B(n16565), .Z(n16563) );
  NANDN U16244 ( .A(n16566), .B(n16567), .Z(n16562) );
  NANDN U16245 ( .A(n16565), .B(n16564), .Z(n16567) );
  ANDN U16246 ( .B(\stack[1][22] ), .A(n5566), .Z(n16334) );
  XNOR U16247 ( .A(n16340), .B(n16568), .Z(n16333) );
  XNOR U16248 ( .A(n16341), .B(n16342), .Z(n16568) );
  AND U16249 ( .A(n16569), .B(n16570), .Z(n16342) );
  NAND U16250 ( .A(n16571), .B(n16572), .Z(n16570) );
  NANDN U16251 ( .A(n16573), .B(n16574), .Z(n16569) );
  OR U16252 ( .A(n16571), .B(n16572), .Z(n16574) );
  ANDN U16253 ( .B(\stack[1][23] ), .A(n5542), .Z(n16341) );
  XNOR U16254 ( .A(n16347), .B(n16575), .Z(n16340) );
  XNOR U16255 ( .A(n16348), .B(n16349), .Z(n16575) );
  AND U16256 ( .A(n16576), .B(n16577), .Z(n16349) );
  NANDN U16257 ( .A(n16578), .B(n16579), .Z(n16577) );
  NANDN U16258 ( .A(n16580), .B(n16581), .Z(n16576) );
  NANDN U16259 ( .A(n16579), .B(n16578), .Z(n16581) );
  ANDN U16260 ( .B(\stack[1][24] ), .A(n5518), .Z(n16348) );
  XNOR U16261 ( .A(n16354), .B(n16582), .Z(n16347) );
  XNOR U16262 ( .A(n16355), .B(n16356), .Z(n16582) );
  AND U16263 ( .A(n16583), .B(n16584), .Z(n16356) );
  NAND U16264 ( .A(n16585), .B(n16586), .Z(n16584) );
  NANDN U16265 ( .A(n16587), .B(n16588), .Z(n16583) );
  OR U16266 ( .A(n16585), .B(n16586), .Z(n16588) );
  ANDN U16267 ( .B(\stack[1][25] ), .A(n5494), .Z(n16355) );
  XNOR U16268 ( .A(n16361), .B(n16589), .Z(n16354) );
  XNOR U16269 ( .A(n16362), .B(n16363), .Z(n16589) );
  AND U16270 ( .A(n16590), .B(n16591), .Z(n16363) );
  NANDN U16271 ( .A(n16592), .B(n16593), .Z(n16591) );
  NANDN U16272 ( .A(n16594), .B(n16595), .Z(n16590) );
  NANDN U16273 ( .A(n16593), .B(n16592), .Z(n16595) );
  ANDN U16274 ( .B(\stack[1][26] ), .A(n5470), .Z(n16362) );
  XNOR U16275 ( .A(n16368), .B(n16596), .Z(n16361) );
  XNOR U16276 ( .A(n16369), .B(n16370), .Z(n16596) );
  AND U16277 ( .A(n16597), .B(n16598), .Z(n16370) );
  NAND U16278 ( .A(n16599), .B(n16600), .Z(n16598) );
  NANDN U16279 ( .A(n16601), .B(n16602), .Z(n16597) );
  OR U16280 ( .A(n16599), .B(n16600), .Z(n16602) );
  ANDN U16281 ( .B(\stack[1][27] ), .A(n5446), .Z(n16369) );
  XNOR U16282 ( .A(n16375), .B(n16603), .Z(n16368) );
  XNOR U16283 ( .A(n16376), .B(n16377), .Z(n16603) );
  AND U16284 ( .A(n16604), .B(n16605), .Z(n16377) );
  NANDN U16285 ( .A(n16606), .B(n16607), .Z(n16605) );
  NANDN U16286 ( .A(n16608), .B(n16609), .Z(n16604) );
  NANDN U16287 ( .A(n16607), .B(n16606), .Z(n16609) );
  ANDN U16288 ( .B(\stack[1][28] ), .A(n5422), .Z(n16376) );
  XNOR U16289 ( .A(n16382), .B(n16610), .Z(n16375) );
  XNOR U16290 ( .A(n16383), .B(n16384), .Z(n16610) );
  AND U16291 ( .A(n16611), .B(n16612), .Z(n16384) );
  NAND U16292 ( .A(n16613), .B(n16614), .Z(n16612) );
  NANDN U16293 ( .A(n16615), .B(n16616), .Z(n16611) );
  OR U16294 ( .A(n16613), .B(n16614), .Z(n16616) );
  ANDN U16295 ( .B(\stack[1][29] ), .A(n5398), .Z(n16383) );
  XNOR U16296 ( .A(n16389), .B(n16617), .Z(n16382) );
  XNOR U16297 ( .A(n16390), .B(n16391), .Z(n16617) );
  AND U16298 ( .A(n16618), .B(n16619), .Z(n16391) );
  NANDN U16299 ( .A(n16620), .B(n16621), .Z(n16619) );
  NANDN U16300 ( .A(n16622), .B(n16623), .Z(n16618) );
  NANDN U16301 ( .A(n16621), .B(n16620), .Z(n16623) );
  ANDN U16302 ( .B(\stack[1][30] ), .A(n5374), .Z(n16390) );
  XNOR U16303 ( .A(n16396), .B(n16624), .Z(n16389) );
  XNOR U16304 ( .A(n16397), .B(n16398), .Z(n16624) );
  AND U16305 ( .A(n16625), .B(n16626), .Z(n16398) );
  NAND U16306 ( .A(n16627), .B(n16628), .Z(n16626) );
  NANDN U16307 ( .A(n16629), .B(n16630), .Z(n16625) );
  OR U16308 ( .A(n16627), .B(n16628), .Z(n16630) );
  ANDN U16309 ( .B(\stack[1][31] ), .A(n5350), .Z(n16397) );
  XNOR U16310 ( .A(n16403), .B(n16631), .Z(n16396) );
  XNOR U16311 ( .A(n16404), .B(n16405), .Z(n16631) );
  AND U16312 ( .A(n16632), .B(n16633), .Z(n16405) );
  NANDN U16313 ( .A(n16634), .B(n16635), .Z(n16633) );
  NANDN U16314 ( .A(n16636), .B(n16637), .Z(n16632) );
  NANDN U16315 ( .A(n16635), .B(n16634), .Z(n16637) );
  ANDN U16316 ( .B(\stack[1][32] ), .A(n5326), .Z(n16404) );
  XNOR U16317 ( .A(n16410), .B(n16638), .Z(n16403) );
  XNOR U16318 ( .A(n16411), .B(n16412), .Z(n16638) );
  AND U16319 ( .A(n16639), .B(n16640), .Z(n16412) );
  NAND U16320 ( .A(n16641), .B(n16642), .Z(n16640) );
  NANDN U16321 ( .A(n16643), .B(n16644), .Z(n16639) );
  OR U16322 ( .A(n16641), .B(n16642), .Z(n16644) );
  ANDN U16323 ( .B(\stack[1][33] ), .A(n5302), .Z(n16411) );
  XNOR U16324 ( .A(n16417), .B(n16645), .Z(n16410) );
  XNOR U16325 ( .A(n16418), .B(n16419), .Z(n16645) );
  AND U16326 ( .A(n16646), .B(n16647), .Z(n16419) );
  NANDN U16327 ( .A(n16648), .B(n16649), .Z(n16647) );
  NANDN U16328 ( .A(n16650), .B(n16651), .Z(n16646) );
  NANDN U16329 ( .A(n16649), .B(n16648), .Z(n16651) );
  ANDN U16330 ( .B(\stack[1][34] ), .A(n5278), .Z(n16418) );
  XNOR U16331 ( .A(n16424), .B(n16652), .Z(n16417) );
  XNOR U16332 ( .A(n16425), .B(n16426), .Z(n16652) );
  AND U16333 ( .A(n16653), .B(n16654), .Z(n16426) );
  NAND U16334 ( .A(n16655), .B(n16656), .Z(n16654) );
  NANDN U16335 ( .A(n16657), .B(n16658), .Z(n16653) );
  OR U16336 ( .A(n16655), .B(n16656), .Z(n16658) );
  ANDN U16337 ( .B(\stack[1][35] ), .A(n5254), .Z(n16425) );
  XNOR U16338 ( .A(n16431), .B(n16659), .Z(n16424) );
  XNOR U16339 ( .A(n16432), .B(n16433), .Z(n16659) );
  AND U16340 ( .A(n16660), .B(n16661), .Z(n16433) );
  NAND U16341 ( .A(n16662), .B(n16663), .Z(n16661) );
  NAND U16342 ( .A(n16664), .B(n16665), .Z(n16660) );
  OR U16343 ( .A(n16662), .B(n16663), .Z(n16664) );
  ANDN U16344 ( .B(\stack[1][36] ), .A(n5230), .Z(n16432) );
  XOR U16345 ( .A(n16438), .B(n16666), .Z(n16431) );
  XNOR U16346 ( .A(n16440), .B(n16441), .Z(n16666) );
  AND U16347 ( .A(\stack[1][37] ), .B(\stack[0][2] ), .Z(n16441) );
  ANDN U16348 ( .B(n16667), .A(n16668), .Z(n16440) );
  ANDN U16349 ( .B(\stack[0][0] ), .A(n6084), .Z(n16667) );
  XNOR U16350 ( .A(n16444), .B(n16669), .Z(n16438) );
  NANDN U16351 ( .A(n5160), .B(\stack[1][39] ), .Z(n16669) );
  NANDN U16352 ( .A(n6084), .B(\stack[0][1] ), .Z(n16444) );
  ANDN U16353 ( .B(\stack[1][5] ), .A(n5974), .Z(n9125) );
  AND U16354 ( .A(n16670), .B(n16671), .Z(n9126) );
  NANDN U16355 ( .A(n9130), .B(n9132), .Z(n16671) );
  NANDN U16356 ( .A(n9133), .B(n16672), .Z(n16670) );
  NANDN U16357 ( .A(n9132), .B(n9130), .Z(n16672) );
  XOR U16358 ( .A(n16452), .B(n16673), .Z(n9130) );
  XNOR U16359 ( .A(n16453), .B(n16454), .Z(n16673) );
  AND U16360 ( .A(n16674), .B(n16675), .Z(n16454) );
  NAND U16361 ( .A(n16676), .B(n16677), .Z(n16675) );
  NANDN U16362 ( .A(n16678), .B(n16679), .Z(n16674) );
  OR U16363 ( .A(n16676), .B(n16677), .Z(n16679) );
  ANDN U16364 ( .B(\stack[0][32] ), .A(n5316), .Z(n16453) );
  XNOR U16365 ( .A(n16459), .B(n16680), .Z(n16452) );
  XNOR U16366 ( .A(n16460), .B(n16461), .Z(n16680) );
  AND U16367 ( .A(n16681), .B(n16682), .Z(n16461) );
  NANDN U16368 ( .A(n16683), .B(n16684), .Z(n16682) );
  NANDN U16369 ( .A(n16685), .B(n16686), .Z(n16681) );
  NANDN U16370 ( .A(n16684), .B(n16683), .Z(n16686) );
  ANDN U16371 ( .B(\stack[0][31] ), .A(n5340), .Z(n16460) );
  XNOR U16372 ( .A(n16466), .B(n16687), .Z(n16459) );
  XNOR U16373 ( .A(n16467), .B(n16468), .Z(n16687) );
  AND U16374 ( .A(n16688), .B(n16689), .Z(n16468) );
  NAND U16375 ( .A(n16690), .B(n16691), .Z(n16689) );
  NANDN U16376 ( .A(n16692), .B(n16693), .Z(n16688) );
  OR U16377 ( .A(n16690), .B(n16691), .Z(n16693) );
  ANDN U16378 ( .B(\stack[0][30] ), .A(n5364), .Z(n16467) );
  XNOR U16379 ( .A(n16473), .B(n16694), .Z(n16466) );
  XNOR U16380 ( .A(n16474), .B(n16475), .Z(n16694) );
  AND U16381 ( .A(n16695), .B(n16696), .Z(n16475) );
  NANDN U16382 ( .A(n16697), .B(n16698), .Z(n16696) );
  NANDN U16383 ( .A(n16699), .B(n16700), .Z(n16695) );
  NANDN U16384 ( .A(n16698), .B(n16697), .Z(n16700) );
  ANDN U16385 ( .B(\stack[0][29] ), .A(n5387), .Z(n16474) );
  XNOR U16386 ( .A(n16480), .B(n16701), .Z(n16473) );
  XNOR U16387 ( .A(n16481), .B(n16482), .Z(n16701) );
  AND U16388 ( .A(n16702), .B(n16703), .Z(n16482) );
  NAND U16389 ( .A(n16704), .B(n16705), .Z(n16703) );
  NANDN U16390 ( .A(n16706), .B(n16707), .Z(n16702) );
  OR U16391 ( .A(n16704), .B(n16705), .Z(n16707) );
  ANDN U16392 ( .B(\stack[1][10] ), .A(n5830), .Z(n16481) );
  XNOR U16393 ( .A(n16487), .B(n16708), .Z(n16480) );
  XNOR U16394 ( .A(n16488), .B(n16489), .Z(n16708) );
  AND U16395 ( .A(n16709), .B(n16710), .Z(n16489) );
  NANDN U16396 ( .A(n16711), .B(n16712), .Z(n16710) );
  NANDN U16397 ( .A(n16713), .B(n16714), .Z(n16709) );
  NANDN U16398 ( .A(n16712), .B(n16711), .Z(n16714) );
  ANDN U16399 ( .B(\stack[1][11] ), .A(n5806), .Z(n16488) );
  XNOR U16400 ( .A(n16494), .B(n16715), .Z(n16487) );
  XNOR U16401 ( .A(n16495), .B(n16496), .Z(n16715) );
  AND U16402 ( .A(n16716), .B(n16717), .Z(n16496) );
  NAND U16403 ( .A(n16718), .B(n16719), .Z(n16717) );
  NANDN U16404 ( .A(n16720), .B(n16721), .Z(n16716) );
  OR U16405 ( .A(n16718), .B(n16719), .Z(n16721) );
  ANDN U16406 ( .B(\stack[1][12] ), .A(n5782), .Z(n16495) );
  XNOR U16407 ( .A(n16501), .B(n16722), .Z(n16494) );
  XNOR U16408 ( .A(n16502), .B(n16503), .Z(n16722) );
  AND U16409 ( .A(n16723), .B(n16724), .Z(n16503) );
  NANDN U16410 ( .A(n16725), .B(n16726), .Z(n16724) );
  NANDN U16411 ( .A(n16727), .B(n16728), .Z(n16723) );
  NANDN U16412 ( .A(n16726), .B(n16725), .Z(n16728) );
  ANDN U16413 ( .B(\stack[1][13] ), .A(n5758), .Z(n16502) );
  XNOR U16414 ( .A(n16508), .B(n16729), .Z(n16501) );
  XNOR U16415 ( .A(n16509), .B(n16510), .Z(n16729) );
  AND U16416 ( .A(n16730), .B(n16731), .Z(n16510) );
  NAND U16417 ( .A(n16732), .B(n16733), .Z(n16731) );
  NANDN U16418 ( .A(n16734), .B(n16735), .Z(n16730) );
  OR U16419 ( .A(n16732), .B(n16733), .Z(n16735) );
  ANDN U16420 ( .B(\stack[1][14] ), .A(n5734), .Z(n16509) );
  XNOR U16421 ( .A(n16515), .B(n16736), .Z(n16508) );
  XNOR U16422 ( .A(n16516), .B(n16517), .Z(n16736) );
  AND U16423 ( .A(n16737), .B(n16738), .Z(n16517) );
  NANDN U16424 ( .A(n16739), .B(n16740), .Z(n16738) );
  NANDN U16425 ( .A(n16741), .B(n16742), .Z(n16737) );
  NANDN U16426 ( .A(n16740), .B(n16739), .Z(n16742) );
  ANDN U16427 ( .B(\stack[1][15] ), .A(n5710), .Z(n16516) );
  XNOR U16428 ( .A(n16522), .B(n16743), .Z(n16515) );
  XNOR U16429 ( .A(n16523), .B(n16524), .Z(n16743) );
  AND U16430 ( .A(n16744), .B(n16745), .Z(n16524) );
  NAND U16431 ( .A(n16746), .B(n16747), .Z(n16745) );
  NANDN U16432 ( .A(n16748), .B(n16749), .Z(n16744) );
  OR U16433 ( .A(n16746), .B(n16747), .Z(n16749) );
  ANDN U16434 ( .B(\stack[1][16] ), .A(n5686), .Z(n16523) );
  XNOR U16435 ( .A(n16529), .B(n16750), .Z(n16522) );
  XNOR U16436 ( .A(n16530), .B(n16531), .Z(n16750) );
  AND U16437 ( .A(n16751), .B(n16752), .Z(n16531) );
  NANDN U16438 ( .A(n16753), .B(n16754), .Z(n16752) );
  NANDN U16439 ( .A(n16755), .B(n16756), .Z(n16751) );
  NANDN U16440 ( .A(n16754), .B(n16753), .Z(n16756) );
  ANDN U16441 ( .B(\stack[1][17] ), .A(n5662), .Z(n16530) );
  XNOR U16442 ( .A(n16536), .B(n16757), .Z(n16529) );
  XNOR U16443 ( .A(n16537), .B(n16538), .Z(n16757) );
  AND U16444 ( .A(n16758), .B(n16759), .Z(n16538) );
  NAND U16445 ( .A(n16760), .B(n16761), .Z(n16759) );
  NANDN U16446 ( .A(n16762), .B(n16763), .Z(n16758) );
  OR U16447 ( .A(n16760), .B(n16761), .Z(n16763) );
  ANDN U16448 ( .B(\stack[1][18] ), .A(n5638), .Z(n16537) );
  XNOR U16449 ( .A(n16543), .B(n16764), .Z(n16536) );
  XNOR U16450 ( .A(n16544), .B(n16545), .Z(n16764) );
  AND U16451 ( .A(n16765), .B(n16766), .Z(n16545) );
  NANDN U16452 ( .A(n16767), .B(n16768), .Z(n16766) );
  NANDN U16453 ( .A(n16769), .B(n16770), .Z(n16765) );
  NANDN U16454 ( .A(n16768), .B(n16767), .Z(n16770) );
  ANDN U16455 ( .B(\stack[1][19] ), .A(n5614), .Z(n16544) );
  XNOR U16456 ( .A(n16550), .B(n16771), .Z(n16543) );
  XNOR U16457 ( .A(n16551), .B(n16552), .Z(n16771) );
  AND U16458 ( .A(n16772), .B(n16773), .Z(n16552) );
  NAND U16459 ( .A(n16774), .B(n16775), .Z(n16773) );
  NANDN U16460 ( .A(n16776), .B(n16777), .Z(n16772) );
  OR U16461 ( .A(n16774), .B(n16775), .Z(n16777) );
  ANDN U16462 ( .B(\stack[1][20] ), .A(n5590), .Z(n16551) );
  XNOR U16463 ( .A(n16557), .B(n16778), .Z(n16550) );
  XNOR U16464 ( .A(n16558), .B(n16559), .Z(n16778) );
  AND U16465 ( .A(n16779), .B(n16780), .Z(n16559) );
  NANDN U16466 ( .A(n16781), .B(n16782), .Z(n16780) );
  NANDN U16467 ( .A(n16783), .B(n16784), .Z(n16779) );
  NANDN U16468 ( .A(n16782), .B(n16781), .Z(n16784) );
  ANDN U16469 ( .B(\stack[1][21] ), .A(n5566), .Z(n16558) );
  XNOR U16470 ( .A(n16564), .B(n16785), .Z(n16557) );
  XNOR U16471 ( .A(n16565), .B(n16566), .Z(n16785) );
  AND U16472 ( .A(n16786), .B(n16787), .Z(n16566) );
  NAND U16473 ( .A(n16788), .B(n16789), .Z(n16787) );
  NANDN U16474 ( .A(n16790), .B(n16791), .Z(n16786) );
  OR U16475 ( .A(n16788), .B(n16789), .Z(n16791) );
  ANDN U16476 ( .B(\stack[1][22] ), .A(n5542), .Z(n16565) );
  XNOR U16477 ( .A(n16571), .B(n16792), .Z(n16564) );
  XNOR U16478 ( .A(n16572), .B(n16573), .Z(n16792) );
  AND U16479 ( .A(n16793), .B(n16794), .Z(n16573) );
  NANDN U16480 ( .A(n16795), .B(n16796), .Z(n16794) );
  NANDN U16481 ( .A(n16797), .B(n16798), .Z(n16793) );
  NANDN U16482 ( .A(n16796), .B(n16795), .Z(n16798) );
  ANDN U16483 ( .B(\stack[1][23] ), .A(n5518), .Z(n16572) );
  XNOR U16484 ( .A(n16578), .B(n16799), .Z(n16571) );
  XNOR U16485 ( .A(n16579), .B(n16580), .Z(n16799) );
  AND U16486 ( .A(n16800), .B(n16801), .Z(n16580) );
  NAND U16487 ( .A(n16802), .B(n16803), .Z(n16801) );
  NANDN U16488 ( .A(n16804), .B(n16805), .Z(n16800) );
  OR U16489 ( .A(n16802), .B(n16803), .Z(n16805) );
  ANDN U16490 ( .B(\stack[1][24] ), .A(n5494), .Z(n16579) );
  XNOR U16491 ( .A(n16585), .B(n16806), .Z(n16578) );
  XNOR U16492 ( .A(n16586), .B(n16587), .Z(n16806) );
  AND U16493 ( .A(n16807), .B(n16808), .Z(n16587) );
  NANDN U16494 ( .A(n16809), .B(n16810), .Z(n16808) );
  NANDN U16495 ( .A(n16811), .B(n16812), .Z(n16807) );
  NANDN U16496 ( .A(n16810), .B(n16809), .Z(n16812) );
  ANDN U16497 ( .B(\stack[1][25] ), .A(n5470), .Z(n16586) );
  XNOR U16498 ( .A(n16592), .B(n16813), .Z(n16585) );
  XNOR U16499 ( .A(n16593), .B(n16594), .Z(n16813) );
  AND U16500 ( .A(n16814), .B(n16815), .Z(n16594) );
  NAND U16501 ( .A(n16816), .B(n16817), .Z(n16815) );
  NANDN U16502 ( .A(n16818), .B(n16819), .Z(n16814) );
  OR U16503 ( .A(n16816), .B(n16817), .Z(n16819) );
  ANDN U16504 ( .B(\stack[1][26] ), .A(n5446), .Z(n16593) );
  XNOR U16505 ( .A(n16599), .B(n16820), .Z(n16592) );
  XNOR U16506 ( .A(n16600), .B(n16601), .Z(n16820) );
  AND U16507 ( .A(n16821), .B(n16822), .Z(n16601) );
  NANDN U16508 ( .A(n16823), .B(n16824), .Z(n16822) );
  NANDN U16509 ( .A(n16825), .B(n16826), .Z(n16821) );
  NANDN U16510 ( .A(n16824), .B(n16823), .Z(n16826) );
  ANDN U16511 ( .B(\stack[1][27] ), .A(n5422), .Z(n16600) );
  XNOR U16512 ( .A(n16606), .B(n16827), .Z(n16599) );
  XNOR U16513 ( .A(n16607), .B(n16608), .Z(n16827) );
  AND U16514 ( .A(n16828), .B(n16829), .Z(n16608) );
  NAND U16515 ( .A(n16830), .B(n16831), .Z(n16829) );
  NANDN U16516 ( .A(n16832), .B(n16833), .Z(n16828) );
  OR U16517 ( .A(n16830), .B(n16831), .Z(n16833) );
  ANDN U16518 ( .B(\stack[1][28] ), .A(n5398), .Z(n16607) );
  XNOR U16519 ( .A(n16613), .B(n16834), .Z(n16606) );
  XNOR U16520 ( .A(n16614), .B(n16615), .Z(n16834) );
  AND U16521 ( .A(n16835), .B(n16836), .Z(n16615) );
  NANDN U16522 ( .A(n16837), .B(n16838), .Z(n16836) );
  NANDN U16523 ( .A(n16839), .B(n16840), .Z(n16835) );
  NANDN U16524 ( .A(n16838), .B(n16837), .Z(n16840) );
  ANDN U16525 ( .B(\stack[1][29] ), .A(n5374), .Z(n16614) );
  XNOR U16526 ( .A(n16620), .B(n16841), .Z(n16613) );
  XNOR U16527 ( .A(n16621), .B(n16622), .Z(n16841) );
  AND U16528 ( .A(n16842), .B(n16843), .Z(n16622) );
  NAND U16529 ( .A(n16844), .B(n16845), .Z(n16843) );
  NANDN U16530 ( .A(n16846), .B(n16847), .Z(n16842) );
  OR U16531 ( .A(n16844), .B(n16845), .Z(n16847) );
  ANDN U16532 ( .B(\stack[1][30] ), .A(n5350), .Z(n16621) );
  XNOR U16533 ( .A(n16627), .B(n16848), .Z(n16620) );
  XNOR U16534 ( .A(n16628), .B(n16629), .Z(n16848) );
  AND U16535 ( .A(n16849), .B(n16850), .Z(n16629) );
  NANDN U16536 ( .A(n16851), .B(n16852), .Z(n16850) );
  NANDN U16537 ( .A(n16853), .B(n16854), .Z(n16849) );
  NANDN U16538 ( .A(n16852), .B(n16851), .Z(n16854) );
  ANDN U16539 ( .B(\stack[1][31] ), .A(n5326), .Z(n16628) );
  XNOR U16540 ( .A(n16634), .B(n16855), .Z(n16627) );
  XNOR U16541 ( .A(n16635), .B(n16636), .Z(n16855) );
  AND U16542 ( .A(n16856), .B(n16857), .Z(n16636) );
  NAND U16543 ( .A(n16858), .B(n16859), .Z(n16857) );
  NANDN U16544 ( .A(n16860), .B(n16861), .Z(n16856) );
  OR U16545 ( .A(n16858), .B(n16859), .Z(n16861) );
  ANDN U16546 ( .B(\stack[1][32] ), .A(n5302), .Z(n16635) );
  XNOR U16547 ( .A(n16641), .B(n16862), .Z(n16634) );
  XNOR U16548 ( .A(n16642), .B(n16643), .Z(n16862) );
  AND U16549 ( .A(n16863), .B(n16864), .Z(n16643) );
  NANDN U16550 ( .A(n16865), .B(n16866), .Z(n16864) );
  NANDN U16551 ( .A(n16867), .B(n16868), .Z(n16863) );
  NANDN U16552 ( .A(n16866), .B(n16865), .Z(n16868) );
  ANDN U16553 ( .B(\stack[1][33] ), .A(n5278), .Z(n16642) );
  XNOR U16554 ( .A(n16648), .B(n16869), .Z(n16641) );
  XNOR U16555 ( .A(n16649), .B(n16650), .Z(n16869) );
  AND U16556 ( .A(n16870), .B(n16871), .Z(n16650) );
  NAND U16557 ( .A(n16872), .B(n16873), .Z(n16871) );
  NANDN U16558 ( .A(n16874), .B(n16875), .Z(n16870) );
  OR U16559 ( .A(n16872), .B(n16873), .Z(n16875) );
  ANDN U16560 ( .B(\stack[1][34] ), .A(n5254), .Z(n16649) );
  XNOR U16561 ( .A(n16655), .B(n16876), .Z(n16648) );
  XNOR U16562 ( .A(n16656), .B(n16657), .Z(n16876) );
  AND U16563 ( .A(n16877), .B(n16878), .Z(n16657) );
  NAND U16564 ( .A(n16879), .B(n16880), .Z(n16878) );
  NAND U16565 ( .A(n16881), .B(n16882), .Z(n16877) );
  OR U16566 ( .A(n16879), .B(n16880), .Z(n16881) );
  ANDN U16567 ( .B(\stack[1][35] ), .A(n5230), .Z(n16656) );
  XNOR U16568 ( .A(n16662), .B(n16883), .Z(n16655) );
  XNOR U16569 ( .A(n16663), .B(n16665), .Z(n16883) );
  ANDN U16570 ( .B(n16884), .A(n16885), .Z(n16665) );
  ANDN U16571 ( .B(\stack[0][0] ), .A(n6060), .Z(n16884) );
  ANDN U16572 ( .B(\stack[1][36] ), .A(n5206), .Z(n16663) );
  XOR U16573 ( .A(n16668), .B(n16886), .Z(n16662) );
  NANDN U16574 ( .A(n5160), .B(\stack[1][38] ), .Z(n16886) );
  NANDN U16575 ( .A(n6060), .B(\stack[0][1] ), .Z(n16668) );
  ANDN U16576 ( .B(\stack[0][33] ), .A(n5292), .Z(n9132) );
  AND U16577 ( .A(n16887), .B(n16888), .Z(n9133) );
  NANDN U16578 ( .A(n9140), .B(n16889), .Z(n16887) );
  NANDN U16579 ( .A(n9139), .B(n9137), .Z(n16889) );
  XNOR U16580 ( .A(n16676), .B(n16890), .Z(n9137) );
  XNOR U16581 ( .A(n16677), .B(n16678), .Z(n16890) );
  AND U16582 ( .A(n16891), .B(n16892), .Z(n16678) );
  NANDN U16583 ( .A(n16893), .B(n16894), .Z(n16892) );
  NANDN U16584 ( .A(n16895), .B(n16896), .Z(n16891) );
  NANDN U16585 ( .A(n16894), .B(n16893), .Z(n16896) );
  ANDN U16586 ( .B(\stack[0][31] ), .A(n5316), .Z(n16677) );
  XNOR U16587 ( .A(n16683), .B(n16897), .Z(n16676) );
  XNOR U16588 ( .A(n16684), .B(n16685), .Z(n16897) );
  AND U16589 ( .A(n16898), .B(n16899), .Z(n16685) );
  NAND U16590 ( .A(n16900), .B(n16901), .Z(n16899) );
  NANDN U16591 ( .A(n16902), .B(n16903), .Z(n16898) );
  OR U16592 ( .A(n16900), .B(n16901), .Z(n16903) );
  ANDN U16593 ( .B(\stack[0][30] ), .A(n5340), .Z(n16684) );
  XNOR U16594 ( .A(n16690), .B(n16904), .Z(n16683) );
  XNOR U16595 ( .A(n16691), .B(n16692), .Z(n16904) );
  AND U16596 ( .A(n16905), .B(n16906), .Z(n16692) );
  NANDN U16597 ( .A(n16907), .B(n16908), .Z(n16906) );
  NANDN U16598 ( .A(n16909), .B(n16910), .Z(n16905) );
  NANDN U16599 ( .A(n16908), .B(n16907), .Z(n16910) );
  ANDN U16600 ( .B(\stack[0][29] ), .A(n5364), .Z(n16691) );
  XNOR U16601 ( .A(n16697), .B(n16911), .Z(n16690) );
  XNOR U16602 ( .A(n16698), .B(n16699), .Z(n16911) );
  AND U16603 ( .A(n16912), .B(n16913), .Z(n16699) );
  NAND U16604 ( .A(n16914), .B(n16915), .Z(n16913) );
  NANDN U16605 ( .A(n16916), .B(n16917), .Z(n16912) );
  OR U16606 ( .A(n16914), .B(n16915), .Z(n16917) );
  ANDN U16607 ( .B(\stack[0][28] ), .A(n5387), .Z(n16698) );
  XNOR U16608 ( .A(n16704), .B(n16918), .Z(n16697) );
  XNOR U16609 ( .A(n16705), .B(n16706), .Z(n16918) );
  AND U16610 ( .A(n16919), .B(n16920), .Z(n16706) );
  NANDN U16611 ( .A(n16921), .B(n16922), .Z(n16920) );
  NANDN U16612 ( .A(n16923), .B(n16924), .Z(n16919) );
  NANDN U16613 ( .A(n16922), .B(n16921), .Z(n16924) );
  ANDN U16614 ( .B(\stack[1][10] ), .A(n5806), .Z(n16705) );
  XNOR U16615 ( .A(n16711), .B(n16925), .Z(n16704) );
  XNOR U16616 ( .A(n16712), .B(n16713), .Z(n16925) );
  AND U16617 ( .A(n16926), .B(n16927), .Z(n16713) );
  NAND U16618 ( .A(n16928), .B(n16929), .Z(n16927) );
  NANDN U16619 ( .A(n16930), .B(n16931), .Z(n16926) );
  OR U16620 ( .A(n16928), .B(n16929), .Z(n16931) );
  ANDN U16621 ( .B(\stack[1][11] ), .A(n5782), .Z(n16712) );
  XNOR U16622 ( .A(n16718), .B(n16932), .Z(n16711) );
  XNOR U16623 ( .A(n16719), .B(n16720), .Z(n16932) );
  AND U16624 ( .A(n16933), .B(n16934), .Z(n16720) );
  NANDN U16625 ( .A(n16935), .B(n16936), .Z(n16934) );
  NANDN U16626 ( .A(n16937), .B(n16938), .Z(n16933) );
  NANDN U16627 ( .A(n16936), .B(n16935), .Z(n16938) );
  ANDN U16628 ( .B(\stack[1][12] ), .A(n5758), .Z(n16719) );
  XNOR U16629 ( .A(n16725), .B(n16939), .Z(n16718) );
  XNOR U16630 ( .A(n16726), .B(n16727), .Z(n16939) );
  AND U16631 ( .A(n16940), .B(n16941), .Z(n16727) );
  NAND U16632 ( .A(n16942), .B(n16943), .Z(n16941) );
  NANDN U16633 ( .A(n16944), .B(n16945), .Z(n16940) );
  OR U16634 ( .A(n16942), .B(n16943), .Z(n16945) );
  ANDN U16635 ( .B(\stack[1][13] ), .A(n5734), .Z(n16726) );
  XNOR U16636 ( .A(n16732), .B(n16946), .Z(n16725) );
  XNOR U16637 ( .A(n16733), .B(n16734), .Z(n16946) );
  AND U16638 ( .A(n16947), .B(n16948), .Z(n16734) );
  NANDN U16639 ( .A(n16949), .B(n16950), .Z(n16948) );
  NANDN U16640 ( .A(n16951), .B(n16952), .Z(n16947) );
  NANDN U16641 ( .A(n16950), .B(n16949), .Z(n16952) );
  ANDN U16642 ( .B(\stack[1][14] ), .A(n5710), .Z(n16733) );
  XNOR U16643 ( .A(n16739), .B(n16953), .Z(n16732) );
  XNOR U16644 ( .A(n16740), .B(n16741), .Z(n16953) );
  AND U16645 ( .A(n16954), .B(n16955), .Z(n16741) );
  NAND U16646 ( .A(n16956), .B(n16957), .Z(n16955) );
  NANDN U16647 ( .A(n16958), .B(n16959), .Z(n16954) );
  OR U16648 ( .A(n16956), .B(n16957), .Z(n16959) );
  ANDN U16649 ( .B(\stack[1][15] ), .A(n5686), .Z(n16740) );
  XNOR U16650 ( .A(n16746), .B(n16960), .Z(n16739) );
  XNOR U16651 ( .A(n16747), .B(n16748), .Z(n16960) );
  AND U16652 ( .A(n16961), .B(n16962), .Z(n16748) );
  NANDN U16653 ( .A(n16963), .B(n16964), .Z(n16962) );
  NANDN U16654 ( .A(n16965), .B(n16966), .Z(n16961) );
  NANDN U16655 ( .A(n16964), .B(n16963), .Z(n16966) );
  ANDN U16656 ( .B(\stack[1][16] ), .A(n5662), .Z(n16747) );
  XNOR U16657 ( .A(n16753), .B(n16967), .Z(n16746) );
  XNOR U16658 ( .A(n16754), .B(n16755), .Z(n16967) );
  AND U16659 ( .A(n16968), .B(n16969), .Z(n16755) );
  NAND U16660 ( .A(n16970), .B(n16971), .Z(n16969) );
  NANDN U16661 ( .A(n16972), .B(n16973), .Z(n16968) );
  OR U16662 ( .A(n16970), .B(n16971), .Z(n16973) );
  ANDN U16663 ( .B(\stack[1][17] ), .A(n5638), .Z(n16754) );
  XNOR U16664 ( .A(n16760), .B(n16974), .Z(n16753) );
  XNOR U16665 ( .A(n16761), .B(n16762), .Z(n16974) );
  AND U16666 ( .A(n16975), .B(n16976), .Z(n16762) );
  NANDN U16667 ( .A(n16977), .B(n16978), .Z(n16976) );
  NANDN U16668 ( .A(n16979), .B(n16980), .Z(n16975) );
  NANDN U16669 ( .A(n16978), .B(n16977), .Z(n16980) );
  ANDN U16670 ( .B(\stack[1][18] ), .A(n5614), .Z(n16761) );
  XNOR U16671 ( .A(n16767), .B(n16981), .Z(n16760) );
  XNOR U16672 ( .A(n16768), .B(n16769), .Z(n16981) );
  AND U16673 ( .A(n16982), .B(n16983), .Z(n16769) );
  NAND U16674 ( .A(n16984), .B(n16985), .Z(n16983) );
  NANDN U16675 ( .A(n16986), .B(n16987), .Z(n16982) );
  OR U16676 ( .A(n16984), .B(n16985), .Z(n16987) );
  ANDN U16677 ( .B(\stack[1][19] ), .A(n5590), .Z(n16768) );
  XNOR U16678 ( .A(n16774), .B(n16988), .Z(n16767) );
  XNOR U16679 ( .A(n16775), .B(n16776), .Z(n16988) );
  AND U16680 ( .A(n16989), .B(n16990), .Z(n16776) );
  NANDN U16681 ( .A(n16991), .B(n16992), .Z(n16990) );
  NANDN U16682 ( .A(n16993), .B(n16994), .Z(n16989) );
  NANDN U16683 ( .A(n16992), .B(n16991), .Z(n16994) );
  ANDN U16684 ( .B(\stack[1][20] ), .A(n5566), .Z(n16775) );
  XNOR U16685 ( .A(n16781), .B(n16995), .Z(n16774) );
  XNOR U16686 ( .A(n16782), .B(n16783), .Z(n16995) );
  AND U16687 ( .A(n16996), .B(n16997), .Z(n16783) );
  NAND U16688 ( .A(n16998), .B(n16999), .Z(n16997) );
  NANDN U16689 ( .A(n17000), .B(n17001), .Z(n16996) );
  OR U16690 ( .A(n16998), .B(n16999), .Z(n17001) );
  ANDN U16691 ( .B(\stack[1][21] ), .A(n5542), .Z(n16782) );
  XNOR U16692 ( .A(n16788), .B(n17002), .Z(n16781) );
  XNOR U16693 ( .A(n16789), .B(n16790), .Z(n17002) );
  AND U16694 ( .A(n17003), .B(n17004), .Z(n16790) );
  NANDN U16695 ( .A(n17005), .B(n17006), .Z(n17004) );
  NANDN U16696 ( .A(n17007), .B(n17008), .Z(n17003) );
  NANDN U16697 ( .A(n17006), .B(n17005), .Z(n17008) );
  ANDN U16698 ( .B(\stack[1][22] ), .A(n5518), .Z(n16789) );
  XNOR U16699 ( .A(n16795), .B(n17009), .Z(n16788) );
  XNOR U16700 ( .A(n16796), .B(n16797), .Z(n17009) );
  AND U16701 ( .A(n17010), .B(n17011), .Z(n16797) );
  NAND U16702 ( .A(n17012), .B(n17013), .Z(n17011) );
  NANDN U16703 ( .A(n17014), .B(n17015), .Z(n17010) );
  OR U16704 ( .A(n17012), .B(n17013), .Z(n17015) );
  ANDN U16705 ( .B(\stack[1][23] ), .A(n5494), .Z(n16796) );
  XNOR U16706 ( .A(n16802), .B(n17016), .Z(n16795) );
  XNOR U16707 ( .A(n16803), .B(n16804), .Z(n17016) );
  AND U16708 ( .A(n17017), .B(n17018), .Z(n16804) );
  NANDN U16709 ( .A(n17019), .B(n17020), .Z(n17018) );
  NANDN U16710 ( .A(n17021), .B(n17022), .Z(n17017) );
  NANDN U16711 ( .A(n17020), .B(n17019), .Z(n17022) );
  ANDN U16712 ( .B(\stack[1][24] ), .A(n5470), .Z(n16803) );
  XNOR U16713 ( .A(n16809), .B(n17023), .Z(n16802) );
  XNOR U16714 ( .A(n16810), .B(n16811), .Z(n17023) );
  AND U16715 ( .A(n17024), .B(n17025), .Z(n16811) );
  NAND U16716 ( .A(n17026), .B(n17027), .Z(n17025) );
  NANDN U16717 ( .A(n17028), .B(n17029), .Z(n17024) );
  OR U16718 ( .A(n17026), .B(n17027), .Z(n17029) );
  ANDN U16719 ( .B(\stack[1][25] ), .A(n5446), .Z(n16810) );
  XNOR U16720 ( .A(n16816), .B(n17030), .Z(n16809) );
  XNOR U16721 ( .A(n16817), .B(n16818), .Z(n17030) );
  AND U16722 ( .A(n17031), .B(n17032), .Z(n16818) );
  NANDN U16723 ( .A(n17033), .B(n17034), .Z(n17032) );
  NANDN U16724 ( .A(n17035), .B(n17036), .Z(n17031) );
  NANDN U16725 ( .A(n17034), .B(n17033), .Z(n17036) );
  ANDN U16726 ( .B(\stack[1][26] ), .A(n5422), .Z(n16817) );
  XNOR U16727 ( .A(n16823), .B(n17037), .Z(n16816) );
  XNOR U16728 ( .A(n16824), .B(n16825), .Z(n17037) );
  AND U16729 ( .A(n17038), .B(n17039), .Z(n16825) );
  NAND U16730 ( .A(n17040), .B(n17041), .Z(n17039) );
  NANDN U16731 ( .A(n17042), .B(n17043), .Z(n17038) );
  OR U16732 ( .A(n17040), .B(n17041), .Z(n17043) );
  ANDN U16733 ( .B(\stack[1][27] ), .A(n5398), .Z(n16824) );
  XNOR U16734 ( .A(n16830), .B(n17044), .Z(n16823) );
  XNOR U16735 ( .A(n16831), .B(n16832), .Z(n17044) );
  AND U16736 ( .A(n17045), .B(n17046), .Z(n16832) );
  NANDN U16737 ( .A(n17047), .B(n17048), .Z(n17046) );
  NANDN U16738 ( .A(n17049), .B(n17050), .Z(n17045) );
  NANDN U16739 ( .A(n17048), .B(n17047), .Z(n17050) );
  ANDN U16740 ( .B(\stack[1][28] ), .A(n5374), .Z(n16831) );
  XNOR U16741 ( .A(n16837), .B(n17051), .Z(n16830) );
  XNOR U16742 ( .A(n16838), .B(n16839), .Z(n17051) );
  AND U16743 ( .A(n17052), .B(n17053), .Z(n16839) );
  NAND U16744 ( .A(n17054), .B(n17055), .Z(n17053) );
  NANDN U16745 ( .A(n17056), .B(n17057), .Z(n17052) );
  OR U16746 ( .A(n17054), .B(n17055), .Z(n17057) );
  ANDN U16747 ( .B(\stack[1][29] ), .A(n5350), .Z(n16838) );
  XNOR U16748 ( .A(n16844), .B(n17058), .Z(n16837) );
  XNOR U16749 ( .A(n16845), .B(n16846), .Z(n17058) );
  AND U16750 ( .A(n17059), .B(n17060), .Z(n16846) );
  NANDN U16751 ( .A(n17061), .B(n17062), .Z(n17060) );
  NANDN U16752 ( .A(n17063), .B(n17064), .Z(n17059) );
  NANDN U16753 ( .A(n17062), .B(n17061), .Z(n17064) );
  ANDN U16754 ( .B(\stack[1][30] ), .A(n5326), .Z(n16845) );
  XNOR U16755 ( .A(n16851), .B(n17065), .Z(n16844) );
  XNOR U16756 ( .A(n16852), .B(n16853), .Z(n17065) );
  AND U16757 ( .A(n17066), .B(n17067), .Z(n16853) );
  NAND U16758 ( .A(n17068), .B(n17069), .Z(n17067) );
  NANDN U16759 ( .A(n17070), .B(n17071), .Z(n17066) );
  OR U16760 ( .A(n17068), .B(n17069), .Z(n17071) );
  ANDN U16761 ( .B(\stack[1][31] ), .A(n5302), .Z(n16852) );
  XNOR U16762 ( .A(n16858), .B(n17072), .Z(n16851) );
  XNOR U16763 ( .A(n16859), .B(n16860), .Z(n17072) );
  AND U16764 ( .A(n17073), .B(n17074), .Z(n16860) );
  NANDN U16765 ( .A(n17075), .B(n17076), .Z(n17074) );
  NANDN U16766 ( .A(n17077), .B(n17078), .Z(n17073) );
  NANDN U16767 ( .A(n17076), .B(n17075), .Z(n17078) );
  ANDN U16768 ( .B(\stack[1][32] ), .A(n5278), .Z(n16859) );
  XNOR U16769 ( .A(n16865), .B(n17079), .Z(n16858) );
  XNOR U16770 ( .A(n16866), .B(n16867), .Z(n17079) );
  AND U16771 ( .A(n17080), .B(n17081), .Z(n16867) );
  NAND U16772 ( .A(n17082), .B(n17083), .Z(n17081) );
  NANDN U16773 ( .A(n17084), .B(n17085), .Z(n17080) );
  OR U16774 ( .A(n17082), .B(n17083), .Z(n17085) );
  ANDN U16775 ( .B(\stack[1][33] ), .A(n5254), .Z(n16866) );
  XNOR U16776 ( .A(n16872), .B(n17086), .Z(n16865) );
  XNOR U16777 ( .A(n16873), .B(n16874), .Z(n17086) );
  AND U16778 ( .A(n17087), .B(n17088), .Z(n16874) );
  NAND U16779 ( .A(n17089), .B(n17090), .Z(n17088) );
  NAND U16780 ( .A(n17091), .B(n17092), .Z(n17087) );
  OR U16781 ( .A(n17089), .B(n17090), .Z(n17091) );
  ANDN U16782 ( .B(\stack[1][34] ), .A(n5230), .Z(n16873) );
  XNOR U16783 ( .A(n16879), .B(n17093), .Z(n16872) );
  XNOR U16784 ( .A(n16880), .B(n16882), .Z(n17093) );
  ANDN U16785 ( .B(n17094), .A(n17095), .Z(n16882) );
  ANDN U16786 ( .B(\stack[0][0] ), .A(n6036), .Z(n17094) );
  ANDN U16787 ( .B(\stack[1][35] ), .A(n5206), .Z(n16880) );
  XOR U16788 ( .A(n16885), .B(n17096), .Z(n16879) );
  NANDN U16789 ( .A(n5160), .B(\stack[1][37] ), .Z(n17096) );
  NANDN U16790 ( .A(n6036), .B(\stack[0][1] ), .Z(n16885) );
  ANDN U16791 ( .B(\stack[1][5] ), .A(n5926), .Z(n9139) );
  AND U16792 ( .A(n17097), .B(n17098), .Z(n9140) );
  NANDN U16793 ( .A(n9144), .B(n9146), .Z(n17098) );
  NANDN U16794 ( .A(n9147), .B(n17099), .Z(n17097) );
  NANDN U16795 ( .A(n9146), .B(n9144), .Z(n17099) );
  XOR U16796 ( .A(n16893), .B(n17100), .Z(n9144) );
  XNOR U16797 ( .A(n16894), .B(n16895), .Z(n17100) );
  AND U16798 ( .A(n17101), .B(n17102), .Z(n16895) );
  NAND U16799 ( .A(n17103), .B(n17104), .Z(n17102) );
  NANDN U16800 ( .A(n17105), .B(n17106), .Z(n17101) );
  OR U16801 ( .A(n17103), .B(n17104), .Z(n17106) );
  ANDN U16802 ( .B(\stack[0][30] ), .A(n5316), .Z(n16894) );
  XNOR U16803 ( .A(n16900), .B(n17107), .Z(n16893) );
  XNOR U16804 ( .A(n16901), .B(n16902), .Z(n17107) );
  AND U16805 ( .A(n17108), .B(n17109), .Z(n16902) );
  NANDN U16806 ( .A(n17110), .B(n17111), .Z(n17109) );
  NANDN U16807 ( .A(n17112), .B(n17113), .Z(n17108) );
  NANDN U16808 ( .A(n17111), .B(n17110), .Z(n17113) );
  ANDN U16809 ( .B(\stack[0][29] ), .A(n5340), .Z(n16901) );
  XNOR U16810 ( .A(n16907), .B(n17114), .Z(n16900) );
  XNOR U16811 ( .A(n16908), .B(n16909), .Z(n17114) );
  AND U16812 ( .A(n17115), .B(n17116), .Z(n16909) );
  NAND U16813 ( .A(n17117), .B(n17118), .Z(n17116) );
  NANDN U16814 ( .A(n17119), .B(n17120), .Z(n17115) );
  OR U16815 ( .A(n17117), .B(n17118), .Z(n17120) );
  ANDN U16816 ( .B(\stack[0][28] ), .A(n5364), .Z(n16908) );
  XNOR U16817 ( .A(n16914), .B(n17121), .Z(n16907) );
  XNOR U16818 ( .A(n16915), .B(n16916), .Z(n17121) );
  AND U16819 ( .A(n17122), .B(n17123), .Z(n16916) );
  NANDN U16820 ( .A(n17124), .B(n17125), .Z(n17123) );
  NANDN U16821 ( .A(n17126), .B(n17127), .Z(n17122) );
  NANDN U16822 ( .A(n17125), .B(n17124), .Z(n17127) );
  ANDN U16823 ( .B(\stack[0][27] ), .A(n5387), .Z(n16915) );
  XNOR U16824 ( .A(n16921), .B(n17128), .Z(n16914) );
  XNOR U16825 ( .A(n16922), .B(n16923), .Z(n17128) );
  AND U16826 ( .A(n17129), .B(n17130), .Z(n16923) );
  NAND U16827 ( .A(n17131), .B(n17132), .Z(n17130) );
  NANDN U16828 ( .A(n17133), .B(n17134), .Z(n17129) );
  OR U16829 ( .A(n17131), .B(n17132), .Z(n17134) );
  ANDN U16830 ( .B(\stack[1][10] ), .A(n5782), .Z(n16922) );
  XNOR U16831 ( .A(n16928), .B(n17135), .Z(n16921) );
  XNOR U16832 ( .A(n16929), .B(n16930), .Z(n17135) );
  AND U16833 ( .A(n17136), .B(n17137), .Z(n16930) );
  NANDN U16834 ( .A(n17138), .B(n17139), .Z(n17137) );
  NANDN U16835 ( .A(n17140), .B(n17141), .Z(n17136) );
  NANDN U16836 ( .A(n17139), .B(n17138), .Z(n17141) );
  ANDN U16837 ( .B(\stack[1][11] ), .A(n5758), .Z(n16929) );
  XNOR U16838 ( .A(n16935), .B(n17142), .Z(n16928) );
  XNOR U16839 ( .A(n16936), .B(n16937), .Z(n17142) );
  AND U16840 ( .A(n17143), .B(n17144), .Z(n16937) );
  NAND U16841 ( .A(n17145), .B(n17146), .Z(n17144) );
  NANDN U16842 ( .A(n17147), .B(n17148), .Z(n17143) );
  OR U16843 ( .A(n17145), .B(n17146), .Z(n17148) );
  ANDN U16844 ( .B(\stack[1][12] ), .A(n5734), .Z(n16936) );
  XNOR U16845 ( .A(n16942), .B(n17149), .Z(n16935) );
  XNOR U16846 ( .A(n16943), .B(n16944), .Z(n17149) );
  AND U16847 ( .A(n17150), .B(n17151), .Z(n16944) );
  NANDN U16848 ( .A(n17152), .B(n17153), .Z(n17151) );
  NANDN U16849 ( .A(n17154), .B(n17155), .Z(n17150) );
  NANDN U16850 ( .A(n17153), .B(n17152), .Z(n17155) );
  ANDN U16851 ( .B(\stack[1][13] ), .A(n5710), .Z(n16943) );
  XNOR U16852 ( .A(n16949), .B(n17156), .Z(n16942) );
  XNOR U16853 ( .A(n16950), .B(n16951), .Z(n17156) );
  AND U16854 ( .A(n17157), .B(n17158), .Z(n16951) );
  NAND U16855 ( .A(n17159), .B(n17160), .Z(n17158) );
  NANDN U16856 ( .A(n17161), .B(n17162), .Z(n17157) );
  OR U16857 ( .A(n17159), .B(n17160), .Z(n17162) );
  ANDN U16858 ( .B(\stack[1][14] ), .A(n5686), .Z(n16950) );
  XNOR U16859 ( .A(n16956), .B(n17163), .Z(n16949) );
  XNOR U16860 ( .A(n16957), .B(n16958), .Z(n17163) );
  AND U16861 ( .A(n17164), .B(n17165), .Z(n16958) );
  NANDN U16862 ( .A(n17166), .B(n17167), .Z(n17165) );
  NANDN U16863 ( .A(n17168), .B(n17169), .Z(n17164) );
  NANDN U16864 ( .A(n17167), .B(n17166), .Z(n17169) );
  ANDN U16865 ( .B(\stack[1][15] ), .A(n5662), .Z(n16957) );
  XNOR U16866 ( .A(n16963), .B(n17170), .Z(n16956) );
  XNOR U16867 ( .A(n16964), .B(n16965), .Z(n17170) );
  AND U16868 ( .A(n17171), .B(n17172), .Z(n16965) );
  NAND U16869 ( .A(n17173), .B(n17174), .Z(n17172) );
  NANDN U16870 ( .A(n17175), .B(n17176), .Z(n17171) );
  OR U16871 ( .A(n17173), .B(n17174), .Z(n17176) );
  ANDN U16872 ( .B(\stack[1][16] ), .A(n5638), .Z(n16964) );
  XNOR U16873 ( .A(n16970), .B(n17177), .Z(n16963) );
  XNOR U16874 ( .A(n16971), .B(n16972), .Z(n17177) );
  AND U16875 ( .A(n17178), .B(n17179), .Z(n16972) );
  NANDN U16876 ( .A(n17180), .B(n17181), .Z(n17179) );
  NANDN U16877 ( .A(n17182), .B(n17183), .Z(n17178) );
  NANDN U16878 ( .A(n17181), .B(n17180), .Z(n17183) );
  ANDN U16879 ( .B(\stack[1][17] ), .A(n5614), .Z(n16971) );
  XNOR U16880 ( .A(n16977), .B(n17184), .Z(n16970) );
  XNOR U16881 ( .A(n16978), .B(n16979), .Z(n17184) );
  AND U16882 ( .A(n17185), .B(n17186), .Z(n16979) );
  NAND U16883 ( .A(n17187), .B(n17188), .Z(n17186) );
  NANDN U16884 ( .A(n17189), .B(n17190), .Z(n17185) );
  OR U16885 ( .A(n17187), .B(n17188), .Z(n17190) );
  ANDN U16886 ( .B(\stack[1][18] ), .A(n5590), .Z(n16978) );
  XNOR U16887 ( .A(n16984), .B(n17191), .Z(n16977) );
  XNOR U16888 ( .A(n16985), .B(n16986), .Z(n17191) );
  AND U16889 ( .A(n17192), .B(n17193), .Z(n16986) );
  NANDN U16890 ( .A(n17194), .B(n17195), .Z(n17193) );
  NANDN U16891 ( .A(n17196), .B(n17197), .Z(n17192) );
  NANDN U16892 ( .A(n17195), .B(n17194), .Z(n17197) );
  ANDN U16893 ( .B(\stack[1][19] ), .A(n5566), .Z(n16985) );
  XNOR U16894 ( .A(n16991), .B(n17198), .Z(n16984) );
  XNOR U16895 ( .A(n16992), .B(n16993), .Z(n17198) );
  AND U16896 ( .A(n17199), .B(n17200), .Z(n16993) );
  NAND U16897 ( .A(n17201), .B(n17202), .Z(n17200) );
  NANDN U16898 ( .A(n17203), .B(n17204), .Z(n17199) );
  OR U16899 ( .A(n17201), .B(n17202), .Z(n17204) );
  ANDN U16900 ( .B(\stack[1][20] ), .A(n5542), .Z(n16992) );
  XNOR U16901 ( .A(n16998), .B(n17205), .Z(n16991) );
  XNOR U16902 ( .A(n16999), .B(n17000), .Z(n17205) );
  AND U16903 ( .A(n17206), .B(n17207), .Z(n17000) );
  NANDN U16904 ( .A(n17208), .B(n17209), .Z(n17207) );
  NANDN U16905 ( .A(n17210), .B(n17211), .Z(n17206) );
  NANDN U16906 ( .A(n17209), .B(n17208), .Z(n17211) );
  ANDN U16907 ( .B(\stack[1][21] ), .A(n5518), .Z(n16999) );
  XNOR U16908 ( .A(n17005), .B(n17212), .Z(n16998) );
  XNOR U16909 ( .A(n17006), .B(n17007), .Z(n17212) );
  AND U16910 ( .A(n17213), .B(n17214), .Z(n17007) );
  NAND U16911 ( .A(n17215), .B(n17216), .Z(n17214) );
  NANDN U16912 ( .A(n17217), .B(n17218), .Z(n17213) );
  OR U16913 ( .A(n17215), .B(n17216), .Z(n17218) );
  ANDN U16914 ( .B(\stack[1][22] ), .A(n5494), .Z(n17006) );
  XNOR U16915 ( .A(n17012), .B(n17219), .Z(n17005) );
  XNOR U16916 ( .A(n17013), .B(n17014), .Z(n17219) );
  AND U16917 ( .A(n17220), .B(n17221), .Z(n17014) );
  NANDN U16918 ( .A(n17222), .B(n17223), .Z(n17221) );
  NANDN U16919 ( .A(n17224), .B(n17225), .Z(n17220) );
  NANDN U16920 ( .A(n17223), .B(n17222), .Z(n17225) );
  ANDN U16921 ( .B(\stack[1][23] ), .A(n5470), .Z(n17013) );
  XNOR U16922 ( .A(n17019), .B(n17226), .Z(n17012) );
  XNOR U16923 ( .A(n17020), .B(n17021), .Z(n17226) );
  AND U16924 ( .A(n17227), .B(n17228), .Z(n17021) );
  NAND U16925 ( .A(n17229), .B(n17230), .Z(n17228) );
  NANDN U16926 ( .A(n17231), .B(n17232), .Z(n17227) );
  OR U16927 ( .A(n17229), .B(n17230), .Z(n17232) );
  ANDN U16928 ( .B(\stack[1][24] ), .A(n5446), .Z(n17020) );
  XNOR U16929 ( .A(n17026), .B(n17233), .Z(n17019) );
  XNOR U16930 ( .A(n17027), .B(n17028), .Z(n17233) );
  AND U16931 ( .A(n17234), .B(n17235), .Z(n17028) );
  NANDN U16932 ( .A(n17236), .B(n17237), .Z(n17235) );
  NANDN U16933 ( .A(n17238), .B(n17239), .Z(n17234) );
  NANDN U16934 ( .A(n17237), .B(n17236), .Z(n17239) );
  ANDN U16935 ( .B(\stack[1][25] ), .A(n5422), .Z(n17027) );
  XNOR U16936 ( .A(n17033), .B(n17240), .Z(n17026) );
  XNOR U16937 ( .A(n17034), .B(n17035), .Z(n17240) );
  AND U16938 ( .A(n17241), .B(n17242), .Z(n17035) );
  NAND U16939 ( .A(n17243), .B(n17244), .Z(n17242) );
  NANDN U16940 ( .A(n17245), .B(n17246), .Z(n17241) );
  OR U16941 ( .A(n17243), .B(n17244), .Z(n17246) );
  ANDN U16942 ( .B(\stack[1][26] ), .A(n5398), .Z(n17034) );
  XNOR U16943 ( .A(n17040), .B(n17247), .Z(n17033) );
  XNOR U16944 ( .A(n17041), .B(n17042), .Z(n17247) );
  AND U16945 ( .A(n17248), .B(n17249), .Z(n17042) );
  NANDN U16946 ( .A(n17250), .B(n17251), .Z(n17249) );
  NANDN U16947 ( .A(n17252), .B(n17253), .Z(n17248) );
  NANDN U16948 ( .A(n17251), .B(n17250), .Z(n17253) );
  ANDN U16949 ( .B(\stack[1][27] ), .A(n5374), .Z(n17041) );
  XNOR U16950 ( .A(n17047), .B(n17254), .Z(n17040) );
  XNOR U16951 ( .A(n17048), .B(n17049), .Z(n17254) );
  AND U16952 ( .A(n17255), .B(n17256), .Z(n17049) );
  NAND U16953 ( .A(n17257), .B(n17258), .Z(n17256) );
  NANDN U16954 ( .A(n17259), .B(n17260), .Z(n17255) );
  OR U16955 ( .A(n17257), .B(n17258), .Z(n17260) );
  ANDN U16956 ( .B(\stack[1][28] ), .A(n5350), .Z(n17048) );
  XNOR U16957 ( .A(n17054), .B(n17261), .Z(n17047) );
  XNOR U16958 ( .A(n17055), .B(n17056), .Z(n17261) );
  AND U16959 ( .A(n17262), .B(n17263), .Z(n17056) );
  NANDN U16960 ( .A(n17264), .B(n17265), .Z(n17263) );
  NANDN U16961 ( .A(n17266), .B(n17267), .Z(n17262) );
  NANDN U16962 ( .A(n17265), .B(n17264), .Z(n17267) );
  ANDN U16963 ( .B(\stack[1][29] ), .A(n5326), .Z(n17055) );
  XNOR U16964 ( .A(n17061), .B(n17268), .Z(n17054) );
  XNOR U16965 ( .A(n17062), .B(n17063), .Z(n17268) );
  AND U16966 ( .A(n17269), .B(n17270), .Z(n17063) );
  NAND U16967 ( .A(n17271), .B(n17272), .Z(n17270) );
  NANDN U16968 ( .A(n17273), .B(n17274), .Z(n17269) );
  OR U16969 ( .A(n17271), .B(n17272), .Z(n17274) );
  ANDN U16970 ( .B(\stack[1][30] ), .A(n5302), .Z(n17062) );
  XNOR U16971 ( .A(n17068), .B(n17275), .Z(n17061) );
  XNOR U16972 ( .A(n17069), .B(n17070), .Z(n17275) );
  AND U16973 ( .A(n17276), .B(n17277), .Z(n17070) );
  NANDN U16974 ( .A(n17278), .B(n17279), .Z(n17277) );
  NANDN U16975 ( .A(n17280), .B(n17281), .Z(n17276) );
  NANDN U16976 ( .A(n17279), .B(n17278), .Z(n17281) );
  ANDN U16977 ( .B(\stack[1][31] ), .A(n5278), .Z(n17069) );
  XNOR U16978 ( .A(n17075), .B(n17282), .Z(n17068) );
  XNOR U16979 ( .A(n17076), .B(n17077), .Z(n17282) );
  AND U16980 ( .A(n17283), .B(n17284), .Z(n17077) );
  NAND U16981 ( .A(n17285), .B(n17286), .Z(n17284) );
  NANDN U16982 ( .A(n17287), .B(n17288), .Z(n17283) );
  OR U16983 ( .A(n17285), .B(n17286), .Z(n17288) );
  ANDN U16984 ( .B(\stack[1][32] ), .A(n5254), .Z(n17076) );
  XNOR U16985 ( .A(n17082), .B(n17289), .Z(n17075) );
  XNOR U16986 ( .A(n17083), .B(n17084), .Z(n17289) );
  AND U16987 ( .A(n17290), .B(n17291), .Z(n17084) );
  NAND U16988 ( .A(n17292), .B(n17293), .Z(n17291) );
  NAND U16989 ( .A(n17294), .B(n17295), .Z(n17290) );
  OR U16990 ( .A(n17292), .B(n17293), .Z(n17294) );
  ANDN U16991 ( .B(\stack[1][33] ), .A(n5230), .Z(n17083) );
  XNOR U16992 ( .A(n17089), .B(n17296), .Z(n17082) );
  XNOR U16993 ( .A(n17090), .B(n17092), .Z(n17296) );
  ANDN U16994 ( .B(n17297), .A(n17298), .Z(n17092) );
  ANDN U16995 ( .B(\stack[0][0] ), .A(n6012), .Z(n17297) );
  ANDN U16996 ( .B(\stack[1][34] ), .A(n5206), .Z(n17090) );
  XOR U16997 ( .A(n17095), .B(n17299), .Z(n17089) );
  NANDN U16998 ( .A(n5160), .B(\stack[1][36] ), .Z(n17299) );
  NANDN U16999 ( .A(n6012), .B(\stack[0][1] ), .Z(n17095) );
  ANDN U17000 ( .B(\stack[0][31] ), .A(n5292), .Z(n9146) );
  AND U17001 ( .A(n17300), .B(n17301), .Z(n9147) );
  NANDN U17002 ( .A(n9154), .B(n17302), .Z(n17300) );
  NANDN U17003 ( .A(n9153), .B(n9151), .Z(n17302) );
  XNOR U17004 ( .A(n17103), .B(n17303), .Z(n9151) );
  XNOR U17005 ( .A(n17104), .B(n17105), .Z(n17303) );
  AND U17006 ( .A(n17304), .B(n17305), .Z(n17105) );
  NANDN U17007 ( .A(n17306), .B(n17307), .Z(n17305) );
  NANDN U17008 ( .A(n17308), .B(n17309), .Z(n17304) );
  NANDN U17009 ( .A(n17307), .B(n17306), .Z(n17309) );
  ANDN U17010 ( .B(\stack[0][29] ), .A(n5316), .Z(n17104) );
  XNOR U17011 ( .A(n17110), .B(n17310), .Z(n17103) );
  XNOR U17012 ( .A(n17111), .B(n17112), .Z(n17310) );
  AND U17013 ( .A(n17311), .B(n17312), .Z(n17112) );
  NAND U17014 ( .A(n17313), .B(n17314), .Z(n17312) );
  NANDN U17015 ( .A(n17315), .B(n17316), .Z(n17311) );
  OR U17016 ( .A(n17313), .B(n17314), .Z(n17316) );
  ANDN U17017 ( .B(\stack[0][28] ), .A(n5340), .Z(n17111) );
  XNOR U17018 ( .A(n17117), .B(n17317), .Z(n17110) );
  XNOR U17019 ( .A(n17118), .B(n17119), .Z(n17317) );
  AND U17020 ( .A(n17318), .B(n17319), .Z(n17119) );
  NANDN U17021 ( .A(n17320), .B(n17321), .Z(n17319) );
  NANDN U17022 ( .A(n17322), .B(n17323), .Z(n17318) );
  NANDN U17023 ( .A(n17321), .B(n17320), .Z(n17323) );
  ANDN U17024 ( .B(\stack[0][27] ), .A(n5364), .Z(n17118) );
  XNOR U17025 ( .A(n17124), .B(n17324), .Z(n17117) );
  XNOR U17026 ( .A(n17125), .B(n17126), .Z(n17324) );
  AND U17027 ( .A(n17325), .B(n17326), .Z(n17126) );
  NAND U17028 ( .A(n17327), .B(n17328), .Z(n17326) );
  NANDN U17029 ( .A(n17329), .B(n17330), .Z(n17325) );
  OR U17030 ( .A(n17327), .B(n17328), .Z(n17330) );
  ANDN U17031 ( .B(\stack[0][26] ), .A(n5387), .Z(n17125) );
  XNOR U17032 ( .A(n17131), .B(n17331), .Z(n17124) );
  XNOR U17033 ( .A(n17132), .B(n17133), .Z(n17331) );
  AND U17034 ( .A(n17332), .B(n17333), .Z(n17133) );
  NANDN U17035 ( .A(n17334), .B(n17335), .Z(n17333) );
  NANDN U17036 ( .A(n17336), .B(n17337), .Z(n17332) );
  NANDN U17037 ( .A(n17335), .B(n17334), .Z(n17337) );
  ANDN U17038 ( .B(\stack[1][10] ), .A(n5758), .Z(n17132) );
  XNOR U17039 ( .A(n17138), .B(n17338), .Z(n17131) );
  XNOR U17040 ( .A(n17139), .B(n17140), .Z(n17338) );
  AND U17041 ( .A(n17339), .B(n17340), .Z(n17140) );
  NAND U17042 ( .A(n17341), .B(n17342), .Z(n17340) );
  NANDN U17043 ( .A(n17343), .B(n17344), .Z(n17339) );
  OR U17044 ( .A(n17341), .B(n17342), .Z(n17344) );
  ANDN U17045 ( .B(\stack[1][11] ), .A(n5734), .Z(n17139) );
  XNOR U17046 ( .A(n17145), .B(n17345), .Z(n17138) );
  XNOR U17047 ( .A(n17146), .B(n17147), .Z(n17345) );
  AND U17048 ( .A(n17346), .B(n17347), .Z(n17147) );
  NANDN U17049 ( .A(n17348), .B(n17349), .Z(n17347) );
  NANDN U17050 ( .A(n17350), .B(n17351), .Z(n17346) );
  NANDN U17051 ( .A(n17349), .B(n17348), .Z(n17351) );
  ANDN U17052 ( .B(\stack[1][12] ), .A(n5710), .Z(n17146) );
  XNOR U17053 ( .A(n17152), .B(n17352), .Z(n17145) );
  XNOR U17054 ( .A(n17153), .B(n17154), .Z(n17352) );
  AND U17055 ( .A(n17353), .B(n17354), .Z(n17154) );
  NAND U17056 ( .A(n17355), .B(n17356), .Z(n17354) );
  NANDN U17057 ( .A(n17357), .B(n17358), .Z(n17353) );
  OR U17058 ( .A(n17355), .B(n17356), .Z(n17358) );
  ANDN U17059 ( .B(\stack[1][13] ), .A(n5686), .Z(n17153) );
  XNOR U17060 ( .A(n17159), .B(n17359), .Z(n17152) );
  XNOR U17061 ( .A(n17160), .B(n17161), .Z(n17359) );
  AND U17062 ( .A(n17360), .B(n17361), .Z(n17161) );
  NANDN U17063 ( .A(n17362), .B(n17363), .Z(n17361) );
  NANDN U17064 ( .A(n17364), .B(n17365), .Z(n17360) );
  NANDN U17065 ( .A(n17363), .B(n17362), .Z(n17365) );
  ANDN U17066 ( .B(\stack[1][14] ), .A(n5662), .Z(n17160) );
  XNOR U17067 ( .A(n17166), .B(n17366), .Z(n17159) );
  XNOR U17068 ( .A(n17167), .B(n17168), .Z(n17366) );
  AND U17069 ( .A(n17367), .B(n17368), .Z(n17168) );
  NAND U17070 ( .A(n17369), .B(n17370), .Z(n17368) );
  NANDN U17071 ( .A(n17371), .B(n17372), .Z(n17367) );
  OR U17072 ( .A(n17369), .B(n17370), .Z(n17372) );
  ANDN U17073 ( .B(\stack[1][15] ), .A(n5638), .Z(n17167) );
  XNOR U17074 ( .A(n17173), .B(n17373), .Z(n17166) );
  XNOR U17075 ( .A(n17174), .B(n17175), .Z(n17373) );
  AND U17076 ( .A(n17374), .B(n17375), .Z(n17175) );
  NANDN U17077 ( .A(n17376), .B(n17377), .Z(n17375) );
  NANDN U17078 ( .A(n17378), .B(n17379), .Z(n17374) );
  NANDN U17079 ( .A(n17377), .B(n17376), .Z(n17379) );
  ANDN U17080 ( .B(\stack[1][16] ), .A(n5614), .Z(n17174) );
  XNOR U17081 ( .A(n17180), .B(n17380), .Z(n17173) );
  XNOR U17082 ( .A(n17181), .B(n17182), .Z(n17380) );
  AND U17083 ( .A(n17381), .B(n17382), .Z(n17182) );
  NAND U17084 ( .A(n17383), .B(n17384), .Z(n17382) );
  NANDN U17085 ( .A(n17385), .B(n17386), .Z(n17381) );
  OR U17086 ( .A(n17383), .B(n17384), .Z(n17386) );
  ANDN U17087 ( .B(\stack[1][17] ), .A(n5590), .Z(n17181) );
  XNOR U17088 ( .A(n17187), .B(n17387), .Z(n17180) );
  XNOR U17089 ( .A(n17188), .B(n17189), .Z(n17387) );
  AND U17090 ( .A(n17388), .B(n17389), .Z(n17189) );
  NANDN U17091 ( .A(n17390), .B(n17391), .Z(n17389) );
  NANDN U17092 ( .A(n17392), .B(n17393), .Z(n17388) );
  NANDN U17093 ( .A(n17391), .B(n17390), .Z(n17393) );
  ANDN U17094 ( .B(\stack[1][18] ), .A(n5566), .Z(n17188) );
  XNOR U17095 ( .A(n17194), .B(n17394), .Z(n17187) );
  XNOR U17096 ( .A(n17195), .B(n17196), .Z(n17394) );
  AND U17097 ( .A(n17395), .B(n17396), .Z(n17196) );
  NAND U17098 ( .A(n17397), .B(n17398), .Z(n17396) );
  NANDN U17099 ( .A(n17399), .B(n17400), .Z(n17395) );
  OR U17100 ( .A(n17397), .B(n17398), .Z(n17400) );
  ANDN U17101 ( .B(\stack[1][19] ), .A(n5542), .Z(n17195) );
  XNOR U17102 ( .A(n17201), .B(n17401), .Z(n17194) );
  XNOR U17103 ( .A(n17202), .B(n17203), .Z(n17401) );
  AND U17104 ( .A(n17402), .B(n17403), .Z(n17203) );
  NANDN U17105 ( .A(n17404), .B(n17405), .Z(n17403) );
  NANDN U17106 ( .A(n17406), .B(n17407), .Z(n17402) );
  NANDN U17107 ( .A(n17405), .B(n17404), .Z(n17407) );
  ANDN U17108 ( .B(\stack[1][20] ), .A(n5518), .Z(n17202) );
  XNOR U17109 ( .A(n17208), .B(n17408), .Z(n17201) );
  XNOR U17110 ( .A(n17209), .B(n17210), .Z(n17408) );
  AND U17111 ( .A(n17409), .B(n17410), .Z(n17210) );
  NAND U17112 ( .A(n17411), .B(n17412), .Z(n17410) );
  NANDN U17113 ( .A(n17413), .B(n17414), .Z(n17409) );
  OR U17114 ( .A(n17411), .B(n17412), .Z(n17414) );
  ANDN U17115 ( .B(\stack[1][21] ), .A(n5494), .Z(n17209) );
  XNOR U17116 ( .A(n17215), .B(n17415), .Z(n17208) );
  XNOR U17117 ( .A(n17216), .B(n17217), .Z(n17415) );
  AND U17118 ( .A(n17416), .B(n17417), .Z(n17217) );
  NANDN U17119 ( .A(n17418), .B(n17419), .Z(n17417) );
  NANDN U17120 ( .A(n17420), .B(n17421), .Z(n17416) );
  NANDN U17121 ( .A(n17419), .B(n17418), .Z(n17421) );
  ANDN U17122 ( .B(\stack[1][22] ), .A(n5470), .Z(n17216) );
  XNOR U17123 ( .A(n17222), .B(n17422), .Z(n17215) );
  XNOR U17124 ( .A(n17223), .B(n17224), .Z(n17422) );
  AND U17125 ( .A(n17423), .B(n17424), .Z(n17224) );
  NAND U17126 ( .A(n17425), .B(n17426), .Z(n17424) );
  NANDN U17127 ( .A(n17427), .B(n17428), .Z(n17423) );
  OR U17128 ( .A(n17425), .B(n17426), .Z(n17428) );
  ANDN U17129 ( .B(\stack[1][23] ), .A(n5446), .Z(n17223) );
  XNOR U17130 ( .A(n17229), .B(n17429), .Z(n17222) );
  XNOR U17131 ( .A(n17230), .B(n17231), .Z(n17429) );
  AND U17132 ( .A(n17430), .B(n17431), .Z(n17231) );
  NANDN U17133 ( .A(n17432), .B(n17433), .Z(n17431) );
  NANDN U17134 ( .A(n17434), .B(n17435), .Z(n17430) );
  NANDN U17135 ( .A(n17433), .B(n17432), .Z(n17435) );
  ANDN U17136 ( .B(\stack[1][24] ), .A(n5422), .Z(n17230) );
  XNOR U17137 ( .A(n17236), .B(n17436), .Z(n17229) );
  XNOR U17138 ( .A(n17237), .B(n17238), .Z(n17436) );
  AND U17139 ( .A(n17437), .B(n17438), .Z(n17238) );
  NAND U17140 ( .A(n17439), .B(n17440), .Z(n17438) );
  NANDN U17141 ( .A(n17441), .B(n17442), .Z(n17437) );
  OR U17142 ( .A(n17439), .B(n17440), .Z(n17442) );
  ANDN U17143 ( .B(\stack[1][25] ), .A(n5398), .Z(n17237) );
  XNOR U17144 ( .A(n17243), .B(n17443), .Z(n17236) );
  XNOR U17145 ( .A(n17244), .B(n17245), .Z(n17443) );
  AND U17146 ( .A(n17444), .B(n17445), .Z(n17245) );
  NANDN U17147 ( .A(n17446), .B(n17447), .Z(n17445) );
  NANDN U17148 ( .A(n17448), .B(n17449), .Z(n17444) );
  NANDN U17149 ( .A(n17447), .B(n17446), .Z(n17449) );
  ANDN U17150 ( .B(\stack[1][26] ), .A(n5374), .Z(n17244) );
  XNOR U17151 ( .A(n17250), .B(n17450), .Z(n17243) );
  XNOR U17152 ( .A(n17251), .B(n17252), .Z(n17450) );
  AND U17153 ( .A(n17451), .B(n17452), .Z(n17252) );
  NAND U17154 ( .A(n17453), .B(n17454), .Z(n17452) );
  NANDN U17155 ( .A(n17455), .B(n17456), .Z(n17451) );
  OR U17156 ( .A(n17453), .B(n17454), .Z(n17456) );
  ANDN U17157 ( .B(\stack[1][27] ), .A(n5350), .Z(n17251) );
  XNOR U17158 ( .A(n17257), .B(n17457), .Z(n17250) );
  XNOR U17159 ( .A(n17258), .B(n17259), .Z(n17457) );
  AND U17160 ( .A(n17458), .B(n17459), .Z(n17259) );
  NANDN U17161 ( .A(n17460), .B(n17461), .Z(n17459) );
  NANDN U17162 ( .A(n17462), .B(n17463), .Z(n17458) );
  NANDN U17163 ( .A(n17461), .B(n17460), .Z(n17463) );
  ANDN U17164 ( .B(\stack[1][28] ), .A(n5326), .Z(n17258) );
  XNOR U17165 ( .A(n17264), .B(n17464), .Z(n17257) );
  XNOR U17166 ( .A(n17265), .B(n17266), .Z(n17464) );
  AND U17167 ( .A(n17465), .B(n17466), .Z(n17266) );
  NAND U17168 ( .A(n17467), .B(n17468), .Z(n17466) );
  NANDN U17169 ( .A(n17469), .B(n17470), .Z(n17465) );
  OR U17170 ( .A(n17467), .B(n17468), .Z(n17470) );
  ANDN U17171 ( .B(\stack[1][29] ), .A(n5302), .Z(n17265) );
  XNOR U17172 ( .A(n17271), .B(n17471), .Z(n17264) );
  XNOR U17173 ( .A(n17272), .B(n17273), .Z(n17471) );
  AND U17174 ( .A(n17472), .B(n17473), .Z(n17273) );
  NANDN U17175 ( .A(n17474), .B(n17475), .Z(n17473) );
  NANDN U17176 ( .A(n17476), .B(n17477), .Z(n17472) );
  NANDN U17177 ( .A(n17475), .B(n17474), .Z(n17477) );
  ANDN U17178 ( .B(\stack[1][30] ), .A(n5278), .Z(n17272) );
  XNOR U17179 ( .A(n17278), .B(n17478), .Z(n17271) );
  XNOR U17180 ( .A(n17279), .B(n17280), .Z(n17478) );
  AND U17181 ( .A(n17479), .B(n17480), .Z(n17280) );
  NAND U17182 ( .A(n17481), .B(n17482), .Z(n17480) );
  NANDN U17183 ( .A(n17483), .B(n17484), .Z(n17479) );
  OR U17184 ( .A(n17481), .B(n17482), .Z(n17484) );
  ANDN U17185 ( .B(\stack[1][31] ), .A(n5254), .Z(n17279) );
  XNOR U17186 ( .A(n17285), .B(n17485), .Z(n17278) );
  XNOR U17187 ( .A(n17286), .B(n17287), .Z(n17485) );
  AND U17188 ( .A(n17486), .B(n17487), .Z(n17287) );
  NAND U17189 ( .A(n17488), .B(n17489), .Z(n17487) );
  NAND U17190 ( .A(n17490), .B(n17491), .Z(n17486) );
  OR U17191 ( .A(n17488), .B(n17489), .Z(n17490) );
  ANDN U17192 ( .B(\stack[1][32] ), .A(n5230), .Z(n17286) );
  XNOR U17193 ( .A(n17292), .B(n17492), .Z(n17285) );
  XNOR U17194 ( .A(n17293), .B(n17295), .Z(n17492) );
  ANDN U17195 ( .B(n17493), .A(n17494), .Z(n17295) );
  ANDN U17196 ( .B(\stack[0][0] ), .A(n5988), .Z(n17493) );
  ANDN U17197 ( .B(\stack[1][33] ), .A(n5206), .Z(n17293) );
  XOR U17198 ( .A(n17298), .B(n17495), .Z(n17292) );
  NANDN U17199 ( .A(n5160), .B(\stack[1][35] ), .Z(n17495) );
  NANDN U17200 ( .A(n5988), .B(\stack[0][1] ), .Z(n17298) );
  ANDN U17201 ( .B(\stack[1][5] ), .A(n5878), .Z(n9153) );
  AND U17202 ( .A(n17496), .B(n17497), .Z(n9154) );
  NANDN U17203 ( .A(n9158), .B(n9160), .Z(n17497) );
  NANDN U17204 ( .A(n9161), .B(n17498), .Z(n17496) );
  NANDN U17205 ( .A(n9160), .B(n9158), .Z(n17498) );
  XOR U17206 ( .A(n17306), .B(n17499), .Z(n9158) );
  XNOR U17207 ( .A(n17307), .B(n17308), .Z(n17499) );
  AND U17208 ( .A(n17500), .B(n17501), .Z(n17308) );
  NAND U17209 ( .A(n17502), .B(n17503), .Z(n17501) );
  NANDN U17210 ( .A(n17504), .B(n17505), .Z(n17500) );
  OR U17211 ( .A(n17502), .B(n17503), .Z(n17505) );
  ANDN U17212 ( .B(\stack[0][28] ), .A(n5316), .Z(n17307) );
  XNOR U17213 ( .A(n17313), .B(n17506), .Z(n17306) );
  XNOR U17214 ( .A(n17314), .B(n17315), .Z(n17506) );
  AND U17215 ( .A(n17507), .B(n17508), .Z(n17315) );
  NANDN U17216 ( .A(n17509), .B(n17510), .Z(n17508) );
  NANDN U17217 ( .A(n17511), .B(n17512), .Z(n17507) );
  NANDN U17218 ( .A(n17510), .B(n17509), .Z(n17512) );
  ANDN U17219 ( .B(\stack[0][27] ), .A(n5340), .Z(n17314) );
  XNOR U17220 ( .A(n17320), .B(n17513), .Z(n17313) );
  XNOR U17221 ( .A(n17321), .B(n17322), .Z(n17513) );
  AND U17222 ( .A(n17514), .B(n17515), .Z(n17322) );
  NAND U17223 ( .A(n17516), .B(n17517), .Z(n17515) );
  NANDN U17224 ( .A(n17518), .B(n17519), .Z(n17514) );
  OR U17225 ( .A(n17516), .B(n17517), .Z(n17519) );
  ANDN U17226 ( .B(\stack[0][26] ), .A(n5364), .Z(n17321) );
  XNOR U17227 ( .A(n17327), .B(n17520), .Z(n17320) );
  XNOR U17228 ( .A(n17328), .B(n17329), .Z(n17520) );
  AND U17229 ( .A(n17521), .B(n17522), .Z(n17329) );
  NANDN U17230 ( .A(n17523), .B(n17524), .Z(n17522) );
  NANDN U17231 ( .A(n17525), .B(n17526), .Z(n17521) );
  NANDN U17232 ( .A(n17524), .B(n17523), .Z(n17526) );
  ANDN U17233 ( .B(\stack[0][25] ), .A(n5387), .Z(n17328) );
  XNOR U17234 ( .A(n17334), .B(n17527), .Z(n17327) );
  XNOR U17235 ( .A(n17335), .B(n17336), .Z(n17527) );
  AND U17236 ( .A(n17528), .B(n17529), .Z(n17336) );
  NAND U17237 ( .A(n17530), .B(n17531), .Z(n17529) );
  NANDN U17238 ( .A(n17532), .B(n17533), .Z(n17528) );
  OR U17239 ( .A(n17530), .B(n17531), .Z(n17533) );
  ANDN U17240 ( .B(\stack[1][10] ), .A(n5734), .Z(n17335) );
  XNOR U17241 ( .A(n17341), .B(n17534), .Z(n17334) );
  XNOR U17242 ( .A(n17342), .B(n17343), .Z(n17534) );
  AND U17243 ( .A(n17535), .B(n17536), .Z(n17343) );
  NANDN U17244 ( .A(n17537), .B(n17538), .Z(n17536) );
  NANDN U17245 ( .A(n17539), .B(n17540), .Z(n17535) );
  NANDN U17246 ( .A(n17538), .B(n17537), .Z(n17540) );
  ANDN U17247 ( .B(\stack[1][11] ), .A(n5710), .Z(n17342) );
  XNOR U17248 ( .A(n17348), .B(n17541), .Z(n17341) );
  XNOR U17249 ( .A(n17349), .B(n17350), .Z(n17541) );
  AND U17250 ( .A(n17542), .B(n17543), .Z(n17350) );
  NAND U17251 ( .A(n17544), .B(n17545), .Z(n17543) );
  NANDN U17252 ( .A(n17546), .B(n17547), .Z(n17542) );
  OR U17253 ( .A(n17544), .B(n17545), .Z(n17547) );
  ANDN U17254 ( .B(\stack[1][12] ), .A(n5686), .Z(n17349) );
  XNOR U17255 ( .A(n17355), .B(n17548), .Z(n17348) );
  XNOR U17256 ( .A(n17356), .B(n17357), .Z(n17548) );
  AND U17257 ( .A(n17549), .B(n17550), .Z(n17357) );
  NANDN U17258 ( .A(n17551), .B(n17552), .Z(n17550) );
  NANDN U17259 ( .A(n17553), .B(n17554), .Z(n17549) );
  NANDN U17260 ( .A(n17552), .B(n17551), .Z(n17554) );
  ANDN U17261 ( .B(\stack[1][13] ), .A(n5662), .Z(n17356) );
  XNOR U17262 ( .A(n17362), .B(n17555), .Z(n17355) );
  XNOR U17263 ( .A(n17363), .B(n17364), .Z(n17555) );
  AND U17264 ( .A(n17556), .B(n17557), .Z(n17364) );
  NAND U17265 ( .A(n17558), .B(n17559), .Z(n17557) );
  NANDN U17266 ( .A(n17560), .B(n17561), .Z(n17556) );
  OR U17267 ( .A(n17558), .B(n17559), .Z(n17561) );
  ANDN U17268 ( .B(\stack[1][14] ), .A(n5638), .Z(n17363) );
  XNOR U17269 ( .A(n17369), .B(n17562), .Z(n17362) );
  XNOR U17270 ( .A(n17370), .B(n17371), .Z(n17562) );
  AND U17271 ( .A(n17563), .B(n17564), .Z(n17371) );
  NANDN U17272 ( .A(n17565), .B(n17566), .Z(n17564) );
  NANDN U17273 ( .A(n17567), .B(n17568), .Z(n17563) );
  NANDN U17274 ( .A(n17566), .B(n17565), .Z(n17568) );
  ANDN U17275 ( .B(\stack[1][15] ), .A(n5614), .Z(n17370) );
  XNOR U17276 ( .A(n17376), .B(n17569), .Z(n17369) );
  XNOR U17277 ( .A(n17377), .B(n17378), .Z(n17569) );
  AND U17278 ( .A(n17570), .B(n17571), .Z(n17378) );
  NAND U17279 ( .A(n17572), .B(n17573), .Z(n17571) );
  NANDN U17280 ( .A(n17574), .B(n17575), .Z(n17570) );
  OR U17281 ( .A(n17572), .B(n17573), .Z(n17575) );
  ANDN U17282 ( .B(\stack[1][16] ), .A(n5590), .Z(n17377) );
  XNOR U17283 ( .A(n17383), .B(n17576), .Z(n17376) );
  XNOR U17284 ( .A(n17384), .B(n17385), .Z(n17576) );
  AND U17285 ( .A(n17577), .B(n17578), .Z(n17385) );
  NANDN U17286 ( .A(n17579), .B(n17580), .Z(n17578) );
  NANDN U17287 ( .A(n17581), .B(n17582), .Z(n17577) );
  NANDN U17288 ( .A(n17580), .B(n17579), .Z(n17582) );
  ANDN U17289 ( .B(\stack[1][17] ), .A(n5566), .Z(n17384) );
  XNOR U17290 ( .A(n17390), .B(n17583), .Z(n17383) );
  XNOR U17291 ( .A(n17391), .B(n17392), .Z(n17583) );
  AND U17292 ( .A(n17584), .B(n17585), .Z(n17392) );
  NAND U17293 ( .A(n17586), .B(n17587), .Z(n17585) );
  NANDN U17294 ( .A(n17588), .B(n17589), .Z(n17584) );
  OR U17295 ( .A(n17586), .B(n17587), .Z(n17589) );
  ANDN U17296 ( .B(\stack[1][18] ), .A(n5542), .Z(n17391) );
  XNOR U17297 ( .A(n17397), .B(n17590), .Z(n17390) );
  XNOR U17298 ( .A(n17398), .B(n17399), .Z(n17590) );
  AND U17299 ( .A(n17591), .B(n17592), .Z(n17399) );
  NANDN U17300 ( .A(n17593), .B(n17594), .Z(n17592) );
  NANDN U17301 ( .A(n17595), .B(n17596), .Z(n17591) );
  NANDN U17302 ( .A(n17594), .B(n17593), .Z(n17596) );
  ANDN U17303 ( .B(\stack[1][19] ), .A(n5518), .Z(n17398) );
  XNOR U17304 ( .A(n17404), .B(n17597), .Z(n17397) );
  XNOR U17305 ( .A(n17405), .B(n17406), .Z(n17597) );
  AND U17306 ( .A(n17598), .B(n17599), .Z(n17406) );
  NAND U17307 ( .A(n17600), .B(n17601), .Z(n17599) );
  NANDN U17308 ( .A(n17602), .B(n17603), .Z(n17598) );
  OR U17309 ( .A(n17600), .B(n17601), .Z(n17603) );
  ANDN U17310 ( .B(\stack[1][20] ), .A(n5494), .Z(n17405) );
  XNOR U17311 ( .A(n17411), .B(n17604), .Z(n17404) );
  XNOR U17312 ( .A(n17412), .B(n17413), .Z(n17604) );
  AND U17313 ( .A(n17605), .B(n17606), .Z(n17413) );
  NANDN U17314 ( .A(n17607), .B(n17608), .Z(n17606) );
  NANDN U17315 ( .A(n17609), .B(n17610), .Z(n17605) );
  NANDN U17316 ( .A(n17608), .B(n17607), .Z(n17610) );
  ANDN U17317 ( .B(\stack[1][21] ), .A(n5470), .Z(n17412) );
  XNOR U17318 ( .A(n17418), .B(n17611), .Z(n17411) );
  XNOR U17319 ( .A(n17419), .B(n17420), .Z(n17611) );
  AND U17320 ( .A(n17612), .B(n17613), .Z(n17420) );
  NAND U17321 ( .A(n17614), .B(n17615), .Z(n17613) );
  NANDN U17322 ( .A(n17616), .B(n17617), .Z(n17612) );
  OR U17323 ( .A(n17614), .B(n17615), .Z(n17617) );
  ANDN U17324 ( .B(\stack[1][22] ), .A(n5446), .Z(n17419) );
  XNOR U17325 ( .A(n17425), .B(n17618), .Z(n17418) );
  XNOR U17326 ( .A(n17426), .B(n17427), .Z(n17618) );
  AND U17327 ( .A(n17619), .B(n17620), .Z(n17427) );
  NANDN U17328 ( .A(n17621), .B(n17622), .Z(n17620) );
  NANDN U17329 ( .A(n17623), .B(n17624), .Z(n17619) );
  NANDN U17330 ( .A(n17622), .B(n17621), .Z(n17624) );
  ANDN U17331 ( .B(\stack[1][23] ), .A(n5422), .Z(n17426) );
  XNOR U17332 ( .A(n17432), .B(n17625), .Z(n17425) );
  XNOR U17333 ( .A(n17433), .B(n17434), .Z(n17625) );
  AND U17334 ( .A(n17626), .B(n17627), .Z(n17434) );
  NAND U17335 ( .A(n17628), .B(n17629), .Z(n17627) );
  NANDN U17336 ( .A(n17630), .B(n17631), .Z(n17626) );
  OR U17337 ( .A(n17628), .B(n17629), .Z(n17631) );
  ANDN U17338 ( .B(\stack[1][24] ), .A(n5398), .Z(n17433) );
  XNOR U17339 ( .A(n17439), .B(n17632), .Z(n17432) );
  XNOR U17340 ( .A(n17440), .B(n17441), .Z(n17632) );
  AND U17341 ( .A(n17633), .B(n17634), .Z(n17441) );
  NANDN U17342 ( .A(n17635), .B(n17636), .Z(n17634) );
  NANDN U17343 ( .A(n17637), .B(n17638), .Z(n17633) );
  NANDN U17344 ( .A(n17636), .B(n17635), .Z(n17638) );
  ANDN U17345 ( .B(\stack[1][25] ), .A(n5374), .Z(n17440) );
  XNOR U17346 ( .A(n17446), .B(n17639), .Z(n17439) );
  XNOR U17347 ( .A(n17447), .B(n17448), .Z(n17639) );
  AND U17348 ( .A(n17640), .B(n17641), .Z(n17448) );
  NAND U17349 ( .A(n17642), .B(n17643), .Z(n17641) );
  NANDN U17350 ( .A(n17644), .B(n17645), .Z(n17640) );
  OR U17351 ( .A(n17642), .B(n17643), .Z(n17645) );
  ANDN U17352 ( .B(\stack[1][26] ), .A(n5350), .Z(n17447) );
  XNOR U17353 ( .A(n17453), .B(n17646), .Z(n17446) );
  XNOR U17354 ( .A(n17454), .B(n17455), .Z(n17646) );
  AND U17355 ( .A(n17647), .B(n17648), .Z(n17455) );
  NANDN U17356 ( .A(n17649), .B(n17650), .Z(n17648) );
  NANDN U17357 ( .A(n17651), .B(n17652), .Z(n17647) );
  NANDN U17358 ( .A(n17650), .B(n17649), .Z(n17652) );
  ANDN U17359 ( .B(\stack[1][27] ), .A(n5326), .Z(n17454) );
  XNOR U17360 ( .A(n17460), .B(n17653), .Z(n17453) );
  XNOR U17361 ( .A(n17461), .B(n17462), .Z(n17653) );
  AND U17362 ( .A(n17654), .B(n17655), .Z(n17462) );
  NAND U17363 ( .A(n17656), .B(n17657), .Z(n17655) );
  NANDN U17364 ( .A(n17658), .B(n17659), .Z(n17654) );
  OR U17365 ( .A(n17656), .B(n17657), .Z(n17659) );
  ANDN U17366 ( .B(\stack[1][28] ), .A(n5302), .Z(n17461) );
  XNOR U17367 ( .A(n17467), .B(n17660), .Z(n17460) );
  XNOR U17368 ( .A(n17468), .B(n17469), .Z(n17660) );
  AND U17369 ( .A(n17661), .B(n17662), .Z(n17469) );
  NANDN U17370 ( .A(n17663), .B(n17664), .Z(n17662) );
  NANDN U17371 ( .A(n17665), .B(n17666), .Z(n17661) );
  NANDN U17372 ( .A(n17664), .B(n17663), .Z(n17666) );
  ANDN U17373 ( .B(\stack[1][29] ), .A(n5278), .Z(n17468) );
  XNOR U17374 ( .A(n17474), .B(n17667), .Z(n17467) );
  XNOR U17375 ( .A(n17475), .B(n17476), .Z(n17667) );
  AND U17376 ( .A(n17668), .B(n17669), .Z(n17476) );
  NAND U17377 ( .A(n17670), .B(n17671), .Z(n17669) );
  NANDN U17378 ( .A(n17672), .B(n17673), .Z(n17668) );
  OR U17379 ( .A(n17670), .B(n17671), .Z(n17673) );
  ANDN U17380 ( .B(\stack[1][30] ), .A(n5254), .Z(n17475) );
  XNOR U17381 ( .A(n17481), .B(n17674), .Z(n17474) );
  XNOR U17382 ( .A(n17482), .B(n17483), .Z(n17674) );
  AND U17383 ( .A(n17675), .B(n17676), .Z(n17483) );
  NAND U17384 ( .A(n17677), .B(n17678), .Z(n17676) );
  NAND U17385 ( .A(n17679), .B(n17680), .Z(n17675) );
  OR U17386 ( .A(n17677), .B(n17678), .Z(n17679) );
  ANDN U17387 ( .B(\stack[1][31] ), .A(n5230), .Z(n17482) );
  XNOR U17388 ( .A(n17488), .B(n17681), .Z(n17481) );
  XNOR U17389 ( .A(n17489), .B(n17491), .Z(n17681) );
  ANDN U17390 ( .B(n17682), .A(n17683), .Z(n17491) );
  ANDN U17391 ( .B(\stack[0][0] ), .A(n5964), .Z(n17682) );
  ANDN U17392 ( .B(\stack[1][32] ), .A(n5206), .Z(n17489) );
  XOR U17393 ( .A(n17494), .B(n17684), .Z(n17488) );
  NANDN U17394 ( .A(n5160), .B(\stack[1][34] ), .Z(n17684) );
  NANDN U17395 ( .A(n5964), .B(\stack[0][1] ), .Z(n17494) );
  ANDN U17396 ( .B(\stack[0][29] ), .A(n5292), .Z(n9160) );
  AND U17397 ( .A(n17685), .B(n17686), .Z(n9161) );
  NANDN U17398 ( .A(n9168), .B(n17687), .Z(n17685) );
  NANDN U17399 ( .A(n9167), .B(n9165), .Z(n17687) );
  XNOR U17400 ( .A(n17502), .B(n17688), .Z(n9165) );
  XNOR U17401 ( .A(n17503), .B(n17504), .Z(n17688) );
  AND U17402 ( .A(n17689), .B(n17690), .Z(n17504) );
  NANDN U17403 ( .A(n17691), .B(n17692), .Z(n17690) );
  NANDN U17404 ( .A(n17693), .B(n17694), .Z(n17689) );
  NANDN U17405 ( .A(n17692), .B(n17691), .Z(n17694) );
  ANDN U17406 ( .B(\stack[0][27] ), .A(n5316), .Z(n17503) );
  XNOR U17407 ( .A(n17509), .B(n17695), .Z(n17502) );
  XNOR U17408 ( .A(n17510), .B(n17511), .Z(n17695) );
  AND U17409 ( .A(n17696), .B(n17697), .Z(n17511) );
  NAND U17410 ( .A(n17698), .B(n17699), .Z(n17697) );
  NANDN U17411 ( .A(n17700), .B(n17701), .Z(n17696) );
  OR U17412 ( .A(n17698), .B(n17699), .Z(n17701) );
  ANDN U17413 ( .B(\stack[0][26] ), .A(n5340), .Z(n17510) );
  XNOR U17414 ( .A(n17516), .B(n17702), .Z(n17509) );
  XNOR U17415 ( .A(n17517), .B(n17518), .Z(n17702) );
  AND U17416 ( .A(n17703), .B(n17704), .Z(n17518) );
  NANDN U17417 ( .A(n17705), .B(n17706), .Z(n17704) );
  NANDN U17418 ( .A(n17707), .B(n17708), .Z(n17703) );
  NANDN U17419 ( .A(n17706), .B(n17705), .Z(n17708) );
  ANDN U17420 ( .B(\stack[0][25] ), .A(n5364), .Z(n17517) );
  XNOR U17421 ( .A(n17523), .B(n17709), .Z(n17516) );
  XNOR U17422 ( .A(n17524), .B(n17525), .Z(n17709) );
  AND U17423 ( .A(n17710), .B(n17711), .Z(n17525) );
  NAND U17424 ( .A(n17712), .B(n17713), .Z(n17711) );
  NANDN U17425 ( .A(n17714), .B(n17715), .Z(n17710) );
  OR U17426 ( .A(n17712), .B(n17713), .Z(n17715) );
  ANDN U17427 ( .B(\stack[0][24] ), .A(n5387), .Z(n17524) );
  XNOR U17428 ( .A(n17530), .B(n17716), .Z(n17523) );
  XNOR U17429 ( .A(n17531), .B(n17532), .Z(n17716) );
  AND U17430 ( .A(n17717), .B(n17718), .Z(n17532) );
  NANDN U17431 ( .A(n17719), .B(n17720), .Z(n17718) );
  NANDN U17432 ( .A(n17721), .B(n17722), .Z(n17717) );
  NANDN U17433 ( .A(n17720), .B(n17719), .Z(n17722) );
  ANDN U17434 ( .B(\stack[1][10] ), .A(n5710), .Z(n17531) );
  XNOR U17435 ( .A(n17537), .B(n17723), .Z(n17530) );
  XNOR U17436 ( .A(n17538), .B(n17539), .Z(n17723) );
  AND U17437 ( .A(n17724), .B(n17725), .Z(n17539) );
  NAND U17438 ( .A(n17726), .B(n17727), .Z(n17725) );
  NANDN U17439 ( .A(n17728), .B(n17729), .Z(n17724) );
  OR U17440 ( .A(n17726), .B(n17727), .Z(n17729) );
  ANDN U17441 ( .B(\stack[1][11] ), .A(n5686), .Z(n17538) );
  XNOR U17442 ( .A(n17544), .B(n17730), .Z(n17537) );
  XNOR U17443 ( .A(n17545), .B(n17546), .Z(n17730) );
  AND U17444 ( .A(n17731), .B(n17732), .Z(n17546) );
  NANDN U17445 ( .A(n17733), .B(n17734), .Z(n17732) );
  NANDN U17446 ( .A(n17735), .B(n17736), .Z(n17731) );
  NANDN U17447 ( .A(n17734), .B(n17733), .Z(n17736) );
  ANDN U17448 ( .B(\stack[1][12] ), .A(n5662), .Z(n17545) );
  XNOR U17449 ( .A(n17551), .B(n17737), .Z(n17544) );
  XNOR U17450 ( .A(n17552), .B(n17553), .Z(n17737) );
  AND U17451 ( .A(n17738), .B(n17739), .Z(n17553) );
  NAND U17452 ( .A(n17740), .B(n17741), .Z(n17739) );
  NANDN U17453 ( .A(n17742), .B(n17743), .Z(n17738) );
  OR U17454 ( .A(n17740), .B(n17741), .Z(n17743) );
  ANDN U17455 ( .B(\stack[1][13] ), .A(n5638), .Z(n17552) );
  XNOR U17456 ( .A(n17558), .B(n17744), .Z(n17551) );
  XNOR U17457 ( .A(n17559), .B(n17560), .Z(n17744) );
  AND U17458 ( .A(n17745), .B(n17746), .Z(n17560) );
  NANDN U17459 ( .A(n17747), .B(n17748), .Z(n17746) );
  NANDN U17460 ( .A(n17749), .B(n17750), .Z(n17745) );
  NANDN U17461 ( .A(n17748), .B(n17747), .Z(n17750) );
  ANDN U17462 ( .B(\stack[1][14] ), .A(n5614), .Z(n17559) );
  XNOR U17463 ( .A(n17565), .B(n17751), .Z(n17558) );
  XNOR U17464 ( .A(n17566), .B(n17567), .Z(n17751) );
  AND U17465 ( .A(n17752), .B(n17753), .Z(n17567) );
  NAND U17466 ( .A(n17754), .B(n17755), .Z(n17753) );
  NANDN U17467 ( .A(n17756), .B(n17757), .Z(n17752) );
  OR U17468 ( .A(n17754), .B(n17755), .Z(n17757) );
  ANDN U17469 ( .B(\stack[1][15] ), .A(n5590), .Z(n17566) );
  XNOR U17470 ( .A(n17572), .B(n17758), .Z(n17565) );
  XNOR U17471 ( .A(n17573), .B(n17574), .Z(n17758) );
  AND U17472 ( .A(n17759), .B(n17760), .Z(n17574) );
  NANDN U17473 ( .A(n17761), .B(n17762), .Z(n17760) );
  NANDN U17474 ( .A(n17763), .B(n17764), .Z(n17759) );
  NANDN U17475 ( .A(n17762), .B(n17761), .Z(n17764) );
  ANDN U17476 ( .B(\stack[1][16] ), .A(n5566), .Z(n17573) );
  XNOR U17477 ( .A(n17579), .B(n17765), .Z(n17572) );
  XNOR U17478 ( .A(n17580), .B(n17581), .Z(n17765) );
  AND U17479 ( .A(n17766), .B(n17767), .Z(n17581) );
  NAND U17480 ( .A(n17768), .B(n17769), .Z(n17767) );
  NANDN U17481 ( .A(n17770), .B(n17771), .Z(n17766) );
  OR U17482 ( .A(n17768), .B(n17769), .Z(n17771) );
  ANDN U17483 ( .B(\stack[1][17] ), .A(n5542), .Z(n17580) );
  XNOR U17484 ( .A(n17586), .B(n17772), .Z(n17579) );
  XNOR U17485 ( .A(n17587), .B(n17588), .Z(n17772) );
  AND U17486 ( .A(n17773), .B(n17774), .Z(n17588) );
  NANDN U17487 ( .A(n17775), .B(n17776), .Z(n17774) );
  NANDN U17488 ( .A(n17777), .B(n17778), .Z(n17773) );
  NANDN U17489 ( .A(n17776), .B(n17775), .Z(n17778) );
  ANDN U17490 ( .B(\stack[1][18] ), .A(n5518), .Z(n17587) );
  XNOR U17491 ( .A(n17593), .B(n17779), .Z(n17586) );
  XNOR U17492 ( .A(n17594), .B(n17595), .Z(n17779) );
  AND U17493 ( .A(n17780), .B(n17781), .Z(n17595) );
  NAND U17494 ( .A(n17782), .B(n17783), .Z(n17781) );
  NANDN U17495 ( .A(n17784), .B(n17785), .Z(n17780) );
  OR U17496 ( .A(n17782), .B(n17783), .Z(n17785) );
  ANDN U17497 ( .B(\stack[1][19] ), .A(n5494), .Z(n17594) );
  XNOR U17498 ( .A(n17600), .B(n17786), .Z(n17593) );
  XNOR U17499 ( .A(n17601), .B(n17602), .Z(n17786) );
  AND U17500 ( .A(n17787), .B(n17788), .Z(n17602) );
  NANDN U17501 ( .A(n17789), .B(n17790), .Z(n17788) );
  NANDN U17502 ( .A(n17791), .B(n17792), .Z(n17787) );
  NANDN U17503 ( .A(n17790), .B(n17789), .Z(n17792) );
  ANDN U17504 ( .B(\stack[1][20] ), .A(n5470), .Z(n17601) );
  XNOR U17505 ( .A(n17607), .B(n17793), .Z(n17600) );
  XNOR U17506 ( .A(n17608), .B(n17609), .Z(n17793) );
  AND U17507 ( .A(n17794), .B(n17795), .Z(n17609) );
  NAND U17508 ( .A(n17796), .B(n17797), .Z(n17795) );
  NANDN U17509 ( .A(n17798), .B(n17799), .Z(n17794) );
  OR U17510 ( .A(n17796), .B(n17797), .Z(n17799) );
  ANDN U17511 ( .B(\stack[1][21] ), .A(n5446), .Z(n17608) );
  XNOR U17512 ( .A(n17614), .B(n17800), .Z(n17607) );
  XNOR U17513 ( .A(n17615), .B(n17616), .Z(n17800) );
  AND U17514 ( .A(n17801), .B(n17802), .Z(n17616) );
  NANDN U17515 ( .A(n17803), .B(n17804), .Z(n17802) );
  NANDN U17516 ( .A(n17805), .B(n17806), .Z(n17801) );
  NANDN U17517 ( .A(n17804), .B(n17803), .Z(n17806) );
  ANDN U17518 ( .B(\stack[1][22] ), .A(n5422), .Z(n17615) );
  XNOR U17519 ( .A(n17621), .B(n17807), .Z(n17614) );
  XNOR U17520 ( .A(n17622), .B(n17623), .Z(n17807) );
  AND U17521 ( .A(n17808), .B(n17809), .Z(n17623) );
  NAND U17522 ( .A(n17810), .B(n17811), .Z(n17809) );
  NANDN U17523 ( .A(n17812), .B(n17813), .Z(n17808) );
  OR U17524 ( .A(n17810), .B(n17811), .Z(n17813) );
  ANDN U17525 ( .B(\stack[1][23] ), .A(n5398), .Z(n17622) );
  XNOR U17526 ( .A(n17628), .B(n17814), .Z(n17621) );
  XNOR U17527 ( .A(n17629), .B(n17630), .Z(n17814) );
  AND U17528 ( .A(n17815), .B(n17816), .Z(n17630) );
  NANDN U17529 ( .A(n17817), .B(n17818), .Z(n17816) );
  NANDN U17530 ( .A(n17819), .B(n17820), .Z(n17815) );
  NANDN U17531 ( .A(n17818), .B(n17817), .Z(n17820) );
  ANDN U17532 ( .B(\stack[1][24] ), .A(n5374), .Z(n17629) );
  XNOR U17533 ( .A(n17635), .B(n17821), .Z(n17628) );
  XNOR U17534 ( .A(n17636), .B(n17637), .Z(n17821) );
  AND U17535 ( .A(n17822), .B(n17823), .Z(n17637) );
  NAND U17536 ( .A(n17824), .B(n17825), .Z(n17823) );
  NANDN U17537 ( .A(n17826), .B(n17827), .Z(n17822) );
  OR U17538 ( .A(n17824), .B(n17825), .Z(n17827) );
  ANDN U17539 ( .B(\stack[1][25] ), .A(n5350), .Z(n17636) );
  XNOR U17540 ( .A(n17642), .B(n17828), .Z(n17635) );
  XNOR U17541 ( .A(n17643), .B(n17644), .Z(n17828) );
  AND U17542 ( .A(n17829), .B(n17830), .Z(n17644) );
  NANDN U17543 ( .A(n17831), .B(n17832), .Z(n17830) );
  NANDN U17544 ( .A(n17833), .B(n17834), .Z(n17829) );
  NANDN U17545 ( .A(n17832), .B(n17831), .Z(n17834) );
  ANDN U17546 ( .B(\stack[1][26] ), .A(n5326), .Z(n17643) );
  XNOR U17547 ( .A(n17649), .B(n17835), .Z(n17642) );
  XNOR U17548 ( .A(n17650), .B(n17651), .Z(n17835) );
  AND U17549 ( .A(n17836), .B(n17837), .Z(n17651) );
  NAND U17550 ( .A(n17838), .B(n17839), .Z(n17837) );
  NANDN U17551 ( .A(n17840), .B(n17841), .Z(n17836) );
  OR U17552 ( .A(n17838), .B(n17839), .Z(n17841) );
  ANDN U17553 ( .B(\stack[1][27] ), .A(n5302), .Z(n17650) );
  XNOR U17554 ( .A(n17656), .B(n17842), .Z(n17649) );
  XNOR U17555 ( .A(n17657), .B(n17658), .Z(n17842) );
  AND U17556 ( .A(n17843), .B(n17844), .Z(n17658) );
  NANDN U17557 ( .A(n17845), .B(n17846), .Z(n17844) );
  NANDN U17558 ( .A(n17847), .B(n17848), .Z(n17843) );
  NANDN U17559 ( .A(n17846), .B(n17845), .Z(n17848) );
  ANDN U17560 ( .B(\stack[1][28] ), .A(n5278), .Z(n17657) );
  XNOR U17561 ( .A(n17663), .B(n17849), .Z(n17656) );
  XNOR U17562 ( .A(n17664), .B(n17665), .Z(n17849) );
  AND U17563 ( .A(n17850), .B(n17851), .Z(n17665) );
  NAND U17564 ( .A(n17852), .B(n17853), .Z(n17851) );
  NANDN U17565 ( .A(n17854), .B(n17855), .Z(n17850) );
  OR U17566 ( .A(n17852), .B(n17853), .Z(n17855) );
  ANDN U17567 ( .B(\stack[1][29] ), .A(n5254), .Z(n17664) );
  XNOR U17568 ( .A(n17670), .B(n17856), .Z(n17663) );
  XNOR U17569 ( .A(n17671), .B(n17672), .Z(n17856) );
  AND U17570 ( .A(n17857), .B(n17858), .Z(n17672) );
  NAND U17571 ( .A(n17859), .B(n17860), .Z(n17858) );
  NAND U17572 ( .A(n17861), .B(n17862), .Z(n17857) );
  OR U17573 ( .A(n17859), .B(n17860), .Z(n17861) );
  ANDN U17574 ( .B(\stack[1][30] ), .A(n5230), .Z(n17671) );
  XNOR U17575 ( .A(n17677), .B(n17863), .Z(n17670) );
  XNOR U17576 ( .A(n17678), .B(n17680), .Z(n17863) );
  ANDN U17577 ( .B(n17864), .A(n17865), .Z(n17680) );
  ANDN U17578 ( .B(\stack[0][0] ), .A(n5940), .Z(n17864) );
  ANDN U17579 ( .B(\stack[1][31] ), .A(n5206), .Z(n17678) );
  XOR U17580 ( .A(n17683), .B(n17866), .Z(n17677) );
  NANDN U17581 ( .A(n5160), .B(\stack[1][33] ), .Z(n17866) );
  NANDN U17582 ( .A(n5940), .B(\stack[0][1] ), .Z(n17683) );
  ANDN U17583 ( .B(\stack[1][5] ), .A(n5830), .Z(n9167) );
  AND U17584 ( .A(n17867), .B(n17868), .Z(n9168) );
  NANDN U17585 ( .A(n9172), .B(n9174), .Z(n17868) );
  NANDN U17586 ( .A(n9175), .B(n17869), .Z(n17867) );
  NANDN U17587 ( .A(n9174), .B(n9172), .Z(n17869) );
  XOR U17588 ( .A(n17691), .B(n17870), .Z(n9172) );
  XNOR U17589 ( .A(n17692), .B(n17693), .Z(n17870) );
  AND U17590 ( .A(n17871), .B(n17872), .Z(n17693) );
  NAND U17591 ( .A(n17873), .B(n17874), .Z(n17872) );
  NANDN U17592 ( .A(n17875), .B(n17876), .Z(n17871) );
  OR U17593 ( .A(n17873), .B(n17874), .Z(n17876) );
  ANDN U17594 ( .B(\stack[0][26] ), .A(n5316), .Z(n17692) );
  XNOR U17595 ( .A(n17698), .B(n17877), .Z(n17691) );
  XNOR U17596 ( .A(n17699), .B(n17700), .Z(n17877) );
  AND U17597 ( .A(n17878), .B(n17879), .Z(n17700) );
  NANDN U17598 ( .A(n17880), .B(n17881), .Z(n17879) );
  NANDN U17599 ( .A(n17882), .B(n17883), .Z(n17878) );
  NANDN U17600 ( .A(n17881), .B(n17880), .Z(n17883) );
  ANDN U17601 ( .B(\stack[0][25] ), .A(n5340), .Z(n17699) );
  XNOR U17602 ( .A(n17705), .B(n17884), .Z(n17698) );
  XNOR U17603 ( .A(n17706), .B(n17707), .Z(n17884) );
  AND U17604 ( .A(n17885), .B(n17886), .Z(n17707) );
  NAND U17605 ( .A(n17887), .B(n17888), .Z(n17886) );
  NANDN U17606 ( .A(n17889), .B(n17890), .Z(n17885) );
  OR U17607 ( .A(n17887), .B(n17888), .Z(n17890) );
  ANDN U17608 ( .B(\stack[0][24] ), .A(n5364), .Z(n17706) );
  XNOR U17609 ( .A(n17712), .B(n17891), .Z(n17705) );
  XNOR U17610 ( .A(n17713), .B(n17714), .Z(n17891) );
  AND U17611 ( .A(n17892), .B(n17893), .Z(n17714) );
  NANDN U17612 ( .A(n17894), .B(n17895), .Z(n17893) );
  NANDN U17613 ( .A(n17896), .B(n17897), .Z(n17892) );
  NANDN U17614 ( .A(n17895), .B(n17894), .Z(n17897) );
  ANDN U17615 ( .B(\stack[0][23] ), .A(n5387), .Z(n17713) );
  XNOR U17616 ( .A(n17719), .B(n17898), .Z(n17712) );
  XNOR U17617 ( .A(n17720), .B(n17721), .Z(n17898) );
  AND U17618 ( .A(n17899), .B(n17900), .Z(n17721) );
  NAND U17619 ( .A(n17901), .B(n17902), .Z(n17900) );
  NANDN U17620 ( .A(n17903), .B(n17904), .Z(n17899) );
  OR U17621 ( .A(n17901), .B(n17902), .Z(n17904) );
  ANDN U17622 ( .B(\stack[1][10] ), .A(n5686), .Z(n17720) );
  XNOR U17623 ( .A(n17726), .B(n17905), .Z(n17719) );
  XNOR U17624 ( .A(n17727), .B(n17728), .Z(n17905) );
  AND U17625 ( .A(n17906), .B(n17907), .Z(n17728) );
  NANDN U17626 ( .A(n17908), .B(n17909), .Z(n17907) );
  NANDN U17627 ( .A(n17910), .B(n17911), .Z(n17906) );
  NANDN U17628 ( .A(n17909), .B(n17908), .Z(n17911) );
  ANDN U17629 ( .B(\stack[1][11] ), .A(n5662), .Z(n17727) );
  XNOR U17630 ( .A(n17733), .B(n17912), .Z(n17726) );
  XNOR U17631 ( .A(n17734), .B(n17735), .Z(n17912) );
  AND U17632 ( .A(n17913), .B(n17914), .Z(n17735) );
  NAND U17633 ( .A(n17915), .B(n17916), .Z(n17914) );
  NANDN U17634 ( .A(n17917), .B(n17918), .Z(n17913) );
  OR U17635 ( .A(n17915), .B(n17916), .Z(n17918) );
  ANDN U17636 ( .B(\stack[1][12] ), .A(n5638), .Z(n17734) );
  XNOR U17637 ( .A(n17740), .B(n17919), .Z(n17733) );
  XNOR U17638 ( .A(n17741), .B(n17742), .Z(n17919) );
  AND U17639 ( .A(n17920), .B(n17921), .Z(n17742) );
  NANDN U17640 ( .A(n17922), .B(n17923), .Z(n17921) );
  NANDN U17641 ( .A(n17924), .B(n17925), .Z(n17920) );
  NANDN U17642 ( .A(n17923), .B(n17922), .Z(n17925) );
  ANDN U17643 ( .B(\stack[1][13] ), .A(n5614), .Z(n17741) );
  XNOR U17644 ( .A(n17747), .B(n17926), .Z(n17740) );
  XNOR U17645 ( .A(n17748), .B(n17749), .Z(n17926) );
  AND U17646 ( .A(n17927), .B(n17928), .Z(n17749) );
  NAND U17647 ( .A(n17929), .B(n17930), .Z(n17928) );
  NANDN U17648 ( .A(n17931), .B(n17932), .Z(n17927) );
  OR U17649 ( .A(n17929), .B(n17930), .Z(n17932) );
  ANDN U17650 ( .B(\stack[1][14] ), .A(n5590), .Z(n17748) );
  XNOR U17651 ( .A(n17754), .B(n17933), .Z(n17747) );
  XNOR U17652 ( .A(n17755), .B(n17756), .Z(n17933) );
  AND U17653 ( .A(n17934), .B(n17935), .Z(n17756) );
  NANDN U17654 ( .A(n17936), .B(n17937), .Z(n17935) );
  NANDN U17655 ( .A(n17938), .B(n17939), .Z(n17934) );
  NANDN U17656 ( .A(n17937), .B(n17936), .Z(n17939) );
  ANDN U17657 ( .B(\stack[1][15] ), .A(n5566), .Z(n17755) );
  XNOR U17658 ( .A(n17761), .B(n17940), .Z(n17754) );
  XNOR U17659 ( .A(n17762), .B(n17763), .Z(n17940) );
  AND U17660 ( .A(n17941), .B(n17942), .Z(n17763) );
  NAND U17661 ( .A(n17943), .B(n17944), .Z(n17942) );
  NANDN U17662 ( .A(n17945), .B(n17946), .Z(n17941) );
  OR U17663 ( .A(n17943), .B(n17944), .Z(n17946) );
  ANDN U17664 ( .B(\stack[1][16] ), .A(n5542), .Z(n17762) );
  XNOR U17665 ( .A(n17768), .B(n17947), .Z(n17761) );
  XNOR U17666 ( .A(n17769), .B(n17770), .Z(n17947) );
  AND U17667 ( .A(n17948), .B(n17949), .Z(n17770) );
  NANDN U17668 ( .A(n17950), .B(n17951), .Z(n17949) );
  NANDN U17669 ( .A(n17952), .B(n17953), .Z(n17948) );
  NANDN U17670 ( .A(n17951), .B(n17950), .Z(n17953) );
  ANDN U17671 ( .B(\stack[1][17] ), .A(n5518), .Z(n17769) );
  XNOR U17672 ( .A(n17775), .B(n17954), .Z(n17768) );
  XNOR U17673 ( .A(n17776), .B(n17777), .Z(n17954) );
  AND U17674 ( .A(n17955), .B(n17956), .Z(n17777) );
  NAND U17675 ( .A(n17957), .B(n17958), .Z(n17956) );
  NANDN U17676 ( .A(n17959), .B(n17960), .Z(n17955) );
  OR U17677 ( .A(n17957), .B(n17958), .Z(n17960) );
  ANDN U17678 ( .B(\stack[1][18] ), .A(n5494), .Z(n17776) );
  XNOR U17679 ( .A(n17782), .B(n17961), .Z(n17775) );
  XNOR U17680 ( .A(n17783), .B(n17784), .Z(n17961) );
  AND U17681 ( .A(n17962), .B(n17963), .Z(n17784) );
  NANDN U17682 ( .A(n17964), .B(n17965), .Z(n17963) );
  NANDN U17683 ( .A(n17966), .B(n17967), .Z(n17962) );
  NANDN U17684 ( .A(n17965), .B(n17964), .Z(n17967) );
  ANDN U17685 ( .B(\stack[1][19] ), .A(n5470), .Z(n17783) );
  XNOR U17686 ( .A(n17789), .B(n17968), .Z(n17782) );
  XNOR U17687 ( .A(n17790), .B(n17791), .Z(n17968) );
  AND U17688 ( .A(n17969), .B(n17970), .Z(n17791) );
  NAND U17689 ( .A(n17971), .B(n17972), .Z(n17970) );
  NANDN U17690 ( .A(n17973), .B(n17974), .Z(n17969) );
  OR U17691 ( .A(n17971), .B(n17972), .Z(n17974) );
  ANDN U17692 ( .B(\stack[1][20] ), .A(n5446), .Z(n17790) );
  XNOR U17693 ( .A(n17796), .B(n17975), .Z(n17789) );
  XNOR U17694 ( .A(n17797), .B(n17798), .Z(n17975) );
  AND U17695 ( .A(n17976), .B(n17977), .Z(n17798) );
  NANDN U17696 ( .A(n17978), .B(n17979), .Z(n17977) );
  NANDN U17697 ( .A(n17980), .B(n17981), .Z(n17976) );
  NANDN U17698 ( .A(n17979), .B(n17978), .Z(n17981) );
  ANDN U17699 ( .B(\stack[1][21] ), .A(n5422), .Z(n17797) );
  XNOR U17700 ( .A(n17803), .B(n17982), .Z(n17796) );
  XNOR U17701 ( .A(n17804), .B(n17805), .Z(n17982) );
  AND U17702 ( .A(n17983), .B(n17984), .Z(n17805) );
  NAND U17703 ( .A(n17985), .B(n17986), .Z(n17984) );
  NANDN U17704 ( .A(n17987), .B(n17988), .Z(n17983) );
  OR U17705 ( .A(n17985), .B(n17986), .Z(n17988) );
  ANDN U17706 ( .B(\stack[1][22] ), .A(n5398), .Z(n17804) );
  XNOR U17707 ( .A(n17810), .B(n17989), .Z(n17803) );
  XNOR U17708 ( .A(n17811), .B(n17812), .Z(n17989) );
  AND U17709 ( .A(n17990), .B(n17991), .Z(n17812) );
  NANDN U17710 ( .A(n17992), .B(n17993), .Z(n17991) );
  NANDN U17711 ( .A(n17994), .B(n17995), .Z(n17990) );
  NANDN U17712 ( .A(n17993), .B(n17992), .Z(n17995) );
  ANDN U17713 ( .B(\stack[1][23] ), .A(n5374), .Z(n17811) );
  XNOR U17714 ( .A(n17817), .B(n17996), .Z(n17810) );
  XNOR U17715 ( .A(n17818), .B(n17819), .Z(n17996) );
  AND U17716 ( .A(n17997), .B(n17998), .Z(n17819) );
  NAND U17717 ( .A(n17999), .B(n18000), .Z(n17998) );
  NANDN U17718 ( .A(n18001), .B(n18002), .Z(n17997) );
  OR U17719 ( .A(n17999), .B(n18000), .Z(n18002) );
  ANDN U17720 ( .B(\stack[1][24] ), .A(n5350), .Z(n17818) );
  XNOR U17721 ( .A(n17824), .B(n18003), .Z(n17817) );
  XNOR U17722 ( .A(n17825), .B(n17826), .Z(n18003) );
  AND U17723 ( .A(n18004), .B(n18005), .Z(n17826) );
  NANDN U17724 ( .A(n18006), .B(n18007), .Z(n18005) );
  NANDN U17725 ( .A(n18008), .B(n18009), .Z(n18004) );
  NANDN U17726 ( .A(n18007), .B(n18006), .Z(n18009) );
  ANDN U17727 ( .B(\stack[1][25] ), .A(n5326), .Z(n17825) );
  XNOR U17728 ( .A(n17831), .B(n18010), .Z(n17824) );
  XNOR U17729 ( .A(n17832), .B(n17833), .Z(n18010) );
  AND U17730 ( .A(n18011), .B(n18012), .Z(n17833) );
  NAND U17731 ( .A(n18013), .B(n18014), .Z(n18012) );
  NANDN U17732 ( .A(n18015), .B(n18016), .Z(n18011) );
  OR U17733 ( .A(n18013), .B(n18014), .Z(n18016) );
  ANDN U17734 ( .B(\stack[1][26] ), .A(n5302), .Z(n17832) );
  XNOR U17735 ( .A(n17838), .B(n18017), .Z(n17831) );
  XNOR U17736 ( .A(n17839), .B(n17840), .Z(n18017) );
  AND U17737 ( .A(n18018), .B(n18019), .Z(n17840) );
  NANDN U17738 ( .A(n18020), .B(n18021), .Z(n18019) );
  NANDN U17739 ( .A(n18022), .B(n18023), .Z(n18018) );
  NANDN U17740 ( .A(n18021), .B(n18020), .Z(n18023) );
  ANDN U17741 ( .B(\stack[1][27] ), .A(n5278), .Z(n17839) );
  XNOR U17742 ( .A(n17845), .B(n18024), .Z(n17838) );
  XNOR U17743 ( .A(n17846), .B(n17847), .Z(n18024) );
  AND U17744 ( .A(n18025), .B(n18026), .Z(n17847) );
  NAND U17745 ( .A(n18027), .B(n18028), .Z(n18026) );
  NANDN U17746 ( .A(n18029), .B(n18030), .Z(n18025) );
  OR U17747 ( .A(n18027), .B(n18028), .Z(n18030) );
  ANDN U17748 ( .B(\stack[1][28] ), .A(n5254), .Z(n17846) );
  XNOR U17749 ( .A(n17852), .B(n18031), .Z(n17845) );
  XNOR U17750 ( .A(n17853), .B(n17854), .Z(n18031) );
  AND U17751 ( .A(n18032), .B(n18033), .Z(n17854) );
  NAND U17752 ( .A(n18034), .B(n18035), .Z(n18033) );
  NAND U17753 ( .A(n18036), .B(n18037), .Z(n18032) );
  OR U17754 ( .A(n18034), .B(n18035), .Z(n18036) );
  ANDN U17755 ( .B(\stack[1][29] ), .A(n5230), .Z(n17853) );
  XNOR U17756 ( .A(n17859), .B(n18038), .Z(n17852) );
  XNOR U17757 ( .A(n17860), .B(n17862), .Z(n18038) );
  ANDN U17758 ( .B(n18039), .A(n18040), .Z(n17862) );
  ANDN U17759 ( .B(\stack[0][0] ), .A(n5915), .Z(n18039) );
  ANDN U17760 ( .B(\stack[1][30] ), .A(n5206), .Z(n17860) );
  XOR U17761 ( .A(n17865), .B(n18041), .Z(n17859) );
  NANDN U17762 ( .A(n5160), .B(\stack[1][32] ), .Z(n18041) );
  NANDN U17763 ( .A(n5915), .B(\stack[0][1] ), .Z(n17865) );
  ANDN U17764 ( .B(\stack[0][27] ), .A(n5292), .Z(n9174) );
  AND U17765 ( .A(n18042), .B(n18043), .Z(n9175) );
  NANDN U17766 ( .A(n9182), .B(n18044), .Z(n18042) );
  NANDN U17767 ( .A(n9181), .B(n9179), .Z(n18044) );
  XNOR U17768 ( .A(n17873), .B(n18045), .Z(n9179) );
  XNOR U17769 ( .A(n17874), .B(n17875), .Z(n18045) );
  AND U17770 ( .A(n18046), .B(n18047), .Z(n17875) );
  NANDN U17771 ( .A(n18048), .B(n18049), .Z(n18047) );
  NANDN U17772 ( .A(n18050), .B(n18051), .Z(n18046) );
  NANDN U17773 ( .A(n18049), .B(n18048), .Z(n18051) );
  ANDN U17774 ( .B(\stack[0][25] ), .A(n5316), .Z(n17874) );
  XNOR U17775 ( .A(n17880), .B(n18052), .Z(n17873) );
  XNOR U17776 ( .A(n17881), .B(n17882), .Z(n18052) );
  AND U17777 ( .A(n18053), .B(n18054), .Z(n17882) );
  NAND U17778 ( .A(n18055), .B(n18056), .Z(n18054) );
  NANDN U17779 ( .A(n18057), .B(n18058), .Z(n18053) );
  OR U17780 ( .A(n18055), .B(n18056), .Z(n18058) );
  ANDN U17781 ( .B(\stack[0][24] ), .A(n5340), .Z(n17881) );
  XNOR U17782 ( .A(n17887), .B(n18059), .Z(n17880) );
  XNOR U17783 ( .A(n17888), .B(n17889), .Z(n18059) );
  AND U17784 ( .A(n18060), .B(n18061), .Z(n17889) );
  NANDN U17785 ( .A(n18062), .B(n18063), .Z(n18061) );
  NANDN U17786 ( .A(n18064), .B(n18065), .Z(n18060) );
  NANDN U17787 ( .A(n18063), .B(n18062), .Z(n18065) );
  ANDN U17788 ( .B(\stack[0][23] ), .A(n5364), .Z(n17888) );
  XNOR U17789 ( .A(n17894), .B(n18066), .Z(n17887) );
  XNOR U17790 ( .A(n17895), .B(n17896), .Z(n18066) );
  AND U17791 ( .A(n18067), .B(n18068), .Z(n17896) );
  NAND U17792 ( .A(n18069), .B(n18070), .Z(n18068) );
  NANDN U17793 ( .A(n18071), .B(n18072), .Z(n18067) );
  OR U17794 ( .A(n18069), .B(n18070), .Z(n18072) );
  ANDN U17795 ( .B(\stack[0][22] ), .A(n5387), .Z(n17895) );
  XNOR U17796 ( .A(n17901), .B(n18073), .Z(n17894) );
  XNOR U17797 ( .A(n17902), .B(n17903), .Z(n18073) );
  AND U17798 ( .A(n18074), .B(n18075), .Z(n17903) );
  NANDN U17799 ( .A(n18076), .B(n18077), .Z(n18075) );
  NANDN U17800 ( .A(n18078), .B(n18079), .Z(n18074) );
  NANDN U17801 ( .A(n18077), .B(n18076), .Z(n18079) );
  ANDN U17802 ( .B(\stack[1][10] ), .A(n5662), .Z(n17902) );
  XNOR U17803 ( .A(n17908), .B(n18080), .Z(n17901) );
  XNOR U17804 ( .A(n17909), .B(n17910), .Z(n18080) );
  AND U17805 ( .A(n18081), .B(n18082), .Z(n17910) );
  NAND U17806 ( .A(n18083), .B(n18084), .Z(n18082) );
  NANDN U17807 ( .A(n18085), .B(n18086), .Z(n18081) );
  OR U17808 ( .A(n18083), .B(n18084), .Z(n18086) );
  ANDN U17809 ( .B(\stack[1][11] ), .A(n5638), .Z(n17909) );
  XNOR U17810 ( .A(n17915), .B(n18087), .Z(n17908) );
  XNOR U17811 ( .A(n17916), .B(n17917), .Z(n18087) );
  AND U17812 ( .A(n18088), .B(n18089), .Z(n17917) );
  NANDN U17813 ( .A(n18090), .B(n18091), .Z(n18089) );
  NANDN U17814 ( .A(n18092), .B(n18093), .Z(n18088) );
  NANDN U17815 ( .A(n18091), .B(n18090), .Z(n18093) );
  ANDN U17816 ( .B(\stack[1][12] ), .A(n5614), .Z(n17916) );
  XNOR U17817 ( .A(n17922), .B(n18094), .Z(n17915) );
  XNOR U17818 ( .A(n17923), .B(n17924), .Z(n18094) );
  AND U17819 ( .A(n18095), .B(n18096), .Z(n17924) );
  NAND U17820 ( .A(n18097), .B(n18098), .Z(n18096) );
  NANDN U17821 ( .A(n18099), .B(n18100), .Z(n18095) );
  OR U17822 ( .A(n18097), .B(n18098), .Z(n18100) );
  ANDN U17823 ( .B(\stack[1][13] ), .A(n5590), .Z(n17923) );
  XNOR U17824 ( .A(n17929), .B(n18101), .Z(n17922) );
  XNOR U17825 ( .A(n17930), .B(n17931), .Z(n18101) );
  AND U17826 ( .A(n18102), .B(n18103), .Z(n17931) );
  NANDN U17827 ( .A(n18104), .B(n18105), .Z(n18103) );
  NANDN U17828 ( .A(n18106), .B(n18107), .Z(n18102) );
  NANDN U17829 ( .A(n18105), .B(n18104), .Z(n18107) );
  ANDN U17830 ( .B(\stack[1][14] ), .A(n5566), .Z(n17930) );
  XNOR U17831 ( .A(n17936), .B(n18108), .Z(n17929) );
  XNOR U17832 ( .A(n17937), .B(n17938), .Z(n18108) );
  AND U17833 ( .A(n18109), .B(n18110), .Z(n17938) );
  NAND U17834 ( .A(n18111), .B(n18112), .Z(n18110) );
  NANDN U17835 ( .A(n18113), .B(n18114), .Z(n18109) );
  OR U17836 ( .A(n18111), .B(n18112), .Z(n18114) );
  ANDN U17837 ( .B(\stack[1][15] ), .A(n5542), .Z(n17937) );
  XNOR U17838 ( .A(n17943), .B(n18115), .Z(n17936) );
  XNOR U17839 ( .A(n17944), .B(n17945), .Z(n18115) );
  AND U17840 ( .A(n18116), .B(n18117), .Z(n17945) );
  NANDN U17841 ( .A(n18118), .B(n18119), .Z(n18117) );
  NANDN U17842 ( .A(n18120), .B(n18121), .Z(n18116) );
  NANDN U17843 ( .A(n18119), .B(n18118), .Z(n18121) );
  ANDN U17844 ( .B(\stack[1][16] ), .A(n5518), .Z(n17944) );
  XNOR U17845 ( .A(n17950), .B(n18122), .Z(n17943) );
  XNOR U17846 ( .A(n17951), .B(n17952), .Z(n18122) );
  AND U17847 ( .A(n18123), .B(n18124), .Z(n17952) );
  NAND U17848 ( .A(n18125), .B(n18126), .Z(n18124) );
  NANDN U17849 ( .A(n18127), .B(n18128), .Z(n18123) );
  OR U17850 ( .A(n18125), .B(n18126), .Z(n18128) );
  ANDN U17851 ( .B(\stack[1][17] ), .A(n5494), .Z(n17951) );
  XNOR U17852 ( .A(n17957), .B(n18129), .Z(n17950) );
  XNOR U17853 ( .A(n17958), .B(n17959), .Z(n18129) );
  AND U17854 ( .A(n18130), .B(n18131), .Z(n17959) );
  NANDN U17855 ( .A(n18132), .B(n18133), .Z(n18131) );
  NANDN U17856 ( .A(n18134), .B(n18135), .Z(n18130) );
  NANDN U17857 ( .A(n18133), .B(n18132), .Z(n18135) );
  ANDN U17858 ( .B(\stack[1][18] ), .A(n5470), .Z(n17958) );
  XNOR U17859 ( .A(n17964), .B(n18136), .Z(n17957) );
  XNOR U17860 ( .A(n17965), .B(n17966), .Z(n18136) );
  AND U17861 ( .A(n18137), .B(n18138), .Z(n17966) );
  NAND U17862 ( .A(n18139), .B(n18140), .Z(n18138) );
  NANDN U17863 ( .A(n18141), .B(n18142), .Z(n18137) );
  OR U17864 ( .A(n18139), .B(n18140), .Z(n18142) );
  ANDN U17865 ( .B(\stack[1][19] ), .A(n5446), .Z(n17965) );
  XNOR U17866 ( .A(n17971), .B(n18143), .Z(n17964) );
  XNOR U17867 ( .A(n17972), .B(n17973), .Z(n18143) );
  AND U17868 ( .A(n18144), .B(n18145), .Z(n17973) );
  NANDN U17869 ( .A(n18146), .B(n18147), .Z(n18145) );
  NANDN U17870 ( .A(n18148), .B(n18149), .Z(n18144) );
  NANDN U17871 ( .A(n18147), .B(n18146), .Z(n18149) );
  ANDN U17872 ( .B(\stack[1][20] ), .A(n5422), .Z(n17972) );
  XNOR U17873 ( .A(n17978), .B(n18150), .Z(n17971) );
  XNOR U17874 ( .A(n17979), .B(n17980), .Z(n18150) );
  AND U17875 ( .A(n18151), .B(n18152), .Z(n17980) );
  NAND U17876 ( .A(n18153), .B(n18154), .Z(n18152) );
  NANDN U17877 ( .A(n18155), .B(n18156), .Z(n18151) );
  OR U17878 ( .A(n18153), .B(n18154), .Z(n18156) );
  ANDN U17879 ( .B(\stack[1][21] ), .A(n5398), .Z(n17979) );
  XNOR U17880 ( .A(n17985), .B(n18157), .Z(n17978) );
  XNOR U17881 ( .A(n17986), .B(n17987), .Z(n18157) );
  AND U17882 ( .A(n18158), .B(n18159), .Z(n17987) );
  NANDN U17883 ( .A(n18160), .B(n18161), .Z(n18159) );
  NANDN U17884 ( .A(n18162), .B(n18163), .Z(n18158) );
  NANDN U17885 ( .A(n18161), .B(n18160), .Z(n18163) );
  ANDN U17886 ( .B(\stack[1][22] ), .A(n5374), .Z(n17986) );
  XNOR U17887 ( .A(n17992), .B(n18164), .Z(n17985) );
  XNOR U17888 ( .A(n17993), .B(n17994), .Z(n18164) );
  AND U17889 ( .A(n18165), .B(n18166), .Z(n17994) );
  NAND U17890 ( .A(n18167), .B(n18168), .Z(n18166) );
  NANDN U17891 ( .A(n18169), .B(n18170), .Z(n18165) );
  OR U17892 ( .A(n18167), .B(n18168), .Z(n18170) );
  ANDN U17893 ( .B(\stack[1][23] ), .A(n5350), .Z(n17993) );
  XNOR U17894 ( .A(n17999), .B(n18171), .Z(n17992) );
  XNOR U17895 ( .A(n18000), .B(n18001), .Z(n18171) );
  AND U17896 ( .A(n18172), .B(n18173), .Z(n18001) );
  NANDN U17897 ( .A(n18174), .B(n18175), .Z(n18173) );
  NANDN U17898 ( .A(n18176), .B(n18177), .Z(n18172) );
  NANDN U17899 ( .A(n18175), .B(n18174), .Z(n18177) );
  ANDN U17900 ( .B(\stack[1][24] ), .A(n5326), .Z(n18000) );
  XNOR U17901 ( .A(n18006), .B(n18178), .Z(n17999) );
  XNOR U17902 ( .A(n18007), .B(n18008), .Z(n18178) );
  AND U17903 ( .A(n18179), .B(n18180), .Z(n18008) );
  NAND U17904 ( .A(n18181), .B(n18182), .Z(n18180) );
  NANDN U17905 ( .A(n18183), .B(n18184), .Z(n18179) );
  OR U17906 ( .A(n18181), .B(n18182), .Z(n18184) );
  ANDN U17907 ( .B(\stack[1][25] ), .A(n5302), .Z(n18007) );
  XNOR U17908 ( .A(n18013), .B(n18185), .Z(n18006) );
  XNOR U17909 ( .A(n18014), .B(n18015), .Z(n18185) );
  AND U17910 ( .A(n18186), .B(n18187), .Z(n18015) );
  NANDN U17911 ( .A(n18188), .B(n18189), .Z(n18187) );
  NANDN U17912 ( .A(n18190), .B(n18191), .Z(n18186) );
  NANDN U17913 ( .A(n18189), .B(n18188), .Z(n18191) );
  ANDN U17914 ( .B(\stack[1][26] ), .A(n5278), .Z(n18014) );
  XNOR U17915 ( .A(n18020), .B(n18192), .Z(n18013) );
  XNOR U17916 ( .A(n18021), .B(n18022), .Z(n18192) );
  AND U17917 ( .A(n18193), .B(n18194), .Z(n18022) );
  NAND U17918 ( .A(n18195), .B(n18196), .Z(n18194) );
  NANDN U17919 ( .A(n18197), .B(n18198), .Z(n18193) );
  OR U17920 ( .A(n18195), .B(n18196), .Z(n18198) );
  ANDN U17921 ( .B(\stack[1][27] ), .A(n5254), .Z(n18021) );
  XNOR U17922 ( .A(n18027), .B(n18199), .Z(n18020) );
  XNOR U17923 ( .A(n18028), .B(n18029), .Z(n18199) );
  AND U17924 ( .A(n18200), .B(n18201), .Z(n18029) );
  NAND U17925 ( .A(n18202), .B(n18203), .Z(n18201) );
  NAND U17926 ( .A(n18204), .B(n18205), .Z(n18200) );
  OR U17927 ( .A(n18202), .B(n18203), .Z(n18204) );
  ANDN U17928 ( .B(\stack[1][28] ), .A(n5230), .Z(n18028) );
  XNOR U17929 ( .A(n18034), .B(n18206), .Z(n18027) );
  XNOR U17930 ( .A(n18035), .B(n18037), .Z(n18206) );
  ANDN U17931 ( .B(n18207), .A(n18208), .Z(n18037) );
  ANDN U17932 ( .B(\stack[0][0] ), .A(n5891), .Z(n18207) );
  ANDN U17933 ( .B(\stack[1][29] ), .A(n5206), .Z(n18035) );
  XOR U17934 ( .A(n18040), .B(n18209), .Z(n18034) );
  NANDN U17935 ( .A(n5160), .B(\stack[1][31] ), .Z(n18209) );
  NANDN U17936 ( .A(n5891), .B(\stack[0][1] ), .Z(n18040) );
  ANDN U17937 ( .B(\stack[1][5] ), .A(n5782), .Z(n9181) );
  AND U17938 ( .A(n18210), .B(n18211), .Z(n9182) );
  NANDN U17939 ( .A(n9186), .B(n9188), .Z(n18211) );
  NANDN U17940 ( .A(n9189), .B(n18212), .Z(n18210) );
  NANDN U17941 ( .A(n9188), .B(n9186), .Z(n18212) );
  XOR U17942 ( .A(n18048), .B(n18213), .Z(n9186) );
  XNOR U17943 ( .A(n18049), .B(n18050), .Z(n18213) );
  AND U17944 ( .A(n18214), .B(n18215), .Z(n18050) );
  NAND U17945 ( .A(n18216), .B(n18217), .Z(n18215) );
  NANDN U17946 ( .A(n18218), .B(n18219), .Z(n18214) );
  OR U17947 ( .A(n18216), .B(n18217), .Z(n18219) );
  ANDN U17948 ( .B(\stack[0][24] ), .A(n5316), .Z(n18049) );
  XNOR U17949 ( .A(n18055), .B(n18220), .Z(n18048) );
  XNOR U17950 ( .A(n18056), .B(n18057), .Z(n18220) );
  AND U17951 ( .A(n18221), .B(n18222), .Z(n18057) );
  NANDN U17952 ( .A(n18223), .B(n18224), .Z(n18222) );
  NANDN U17953 ( .A(n18225), .B(n18226), .Z(n18221) );
  NANDN U17954 ( .A(n18224), .B(n18223), .Z(n18226) );
  ANDN U17955 ( .B(\stack[0][23] ), .A(n5340), .Z(n18056) );
  XNOR U17956 ( .A(n18062), .B(n18227), .Z(n18055) );
  XNOR U17957 ( .A(n18063), .B(n18064), .Z(n18227) );
  AND U17958 ( .A(n18228), .B(n18229), .Z(n18064) );
  NAND U17959 ( .A(n18230), .B(n18231), .Z(n18229) );
  NANDN U17960 ( .A(n18232), .B(n18233), .Z(n18228) );
  OR U17961 ( .A(n18230), .B(n18231), .Z(n18233) );
  ANDN U17962 ( .B(\stack[0][22] ), .A(n5364), .Z(n18063) );
  XNOR U17963 ( .A(n18069), .B(n18234), .Z(n18062) );
  XNOR U17964 ( .A(n18070), .B(n18071), .Z(n18234) );
  AND U17965 ( .A(n18235), .B(n18236), .Z(n18071) );
  NANDN U17966 ( .A(n18237), .B(n18238), .Z(n18236) );
  NANDN U17967 ( .A(n18239), .B(n18240), .Z(n18235) );
  NANDN U17968 ( .A(n18238), .B(n18237), .Z(n18240) );
  ANDN U17969 ( .B(\stack[0][21] ), .A(n5387), .Z(n18070) );
  XNOR U17970 ( .A(n18076), .B(n18241), .Z(n18069) );
  XNOR U17971 ( .A(n18077), .B(n18078), .Z(n18241) );
  AND U17972 ( .A(n18242), .B(n18243), .Z(n18078) );
  NAND U17973 ( .A(n18244), .B(n18245), .Z(n18243) );
  NANDN U17974 ( .A(n18246), .B(n18247), .Z(n18242) );
  OR U17975 ( .A(n18244), .B(n18245), .Z(n18247) );
  ANDN U17976 ( .B(\stack[1][10] ), .A(n5638), .Z(n18077) );
  XNOR U17977 ( .A(n18083), .B(n18248), .Z(n18076) );
  XNOR U17978 ( .A(n18084), .B(n18085), .Z(n18248) );
  AND U17979 ( .A(n18249), .B(n18250), .Z(n18085) );
  NANDN U17980 ( .A(n18251), .B(n18252), .Z(n18250) );
  NANDN U17981 ( .A(n18253), .B(n18254), .Z(n18249) );
  NANDN U17982 ( .A(n18252), .B(n18251), .Z(n18254) );
  ANDN U17983 ( .B(\stack[1][11] ), .A(n5614), .Z(n18084) );
  XNOR U17984 ( .A(n18090), .B(n18255), .Z(n18083) );
  XNOR U17985 ( .A(n18091), .B(n18092), .Z(n18255) );
  AND U17986 ( .A(n18256), .B(n18257), .Z(n18092) );
  NAND U17987 ( .A(n18258), .B(n18259), .Z(n18257) );
  NANDN U17988 ( .A(n18260), .B(n18261), .Z(n18256) );
  OR U17989 ( .A(n18258), .B(n18259), .Z(n18261) );
  ANDN U17990 ( .B(\stack[1][12] ), .A(n5590), .Z(n18091) );
  XNOR U17991 ( .A(n18097), .B(n18262), .Z(n18090) );
  XNOR U17992 ( .A(n18098), .B(n18099), .Z(n18262) );
  AND U17993 ( .A(n18263), .B(n18264), .Z(n18099) );
  NANDN U17994 ( .A(n18265), .B(n18266), .Z(n18264) );
  NANDN U17995 ( .A(n18267), .B(n18268), .Z(n18263) );
  NANDN U17996 ( .A(n18266), .B(n18265), .Z(n18268) );
  ANDN U17997 ( .B(\stack[1][13] ), .A(n5566), .Z(n18098) );
  XNOR U17998 ( .A(n18104), .B(n18269), .Z(n18097) );
  XNOR U17999 ( .A(n18105), .B(n18106), .Z(n18269) );
  AND U18000 ( .A(n18270), .B(n18271), .Z(n18106) );
  NAND U18001 ( .A(n18272), .B(n18273), .Z(n18271) );
  NANDN U18002 ( .A(n18274), .B(n18275), .Z(n18270) );
  OR U18003 ( .A(n18272), .B(n18273), .Z(n18275) );
  ANDN U18004 ( .B(\stack[1][14] ), .A(n5542), .Z(n18105) );
  XNOR U18005 ( .A(n18111), .B(n18276), .Z(n18104) );
  XNOR U18006 ( .A(n18112), .B(n18113), .Z(n18276) );
  AND U18007 ( .A(n18277), .B(n18278), .Z(n18113) );
  NANDN U18008 ( .A(n18279), .B(n18280), .Z(n18278) );
  NANDN U18009 ( .A(n18281), .B(n18282), .Z(n18277) );
  NANDN U18010 ( .A(n18280), .B(n18279), .Z(n18282) );
  ANDN U18011 ( .B(\stack[1][15] ), .A(n5518), .Z(n18112) );
  XNOR U18012 ( .A(n18118), .B(n18283), .Z(n18111) );
  XNOR U18013 ( .A(n18119), .B(n18120), .Z(n18283) );
  AND U18014 ( .A(n18284), .B(n18285), .Z(n18120) );
  NAND U18015 ( .A(n18286), .B(n18287), .Z(n18285) );
  NANDN U18016 ( .A(n18288), .B(n18289), .Z(n18284) );
  OR U18017 ( .A(n18286), .B(n18287), .Z(n18289) );
  ANDN U18018 ( .B(\stack[1][16] ), .A(n5494), .Z(n18119) );
  XNOR U18019 ( .A(n18125), .B(n18290), .Z(n18118) );
  XNOR U18020 ( .A(n18126), .B(n18127), .Z(n18290) );
  AND U18021 ( .A(n18291), .B(n18292), .Z(n18127) );
  NANDN U18022 ( .A(n18293), .B(n18294), .Z(n18292) );
  NANDN U18023 ( .A(n18295), .B(n18296), .Z(n18291) );
  NANDN U18024 ( .A(n18294), .B(n18293), .Z(n18296) );
  ANDN U18025 ( .B(\stack[1][17] ), .A(n5470), .Z(n18126) );
  XNOR U18026 ( .A(n18132), .B(n18297), .Z(n18125) );
  XNOR U18027 ( .A(n18133), .B(n18134), .Z(n18297) );
  AND U18028 ( .A(n18298), .B(n18299), .Z(n18134) );
  NAND U18029 ( .A(n18300), .B(n18301), .Z(n18299) );
  NANDN U18030 ( .A(n18302), .B(n18303), .Z(n18298) );
  OR U18031 ( .A(n18300), .B(n18301), .Z(n18303) );
  ANDN U18032 ( .B(\stack[1][18] ), .A(n5446), .Z(n18133) );
  XNOR U18033 ( .A(n18139), .B(n18304), .Z(n18132) );
  XNOR U18034 ( .A(n18140), .B(n18141), .Z(n18304) );
  AND U18035 ( .A(n18305), .B(n18306), .Z(n18141) );
  NANDN U18036 ( .A(n18307), .B(n18308), .Z(n18306) );
  NANDN U18037 ( .A(n18309), .B(n18310), .Z(n18305) );
  NANDN U18038 ( .A(n18308), .B(n18307), .Z(n18310) );
  ANDN U18039 ( .B(\stack[1][19] ), .A(n5422), .Z(n18140) );
  XNOR U18040 ( .A(n18146), .B(n18311), .Z(n18139) );
  XNOR U18041 ( .A(n18147), .B(n18148), .Z(n18311) );
  AND U18042 ( .A(n18312), .B(n18313), .Z(n18148) );
  NAND U18043 ( .A(n18314), .B(n18315), .Z(n18313) );
  NANDN U18044 ( .A(n18316), .B(n18317), .Z(n18312) );
  OR U18045 ( .A(n18314), .B(n18315), .Z(n18317) );
  ANDN U18046 ( .B(\stack[1][20] ), .A(n5398), .Z(n18147) );
  XNOR U18047 ( .A(n18153), .B(n18318), .Z(n18146) );
  XNOR U18048 ( .A(n18154), .B(n18155), .Z(n18318) );
  AND U18049 ( .A(n18319), .B(n18320), .Z(n18155) );
  NANDN U18050 ( .A(n18321), .B(n18322), .Z(n18320) );
  NANDN U18051 ( .A(n18323), .B(n18324), .Z(n18319) );
  NANDN U18052 ( .A(n18322), .B(n18321), .Z(n18324) );
  ANDN U18053 ( .B(\stack[1][21] ), .A(n5374), .Z(n18154) );
  XNOR U18054 ( .A(n18160), .B(n18325), .Z(n18153) );
  XNOR U18055 ( .A(n18161), .B(n18162), .Z(n18325) );
  AND U18056 ( .A(n18326), .B(n18327), .Z(n18162) );
  NAND U18057 ( .A(n18328), .B(n18329), .Z(n18327) );
  NANDN U18058 ( .A(n18330), .B(n18331), .Z(n18326) );
  OR U18059 ( .A(n18328), .B(n18329), .Z(n18331) );
  ANDN U18060 ( .B(\stack[1][22] ), .A(n5350), .Z(n18161) );
  XNOR U18061 ( .A(n18167), .B(n18332), .Z(n18160) );
  XNOR U18062 ( .A(n18168), .B(n18169), .Z(n18332) );
  AND U18063 ( .A(n18333), .B(n18334), .Z(n18169) );
  NANDN U18064 ( .A(n18335), .B(n18336), .Z(n18334) );
  NANDN U18065 ( .A(n18337), .B(n18338), .Z(n18333) );
  NANDN U18066 ( .A(n18336), .B(n18335), .Z(n18338) );
  ANDN U18067 ( .B(\stack[1][23] ), .A(n5326), .Z(n18168) );
  XNOR U18068 ( .A(n18174), .B(n18339), .Z(n18167) );
  XNOR U18069 ( .A(n18175), .B(n18176), .Z(n18339) );
  AND U18070 ( .A(n18340), .B(n18341), .Z(n18176) );
  NAND U18071 ( .A(n18342), .B(n18343), .Z(n18341) );
  NANDN U18072 ( .A(n18344), .B(n18345), .Z(n18340) );
  OR U18073 ( .A(n18342), .B(n18343), .Z(n18345) );
  ANDN U18074 ( .B(\stack[1][24] ), .A(n5302), .Z(n18175) );
  XNOR U18075 ( .A(n18181), .B(n18346), .Z(n18174) );
  XNOR U18076 ( .A(n18182), .B(n18183), .Z(n18346) );
  AND U18077 ( .A(n18347), .B(n18348), .Z(n18183) );
  NANDN U18078 ( .A(n18349), .B(n18350), .Z(n18348) );
  NANDN U18079 ( .A(n18351), .B(n18352), .Z(n18347) );
  NANDN U18080 ( .A(n18350), .B(n18349), .Z(n18352) );
  ANDN U18081 ( .B(\stack[1][25] ), .A(n5278), .Z(n18182) );
  XNOR U18082 ( .A(n18188), .B(n18353), .Z(n18181) );
  XNOR U18083 ( .A(n18189), .B(n18190), .Z(n18353) );
  AND U18084 ( .A(n18354), .B(n18355), .Z(n18190) );
  NAND U18085 ( .A(n18356), .B(n18357), .Z(n18355) );
  NANDN U18086 ( .A(n18358), .B(n18359), .Z(n18354) );
  OR U18087 ( .A(n18356), .B(n18357), .Z(n18359) );
  ANDN U18088 ( .B(\stack[1][26] ), .A(n5254), .Z(n18189) );
  XNOR U18089 ( .A(n18195), .B(n18360), .Z(n18188) );
  XNOR U18090 ( .A(n18196), .B(n18197), .Z(n18360) );
  AND U18091 ( .A(n18361), .B(n18362), .Z(n18197) );
  NAND U18092 ( .A(n18363), .B(n18364), .Z(n18362) );
  NAND U18093 ( .A(n18365), .B(n18366), .Z(n18361) );
  OR U18094 ( .A(n18363), .B(n18364), .Z(n18365) );
  ANDN U18095 ( .B(\stack[1][27] ), .A(n5230), .Z(n18196) );
  XNOR U18096 ( .A(n18202), .B(n18367), .Z(n18195) );
  XNOR U18097 ( .A(n18203), .B(n18205), .Z(n18367) );
  ANDN U18098 ( .B(n18368), .A(n18369), .Z(n18205) );
  ANDN U18099 ( .B(\stack[0][0] ), .A(n5867), .Z(n18368) );
  ANDN U18100 ( .B(\stack[1][28] ), .A(n5206), .Z(n18203) );
  XOR U18101 ( .A(n18208), .B(n18370), .Z(n18202) );
  NANDN U18102 ( .A(n5160), .B(\stack[1][30] ), .Z(n18370) );
  NANDN U18103 ( .A(n5867), .B(\stack[0][1] ), .Z(n18208) );
  ANDN U18104 ( .B(\stack[0][25] ), .A(n5292), .Z(n9188) );
  AND U18105 ( .A(n18371), .B(n18372), .Z(n9189) );
  NANDN U18106 ( .A(n9196), .B(n18373), .Z(n18371) );
  NANDN U18107 ( .A(n9195), .B(n9193), .Z(n18373) );
  XNOR U18108 ( .A(n18216), .B(n18374), .Z(n9193) );
  XNOR U18109 ( .A(n18217), .B(n18218), .Z(n18374) );
  AND U18110 ( .A(n18375), .B(n18376), .Z(n18218) );
  NANDN U18111 ( .A(n18377), .B(n18378), .Z(n18376) );
  NANDN U18112 ( .A(n18379), .B(n18380), .Z(n18375) );
  NANDN U18113 ( .A(n18378), .B(n18377), .Z(n18380) );
  ANDN U18114 ( .B(\stack[0][23] ), .A(n5316), .Z(n18217) );
  XNOR U18115 ( .A(n18223), .B(n18381), .Z(n18216) );
  XNOR U18116 ( .A(n18224), .B(n18225), .Z(n18381) );
  AND U18117 ( .A(n18382), .B(n18383), .Z(n18225) );
  NAND U18118 ( .A(n18384), .B(n18385), .Z(n18383) );
  NANDN U18119 ( .A(n18386), .B(n18387), .Z(n18382) );
  OR U18120 ( .A(n18384), .B(n18385), .Z(n18387) );
  ANDN U18121 ( .B(\stack[0][22] ), .A(n5340), .Z(n18224) );
  XNOR U18122 ( .A(n18230), .B(n18388), .Z(n18223) );
  XNOR U18123 ( .A(n18231), .B(n18232), .Z(n18388) );
  AND U18124 ( .A(n18389), .B(n18390), .Z(n18232) );
  NANDN U18125 ( .A(n18391), .B(n18392), .Z(n18390) );
  NANDN U18126 ( .A(n18393), .B(n18394), .Z(n18389) );
  NANDN U18127 ( .A(n18392), .B(n18391), .Z(n18394) );
  ANDN U18128 ( .B(\stack[0][21] ), .A(n5364), .Z(n18231) );
  XNOR U18129 ( .A(n18237), .B(n18395), .Z(n18230) );
  XNOR U18130 ( .A(n18238), .B(n18239), .Z(n18395) );
  AND U18131 ( .A(n18396), .B(n18397), .Z(n18239) );
  NAND U18132 ( .A(n18398), .B(n18399), .Z(n18397) );
  NANDN U18133 ( .A(n18400), .B(n18401), .Z(n18396) );
  OR U18134 ( .A(n18398), .B(n18399), .Z(n18401) );
  ANDN U18135 ( .B(\stack[0][20] ), .A(n5387), .Z(n18238) );
  XNOR U18136 ( .A(n18244), .B(n18402), .Z(n18237) );
  XNOR U18137 ( .A(n18245), .B(n18246), .Z(n18402) );
  AND U18138 ( .A(n18403), .B(n18404), .Z(n18246) );
  NANDN U18139 ( .A(n18405), .B(n18406), .Z(n18404) );
  NANDN U18140 ( .A(n18407), .B(n18408), .Z(n18403) );
  NANDN U18141 ( .A(n18406), .B(n18405), .Z(n18408) );
  ANDN U18142 ( .B(\stack[1][10] ), .A(n5614), .Z(n18245) );
  XNOR U18143 ( .A(n18251), .B(n18409), .Z(n18244) );
  XNOR U18144 ( .A(n18252), .B(n18253), .Z(n18409) );
  AND U18145 ( .A(n18410), .B(n18411), .Z(n18253) );
  NAND U18146 ( .A(n18412), .B(n18413), .Z(n18411) );
  NANDN U18147 ( .A(n18414), .B(n18415), .Z(n18410) );
  OR U18148 ( .A(n18412), .B(n18413), .Z(n18415) );
  ANDN U18149 ( .B(\stack[1][11] ), .A(n5590), .Z(n18252) );
  XNOR U18150 ( .A(n18258), .B(n18416), .Z(n18251) );
  XNOR U18151 ( .A(n18259), .B(n18260), .Z(n18416) );
  AND U18152 ( .A(n18417), .B(n18418), .Z(n18260) );
  NANDN U18153 ( .A(n18419), .B(n18420), .Z(n18418) );
  NANDN U18154 ( .A(n18421), .B(n18422), .Z(n18417) );
  NANDN U18155 ( .A(n18420), .B(n18419), .Z(n18422) );
  ANDN U18156 ( .B(\stack[1][12] ), .A(n5566), .Z(n18259) );
  XNOR U18157 ( .A(n18265), .B(n18423), .Z(n18258) );
  XNOR U18158 ( .A(n18266), .B(n18267), .Z(n18423) );
  AND U18159 ( .A(n18424), .B(n18425), .Z(n18267) );
  NAND U18160 ( .A(n18426), .B(n18427), .Z(n18425) );
  NANDN U18161 ( .A(n18428), .B(n18429), .Z(n18424) );
  OR U18162 ( .A(n18426), .B(n18427), .Z(n18429) );
  ANDN U18163 ( .B(\stack[1][13] ), .A(n5542), .Z(n18266) );
  XNOR U18164 ( .A(n18272), .B(n18430), .Z(n18265) );
  XNOR U18165 ( .A(n18273), .B(n18274), .Z(n18430) );
  AND U18166 ( .A(n18431), .B(n18432), .Z(n18274) );
  NANDN U18167 ( .A(n18433), .B(n18434), .Z(n18432) );
  NANDN U18168 ( .A(n18435), .B(n18436), .Z(n18431) );
  NANDN U18169 ( .A(n18434), .B(n18433), .Z(n18436) );
  ANDN U18170 ( .B(\stack[1][14] ), .A(n5518), .Z(n18273) );
  XNOR U18171 ( .A(n18279), .B(n18437), .Z(n18272) );
  XNOR U18172 ( .A(n18280), .B(n18281), .Z(n18437) );
  AND U18173 ( .A(n18438), .B(n18439), .Z(n18281) );
  NAND U18174 ( .A(n18440), .B(n18441), .Z(n18439) );
  NANDN U18175 ( .A(n18442), .B(n18443), .Z(n18438) );
  OR U18176 ( .A(n18440), .B(n18441), .Z(n18443) );
  ANDN U18177 ( .B(\stack[1][15] ), .A(n5494), .Z(n18280) );
  XNOR U18178 ( .A(n18286), .B(n18444), .Z(n18279) );
  XNOR U18179 ( .A(n18287), .B(n18288), .Z(n18444) );
  AND U18180 ( .A(n18445), .B(n18446), .Z(n18288) );
  NANDN U18181 ( .A(n18447), .B(n18448), .Z(n18446) );
  NANDN U18182 ( .A(n18449), .B(n18450), .Z(n18445) );
  NANDN U18183 ( .A(n18448), .B(n18447), .Z(n18450) );
  ANDN U18184 ( .B(\stack[1][16] ), .A(n5470), .Z(n18287) );
  XNOR U18185 ( .A(n18293), .B(n18451), .Z(n18286) );
  XNOR U18186 ( .A(n18294), .B(n18295), .Z(n18451) );
  AND U18187 ( .A(n18452), .B(n18453), .Z(n18295) );
  NAND U18188 ( .A(n18454), .B(n18455), .Z(n18453) );
  NANDN U18189 ( .A(n18456), .B(n18457), .Z(n18452) );
  OR U18190 ( .A(n18454), .B(n18455), .Z(n18457) );
  ANDN U18191 ( .B(\stack[1][17] ), .A(n5446), .Z(n18294) );
  XNOR U18192 ( .A(n18300), .B(n18458), .Z(n18293) );
  XNOR U18193 ( .A(n18301), .B(n18302), .Z(n18458) );
  AND U18194 ( .A(n18459), .B(n18460), .Z(n18302) );
  NANDN U18195 ( .A(n18461), .B(n18462), .Z(n18460) );
  NANDN U18196 ( .A(n18463), .B(n18464), .Z(n18459) );
  NANDN U18197 ( .A(n18462), .B(n18461), .Z(n18464) );
  ANDN U18198 ( .B(\stack[1][18] ), .A(n5422), .Z(n18301) );
  XNOR U18199 ( .A(n18307), .B(n18465), .Z(n18300) );
  XNOR U18200 ( .A(n18308), .B(n18309), .Z(n18465) );
  AND U18201 ( .A(n18466), .B(n18467), .Z(n18309) );
  NAND U18202 ( .A(n18468), .B(n18469), .Z(n18467) );
  NANDN U18203 ( .A(n18470), .B(n18471), .Z(n18466) );
  OR U18204 ( .A(n18468), .B(n18469), .Z(n18471) );
  ANDN U18205 ( .B(\stack[1][19] ), .A(n5398), .Z(n18308) );
  XNOR U18206 ( .A(n18314), .B(n18472), .Z(n18307) );
  XNOR U18207 ( .A(n18315), .B(n18316), .Z(n18472) );
  AND U18208 ( .A(n18473), .B(n18474), .Z(n18316) );
  NANDN U18209 ( .A(n18475), .B(n18476), .Z(n18474) );
  NANDN U18210 ( .A(n18477), .B(n18478), .Z(n18473) );
  NANDN U18211 ( .A(n18476), .B(n18475), .Z(n18478) );
  ANDN U18212 ( .B(\stack[1][20] ), .A(n5374), .Z(n18315) );
  XNOR U18213 ( .A(n18321), .B(n18479), .Z(n18314) );
  XNOR U18214 ( .A(n18322), .B(n18323), .Z(n18479) );
  AND U18215 ( .A(n18480), .B(n18481), .Z(n18323) );
  NAND U18216 ( .A(n18482), .B(n18483), .Z(n18481) );
  NANDN U18217 ( .A(n18484), .B(n18485), .Z(n18480) );
  OR U18218 ( .A(n18482), .B(n18483), .Z(n18485) );
  ANDN U18219 ( .B(\stack[1][21] ), .A(n5350), .Z(n18322) );
  XNOR U18220 ( .A(n18328), .B(n18486), .Z(n18321) );
  XNOR U18221 ( .A(n18329), .B(n18330), .Z(n18486) );
  AND U18222 ( .A(n18487), .B(n18488), .Z(n18330) );
  NANDN U18223 ( .A(n18489), .B(n18490), .Z(n18488) );
  NANDN U18224 ( .A(n18491), .B(n18492), .Z(n18487) );
  NANDN U18225 ( .A(n18490), .B(n18489), .Z(n18492) );
  ANDN U18226 ( .B(\stack[1][22] ), .A(n5326), .Z(n18329) );
  XNOR U18227 ( .A(n18335), .B(n18493), .Z(n18328) );
  XNOR U18228 ( .A(n18336), .B(n18337), .Z(n18493) );
  AND U18229 ( .A(n18494), .B(n18495), .Z(n18337) );
  NAND U18230 ( .A(n18496), .B(n18497), .Z(n18495) );
  NANDN U18231 ( .A(n18498), .B(n18499), .Z(n18494) );
  OR U18232 ( .A(n18496), .B(n18497), .Z(n18499) );
  ANDN U18233 ( .B(\stack[1][23] ), .A(n5302), .Z(n18336) );
  XNOR U18234 ( .A(n18342), .B(n18500), .Z(n18335) );
  XNOR U18235 ( .A(n18343), .B(n18344), .Z(n18500) );
  AND U18236 ( .A(n18501), .B(n18502), .Z(n18344) );
  NANDN U18237 ( .A(n18503), .B(n18504), .Z(n18502) );
  NANDN U18238 ( .A(n18505), .B(n18506), .Z(n18501) );
  NANDN U18239 ( .A(n18504), .B(n18503), .Z(n18506) );
  ANDN U18240 ( .B(\stack[1][24] ), .A(n5278), .Z(n18343) );
  XNOR U18241 ( .A(n18349), .B(n18507), .Z(n18342) );
  XNOR U18242 ( .A(n18350), .B(n18351), .Z(n18507) );
  AND U18243 ( .A(n18508), .B(n18509), .Z(n18351) );
  NAND U18244 ( .A(n18510), .B(n18511), .Z(n18509) );
  NANDN U18245 ( .A(n18512), .B(n18513), .Z(n18508) );
  OR U18246 ( .A(n18510), .B(n18511), .Z(n18513) );
  ANDN U18247 ( .B(\stack[1][25] ), .A(n5254), .Z(n18350) );
  XNOR U18248 ( .A(n18356), .B(n18514), .Z(n18349) );
  XNOR U18249 ( .A(n18357), .B(n18358), .Z(n18514) );
  AND U18250 ( .A(n18515), .B(n18516), .Z(n18358) );
  NAND U18251 ( .A(n18517), .B(n18518), .Z(n18516) );
  NAND U18252 ( .A(n18519), .B(n18520), .Z(n18515) );
  OR U18253 ( .A(n18517), .B(n18518), .Z(n18519) );
  ANDN U18254 ( .B(\stack[1][26] ), .A(n5230), .Z(n18357) );
  XNOR U18255 ( .A(n18363), .B(n18521), .Z(n18356) );
  XNOR U18256 ( .A(n18364), .B(n18366), .Z(n18521) );
  ANDN U18257 ( .B(n18522), .A(n18523), .Z(n18366) );
  ANDN U18258 ( .B(\stack[0][0] ), .A(n5843), .Z(n18522) );
  ANDN U18259 ( .B(\stack[1][27] ), .A(n5206), .Z(n18364) );
  XOR U18260 ( .A(n18369), .B(n18524), .Z(n18363) );
  NANDN U18261 ( .A(n5160), .B(\stack[1][29] ), .Z(n18524) );
  NANDN U18262 ( .A(n5843), .B(\stack[0][1] ), .Z(n18369) );
  ANDN U18263 ( .B(\stack[1][5] ), .A(n5734), .Z(n9195) );
  AND U18264 ( .A(n18525), .B(n18526), .Z(n9196) );
  NANDN U18265 ( .A(n9200), .B(n9202), .Z(n18526) );
  NANDN U18266 ( .A(n9203), .B(n18527), .Z(n18525) );
  NANDN U18267 ( .A(n9202), .B(n9200), .Z(n18527) );
  XOR U18268 ( .A(n18377), .B(n18528), .Z(n9200) );
  XNOR U18269 ( .A(n18378), .B(n18379), .Z(n18528) );
  AND U18270 ( .A(n18529), .B(n18530), .Z(n18379) );
  NAND U18271 ( .A(n18531), .B(n18532), .Z(n18530) );
  NANDN U18272 ( .A(n18533), .B(n18534), .Z(n18529) );
  OR U18273 ( .A(n18531), .B(n18532), .Z(n18534) );
  ANDN U18274 ( .B(\stack[0][22] ), .A(n5316), .Z(n18378) );
  XNOR U18275 ( .A(n18384), .B(n18535), .Z(n18377) );
  XNOR U18276 ( .A(n18385), .B(n18386), .Z(n18535) );
  AND U18277 ( .A(n18536), .B(n18537), .Z(n18386) );
  NANDN U18278 ( .A(n18538), .B(n18539), .Z(n18537) );
  NANDN U18279 ( .A(n18540), .B(n18541), .Z(n18536) );
  NANDN U18280 ( .A(n18539), .B(n18538), .Z(n18541) );
  ANDN U18281 ( .B(\stack[0][21] ), .A(n5340), .Z(n18385) );
  XNOR U18282 ( .A(n18391), .B(n18542), .Z(n18384) );
  XNOR U18283 ( .A(n18392), .B(n18393), .Z(n18542) );
  AND U18284 ( .A(n18543), .B(n18544), .Z(n18393) );
  NAND U18285 ( .A(n18545), .B(n18546), .Z(n18544) );
  NANDN U18286 ( .A(n18547), .B(n18548), .Z(n18543) );
  OR U18287 ( .A(n18545), .B(n18546), .Z(n18548) );
  ANDN U18288 ( .B(\stack[0][20] ), .A(n5364), .Z(n18392) );
  XNOR U18289 ( .A(n18398), .B(n18549), .Z(n18391) );
  XNOR U18290 ( .A(n18399), .B(n18400), .Z(n18549) );
  AND U18291 ( .A(n18550), .B(n18551), .Z(n18400) );
  NANDN U18292 ( .A(n18552), .B(n18553), .Z(n18551) );
  NANDN U18293 ( .A(n18554), .B(n18555), .Z(n18550) );
  NANDN U18294 ( .A(n18553), .B(n18552), .Z(n18555) );
  ANDN U18295 ( .B(\stack[0][19] ), .A(n5387), .Z(n18399) );
  XNOR U18296 ( .A(n18405), .B(n18556), .Z(n18398) );
  XNOR U18297 ( .A(n18406), .B(n18407), .Z(n18556) );
  AND U18298 ( .A(n18557), .B(n18558), .Z(n18407) );
  NAND U18299 ( .A(n18559), .B(n18560), .Z(n18558) );
  NANDN U18300 ( .A(n18561), .B(n18562), .Z(n18557) );
  OR U18301 ( .A(n18559), .B(n18560), .Z(n18562) );
  ANDN U18302 ( .B(\stack[1][10] ), .A(n5590), .Z(n18406) );
  XNOR U18303 ( .A(n18412), .B(n18563), .Z(n18405) );
  XNOR U18304 ( .A(n18413), .B(n18414), .Z(n18563) );
  AND U18305 ( .A(n18564), .B(n18565), .Z(n18414) );
  NANDN U18306 ( .A(n18566), .B(n18567), .Z(n18565) );
  NANDN U18307 ( .A(n18568), .B(n18569), .Z(n18564) );
  NANDN U18308 ( .A(n18567), .B(n18566), .Z(n18569) );
  ANDN U18309 ( .B(\stack[1][11] ), .A(n5566), .Z(n18413) );
  XNOR U18310 ( .A(n18419), .B(n18570), .Z(n18412) );
  XNOR U18311 ( .A(n18420), .B(n18421), .Z(n18570) );
  AND U18312 ( .A(n18571), .B(n18572), .Z(n18421) );
  NAND U18313 ( .A(n18573), .B(n18574), .Z(n18572) );
  NANDN U18314 ( .A(n18575), .B(n18576), .Z(n18571) );
  OR U18315 ( .A(n18573), .B(n18574), .Z(n18576) );
  ANDN U18316 ( .B(\stack[1][12] ), .A(n5542), .Z(n18420) );
  XNOR U18317 ( .A(n18426), .B(n18577), .Z(n18419) );
  XNOR U18318 ( .A(n18427), .B(n18428), .Z(n18577) );
  AND U18319 ( .A(n18578), .B(n18579), .Z(n18428) );
  NANDN U18320 ( .A(n18580), .B(n18581), .Z(n18579) );
  NANDN U18321 ( .A(n18582), .B(n18583), .Z(n18578) );
  NANDN U18322 ( .A(n18581), .B(n18580), .Z(n18583) );
  ANDN U18323 ( .B(\stack[1][13] ), .A(n5518), .Z(n18427) );
  XNOR U18324 ( .A(n18433), .B(n18584), .Z(n18426) );
  XNOR U18325 ( .A(n18434), .B(n18435), .Z(n18584) );
  AND U18326 ( .A(n18585), .B(n18586), .Z(n18435) );
  NAND U18327 ( .A(n18587), .B(n18588), .Z(n18586) );
  NANDN U18328 ( .A(n18589), .B(n18590), .Z(n18585) );
  OR U18329 ( .A(n18587), .B(n18588), .Z(n18590) );
  ANDN U18330 ( .B(\stack[1][14] ), .A(n5494), .Z(n18434) );
  XNOR U18331 ( .A(n18440), .B(n18591), .Z(n18433) );
  XNOR U18332 ( .A(n18441), .B(n18442), .Z(n18591) );
  AND U18333 ( .A(n18592), .B(n18593), .Z(n18442) );
  NANDN U18334 ( .A(n18594), .B(n18595), .Z(n18593) );
  NANDN U18335 ( .A(n18596), .B(n18597), .Z(n18592) );
  NANDN U18336 ( .A(n18595), .B(n18594), .Z(n18597) );
  ANDN U18337 ( .B(\stack[1][15] ), .A(n5470), .Z(n18441) );
  XNOR U18338 ( .A(n18447), .B(n18598), .Z(n18440) );
  XNOR U18339 ( .A(n18448), .B(n18449), .Z(n18598) );
  AND U18340 ( .A(n18599), .B(n18600), .Z(n18449) );
  NAND U18341 ( .A(n18601), .B(n18602), .Z(n18600) );
  NANDN U18342 ( .A(n18603), .B(n18604), .Z(n18599) );
  OR U18343 ( .A(n18601), .B(n18602), .Z(n18604) );
  ANDN U18344 ( .B(\stack[1][16] ), .A(n5446), .Z(n18448) );
  XNOR U18345 ( .A(n18454), .B(n18605), .Z(n18447) );
  XNOR U18346 ( .A(n18455), .B(n18456), .Z(n18605) );
  AND U18347 ( .A(n18606), .B(n18607), .Z(n18456) );
  NANDN U18348 ( .A(n18608), .B(n18609), .Z(n18607) );
  NANDN U18349 ( .A(n18610), .B(n18611), .Z(n18606) );
  NANDN U18350 ( .A(n18609), .B(n18608), .Z(n18611) );
  ANDN U18351 ( .B(\stack[1][17] ), .A(n5422), .Z(n18455) );
  XNOR U18352 ( .A(n18461), .B(n18612), .Z(n18454) );
  XNOR U18353 ( .A(n18462), .B(n18463), .Z(n18612) );
  AND U18354 ( .A(n18613), .B(n18614), .Z(n18463) );
  NAND U18355 ( .A(n18615), .B(n18616), .Z(n18614) );
  NANDN U18356 ( .A(n18617), .B(n18618), .Z(n18613) );
  OR U18357 ( .A(n18615), .B(n18616), .Z(n18618) );
  ANDN U18358 ( .B(\stack[1][18] ), .A(n5398), .Z(n18462) );
  XNOR U18359 ( .A(n18468), .B(n18619), .Z(n18461) );
  XNOR U18360 ( .A(n18469), .B(n18470), .Z(n18619) );
  AND U18361 ( .A(n18620), .B(n18621), .Z(n18470) );
  NANDN U18362 ( .A(n18622), .B(n18623), .Z(n18621) );
  NANDN U18363 ( .A(n18624), .B(n18625), .Z(n18620) );
  NANDN U18364 ( .A(n18623), .B(n18622), .Z(n18625) );
  ANDN U18365 ( .B(\stack[1][19] ), .A(n5374), .Z(n18469) );
  XNOR U18366 ( .A(n18475), .B(n18626), .Z(n18468) );
  XNOR U18367 ( .A(n18476), .B(n18477), .Z(n18626) );
  AND U18368 ( .A(n18627), .B(n18628), .Z(n18477) );
  NAND U18369 ( .A(n18629), .B(n18630), .Z(n18628) );
  NANDN U18370 ( .A(n18631), .B(n18632), .Z(n18627) );
  OR U18371 ( .A(n18629), .B(n18630), .Z(n18632) );
  ANDN U18372 ( .B(\stack[1][20] ), .A(n5350), .Z(n18476) );
  XNOR U18373 ( .A(n18482), .B(n18633), .Z(n18475) );
  XNOR U18374 ( .A(n18483), .B(n18484), .Z(n18633) );
  AND U18375 ( .A(n18634), .B(n18635), .Z(n18484) );
  NANDN U18376 ( .A(n18636), .B(n18637), .Z(n18635) );
  NANDN U18377 ( .A(n18638), .B(n18639), .Z(n18634) );
  NANDN U18378 ( .A(n18637), .B(n18636), .Z(n18639) );
  ANDN U18379 ( .B(\stack[1][21] ), .A(n5326), .Z(n18483) );
  XNOR U18380 ( .A(n18489), .B(n18640), .Z(n18482) );
  XNOR U18381 ( .A(n18490), .B(n18491), .Z(n18640) );
  AND U18382 ( .A(n18641), .B(n18642), .Z(n18491) );
  NAND U18383 ( .A(n18643), .B(n18644), .Z(n18642) );
  NANDN U18384 ( .A(n18645), .B(n18646), .Z(n18641) );
  OR U18385 ( .A(n18643), .B(n18644), .Z(n18646) );
  ANDN U18386 ( .B(\stack[1][22] ), .A(n5302), .Z(n18490) );
  XNOR U18387 ( .A(n18496), .B(n18647), .Z(n18489) );
  XNOR U18388 ( .A(n18497), .B(n18498), .Z(n18647) );
  AND U18389 ( .A(n18648), .B(n18649), .Z(n18498) );
  NANDN U18390 ( .A(n18650), .B(n18651), .Z(n18649) );
  NANDN U18391 ( .A(n18652), .B(n18653), .Z(n18648) );
  NANDN U18392 ( .A(n18651), .B(n18650), .Z(n18653) );
  ANDN U18393 ( .B(\stack[1][23] ), .A(n5278), .Z(n18497) );
  XNOR U18394 ( .A(n18503), .B(n18654), .Z(n18496) );
  XNOR U18395 ( .A(n18504), .B(n18505), .Z(n18654) );
  AND U18396 ( .A(n18655), .B(n18656), .Z(n18505) );
  NAND U18397 ( .A(n18657), .B(n18658), .Z(n18656) );
  NANDN U18398 ( .A(n18659), .B(n18660), .Z(n18655) );
  OR U18399 ( .A(n18657), .B(n18658), .Z(n18660) );
  ANDN U18400 ( .B(\stack[1][24] ), .A(n5254), .Z(n18504) );
  XNOR U18401 ( .A(n18510), .B(n18661), .Z(n18503) );
  XNOR U18402 ( .A(n18511), .B(n18512), .Z(n18661) );
  AND U18403 ( .A(n18662), .B(n18663), .Z(n18512) );
  NAND U18404 ( .A(n18664), .B(n18665), .Z(n18663) );
  NAND U18405 ( .A(n18666), .B(n18667), .Z(n18662) );
  OR U18406 ( .A(n18664), .B(n18665), .Z(n18666) );
  ANDN U18407 ( .B(\stack[1][25] ), .A(n5230), .Z(n18511) );
  XNOR U18408 ( .A(n18517), .B(n18668), .Z(n18510) );
  XNOR U18409 ( .A(n18518), .B(n18520), .Z(n18668) );
  ANDN U18410 ( .B(n18669), .A(n18670), .Z(n18520) );
  ANDN U18411 ( .B(\stack[0][0] ), .A(n5819), .Z(n18669) );
  ANDN U18412 ( .B(\stack[1][26] ), .A(n5206), .Z(n18518) );
  XOR U18413 ( .A(n18523), .B(n18671), .Z(n18517) );
  NANDN U18414 ( .A(n5160), .B(\stack[1][28] ), .Z(n18671) );
  NANDN U18415 ( .A(n5819), .B(\stack[0][1] ), .Z(n18523) );
  ANDN U18416 ( .B(\stack[0][23] ), .A(n5292), .Z(n9202) );
  AND U18417 ( .A(n18672), .B(n18673), .Z(n9203) );
  NANDN U18418 ( .A(n9210), .B(n18674), .Z(n18672) );
  NANDN U18419 ( .A(n9209), .B(n9207), .Z(n18674) );
  XNOR U18420 ( .A(n18531), .B(n18675), .Z(n9207) );
  XNOR U18421 ( .A(n18532), .B(n18533), .Z(n18675) );
  AND U18422 ( .A(n18676), .B(n18677), .Z(n18533) );
  NANDN U18423 ( .A(n18678), .B(n18679), .Z(n18677) );
  NANDN U18424 ( .A(n18680), .B(n18681), .Z(n18676) );
  NANDN U18425 ( .A(n18679), .B(n18678), .Z(n18681) );
  ANDN U18426 ( .B(\stack[0][21] ), .A(n5316), .Z(n18532) );
  XNOR U18427 ( .A(n18538), .B(n18682), .Z(n18531) );
  XNOR U18428 ( .A(n18539), .B(n18540), .Z(n18682) );
  AND U18429 ( .A(n18683), .B(n18684), .Z(n18540) );
  NAND U18430 ( .A(n18685), .B(n18686), .Z(n18684) );
  NANDN U18431 ( .A(n18687), .B(n18688), .Z(n18683) );
  OR U18432 ( .A(n18685), .B(n18686), .Z(n18688) );
  ANDN U18433 ( .B(\stack[0][20] ), .A(n5340), .Z(n18539) );
  XNOR U18434 ( .A(n18545), .B(n18689), .Z(n18538) );
  XNOR U18435 ( .A(n18546), .B(n18547), .Z(n18689) );
  AND U18436 ( .A(n18690), .B(n18691), .Z(n18547) );
  NANDN U18437 ( .A(n18692), .B(n18693), .Z(n18691) );
  NANDN U18438 ( .A(n18694), .B(n18695), .Z(n18690) );
  NANDN U18439 ( .A(n18693), .B(n18692), .Z(n18695) );
  ANDN U18440 ( .B(\stack[0][19] ), .A(n5364), .Z(n18546) );
  XNOR U18441 ( .A(n18552), .B(n18696), .Z(n18545) );
  XNOR U18442 ( .A(n18553), .B(n18554), .Z(n18696) );
  AND U18443 ( .A(n18697), .B(n18698), .Z(n18554) );
  NAND U18444 ( .A(n18699), .B(n18700), .Z(n18698) );
  NANDN U18445 ( .A(n18701), .B(n18702), .Z(n18697) );
  OR U18446 ( .A(n18699), .B(n18700), .Z(n18702) );
  ANDN U18447 ( .B(\stack[0][18] ), .A(n5387), .Z(n18553) );
  XNOR U18448 ( .A(n18559), .B(n18703), .Z(n18552) );
  XNOR U18449 ( .A(n18560), .B(n18561), .Z(n18703) );
  AND U18450 ( .A(n18704), .B(n18705), .Z(n18561) );
  NANDN U18451 ( .A(n18706), .B(n18707), .Z(n18705) );
  NANDN U18452 ( .A(n18708), .B(n18709), .Z(n18704) );
  NANDN U18453 ( .A(n18707), .B(n18706), .Z(n18709) );
  ANDN U18454 ( .B(\stack[1][10] ), .A(n5566), .Z(n18560) );
  XNOR U18455 ( .A(n18566), .B(n18710), .Z(n18559) );
  XNOR U18456 ( .A(n18567), .B(n18568), .Z(n18710) );
  AND U18457 ( .A(n18711), .B(n18712), .Z(n18568) );
  NAND U18458 ( .A(n18713), .B(n18714), .Z(n18712) );
  NANDN U18459 ( .A(n18715), .B(n18716), .Z(n18711) );
  OR U18460 ( .A(n18713), .B(n18714), .Z(n18716) );
  ANDN U18461 ( .B(\stack[1][11] ), .A(n5542), .Z(n18567) );
  XNOR U18462 ( .A(n18573), .B(n18717), .Z(n18566) );
  XNOR U18463 ( .A(n18574), .B(n18575), .Z(n18717) );
  AND U18464 ( .A(n18718), .B(n18719), .Z(n18575) );
  NANDN U18465 ( .A(n18720), .B(n18721), .Z(n18719) );
  NANDN U18466 ( .A(n18722), .B(n18723), .Z(n18718) );
  NANDN U18467 ( .A(n18721), .B(n18720), .Z(n18723) );
  ANDN U18468 ( .B(\stack[1][12] ), .A(n5518), .Z(n18574) );
  XNOR U18469 ( .A(n18580), .B(n18724), .Z(n18573) );
  XNOR U18470 ( .A(n18581), .B(n18582), .Z(n18724) );
  AND U18471 ( .A(n18725), .B(n18726), .Z(n18582) );
  NAND U18472 ( .A(n18727), .B(n18728), .Z(n18726) );
  NANDN U18473 ( .A(n18729), .B(n18730), .Z(n18725) );
  OR U18474 ( .A(n18727), .B(n18728), .Z(n18730) );
  ANDN U18475 ( .B(\stack[1][13] ), .A(n5494), .Z(n18581) );
  XNOR U18476 ( .A(n18587), .B(n18731), .Z(n18580) );
  XNOR U18477 ( .A(n18588), .B(n18589), .Z(n18731) );
  AND U18478 ( .A(n18732), .B(n18733), .Z(n18589) );
  NANDN U18479 ( .A(n18734), .B(n18735), .Z(n18733) );
  NANDN U18480 ( .A(n18736), .B(n18737), .Z(n18732) );
  NANDN U18481 ( .A(n18735), .B(n18734), .Z(n18737) );
  ANDN U18482 ( .B(\stack[1][14] ), .A(n5470), .Z(n18588) );
  XNOR U18483 ( .A(n18594), .B(n18738), .Z(n18587) );
  XNOR U18484 ( .A(n18595), .B(n18596), .Z(n18738) );
  AND U18485 ( .A(n18739), .B(n18740), .Z(n18596) );
  NAND U18486 ( .A(n18741), .B(n18742), .Z(n18740) );
  NANDN U18487 ( .A(n18743), .B(n18744), .Z(n18739) );
  OR U18488 ( .A(n18741), .B(n18742), .Z(n18744) );
  ANDN U18489 ( .B(\stack[1][15] ), .A(n5446), .Z(n18595) );
  XNOR U18490 ( .A(n18601), .B(n18745), .Z(n18594) );
  XNOR U18491 ( .A(n18602), .B(n18603), .Z(n18745) );
  AND U18492 ( .A(n18746), .B(n18747), .Z(n18603) );
  NANDN U18493 ( .A(n18748), .B(n18749), .Z(n18747) );
  NANDN U18494 ( .A(n18750), .B(n18751), .Z(n18746) );
  NANDN U18495 ( .A(n18749), .B(n18748), .Z(n18751) );
  ANDN U18496 ( .B(\stack[1][16] ), .A(n5422), .Z(n18602) );
  XNOR U18497 ( .A(n18608), .B(n18752), .Z(n18601) );
  XNOR U18498 ( .A(n18609), .B(n18610), .Z(n18752) );
  AND U18499 ( .A(n18753), .B(n18754), .Z(n18610) );
  NAND U18500 ( .A(n18755), .B(n18756), .Z(n18754) );
  NANDN U18501 ( .A(n18757), .B(n18758), .Z(n18753) );
  OR U18502 ( .A(n18755), .B(n18756), .Z(n18758) );
  ANDN U18503 ( .B(\stack[1][17] ), .A(n5398), .Z(n18609) );
  XNOR U18504 ( .A(n18615), .B(n18759), .Z(n18608) );
  XNOR U18505 ( .A(n18616), .B(n18617), .Z(n18759) );
  AND U18506 ( .A(n18760), .B(n18761), .Z(n18617) );
  NANDN U18507 ( .A(n18762), .B(n18763), .Z(n18761) );
  NANDN U18508 ( .A(n18764), .B(n18765), .Z(n18760) );
  NANDN U18509 ( .A(n18763), .B(n18762), .Z(n18765) );
  ANDN U18510 ( .B(\stack[1][18] ), .A(n5374), .Z(n18616) );
  XNOR U18511 ( .A(n18622), .B(n18766), .Z(n18615) );
  XNOR U18512 ( .A(n18623), .B(n18624), .Z(n18766) );
  AND U18513 ( .A(n18767), .B(n18768), .Z(n18624) );
  NAND U18514 ( .A(n18769), .B(n18770), .Z(n18768) );
  NANDN U18515 ( .A(n18771), .B(n18772), .Z(n18767) );
  OR U18516 ( .A(n18769), .B(n18770), .Z(n18772) );
  ANDN U18517 ( .B(\stack[1][19] ), .A(n5350), .Z(n18623) );
  XNOR U18518 ( .A(n18629), .B(n18773), .Z(n18622) );
  XNOR U18519 ( .A(n18630), .B(n18631), .Z(n18773) );
  AND U18520 ( .A(n18774), .B(n18775), .Z(n18631) );
  NANDN U18521 ( .A(n18776), .B(n18777), .Z(n18775) );
  NANDN U18522 ( .A(n18778), .B(n18779), .Z(n18774) );
  NANDN U18523 ( .A(n18777), .B(n18776), .Z(n18779) );
  ANDN U18524 ( .B(\stack[1][20] ), .A(n5326), .Z(n18630) );
  XNOR U18525 ( .A(n18636), .B(n18780), .Z(n18629) );
  XNOR U18526 ( .A(n18637), .B(n18638), .Z(n18780) );
  AND U18527 ( .A(n18781), .B(n18782), .Z(n18638) );
  NAND U18528 ( .A(n18783), .B(n18784), .Z(n18782) );
  NANDN U18529 ( .A(n18785), .B(n18786), .Z(n18781) );
  OR U18530 ( .A(n18783), .B(n18784), .Z(n18786) );
  ANDN U18531 ( .B(\stack[1][21] ), .A(n5302), .Z(n18637) );
  XNOR U18532 ( .A(n18643), .B(n18787), .Z(n18636) );
  XNOR U18533 ( .A(n18644), .B(n18645), .Z(n18787) );
  AND U18534 ( .A(n18788), .B(n18789), .Z(n18645) );
  NANDN U18535 ( .A(n18790), .B(n18791), .Z(n18789) );
  NANDN U18536 ( .A(n18792), .B(n18793), .Z(n18788) );
  NANDN U18537 ( .A(n18791), .B(n18790), .Z(n18793) );
  ANDN U18538 ( .B(\stack[1][22] ), .A(n5278), .Z(n18644) );
  XNOR U18539 ( .A(n18650), .B(n18794), .Z(n18643) );
  XNOR U18540 ( .A(n18651), .B(n18652), .Z(n18794) );
  AND U18541 ( .A(n18795), .B(n18796), .Z(n18652) );
  NAND U18542 ( .A(n18797), .B(n18798), .Z(n18796) );
  NANDN U18543 ( .A(n18799), .B(n18800), .Z(n18795) );
  OR U18544 ( .A(n18797), .B(n18798), .Z(n18800) );
  ANDN U18545 ( .B(\stack[1][23] ), .A(n5254), .Z(n18651) );
  XNOR U18546 ( .A(n18657), .B(n18801), .Z(n18650) );
  XNOR U18547 ( .A(n18658), .B(n18659), .Z(n18801) );
  AND U18548 ( .A(n18802), .B(n18803), .Z(n18659) );
  NAND U18549 ( .A(n18804), .B(n18805), .Z(n18803) );
  NAND U18550 ( .A(n18806), .B(n18807), .Z(n18802) );
  OR U18551 ( .A(n18804), .B(n18805), .Z(n18806) );
  ANDN U18552 ( .B(\stack[1][24] ), .A(n5230), .Z(n18658) );
  XNOR U18553 ( .A(n18664), .B(n18808), .Z(n18657) );
  XNOR U18554 ( .A(n18665), .B(n18667), .Z(n18808) );
  ANDN U18555 ( .B(n18809), .A(n18810), .Z(n18667) );
  ANDN U18556 ( .B(\stack[0][0] ), .A(n5795), .Z(n18809) );
  ANDN U18557 ( .B(\stack[1][25] ), .A(n5206), .Z(n18665) );
  XOR U18558 ( .A(n18670), .B(n18811), .Z(n18664) );
  NANDN U18559 ( .A(n5160), .B(\stack[1][27] ), .Z(n18811) );
  NANDN U18560 ( .A(n5795), .B(\stack[0][1] ), .Z(n18670) );
  ANDN U18561 ( .B(\stack[1][5] ), .A(n5686), .Z(n9209) );
  AND U18562 ( .A(n18812), .B(n18813), .Z(n9210) );
  NANDN U18563 ( .A(n9214), .B(n9216), .Z(n18813) );
  NANDN U18564 ( .A(n9217), .B(n18814), .Z(n18812) );
  NANDN U18565 ( .A(n9216), .B(n9214), .Z(n18814) );
  XOR U18566 ( .A(n18678), .B(n18815), .Z(n9214) );
  XNOR U18567 ( .A(n18679), .B(n18680), .Z(n18815) );
  AND U18568 ( .A(n18816), .B(n18817), .Z(n18680) );
  NAND U18569 ( .A(n18818), .B(n18819), .Z(n18817) );
  NANDN U18570 ( .A(n18820), .B(n18821), .Z(n18816) );
  OR U18571 ( .A(n18818), .B(n18819), .Z(n18821) );
  ANDN U18572 ( .B(\stack[0][20] ), .A(n5316), .Z(n18679) );
  XNOR U18573 ( .A(n18685), .B(n18822), .Z(n18678) );
  XNOR U18574 ( .A(n18686), .B(n18687), .Z(n18822) );
  AND U18575 ( .A(n18823), .B(n18824), .Z(n18687) );
  NANDN U18576 ( .A(n18825), .B(n18826), .Z(n18824) );
  NANDN U18577 ( .A(n18827), .B(n18828), .Z(n18823) );
  NANDN U18578 ( .A(n18826), .B(n18825), .Z(n18828) );
  ANDN U18579 ( .B(\stack[0][19] ), .A(n5340), .Z(n18686) );
  XNOR U18580 ( .A(n18692), .B(n18829), .Z(n18685) );
  XNOR U18581 ( .A(n18693), .B(n18694), .Z(n18829) );
  AND U18582 ( .A(n18830), .B(n18831), .Z(n18694) );
  NAND U18583 ( .A(n18832), .B(n18833), .Z(n18831) );
  NANDN U18584 ( .A(n18834), .B(n18835), .Z(n18830) );
  OR U18585 ( .A(n18832), .B(n18833), .Z(n18835) );
  ANDN U18586 ( .B(\stack[0][18] ), .A(n5364), .Z(n18693) );
  XNOR U18587 ( .A(n18699), .B(n18836), .Z(n18692) );
  XNOR U18588 ( .A(n18700), .B(n18701), .Z(n18836) );
  AND U18589 ( .A(n18837), .B(n18838), .Z(n18701) );
  NANDN U18590 ( .A(n18839), .B(n18840), .Z(n18838) );
  NANDN U18591 ( .A(n18841), .B(n18842), .Z(n18837) );
  NANDN U18592 ( .A(n18840), .B(n18839), .Z(n18842) );
  ANDN U18593 ( .B(\stack[0][17] ), .A(n5387), .Z(n18700) );
  XNOR U18594 ( .A(n18706), .B(n18843), .Z(n18699) );
  XNOR U18595 ( .A(n18707), .B(n18708), .Z(n18843) );
  AND U18596 ( .A(n18844), .B(n18845), .Z(n18708) );
  NAND U18597 ( .A(n18846), .B(n18847), .Z(n18845) );
  NANDN U18598 ( .A(n18848), .B(n18849), .Z(n18844) );
  OR U18599 ( .A(n18846), .B(n18847), .Z(n18849) );
  ANDN U18600 ( .B(\stack[1][10] ), .A(n5542), .Z(n18707) );
  XNOR U18601 ( .A(n18713), .B(n18850), .Z(n18706) );
  XNOR U18602 ( .A(n18714), .B(n18715), .Z(n18850) );
  AND U18603 ( .A(n18851), .B(n18852), .Z(n18715) );
  NANDN U18604 ( .A(n18853), .B(n18854), .Z(n18852) );
  NANDN U18605 ( .A(n18855), .B(n18856), .Z(n18851) );
  NANDN U18606 ( .A(n18854), .B(n18853), .Z(n18856) );
  ANDN U18607 ( .B(\stack[1][11] ), .A(n5518), .Z(n18714) );
  XNOR U18608 ( .A(n18720), .B(n18857), .Z(n18713) );
  XNOR U18609 ( .A(n18721), .B(n18722), .Z(n18857) );
  AND U18610 ( .A(n18858), .B(n18859), .Z(n18722) );
  NAND U18611 ( .A(n18860), .B(n18861), .Z(n18859) );
  NANDN U18612 ( .A(n18862), .B(n18863), .Z(n18858) );
  OR U18613 ( .A(n18860), .B(n18861), .Z(n18863) );
  ANDN U18614 ( .B(\stack[1][12] ), .A(n5494), .Z(n18721) );
  XNOR U18615 ( .A(n18727), .B(n18864), .Z(n18720) );
  XNOR U18616 ( .A(n18728), .B(n18729), .Z(n18864) );
  AND U18617 ( .A(n18865), .B(n18866), .Z(n18729) );
  NANDN U18618 ( .A(n18867), .B(n18868), .Z(n18866) );
  NANDN U18619 ( .A(n18869), .B(n18870), .Z(n18865) );
  NANDN U18620 ( .A(n18868), .B(n18867), .Z(n18870) );
  ANDN U18621 ( .B(\stack[1][13] ), .A(n5470), .Z(n18728) );
  XNOR U18622 ( .A(n18734), .B(n18871), .Z(n18727) );
  XNOR U18623 ( .A(n18735), .B(n18736), .Z(n18871) );
  AND U18624 ( .A(n18872), .B(n18873), .Z(n18736) );
  NAND U18625 ( .A(n18874), .B(n18875), .Z(n18873) );
  NANDN U18626 ( .A(n18876), .B(n18877), .Z(n18872) );
  OR U18627 ( .A(n18874), .B(n18875), .Z(n18877) );
  ANDN U18628 ( .B(\stack[1][14] ), .A(n5446), .Z(n18735) );
  XNOR U18629 ( .A(n18741), .B(n18878), .Z(n18734) );
  XNOR U18630 ( .A(n18742), .B(n18743), .Z(n18878) );
  AND U18631 ( .A(n18879), .B(n18880), .Z(n18743) );
  NANDN U18632 ( .A(n18881), .B(n18882), .Z(n18880) );
  NANDN U18633 ( .A(n18883), .B(n18884), .Z(n18879) );
  NANDN U18634 ( .A(n18882), .B(n18881), .Z(n18884) );
  ANDN U18635 ( .B(\stack[1][15] ), .A(n5422), .Z(n18742) );
  XNOR U18636 ( .A(n18748), .B(n18885), .Z(n18741) );
  XNOR U18637 ( .A(n18749), .B(n18750), .Z(n18885) );
  AND U18638 ( .A(n18886), .B(n18887), .Z(n18750) );
  NAND U18639 ( .A(n18888), .B(n18889), .Z(n18887) );
  NANDN U18640 ( .A(n18890), .B(n18891), .Z(n18886) );
  OR U18641 ( .A(n18888), .B(n18889), .Z(n18891) );
  ANDN U18642 ( .B(\stack[1][16] ), .A(n5398), .Z(n18749) );
  XNOR U18643 ( .A(n18755), .B(n18892), .Z(n18748) );
  XNOR U18644 ( .A(n18756), .B(n18757), .Z(n18892) );
  AND U18645 ( .A(n18893), .B(n18894), .Z(n18757) );
  NANDN U18646 ( .A(n18895), .B(n18896), .Z(n18894) );
  NANDN U18647 ( .A(n18897), .B(n18898), .Z(n18893) );
  NANDN U18648 ( .A(n18896), .B(n18895), .Z(n18898) );
  ANDN U18649 ( .B(\stack[1][17] ), .A(n5374), .Z(n18756) );
  XNOR U18650 ( .A(n18762), .B(n18899), .Z(n18755) );
  XNOR U18651 ( .A(n18763), .B(n18764), .Z(n18899) );
  AND U18652 ( .A(n18900), .B(n18901), .Z(n18764) );
  NAND U18653 ( .A(n18902), .B(n18903), .Z(n18901) );
  NANDN U18654 ( .A(n18904), .B(n18905), .Z(n18900) );
  OR U18655 ( .A(n18902), .B(n18903), .Z(n18905) );
  ANDN U18656 ( .B(\stack[1][18] ), .A(n5350), .Z(n18763) );
  XNOR U18657 ( .A(n18769), .B(n18906), .Z(n18762) );
  XNOR U18658 ( .A(n18770), .B(n18771), .Z(n18906) );
  AND U18659 ( .A(n18907), .B(n18908), .Z(n18771) );
  NANDN U18660 ( .A(n18909), .B(n18910), .Z(n18908) );
  NANDN U18661 ( .A(n18911), .B(n18912), .Z(n18907) );
  NANDN U18662 ( .A(n18910), .B(n18909), .Z(n18912) );
  ANDN U18663 ( .B(\stack[1][19] ), .A(n5326), .Z(n18770) );
  XNOR U18664 ( .A(n18776), .B(n18913), .Z(n18769) );
  XNOR U18665 ( .A(n18777), .B(n18778), .Z(n18913) );
  AND U18666 ( .A(n18914), .B(n18915), .Z(n18778) );
  NAND U18667 ( .A(n18916), .B(n18917), .Z(n18915) );
  NANDN U18668 ( .A(n18918), .B(n18919), .Z(n18914) );
  OR U18669 ( .A(n18916), .B(n18917), .Z(n18919) );
  ANDN U18670 ( .B(\stack[1][20] ), .A(n5302), .Z(n18777) );
  XNOR U18671 ( .A(n18783), .B(n18920), .Z(n18776) );
  XNOR U18672 ( .A(n18784), .B(n18785), .Z(n18920) );
  AND U18673 ( .A(n18921), .B(n18922), .Z(n18785) );
  NANDN U18674 ( .A(n18923), .B(n18924), .Z(n18922) );
  NANDN U18675 ( .A(n18925), .B(n18926), .Z(n18921) );
  NANDN U18676 ( .A(n18924), .B(n18923), .Z(n18926) );
  ANDN U18677 ( .B(\stack[1][21] ), .A(n5278), .Z(n18784) );
  XNOR U18678 ( .A(n18790), .B(n18927), .Z(n18783) );
  XNOR U18679 ( .A(n18791), .B(n18792), .Z(n18927) );
  AND U18680 ( .A(n18928), .B(n18929), .Z(n18792) );
  NAND U18681 ( .A(n18930), .B(n18931), .Z(n18929) );
  NANDN U18682 ( .A(n18932), .B(n18933), .Z(n18928) );
  OR U18683 ( .A(n18930), .B(n18931), .Z(n18933) );
  ANDN U18684 ( .B(\stack[1][22] ), .A(n5254), .Z(n18791) );
  XNOR U18685 ( .A(n18797), .B(n18934), .Z(n18790) );
  XNOR U18686 ( .A(n18798), .B(n18799), .Z(n18934) );
  AND U18687 ( .A(n18935), .B(n18936), .Z(n18799) );
  NAND U18688 ( .A(n18937), .B(n18938), .Z(n18936) );
  NAND U18689 ( .A(n18939), .B(n18940), .Z(n18935) );
  OR U18690 ( .A(n18937), .B(n18938), .Z(n18939) );
  ANDN U18691 ( .B(\stack[1][23] ), .A(n5230), .Z(n18798) );
  XNOR U18692 ( .A(n18804), .B(n18941), .Z(n18797) );
  XNOR U18693 ( .A(n18805), .B(n18807), .Z(n18941) );
  ANDN U18694 ( .B(n18942), .A(n18943), .Z(n18807) );
  ANDN U18695 ( .B(\stack[0][0] ), .A(n5771), .Z(n18942) );
  ANDN U18696 ( .B(\stack[1][24] ), .A(n5206), .Z(n18805) );
  XOR U18697 ( .A(n18810), .B(n18944), .Z(n18804) );
  NANDN U18698 ( .A(n5160), .B(\stack[1][26] ), .Z(n18944) );
  NANDN U18699 ( .A(n5771), .B(\stack[0][1] ), .Z(n18810) );
  ANDN U18700 ( .B(\stack[0][21] ), .A(n5292), .Z(n9216) );
  AND U18701 ( .A(n18945), .B(n18946), .Z(n9217) );
  NANDN U18702 ( .A(n9224), .B(n18947), .Z(n18945) );
  NANDN U18703 ( .A(n9223), .B(n9221), .Z(n18947) );
  XNOR U18704 ( .A(n18818), .B(n18948), .Z(n9221) );
  XNOR U18705 ( .A(n18819), .B(n18820), .Z(n18948) );
  AND U18706 ( .A(n18949), .B(n18950), .Z(n18820) );
  NANDN U18707 ( .A(n18951), .B(n18952), .Z(n18950) );
  NANDN U18708 ( .A(n18953), .B(n18954), .Z(n18949) );
  NANDN U18709 ( .A(n18952), .B(n18951), .Z(n18954) );
  ANDN U18710 ( .B(\stack[0][19] ), .A(n5316), .Z(n18819) );
  XNOR U18711 ( .A(n18825), .B(n18955), .Z(n18818) );
  XNOR U18712 ( .A(n18826), .B(n18827), .Z(n18955) );
  AND U18713 ( .A(n18956), .B(n18957), .Z(n18827) );
  NAND U18714 ( .A(n18958), .B(n18959), .Z(n18957) );
  NANDN U18715 ( .A(n18960), .B(n18961), .Z(n18956) );
  OR U18716 ( .A(n18958), .B(n18959), .Z(n18961) );
  ANDN U18717 ( .B(\stack[0][18] ), .A(n5340), .Z(n18826) );
  XNOR U18718 ( .A(n18832), .B(n18962), .Z(n18825) );
  XNOR U18719 ( .A(n18833), .B(n18834), .Z(n18962) );
  AND U18720 ( .A(n18963), .B(n18964), .Z(n18834) );
  NANDN U18721 ( .A(n18965), .B(n18966), .Z(n18964) );
  NANDN U18722 ( .A(n18967), .B(n18968), .Z(n18963) );
  NANDN U18723 ( .A(n18966), .B(n18965), .Z(n18968) );
  ANDN U18724 ( .B(\stack[0][17] ), .A(n5364), .Z(n18833) );
  XNOR U18725 ( .A(n18839), .B(n18969), .Z(n18832) );
  XNOR U18726 ( .A(n18840), .B(n18841), .Z(n18969) );
  AND U18727 ( .A(n18970), .B(n18971), .Z(n18841) );
  NAND U18728 ( .A(n18972), .B(n18973), .Z(n18971) );
  NANDN U18729 ( .A(n18974), .B(n18975), .Z(n18970) );
  OR U18730 ( .A(n18972), .B(n18973), .Z(n18975) );
  ANDN U18731 ( .B(\stack[0][16] ), .A(n5387), .Z(n18840) );
  XNOR U18732 ( .A(n18846), .B(n18976), .Z(n18839) );
  XNOR U18733 ( .A(n18847), .B(n18848), .Z(n18976) );
  AND U18734 ( .A(n18977), .B(n18978), .Z(n18848) );
  NANDN U18735 ( .A(n18979), .B(n18980), .Z(n18978) );
  NANDN U18736 ( .A(n18981), .B(n18982), .Z(n18977) );
  NANDN U18737 ( .A(n18980), .B(n18979), .Z(n18982) );
  ANDN U18738 ( .B(\stack[1][10] ), .A(n5518), .Z(n18847) );
  XNOR U18739 ( .A(n18853), .B(n18983), .Z(n18846) );
  XNOR U18740 ( .A(n18854), .B(n18855), .Z(n18983) );
  AND U18741 ( .A(n18984), .B(n18985), .Z(n18855) );
  NAND U18742 ( .A(n18986), .B(n18987), .Z(n18985) );
  NANDN U18743 ( .A(n18988), .B(n18989), .Z(n18984) );
  OR U18744 ( .A(n18986), .B(n18987), .Z(n18989) );
  ANDN U18745 ( .B(\stack[1][11] ), .A(n5494), .Z(n18854) );
  XNOR U18746 ( .A(n18860), .B(n18990), .Z(n18853) );
  XNOR U18747 ( .A(n18861), .B(n18862), .Z(n18990) );
  AND U18748 ( .A(n18991), .B(n18992), .Z(n18862) );
  NANDN U18749 ( .A(n18993), .B(n18994), .Z(n18992) );
  NANDN U18750 ( .A(n18995), .B(n18996), .Z(n18991) );
  NANDN U18751 ( .A(n18994), .B(n18993), .Z(n18996) );
  ANDN U18752 ( .B(\stack[1][12] ), .A(n5470), .Z(n18861) );
  XNOR U18753 ( .A(n18867), .B(n18997), .Z(n18860) );
  XNOR U18754 ( .A(n18868), .B(n18869), .Z(n18997) );
  AND U18755 ( .A(n18998), .B(n18999), .Z(n18869) );
  NAND U18756 ( .A(n19000), .B(n19001), .Z(n18999) );
  NANDN U18757 ( .A(n19002), .B(n19003), .Z(n18998) );
  OR U18758 ( .A(n19000), .B(n19001), .Z(n19003) );
  ANDN U18759 ( .B(\stack[1][13] ), .A(n5446), .Z(n18868) );
  XNOR U18760 ( .A(n18874), .B(n19004), .Z(n18867) );
  XNOR U18761 ( .A(n18875), .B(n18876), .Z(n19004) );
  AND U18762 ( .A(n19005), .B(n19006), .Z(n18876) );
  NANDN U18763 ( .A(n19007), .B(n19008), .Z(n19006) );
  NANDN U18764 ( .A(n19009), .B(n19010), .Z(n19005) );
  NANDN U18765 ( .A(n19008), .B(n19007), .Z(n19010) );
  ANDN U18766 ( .B(\stack[1][14] ), .A(n5422), .Z(n18875) );
  XNOR U18767 ( .A(n18881), .B(n19011), .Z(n18874) );
  XNOR U18768 ( .A(n18882), .B(n18883), .Z(n19011) );
  AND U18769 ( .A(n19012), .B(n19013), .Z(n18883) );
  NAND U18770 ( .A(n19014), .B(n19015), .Z(n19013) );
  NANDN U18771 ( .A(n19016), .B(n19017), .Z(n19012) );
  OR U18772 ( .A(n19014), .B(n19015), .Z(n19017) );
  ANDN U18773 ( .B(\stack[1][15] ), .A(n5398), .Z(n18882) );
  XNOR U18774 ( .A(n18888), .B(n19018), .Z(n18881) );
  XNOR U18775 ( .A(n18889), .B(n18890), .Z(n19018) );
  AND U18776 ( .A(n19019), .B(n19020), .Z(n18890) );
  NANDN U18777 ( .A(n19021), .B(n19022), .Z(n19020) );
  NANDN U18778 ( .A(n19023), .B(n19024), .Z(n19019) );
  NANDN U18779 ( .A(n19022), .B(n19021), .Z(n19024) );
  ANDN U18780 ( .B(\stack[1][16] ), .A(n5374), .Z(n18889) );
  XNOR U18781 ( .A(n18895), .B(n19025), .Z(n18888) );
  XNOR U18782 ( .A(n18896), .B(n18897), .Z(n19025) );
  AND U18783 ( .A(n19026), .B(n19027), .Z(n18897) );
  NAND U18784 ( .A(n19028), .B(n19029), .Z(n19027) );
  NANDN U18785 ( .A(n19030), .B(n19031), .Z(n19026) );
  OR U18786 ( .A(n19028), .B(n19029), .Z(n19031) );
  ANDN U18787 ( .B(\stack[1][17] ), .A(n5350), .Z(n18896) );
  XNOR U18788 ( .A(n18902), .B(n19032), .Z(n18895) );
  XNOR U18789 ( .A(n18903), .B(n18904), .Z(n19032) );
  AND U18790 ( .A(n19033), .B(n19034), .Z(n18904) );
  NANDN U18791 ( .A(n19035), .B(n19036), .Z(n19034) );
  NANDN U18792 ( .A(n19037), .B(n19038), .Z(n19033) );
  NANDN U18793 ( .A(n19036), .B(n19035), .Z(n19038) );
  ANDN U18794 ( .B(\stack[1][18] ), .A(n5326), .Z(n18903) );
  XNOR U18795 ( .A(n18909), .B(n19039), .Z(n18902) );
  XNOR U18796 ( .A(n18910), .B(n18911), .Z(n19039) );
  AND U18797 ( .A(n19040), .B(n19041), .Z(n18911) );
  NAND U18798 ( .A(n19042), .B(n19043), .Z(n19041) );
  NANDN U18799 ( .A(n19044), .B(n19045), .Z(n19040) );
  OR U18800 ( .A(n19042), .B(n19043), .Z(n19045) );
  ANDN U18801 ( .B(\stack[1][19] ), .A(n5302), .Z(n18910) );
  XNOR U18802 ( .A(n18916), .B(n19046), .Z(n18909) );
  XNOR U18803 ( .A(n18917), .B(n18918), .Z(n19046) );
  AND U18804 ( .A(n19047), .B(n19048), .Z(n18918) );
  NANDN U18805 ( .A(n19049), .B(n19050), .Z(n19048) );
  NANDN U18806 ( .A(n19051), .B(n19052), .Z(n19047) );
  NANDN U18807 ( .A(n19050), .B(n19049), .Z(n19052) );
  ANDN U18808 ( .B(\stack[1][20] ), .A(n5278), .Z(n18917) );
  XNOR U18809 ( .A(n18923), .B(n19053), .Z(n18916) );
  XNOR U18810 ( .A(n18924), .B(n18925), .Z(n19053) );
  AND U18811 ( .A(n19054), .B(n19055), .Z(n18925) );
  NAND U18812 ( .A(n19056), .B(n19057), .Z(n19055) );
  NANDN U18813 ( .A(n19058), .B(n19059), .Z(n19054) );
  OR U18814 ( .A(n19056), .B(n19057), .Z(n19059) );
  ANDN U18815 ( .B(\stack[1][21] ), .A(n5254), .Z(n18924) );
  XNOR U18816 ( .A(n18930), .B(n19060), .Z(n18923) );
  XNOR U18817 ( .A(n18931), .B(n18932), .Z(n19060) );
  AND U18818 ( .A(n19061), .B(n19062), .Z(n18932) );
  NAND U18819 ( .A(n19063), .B(n19064), .Z(n19062) );
  NAND U18820 ( .A(n19065), .B(n19066), .Z(n19061) );
  OR U18821 ( .A(n19063), .B(n19064), .Z(n19065) );
  ANDN U18822 ( .B(\stack[1][22] ), .A(n5230), .Z(n18931) );
  XNOR U18823 ( .A(n18937), .B(n19067), .Z(n18930) );
  XNOR U18824 ( .A(n18938), .B(n18940), .Z(n19067) );
  ANDN U18825 ( .B(n19068), .A(n19069), .Z(n18940) );
  ANDN U18826 ( .B(\stack[0][0] ), .A(n5747), .Z(n19068) );
  ANDN U18827 ( .B(\stack[1][23] ), .A(n5206), .Z(n18938) );
  XOR U18828 ( .A(n18943), .B(n19070), .Z(n18937) );
  NANDN U18829 ( .A(n5160), .B(\stack[1][25] ), .Z(n19070) );
  NANDN U18830 ( .A(n5747), .B(\stack[0][1] ), .Z(n18943) );
  ANDN U18831 ( .B(\stack[1][5] ), .A(n5638), .Z(n9223) );
  AND U18832 ( .A(n19071), .B(n19072), .Z(n9224) );
  NANDN U18833 ( .A(n9228), .B(n9230), .Z(n19072) );
  NANDN U18834 ( .A(n9231), .B(n19073), .Z(n19071) );
  NANDN U18835 ( .A(n9230), .B(n9228), .Z(n19073) );
  XOR U18836 ( .A(n18951), .B(n19074), .Z(n9228) );
  XNOR U18837 ( .A(n18952), .B(n18953), .Z(n19074) );
  AND U18838 ( .A(n19075), .B(n19076), .Z(n18953) );
  NAND U18839 ( .A(n19077), .B(n19078), .Z(n19076) );
  NANDN U18840 ( .A(n19079), .B(n19080), .Z(n19075) );
  OR U18841 ( .A(n19077), .B(n19078), .Z(n19080) );
  ANDN U18842 ( .B(\stack[0][18] ), .A(n5316), .Z(n18952) );
  XNOR U18843 ( .A(n18958), .B(n19081), .Z(n18951) );
  XNOR U18844 ( .A(n18959), .B(n18960), .Z(n19081) );
  AND U18845 ( .A(n19082), .B(n19083), .Z(n18960) );
  NANDN U18846 ( .A(n19084), .B(n19085), .Z(n19083) );
  NANDN U18847 ( .A(n19086), .B(n19087), .Z(n19082) );
  NANDN U18848 ( .A(n19085), .B(n19084), .Z(n19087) );
  ANDN U18849 ( .B(\stack[0][17] ), .A(n5340), .Z(n18959) );
  XNOR U18850 ( .A(n18965), .B(n19088), .Z(n18958) );
  XNOR U18851 ( .A(n18966), .B(n18967), .Z(n19088) );
  AND U18852 ( .A(n19089), .B(n19090), .Z(n18967) );
  NAND U18853 ( .A(n19091), .B(n19092), .Z(n19090) );
  NANDN U18854 ( .A(n19093), .B(n19094), .Z(n19089) );
  OR U18855 ( .A(n19091), .B(n19092), .Z(n19094) );
  ANDN U18856 ( .B(\stack[0][16] ), .A(n5364), .Z(n18966) );
  XNOR U18857 ( .A(n18972), .B(n19095), .Z(n18965) );
  XNOR U18858 ( .A(n18973), .B(n18974), .Z(n19095) );
  AND U18859 ( .A(n19096), .B(n19097), .Z(n18974) );
  NANDN U18860 ( .A(n19098), .B(n19099), .Z(n19097) );
  NANDN U18861 ( .A(n19100), .B(n19101), .Z(n19096) );
  NANDN U18862 ( .A(n19099), .B(n19098), .Z(n19101) );
  ANDN U18863 ( .B(\stack[0][15] ), .A(n5387), .Z(n18973) );
  XNOR U18864 ( .A(n18979), .B(n19102), .Z(n18972) );
  XNOR U18865 ( .A(n18980), .B(n18981), .Z(n19102) );
  AND U18866 ( .A(n19103), .B(n19104), .Z(n18981) );
  NAND U18867 ( .A(n19105), .B(n19106), .Z(n19104) );
  NANDN U18868 ( .A(n19107), .B(n19108), .Z(n19103) );
  OR U18869 ( .A(n19105), .B(n19106), .Z(n19108) );
  ANDN U18870 ( .B(\stack[1][10] ), .A(n5494), .Z(n18980) );
  XNOR U18871 ( .A(n18986), .B(n19109), .Z(n18979) );
  XNOR U18872 ( .A(n18987), .B(n18988), .Z(n19109) );
  AND U18873 ( .A(n19110), .B(n19111), .Z(n18988) );
  NANDN U18874 ( .A(n19112), .B(n19113), .Z(n19111) );
  NANDN U18875 ( .A(n19114), .B(n19115), .Z(n19110) );
  NANDN U18876 ( .A(n19113), .B(n19112), .Z(n19115) );
  ANDN U18877 ( .B(\stack[1][11] ), .A(n5470), .Z(n18987) );
  XNOR U18878 ( .A(n18993), .B(n19116), .Z(n18986) );
  XNOR U18879 ( .A(n18994), .B(n18995), .Z(n19116) );
  AND U18880 ( .A(n19117), .B(n19118), .Z(n18995) );
  NAND U18881 ( .A(n19119), .B(n19120), .Z(n19118) );
  NANDN U18882 ( .A(n19121), .B(n19122), .Z(n19117) );
  OR U18883 ( .A(n19119), .B(n19120), .Z(n19122) );
  ANDN U18884 ( .B(\stack[1][12] ), .A(n5446), .Z(n18994) );
  XNOR U18885 ( .A(n19000), .B(n19123), .Z(n18993) );
  XNOR U18886 ( .A(n19001), .B(n19002), .Z(n19123) );
  AND U18887 ( .A(n19124), .B(n19125), .Z(n19002) );
  NANDN U18888 ( .A(n19126), .B(n19127), .Z(n19125) );
  NANDN U18889 ( .A(n19128), .B(n19129), .Z(n19124) );
  NANDN U18890 ( .A(n19127), .B(n19126), .Z(n19129) );
  ANDN U18891 ( .B(\stack[1][13] ), .A(n5422), .Z(n19001) );
  XNOR U18892 ( .A(n19007), .B(n19130), .Z(n19000) );
  XNOR U18893 ( .A(n19008), .B(n19009), .Z(n19130) );
  AND U18894 ( .A(n19131), .B(n19132), .Z(n19009) );
  NAND U18895 ( .A(n19133), .B(n19134), .Z(n19132) );
  NANDN U18896 ( .A(n19135), .B(n19136), .Z(n19131) );
  OR U18897 ( .A(n19133), .B(n19134), .Z(n19136) );
  ANDN U18898 ( .B(\stack[1][14] ), .A(n5398), .Z(n19008) );
  XNOR U18899 ( .A(n19014), .B(n19137), .Z(n19007) );
  XNOR U18900 ( .A(n19015), .B(n19016), .Z(n19137) );
  AND U18901 ( .A(n19138), .B(n19139), .Z(n19016) );
  NANDN U18902 ( .A(n19140), .B(n19141), .Z(n19139) );
  NANDN U18903 ( .A(n19142), .B(n19143), .Z(n19138) );
  NANDN U18904 ( .A(n19141), .B(n19140), .Z(n19143) );
  ANDN U18905 ( .B(\stack[1][15] ), .A(n5374), .Z(n19015) );
  XNOR U18906 ( .A(n19021), .B(n19144), .Z(n19014) );
  XNOR U18907 ( .A(n19022), .B(n19023), .Z(n19144) );
  AND U18908 ( .A(n19145), .B(n19146), .Z(n19023) );
  NAND U18909 ( .A(n19147), .B(n19148), .Z(n19146) );
  NANDN U18910 ( .A(n19149), .B(n19150), .Z(n19145) );
  OR U18911 ( .A(n19147), .B(n19148), .Z(n19150) );
  ANDN U18912 ( .B(\stack[1][16] ), .A(n5350), .Z(n19022) );
  XNOR U18913 ( .A(n19028), .B(n19151), .Z(n19021) );
  XNOR U18914 ( .A(n19029), .B(n19030), .Z(n19151) );
  AND U18915 ( .A(n19152), .B(n19153), .Z(n19030) );
  NANDN U18916 ( .A(n19154), .B(n19155), .Z(n19153) );
  NANDN U18917 ( .A(n19156), .B(n19157), .Z(n19152) );
  NANDN U18918 ( .A(n19155), .B(n19154), .Z(n19157) );
  ANDN U18919 ( .B(\stack[1][17] ), .A(n5326), .Z(n19029) );
  XNOR U18920 ( .A(n19035), .B(n19158), .Z(n19028) );
  XNOR U18921 ( .A(n19036), .B(n19037), .Z(n19158) );
  AND U18922 ( .A(n19159), .B(n19160), .Z(n19037) );
  NAND U18923 ( .A(n19161), .B(n19162), .Z(n19160) );
  NANDN U18924 ( .A(n19163), .B(n19164), .Z(n19159) );
  OR U18925 ( .A(n19161), .B(n19162), .Z(n19164) );
  ANDN U18926 ( .B(\stack[1][18] ), .A(n5302), .Z(n19036) );
  XNOR U18927 ( .A(n19042), .B(n19165), .Z(n19035) );
  XNOR U18928 ( .A(n19043), .B(n19044), .Z(n19165) );
  AND U18929 ( .A(n19166), .B(n19167), .Z(n19044) );
  NANDN U18930 ( .A(n19168), .B(n19169), .Z(n19167) );
  NANDN U18931 ( .A(n19170), .B(n19171), .Z(n19166) );
  NANDN U18932 ( .A(n19169), .B(n19168), .Z(n19171) );
  ANDN U18933 ( .B(\stack[1][19] ), .A(n5278), .Z(n19043) );
  XNOR U18934 ( .A(n19049), .B(n19172), .Z(n19042) );
  XNOR U18935 ( .A(n19050), .B(n19051), .Z(n19172) );
  AND U18936 ( .A(n19173), .B(n19174), .Z(n19051) );
  NAND U18937 ( .A(n19175), .B(n19176), .Z(n19174) );
  NANDN U18938 ( .A(n19177), .B(n19178), .Z(n19173) );
  OR U18939 ( .A(n19175), .B(n19176), .Z(n19178) );
  ANDN U18940 ( .B(\stack[1][20] ), .A(n5254), .Z(n19050) );
  XNOR U18941 ( .A(n19056), .B(n19179), .Z(n19049) );
  XNOR U18942 ( .A(n19057), .B(n19058), .Z(n19179) );
  AND U18943 ( .A(n19180), .B(n19181), .Z(n19058) );
  NAND U18944 ( .A(n19182), .B(n19183), .Z(n19181) );
  NAND U18945 ( .A(n19184), .B(n19185), .Z(n19180) );
  OR U18946 ( .A(n19182), .B(n19183), .Z(n19184) );
  ANDN U18947 ( .B(\stack[1][21] ), .A(n5230), .Z(n19057) );
  XNOR U18948 ( .A(n19063), .B(n19186), .Z(n19056) );
  XNOR U18949 ( .A(n19064), .B(n19066), .Z(n19186) );
  ANDN U18950 ( .B(n19187), .A(n19188), .Z(n19066) );
  ANDN U18951 ( .B(\stack[0][0] ), .A(n5723), .Z(n19187) );
  ANDN U18952 ( .B(\stack[1][22] ), .A(n5206), .Z(n19064) );
  XOR U18953 ( .A(n19069), .B(n19189), .Z(n19063) );
  NANDN U18954 ( .A(n5160), .B(\stack[1][24] ), .Z(n19189) );
  NANDN U18955 ( .A(n5723), .B(\stack[0][1] ), .Z(n19069) );
  ANDN U18956 ( .B(\stack[0][19] ), .A(n5292), .Z(n9230) );
  AND U18957 ( .A(n19190), .B(n19191), .Z(n9231) );
  NANDN U18958 ( .A(n9238), .B(n19192), .Z(n19190) );
  NANDN U18959 ( .A(n9237), .B(n9235), .Z(n19192) );
  XNOR U18960 ( .A(n19077), .B(n19193), .Z(n9235) );
  XNOR U18961 ( .A(n19078), .B(n19079), .Z(n19193) );
  AND U18962 ( .A(n19194), .B(n19195), .Z(n19079) );
  NANDN U18963 ( .A(n19196), .B(n19197), .Z(n19195) );
  NANDN U18964 ( .A(n19198), .B(n19199), .Z(n19194) );
  NANDN U18965 ( .A(n19197), .B(n19196), .Z(n19199) );
  ANDN U18966 ( .B(\stack[0][17] ), .A(n5316), .Z(n19078) );
  XNOR U18967 ( .A(n19084), .B(n19200), .Z(n19077) );
  XNOR U18968 ( .A(n19085), .B(n19086), .Z(n19200) );
  AND U18969 ( .A(n19201), .B(n19202), .Z(n19086) );
  NAND U18970 ( .A(n19203), .B(n19204), .Z(n19202) );
  NANDN U18971 ( .A(n19205), .B(n19206), .Z(n19201) );
  OR U18972 ( .A(n19203), .B(n19204), .Z(n19206) );
  ANDN U18973 ( .B(\stack[0][16] ), .A(n5340), .Z(n19085) );
  XNOR U18974 ( .A(n19091), .B(n19207), .Z(n19084) );
  XNOR U18975 ( .A(n19092), .B(n19093), .Z(n19207) );
  AND U18976 ( .A(n19208), .B(n19209), .Z(n19093) );
  NANDN U18977 ( .A(n19210), .B(n19211), .Z(n19209) );
  NANDN U18978 ( .A(n19212), .B(n19213), .Z(n19208) );
  NANDN U18979 ( .A(n19211), .B(n19210), .Z(n19213) );
  ANDN U18980 ( .B(\stack[0][15] ), .A(n5364), .Z(n19092) );
  XNOR U18981 ( .A(n19098), .B(n19214), .Z(n19091) );
  XNOR U18982 ( .A(n19099), .B(n19100), .Z(n19214) );
  AND U18983 ( .A(n19215), .B(n19216), .Z(n19100) );
  NAND U18984 ( .A(n19217), .B(n19218), .Z(n19216) );
  NANDN U18985 ( .A(n19219), .B(n19220), .Z(n19215) );
  OR U18986 ( .A(n19217), .B(n19218), .Z(n19220) );
  ANDN U18987 ( .B(\stack[0][14] ), .A(n5387), .Z(n19099) );
  XNOR U18988 ( .A(n19105), .B(n19221), .Z(n19098) );
  XNOR U18989 ( .A(n19106), .B(n19107), .Z(n19221) );
  AND U18990 ( .A(n19222), .B(n19223), .Z(n19107) );
  NANDN U18991 ( .A(n19224), .B(n19225), .Z(n19223) );
  NANDN U18992 ( .A(n19226), .B(n19227), .Z(n19222) );
  NANDN U18993 ( .A(n19225), .B(n19224), .Z(n19227) );
  ANDN U18994 ( .B(\stack[1][10] ), .A(n5470), .Z(n19106) );
  XNOR U18995 ( .A(n19112), .B(n19228), .Z(n19105) );
  XNOR U18996 ( .A(n19113), .B(n19114), .Z(n19228) );
  AND U18997 ( .A(n19229), .B(n19230), .Z(n19114) );
  NAND U18998 ( .A(n19231), .B(n19232), .Z(n19230) );
  NANDN U18999 ( .A(n19233), .B(n19234), .Z(n19229) );
  OR U19000 ( .A(n19231), .B(n19232), .Z(n19234) );
  ANDN U19001 ( .B(\stack[1][11] ), .A(n5446), .Z(n19113) );
  XNOR U19002 ( .A(n19119), .B(n19235), .Z(n19112) );
  XNOR U19003 ( .A(n19120), .B(n19121), .Z(n19235) );
  AND U19004 ( .A(n19236), .B(n19237), .Z(n19121) );
  NANDN U19005 ( .A(n19238), .B(n19239), .Z(n19237) );
  NANDN U19006 ( .A(n19240), .B(n19241), .Z(n19236) );
  NANDN U19007 ( .A(n19239), .B(n19238), .Z(n19241) );
  ANDN U19008 ( .B(\stack[1][12] ), .A(n5422), .Z(n19120) );
  XNOR U19009 ( .A(n19126), .B(n19242), .Z(n19119) );
  XNOR U19010 ( .A(n19127), .B(n19128), .Z(n19242) );
  AND U19011 ( .A(n19243), .B(n19244), .Z(n19128) );
  NAND U19012 ( .A(n19245), .B(n19246), .Z(n19244) );
  NANDN U19013 ( .A(n19247), .B(n19248), .Z(n19243) );
  OR U19014 ( .A(n19245), .B(n19246), .Z(n19248) );
  ANDN U19015 ( .B(\stack[1][13] ), .A(n5398), .Z(n19127) );
  XNOR U19016 ( .A(n19133), .B(n19249), .Z(n19126) );
  XNOR U19017 ( .A(n19134), .B(n19135), .Z(n19249) );
  AND U19018 ( .A(n19250), .B(n19251), .Z(n19135) );
  NANDN U19019 ( .A(n19252), .B(n19253), .Z(n19251) );
  NANDN U19020 ( .A(n19254), .B(n19255), .Z(n19250) );
  NANDN U19021 ( .A(n19253), .B(n19252), .Z(n19255) );
  ANDN U19022 ( .B(\stack[1][14] ), .A(n5374), .Z(n19134) );
  XNOR U19023 ( .A(n19140), .B(n19256), .Z(n19133) );
  XNOR U19024 ( .A(n19141), .B(n19142), .Z(n19256) );
  AND U19025 ( .A(n19257), .B(n19258), .Z(n19142) );
  NAND U19026 ( .A(n19259), .B(n19260), .Z(n19258) );
  NANDN U19027 ( .A(n19261), .B(n19262), .Z(n19257) );
  OR U19028 ( .A(n19259), .B(n19260), .Z(n19262) );
  ANDN U19029 ( .B(\stack[1][15] ), .A(n5350), .Z(n19141) );
  XNOR U19030 ( .A(n19147), .B(n19263), .Z(n19140) );
  XNOR U19031 ( .A(n19148), .B(n19149), .Z(n19263) );
  AND U19032 ( .A(n19264), .B(n19265), .Z(n19149) );
  NANDN U19033 ( .A(n19266), .B(n19267), .Z(n19265) );
  NANDN U19034 ( .A(n19268), .B(n19269), .Z(n19264) );
  NANDN U19035 ( .A(n19267), .B(n19266), .Z(n19269) );
  ANDN U19036 ( .B(\stack[1][16] ), .A(n5326), .Z(n19148) );
  XNOR U19037 ( .A(n19154), .B(n19270), .Z(n19147) );
  XNOR U19038 ( .A(n19155), .B(n19156), .Z(n19270) );
  AND U19039 ( .A(n19271), .B(n19272), .Z(n19156) );
  NAND U19040 ( .A(n19273), .B(n19274), .Z(n19272) );
  NANDN U19041 ( .A(n19275), .B(n19276), .Z(n19271) );
  OR U19042 ( .A(n19273), .B(n19274), .Z(n19276) );
  ANDN U19043 ( .B(\stack[1][17] ), .A(n5302), .Z(n19155) );
  XNOR U19044 ( .A(n19161), .B(n19277), .Z(n19154) );
  XNOR U19045 ( .A(n19162), .B(n19163), .Z(n19277) );
  AND U19046 ( .A(n19278), .B(n19279), .Z(n19163) );
  NANDN U19047 ( .A(n19280), .B(n19281), .Z(n19279) );
  NANDN U19048 ( .A(n19282), .B(n19283), .Z(n19278) );
  NANDN U19049 ( .A(n19281), .B(n19280), .Z(n19283) );
  ANDN U19050 ( .B(\stack[1][18] ), .A(n5278), .Z(n19162) );
  XNOR U19051 ( .A(n19168), .B(n19284), .Z(n19161) );
  XNOR U19052 ( .A(n19169), .B(n19170), .Z(n19284) );
  AND U19053 ( .A(n19285), .B(n19286), .Z(n19170) );
  NAND U19054 ( .A(n19287), .B(n19288), .Z(n19286) );
  NANDN U19055 ( .A(n19289), .B(n19290), .Z(n19285) );
  OR U19056 ( .A(n19287), .B(n19288), .Z(n19290) );
  ANDN U19057 ( .B(\stack[1][19] ), .A(n5254), .Z(n19169) );
  XNOR U19058 ( .A(n19175), .B(n19291), .Z(n19168) );
  XNOR U19059 ( .A(n19176), .B(n19177), .Z(n19291) );
  AND U19060 ( .A(n19292), .B(n19293), .Z(n19177) );
  NAND U19061 ( .A(n19294), .B(n19295), .Z(n19293) );
  NAND U19062 ( .A(n19296), .B(n19297), .Z(n19292) );
  OR U19063 ( .A(n19294), .B(n19295), .Z(n19296) );
  ANDN U19064 ( .B(\stack[1][20] ), .A(n5230), .Z(n19176) );
  XNOR U19065 ( .A(n19182), .B(n19298), .Z(n19175) );
  XNOR U19066 ( .A(n19183), .B(n19185), .Z(n19298) );
  ANDN U19067 ( .B(n19299), .A(n19300), .Z(n19185) );
  ANDN U19068 ( .B(\stack[0][0] ), .A(n5699), .Z(n19299) );
  ANDN U19069 ( .B(\stack[1][21] ), .A(n5206), .Z(n19183) );
  XOR U19070 ( .A(n19188), .B(n19301), .Z(n19182) );
  NANDN U19071 ( .A(n5160), .B(\stack[1][23] ), .Z(n19301) );
  NANDN U19072 ( .A(n5699), .B(\stack[0][1] ), .Z(n19188) );
  ANDN U19073 ( .B(\stack[1][5] ), .A(n5590), .Z(n9237) );
  AND U19074 ( .A(n19302), .B(n19303), .Z(n9238) );
  NANDN U19075 ( .A(n9242), .B(n9244), .Z(n19303) );
  NANDN U19076 ( .A(n9245), .B(n19304), .Z(n19302) );
  NANDN U19077 ( .A(n9244), .B(n9242), .Z(n19304) );
  XOR U19078 ( .A(n19196), .B(n19305), .Z(n9242) );
  XNOR U19079 ( .A(n19197), .B(n19198), .Z(n19305) );
  AND U19080 ( .A(n19306), .B(n19307), .Z(n19198) );
  NAND U19081 ( .A(n19308), .B(n19309), .Z(n19307) );
  NANDN U19082 ( .A(n19310), .B(n19311), .Z(n19306) );
  OR U19083 ( .A(n19308), .B(n19309), .Z(n19311) );
  ANDN U19084 ( .B(\stack[0][16] ), .A(n5316), .Z(n19197) );
  XNOR U19085 ( .A(n19203), .B(n19312), .Z(n19196) );
  XNOR U19086 ( .A(n19204), .B(n19205), .Z(n19312) );
  AND U19087 ( .A(n19313), .B(n19314), .Z(n19205) );
  NANDN U19088 ( .A(n19315), .B(n19316), .Z(n19314) );
  NANDN U19089 ( .A(n19317), .B(n19318), .Z(n19313) );
  NANDN U19090 ( .A(n19316), .B(n19315), .Z(n19318) );
  ANDN U19091 ( .B(\stack[0][15] ), .A(n5340), .Z(n19204) );
  XNOR U19092 ( .A(n19210), .B(n19319), .Z(n19203) );
  XNOR U19093 ( .A(n19211), .B(n19212), .Z(n19319) );
  AND U19094 ( .A(n19320), .B(n19321), .Z(n19212) );
  NAND U19095 ( .A(n19322), .B(n19323), .Z(n19321) );
  NANDN U19096 ( .A(n19324), .B(n19325), .Z(n19320) );
  OR U19097 ( .A(n19322), .B(n19323), .Z(n19325) );
  ANDN U19098 ( .B(\stack[0][14] ), .A(n5364), .Z(n19211) );
  XNOR U19099 ( .A(n19217), .B(n19326), .Z(n19210) );
  XNOR U19100 ( .A(n19218), .B(n19219), .Z(n19326) );
  AND U19101 ( .A(n19327), .B(n19328), .Z(n19219) );
  NANDN U19102 ( .A(n19329), .B(n19330), .Z(n19328) );
  NANDN U19103 ( .A(n19331), .B(n19332), .Z(n19327) );
  NANDN U19104 ( .A(n19330), .B(n19329), .Z(n19332) );
  ANDN U19105 ( .B(\stack[0][13] ), .A(n5387), .Z(n19218) );
  XNOR U19106 ( .A(n19224), .B(n19333), .Z(n19217) );
  XNOR U19107 ( .A(n19225), .B(n19226), .Z(n19333) );
  AND U19108 ( .A(n19334), .B(n19335), .Z(n19226) );
  NAND U19109 ( .A(n19336), .B(n19337), .Z(n19335) );
  NANDN U19110 ( .A(n19338), .B(n19339), .Z(n19334) );
  OR U19111 ( .A(n19336), .B(n19337), .Z(n19339) );
  ANDN U19112 ( .B(\stack[1][10] ), .A(n5446), .Z(n19225) );
  XNOR U19113 ( .A(n19231), .B(n19340), .Z(n19224) );
  XNOR U19114 ( .A(n19232), .B(n19233), .Z(n19340) );
  AND U19115 ( .A(n19341), .B(n19342), .Z(n19233) );
  NANDN U19116 ( .A(n19343), .B(n19344), .Z(n19342) );
  NANDN U19117 ( .A(n19345), .B(n19346), .Z(n19341) );
  NANDN U19118 ( .A(n19344), .B(n19343), .Z(n19346) );
  ANDN U19119 ( .B(\stack[1][11] ), .A(n5422), .Z(n19232) );
  XNOR U19120 ( .A(n19238), .B(n19347), .Z(n19231) );
  XNOR U19121 ( .A(n19239), .B(n19240), .Z(n19347) );
  AND U19122 ( .A(n19348), .B(n19349), .Z(n19240) );
  NAND U19123 ( .A(n19350), .B(n19351), .Z(n19349) );
  NANDN U19124 ( .A(n19352), .B(n19353), .Z(n19348) );
  OR U19125 ( .A(n19350), .B(n19351), .Z(n19353) );
  ANDN U19126 ( .B(\stack[1][12] ), .A(n5398), .Z(n19239) );
  XNOR U19127 ( .A(n19245), .B(n19354), .Z(n19238) );
  XNOR U19128 ( .A(n19246), .B(n19247), .Z(n19354) );
  AND U19129 ( .A(n19355), .B(n19356), .Z(n19247) );
  NANDN U19130 ( .A(n19357), .B(n19358), .Z(n19356) );
  NANDN U19131 ( .A(n19359), .B(n19360), .Z(n19355) );
  NANDN U19132 ( .A(n19358), .B(n19357), .Z(n19360) );
  ANDN U19133 ( .B(\stack[1][13] ), .A(n5374), .Z(n19246) );
  XNOR U19134 ( .A(n19252), .B(n19361), .Z(n19245) );
  XNOR U19135 ( .A(n19253), .B(n19254), .Z(n19361) );
  AND U19136 ( .A(n19362), .B(n19363), .Z(n19254) );
  NAND U19137 ( .A(n19364), .B(n19365), .Z(n19363) );
  NANDN U19138 ( .A(n19366), .B(n19367), .Z(n19362) );
  OR U19139 ( .A(n19364), .B(n19365), .Z(n19367) );
  ANDN U19140 ( .B(\stack[1][14] ), .A(n5350), .Z(n19253) );
  XNOR U19141 ( .A(n19259), .B(n19368), .Z(n19252) );
  XNOR U19142 ( .A(n19260), .B(n19261), .Z(n19368) );
  AND U19143 ( .A(n19369), .B(n19370), .Z(n19261) );
  NANDN U19144 ( .A(n19371), .B(n19372), .Z(n19370) );
  NANDN U19145 ( .A(n19373), .B(n19374), .Z(n19369) );
  NANDN U19146 ( .A(n19372), .B(n19371), .Z(n19374) );
  ANDN U19147 ( .B(\stack[1][15] ), .A(n5326), .Z(n19260) );
  XNOR U19148 ( .A(n19266), .B(n19375), .Z(n19259) );
  XNOR U19149 ( .A(n19267), .B(n19268), .Z(n19375) );
  AND U19150 ( .A(n19376), .B(n19377), .Z(n19268) );
  NAND U19151 ( .A(n19378), .B(n19379), .Z(n19377) );
  NANDN U19152 ( .A(n19380), .B(n19381), .Z(n19376) );
  OR U19153 ( .A(n19378), .B(n19379), .Z(n19381) );
  ANDN U19154 ( .B(\stack[1][16] ), .A(n5302), .Z(n19267) );
  XNOR U19155 ( .A(n19273), .B(n19382), .Z(n19266) );
  XNOR U19156 ( .A(n19274), .B(n19275), .Z(n19382) );
  AND U19157 ( .A(n19383), .B(n19384), .Z(n19275) );
  NANDN U19158 ( .A(n19385), .B(n19386), .Z(n19384) );
  NANDN U19159 ( .A(n19387), .B(n19388), .Z(n19383) );
  NANDN U19160 ( .A(n19386), .B(n19385), .Z(n19388) );
  ANDN U19161 ( .B(\stack[1][17] ), .A(n5278), .Z(n19274) );
  XNOR U19162 ( .A(n19280), .B(n19389), .Z(n19273) );
  XNOR U19163 ( .A(n19281), .B(n19282), .Z(n19389) );
  AND U19164 ( .A(n19390), .B(n19391), .Z(n19282) );
  NAND U19165 ( .A(n19392), .B(n19393), .Z(n19391) );
  NANDN U19166 ( .A(n19394), .B(n19395), .Z(n19390) );
  OR U19167 ( .A(n19392), .B(n19393), .Z(n19395) );
  ANDN U19168 ( .B(\stack[1][18] ), .A(n5254), .Z(n19281) );
  XNOR U19169 ( .A(n19287), .B(n19396), .Z(n19280) );
  XNOR U19170 ( .A(n19288), .B(n19289), .Z(n19396) );
  AND U19171 ( .A(n19397), .B(n19398), .Z(n19289) );
  NAND U19172 ( .A(n19399), .B(n19400), .Z(n19398) );
  NAND U19173 ( .A(n19401), .B(n19402), .Z(n19397) );
  OR U19174 ( .A(n19399), .B(n19400), .Z(n19401) );
  ANDN U19175 ( .B(\stack[1][19] ), .A(n5230), .Z(n19288) );
  XNOR U19176 ( .A(n19294), .B(n19403), .Z(n19287) );
  XNOR U19177 ( .A(n19295), .B(n19297), .Z(n19403) );
  ANDN U19178 ( .B(n19404), .A(n19405), .Z(n19297) );
  ANDN U19179 ( .B(\stack[0][0] ), .A(n5675), .Z(n19404) );
  ANDN U19180 ( .B(\stack[1][20] ), .A(n5206), .Z(n19295) );
  XOR U19181 ( .A(n19300), .B(n19406), .Z(n19294) );
  NANDN U19182 ( .A(n5160), .B(\stack[1][22] ), .Z(n19406) );
  NANDN U19183 ( .A(n5675), .B(\stack[0][1] ), .Z(n19300) );
  ANDN U19184 ( .B(\stack[0][17] ), .A(n5292), .Z(n9244) );
  AND U19185 ( .A(n19407), .B(n19408), .Z(n9245) );
  NANDN U19186 ( .A(n9252), .B(n19409), .Z(n19407) );
  NANDN U19187 ( .A(n9251), .B(n9249), .Z(n19409) );
  XNOR U19188 ( .A(n19308), .B(n19410), .Z(n9249) );
  XNOR U19189 ( .A(n19309), .B(n19310), .Z(n19410) );
  AND U19190 ( .A(n19411), .B(n19412), .Z(n19310) );
  NANDN U19191 ( .A(n19413), .B(n19414), .Z(n19412) );
  NANDN U19192 ( .A(n19415), .B(n19416), .Z(n19411) );
  NANDN U19193 ( .A(n19414), .B(n19413), .Z(n19416) );
  ANDN U19194 ( .B(\stack[0][15] ), .A(n5316), .Z(n19309) );
  XNOR U19195 ( .A(n19315), .B(n19417), .Z(n19308) );
  XNOR U19196 ( .A(n19316), .B(n19317), .Z(n19417) );
  AND U19197 ( .A(n19418), .B(n19419), .Z(n19317) );
  NAND U19198 ( .A(n19420), .B(n19421), .Z(n19419) );
  NANDN U19199 ( .A(n19422), .B(n19423), .Z(n19418) );
  OR U19200 ( .A(n19420), .B(n19421), .Z(n19423) );
  ANDN U19201 ( .B(\stack[0][14] ), .A(n5340), .Z(n19316) );
  XNOR U19202 ( .A(n19322), .B(n19424), .Z(n19315) );
  XNOR U19203 ( .A(n19323), .B(n19324), .Z(n19424) );
  AND U19204 ( .A(n19425), .B(n19426), .Z(n19324) );
  NANDN U19205 ( .A(n19427), .B(n19428), .Z(n19426) );
  NANDN U19206 ( .A(n19429), .B(n19430), .Z(n19425) );
  NANDN U19207 ( .A(n19428), .B(n19427), .Z(n19430) );
  ANDN U19208 ( .B(\stack[0][13] ), .A(n5364), .Z(n19323) );
  XNOR U19209 ( .A(n19329), .B(n19431), .Z(n19322) );
  XNOR U19210 ( .A(n19330), .B(n19331), .Z(n19431) );
  AND U19211 ( .A(n19432), .B(n19433), .Z(n19331) );
  NAND U19212 ( .A(n19434), .B(n19435), .Z(n19433) );
  NANDN U19213 ( .A(n19436), .B(n19437), .Z(n19432) );
  OR U19214 ( .A(n19434), .B(n19435), .Z(n19437) );
  ANDN U19215 ( .B(\stack[0][12] ), .A(n5387), .Z(n19330) );
  XNOR U19216 ( .A(n19336), .B(n19438), .Z(n19329) );
  XNOR U19217 ( .A(n19337), .B(n19338), .Z(n19438) );
  AND U19218 ( .A(n19439), .B(n19440), .Z(n19338) );
  NANDN U19219 ( .A(n19441), .B(n19442), .Z(n19440) );
  NANDN U19220 ( .A(n19443), .B(n19444), .Z(n19439) );
  NANDN U19221 ( .A(n19442), .B(n19441), .Z(n19444) );
  ANDN U19222 ( .B(\stack[1][10] ), .A(n5422), .Z(n19337) );
  XNOR U19223 ( .A(n19343), .B(n19445), .Z(n19336) );
  XNOR U19224 ( .A(n19344), .B(n19345), .Z(n19445) );
  AND U19225 ( .A(n19446), .B(n19447), .Z(n19345) );
  NAND U19226 ( .A(n19448), .B(n19449), .Z(n19447) );
  NANDN U19227 ( .A(n19450), .B(n19451), .Z(n19446) );
  OR U19228 ( .A(n19448), .B(n19449), .Z(n19451) );
  ANDN U19229 ( .B(\stack[1][11] ), .A(n5398), .Z(n19344) );
  XNOR U19230 ( .A(n19350), .B(n19452), .Z(n19343) );
  XNOR U19231 ( .A(n19351), .B(n19352), .Z(n19452) );
  AND U19232 ( .A(n19453), .B(n19454), .Z(n19352) );
  NANDN U19233 ( .A(n19455), .B(n19456), .Z(n19454) );
  NANDN U19234 ( .A(n19457), .B(n19458), .Z(n19453) );
  NANDN U19235 ( .A(n19456), .B(n19455), .Z(n19458) );
  ANDN U19236 ( .B(\stack[1][12] ), .A(n5374), .Z(n19351) );
  XNOR U19237 ( .A(n19357), .B(n19459), .Z(n19350) );
  XNOR U19238 ( .A(n19358), .B(n19359), .Z(n19459) );
  AND U19239 ( .A(n19460), .B(n19461), .Z(n19359) );
  NAND U19240 ( .A(n19462), .B(n19463), .Z(n19461) );
  NANDN U19241 ( .A(n19464), .B(n19465), .Z(n19460) );
  OR U19242 ( .A(n19462), .B(n19463), .Z(n19465) );
  ANDN U19243 ( .B(\stack[1][13] ), .A(n5350), .Z(n19358) );
  XNOR U19244 ( .A(n19364), .B(n19466), .Z(n19357) );
  XNOR U19245 ( .A(n19365), .B(n19366), .Z(n19466) );
  AND U19246 ( .A(n19467), .B(n19468), .Z(n19366) );
  NANDN U19247 ( .A(n19469), .B(n19470), .Z(n19468) );
  NANDN U19248 ( .A(n19471), .B(n19472), .Z(n19467) );
  NANDN U19249 ( .A(n19470), .B(n19469), .Z(n19472) );
  ANDN U19250 ( .B(\stack[1][14] ), .A(n5326), .Z(n19365) );
  XNOR U19251 ( .A(n19371), .B(n19473), .Z(n19364) );
  XNOR U19252 ( .A(n19372), .B(n19373), .Z(n19473) );
  AND U19253 ( .A(n19474), .B(n19475), .Z(n19373) );
  NAND U19254 ( .A(n19476), .B(n19477), .Z(n19475) );
  NANDN U19255 ( .A(n19478), .B(n19479), .Z(n19474) );
  OR U19256 ( .A(n19476), .B(n19477), .Z(n19479) );
  ANDN U19257 ( .B(\stack[1][15] ), .A(n5302), .Z(n19372) );
  XNOR U19258 ( .A(n19378), .B(n19480), .Z(n19371) );
  XNOR U19259 ( .A(n19379), .B(n19380), .Z(n19480) );
  AND U19260 ( .A(n19481), .B(n19482), .Z(n19380) );
  NANDN U19261 ( .A(n19483), .B(n19484), .Z(n19482) );
  NANDN U19262 ( .A(n19485), .B(n19486), .Z(n19481) );
  NANDN U19263 ( .A(n19484), .B(n19483), .Z(n19486) );
  ANDN U19264 ( .B(\stack[1][16] ), .A(n5278), .Z(n19379) );
  XNOR U19265 ( .A(n19385), .B(n19487), .Z(n19378) );
  XNOR U19266 ( .A(n19386), .B(n19387), .Z(n19487) );
  AND U19267 ( .A(n19488), .B(n19489), .Z(n19387) );
  NAND U19268 ( .A(n19490), .B(n19491), .Z(n19489) );
  NANDN U19269 ( .A(n19492), .B(n19493), .Z(n19488) );
  OR U19270 ( .A(n19490), .B(n19491), .Z(n19493) );
  ANDN U19271 ( .B(\stack[1][17] ), .A(n5254), .Z(n19386) );
  XNOR U19272 ( .A(n19392), .B(n19494), .Z(n19385) );
  XNOR U19273 ( .A(n19393), .B(n19394), .Z(n19494) );
  AND U19274 ( .A(n19495), .B(n19496), .Z(n19394) );
  NAND U19275 ( .A(n19497), .B(n19498), .Z(n19496) );
  NAND U19276 ( .A(n19499), .B(n19500), .Z(n19495) );
  OR U19277 ( .A(n19497), .B(n19498), .Z(n19499) );
  ANDN U19278 ( .B(\stack[1][18] ), .A(n5230), .Z(n19393) );
  XNOR U19279 ( .A(n19399), .B(n19501), .Z(n19392) );
  XNOR U19280 ( .A(n19400), .B(n19402), .Z(n19501) );
  ANDN U19281 ( .B(n19502), .A(n19503), .Z(n19402) );
  ANDN U19282 ( .B(\stack[0][0] ), .A(n5651), .Z(n19502) );
  ANDN U19283 ( .B(\stack[1][19] ), .A(n5206), .Z(n19400) );
  XOR U19284 ( .A(n19405), .B(n19504), .Z(n19399) );
  NANDN U19285 ( .A(n5160), .B(\stack[1][21] ), .Z(n19504) );
  NANDN U19286 ( .A(n5651), .B(\stack[0][1] ), .Z(n19405) );
  ANDN U19287 ( .B(\stack[1][5] ), .A(n5542), .Z(n9251) );
  AND U19288 ( .A(n19505), .B(n19506), .Z(n9252) );
  NANDN U19289 ( .A(n9256), .B(n9258), .Z(n19506) );
  NANDN U19290 ( .A(n9259), .B(n19507), .Z(n19505) );
  NANDN U19291 ( .A(n9258), .B(n9256), .Z(n19507) );
  XOR U19292 ( .A(n19413), .B(n19508), .Z(n9256) );
  XNOR U19293 ( .A(n19414), .B(n19415), .Z(n19508) );
  AND U19294 ( .A(n19509), .B(n19510), .Z(n19415) );
  NAND U19295 ( .A(n19511), .B(n19512), .Z(n19510) );
  NANDN U19296 ( .A(n19513), .B(n19514), .Z(n19509) );
  OR U19297 ( .A(n19511), .B(n19512), .Z(n19514) );
  ANDN U19298 ( .B(\stack[0][14] ), .A(n5316), .Z(n19414) );
  XNOR U19299 ( .A(n19420), .B(n19515), .Z(n19413) );
  XNOR U19300 ( .A(n19421), .B(n19422), .Z(n19515) );
  AND U19301 ( .A(n19516), .B(n19517), .Z(n19422) );
  NANDN U19302 ( .A(n19518), .B(n19519), .Z(n19517) );
  NANDN U19303 ( .A(n19520), .B(n19521), .Z(n19516) );
  NANDN U19304 ( .A(n19519), .B(n19518), .Z(n19521) );
  ANDN U19305 ( .B(\stack[0][13] ), .A(n5340), .Z(n19421) );
  XNOR U19306 ( .A(n19427), .B(n19522), .Z(n19420) );
  XNOR U19307 ( .A(n19428), .B(n19429), .Z(n19522) );
  AND U19308 ( .A(n19523), .B(n19524), .Z(n19429) );
  NAND U19309 ( .A(n19525), .B(n19526), .Z(n19524) );
  NANDN U19310 ( .A(n19527), .B(n19528), .Z(n19523) );
  OR U19311 ( .A(n19525), .B(n19526), .Z(n19528) );
  ANDN U19312 ( .B(\stack[0][12] ), .A(n5364), .Z(n19428) );
  XNOR U19313 ( .A(n19434), .B(n19529), .Z(n19427) );
  XNOR U19314 ( .A(n19435), .B(n19436), .Z(n19529) );
  AND U19315 ( .A(n19530), .B(n19531), .Z(n19436) );
  NANDN U19316 ( .A(n19532), .B(n19533), .Z(n19531) );
  NANDN U19317 ( .A(n19534), .B(n19535), .Z(n19530) );
  NANDN U19318 ( .A(n19533), .B(n19532), .Z(n19535) );
  ANDN U19319 ( .B(\stack[0][11] ), .A(n5387), .Z(n19435) );
  XNOR U19320 ( .A(n19441), .B(n19536), .Z(n19434) );
  XNOR U19321 ( .A(n19442), .B(n19443), .Z(n19536) );
  AND U19322 ( .A(n19537), .B(n19538), .Z(n19443) );
  NAND U19323 ( .A(n19539), .B(n19540), .Z(n19538) );
  NANDN U19324 ( .A(n19541), .B(n19542), .Z(n19537) );
  OR U19325 ( .A(n19539), .B(n19540), .Z(n19542) );
  ANDN U19326 ( .B(\stack[1][10] ), .A(n5398), .Z(n19442) );
  XNOR U19327 ( .A(n19448), .B(n19543), .Z(n19441) );
  XNOR U19328 ( .A(n19449), .B(n19450), .Z(n19543) );
  AND U19329 ( .A(n19544), .B(n19545), .Z(n19450) );
  NANDN U19330 ( .A(n19546), .B(n19547), .Z(n19545) );
  NANDN U19331 ( .A(n19548), .B(n19549), .Z(n19544) );
  NANDN U19332 ( .A(n19547), .B(n19546), .Z(n19549) );
  ANDN U19333 ( .B(\stack[1][11] ), .A(n5374), .Z(n19449) );
  XNOR U19334 ( .A(n19455), .B(n19550), .Z(n19448) );
  XNOR U19335 ( .A(n19456), .B(n19457), .Z(n19550) );
  AND U19336 ( .A(n19551), .B(n19552), .Z(n19457) );
  NAND U19337 ( .A(n19553), .B(n19554), .Z(n19552) );
  NANDN U19338 ( .A(n19555), .B(n19556), .Z(n19551) );
  OR U19339 ( .A(n19553), .B(n19554), .Z(n19556) );
  ANDN U19340 ( .B(\stack[1][12] ), .A(n5350), .Z(n19456) );
  XNOR U19341 ( .A(n19462), .B(n19557), .Z(n19455) );
  XNOR U19342 ( .A(n19463), .B(n19464), .Z(n19557) );
  AND U19343 ( .A(n19558), .B(n19559), .Z(n19464) );
  NANDN U19344 ( .A(n19560), .B(n19561), .Z(n19559) );
  NANDN U19345 ( .A(n19562), .B(n19563), .Z(n19558) );
  NANDN U19346 ( .A(n19561), .B(n19560), .Z(n19563) );
  ANDN U19347 ( .B(\stack[1][13] ), .A(n5326), .Z(n19463) );
  XNOR U19348 ( .A(n19469), .B(n19564), .Z(n19462) );
  XNOR U19349 ( .A(n19470), .B(n19471), .Z(n19564) );
  AND U19350 ( .A(n19565), .B(n19566), .Z(n19471) );
  NAND U19351 ( .A(n19567), .B(n19568), .Z(n19566) );
  NANDN U19352 ( .A(n19569), .B(n19570), .Z(n19565) );
  OR U19353 ( .A(n19567), .B(n19568), .Z(n19570) );
  ANDN U19354 ( .B(\stack[1][14] ), .A(n5302), .Z(n19470) );
  XNOR U19355 ( .A(n19476), .B(n19571), .Z(n19469) );
  XNOR U19356 ( .A(n19477), .B(n19478), .Z(n19571) );
  AND U19357 ( .A(n19572), .B(n19573), .Z(n19478) );
  NANDN U19358 ( .A(n19574), .B(n19575), .Z(n19573) );
  NANDN U19359 ( .A(n19576), .B(n19577), .Z(n19572) );
  NANDN U19360 ( .A(n19575), .B(n19574), .Z(n19577) );
  ANDN U19361 ( .B(\stack[1][15] ), .A(n5278), .Z(n19477) );
  XNOR U19362 ( .A(n19483), .B(n19578), .Z(n19476) );
  XNOR U19363 ( .A(n19484), .B(n19485), .Z(n19578) );
  AND U19364 ( .A(n19579), .B(n19580), .Z(n19485) );
  NAND U19365 ( .A(n19581), .B(n19582), .Z(n19580) );
  NANDN U19366 ( .A(n19583), .B(n19584), .Z(n19579) );
  OR U19367 ( .A(n19581), .B(n19582), .Z(n19584) );
  ANDN U19368 ( .B(\stack[1][16] ), .A(n5254), .Z(n19484) );
  XNOR U19369 ( .A(n19490), .B(n19585), .Z(n19483) );
  XNOR U19370 ( .A(n19491), .B(n19492), .Z(n19585) );
  AND U19371 ( .A(n19586), .B(n19587), .Z(n19492) );
  NAND U19372 ( .A(n19588), .B(n19589), .Z(n19587) );
  NAND U19373 ( .A(n19590), .B(n19591), .Z(n19586) );
  OR U19374 ( .A(n19588), .B(n19589), .Z(n19590) );
  ANDN U19375 ( .B(\stack[1][17] ), .A(n5230), .Z(n19491) );
  XNOR U19376 ( .A(n19497), .B(n19592), .Z(n19490) );
  XNOR U19377 ( .A(n19498), .B(n19500), .Z(n19592) );
  ANDN U19378 ( .B(n19593), .A(n19594), .Z(n19500) );
  ANDN U19379 ( .B(\stack[0][0] ), .A(n5627), .Z(n19593) );
  ANDN U19380 ( .B(\stack[1][18] ), .A(n5206), .Z(n19498) );
  XOR U19381 ( .A(n19503), .B(n19595), .Z(n19497) );
  NANDN U19382 ( .A(n5160), .B(\stack[1][20] ), .Z(n19595) );
  NANDN U19383 ( .A(n5627), .B(\stack[0][1] ), .Z(n19503) );
  ANDN U19384 ( .B(\stack[0][15] ), .A(n5292), .Z(n9258) );
  AND U19385 ( .A(n19596), .B(n19597), .Z(n9259) );
  NANDN U19386 ( .A(n9266), .B(n19598), .Z(n19596) );
  NANDN U19387 ( .A(n9265), .B(n9263), .Z(n19598) );
  XNOR U19388 ( .A(n19511), .B(n19599), .Z(n9263) );
  XNOR U19389 ( .A(n19512), .B(n19513), .Z(n19599) );
  AND U19390 ( .A(n19600), .B(n19601), .Z(n19513) );
  NANDN U19391 ( .A(n19602), .B(n19603), .Z(n19601) );
  NANDN U19392 ( .A(n19604), .B(n19605), .Z(n19600) );
  NANDN U19393 ( .A(n19603), .B(n19602), .Z(n19605) );
  ANDN U19394 ( .B(\stack[0][13] ), .A(n5316), .Z(n19512) );
  XNOR U19395 ( .A(n19518), .B(n19606), .Z(n19511) );
  XNOR U19396 ( .A(n19519), .B(n19520), .Z(n19606) );
  AND U19397 ( .A(n19607), .B(n19608), .Z(n19520) );
  NAND U19398 ( .A(n19609), .B(n19610), .Z(n19608) );
  NANDN U19399 ( .A(n19611), .B(n19612), .Z(n19607) );
  OR U19400 ( .A(n19609), .B(n19610), .Z(n19612) );
  ANDN U19401 ( .B(\stack[0][12] ), .A(n5340), .Z(n19519) );
  XNOR U19402 ( .A(n19525), .B(n19613), .Z(n19518) );
  XNOR U19403 ( .A(n19526), .B(n19527), .Z(n19613) );
  AND U19404 ( .A(n19614), .B(n19615), .Z(n19527) );
  NANDN U19405 ( .A(n19616), .B(n19617), .Z(n19615) );
  NANDN U19406 ( .A(n19618), .B(n19619), .Z(n19614) );
  NANDN U19407 ( .A(n19617), .B(n19616), .Z(n19619) );
  ANDN U19408 ( .B(\stack[0][11] ), .A(n5364), .Z(n19526) );
  XNOR U19409 ( .A(n19532), .B(n19620), .Z(n19525) );
  XNOR U19410 ( .A(n19533), .B(n19534), .Z(n19620) );
  AND U19411 ( .A(n19621), .B(n19622), .Z(n19534) );
  NAND U19412 ( .A(n19623), .B(n19624), .Z(n19622) );
  NANDN U19413 ( .A(n19625), .B(n19626), .Z(n19621) );
  OR U19414 ( .A(n19623), .B(n19624), .Z(n19626) );
  ANDN U19415 ( .B(\stack[0][10] ), .A(n5387), .Z(n19533) );
  XNOR U19416 ( .A(n19539), .B(n19627), .Z(n19532) );
  XNOR U19417 ( .A(n19540), .B(n19541), .Z(n19627) );
  AND U19418 ( .A(n19628), .B(n19629), .Z(n19541) );
  NANDN U19419 ( .A(n19630), .B(n19631), .Z(n19629) );
  NANDN U19420 ( .A(n19632), .B(n19633), .Z(n19628) );
  NANDN U19421 ( .A(n19631), .B(n19630), .Z(n19633) );
  ANDN U19422 ( .B(\stack[1][10] ), .A(n5374), .Z(n19540) );
  XNOR U19423 ( .A(n19546), .B(n19634), .Z(n19539) );
  XNOR U19424 ( .A(n19547), .B(n19548), .Z(n19634) );
  AND U19425 ( .A(n19635), .B(n19636), .Z(n19548) );
  NAND U19426 ( .A(n19637), .B(n19638), .Z(n19636) );
  NANDN U19427 ( .A(n19639), .B(n19640), .Z(n19635) );
  OR U19428 ( .A(n19637), .B(n19638), .Z(n19640) );
  ANDN U19429 ( .B(\stack[1][11] ), .A(n5350), .Z(n19547) );
  XNOR U19430 ( .A(n19553), .B(n19641), .Z(n19546) );
  XNOR U19431 ( .A(n19554), .B(n19555), .Z(n19641) );
  AND U19432 ( .A(n19642), .B(n19643), .Z(n19555) );
  NANDN U19433 ( .A(n19644), .B(n19645), .Z(n19643) );
  NANDN U19434 ( .A(n19646), .B(n19647), .Z(n19642) );
  NANDN U19435 ( .A(n19645), .B(n19644), .Z(n19647) );
  ANDN U19436 ( .B(\stack[1][12] ), .A(n5326), .Z(n19554) );
  XNOR U19437 ( .A(n19560), .B(n19648), .Z(n19553) );
  XNOR U19438 ( .A(n19561), .B(n19562), .Z(n19648) );
  AND U19439 ( .A(n19649), .B(n19650), .Z(n19562) );
  NAND U19440 ( .A(n19651), .B(n19652), .Z(n19650) );
  NANDN U19441 ( .A(n19653), .B(n19654), .Z(n19649) );
  OR U19442 ( .A(n19651), .B(n19652), .Z(n19654) );
  ANDN U19443 ( .B(\stack[1][13] ), .A(n5302), .Z(n19561) );
  XNOR U19444 ( .A(n19567), .B(n19655), .Z(n19560) );
  XNOR U19445 ( .A(n19568), .B(n19569), .Z(n19655) );
  AND U19446 ( .A(n19656), .B(n19657), .Z(n19569) );
  NANDN U19447 ( .A(n19658), .B(n19659), .Z(n19657) );
  NANDN U19448 ( .A(n19660), .B(n19661), .Z(n19656) );
  NANDN U19449 ( .A(n19659), .B(n19658), .Z(n19661) );
  ANDN U19450 ( .B(\stack[1][14] ), .A(n5278), .Z(n19568) );
  XNOR U19451 ( .A(n19574), .B(n19662), .Z(n19567) );
  XNOR U19452 ( .A(n19575), .B(n19576), .Z(n19662) );
  AND U19453 ( .A(n19663), .B(n19664), .Z(n19576) );
  NAND U19454 ( .A(n19665), .B(n19666), .Z(n19664) );
  NANDN U19455 ( .A(n19667), .B(n19668), .Z(n19663) );
  OR U19456 ( .A(n19665), .B(n19666), .Z(n19668) );
  ANDN U19457 ( .B(\stack[1][15] ), .A(n5254), .Z(n19575) );
  XNOR U19458 ( .A(n19581), .B(n19669), .Z(n19574) );
  XNOR U19459 ( .A(n19582), .B(n19583), .Z(n19669) );
  AND U19460 ( .A(n19670), .B(n19671), .Z(n19583) );
  NAND U19461 ( .A(n19672), .B(n19673), .Z(n19671) );
  NAND U19462 ( .A(n19674), .B(n19675), .Z(n19670) );
  OR U19463 ( .A(n19672), .B(n19673), .Z(n19674) );
  ANDN U19464 ( .B(\stack[1][16] ), .A(n5230), .Z(n19582) );
  XNOR U19465 ( .A(n19588), .B(n19676), .Z(n19581) );
  XNOR U19466 ( .A(n19589), .B(n19591), .Z(n19676) );
  ANDN U19467 ( .B(n19677), .A(n19678), .Z(n19591) );
  ANDN U19468 ( .B(\stack[0][0] ), .A(n5603), .Z(n19677) );
  ANDN U19469 ( .B(\stack[1][17] ), .A(n5206), .Z(n19589) );
  XOR U19470 ( .A(n19594), .B(n19679), .Z(n19588) );
  NANDN U19471 ( .A(n5160), .B(\stack[1][19] ), .Z(n19679) );
  NANDN U19472 ( .A(n5603), .B(\stack[0][1] ), .Z(n19594) );
  ANDN U19473 ( .B(\stack[1][5] ), .A(n5494), .Z(n9265) );
  AND U19474 ( .A(n19680), .B(n19681), .Z(n9266) );
  NANDN U19475 ( .A(n9270), .B(n9272), .Z(n19681) );
  NANDN U19476 ( .A(n9273), .B(n19682), .Z(n19680) );
  NANDN U19477 ( .A(n9272), .B(n9270), .Z(n19682) );
  XOR U19478 ( .A(n19602), .B(n19683), .Z(n9270) );
  XNOR U19479 ( .A(n19603), .B(n19604), .Z(n19683) );
  AND U19480 ( .A(n19684), .B(n19685), .Z(n19604) );
  NAND U19481 ( .A(n19686), .B(n19687), .Z(n19685) );
  NANDN U19482 ( .A(n19688), .B(n19689), .Z(n19684) );
  OR U19483 ( .A(n19686), .B(n19687), .Z(n19689) );
  ANDN U19484 ( .B(\stack[0][12] ), .A(n5316), .Z(n19603) );
  XNOR U19485 ( .A(n19609), .B(n19690), .Z(n19602) );
  XNOR U19486 ( .A(n19610), .B(n19611), .Z(n19690) );
  AND U19487 ( .A(n19691), .B(n19692), .Z(n19611) );
  NANDN U19488 ( .A(n19693), .B(n19694), .Z(n19692) );
  NANDN U19489 ( .A(n19695), .B(n19696), .Z(n19691) );
  NANDN U19490 ( .A(n19694), .B(n19693), .Z(n19696) );
  ANDN U19491 ( .B(\stack[0][11] ), .A(n5340), .Z(n19610) );
  XNOR U19492 ( .A(n19616), .B(n19697), .Z(n19609) );
  XNOR U19493 ( .A(n19617), .B(n19618), .Z(n19697) );
  AND U19494 ( .A(n19698), .B(n19699), .Z(n19618) );
  NAND U19495 ( .A(n19700), .B(n19701), .Z(n19699) );
  NANDN U19496 ( .A(n19702), .B(n19703), .Z(n19698) );
  OR U19497 ( .A(n19700), .B(n19701), .Z(n19703) );
  ANDN U19498 ( .B(\stack[0][10] ), .A(n5364), .Z(n19617) );
  XNOR U19499 ( .A(n19623), .B(n19704), .Z(n19616) );
  XNOR U19500 ( .A(n19624), .B(n19625), .Z(n19704) );
  AND U19501 ( .A(n19705), .B(n19706), .Z(n19625) );
  NANDN U19502 ( .A(n19707), .B(n19708), .Z(n19706) );
  NANDN U19503 ( .A(n19709), .B(n19710), .Z(n19705) );
  NANDN U19504 ( .A(n19708), .B(n19707), .Z(n19710) );
  ANDN U19505 ( .B(\stack[1][9] ), .A(n5374), .Z(n19624) );
  XNOR U19506 ( .A(n19630), .B(n19711), .Z(n19623) );
  XNOR U19507 ( .A(n19631), .B(n19632), .Z(n19711) );
  AND U19508 ( .A(n19712), .B(n19713), .Z(n19632) );
  NAND U19509 ( .A(n19714), .B(n19715), .Z(n19713) );
  NANDN U19510 ( .A(n19716), .B(n19717), .Z(n19712) );
  OR U19511 ( .A(n19714), .B(n19715), .Z(n19717) );
  ANDN U19512 ( .B(\stack[1][10] ), .A(n5350), .Z(n19631) );
  XNOR U19513 ( .A(n19637), .B(n19718), .Z(n19630) );
  XNOR U19514 ( .A(n19638), .B(n19639), .Z(n19718) );
  AND U19515 ( .A(n19719), .B(n19720), .Z(n19639) );
  NANDN U19516 ( .A(n19721), .B(n19722), .Z(n19720) );
  NANDN U19517 ( .A(n19723), .B(n19724), .Z(n19719) );
  NANDN U19518 ( .A(n19722), .B(n19721), .Z(n19724) );
  ANDN U19519 ( .B(\stack[1][11] ), .A(n5326), .Z(n19638) );
  XNOR U19520 ( .A(n19644), .B(n19725), .Z(n19637) );
  XNOR U19521 ( .A(n19645), .B(n19646), .Z(n19725) );
  AND U19522 ( .A(n19726), .B(n19727), .Z(n19646) );
  NAND U19523 ( .A(n19728), .B(n19729), .Z(n19727) );
  NANDN U19524 ( .A(n19730), .B(n19731), .Z(n19726) );
  OR U19525 ( .A(n19728), .B(n19729), .Z(n19731) );
  ANDN U19526 ( .B(\stack[1][12] ), .A(n5302), .Z(n19645) );
  XNOR U19527 ( .A(n19651), .B(n19732), .Z(n19644) );
  XNOR U19528 ( .A(n19652), .B(n19653), .Z(n19732) );
  AND U19529 ( .A(n19733), .B(n19734), .Z(n19653) );
  NANDN U19530 ( .A(n19735), .B(n19736), .Z(n19734) );
  NANDN U19531 ( .A(n19737), .B(n19738), .Z(n19733) );
  NANDN U19532 ( .A(n19736), .B(n19735), .Z(n19738) );
  ANDN U19533 ( .B(\stack[1][13] ), .A(n5278), .Z(n19652) );
  XNOR U19534 ( .A(n19658), .B(n19739), .Z(n19651) );
  XNOR U19535 ( .A(n19659), .B(n19660), .Z(n19739) );
  AND U19536 ( .A(n19740), .B(n19741), .Z(n19660) );
  NAND U19537 ( .A(n19742), .B(n19743), .Z(n19741) );
  NANDN U19538 ( .A(n19744), .B(n19745), .Z(n19740) );
  OR U19539 ( .A(n19742), .B(n19743), .Z(n19745) );
  ANDN U19540 ( .B(\stack[1][14] ), .A(n5254), .Z(n19659) );
  XNOR U19541 ( .A(n19665), .B(n19746), .Z(n19658) );
  XNOR U19542 ( .A(n19666), .B(n19667), .Z(n19746) );
  AND U19543 ( .A(n19747), .B(n19748), .Z(n19667) );
  NAND U19544 ( .A(n19749), .B(n19750), .Z(n19748) );
  NAND U19545 ( .A(n19751), .B(n19752), .Z(n19747) );
  OR U19546 ( .A(n19749), .B(n19750), .Z(n19751) );
  ANDN U19547 ( .B(\stack[1][15] ), .A(n5230), .Z(n19666) );
  XNOR U19548 ( .A(n19672), .B(n19753), .Z(n19665) );
  XNOR U19549 ( .A(n19673), .B(n19675), .Z(n19753) );
  ANDN U19550 ( .B(n19754), .A(n19755), .Z(n19675) );
  ANDN U19551 ( .B(\stack[0][0] ), .A(n5579), .Z(n19754) );
  ANDN U19552 ( .B(\stack[1][16] ), .A(n5206), .Z(n19673) );
  XOR U19553 ( .A(n19678), .B(n19756), .Z(n19672) );
  NANDN U19554 ( .A(n5160), .B(\stack[1][18] ), .Z(n19756) );
  NANDN U19555 ( .A(n5579), .B(\stack[0][1] ), .Z(n19678) );
  ANDN U19556 ( .B(\stack[0][13] ), .A(n5292), .Z(n9272) );
  AND U19557 ( .A(n19757), .B(n19758), .Z(n9273) );
  NANDN U19558 ( .A(n9280), .B(n19759), .Z(n19757) );
  NANDN U19559 ( .A(n9279), .B(n9277), .Z(n19759) );
  XNOR U19560 ( .A(n19686), .B(n19760), .Z(n9277) );
  XNOR U19561 ( .A(n19687), .B(n19688), .Z(n19760) );
  AND U19562 ( .A(n19761), .B(n19762), .Z(n19688) );
  NANDN U19563 ( .A(n19763), .B(n19764), .Z(n19762) );
  NANDN U19564 ( .A(n19765), .B(n19766), .Z(n19761) );
  NANDN U19565 ( .A(n19764), .B(n19763), .Z(n19766) );
  ANDN U19566 ( .B(\stack[0][11] ), .A(n5316), .Z(n19687) );
  XNOR U19567 ( .A(n19693), .B(n19767), .Z(n19686) );
  XNOR U19568 ( .A(n19694), .B(n19695), .Z(n19767) );
  AND U19569 ( .A(n19768), .B(n19769), .Z(n19695) );
  NAND U19570 ( .A(n19770), .B(n19771), .Z(n19769) );
  NANDN U19571 ( .A(n19772), .B(n19773), .Z(n19768) );
  OR U19572 ( .A(n19770), .B(n19771), .Z(n19773) );
  ANDN U19573 ( .B(\stack[0][10] ), .A(n5340), .Z(n19694) );
  XNOR U19574 ( .A(n19700), .B(n19774), .Z(n19693) );
  XNOR U19575 ( .A(n19701), .B(n19702), .Z(n19774) );
  AND U19576 ( .A(n19775), .B(n19776), .Z(n19702) );
  NANDN U19577 ( .A(n19777), .B(n19778), .Z(n19776) );
  NANDN U19578 ( .A(n19779), .B(n19780), .Z(n19775) );
  NANDN U19579 ( .A(n19778), .B(n19777), .Z(n19780) );
  ANDN U19580 ( .B(\stack[1][8] ), .A(n5374), .Z(n19701) );
  XNOR U19581 ( .A(n19707), .B(n19781), .Z(n19700) );
  XNOR U19582 ( .A(n19708), .B(n19709), .Z(n19781) );
  AND U19583 ( .A(n19782), .B(n19783), .Z(n19709) );
  NAND U19584 ( .A(n19784), .B(n19785), .Z(n19783) );
  NANDN U19585 ( .A(n19786), .B(n19787), .Z(n19782) );
  OR U19586 ( .A(n19784), .B(n19785), .Z(n19787) );
  ANDN U19587 ( .B(\stack[0][8] ), .A(n5387), .Z(n19708) );
  XNOR U19588 ( .A(n19714), .B(n19788), .Z(n19707) );
  XNOR U19589 ( .A(n19715), .B(n19716), .Z(n19788) );
  AND U19590 ( .A(n19789), .B(n19790), .Z(n19716) );
  NANDN U19591 ( .A(n19791), .B(n19792), .Z(n19790) );
  NANDN U19592 ( .A(n19793), .B(n19794), .Z(n19789) );
  NANDN U19593 ( .A(n19792), .B(n19791), .Z(n19794) );
  ANDN U19594 ( .B(\stack[1][10] ), .A(n5326), .Z(n19715) );
  XNOR U19595 ( .A(n19721), .B(n19795), .Z(n19714) );
  XNOR U19596 ( .A(n19722), .B(n19723), .Z(n19795) );
  AND U19597 ( .A(n19796), .B(n19797), .Z(n19723) );
  NAND U19598 ( .A(n19798), .B(n19799), .Z(n19797) );
  NANDN U19599 ( .A(n19800), .B(n19801), .Z(n19796) );
  OR U19600 ( .A(n19798), .B(n19799), .Z(n19801) );
  ANDN U19601 ( .B(\stack[1][11] ), .A(n5302), .Z(n19722) );
  XNOR U19602 ( .A(n19728), .B(n19802), .Z(n19721) );
  XNOR U19603 ( .A(n19729), .B(n19730), .Z(n19802) );
  AND U19604 ( .A(n19803), .B(n19804), .Z(n19730) );
  NANDN U19605 ( .A(n19805), .B(n19806), .Z(n19804) );
  NANDN U19606 ( .A(n19807), .B(n19808), .Z(n19803) );
  NANDN U19607 ( .A(n19806), .B(n19805), .Z(n19808) );
  ANDN U19608 ( .B(\stack[1][12] ), .A(n5278), .Z(n19729) );
  XNOR U19609 ( .A(n19735), .B(n19809), .Z(n19728) );
  XNOR U19610 ( .A(n19736), .B(n19737), .Z(n19809) );
  AND U19611 ( .A(n19810), .B(n19811), .Z(n19737) );
  NAND U19612 ( .A(n19812), .B(n19813), .Z(n19811) );
  NANDN U19613 ( .A(n19814), .B(n19815), .Z(n19810) );
  OR U19614 ( .A(n19812), .B(n19813), .Z(n19815) );
  ANDN U19615 ( .B(\stack[1][13] ), .A(n5254), .Z(n19736) );
  XNOR U19616 ( .A(n19742), .B(n19816), .Z(n19735) );
  XNOR U19617 ( .A(n19743), .B(n19744), .Z(n19816) );
  AND U19618 ( .A(n19817), .B(n19818), .Z(n19744) );
  NAND U19619 ( .A(n19819), .B(n19820), .Z(n19818) );
  NAND U19620 ( .A(n19821), .B(n19822), .Z(n19817) );
  OR U19621 ( .A(n19819), .B(n19820), .Z(n19821) );
  ANDN U19622 ( .B(\stack[1][14] ), .A(n5230), .Z(n19743) );
  XNOR U19623 ( .A(n19749), .B(n19823), .Z(n19742) );
  XNOR U19624 ( .A(n19750), .B(n19752), .Z(n19823) );
  ANDN U19625 ( .B(n19824), .A(n19825), .Z(n19752) );
  ANDN U19626 ( .B(\stack[0][0] ), .A(n5555), .Z(n19824) );
  ANDN U19627 ( .B(\stack[1][15] ), .A(n5206), .Z(n19750) );
  XOR U19628 ( .A(n19755), .B(n19826), .Z(n19749) );
  NANDN U19629 ( .A(n5160), .B(\stack[1][17] ), .Z(n19826) );
  NANDN U19630 ( .A(n5555), .B(\stack[0][1] ), .Z(n19755) );
  ANDN U19631 ( .B(\stack[1][5] ), .A(n5446), .Z(n9279) );
  AND U19632 ( .A(n19827), .B(n19828), .Z(n9280) );
  NANDN U19633 ( .A(n9284), .B(n9286), .Z(n19828) );
  NANDN U19634 ( .A(n9287), .B(n19829), .Z(n19827) );
  NANDN U19635 ( .A(n9286), .B(n9284), .Z(n19829) );
  XOR U19636 ( .A(n19763), .B(n19830), .Z(n9284) );
  XNOR U19637 ( .A(n19764), .B(n19765), .Z(n19830) );
  AND U19638 ( .A(n19831), .B(n19832), .Z(n19765) );
  NAND U19639 ( .A(n19833), .B(n19834), .Z(n19832) );
  NANDN U19640 ( .A(n19835), .B(n19836), .Z(n19831) );
  OR U19641 ( .A(n19833), .B(n19834), .Z(n19836) );
  ANDN U19642 ( .B(\stack[0][10] ), .A(n5316), .Z(n19764) );
  XNOR U19643 ( .A(n19770), .B(n19837), .Z(n19763) );
  XNOR U19644 ( .A(n19771), .B(n19772), .Z(n19837) );
  AND U19645 ( .A(n19838), .B(n19839), .Z(n19772) );
  NANDN U19646 ( .A(n19840), .B(n19841), .Z(n19839) );
  NANDN U19647 ( .A(n19842), .B(n19843), .Z(n19838) );
  NANDN U19648 ( .A(n19841), .B(n19840), .Z(n19843) );
  ANDN U19649 ( .B(\stack[1][7] ), .A(n5374), .Z(n19771) );
  XNOR U19650 ( .A(n19777), .B(n19844), .Z(n19770) );
  XNOR U19651 ( .A(n19778), .B(n19779), .Z(n19844) );
  AND U19652 ( .A(n19845), .B(n19846), .Z(n19779) );
  NAND U19653 ( .A(n19847), .B(n19848), .Z(n19846) );
  NANDN U19654 ( .A(n19849), .B(n19850), .Z(n19845) );
  OR U19655 ( .A(n19847), .B(n19848), .Z(n19850) );
  ANDN U19656 ( .B(\stack[0][8] ), .A(n5364), .Z(n19778) );
  XNOR U19657 ( .A(n19784), .B(n19851), .Z(n19777) );
  XNOR U19658 ( .A(n19785), .B(n19786), .Z(n19851) );
  AND U19659 ( .A(n19852), .B(n19853), .Z(n19786) );
  NANDN U19660 ( .A(n19854), .B(n19855), .Z(n19853) );
  NANDN U19661 ( .A(n19856), .B(n19857), .Z(n19852) );
  NANDN U19662 ( .A(n19855), .B(n19854), .Z(n19857) );
  ANDN U19663 ( .B(\stack[0][7] ), .A(n5387), .Z(n19785) );
  XNOR U19664 ( .A(n19791), .B(n19858), .Z(n19784) );
  XNOR U19665 ( .A(n19792), .B(n19793), .Z(n19858) );
  AND U19666 ( .A(n19859), .B(n19860), .Z(n19793) );
  NAND U19667 ( .A(n19861), .B(n19862), .Z(n19860) );
  NANDN U19668 ( .A(n19863), .B(n19864), .Z(n19859) );
  OR U19669 ( .A(n19861), .B(n19862), .Z(n19864) );
  ANDN U19670 ( .B(\stack[1][10] ), .A(n5302), .Z(n19792) );
  XNOR U19671 ( .A(n19798), .B(n19865), .Z(n19791) );
  XNOR U19672 ( .A(n19799), .B(n19800), .Z(n19865) );
  AND U19673 ( .A(n19866), .B(n19867), .Z(n19800) );
  NANDN U19674 ( .A(n19868), .B(n19869), .Z(n19867) );
  NANDN U19675 ( .A(n19870), .B(n19871), .Z(n19866) );
  NANDN U19676 ( .A(n19869), .B(n19868), .Z(n19871) );
  ANDN U19677 ( .B(\stack[1][11] ), .A(n5278), .Z(n19799) );
  XNOR U19678 ( .A(n19805), .B(n19872), .Z(n19798) );
  XNOR U19679 ( .A(n19806), .B(n19807), .Z(n19872) );
  AND U19680 ( .A(n19873), .B(n19874), .Z(n19807) );
  NAND U19681 ( .A(n19875), .B(n19876), .Z(n19874) );
  NANDN U19682 ( .A(n19877), .B(n19878), .Z(n19873) );
  OR U19683 ( .A(n19875), .B(n19876), .Z(n19878) );
  ANDN U19684 ( .B(\stack[1][12] ), .A(n5254), .Z(n19806) );
  XNOR U19685 ( .A(n19812), .B(n19879), .Z(n19805) );
  XNOR U19686 ( .A(n19813), .B(n19814), .Z(n19879) );
  AND U19687 ( .A(n19880), .B(n19881), .Z(n19814) );
  NAND U19688 ( .A(n19882), .B(n19883), .Z(n19881) );
  NAND U19689 ( .A(n19884), .B(n19885), .Z(n19880) );
  OR U19690 ( .A(n19882), .B(n19883), .Z(n19884) );
  ANDN U19691 ( .B(\stack[1][13] ), .A(n5230), .Z(n19813) );
  XNOR U19692 ( .A(n19819), .B(n19886), .Z(n19812) );
  XNOR U19693 ( .A(n19820), .B(n19822), .Z(n19886) );
  ANDN U19694 ( .B(n19887), .A(n19888), .Z(n19822) );
  ANDN U19695 ( .B(\stack[0][0] ), .A(n5531), .Z(n19887) );
  ANDN U19696 ( .B(\stack[1][14] ), .A(n5206), .Z(n19820) );
  XOR U19697 ( .A(n19825), .B(n19889), .Z(n19819) );
  NANDN U19698 ( .A(n5160), .B(\stack[1][16] ), .Z(n19889) );
  NANDN U19699 ( .A(n5531), .B(\stack[0][1] ), .Z(n19825) );
  ANDN U19700 ( .B(\stack[0][11] ), .A(n5292), .Z(n9286) );
  AND U19701 ( .A(n19890), .B(n19891), .Z(n9287) );
  NANDN U19702 ( .A(n9294), .B(n19892), .Z(n19890) );
  NANDN U19703 ( .A(n9293), .B(n9291), .Z(n19892) );
  XNOR U19704 ( .A(n19833), .B(n19893), .Z(n9291) );
  XNOR U19705 ( .A(n19834), .B(n19835), .Z(n19893) );
  AND U19706 ( .A(n19894), .B(n19895), .Z(n19835) );
  NANDN U19707 ( .A(n19896), .B(n19897), .Z(n19895) );
  NANDN U19708 ( .A(n19898), .B(n19899), .Z(n19894) );
  NANDN U19709 ( .A(n19897), .B(n19896), .Z(n19899) );
  ANDN U19710 ( .B(\stack[1][6] ), .A(n5374), .Z(n19834) );
  XNOR U19711 ( .A(n19840), .B(n19900), .Z(n19833) );
  XNOR U19712 ( .A(n19841), .B(n19842), .Z(n19900) );
  AND U19713 ( .A(n19901), .B(n19902), .Z(n19842) );
  NAND U19714 ( .A(n19903), .B(n19904), .Z(n19902) );
  NANDN U19715 ( .A(n19905), .B(n19906), .Z(n19901) );
  OR U19716 ( .A(n19903), .B(n19904), .Z(n19906) );
  ANDN U19717 ( .B(\stack[0][8] ), .A(n5340), .Z(n19841) );
  XNOR U19718 ( .A(n19847), .B(n19907), .Z(n19840) );
  XNOR U19719 ( .A(n19848), .B(n19849), .Z(n19907) );
  AND U19720 ( .A(n19908), .B(n19909), .Z(n19849) );
  NANDN U19721 ( .A(n19910), .B(n19911), .Z(n19909) );
  NANDN U19722 ( .A(n19912), .B(n19913), .Z(n19908) );
  NANDN U19723 ( .A(n19911), .B(n19910), .Z(n19913) );
  ANDN U19724 ( .B(\stack[0][7] ), .A(n5364), .Z(n19848) );
  XNOR U19725 ( .A(n19854), .B(n19914), .Z(n19847) );
  XNOR U19726 ( .A(n19855), .B(n19856), .Z(n19914) );
  AND U19727 ( .A(n19915), .B(n19916), .Z(n19856) );
  NAND U19728 ( .A(n19917), .B(n19918), .Z(n19916) );
  NANDN U19729 ( .A(n19919), .B(n19920), .Z(n19915) );
  OR U19730 ( .A(n19917), .B(n19918), .Z(n19920) );
  ANDN U19731 ( .B(\stack[0][6] ), .A(n5387), .Z(n19855) );
  XNOR U19732 ( .A(n19861), .B(n19921), .Z(n19854) );
  XNOR U19733 ( .A(n19862), .B(n19863), .Z(n19921) );
  AND U19734 ( .A(n19922), .B(n19923), .Z(n19863) );
  NANDN U19735 ( .A(n19924), .B(n19925), .Z(n19923) );
  NANDN U19736 ( .A(n19926), .B(n19927), .Z(n19922) );
  NANDN U19737 ( .A(n19925), .B(n19924), .Z(n19927) );
  ANDN U19738 ( .B(\stack[1][10] ), .A(n5278), .Z(n19862) );
  XNOR U19739 ( .A(n19868), .B(n19928), .Z(n19861) );
  XNOR U19740 ( .A(n19869), .B(n19870), .Z(n19928) );
  AND U19741 ( .A(n19929), .B(n19930), .Z(n19870) );
  NAND U19742 ( .A(n19931), .B(n19932), .Z(n19930) );
  NANDN U19743 ( .A(n19933), .B(n19934), .Z(n19929) );
  OR U19744 ( .A(n19931), .B(n19932), .Z(n19934) );
  ANDN U19745 ( .B(\stack[1][11] ), .A(n5254), .Z(n19869) );
  XNOR U19746 ( .A(n19875), .B(n19935), .Z(n19868) );
  XNOR U19747 ( .A(n19876), .B(n19877), .Z(n19935) );
  AND U19748 ( .A(n19936), .B(n19937), .Z(n19877) );
  NAND U19749 ( .A(n19938), .B(n19939), .Z(n19937) );
  NAND U19750 ( .A(n19940), .B(n19941), .Z(n19936) );
  OR U19751 ( .A(n19938), .B(n19939), .Z(n19940) );
  ANDN U19752 ( .B(\stack[1][12] ), .A(n5230), .Z(n19876) );
  XNOR U19753 ( .A(n19882), .B(n19942), .Z(n19875) );
  XNOR U19754 ( .A(n19883), .B(n19885), .Z(n19942) );
  ANDN U19755 ( .B(n19943), .A(n19944), .Z(n19885) );
  ANDN U19756 ( .B(\stack[0][0] ), .A(n5507), .Z(n19943) );
  ANDN U19757 ( .B(\stack[1][13] ), .A(n5206), .Z(n19883) );
  XOR U19758 ( .A(n19888), .B(n19945), .Z(n19882) );
  NANDN U19759 ( .A(n5160), .B(\stack[1][15] ), .Z(n19945) );
  NANDN U19760 ( .A(n5507), .B(\stack[0][1] ), .Z(n19888) );
  ANDN U19761 ( .B(\stack[1][5] ), .A(n5398), .Z(n9293) );
  AND U19762 ( .A(n19946), .B(n19947), .Z(n9294) );
  NANDN U19763 ( .A(n9298), .B(n9300), .Z(n19947) );
  NANDN U19764 ( .A(n9301), .B(n19948), .Z(n19946) );
  NANDN U19765 ( .A(n9300), .B(n9298), .Z(n19948) );
  XOR U19766 ( .A(n19896), .B(n19949), .Z(n9298) );
  XNOR U19767 ( .A(n19897), .B(n19898), .Z(n19949) );
  AND U19768 ( .A(n19950), .B(n19951), .Z(n19898) );
  NAND U19769 ( .A(n19952), .B(n19953), .Z(n19951) );
  NANDN U19770 ( .A(n19954), .B(n19955), .Z(n19950) );
  OR U19771 ( .A(n19952), .B(n19953), .Z(n19955) );
  ANDN U19772 ( .B(\stack[0][8] ), .A(n5316), .Z(n19897) );
  XNOR U19773 ( .A(n19903), .B(n19956), .Z(n19896) );
  XNOR U19774 ( .A(n19904), .B(n19905), .Z(n19956) );
  AND U19775 ( .A(n19957), .B(n19958), .Z(n19905) );
  NANDN U19776 ( .A(n19959), .B(n19960), .Z(n19958) );
  NANDN U19777 ( .A(n19961), .B(n19962), .Z(n19957) );
  NANDN U19778 ( .A(n19960), .B(n19959), .Z(n19962) );
  ANDN U19779 ( .B(\stack[0][7] ), .A(n5340), .Z(n19904) );
  XNOR U19780 ( .A(n19910), .B(n19963), .Z(n19903) );
  XNOR U19781 ( .A(n19911), .B(n19912), .Z(n19963) );
  AND U19782 ( .A(n19964), .B(n19965), .Z(n19912) );
  NAND U19783 ( .A(n19966), .B(n19967), .Z(n19965) );
  NANDN U19784 ( .A(n19968), .B(n19969), .Z(n19964) );
  OR U19785 ( .A(n19966), .B(n19967), .Z(n19969) );
  ANDN U19786 ( .B(\stack[0][6] ), .A(n5364), .Z(n19911) );
  XNOR U19787 ( .A(n19917), .B(n19970), .Z(n19910) );
  XNOR U19788 ( .A(n19918), .B(n19919), .Z(n19970) );
  AND U19789 ( .A(n19971), .B(n19972), .Z(n19919) );
  NANDN U19790 ( .A(n19973), .B(n19974), .Z(n19972) );
  NANDN U19791 ( .A(n19975), .B(n19976), .Z(n19971) );
  NANDN U19792 ( .A(n19974), .B(n19973), .Z(n19976) );
  ANDN U19793 ( .B(\stack[0][5] ), .A(n5387), .Z(n19918) );
  XNOR U19794 ( .A(n19924), .B(n19977), .Z(n19917) );
  XNOR U19795 ( .A(n19925), .B(n19926), .Z(n19977) );
  AND U19796 ( .A(n19978), .B(n19979), .Z(n19926) );
  NAND U19797 ( .A(n19980), .B(n19981), .Z(n19979) );
  NANDN U19798 ( .A(n19982), .B(n19983), .Z(n19978) );
  OR U19799 ( .A(n19980), .B(n19981), .Z(n19983) );
  ANDN U19800 ( .B(\stack[1][10] ), .A(n5254), .Z(n19925) );
  XNOR U19801 ( .A(n19931), .B(n19984), .Z(n19924) );
  XNOR U19802 ( .A(n19932), .B(n19933), .Z(n19984) );
  AND U19803 ( .A(n19985), .B(n19986), .Z(n19933) );
  NAND U19804 ( .A(n19987), .B(n19988), .Z(n19986) );
  NAND U19805 ( .A(n19989), .B(n19990), .Z(n19985) );
  OR U19806 ( .A(n19987), .B(n19988), .Z(n19989) );
  ANDN U19807 ( .B(\stack[1][11] ), .A(n5230), .Z(n19932) );
  XNOR U19808 ( .A(n19938), .B(n19991), .Z(n19931) );
  XNOR U19809 ( .A(n19939), .B(n19941), .Z(n19991) );
  ANDN U19810 ( .B(n19992), .A(n19993), .Z(n19941) );
  ANDN U19811 ( .B(\stack[0][0] ), .A(n5483), .Z(n19992) );
  ANDN U19812 ( .B(\stack[1][12] ), .A(n5206), .Z(n19939) );
  XOR U19813 ( .A(n19944), .B(n19994), .Z(n19938) );
  NANDN U19814 ( .A(n5160), .B(\stack[1][14] ), .Z(n19994) );
  NANDN U19815 ( .A(n5483), .B(\stack[0][1] ), .Z(n19944) );
  ANDN U19816 ( .B(\stack[1][5] ), .A(n5374), .Z(n9300) );
  AND U19817 ( .A(n19995), .B(n19996), .Z(n9301) );
  NANDN U19818 ( .A(n9308), .B(n19997), .Z(n19995) );
  NANDN U19819 ( .A(n9307), .B(n9305), .Z(n19997) );
  XNOR U19820 ( .A(n19952), .B(n19998), .Z(n9305) );
  XNOR U19821 ( .A(n19953), .B(n19954), .Z(n19998) );
  AND U19822 ( .A(n19999), .B(n20000), .Z(n19954) );
  NANDN U19823 ( .A(n20001), .B(n20002), .Z(n20000) );
  NANDN U19824 ( .A(n20003), .B(n20004), .Z(n19999) );
  NANDN U19825 ( .A(n20002), .B(n20001), .Z(n20004) );
  ANDN U19826 ( .B(\stack[0][7] ), .A(n5316), .Z(n19953) );
  XNOR U19827 ( .A(n19959), .B(n20005), .Z(n19952) );
  XNOR U19828 ( .A(n19960), .B(n19961), .Z(n20005) );
  AND U19829 ( .A(n20006), .B(n20007), .Z(n19961) );
  NAND U19830 ( .A(n20008), .B(n20009), .Z(n20007) );
  NANDN U19831 ( .A(n20010), .B(n20011), .Z(n20006) );
  OR U19832 ( .A(n20008), .B(n20009), .Z(n20011) );
  ANDN U19833 ( .B(\stack[0][6] ), .A(n5340), .Z(n19960) );
  XNOR U19834 ( .A(n19966), .B(n20012), .Z(n19959) );
  XNOR U19835 ( .A(n19967), .B(n19968), .Z(n20012) );
  AND U19836 ( .A(n20013), .B(n20014), .Z(n19968) );
  NANDN U19837 ( .A(n20015), .B(n20016), .Z(n20014) );
  NANDN U19838 ( .A(n20017), .B(n20018), .Z(n20013) );
  NANDN U19839 ( .A(n20016), .B(n20015), .Z(n20018) );
  ANDN U19840 ( .B(\stack[0][5] ), .A(n5364), .Z(n19967) );
  XNOR U19841 ( .A(n19973), .B(n20019), .Z(n19966) );
  XNOR U19842 ( .A(n19974), .B(n19975), .Z(n20019) );
  AND U19843 ( .A(n20020), .B(n20021), .Z(n19975) );
  NAND U19844 ( .A(n20022), .B(n20023), .Z(n20021) );
  NANDN U19845 ( .A(n20024), .B(n20025), .Z(n20020) );
  OR U19846 ( .A(n20022), .B(n20023), .Z(n20025) );
  ANDN U19847 ( .B(\stack[0][4] ), .A(n5387), .Z(n19974) );
  XNOR U19848 ( .A(n19980), .B(n20026), .Z(n19973) );
  XNOR U19849 ( .A(n19981), .B(n19982), .Z(n20026) );
  AND U19850 ( .A(n20027), .B(n20028), .Z(n19982) );
  NAND U19851 ( .A(n20029), .B(n20030), .Z(n20028) );
  NAND U19852 ( .A(n20031), .B(n20032), .Z(n20027) );
  OR U19853 ( .A(n20029), .B(n20030), .Z(n20031) );
  ANDN U19854 ( .B(\stack[1][10] ), .A(n5230), .Z(n19981) );
  XNOR U19855 ( .A(n19987), .B(n20033), .Z(n19980) );
  XNOR U19856 ( .A(n19988), .B(n19990), .Z(n20033) );
  ANDN U19857 ( .B(n20034), .A(n20035), .Z(n19990) );
  ANDN U19858 ( .B(\stack[0][0] ), .A(n5459), .Z(n20034) );
  ANDN U19859 ( .B(\stack[1][11] ), .A(n5206), .Z(n19988) );
  XOR U19860 ( .A(n19993), .B(n20036), .Z(n19987) );
  NANDN U19861 ( .A(n5160), .B(\stack[1][13] ), .Z(n20036) );
  NANDN U19862 ( .A(n5459), .B(\stack[0][1] ), .Z(n19993) );
  ANDN U19863 ( .B(\stack[1][5] ), .A(n5350), .Z(n9307) );
  AND U19864 ( .A(n20037), .B(n20038), .Z(n9308) );
  NANDN U19865 ( .A(n9312), .B(n9314), .Z(n20038) );
  NANDN U19866 ( .A(n9315), .B(n20039), .Z(n20037) );
  NANDN U19867 ( .A(n9314), .B(n9312), .Z(n20039) );
  XOR U19868 ( .A(n20001), .B(n20040), .Z(n9312) );
  XNOR U19869 ( .A(n20002), .B(n20003), .Z(n20040) );
  AND U19870 ( .A(n20041), .B(n20042), .Z(n20003) );
  NAND U19871 ( .A(n20043), .B(n20044), .Z(n20042) );
  NANDN U19872 ( .A(n20045), .B(n20046), .Z(n20041) );
  OR U19873 ( .A(n20043), .B(n20044), .Z(n20046) );
  ANDN U19874 ( .B(\stack[0][6] ), .A(n5316), .Z(n20002) );
  XNOR U19875 ( .A(n20008), .B(n20047), .Z(n20001) );
  XNOR U19876 ( .A(n20009), .B(n20010), .Z(n20047) );
  AND U19877 ( .A(n20048), .B(n20049), .Z(n20010) );
  NANDN U19878 ( .A(n20050), .B(n20051), .Z(n20049) );
  NANDN U19879 ( .A(n20052), .B(n20053), .Z(n20048) );
  NANDN U19880 ( .A(n20051), .B(n20050), .Z(n20053) );
  ANDN U19881 ( .B(\stack[0][5] ), .A(n5340), .Z(n20009) );
  XNOR U19882 ( .A(n20015), .B(n20054), .Z(n20008) );
  XNOR U19883 ( .A(n20016), .B(n20017), .Z(n20054) );
  AND U19884 ( .A(n20055), .B(n20056), .Z(n20017) );
  NAND U19885 ( .A(n20057), .B(n20058), .Z(n20056) );
  NANDN U19886 ( .A(n20059), .B(n20060), .Z(n20055) );
  OR U19887 ( .A(n20057), .B(n20058), .Z(n20060) );
  ANDN U19888 ( .B(\stack[0][4] ), .A(n5364), .Z(n20016) );
  XNOR U19889 ( .A(n20022), .B(n20061), .Z(n20015) );
  XNOR U19890 ( .A(n20023), .B(n20024), .Z(n20061) );
  AND U19891 ( .A(n20062), .B(n20063), .Z(n20024) );
  NAND U19892 ( .A(n20064), .B(n20065), .Z(n20063) );
  NAND U19893 ( .A(n20066), .B(n20067), .Z(n20062) );
  OR U19894 ( .A(n20064), .B(n20065), .Z(n20066) );
  ANDN U19895 ( .B(\stack[0][3] ), .A(n5387), .Z(n20023) );
  XNOR U19896 ( .A(n20029), .B(n20068), .Z(n20022) );
  XNOR U19897 ( .A(n20030), .B(n20032), .Z(n20068) );
  ANDN U19898 ( .B(n20069), .A(n20070), .Z(n20032) );
  ANDN U19899 ( .B(\stack[0][0] ), .A(n5435), .Z(n20069) );
  ANDN U19900 ( .B(\stack[1][10] ), .A(n5206), .Z(n20030) );
  XOR U19901 ( .A(n20035), .B(n20071), .Z(n20029) );
  NANDN U19902 ( .A(n5160), .B(\stack[1][12] ), .Z(n20071) );
  NANDN U19903 ( .A(n5435), .B(\stack[0][1] ), .Z(n20035) );
  ANDN U19904 ( .B(\stack[0][7] ), .A(n5292), .Z(n9314) );
  AND U19905 ( .A(n20072), .B(n20073), .Z(n9315) );
  NANDN U19906 ( .A(n9322), .B(n20074), .Z(n20072) );
  NANDN U19907 ( .A(n9321), .B(n9319), .Z(n20074) );
  XNOR U19908 ( .A(n20043), .B(n20075), .Z(n9319) );
  XNOR U19909 ( .A(n20044), .B(n20045), .Z(n20075) );
  AND U19910 ( .A(n20076), .B(n20077), .Z(n20045) );
  NANDN U19911 ( .A(n20078), .B(n20079), .Z(n20077) );
  NANDN U19912 ( .A(n20080), .B(n20081), .Z(n20076) );
  NANDN U19913 ( .A(n20079), .B(n20078), .Z(n20081) );
  ANDN U19914 ( .B(\stack[0][5] ), .A(n5316), .Z(n20044) );
  XNOR U19915 ( .A(n20050), .B(n20082), .Z(n20043) );
  XNOR U19916 ( .A(n20051), .B(n20052), .Z(n20082) );
  AND U19917 ( .A(n20083), .B(n20084), .Z(n20052) );
  NAND U19918 ( .A(n20085), .B(n20086), .Z(n20084) );
  NANDN U19919 ( .A(n20087), .B(n20088), .Z(n20083) );
  OR U19920 ( .A(n20085), .B(n20086), .Z(n20088) );
  ANDN U19921 ( .B(\stack[0][4] ), .A(n5340), .Z(n20051) );
  XNOR U19922 ( .A(n20057), .B(n20089), .Z(n20050) );
  XNOR U19923 ( .A(n20058), .B(n20059), .Z(n20089) );
  AND U19924 ( .A(n20090), .B(n20091), .Z(n20059) );
  NAND U19925 ( .A(n20092), .B(n20093), .Z(n20091) );
  NAND U19926 ( .A(n20094), .B(n20095), .Z(n20090) );
  OR U19927 ( .A(n20092), .B(n20093), .Z(n20094) );
  ANDN U19928 ( .B(\stack[0][3] ), .A(n5364), .Z(n20058) );
  XNOR U19929 ( .A(n20064), .B(n20096), .Z(n20057) );
  XNOR U19930 ( .A(n20065), .B(n20067), .Z(n20096) );
  ANDN U19931 ( .B(n20097), .A(n20098), .Z(n20067) );
  ANDN U19932 ( .B(\stack[0][0] ), .A(n5411), .Z(n20097) );
  ANDN U19933 ( .B(\stack[0][2] ), .A(n5387), .Z(n20065) );
  XOR U19934 ( .A(n20070), .B(n20099), .Z(n20064) );
  NANDN U19935 ( .A(n5160), .B(\stack[1][11] ), .Z(n20099) );
  NANDN U19936 ( .A(n5411), .B(\stack[0][1] ), .Z(n20070) );
  ANDN U19937 ( .B(\stack[1][5] ), .A(n5302), .Z(n9321) );
  AND U19938 ( .A(n20100), .B(n20101), .Z(n9322) );
  NANDN U19939 ( .A(n9326), .B(n9328), .Z(n20101) );
  NANDN U19940 ( .A(n9329), .B(n20102), .Z(n20100) );
  NANDN U19941 ( .A(n9328), .B(n9326), .Z(n20102) );
  XOR U19942 ( .A(n20078), .B(n20103), .Z(n9326) );
  XNOR U19943 ( .A(n20079), .B(n20080), .Z(n20103) );
  AND U19944 ( .A(n20104), .B(n20105), .Z(n20080) );
  NANDN U19945 ( .A(n20106), .B(n20107), .Z(n20105) );
  NANDN U19946 ( .A(n20108), .B(n20109), .Z(n20104) );
  OR U19947 ( .A(n20107), .B(n20110), .Z(n20109) );
  ANDN U19948 ( .B(\stack[0][4] ), .A(n5316), .Z(n20079) );
  XNOR U19949 ( .A(n20085), .B(n20111), .Z(n20078) );
  XNOR U19950 ( .A(n20086), .B(n20087), .Z(n20111) );
  AND U19951 ( .A(n20112), .B(n20113), .Z(n20087) );
  NAND U19952 ( .A(n20114), .B(n20115), .Z(n20113) );
  NANDN U19953 ( .A(n20116), .B(n20117), .Z(n20112) );
  OR U19954 ( .A(n20114), .B(n20115), .Z(n20117) );
  ANDN U19955 ( .B(\stack[0][3] ), .A(n5340), .Z(n20086) );
  XNOR U19956 ( .A(n20092), .B(n20118), .Z(n20085) );
  XNOR U19957 ( .A(n20093), .B(n20095), .Z(n20118) );
  ANDN U19958 ( .B(n20119), .A(n20120), .Z(n20095) );
  ANDN U19959 ( .B(\stack[1][9] ), .A(n5160), .Z(n20119) );
  ANDN U19960 ( .B(\stack[0][2] ), .A(n5364), .Z(n20093) );
  XOR U19961 ( .A(n20098), .B(n20121), .Z(n20092) );
  NANDN U19962 ( .A(n5160), .B(\stack[1][10] ), .Z(n20121) );
  NANDN U19963 ( .A(n5387), .B(\stack[0][1] ), .Z(n20098) );
  ANDN U19964 ( .B(\stack[0][5] ), .A(n5292), .Z(n9328) );
  AND U19965 ( .A(n20122), .B(n20123), .Z(n9329) );
  NANDN U19966 ( .A(n9334), .B(n9336), .Z(n20123) );
  NANDN U19967 ( .A(n9337), .B(n20124), .Z(n20122) );
  NANDN U19968 ( .A(n9336), .B(n9334), .Z(n20124) );
  XNOR U19969 ( .A(n20107), .B(n20125), .Z(n9334) );
  XOR U19970 ( .A(n20106), .B(n20108), .Z(n20125) );
  AND U19971 ( .A(n20126), .B(n20127), .Z(n20108) );
  NANDN U19972 ( .A(n20128), .B(n20129), .Z(n20127) );
  NAND U19973 ( .A(n20130), .B(n20131), .Z(n20126) );
  NANDN U19974 ( .A(n20129), .B(n20128), .Z(n20130) );
  IV U19975 ( .A(n20110), .Z(n20106) );
  ANDN U19976 ( .B(\stack[0][3] ), .A(n5316), .Z(n20110) );
  XNOR U19977 ( .A(n20114), .B(n20132), .Z(n20107) );
  XOR U19978 ( .A(n20116), .B(n20115), .Z(n20132) );
  ANDN U19979 ( .B(\stack[0][2] ), .A(n5340), .Z(n20115) );
  NANDN U19980 ( .A(n20133), .B(n20134), .Z(n20116) );
  ANDN U19981 ( .B(\stack[1][8] ), .A(n5160), .Z(n20134) );
  XOR U19982 ( .A(n20120), .B(n20135), .Z(n20114) );
  NANDN U19983 ( .A(n5387), .B(\stack[0][0] ), .Z(n20135) );
  NANDN U19984 ( .A(n5364), .B(\stack[0][1] ), .Z(n20120) );
  AND U19985 ( .A(\stack[0][4] ), .B(\stack[1][5] ), .Z(n9336) );
  AND U19986 ( .A(n20136), .B(n20137), .Z(n9337) );
  NANDN U19987 ( .A(n9341), .B(n9343), .Z(n20137) );
  NANDN U19988 ( .A(n9344), .B(n20138), .Z(n20136) );
  NANDN U19989 ( .A(n9343), .B(n9341), .Z(n20138) );
  XNOR U19990 ( .A(n20128), .B(n20139), .Z(n9341) );
  XNOR U19991 ( .A(n20129), .B(n20131), .Z(n20139) );
  ANDN U19992 ( .B(n20140), .A(n20141), .Z(n20131) );
  ANDN U19993 ( .B(\stack[0][0] ), .A(n5340), .Z(n20140) );
  ANDN U19994 ( .B(\stack[1][6] ), .A(n5206), .Z(n20129) );
  XNOR U19995 ( .A(n20133), .B(n20142), .Z(n20128) );
  NANDN U19996 ( .A(n5364), .B(\stack[0][0] ), .Z(n20142) );
  NANDN U19997 ( .A(n5340), .B(\stack[0][1] ), .Z(n20133) );
  ANDN U19998 ( .B(\stack[1][5] ), .A(n5230), .Z(n9343) );
  AND U19999 ( .A(n20143), .B(n20144), .Z(n9344) );
  NANDN U20000 ( .A(n9348), .B(n9350), .Z(n20144) );
  NAND U20001 ( .A(n20145), .B(n9351), .Z(n20143) );
  ANDN U20002 ( .B(n20146), .A(n9356), .Z(n9351) );
  NANDN U20003 ( .A(n5292), .B(\stack[0][1] ), .Z(n9356) );
  ANDN U20004 ( .B(\stack[0][0] ), .A(n5316), .Z(n20146) );
  NANDN U20005 ( .A(n9350), .B(n9348), .Z(n20145) );
  XNOR U20006 ( .A(n20141), .B(n20147), .Z(n9348) );
  NANDN U20007 ( .A(n5160), .B(\stack[1][7] ), .Z(n20147) );
  NANDN U20008 ( .A(n5316), .B(\stack[0][1] ), .Z(n20141) );
  ANDN U20009 ( .B(\stack[1][5] ), .A(n5206), .Z(n9350) );
  ANDN U20010 ( .B(\stack[1][5] ), .A(n6550), .Z(n9358) );
  XNOR U20011 ( .A(n6684), .B(\stack[0][63] ), .Z(n6685) );
  AND U20012 ( .A(n20148), .B(n20149), .Z(n6677) );
  NANDN U20013 ( .A(n6684), .B(n20150), .Z(n20149) );
  NOR U20014 ( .A(n6670), .B(n5173), .Z(n20150) );
  NANDN U20015 ( .A(opcode[0]), .B(opcode[2]), .Z(n5173) );
  NAND U20016 ( .A(n20151), .B(n5175), .Z(n20148) );
  NOR U20017 ( .A(n20152), .B(n20153), .Z(n5175) );
  NANDN U20018 ( .A(\stack[0][63] ), .B(n6684), .Z(n20151) );
  AND U20019 ( .A(n20154), .B(n20155), .Z(n6675) );
  NANDN U20020 ( .A(n6670), .B(n5178), .Z(n20155) );
  AND U20021 ( .A(n20156), .B(n20152), .Z(n5178) );
  XOR U20022 ( .A(n20157), .B(n20158), .Z(n20154) );
  XOR U20023 ( .A(n20159), .B(n20160), .Z(n20158) );
  NAND U20024 ( .A(n20161), .B(n20162), .Z(n20160) );
  NANDN U20025 ( .A(n6667), .B(n20163), .Z(n20162) );
  OR U20026 ( .A(n6666), .B(n6664), .Z(n20163) );
  AND U20027 ( .A(n20164), .B(n20165), .Z(n6667) );
  NANDN U20028 ( .A(n6646), .B(n20166), .Z(n20165) );
  NANDN U20029 ( .A(n6646), .B(n20167), .Z(n20164) );
  NAND U20030 ( .A(n6666), .B(n6664), .Z(n20161) );
  XNOR U20031 ( .A(n20168), .B(n20169), .Z(n6664) );
  NAND U20032 ( .A(n20170), .B(n20171), .Z(n20169) );
  NANDN U20033 ( .A(n6659), .B(n20167), .Z(n20171) );
  AND U20034 ( .A(n20172), .B(n20173), .Z(n20170) );
  NANDN U20035 ( .A(n6646), .B(n6673), .Z(n20173) );
  IV U20036 ( .A(\stack[0][62] ), .Z(n6646) );
  NANDN U20037 ( .A(n6659), .B(n20166), .Z(n20172) );
  NAND U20038 ( .A(n20174), .B(n20175), .Z(n6666) );
  OR U20039 ( .A(n6642), .B(n20176), .Z(n20175) );
  NANDN U20040 ( .A(n6643), .B(n20177), .Z(n20174) );
  NANDN U20041 ( .A(n6640), .B(n6642), .Z(n20177) );
  AND U20042 ( .A(n20178), .B(n20179), .Z(n6642) );
  OR U20043 ( .A(n6618), .B(n20180), .Z(n20179) );
  NANDN U20044 ( .A(n6619), .B(n20181), .Z(n20178) );
  NANDN U20045 ( .A(n6616), .B(n6618), .Z(n20181) );
  AND U20046 ( .A(n20182), .B(n20183), .Z(n6618) );
  OR U20047 ( .A(n6594), .B(n20184), .Z(n20183) );
  NANDN U20048 ( .A(n6595), .B(n20185), .Z(n20182) );
  NANDN U20049 ( .A(n6592), .B(n6594), .Z(n20185) );
  AND U20050 ( .A(n20186), .B(n20187), .Z(n6594) );
  OR U20051 ( .A(n6570), .B(n20188), .Z(n20187) );
  NANDN U20052 ( .A(n6571), .B(n20189), .Z(n20186) );
  NANDN U20053 ( .A(n6568), .B(n6570), .Z(n20189) );
  AND U20054 ( .A(n20190), .B(n20191), .Z(n6570) );
  OR U20055 ( .A(n6546), .B(n20192), .Z(n20191) );
  NANDN U20056 ( .A(n6547), .B(n20193), .Z(n20190) );
  NANDN U20057 ( .A(n6544), .B(n6546), .Z(n20193) );
  AND U20058 ( .A(n20194), .B(n20195), .Z(n6546) );
  OR U20059 ( .A(n6522), .B(n20196), .Z(n20195) );
  NANDN U20060 ( .A(n6523), .B(n20197), .Z(n20194) );
  NANDN U20061 ( .A(n6520), .B(n6522), .Z(n20197) );
  AND U20062 ( .A(n20198), .B(n20199), .Z(n6522) );
  OR U20063 ( .A(n6498), .B(n20200), .Z(n20199) );
  NANDN U20064 ( .A(n6499), .B(n20201), .Z(n20198) );
  NANDN U20065 ( .A(n6496), .B(n6498), .Z(n20201) );
  AND U20066 ( .A(n20202), .B(n20203), .Z(n6498) );
  OR U20067 ( .A(n6474), .B(n20204), .Z(n20203) );
  NANDN U20068 ( .A(n6475), .B(n20205), .Z(n20202) );
  NANDN U20069 ( .A(n6472), .B(n6474), .Z(n20205) );
  AND U20070 ( .A(n20206), .B(n20207), .Z(n6474) );
  OR U20071 ( .A(n6450), .B(n20208), .Z(n20207) );
  NANDN U20072 ( .A(n6451), .B(n20209), .Z(n20206) );
  NANDN U20073 ( .A(n6448), .B(n6450), .Z(n20209) );
  AND U20074 ( .A(n20210), .B(n20211), .Z(n6450) );
  OR U20075 ( .A(n6426), .B(n20212), .Z(n20211) );
  NANDN U20076 ( .A(n6427), .B(n20213), .Z(n20210) );
  NANDN U20077 ( .A(n6424), .B(n6426), .Z(n20213) );
  AND U20078 ( .A(n20214), .B(n20215), .Z(n6426) );
  OR U20079 ( .A(n6402), .B(n20216), .Z(n20215) );
  NANDN U20080 ( .A(n6403), .B(n20217), .Z(n20214) );
  NANDN U20081 ( .A(n6400), .B(n6402), .Z(n20217) );
  AND U20082 ( .A(n20218), .B(n20219), .Z(n6402) );
  OR U20083 ( .A(n6378), .B(n20220), .Z(n20219) );
  NANDN U20084 ( .A(n6379), .B(n20221), .Z(n20218) );
  NANDN U20085 ( .A(n6376), .B(n6378), .Z(n20221) );
  AND U20086 ( .A(n20222), .B(n20223), .Z(n6378) );
  OR U20087 ( .A(n6354), .B(n20224), .Z(n20223) );
  NANDN U20088 ( .A(n6355), .B(n20225), .Z(n20222) );
  NANDN U20089 ( .A(n6352), .B(n6354), .Z(n20225) );
  AND U20090 ( .A(n20226), .B(n20227), .Z(n6354) );
  OR U20091 ( .A(n6330), .B(n20228), .Z(n20227) );
  NANDN U20092 ( .A(n6331), .B(n20229), .Z(n20226) );
  NANDN U20093 ( .A(n6328), .B(n6330), .Z(n20229) );
  AND U20094 ( .A(n20230), .B(n20231), .Z(n6330) );
  OR U20095 ( .A(n6306), .B(n20232), .Z(n20231) );
  NANDN U20096 ( .A(n6307), .B(n20233), .Z(n20230) );
  NANDN U20097 ( .A(n6304), .B(n6306), .Z(n20233) );
  AND U20098 ( .A(n20234), .B(n20235), .Z(n6306) );
  OR U20099 ( .A(n6282), .B(n20236), .Z(n20235) );
  NANDN U20100 ( .A(n6283), .B(n20237), .Z(n20234) );
  NANDN U20101 ( .A(n6280), .B(n6282), .Z(n20237) );
  AND U20102 ( .A(n20238), .B(n20239), .Z(n6282) );
  OR U20103 ( .A(n6258), .B(n20240), .Z(n20239) );
  NANDN U20104 ( .A(n6259), .B(n20241), .Z(n20238) );
  NANDN U20105 ( .A(n6256), .B(n6258), .Z(n20241) );
  AND U20106 ( .A(n20242), .B(n20243), .Z(n6258) );
  OR U20107 ( .A(n6234), .B(n20244), .Z(n20243) );
  NANDN U20108 ( .A(n6235), .B(n20245), .Z(n20242) );
  NANDN U20109 ( .A(n6232), .B(n6234), .Z(n20245) );
  AND U20110 ( .A(n20246), .B(n20247), .Z(n6234) );
  OR U20111 ( .A(n6210), .B(n20248), .Z(n20247) );
  NANDN U20112 ( .A(n6211), .B(n20249), .Z(n20246) );
  NANDN U20113 ( .A(n6208), .B(n6210), .Z(n20249) );
  AND U20114 ( .A(n20250), .B(n20251), .Z(n6210) );
  OR U20115 ( .A(n6186), .B(n20252), .Z(n20251) );
  NANDN U20116 ( .A(n6187), .B(n20253), .Z(n20250) );
  NANDN U20117 ( .A(n6184), .B(n6186), .Z(n20253) );
  AND U20118 ( .A(n20254), .B(n20255), .Z(n6186) );
  OR U20119 ( .A(n6162), .B(n20256), .Z(n20255) );
  NANDN U20120 ( .A(n6163), .B(n20257), .Z(n20254) );
  NANDN U20121 ( .A(n6160), .B(n6162), .Z(n20257) );
  AND U20122 ( .A(n20258), .B(n20259), .Z(n6162) );
  OR U20123 ( .A(n6138), .B(n20260), .Z(n20259) );
  NANDN U20124 ( .A(n6139), .B(n20261), .Z(n20258) );
  NANDN U20125 ( .A(n6136), .B(n6138), .Z(n20261) );
  AND U20126 ( .A(n20262), .B(n20263), .Z(n6138) );
  OR U20127 ( .A(n6114), .B(n20264), .Z(n20263) );
  NANDN U20128 ( .A(n6115), .B(n20265), .Z(n20262) );
  NANDN U20129 ( .A(n6112), .B(n6114), .Z(n20265) );
  AND U20130 ( .A(n20266), .B(n20267), .Z(n6114) );
  OR U20131 ( .A(n6090), .B(n20268), .Z(n20267) );
  NANDN U20132 ( .A(n6091), .B(n20269), .Z(n20266) );
  NANDN U20133 ( .A(n6088), .B(n6090), .Z(n20269) );
  AND U20134 ( .A(n20270), .B(n20271), .Z(n6090) );
  OR U20135 ( .A(n6066), .B(n20272), .Z(n20271) );
  NANDN U20136 ( .A(n6067), .B(n20273), .Z(n20270) );
  NANDN U20137 ( .A(n6064), .B(n6066), .Z(n20273) );
  AND U20138 ( .A(n20274), .B(n20275), .Z(n6066) );
  OR U20139 ( .A(n6042), .B(n20276), .Z(n20275) );
  NANDN U20140 ( .A(n6043), .B(n20277), .Z(n20274) );
  NANDN U20141 ( .A(n6040), .B(n6042), .Z(n20277) );
  AND U20142 ( .A(n20278), .B(n20279), .Z(n6042) );
  OR U20143 ( .A(n6018), .B(n20280), .Z(n20279) );
  NANDN U20144 ( .A(n6019), .B(n20281), .Z(n20278) );
  NANDN U20145 ( .A(n6016), .B(n6018), .Z(n20281) );
  AND U20146 ( .A(n20282), .B(n20283), .Z(n6018) );
  OR U20147 ( .A(n5994), .B(n20284), .Z(n20283) );
  NANDN U20148 ( .A(n5995), .B(n20285), .Z(n20282) );
  NANDN U20149 ( .A(n5992), .B(n5994), .Z(n20285) );
  AND U20150 ( .A(n20286), .B(n20287), .Z(n5994) );
  OR U20151 ( .A(n5970), .B(n20288), .Z(n20287) );
  NANDN U20152 ( .A(n5971), .B(n20289), .Z(n20286) );
  NANDN U20153 ( .A(n5968), .B(n5970), .Z(n20289) );
  AND U20154 ( .A(n20290), .B(n20291), .Z(n5970) );
  OR U20155 ( .A(n5946), .B(n20292), .Z(n20291) );
  NANDN U20156 ( .A(n5947), .B(n20293), .Z(n20290) );
  NANDN U20157 ( .A(n5944), .B(n5946), .Z(n20293) );
  AND U20158 ( .A(n20294), .B(n20295), .Z(n5946) );
  OR U20159 ( .A(n5922), .B(n20296), .Z(n20295) );
  NANDN U20160 ( .A(n5923), .B(n20297), .Z(n20294) );
  NANDN U20161 ( .A(n5920), .B(n5922), .Z(n20297) );
  AND U20162 ( .A(n20298), .B(n20299), .Z(n5922) );
  OR U20163 ( .A(n5898), .B(n20300), .Z(n20299) );
  NANDN U20164 ( .A(n5899), .B(n20301), .Z(n20298) );
  NANDN U20165 ( .A(n5896), .B(n5898), .Z(n20301) );
  AND U20166 ( .A(n20302), .B(n20303), .Z(n5898) );
  OR U20167 ( .A(n5874), .B(n20304), .Z(n20303) );
  NANDN U20168 ( .A(n5875), .B(n20305), .Z(n20302) );
  NANDN U20169 ( .A(n5872), .B(n5874), .Z(n20305) );
  AND U20170 ( .A(n20306), .B(n20307), .Z(n5874) );
  OR U20171 ( .A(n5850), .B(n20308), .Z(n20307) );
  NANDN U20172 ( .A(n5851), .B(n20309), .Z(n20306) );
  NANDN U20173 ( .A(n5848), .B(n5850), .Z(n20309) );
  AND U20174 ( .A(n20310), .B(n20311), .Z(n5850) );
  OR U20175 ( .A(n5826), .B(n20312), .Z(n20311) );
  NANDN U20176 ( .A(n5827), .B(n20313), .Z(n20310) );
  NANDN U20177 ( .A(n5824), .B(n5826), .Z(n20313) );
  AND U20178 ( .A(n20314), .B(n20315), .Z(n5826) );
  OR U20179 ( .A(n5802), .B(n20316), .Z(n20315) );
  NANDN U20180 ( .A(n5803), .B(n20317), .Z(n20314) );
  NANDN U20181 ( .A(n5800), .B(n5802), .Z(n20317) );
  AND U20182 ( .A(n20318), .B(n20319), .Z(n5802) );
  OR U20183 ( .A(n5778), .B(n20320), .Z(n20319) );
  NANDN U20184 ( .A(n5779), .B(n20321), .Z(n20318) );
  NANDN U20185 ( .A(n5776), .B(n5778), .Z(n20321) );
  AND U20186 ( .A(n20322), .B(n20323), .Z(n5778) );
  OR U20187 ( .A(n5754), .B(n20324), .Z(n20323) );
  NANDN U20188 ( .A(n5755), .B(n20325), .Z(n20322) );
  NANDN U20189 ( .A(n5752), .B(n5754), .Z(n20325) );
  AND U20190 ( .A(n20326), .B(n20327), .Z(n5754) );
  OR U20191 ( .A(n5730), .B(n20328), .Z(n20327) );
  NANDN U20192 ( .A(n5731), .B(n20329), .Z(n20326) );
  NANDN U20193 ( .A(n5728), .B(n5730), .Z(n20329) );
  AND U20194 ( .A(n20330), .B(n20331), .Z(n5730) );
  OR U20195 ( .A(n5706), .B(n20332), .Z(n20331) );
  NANDN U20196 ( .A(n5707), .B(n20333), .Z(n20330) );
  NANDN U20197 ( .A(n5704), .B(n5706), .Z(n20333) );
  AND U20198 ( .A(n20334), .B(n20335), .Z(n5706) );
  OR U20199 ( .A(n5682), .B(n20336), .Z(n20335) );
  NANDN U20200 ( .A(n5683), .B(n20337), .Z(n20334) );
  NANDN U20201 ( .A(n5680), .B(n5682), .Z(n20337) );
  AND U20202 ( .A(n20338), .B(n20339), .Z(n5682) );
  OR U20203 ( .A(n5658), .B(n20340), .Z(n20339) );
  NANDN U20204 ( .A(n5659), .B(n20341), .Z(n20338) );
  NANDN U20205 ( .A(n5656), .B(n5658), .Z(n20341) );
  AND U20206 ( .A(n20342), .B(n20343), .Z(n5658) );
  OR U20207 ( .A(n5634), .B(n20344), .Z(n20343) );
  NANDN U20208 ( .A(n5635), .B(n20345), .Z(n20342) );
  NANDN U20209 ( .A(n5632), .B(n5634), .Z(n20345) );
  AND U20210 ( .A(n20346), .B(n20347), .Z(n5634) );
  OR U20211 ( .A(n5610), .B(n20348), .Z(n20347) );
  NANDN U20212 ( .A(n5611), .B(n20349), .Z(n20346) );
  NANDN U20213 ( .A(n5608), .B(n5610), .Z(n20349) );
  AND U20214 ( .A(n20350), .B(n20351), .Z(n5610) );
  OR U20215 ( .A(n5586), .B(n20352), .Z(n20351) );
  NANDN U20216 ( .A(n5587), .B(n20353), .Z(n20350) );
  NANDN U20217 ( .A(n5584), .B(n5586), .Z(n20353) );
  AND U20218 ( .A(n20354), .B(n20355), .Z(n5586) );
  OR U20219 ( .A(n5562), .B(n20356), .Z(n20355) );
  NANDN U20220 ( .A(n5563), .B(n20357), .Z(n20354) );
  NANDN U20221 ( .A(n5560), .B(n5562), .Z(n20357) );
  AND U20222 ( .A(n20358), .B(n20359), .Z(n5562) );
  OR U20223 ( .A(n5538), .B(n20360), .Z(n20359) );
  NANDN U20224 ( .A(n5539), .B(n20361), .Z(n20358) );
  NANDN U20225 ( .A(n5536), .B(n5538), .Z(n20361) );
  AND U20226 ( .A(n20362), .B(n20363), .Z(n5538) );
  OR U20227 ( .A(n5514), .B(n20364), .Z(n20363) );
  NANDN U20228 ( .A(n5515), .B(n20365), .Z(n20362) );
  NANDN U20229 ( .A(n5512), .B(n5514), .Z(n20365) );
  AND U20230 ( .A(n20366), .B(n20367), .Z(n5514) );
  OR U20231 ( .A(n5490), .B(n20368), .Z(n20367) );
  NANDN U20232 ( .A(n5491), .B(n20369), .Z(n20366) );
  NANDN U20233 ( .A(n5488), .B(n5490), .Z(n20369) );
  AND U20234 ( .A(n20370), .B(n20371), .Z(n5490) );
  OR U20235 ( .A(n5466), .B(n20372), .Z(n20371) );
  NANDN U20236 ( .A(n5467), .B(n20373), .Z(n20370) );
  NANDN U20237 ( .A(n5464), .B(n5466), .Z(n20373) );
  AND U20238 ( .A(n20374), .B(n20375), .Z(n5466) );
  OR U20239 ( .A(n5442), .B(n20376), .Z(n20375) );
  NANDN U20240 ( .A(n5443), .B(n20377), .Z(n20374) );
  NANDN U20241 ( .A(n5440), .B(n5442), .Z(n20377) );
  AND U20242 ( .A(n20378), .B(n20379), .Z(n5442) );
  OR U20243 ( .A(n5418), .B(n20380), .Z(n20379) );
  NANDN U20244 ( .A(n5419), .B(n20381), .Z(n20378) );
  NANDN U20245 ( .A(n5416), .B(n5418), .Z(n20381) );
  AND U20246 ( .A(n20382), .B(n20383), .Z(n5418) );
  OR U20247 ( .A(n5394), .B(n5392), .Z(n20383) );
  NANDN U20248 ( .A(n5395), .B(n20384), .Z(n20382) );
  AND U20249 ( .A(n20385), .B(n20386), .Z(n5394) );
  OR U20250 ( .A(n5370), .B(n20387), .Z(n20386) );
  NANDN U20251 ( .A(n5371), .B(n20388), .Z(n20385) );
  NANDN U20252 ( .A(n5368), .B(n5370), .Z(n20388) );
  AND U20253 ( .A(n20389), .B(n20390), .Z(n5370) );
  OR U20254 ( .A(n5346), .B(n20391), .Z(n20390) );
  NANDN U20255 ( .A(n5347), .B(n20392), .Z(n20389) );
  NANDN U20256 ( .A(n5344), .B(n5346), .Z(n20392) );
  AND U20257 ( .A(n20393), .B(n20394), .Z(n5346) );
  OR U20258 ( .A(n5322), .B(n20395), .Z(n20394) );
  NANDN U20259 ( .A(n5323), .B(n20396), .Z(n20393) );
  NANDN U20260 ( .A(n5320), .B(n5322), .Z(n20396) );
  AND U20261 ( .A(n20397), .B(n20398), .Z(n5322) );
  OR U20262 ( .A(n5298), .B(n20399), .Z(n20398) );
  NANDN U20263 ( .A(n5299), .B(n20400), .Z(n20397) );
  NANDN U20264 ( .A(n5296), .B(n5298), .Z(n20400) );
  AND U20265 ( .A(n20401), .B(n20402), .Z(n5298) );
  OR U20266 ( .A(n5274), .B(n20403), .Z(n20402) );
  NANDN U20267 ( .A(n5275), .B(n20404), .Z(n20401) );
  NANDN U20268 ( .A(n5272), .B(n5274), .Z(n20404) );
  AND U20269 ( .A(n20405), .B(n20406), .Z(n5274) );
  OR U20270 ( .A(n5250), .B(n20407), .Z(n20406) );
  NANDN U20271 ( .A(n5251), .B(n20408), .Z(n20405) );
  NANDN U20272 ( .A(n5248), .B(n5250), .Z(n20408) );
  AND U20273 ( .A(n20409), .B(n20410), .Z(n5250) );
  OR U20274 ( .A(n5226), .B(n20411), .Z(n20410) );
  NANDN U20275 ( .A(n5227), .B(n20412), .Z(n20409) );
  NANDN U20276 ( .A(n5224), .B(n5226), .Z(n20412) );
  AND U20277 ( .A(n20413), .B(n20414), .Z(n5226) );
  OR U20278 ( .A(n5202), .B(n20415), .Z(n20414) );
  NANDN U20279 ( .A(n5203), .B(n20416), .Z(n20413) );
  NANDN U20280 ( .A(n5200), .B(n5202), .Z(n20416) );
  AND U20281 ( .A(n20417), .B(n20418), .Z(n5202) );
  NANDN U20282 ( .A(n20168), .B(n20419), .Z(n20418) );
  NANDN U20283 ( .A(n5182), .B(n20420), .Z(n20417) );
  NANDN U20284 ( .A(n20419), .B(n20168), .Z(n20420) );
  IV U20285 ( .A(n5179), .Z(n20419) );
  XOR U20286 ( .A(n20168), .B(n20421), .Z(n5179) );
  NAND U20287 ( .A(n20422), .B(n20423), .Z(n20421) );
  NANDN U20288 ( .A(n5169), .B(n20167), .Z(n20423) );
  AND U20289 ( .A(n20424), .B(n20425), .Z(n20422) );
  NANDN U20290 ( .A(n5160), .B(n6673), .Z(n20425) );
  NANDN U20291 ( .A(n5169), .B(n20166), .Z(n20424) );
  AND U20292 ( .A(n20426), .B(n20427), .Z(n5182) );
  NANDN U20293 ( .A(n5160), .B(n20166), .Z(n20427) );
  NANDN U20294 ( .A(n5160), .B(n20167), .Z(n20426) );
  IV U20295 ( .A(n20415), .Z(n5200) );
  XOR U20296 ( .A(n20168), .B(n20428), .Z(n20415) );
  NAND U20297 ( .A(n20429), .B(n20430), .Z(n20428) );
  NANDN U20298 ( .A(n5195), .B(n20167), .Z(n20430) );
  AND U20299 ( .A(n20431), .B(n20432), .Z(n20429) );
  NAND U20300 ( .A(\stack[0][1] ), .B(n6673), .Z(n20432) );
  NANDN U20301 ( .A(n5195), .B(n20166), .Z(n20431) );
  AND U20302 ( .A(n20433), .B(n20434), .Z(n5203) );
  NAND U20303 ( .A(\stack[0][1] ), .B(n20166), .Z(n20434) );
  NAND U20304 ( .A(\stack[0][1] ), .B(n20167), .Z(n20433) );
  IV U20305 ( .A(n20411), .Z(n5224) );
  XOR U20306 ( .A(n20168), .B(n20435), .Z(n20411) );
  NAND U20307 ( .A(n20436), .B(n20437), .Z(n20435) );
  NANDN U20308 ( .A(n5219), .B(n20167), .Z(n20437) );
  AND U20309 ( .A(n20438), .B(n20439), .Z(n20436) );
  NANDN U20310 ( .A(n5206), .B(n6673), .Z(n20439) );
  NANDN U20311 ( .A(n5219), .B(n20166), .Z(n20438) );
  AND U20312 ( .A(n20440), .B(n20441), .Z(n5227) );
  NANDN U20313 ( .A(n5206), .B(n20166), .Z(n20441) );
  NANDN U20314 ( .A(n5206), .B(n20167), .Z(n20440) );
  IV U20315 ( .A(n20407), .Z(n5248) );
  XOR U20316 ( .A(n20168), .B(n20442), .Z(n20407) );
  NAND U20317 ( .A(n20443), .B(n20444), .Z(n20442) );
  NANDN U20318 ( .A(n5243), .B(n20167), .Z(n20444) );
  AND U20319 ( .A(n20445), .B(n20446), .Z(n20443) );
  NANDN U20320 ( .A(n5230), .B(n6673), .Z(n20446) );
  NANDN U20321 ( .A(n5243), .B(n20166), .Z(n20445) );
  AND U20322 ( .A(n20447), .B(n20448), .Z(n5251) );
  NANDN U20323 ( .A(n5230), .B(n20166), .Z(n20448) );
  NANDN U20324 ( .A(n5230), .B(n20167), .Z(n20447) );
  IV U20325 ( .A(n20403), .Z(n5272) );
  XOR U20326 ( .A(n20168), .B(n20449), .Z(n20403) );
  NAND U20327 ( .A(n20450), .B(n20451), .Z(n20449) );
  NANDN U20328 ( .A(n5267), .B(n20167), .Z(n20451) );
  AND U20329 ( .A(n20452), .B(n20453), .Z(n20450) );
  NANDN U20330 ( .A(n5254), .B(n6673), .Z(n20453) );
  NANDN U20331 ( .A(n5267), .B(n20166), .Z(n20452) );
  AND U20332 ( .A(n20454), .B(n20455), .Z(n5275) );
  NANDN U20333 ( .A(n5254), .B(n20166), .Z(n20455) );
  NANDN U20334 ( .A(n5254), .B(n20167), .Z(n20454) );
  IV U20335 ( .A(n20399), .Z(n5296) );
  XOR U20336 ( .A(n20168), .B(n20456), .Z(n20399) );
  NAND U20337 ( .A(n20457), .B(n20458), .Z(n20456) );
  NANDN U20338 ( .A(n5292), .B(n20167), .Z(n20458) );
  AND U20339 ( .A(n20459), .B(n20460), .Z(n20457) );
  NANDN U20340 ( .A(n5278), .B(n6673), .Z(n20460) );
  NANDN U20341 ( .A(n5292), .B(n20166), .Z(n20459) );
  AND U20342 ( .A(n20461), .B(n20462), .Z(n5299) );
  NANDN U20343 ( .A(n5278), .B(n20166), .Z(n20462) );
  NANDN U20344 ( .A(n5278), .B(n20167), .Z(n20461) );
  IV U20345 ( .A(n20395), .Z(n5320) );
  XOR U20346 ( .A(n20168), .B(n20463), .Z(n20395) );
  NAND U20347 ( .A(n20464), .B(n20465), .Z(n20463) );
  NANDN U20348 ( .A(n5316), .B(n20167), .Z(n20465) );
  AND U20349 ( .A(n20466), .B(n20467), .Z(n20464) );
  NANDN U20350 ( .A(n5302), .B(n6673), .Z(n20467) );
  NANDN U20351 ( .A(n5316), .B(n20166), .Z(n20466) );
  AND U20352 ( .A(n20468), .B(n20469), .Z(n5323) );
  NANDN U20353 ( .A(n5302), .B(n20166), .Z(n20469) );
  NANDN U20354 ( .A(n5302), .B(n20167), .Z(n20468) );
  IV U20355 ( .A(n20391), .Z(n5344) );
  XOR U20356 ( .A(n20168), .B(n20470), .Z(n20391) );
  NAND U20357 ( .A(n20471), .B(n20472), .Z(n20470) );
  NANDN U20358 ( .A(n5340), .B(n20167), .Z(n20472) );
  AND U20359 ( .A(n20473), .B(n20474), .Z(n20471) );
  NANDN U20360 ( .A(n5326), .B(n6673), .Z(n20474) );
  NANDN U20361 ( .A(n5340), .B(n20166), .Z(n20473) );
  AND U20362 ( .A(n20475), .B(n20476), .Z(n5347) );
  NANDN U20363 ( .A(n5326), .B(n20166), .Z(n20476) );
  NANDN U20364 ( .A(n5326), .B(n20167), .Z(n20475) );
  IV U20365 ( .A(n20387), .Z(n5368) );
  XOR U20366 ( .A(n20168), .B(n20477), .Z(n20387) );
  NAND U20367 ( .A(n20478), .B(n20479), .Z(n20477) );
  NANDN U20368 ( .A(n5364), .B(n20167), .Z(n20479) );
  AND U20369 ( .A(n20480), .B(n20481), .Z(n20478) );
  NANDN U20370 ( .A(n5350), .B(n6673), .Z(n20481) );
  NANDN U20371 ( .A(n5364), .B(n20166), .Z(n20480) );
  AND U20372 ( .A(n20482), .B(n20483), .Z(n5371) );
  NANDN U20373 ( .A(n5350), .B(n20166), .Z(n20483) );
  NANDN U20374 ( .A(n5350), .B(n20167), .Z(n20482) );
  XOR U20375 ( .A(n20484), .B(n5181), .Z(n5392) );
  AND U20376 ( .A(n20485), .B(n20486), .Z(n20484) );
  NANDN U20377 ( .A(n5387), .B(n20167), .Z(n20486) );
  AND U20378 ( .A(n20487), .B(n20488), .Z(n20485) );
  NANDN U20379 ( .A(n5374), .B(n6673), .Z(n20488) );
  NANDN U20380 ( .A(n5387), .B(n20166), .Z(n20487) );
  AND U20381 ( .A(n20489), .B(n20490), .Z(n5395) );
  NANDN U20382 ( .A(n5374), .B(n20166), .Z(n20490) );
  NANDN U20383 ( .A(n5374), .B(n20167), .Z(n20489) );
  IV U20384 ( .A(n20380), .Z(n5416) );
  XOR U20385 ( .A(n20168), .B(n20491), .Z(n20380) );
  NAND U20386 ( .A(n20492), .B(n20493), .Z(n20491) );
  NANDN U20387 ( .A(n5411), .B(n20167), .Z(n20493) );
  AND U20388 ( .A(n20494), .B(n20495), .Z(n20492) );
  NANDN U20389 ( .A(n5398), .B(n6673), .Z(n20495) );
  NANDN U20390 ( .A(n5411), .B(n20166), .Z(n20494) );
  AND U20391 ( .A(n20496), .B(n20497), .Z(n5419) );
  NANDN U20392 ( .A(n5398), .B(n20166), .Z(n20497) );
  NANDN U20393 ( .A(n5398), .B(n20167), .Z(n20496) );
  IV U20394 ( .A(\stack[0][10] ), .Z(n5398) );
  IV U20395 ( .A(n20376), .Z(n5440) );
  XOR U20396 ( .A(n20168), .B(n20498), .Z(n20376) );
  NAND U20397 ( .A(n20499), .B(n20500), .Z(n20498) );
  NANDN U20398 ( .A(n5435), .B(n20167), .Z(n20500) );
  AND U20399 ( .A(n20501), .B(n20502), .Z(n20499) );
  NANDN U20400 ( .A(n5422), .B(n6673), .Z(n20502) );
  NANDN U20401 ( .A(n5435), .B(n20166), .Z(n20501) );
  AND U20402 ( .A(n20503), .B(n20504), .Z(n5443) );
  NANDN U20403 ( .A(n5422), .B(n20166), .Z(n20504) );
  NANDN U20404 ( .A(n5422), .B(n20167), .Z(n20503) );
  IV U20405 ( .A(\stack[0][11] ), .Z(n5422) );
  IV U20406 ( .A(n20372), .Z(n5464) );
  XOR U20407 ( .A(n20168), .B(n20505), .Z(n20372) );
  NAND U20408 ( .A(n20506), .B(n20507), .Z(n20505) );
  NANDN U20409 ( .A(n5459), .B(n20167), .Z(n20507) );
  AND U20410 ( .A(n20508), .B(n20509), .Z(n20506) );
  NANDN U20411 ( .A(n5446), .B(n6673), .Z(n20509) );
  NANDN U20412 ( .A(n5459), .B(n20166), .Z(n20508) );
  AND U20413 ( .A(n20510), .B(n20511), .Z(n5467) );
  NANDN U20414 ( .A(n5446), .B(n20166), .Z(n20511) );
  NANDN U20415 ( .A(n5446), .B(n20167), .Z(n20510) );
  IV U20416 ( .A(\stack[0][12] ), .Z(n5446) );
  IV U20417 ( .A(n20368), .Z(n5488) );
  XOR U20418 ( .A(n20168), .B(n20512), .Z(n20368) );
  NAND U20419 ( .A(n20513), .B(n20514), .Z(n20512) );
  NANDN U20420 ( .A(n5483), .B(n20167), .Z(n20514) );
  AND U20421 ( .A(n20515), .B(n20516), .Z(n20513) );
  NANDN U20422 ( .A(n5470), .B(n6673), .Z(n20516) );
  NANDN U20423 ( .A(n5483), .B(n20166), .Z(n20515) );
  AND U20424 ( .A(n20517), .B(n20518), .Z(n5491) );
  NANDN U20425 ( .A(n5470), .B(n20166), .Z(n20518) );
  NANDN U20426 ( .A(n5470), .B(n20167), .Z(n20517) );
  IV U20427 ( .A(\stack[0][13] ), .Z(n5470) );
  IV U20428 ( .A(n20364), .Z(n5512) );
  XOR U20429 ( .A(n20168), .B(n20519), .Z(n20364) );
  NAND U20430 ( .A(n20520), .B(n20521), .Z(n20519) );
  NANDN U20431 ( .A(n5507), .B(n20167), .Z(n20521) );
  AND U20432 ( .A(n20522), .B(n20523), .Z(n20520) );
  NANDN U20433 ( .A(n5494), .B(n6673), .Z(n20523) );
  NANDN U20434 ( .A(n5507), .B(n20166), .Z(n20522) );
  AND U20435 ( .A(n20524), .B(n20525), .Z(n5515) );
  NANDN U20436 ( .A(n5494), .B(n20166), .Z(n20525) );
  NANDN U20437 ( .A(n5494), .B(n20167), .Z(n20524) );
  IV U20438 ( .A(\stack[0][14] ), .Z(n5494) );
  IV U20439 ( .A(n20360), .Z(n5536) );
  XOR U20440 ( .A(n20168), .B(n20526), .Z(n20360) );
  NAND U20441 ( .A(n20527), .B(n20528), .Z(n20526) );
  NANDN U20442 ( .A(n5531), .B(n20167), .Z(n20528) );
  AND U20443 ( .A(n20529), .B(n20530), .Z(n20527) );
  NANDN U20444 ( .A(n5518), .B(n6673), .Z(n20530) );
  NANDN U20445 ( .A(n5531), .B(n20166), .Z(n20529) );
  AND U20446 ( .A(n20531), .B(n20532), .Z(n5539) );
  NANDN U20447 ( .A(n5518), .B(n20166), .Z(n20532) );
  NANDN U20448 ( .A(n5518), .B(n20167), .Z(n20531) );
  IV U20449 ( .A(\stack[0][15] ), .Z(n5518) );
  IV U20450 ( .A(n20356), .Z(n5560) );
  XOR U20451 ( .A(n20168), .B(n20533), .Z(n20356) );
  NAND U20452 ( .A(n20534), .B(n20535), .Z(n20533) );
  NANDN U20453 ( .A(n5555), .B(n20167), .Z(n20535) );
  AND U20454 ( .A(n20536), .B(n20537), .Z(n20534) );
  NANDN U20455 ( .A(n5542), .B(n6673), .Z(n20537) );
  NANDN U20456 ( .A(n5555), .B(n20166), .Z(n20536) );
  AND U20457 ( .A(n20538), .B(n20539), .Z(n5563) );
  NANDN U20458 ( .A(n5542), .B(n20166), .Z(n20539) );
  NANDN U20459 ( .A(n5542), .B(n20167), .Z(n20538) );
  IV U20460 ( .A(\stack[0][16] ), .Z(n5542) );
  IV U20461 ( .A(n20352), .Z(n5584) );
  XOR U20462 ( .A(n20168), .B(n20540), .Z(n20352) );
  NAND U20463 ( .A(n20541), .B(n20542), .Z(n20540) );
  NANDN U20464 ( .A(n5579), .B(n20167), .Z(n20542) );
  AND U20465 ( .A(n20543), .B(n20544), .Z(n20541) );
  NANDN U20466 ( .A(n5566), .B(n6673), .Z(n20544) );
  NANDN U20467 ( .A(n5579), .B(n20166), .Z(n20543) );
  AND U20468 ( .A(n20545), .B(n20546), .Z(n5587) );
  NANDN U20469 ( .A(n5566), .B(n20166), .Z(n20546) );
  NANDN U20470 ( .A(n5566), .B(n20167), .Z(n20545) );
  IV U20471 ( .A(\stack[0][17] ), .Z(n5566) );
  IV U20472 ( .A(n20348), .Z(n5608) );
  XOR U20473 ( .A(n20168), .B(n20547), .Z(n20348) );
  NAND U20474 ( .A(n20548), .B(n20549), .Z(n20547) );
  NANDN U20475 ( .A(n5603), .B(n20167), .Z(n20549) );
  AND U20476 ( .A(n20550), .B(n20551), .Z(n20548) );
  NANDN U20477 ( .A(n5590), .B(n6673), .Z(n20551) );
  NANDN U20478 ( .A(n5603), .B(n20166), .Z(n20550) );
  AND U20479 ( .A(n20552), .B(n20553), .Z(n5611) );
  NANDN U20480 ( .A(n5590), .B(n20166), .Z(n20553) );
  NANDN U20481 ( .A(n5590), .B(n20167), .Z(n20552) );
  IV U20482 ( .A(\stack[0][18] ), .Z(n5590) );
  IV U20483 ( .A(n20344), .Z(n5632) );
  XOR U20484 ( .A(n20168), .B(n20554), .Z(n20344) );
  NAND U20485 ( .A(n20555), .B(n20556), .Z(n20554) );
  NANDN U20486 ( .A(n5627), .B(n20167), .Z(n20556) );
  AND U20487 ( .A(n20557), .B(n20558), .Z(n20555) );
  NANDN U20488 ( .A(n5614), .B(n6673), .Z(n20558) );
  NANDN U20489 ( .A(n5627), .B(n20166), .Z(n20557) );
  AND U20490 ( .A(n20559), .B(n20560), .Z(n5635) );
  NANDN U20491 ( .A(n5614), .B(n20166), .Z(n20560) );
  NANDN U20492 ( .A(n5614), .B(n20167), .Z(n20559) );
  IV U20493 ( .A(\stack[0][19] ), .Z(n5614) );
  IV U20494 ( .A(n20340), .Z(n5656) );
  XOR U20495 ( .A(n20168), .B(n20561), .Z(n20340) );
  NAND U20496 ( .A(n20562), .B(n20563), .Z(n20561) );
  NANDN U20497 ( .A(n5651), .B(n20167), .Z(n20563) );
  AND U20498 ( .A(n20564), .B(n20565), .Z(n20562) );
  NANDN U20499 ( .A(n5638), .B(n6673), .Z(n20565) );
  NANDN U20500 ( .A(n5651), .B(n20166), .Z(n20564) );
  AND U20501 ( .A(n20566), .B(n20567), .Z(n5659) );
  NANDN U20502 ( .A(n5638), .B(n20166), .Z(n20567) );
  NANDN U20503 ( .A(n5638), .B(n20167), .Z(n20566) );
  IV U20504 ( .A(\stack[0][20] ), .Z(n5638) );
  IV U20505 ( .A(n20336), .Z(n5680) );
  XOR U20506 ( .A(n20168), .B(n20568), .Z(n20336) );
  NAND U20507 ( .A(n20569), .B(n20570), .Z(n20568) );
  NANDN U20508 ( .A(n5675), .B(n20167), .Z(n20570) );
  AND U20509 ( .A(n20571), .B(n20572), .Z(n20569) );
  NANDN U20510 ( .A(n5662), .B(n6673), .Z(n20572) );
  NANDN U20511 ( .A(n5675), .B(n20166), .Z(n20571) );
  AND U20512 ( .A(n20573), .B(n20574), .Z(n5683) );
  NANDN U20513 ( .A(n5662), .B(n20166), .Z(n20574) );
  NANDN U20514 ( .A(n5662), .B(n20167), .Z(n20573) );
  IV U20515 ( .A(\stack[0][21] ), .Z(n5662) );
  IV U20516 ( .A(n20332), .Z(n5704) );
  XOR U20517 ( .A(n20168), .B(n20575), .Z(n20332) );
  NAND U20518 ( .A(n20576), .B(n20577), .Z(n20575) );
  NANDN U20519 ( .A(n5699), .B(n20167), .Z(n20577) );
  AND U20520 ( .A(n20578), .B(n20579), .Z(n20576) );
  NANDN U20521 ( .A(n5686), .B(n6673), .Z(n20579) );
  NANDN U20522 ( .A(n5699), .B(n20166), .Z(n20578) );
  AND U20523 ( .A(n20580), .B(n20581), .Z(n5707) );
  NANDN U20524 ( .A(n5686), .B(n20166), .Z(n20581) );
  NANDN U20525 ( .A(n5686), .B(n20167), .Z(n20580) );
  IV U20526 ( .A(\stack[0][22] ), .Z(n5686) );
  IV U20527 ( .A(n20328), .Z(n5728) );
  XOR U20528 ( .A(n20168), .B(n20582), .Z(n20328) );
  NAND U20529 ( .A(n20583), .B(n20584), .Z(n20582) );
  NANDN U20530 ( .A(n5723), .B(n20167), .Z(n20584) );
  AND U20531 ( .A(n20585), .B(n20586), .Z(n20583) );
  NANDN U20532 ( .A(n5710), .B(n6673), .Z(n20586) );
  NANDN U20533 ( .A(n5723), .B(n20166), .Z(n20585) );
  AND U20534 ( .A(n20587), .B(n20588), .Z(n5731) );
  NANDN U20535 ( .A(n5710), .B(n20166), .Z(n20588) );
  NANDN U20536 ( .A(n5710), .B(n20167), .Z(n20587) );
  IV U20537 ( .A(\stack[0][23] ), .Z(n5710) );
  IV U20538 ( .A(n20324), .Z(n5752) );
  XOR U20539 ( .A(n20168), .B(n20589), .Z(n20324) );
  NAND U20540 ( .A(n20590), .B(n20591), .Z(n20589) );
  NANDN U20541 ( .A(n5747), .B(n20167), .Z(n20591) );
  AND U20542 ( .A(n20592), .B(n20593), .Z(n20590) );
  NANDN U20543 ( .A(n5734), .B(n6673), .Z(n20593) );
  NANDN U20544 ( .A(n5747), .B(n20166), .Z(n20592) );
  AND U20545 ( .A(n20594), .B(n20595), .Z(n5755) );
  NANDN U20546 ( .A(n5734), .B(n20166), .Z(n20595) );
  NANDN U20547 ( .A(n5734), .B(n20167), .Z(n20594) );
  IV U20548 ( .A(\stack[0][24] ), .Z(n5734) );
  IV U20549 ( .A(n20320), .Z(n5776) );
  XOR U20550 ( .A(n20168), .B(n20596), .Z(n20320) );
  NAND U20551 ( .A(n20597), .B(n20598), .Z(n20596) );
  NANDN U20552 ( .A(n5771), .B(n20167), .Z(n20598) );
  AND U20553 ( .A(n20599), .B(n20600), .Z(n20597) );
  NANDN U20554 ( .A(n5758), .B(n6673), .Z(n20600) );
  NANDN U20555 ( .A(n5771), .B(n20166), .Z(n20599) );
  AND U20556 ( .A(n20601), .B(n20602), .Z(n5779) );
  NANDN U20557 ( .A(n5758), .B(n20166), .Z(n20602) );
  NANDN U20558 ( .A(n5758), .B(n20167), .Z(n20601) );
  IV U20559 ( .A(\stack[0][25] ), .Z(n5758) );
  IV U20560 ( .A(n20316), .Z(n5800) );
  XOR U20561 ( .A(n20168), .B(n20603), .Z(n20316) );
  NAND U20562 ( .A(n20604), .B(n20605), .Z(n20603) );
  NANDN U20563 ( .A(n5795), .B(n20167), .Z(n20605) );
  AND U20564 ( .A(n20606), .B(n20607), .Z(n20604) );
  NANDN U20565 ( .A(n5782), .B(n6673), .Z(n20607) );
  NANDN U20566 ( .A(n5795), .B(n20166), .Z(n20606) );
  AND U20567 ( .A(n20608), .B(n20609), .Z(n5803) );
  NANDN U20568 ( .A(n5782), .B(n20166), .Z(n20609) );
  NANDN U20569 ( .A(n5782), .B(n20167), .Z(n20608) );
  IV U20570 ( .A(\stack[0][26] ), .Z(n5782) );
  IV U20571 ( .A(n20312), .Z(n5824) );
  XOR U20572 ( .A(n20168), .B(n20610), .Z(n20312) );
  NAND U20573 ( .A(n20611), .B(n20612), .Z(n20610) );
  NANDN U20574 ( .A(n5819), .B(n20167), .Z(n20612) );
  AND U20575 ( .A(n20613), .B(n20614), .Z(n20611) );
  NANDN U20576 ( .A(n5806), .B(n6673), .Z(n20614) );
  NANDN U20577 ( .A(n5819), .B(n20166), .Z(n20613) );
  AND U20578 ( .A(n20615), .B(n20616), .Z(n5827) );
  NANDN U20579 ( .A(n5806), .B(n20166), .Z(n20616) );
  NANDN U20580 ( .A(n5806), .B(n20167), .Z(n20615) );
  IV U20581 ( .A(\stack[0][27] ), .Z(n5806) );
  IV U20582 ( .A(n20308), .Z(n5848) );
  XOR U20583 ( .A(n20168), .B(n20617), .Z(n20308) );
  NAND U20584 ( .A(n20618), .B(n20619), .Z(n20617) );
  NANDN U20585 ( .A(n5843), .B(n20167), .Z(n20619) );
  AND U20586 ( .A(n20620), .B(n20621), .Z(n20618) );
  NANDN U20587 ( .A(n5830), .B(n6673), .Z(n20621) );
  NANDN U20588 ( .A(n5843), .B(n20166), .Z(n20620) );
  AND U20589 ( .A(n20622), .B(n20623), .Z(n5851) );
  NANDN U20590 ( .A(n5830), .B(n20166), .Z(n20623) );
  NANDN U20591 ( .A(n5830), .B(n20167), .Z(n20622) );
  IV U20592 ( .A(\stack[0][28] ), .Z(n5830) );
  IV U20593 ( .A(n20304), .Z(n5872) );
  XOR U20594 ( .A(n20168), .B(n20624), .Z(n20304) );
  NAND U20595 ( .A(n20625), .B(n20626), .Z(n20624) );
  NANDN U20596 ( .A(n5867), .B(n20167), .Z(n20626) );
  AND U20597 ( .A(n20627), .B(n20628), .Z(n20625) );
  NANDN U20598 ( .A(n5854), .B(n6673), .Z(n20628) );
  NANDN U20599 ( .A(n5867), .B(n20166), .Z(n20627) );
  AND U20600 ( .A(n20629), .B(n20630), .Z(n5875) );
  NANDN U20601 ( .A(n5854), .B(n20166), .Z(n20630) );
  NANDN U20602 ( .A(n5854), .B(n20167), .Z(n20629) );
  IV U20603 ( .A(\stack[0][29] ), .Z(n5854) );
  IV U20604 ( .A(n20300), .Z(n5896) );
  XOR U20605 ( .A(n20168), .B(n20631), .Z(n20300) );
  NAND U20606 ( .A(n20632), .B(n20633), .Z(n20631) );
  NANDN U20607 ( .A(n5891), .B(n20167), .Z(n20633) );
  AND U20608 ( .A(n20634), .B(n20635), .Z(n20632) );
  NANDN U20609 ( .A(n5878), .B(n6673), .Z(n20635) );
  NANDN U20610 ( .A(n5891), .B(n20166), .Z(n20634) );
  AND U20611 ( .A(n20636), .B(n20637), .Z(n5899) );
  NANDN U20612 ( .A(n5878), .B(n20166), .Z(n20637) );
  NANDN U20613 ( .A(n5878), .B(n20167), .Z(n20636) );
  IV U20614 ( .A(\stack[0][30] ), .Z(n5878) );
  IV U20615 ( .A(n20296), .Z(n5920) );
  XOR U20616 ( .A(n20168), .B(n20638), .Z(n20296) );
  NAND U20617 ( .A(n20639), .B(n20640), .Z(n20638) );
  NANDN U20618 ( .A(n5915), .B(n20167), .Z(n20640) );
  AND U20619 ( .A(n20641), .B(n20642), .Z(n20639) );
  NANDN U20620 ( .A(n5902), .B(n6673), .Z(n20642) );
  NANDN U20621 ( .A(n5915), .B(n20166), .Z(n20641) );
  AND U20622 ( .A(n20643), .B(n20644), .Z(n5923) );
  NANDN U20623 ( .A(n5902), .B(n20166), .Z(n20644) );
  NANDN U20624 ( .A(n5902), .B(n20167), .Z(n20643) );
  IV U20625 ( .A(\stack[0][31] ), .Z(n5902) );
  IV U20626 ( .A(n20292), .Z(n5944) );
  XOR U20627 ( .A(n20168), .B(n20645), .Z(n20292) );
  NAND U20628 ( .A(n20646), .B(n20647), .Z(n20645) );
  NANDN U20629 ( .A(n5940), .B(n20167), .Z(n20647) );
  AND U20630 ( .A(n20648), .B(n20649), .Z(n20646) );
  NANDN U20631 ( .A(n5926), .B(n6673), .Z(n20649) );
  NANDN U20632 ( .A(n5940), .B(n20166), .Z(n20648) );
  AND U20633 ( .A(n20650), .B(n20651), .Z(n5947) );
  NANDN U20634 ( .A(n5926), .B(n20166), .Z(n20651) );
  NANDN U20635 ( .A(n5926), .B(n20167), .Z(n20650) );
  IV U20636 ( .A(\stack[0][32] ), .Z(n5926) );
  IV U20637 ( .A(n20288), .Z(n5968) );
  XOR U20638 ( .A(n20168), .B(n20652), .Z(n20288) );
  NAND U20639 ( .A(n20653), .B(n20654), .Z(n20652) );
  NANDN U20640 ( .A(n5964), .B(n20167), .Z(n20654) );
  AND U20641 ( .A(n20655), .B(n20656), .Z(n20653) );
  NANDN U20642 ( .A(n5950), .B(n6673), .Z(n20656) );
  NANDN U20643 ( .A(n5964), .B(n20166), .Z(n20655) );
  AND U20644 ( .A(n20657), .B(n20658), .Z(n5971) );
  NANDN U20645 ( .A(n5950), .B(n20166), .Z(n20658) );
  NANDN U20646 ( .A(n5950), .B(n20167), .Z(n20657) );
  IV U20647 ( .A(\stack[0][33] ), .Z(n5950) );
  IV U20648 ( .A(n20284), .Z(n5992) );
  XOR U20649 ( .A(n20168), .B(n20659), .Z(n20284) );
  NAND U20650 ( .A(n20660), .B(n20661), .Z(n20659) );
  NANDN U20651 ( .A(n5988), .B(n20167), .Z(n20661) );
  AND U20652 ( .A(n20662), .B(n20663), .Z(n20660) );
  NANDN U20653 ( .A(n5974), .B(n6673), .Z(n20663) );
  NANDN U20654 ( .A(n5988), .B(n20166), .Z(n20662) );
  AND U20655 ( .A(n20664), .B(n20665), .Z(n5995) );
  NANDN U20656 ( .A(n5974), .B(n20166), .Z(n20665) );
  NANDN U20657 ( .A(n5974), .B(n20167), .Z(n20664) );
  IV U20658 ( .A(\stack[0][34] ), .Z(n5974) );
  IV U20659 ( .A(n20280), .Z(n6016) );
  XOR U20660 ( .A(n20168), .B(n20666), .Z(n20280) );
  NAND U20661 ( .A(n20667), .B(n20668), .Z(n20666) );
  NANDN U20662 ( .A(n6012), .B(n20167), .Z(n20668) );
  AND U20663 ( .A(n20669), .B(n20670), .Z(n20667) );
  NANDN U20664 ( .A(n5998), .B(n6673), .Z(n20670) );
  NANDN U20665 ( .A(n6012), .B(n20166), .Z(n20669) );
  AND U20666 ( .A(n20671), .B(n20672), .Z(n6019) );
  NANDN U20667 ( .A(n5998), .B(n20166), .Z(n20672) );
  NANDN U20668 ( .A(n5998), .B(n20167), .Z(n20671) );
  IV U20669 ( .A(\stack[0][35] ), .Z(n5998) );
  IV U20670 ( .A(n20276), .Z(n6040) );
  XOR U20671 ( .A(n20168), .B(n20673), .Z(n20276) );
  NAND U20672 ( .A(n20674), .B(n20675), .Z(n20673) );
  NANDN U20673 ( .A(n6036), .B(n20167), .Z(n20675) );
  AND U20674 ( .A(n20676), .B(n20677), .Z(n20674) );
  NANDN U20675 ( .A(n6022), .B(n6673), .Z(n20677) );
  NANDN U20676 ( .A(n6036), .B(n20166), .Z(n20676) );
  AND U20677 ( .A(n20678), .B(n20679), .Z(n6043) );
  NANDN U20678 ( .A(n6022), .B(n20166), .Z(n20679) );
  NANDN U20679 ( .A(n6022), .B(n20167), .Z(n20678) );
  IV U20680 ( .A(\stack[0][36] ), .Z(n6022) );
  IV U20681 ( .A(n20272), .Z(n6064) );
  XOR U20682 ( .A(n20168), .B(n20680), .Z(n20272) );
  NAND U20683 ( .A(n20681), .B(n20682), .Z(n20680) );
  NANDN U20684 ( .A(n6060), .B(n20167), .Z(n20682) );
  AND U20685 ( .A(n20683), .B(n20684), .Z(n20681) );
  NANDN U20686 ( .A(n6046), .B(n6673), .Z(n20684) );
  NANDN U20687 ( .A(n6060), .B(n20166), .Z(n20683) );
  AND U20688 ( .A(n20685), .B(n20686), .Z(n6067) );
  NANDN U20689 ( .A(n6046), .B(n20166), .Z(n20686) );
  NANDN U20690 ( .A(n6046), .B(n20167), .Z(n20685) );
  IV U20691 ( .A(\stack[0][37] ), .Z(n6046) );
  IV U20692 ( .A(n20268), .Z(n6088) );
  XOR U20693 ( .A(n20168), .B(n20687), .Z(n20268) );
  NAND U20694 ( .A(n20688), .B(n20689), .Z(n20687) );
  NANDN U20695 ( .A(n6084), .B(n20167), .Z(n20689) );
  AND U20696 ( .A(n20690), .B(n20691), .Z(n20688) );
  NANDN U20697 ( .A(n6070), .B(n6673), .Z(n20691) );
  NANDN U20698 ( .A(n6084), .B(n20166), .Z(n20690) );
  AND U20699 ( .A(n20692), .B(n20693), .Z(n6091) );
  NANDN U20700 ( .A(n6070), .B(n20166), .Z(n20693) );
  NANDN U20701 ( .A(n6070), .B(n20167), .Z(n20692) );
  IV U20702 ( .A(\stack[0][38] ), .Z(n6070) );
  IV U20703 ( .A(n20264), .Z(n6112) );
  XOR U20704 ( .A(n20168), .B(n20694), .Z(n20264) );
  NAND U20705 ( .A(n20695), .B(n20696), .Z(n20694) );
  NANDN U20706 ( .A(n6108), .B(n20167), .Z(n20696) );
  AND U20707 ( .A(n20697), .B(n20698), .Z(n20695) );
  NANDN U20708 ( .A(n6094), .B(n6673), .Z(n20698) );
  NANDN U20709 ( .A(n6108), .B(n20166), .Z(n20697) );
  AND U20710 ( .A(n20699), .B(n20700), .Z(n6115) );
  NANDN U20711 ( .A(n6094), .B(n20166), .Z(n20700) );
  NANDN U20712 ( .A(n6094), .B(n20167), .Z(n20699) );
  IV U20713 ( .A(\stack[0][39] ), .Z(n6094) );
  IV U20714 ( .A(n20260), .Z(n6136) );
  XOR U20715 ( .A(n20168), .B(n20701), .Z(n20260) );
  NAND U20716 ( .A(n20702), .B(n20703), .Z(n20701) );
  NANDN U20717 ( .A(n6132), .B(n20167), .Z(n20703) );
  AND U20718 ( .A(n20704), .B(n20705), .Z(n20702) );
  NANDN U20719 ( .A(n6118), .B(n6673), .Z(n20705) );
  NANDN U20720 ( .A(n6132), .B(n20166), .Z(n20704) );
  AND U20721 ( .A(n20706), .B(n20707), .Z(n6139) );
  NANDN U20722 ( .A(n6118), .B(n20166), .Z(n20707) );
  NANDN U20723 ( .A(n6118), .B(n20167), .Z(n20706) );
  IV U20724 ( .A(\stack[0][40] ), .Z(n6118) );
  IV U20725 ( .A(n20256), .Z(n6160) );
  XOR U20726 ( .A(n20168), .B(n20708), .Z(n20256) );
  NAND U20727 ( .A(n20709), .B(n20710), .Z(n20708) );
  NANDN U20728 ( .A(n6156), .B(n20167), .Z(n20710) );
  AND U20729 ( .A(n20711), .B(n20712), .Z(n20709) );
  NANDN U20730 ( .A(n6142), .B(n6673), .Z(n20712) );
  NANDN U20731 ( .A(n6156), .B(n20166), .Z(n20711) );
  AND U20732 ( .A(n20713), .B(n20714), .Z(n6163) );
  NANDN U20733 ( .A(n6142), .B(n20166), .Z(n20714) );
  NANDN U20734 ( .A(n6142), .B(n20167), .Z(n20713) );
  IV U20735 ( .A(\stack[0][41] ), .Z(n6142) );
  IV U20736 ( .A(n20252), .Z(n6184) );
  XOR U20737 ( .A(n20168), .B(n20715), .Z(n20252) );
  NAND U20738 ( .A(n20716), .B(n20717), .Z(n20715) );
  NANDN U20739 ( .A(n6180), .B(n20167), .Z(n20717) );
  AND U20740 ( .A(n20718), .B(n20719), .Z(n20716) );
  NANDN U20741 ( .A(n6166), .B(n6673), .Z(n20719) );
  NANDN U20742 ( .A(n6180), .B(n20166), .Z(n20718) );
  AND U20743 ( .A(n20720), .B(n20721), .Z(n6187) );
  NANDN U20744 ( .A(n6166), .B(n20166), .Z(n20721) );
  NANDN U20745 ( .A(n6166), .B(n20167), .Z(n20720) );
  IV U20746 ( .A(\stack[0][42] ), .Z(n6166) );
  IV U20747 ( .A(n20248), .Z(n6208) );
  XOR U20748 ( .A(n20168), .B(n20722), .Z(n20248) );
  NAND U20749 ( .A(n20723), .B(n20724), .Z(n20722) );
  NANDN U20750 ( .A(n6204), .B(n20167), .Z(n20724) );
  AND U20751 ( .A(n20725), .B(n20726), .Z(n20723) );
  NANDN U20752 ( .A(n6190), .B(n6673), .Z(n20726) );
  NANDN U20753 ( .A(n6204), .B(n20166), .Z(n20725) );
  AND U20754 ( .A(n20727), .B(n20728), .Z(n6211) );
  NANDN U20755 ( .A(n6190), .B(n20166), .Z(n20728) );
  NANDN U20756 ( .A(n6190), .B(n20167), .Z(n20727) );
  IV U20757 ( .A(\stack[0][43] ), .Z(n6190) );
  IV U20758 ( .A(n20244), .Z(n6232) );
  XOR U20759 ( .A(n20168), .B(n20729), .Z(n20244) );
  NAND U20760 ( .A(n20730), .B(n20731), .Z(n20729) );
  NANDN U20761 ( .A(n6228), .B(n20167), .Z(n20731) );
  AND U20762 ( .A(n20732), .B(n20733), .Z(n20730) );
  NANDN U20763 ( .A(n6214), .B(n6673), .Z(n20733) );
  NANDN U20764 ( .A(n6228), .B(n20166), .Z(n20732) );
  AND U20765 ( .A(n20734), .B(n20735), .Z(n6235) );
  NANDN U20766 ( .A(n6214), .B(n20166), .Z(n20735) );
  NANDN U20767 ( .A(n6214), .B(n20167), .Z(n20734) );
  IV U20768 ( .A(\stack[0][44] ), .Z(n6214) );
  IV U20769 ( .A(n20240), .Z(n6256) );
  XOR U20770 ( .A(n20168), .B(n20736), .Z(n20240) );
  NAND U20771 ( .A(n20737), .B(n20738), .Z(n20736) );
  NANDN U20772 ( .A(n6252), .B(n20167), .Z(n20738) );
  AND U20773 ( .A(n20739), .B(n20740), .Z(n20737) );
  NANDN U20774 ( .A(n6238), .B(n6673), .Z(n20740) );
  NANDN U20775 ( .A(n6252), .B(n20166), .Z(n20739) );
  AND U20776 ( .A(n20741), .B(n20742), .Z(n6259) );
  NANDN U20777 ( .A(n6238), .B(n20166), .Z(n20742) );
  NANDN U20778 ( .A(n6238), .B(n20167), .Z(n20741) );
  IV U20779 ( .A(\stack[0][45] ), .Z(n6238) );
  IV U20780 ( .A(n20236), .Z(n6280) );
  XOR U20781 ( .A(n20168), .B(n20743), .Z(n20236) );
  NAND U20782 ( .A(n20744), .B(n20745), .Z(n20743) );
  NANDN U20783 ( .A(n6276), .B(n20167), .Z(n20745) );
  AND U20784 ( .A(n20746), .B(n20747), .Z(n20744) );
  NANDN U20785 ( .A(n6262), .B(n6673), .Z(n20747) );
  NANDN U20786 ( .A(n6276), .B(n20166), .Z(n20746) );
  AND U20787 ( .A(n20748), .B(n20749), .Z(n6283) );
  NANDN U20788 ( .A(n6262), .B(n20166), .Z(n20749) );
  NANDN U20789 ( .A(n6262), .B(n20167), .Z(n20748) );
  IV U20790 ( .A(\stack[0][46] ), .Z(n6262) );
  IV U20791 ( .A(n20232), .Z(n6304) );
  XOR U20792 ( .A(n20168), .B(n20750), .Z(n20232) );
  NAND U20793 ( .A(n20751), .B(n20752), .Z(n20750) );
  NANDN U20794 ( .A(n6300), .B(n20167), .Z(n20752) );
  AND U20795 ( .A(n20753), .B(n20754), .Z(n20751) );
  NANDN U20796 ( .A(n6286), .B(n6673), .Z(n20754) );
  NANDN U20797 ( .A(n6300), .B(n20166), .Z(n20753) );
  AND U20798 ( .A(n20755), .B(n20756), .Z(n6307) );
  NANDN U20799 ( .A(n6286), .B(n20166), .Z(n20756) );
  NANDN U20800 ( .A(n6286), .B(n20167), .Z(n20755) );
  IV U20801 ( .A(\stack[0][47] ), .Z(n6286) );
  IV U20802 ( .A(n20228), .Z(n6328) );
  XOR U20803 ( .A(n20168), .B(n20757), .Z(n20228) );
  NAND U20804 ( .A(n20758), .B(n20759), .Z(n20757) );
  NANDN U20805 ( .A(n6324), .B(n20167), .Z(n20759) );
  AND U20806 ( .A(n20760), .B(n20761), .Z(n20758) );
  NANDN U20807 ( .A(n6310), .B(n6673), .Z(n20761) );
  NANDN U20808 ( .A(n6324), .B(n20166), .Z(n20760) );
  AND U20809 ( .A(n20762), .B(n20763), .Z(n6331) );
  NANDN U20810 ( .A(n6310), .B(n20166), .Z(n20763) );
  NANDN U20811 ( .A(n6310), .B(n20167), .Z(n20762) );
  IV U20812 ( .A(\stack[0][48] ), .Z(n6310) );
  IV U20813 ( .A(n20224), .Z(n6352) );
  XOR U20814 ( .A(n20168), .B(n20764), .Z(n20224) );
  NAND U20815 ( .A(n20765), .B(n20766), .Z(n20764) );
  NANDN U20816 ( .A(n6348), .B(n20167), .Z(n20766) );
  AND U20817 ( .A(n20767), .B(n20768), .Z(n20765) );
  NANDN U20818 ( .A(n6334), .B(n6673), .Z(n20768) );
  NANDN U20819 ( .A(n6348), .B(n20166), .Z(n20767) );
  AND U20820 ( .A(n20769), .B(n20770), .Z(n6355) );
  NANDN U20821 ( .A(n6334), .B(n20166), .Z(n20770) );
  NANDN U20822 ( .A(n6334), .B(n20167), .Z(n20769) );
  IV U20823 ( .A(\stack[0][49] ), .Z(n6334) );
  IV U20824 ( .A(n20220), .Z(n6376) );
  XOR U20825 ( .A(n20168), .B(n20771), .Z(n20220) );
  NAND U20826 ( .A(n20772), .B(n20773), .Z(n20771) );
  NANDN U20827 ( .A(n6372), .B(n20167), .Z(n20773) );
  AND U20828 ( .A(n20774), .B(n20775), .Z(n20772) );
  NANDN U20829 ( .A(n6358), .B(n6673), .Z(n20775) );
  NANDN U20830 ( .A(n6372), .B(n20166), .Z(n20774) );
  AND U20831 ( .A(n20776), .B(n20777), .Z(n6379) );
  NANDN U20832 ( .A(n6358), .B(n20166), .Z(n20777) );
  NANDN U20833 ( .A(n6358), .B(n20167), .Z(n20776) );
  IV U20834 ( .A(\stack[0][50] ), .Z(n6358) );
  IV U20835 ( .A(n20216), .Z(n6400) );
  XOR U20836 ( .A(n20168), .B(n20778), .Z(n20216) );
  NAND U20837 ( .A(n20779), .B(n20780), .Z(n20778) );
  NANDN U20838 ( .A(n6396), .B(n20167), .Z(n20780) );
  AND U20839 ( .A(n20781), .B(n20782), .Z(n20779) );
  NANDN U20840 ( .A(n6382), .B(n6673), .Z(n20782) );
  NANDN U20841 ( .A(n6396), .B(n20166), .Z(n20781) );
  AND U20842 ( .A(n20783), .B(n20784), .Z(n6403) );
  NANDN U20843 ( .A(n6382), .B(n20166), .Z(n20784) );
  NANDN U20844 ( .A(n6382), .B(n20167), .Z(n20783) );
  IV U20845 ( .A(\stack[0][51] ), .Z(n6382) );
  IV U20846 ( .A(n20212), .Z(n6424) );
  XOR U20847 ( .A(n20168), .B(n20785), .Z(n20212) );
  NAND U20848 ( .A(n20786), .B(n20787), .Z(n20785) );
  NANDN U20849 ( .A(n6420), .B(n20167), .Z(n20787) );
  AND U20850 ( .A(n20788), .B(n20789), .Z(n20786) );
  NANDN U20851 ( .A(n6406), .B(n6673), .Z(n20789) );
  NANDN U20852 ( .A(n6420), .B(n20166), .Z(n20788) );
  AND U20853 ( .A(n20790), .B(n20791), .Z(n6427) );
  NANDN U20854 ( .A(n6406), .B(n20166), .Z(n20791) );
  NANDN U20855 ( .A(n6406), .B(n20167), .Z(n20790) );
  IV U20856 ( .A(\stack[0][52] ), .Z(n6406) );
  IV U20857 ( .A(n20208), .Z(n6448) );
  XOR U20858 ( .A(n20168), .B(n20792), .Z(n20208) );
  NAND U20859 ( .A(n20793), .B(n20794), .Z(n20792) );
  NANDN U20860 ( .A(n6444), .B(n20167), .Z(n20794) );
  AND U20861 ( .A(n20795), .B(n20796), .Z(n20793) );
  NANDN U20862 ( .A(n6430), .B(n6673), .Z(n20796) );
  NANDN U20863 ( .A(n6444), .B(n20166), .Z(n20795) );
  AND U20864 ( .A(n20797), .B(n20798), .Z(n6451) );
  NANDN U20865 ( .A(n6430), .B(n20166), .Z(n20798) );
  NANDN U20866 ( .A(n6430), .B(n20167), .Z(n20797) );
  IV U20867 ( .A(\stack[0][53] ), .Z(n6430) );
  IV U20868 ( .A(n20204), .Z(n6472) );
  XOR U20869 ( .A(n20168), .B(n20799), .Z(n20204) );
  NAND U20870 ( .A(n20800), .B(n20801), .Z(n20799) );
  NANDN U20871 ( .A(n6468), .B(n20167), .Z(n20801) );
  AND U20872 ( .A(n20802), .B(n20803), .Z(n20800) );
  NANDN U20873 ( .A(n6454), .B(n6673), .Z(n20803) );
  NANDN U20874 ( .A(n6468), .B(n20166), .Z(n20802) );
  AND U20875 ( .A(n20804), .B(n20805), .Z(n6475) );
  NANDN U20876 ( .A(n6454), .B(n20166), .Z(n20805) );
  NANDN U20877 ( .A(n6454), .B(n20167), .Z(n20804) );
  IV U20878 ( .A(\stack[0][54] ), .Z(n6454) );
  IV U20879 ( .A(n20200), .Z(n6496) );
  XOR U20880 ( .A(n20168), .B(n20806), .Z(n20200) );
  NAND U20881 ( .A(n20807), .B(n20808), .Z(n20806) );
  NANDN U20882 ( .A(n6492), .B(n20167), .Z(n20808) );
  AND U20883 ( .A(n20809), .B(n20810), .Z(n20807) );
  NANDN U20884 ( .A(n6478), .B(n6673), .Z(n20810) );
  NANDN U20885 ( .A(n6492), .B(n20166), .Z(n20809) );
  AND U20886 ( .A(n20811), .B(n20812), .Z(n6499) );
  NANDN U20887 ( .A(n6478), .B(n20166), .Z(n20812) );
  NANDN U20888 ( .A(n6478), .B(n20167), .Z(n20811) );
  IV U20889 ( .A(\stack[0][55] ), .Z(n6478) );
  IV U20890 ( .A(n20196), .Z(n6520) );
  XOR U20891 ( .A(n20168), .B(n20813), .Z(n20196) );
  NAND U20892 ( .A(n20814), .B(n20815), .Z(n20813) );
  NANDN U20893 ( .A(n6516), .B(n20167), .Z(n20815) );
  AND U20894 ( .A(n20816), .B(n20817), .Z(n20814) );
  NANDN U20895 ( .A(n6502), .B(n6673), .Z(n20817) );
  NANDN U20896 ( .A(n6516), .B(n20166), .Z(n20816) );
  AND U20897 ( .A(n20818), .B(n20819), .Z(n6523) );
  NANDN U20898 ( .A(n6502), .B(n20166), .Z(n20819) );
  NANDN U20899 ( .A(n6502), .B(n20167), .Z(n20818) );
  IV U20900 ( .A(\stack[0][56] ), .Z(n6502) );
  IV U20901 ( .A(n20192), .Z(n6544) );
  XOR U20902 ( .A(n20168), .B(n20820), .Z(n20192) );
  NAND U20903 ( .A(n20821), .B(n20822), .Z(n20820) );
  NANDN U20904 ( .A(n6540), .B(n20167), .Z(n20822) );
  AND U20905 ( .A(n20823), .B(n20824), .Z(n20821) );
  NANDN U20906 ( .A(n6526), .B(n6673), .Z(n20824) );
  NANDN U20907 ( .A(n6540), .B(n20166), .Z(n20823) );
  AND U20908 ( .A(n20825), .B(n20826), .Z(n6547) );
  NANDN U20909 ( .A(n6526), .B(n20166), .Z(n20826) );
  NANDN U20910 ( .A(n6526), .B(n20167), .Z(n20825) );
  IV U20911 ( .A(\stack[0][57] ), .Z(n6526) );
  IV U20912 ( .A(n20188), .Z(n6568) );
  XOR U20913 ( .A(n20168), .B(n20827), .Z(n20188) );
  NAND U20914 ( .A(n20828), .B(n20829), .Z(n20827) );
  NANDN U20915 ( .A(n6564), .B(n20167), .Z(n20829) );
  AND U20916 ( .A(n20830), .B(n20831), .Z(n20828) );
  NANDN U20917 ( .A(n6550), .B(n6673), .Z(n20831) );
  NANDN U20918 ( .A(n6564), .B(n20166), .Z(n20830) );
  AND U20919 ( .A(n20832), .B(n20833), .Z(n6571) );
  NANDN U20920 ( .A(n6550), .B(n20166), .Z(n20833) );
  NANDN U20921 ( .A(n6550), .B(n20167), .Z(n20832) );
  IV U20922 ( .A(\stack[0][58] ), .Z(n6550) );
  IV U20923 ( .A(n20184), .Z(n6592) );
  XOR U20924 ( .A(n20168), .B(n20834), .Z(n20184) );
  NAND U20925 ( .A(n20835), .B(n20836), .Z(n20834) );
  NANDN U20926 ( .A(n6588), .B(n20167), .Z(n20836) );
  AND U20927 ( .A(n20837), .B(n20838), .Z(n20835) );
  NANDN U20928 ( .A(n6574), .B(n6673), .Z(n20838) );
  NANDN U20929 ( .A(n6588), .B(n20166), .Z(n20837) );
  AND U20930 ( .A(n20839), .B(n20840), .Z(n6595) );
  NANDN U20931 ( .A(n6574), .B(n20166), .Z(n20840) );
  NANDN U20932 ( .A(n6574), .B(n20167), .Z(n20839) );
  IV U20933 ( .A(\stack[0][59] ), .Z(n6574) );
  IV U20934 ( .A(n20180), .Z(n6616) );
  XOR U20935 ( .A(n20168), .B(n20841), .Z(n20180) );
  NAND U20936 ( .A(n20842), .B(n20843), .Z(n20841) );
  NANDN U20937 ( .A(n6612), .B(n20167), .Z(n20843) );
  AND U20938 ( .A(n20844), .B(n20845), .Z(n20842) );
  NANDN U20939 ( .A(n6598), .B(n6673), .Z(n20845) );
  NANDN U20940 ( .A(n6612), .B(n20166), .Z(n20844) );
  AND U20941 ( .A(n20846), .B(n20847), .Z(n6619) );
  NANDN U20942 ( .A(n6598), .B(n20166), .Z(n20847) );
  NANDN U20943 ( .A(n6598), .B(n20167), .Z(n20846) );
  IV U20944 ( .A(\stack[0][60] ), .Z(n6598) );
  IV U20945 ( .A(n20176), .Z(n6640) );
  XOR U20946 ( .A(n20168), .B(n20848), .Z(n20176) );
  NAND U20947 ( .A(n20849), .B(n20850), .Z(n20848) );
  NANDN U20948 ( .A(n6636), .B(n20167), .Z(n20850) );
  AND U20949 ( .A(n20851), .B(n20852), .Z(n20849) );
  NANDN U20950 ( .A(n6622), .B(n6673), .Z(n20852) );
  NANDN U20951 ( .A(n6636), .B(n20166), .Z(n20851) );
  IV U20952 ( .A(n5181), .Z(n20168) );
  AND U20953 ( .A(n20853), .B(n20854), .Z(n6643) );
  NANDN U20954 ( .A(n6622), .B(n20166), .Z(n20854) );
  NANDN U20955 ( .A(n6622), .B(n20167), .Z(n20853) );
  IV U20956 ( .A(\stack[0][61] ), .Z(n6622) );
  AND U20957 ( .A(n20855), .B(n20856), .Z(n20159) );
  NANDN U20958 ( .A(n6670), .B(n20166), .Z(n20856) );
  NANDN U20959 ( .A(n6670), .B(n20167), .Z(n20855) );
  XNOR U20960 ( .A(n5181), .B(n20857), .Z(n20157) );
  AND U20961 ( .A(n20858), .B(n20859), .Z(n20857) );
  NANDN U20962 ( .A(n6684), .B(n20167), .Z(n20859) );
  AND U20963 ( .A(n20860), .B(n20861), .Z(n20858) );
  NANDN U20964 ( .A(n6670), .B(n6673), .Z(n20861) );
  IV U20965 ( .A(\stack[0][63] ), .Z(n6670) );
  NANDN U20966 ( .A(n6684), .B(n20166), .Z(n20860) );
  OR U20967 ( .A(n6673), .B(n20167), .Z(n5181) );
  AND U20968 ( .A(n20862), .B(opcode[0]), .Z(n6673) );
  ANDN U20969 ( .B(n20156), .A(n20863), .Z(n20862) );
  NAND U20970 ( .A(n20864), .B(n20865), .Z(n4899) );
  NANDN U20971 ( .A(n5169), .B(n20866), .Z(n20865) );
  NANDN U20972 ( .A(n20866), .B(n20867), .Z(n20864) );
  NAND U20973 ( .A(n20868), .B(n20869), .Z(n20867) );
  NANDN U20974 ( .A(n4967), .B(\stack[2][0] ), .Z(n20869) );
  NANDN U20975 ( .A(n5160), .B(n4967), .Z(n20868) );
  IV U20976 ( .A(\stack[0][0] ), .Z(n5160) );
  NAND U20977 ( .A(n20870), .B(n20871), .Z(n4898) );
  NANDN U20978 ( .A(n5195), .B(n20866), .Z(n20871) );
  NANDN U20979 ( .A(n20866), .B(n20872), .Z(n20870) );
  NAND U20980 ( .A(n20873), .B(n20874), .Z(n20872) );
  NANDN U20981 ( .A(n4967), .B(\stack[2][1] ), .Z(n20874) );
  NANDN U20982 ( .A(n20875), .B(\stack[0][1] ), .Z(n20873) );
  NAND U20983 ( .A(n20876), .B(n20877), .Z(n4897) );
  NANDN U20984 ( .A(n5219), .B(n20866), .Z(n20877) );
  NANDN U20985 ( .A(n20866), .B(n20878), .Z(n20876) );
  NAND U20986 ( .A(n20879), .B(n20880), .Z(n20878) );
  NANDN U20987 ( .A(n4967), .B(\stack[2][2] ), .Z(n20880) );
  NANDN U20988 ( .A(n5206), .B(n4967), .Z(n20879) );
  IV U20989 ( .A(\stack[0][2] ), .Z(n5206) );
  NAND U20990 ( .A(n20881), .B(n20882), .Z(n4896) );
  NANDN U20991 ( .A(n5243), .B(n20866), .Z(n20882) );
  NANDN U20992 ( .A(n20866), .B(n20883), .Z(n20881) );
  NAND U20993 ( .A(n20884), .B(n20885), .Z(n20883) );
  NANDN U20994 ( .A(n4967), .B(\stack[2][3] ), .Z(n20885) );
  NANDN U20995 ( .A(n5230), .B(n4967), .Z(n20884) );
  IV U20996 ( .A(\stack[0][3] ), .Z(n5230) );
  NAND U20997 ( .A(n20886), .B(n20887), .Z(n4895) );
  NANDN U20998 ( .A(n5267), .B(n20866), .Z(n20887) );
  NANDN U20999 ( .A(n20866), .B(n20888), .Z(n20886) );
  NAND U21000 ( .A(n20889), .B(n20890), .Z(n20888) );
  NANDN U21001 ( .A(n4967), .B(\stack[2][4] ), .Z(n20890) );
  NANDN U21002 ( .A(n5254), .B(n4967), .Z(n20889) );
  IV U21003 ( .A(\stack[0][4] ), .Z(n5254) );
  NAND U21004 ( .A(n20891), .B(n20892), .Z(n4894) );
  NANDN U21005 ( .A(n5292), .B(n20866), .Z(n20892) );
  NANDN U21006 ( .A(n20866), .B(n20893), .Z(n20891) );
  NAND U21007 ( .A(n20894), .B(n20895), .Z(n20893) );
  NANDN U21008 ( .A(n4967), .B(\stack[2][5] ), .Z(n20895) );
  NANDN U21009 ( .A(n5278), .B(n4967), .Z(n20894) );
  IV U21010 ( .A(\stack[0][5] ), .Z(n5278) );
  NAND U21011 ( .A(n20896), .B(n20897), .Z(n4893) );
  NANDN U21012 ( .A(n5316), .B(n20866), .Z(n20897) );
  NANDN U21013 ( .A(n20866), .B(n20898), .Z(n20896) );
  NAND U21014 ( .A(n20899), .B(n20900), .Z(n20898) );
  NANDN U21015 ( .A(n4967), .B(\stack[2][6] ), .Z(n20900) );
  NANDN U21016 ( .A(n5302), .B(n4967), .Z(n20899) );
  IV U21017 ( .A(\stack[0][6] ), .Z(n5302) );
  NAND U21018 ( .A(n20901), .B(n20902), .Z(n4892) );
  NANDN U21019 ( .A(n5340), .B(n20866), .Z(n20902) );
  NANDN U21020 ( .A(n20866), .B(n20903), .Z(n20901) );
  NAND U21021 ( .A(n20904), .B(n20905), .Z(n20903) );
  NANDN U21022 ( .A(n4967), .B(\stack[2][7] ), .Z(n20905) );
  NANDN U21023 ( .A(n5326), .B(n4967), .Z(n20904) );
  IV U21024 ( .A(\stack[0][7] ), .Z(n5326) );
  NAND U21025 ( .A(n20906), .B(n20907), .Z(n4891) );
  NANDN U21026 ( .A(n5364), .B(n20866), .Z(n20907) );
  NANDN U21027 ( .A(n20866), .B(n20908), .Z(n20906) );
  NAND U21028 ( .A(n20909), .B(n20910), .Z(n20908) );
  NANDN U21029 ( .A(n4967), .B(\stack[2][8] ), .Z(n20910) );
  NANDN U21030 ( .A(n5350), .B(n4967), .Z(n20909) );
  IV U21031 ( .A(\stack[0][8] ), .Z(n5350) );
  NAND U21032 ( .A(n20911), .B(n20912), .Z(n4890) );
  NANDN U21033 ( .A(n5387), .B(n20866), .Z(n20912) );
  NANDN U21034 ( .A(n20866), .B(n20913), .Z(n20911) );
  NAND U21035 ( .A(n20914), .B(n20915), .Z(n20913) );
  NANDN U21036 ( .A(n4967), .B(\stack[2][9] ), .Z(n20915) );
  NANDN U21037 ( .A(n5374), .B(n4967), .Z(n20914) );
  IV U21038 ( .A(\stack[0][9] ), .Z(n5374) );
  NAND U21039 ( .A(n20916), .B(n20917), .Z(n4889) );
  NANDN U21040 ( .A(n5411), .B(n20866), .Z(n20917) );
  IV U21041 ( .A(\stack[1][10] ), .Z(n5411) );
  NANDN U21042 ( .A(n20866), .B(n20918), .Z(n20916) );
  NAND U21043 ( .A(n20919), .B(n20920), .Z(n20918) );
  NANDN U21044 ( .A(n4967), .B(\stack[2][10] ), .Z(n20920) );
  NANDN U21045 ( .A(n20875), .B(\stack[0][10] ), .Z(n20919) );
  NAND U21046 ( .A(n20921), .B(n20922), .Z(n4888) );
  NANDN U21047 ( .A(n5435), .B(n20866), .Z(n20922) );
  IV U21048 ( .A(\stack[1][11] ), .Z(n5435) );
  NANDN U21049 ( .A(n20866), .B(n20923), .Z(n20921) );
  NAND U21050 ( .A(n20924), .B(n20925), .Z(n20923) );
  NANDN U21051 ( .A(n4967), .B(\stack[2][11] ), .Z(n20925) );
  NANDN U21052 ( .A(n20875), .B(\stack[0][11] ), .Z(n20924) );
  NAND U21053 ( .A(n20926), .B(n20927), .Z(n4887) );
  NANDN U21054 ( .A(n5459), .B(n20866), .Z(n20927) );
  IV U21055 ( .A(\stack[1][12] ), .Z(n5459) );
  NANDN U21056 ( .A(n20866), .B(n20928), .Z(n20926) );
  NAND U21057 ( .A(n20929), .B(n20930), .Z(n20928) );
  NANDN U21058 ( .A(n4967), .B(\stack[2][12] ), .Z(n20930) );
  NANDN U21059 ( .A(n20875), .B(\stack[0][12] ), .Z(n20929) );
  NAND U21060 ( .A(n20931), .B(n20932), .Z(n4886) );
  NANDN U21061 ( .A(n5483), .B(n20866), .Z(n20932) );
  IV U21062 ( .A(\stack[1][13] ), .Z(n5483) );
  NANDN U21063 ( .A(n20866), .B(n20933), .Z(n20931) );
  NAND U21064 ( .A(n20934), .B(n20935), .Z(n20933) );
  NANDN U21065 ( .A(n4967), .B(\stack[2][13] ), .Z(n20935) );
  NANDN U21066 ( .A(n20875), .B(\stack[0][13] ), .Z(n20934) );
  NAND U21067 ( .A(n20936), .B(n20937), .Z(n4885) );
  NANDN U21068 ( .A(n5507), .B(n20866), .Z(n20937) );
  IV U21069 ( .A(\stack[1][14] ), .Z(n5507) );
  NANDN U21070 ( .A(n20866), .B(n20938), .Z(n20936) );
  NAND U21071 ( .A(n20939), .B(n20940), .Z(n20938) );
  NANDN U21072 ( .A(n4967), .B(\stack[2][14] ), .Z(n20940) );
  NANDN U21073 ( .A(n20875), .B(\stack[0][14] ), .Z(n20939) );
  NAND U21074 ( .A(n20941), .B(n20942), .Z(n4884) );
  NANDN U21075 ( .A(n5531), .B(n20866), .Z(n20942) );
  IV U21076 ( .A(\stack[1][15] ), .Z(n5531) );
  NANDN U21077 ( .A(n20866), .B(n20943), .Z(n20941) );
  NAND U21078 ( .A(n20944), .B(n20945), .Z(n20943) );
  NANDN U21079 ( .A(n4967), .B(\stack[2][15] ), .Z(n20945) );
  NANDN U21080 ( .A(n20875), .B(\stack[0][15] ), .Z(n20944) );
  NAND U21081 ( .A(n20946), .B(n20947), .Z(n4883) );
  NANDN U21082 ( .A(n5555), .B(n20866), .Z(n20947) );
  IV U21083 ( .A(\stack[1][16] ), .Z(n5555) );
  NANDN U21084 ( .A(n20866), .B(n20948), .Z(n20946) );
  NAND U21085 ( .A(n20949), .B(n20950), .Z(n20948) );
  NANDN U21086 ( .A(n4967), .B(\stack[2][16] ), .Z(n20950) );
  NANDN U21087 ( .A(n20875), .B(\stack[0][16] ), .Z(n20949) );
  NAND U21088 ( .A(n20951), .B(n20952), .Z(n4882) );
  NANDN U21089 ( .A(n5579), .B(n20866), .Z(n20952) );
  IV U21090 ( .A(\stack[1][17] ), .Z(n5579) );
  NANDN U21091 ( .A(n20866), .B(n20953), .Z(n20951) );
  NAND U21092 ( .A(n20954), .B(n20955), .Z(n20953) );
  NANDN U21093 ( .A(n4967), .B(\stack[2][17] ), .Z(n20955) );
  NANDN U21094 ( .A(n20875), .B(\stack[0][17] ), .Z(n20954) );
  NAND U21095 ( .A(n20956), .B(n20957), .Z(n4881) );
  NANDN U21096 ( .A(n5603), .B(n20866), .Z(n20957) );
  IV U21097 ( .A(\stack[1][18] ), .Z(n5603) );
  NANDN U21098 ( .A(n20866), .B(n20958), .Z(n20956) );
  NAND U21099 ( .A(n20959), .B(n20960), .Z(n20958) );
  NANDN U21100 ( .A(n4967), .B(\stack[2][18] ), .Z(n20960) );
  NANDN U21101 ( .A(n20875), .B(\stack[0][18] ), .Z(n20959) );
  NAND U21102 ( .A(n20961), .B(n20962), .Z(n4880) );
  NANDN U21103 ( .A(n5627), .B(n20866), .Z(n20962) );
  IV U21104 ( .A(\stack[1][19] ), .Z(n5627) );
  NANDN U21105 ( .A(n20866), .B(n20963), .Z(n20961) );
  NAND U21106 ( .A(n20964), .B(n20965), .Z(n20963) );
  NANDN U21107 ( .A(n4967), .B(\stack[2][19] ), .Z(n20965) );
  NANDN U21108 ( .A(n20875), .B(\stack[0][19] ), .Z(n20964) );
  NAND U21109 ( .A(n20966), .B(n20967), .Z(n4879) );
  NANDN U21110 ( .A(n5651), .B(n20866), .Z(n20967) );
  IV U21111 ( .A(\stack[1][20] ), .Z(n5651) );
  NANDN U21112 ( .A(n20866), .B(n20968), .Z(n20966) );
  NAND U21113 ( .A(n20969), .B(n20970), .Z(n20968) );
  NANDN U21114 ( .A(n4967), .B(\stack[2][20] ), .Z(n20970) );
  NANDN U21115 ( .A(n20875), .B(\stack[0][20] ), .Z(n20969) );
  NAND U21116 ( .A(n20971), .B(n20972), .Z(n4878) );
  NANDN U21117 ( .A(n5675), .B(n20866), .Z(n20972) );
  IV U21118 ( .A(\stack[1][21] ), .Z(n5675) );
  NANDN U21119 ( .A(n20866), .B(n20973), .Z(n20971) );
  NAND U21120 ( .A(n20974), .B(n20975), .Z(n20973) );
  NANDN U21121 ( .A(n4967), .B(\stack[2][21] ), .Z(n20975) );
  NANDN U21122 ( .A(n20875), .B(\stack[0][21] ), .Z(n20974) );
  NAND U21123 ( .A(n20976), .B(n20977), .Z(n4877) );
  NANDN U21124 ( .A(n5699), .B(n20866), .Z(n20977) );
  IV U21125 ( .A(\stack[1][22] ), .Z(n5699) );
  NANDN U21126 ( .A(n20866), .B(n20978), .Z(n20976) );
  NAND U21127 ( .A(n20979), .B(n20980), .Z(n20978) );
  NANDN U21128 ( .A(n4967), .B(\stack[2][22] ), .Z(n20980) );
  NANDN U21129 ( .A(n20875), .B(\stack[0][22] ), .Z(n20979) );
  NAND U21130 ( .A(n20981), .B(n20982), .Z(n4876) );
  NANDN U21131 ( .A(n5723), .B(n20866), .Z(n20982) );
  IV U21132 ( .A(\stack[1][23] ), .Z(n5723) );
  NANDN U21133 ( .A(n20866), .B(n20983), .Z(n20981) );
  NAND U21134 ( .A(n20984), .B(n20985), .Z(n20983) );
  NANDN U21135 ( .A(n4967), .B(\stack[2][23] ), .Z(n20985) );
  NANDN U21136 ( .A(n20875), .B(\stack[0][23] ), .Z(n20984) );
  NAND U21137 ( .A(n20986), .B(n20987), .Z(n4875) );
  NANDN U21138 ( .A(n5747), .B(n20866), .Z(n20987) );
  IV U21139 ( .A(\stack[1][24] ), .Z(n5747) );
  NANDN U21140 ( .A(n20866), .B(n20988), .Z(n20986) );
  NAND U21141 ( .A(n20989), .B(n20990), .Z(n20988) );
  NANDN U21142 ( .A(n4967), .B(\stack[2][24] ), .Z(n20990) );
  NANDN U21143 ( .A(n20875), .B(\stack[0][24] ), .Z(n20989) );
  NAND U21144 ( .A(n20991), .B(n20992), .Z(n4874) );
  NANDN U21145 ( .A(n5771), .B(n20866), .Z(n20992) );
  IV U21146 ( .A(\stack[1][25] ), .Z(n5771) );
  NANDN U21147 ( .A(n20866), .B(n20993), .Z(n20991) );
  NAND U21148 ( .A(n20994), .B(n20995), .Z(n20993) );
  NANDN U21149 ( .A(n4967), .B(\stack[2][25] ), .Z(n20995) );
  NANDN U21150 ( .A(n20875), .B(\stack[0][25] ), .Z(n20994) );
  NAND U21151 ( .A(n20996), .B(n20997), .Z(n4873) );
  NANDN U21152 ( .A(n5795), .B(n20866), .Z(n20997) );
  IV U21153 ( .A(\stack[1][26] ), .Z(n5795) );
  NANDN U21154 ( .A(n20866), .B(n20998), .Z(n20996) );
  NAND U21155 ( .A(n20999), .B(n21000), .Z(n20998) );
  NANDN U21156 ( .A(n4967), .B(\stack[2][26] ), .Z(n21000) );
  NANDN U21157 ( .A(n20875), .B(\stack[0][26] ), .Z(n20999) );
  NAND U21158 ( .A(n21001), .B(n21002), .Z(n4872) );
  NANDN U21159 ( .A(n5819), .B(n20866), .Z(n21002) );
  IV U21160 ( .A(\stack[1][27] ), .Z(n5819) );
  NANDN U21161 ( .A(n20866), .B(n21003), .Z(n21001) );
  NAND U21162 ( .A(n21004), .B(n21005), .Z(n21003) );
  NANDN U21163 ( .A(n4967), .B(\stack[2][27] ), .Z(n21005) );
  NANDN U21164 ( .A(n20875), .B(\stack[0][27] ), .Z(n21004) );
  NAND U21165 ( .A(n21006), .B(n21007), .Z(n4871) );
  NANDN U21166 ( .A(n5843), .B(n20866), .Z(n21007) );
  IV U21167 ( .A(\stack[1][28] ), .Z(n5843) );
  NANDN U21168 ( .A(n20866), .B(n21008), .Z(n21006) );
  NAND U21169 ( .A(n21009), .B(n21010), .Z(n21008) );
  NANDN U21170 ( .A(n4967), .B(\stack[2][28] ), .Z(n21010) );
  NANDN U21171 ( .A(n20875), .B(\stack[0][28] ), .Z(n21009) );
  NAND U21172 ( .A(n21011), .B(n21012), .Z(n4870) );
  NANDN U21173 ( .A(n5867), .B(n20866), .Z(n21012) );
  IV U21174 ( .A(\stack[1][29] ), .Z(n5867) );
  NANDN U21175 ( .A(n20866), .B(n21013), .Z(n21011) );
  NAND U21176 ( .A(n21014), .B(n21015), .Z(n21013) );
  NANDN U21177 ( .A(n4967), .B(\stack[2][29] ), .Z(n21015) );
  NANDN U21178 ( .A(n20875), .B(\stack[0][29] ), .Z(n21014) );
  NAND U21179 ( .A(n21016), .B(n21017), .Z(n4869) );
  NANDN U21180 ( .A(n5891), .B(n20866), .Z(n21017) );
  IV U21181 ( .A(\stack[1][30] ), .Z(n5891) );
  NANDN U21182 ( .A(n20866), .B(n21018), .Z(n21016) );
  NAND U21183 ( .A(n21019), .B(n21020), .Z(n21018) );
  NANDN U21184 ( .A(n4967), .B(\stack[2][30] ), .Z(n21020) );
  NANDN U21185 ( .A(n20875), .B(\stack[0][30] ), .Z(n21019) );
  NAND U21186 ( .A(n21021), .B(n21022), .Z(n4868) );
  NANDN U21187 ( .A(n5915), .B(n20866), .Z(n21022) );
  IV U21188 ( .A(\stack[1][31] ), .Z(n5915) );
  NANDN U21189 ( .A(n20866), .B(n21023), .Z(n21021) );
  NAND U21190 ( .A(n21024), .B(n21025), .Z(n21023) );
  NANDN U21191 ( .A(n4967), .B(\stack[2][31] ), .Z(n21025) );
  NANDN U21192 ( .A(n20875), .B(\stack[0][31] ), .Z(n21024) );
  NAND U21193 ( .A(n21026), .B(n21027), .Z(n4867) );
  NANDN U21194 ( .A(n5940), .B(n20866), .Z(n21027) );
  IV U21195 ( .A(\stack[1][32] ), .Z(n5940) );
  NANDN U21196 ( .A(n20866), .B(n21028), .Z(n21026) );
  NAND U21197 ( .A(n21029), .B(n21030), .Z(n21028) );
  NANDN U21198 ( .A(n4967), .B(\stack[2][32] ), .Z(n21030) );
  NANDN U21199 ( .A(n20875), .B(\stack[0][32] ), .Z(n21029) );
  NAND U21200 ( .A(n21031), .B(n21032), .Z(n4866) );
  NANDN U21201 ( .A(n5964), .B(n20866), .Z(n21032) );
  IV U21202 ( .A(\stack[1][33] ), .Z(n5964) );
  NANDN U21203 ( .A(n20866), .B(n21033), .Z(n21031) );
  NAND U21204 ( .A(n21034), .B(n21035), .Z(n21033) );
  NANDN U21205 ( .A(n4967), .B(\stack[2][33] ), .Z(n21035) );
  NANDN U21206 ( .A(n20875), .B(\stack[0][33] ), .Z(n21034) );
  NAND U21207 ( .A(n21036), .B(n21037), .Z(n4865) );
  NANDN U21208 ( .A(n5988), .B(n20866), .Z(n21037) );
  IV U21209 ( .A(\stack[1][34] ), .Z(n5988) );
  NANDN U21210 ( .A(n20866), .B(n21038), .Z(n21036) );
  NAND U21211 ( .A(n21039), .B(n21040), .Z(n21038) );
  NANDN U21212 ( .A(n4967), .B(\stack[2][34] ), .Z(n21040) );
  NANDN U21213 ( .A(n20875), .B(\stack[0][34] ), .Z(n21039) );
  NAND U21214 ( .A(n21041), .B(n21042), .Z(n4864) );
  NANDN U21215 ( .A(n6012), .B(n20866), .Z(n21042) );
  IV U21216 ( .A(\stack[1][35] ), .Z(n6012) );
  NANDN U21217 ( .A(n20866), .B(n21043), .Z(n21041) );
  NAND U21218 ( .A(n21044), .B(n21045), .Z(n21043) );
  NANDN U21219 ( .A(n4967), .B(\stack[2][35] ), .Z(n21045) );
  NANDN U21220 ( .A(n20875), .B(\stack[0][35] ), .Z(n21044) );
  NAND U21221 ( .A(n21046), .B(n21047), .Z(n4863) );
  NANDN U21222 ( .A(n6036), .B(n20866), .Z(n21047) );
  IV U21223 ( .A(\stack[1][36] ), .Z(n6036) );
  NANDN U21224 ( .A(n20866), .B(n21048), .Z(n21046) );
  NAND U21225 ( .A(n21049), .B(n21050), .Z(n21048) );
  NANDN U21226 ( .A(n4967), .B(\stack[2][36] ), .Z(n21050) );
  NANDN U21227 ( .A(n20875), .B(\stack[0][36] ), .Z(n21049) );
  NAND U21228 ( .A(n21051), .B(n21052), .Z(n4862) );
  NANDN U21229 ( .A(n6060), .B(n20866), .Z(n21052) );
  IV U21230 ( .A(\stack[1][37] ), .Z(n6060) );
  NANDN U21231 ( .A(n20866), .B(n21053), .Z(n21051) );
  NAND U21232 ( .A(n21054), .B(n21055), .Z(n21053) );
  NANDN U21233 ( .A(n4967), .B(\stack[2][37] ), .Z(n21055) );
  NANDN U21234 ( .A(n20875), .B(\stack[0][37] ), .Z(n21054) );
  NAND U21235 ( .A(n21056), .B(n21057), .Z(n4861) );
  NANDN U21236 ( .A(n6084), .B(n20866), .Z(n21057) );
  IV U21237 ( .A(\stack[1][38] ), .Z(n6084) );
  NANDN U21238 ( .A(n20866), .B(n21058), .Z(n21056) );
  NAND U21239 ( .A(n21059), .B(n21060), .Z(n21058) );
  NANDN U21240 ( .A(n4967), .B(\stack[2][38] ), .Z(n21060) );
  NANDN U21241 ( .A(n20875), .B(\stack[0][38] ), .Z(n21059) );
  NAND U21242 ( .A(n21061), .B(n21062), .Z(n4860) );
  NANDN U21243 ( .A(n6108), .B(n20866), .Z(n21062) );
  IV U21244 ( .A(\stack[1][39] ), .Z(n6108) );
  NANDN U21245 ( .A(n20866), .B(n21063), .Z(n21061) );
  NAND U21246 ( .A(n21064), .B(n21065), .Z(n21063) );
  NANDN U21247 ( .A(n4967), .B(\stack[2][39] ), .Z(n21065) );
  NANDN U21248 ( .A(n20875), .B(\stack[0][39] ), .Z(n21064) );
  NAND U21249 ( .A(n21066), .B(n21067), .Z(n4859) );
  NANDN U21250 ( .A(n6132), .B(n20866), .Z(n21067) );
  IV U21251 ( .A(\stack[1][40] ), .Z(n6132) );
  NANDN U21252 ( .A(n20866), .B(n21068), .Z(n21066) );
  NAND U21253 ( .A(n21069), .B(n21070), .Z(n21068) );
  NANDN U21254 ( .A(n4967), .B(\stack[2][40] ), .Z(n21070) );
  NANDN U21255 ( .A(n20875), .B(\stack[0][40] ), .Z(n21069) );
  NAND U21256 ( .A(n21071), .B(n21072), .Z(n4858) );
  NANDN U21257 ( .A(n6156), .B(n20866), .Z(n21072) );
  IV U21258 ( .A(\stack[1][41] ), .Z(n6156) );
  NANDN U21259 ( .A(n20866), .B(n21073), .Z(n21071) );
  NAND U21260 ( .A(n21074), .B(n21075), .Z(n21073) );
  NANDN U21261 ( .A(n4967), .B(\stack[2][41] ), .Z(n21075) );
  NANDN U21262 ( .A(n20875), .B(\stack[0][41] ), .Z(n21074) );
  NAND U21263 ( .A(n21076), .B(n21077), .Z(n4857) );
  NANDN U21264 ( .A(n6180), .B(n20866), .Z(n21077) );
  IV U21265 ( .A(\stack[1][42] ), .Z(n6180) );
  NANDN U21266 ( .A(n20866), .B(n21078), .Z(n21076) );
  NAND U21267 ( .A(n21079), .B(n21080), .Z(n21078) );
  NANDN U21268 ( .A(n4967), .B(\stack[2][42] ), .Z(n21080) );
  NANDN U21269 ( .A(n20875), .B(\stack[0][42] ), .Z(n21079) );
  NAND U21270 ( .A(n21081), .B(n21082), .Z(n4856) );
  NANDN U21271 ( .A(n6204), .B(n20866), .Z(n21082) );
  IV U21272 ( .A(\stack[1][43] ), .Z(n6204) );
  NANDN U21273 ( .A(n20866), .B(n21083), .Z(n21081) );
  NAND U21274 ( .A(n21084), .B(n21085), .Z(n21083) );
  NANDN U21275 ( .A(n4967), .B(\stack[2][43] ), .Z(n21085) );
  NANDN U21276 ( .A(n20875), .B(\stack[0][43] ), .Z(n21084) );
  NAND U21277 ( .A(n21086), .B(n21087), .Z(n4855) );
  NANDN U21278 ( .A(n6228), .B(n20866), .Z(n21087) );
  IV U21279 ( .A(\stack[1][44] ), .Z(n6228) );
  NANDN U21280 ( .A(n20866), .B(n21088), .Z(n21086) );
  NAND U21281 ( .A(n21089), .B(n21090), .Z(n21088) );
  NANDN U21282 ( .A(n4967), .B(\stack[2][44] ), .Z(n21090) );
  NANDN U21283 ( .A(n20875), .B(\stack[0][44] ), .Z(n21089) );
  NAND U21284 ( .A(n21091), .B(n21092), .Z(n4854) );
  NANDN U21285 ( .A(n6252), .B(n20866), .Z(n21092) );
  IV U21286 ( .A(\stack[1][45] ), .Z(n6252) );
  NANDN U21287 ( .A(n20866), .B(n21093), .Z(n21091) );
  NAND U21288 ( .A(n21094), .B(n21095), .Z(n21093) );
  NANDN U21289 ( .A(n4967), .B(\stack[2][45] ), .Z(n21095) );
  NANDN U21290 ( .A(n20875), .B(\stack[0][45] ), .Z(n21094) );
  NAND U21291 ( .A(n21096), .B(n21097), .Z(n4853) );
  NANDN U21292 ( .A(n6276), .B(n20866), .Z(n21097) );
  IV U21293 ( .A(\stack[1][46] ), .Z(n6276) );
  NANDN U21294 ( .A(n20866), .B(n21098), .Z(n21096) );
  NAND U21295 ( .A(n21099), .B(n21100), .Z(n21098) );
  NANDN U21296 ( .A(n4967), .B(\stack[2][46] ), .Z(n21100) );
  NANDN U21297 ( .A(n20875), .B(\stack[0][46] ), .Z(n21099) );
  NAND U21298 ( .A(n21101), .B(n21102), .Z(n4852) );
  NANDN U21299 ( .A(n6300), .B(n20866), .Z(n21102) );
  IV U21300 ( .A(\stack[1][47] ), .Z(n6300) );
  NANDN U21301 ( .A(n20866), .B(n21103), .Z(n21101) );
  NAND U21302 ( .A(n21104), .B(n21105), .Z(n21103) );
  NANDN U21303 ( .A(n4967), .B(\stack[2][47] ), .Z(n21105) );
  NANDN U21304 ( .A(n20875), .B(\stack[0][47] ), .Z(n21104) );
  NAND U21305 ( .A(n21106), .B(n21107), .Z(n4851) );
  NANDN U21306 ( .A(n6324), .B(n20866), .Z(n21107) );
  IV U21307 ( .A(\stack[1][48] ), .Z(n6324) );
  NANDN U21308 ( .A(n20866), .B(n21108), .Z(n21106) );
  NAND U21309 ( .A(n21109), .B(n21110), .Z(n21108) );
  NANDN U21310 ( .A(n4967), .B(\stack[2][48] ), .Z(n21110) );
  NANDN U21311 ( .A(n20875), .B(\stack[0][48] ), .Z(n21109) );
  NAND U21312 ( .A(n21111), .B(n21112), .Z(n4850) );
  NANDN U21313 ( .A(n6348), .B(n20866), .Z(n21112) );
  IV U21314 ( .A(\stack[1][49] ), .Z(n6348) );
  NANDN U21315 ( .A(n20866), .B(n21113), .Z(n21111) );
  NAND U21316 ( .A(n21114), .B(n21115), .Z(n21113) );
  NANDN U21317 ( .A(n4967), .B(\stack[2][49] ), .Z(n21115) );
  NANDN U21318 ( .A(n20875), .B(\stack[0][49] ), .Z(n21114) );
  NAND U21319 ( .A(n21116), .B(n21117), .Z(n4849) );
  NANDN U21320 ( .A(n6372), .B(n20866), .Z(n21117) );
  IV U21321 ( .A(\stack[1][50] ), .Z(n6372) );
  NANDN U21322 ( .A(n20866), .B(n21118), .Z(n21116) );
  NAND U21323 ( .A(n21119), .B(n21120), .Z(n21118) );
  NANDN U21324 ( .A(n4967), .B(\stack[2][50] ), .Z(n21120) );
  NANDN U21325 ( .A(n20875), .B(\stack[0][50] ), .Z(n21119) );
  NAND U21326 ( .A(n21121), .B(n21122), .Z(n4848) );
  NANDN U21327 ( .A(n6396), .B(n20866), .Z(n21122) );
  IV U21328 ( .A(\stack[1][51] ), .Z(n6396) );
  NANDN U21329 ( .A(n20866), .B(n21123), .Z(n21121) );
  NAND U21330 ( .A(n21124), .B(n21125), .Z(n21123) );
  NANDN U21331 ( .A(n4967), .B(\stack[2][51] ), .Z(n21125) );
  NANDN U21332 ( .A(n20875), .B(\stack[0][51] ), .Z(n21124) );
  NAND U21333 ( .A(n21126), .B(n21127), .Z(n4847) );
  NANDN U21334 ( .A(n6420), .B(n20866), .Z(n21127) );
  IV U21335 ( .A(\stack[1][52] ), .Z(n6420) );
  NANDN U21336 ( .A(n20866), .B(n21128), .Z(n21126) );
  NAND U21337 ( .A(n21129), .B(n21130), .Z(n21128) );
  NANDN U21338 ( .A(n4967), .B(\stack[2][52] ), .Z(n21130) );
  NANDN U21339 ( .A(n20875), .B(\stack[0][52] ), .Z(n21129) );
  NAND U21340 ( .A(n21131), .B(n21132), .Z(n4846) );
  NANDN U21341 ( .A(n6444), .B(n20866), .Z(n21132) );
  IV U21342 ( .A(\stack[1][53] ), .Z(n6444) );
  NANDN U21343 ( .A(n20866), .B(n21133), .Z(n21131) );
  NAND U21344 ( .A(n21134), .B(n21135), .Z(n21133) );
  NANDN U21345 ( .A(n4967), .B(\stack[2][53] ), .Z(n21135) );
  NANDN U21346 ( .A(n20875), .B(\stack[0][53] ), .Z(n21134) );
  NAND U21347 ( .A(n21136), .B(n21137), .Z(n4845) );
  NANDN U21348 ( .A(n6468), .B(n20866), .Z(n21137) );
  IV U21349 ( .A(\stack[1][54] ), .Z(n6468) );
  NANDN U21350 ( .A(n20866), .B(n21138), .Z(n21136) );
  NAND U21351 ( .A(n21139), .B(n21140), .Z(n21138) );
  NANDN U21352 ( .A(n4967), .B(\stack[2][54] ), .Z(n21140) );
  NANDN U21353 ( .A(n20875), .B(\stack[0][54] ), .Z(n21139) );
  NAND U21354 ( .A(n21141), .B(n21142), .Z(n4844) );
  NANDN U21355 ( .A(n6492), .B(n20866), .Z(n21142) );
  IV U21356 ( .A(\stack[1][55] ), .Z(n6492) );
  NANDN U21357 ( .A(n20866), .B(n21143), .Z(n21141) );
  NAND U21358 ( .A(n21144), .B(n21145), .Z(n21143) );
  NANDN U21359 ( .A(n4967), .B(\stack[2][55] ), .Z(n21145) );
  NANDN U21360 ( .A(n20875), .B(\stack[0][55] ), .Z(n21144) );
  NAND U21361 ( .A(n21146), .B(n21147), .Z(n4843) );
  NANDN U21362 ( .A(n6516), .B(n20866), .Z(n21147) );
  IV U21363 ( .A(\stack[1][56] ), .Z(n6516) );
  NANDN U21364 ( .A(n20866), .B(n21148), .Z(n21146) );
  NAND U21365 ( .A(n21149), .B(n21150), .Z(n21148) );
  NANDN U21366 ( .A(n4967), .B(\stack[2][56] ), .Z(n21150) );
  NANDN U21367 ( .A(n20875), .B(\stack[0][56] ), .Z(n21149) );
  NAND U21368 ( .A(n21151), .B(n21152), .Z(n4842) );
  NANDN U21369 ( .A(n6540), .B(n20866), .Z(n21152) );
  IV U21370 ( .A(\stack[1][57] ), .Z(n6540) );
  NANDN U21371 ( .A(n20866), .B(n21153), .Z(n21151) );
  NAND U21372 ( .A(n21154), .B(n21155), .Z(n21153) );
  NANDN U21373 ( .A(n4967), .B(\stack[2][57] ), .Z(n21155) );
  NANDN U21374 ( .A(n20875), .B(\stack[0][57] ), .Z(n21154) );
  NAND U21375 ( .A(n21156), .B(n21157), .Z(n4841) );
  NANDN U21376 ( .A(n6564), .B(n20866), .Z(n21157) );
  IV U21377 ( .A(\stack[1][58] ), .Z(n6564) );
  NANDN U21378 ( .A(n20866), .B(n21158), .Z(n21156) );
  NAND U21379 ( .A(n21159), .B(n21160), .Z(n21158) );
  NANDN U21380 ( .A(n4967), .B(\stack[2][58] ), .Z(n21160) );
  NANDN U21381 ( .A(n20875), .B(\stack[0][58] ), .Z(n21159) );
  NAND U21382 ( .A(n21161), .B(n21162), .Z(n4840) );
  NANDN U21383 ( .A(n6588), .B(n20866), .Z(n21162) );
  IV U21384 ( .A(\stack[1][59] ), .Z(n6588) );
  NANDN U21385 ( .A(n20866), .B(n21163), .Z(n21161) );
  NAND U21386 ( .A(n21164), .B(n21165), .Z(n21163) );
  NANDN U21387 ( .A(n4967), .B(\stack[2][59] ), .Z(n21165) );
  NANDN U21388 ( .A(n20875), .B(\stack[0][59] ), .Z(n21164) );
  NAND U21389 ( .A(n21166), .B(n21167), .Z(n4839) );
  NANDN U21390 ( .A(n6612), .B(n20866), .Z(n21167) );
  IV U21391 ( .A(\stack[1][60] ), .Z(n6612) );
  NANDN U21392 ( .A(n20866), .B(n21168), .Z(n21166) );
  NAND U21393 ( .A(n21169), .B(n21170), .Z(n21168) );
  NANDN U21394 ( .A(n4967), .B(\stack[2][60] ), .Z(n21170) );
  NANDN U21395 ( .A(n20875), .B(\stack[0][60] ), .Z(n21169) );
  NAND U21396 ( .A(n21171), .B(n21172), .Z(n4838) );
  NANDN U21397 ( .A(n6636), .B(n20866), .Z(n21172) );
  IV U21398 ( .A(\stack[1][61] ), .Z(n6636) );
  NANDN U21399 ( .A(n20866), .B(n21173), .Z(n21171) );
  NAND U21400 ( .A(n21174), .B(n21175), .Z(n21173) );
  NANDN U21401 ( .A(n4967), .B(\stack[2][61] ), .Z(n21175) );
  NANDN U21402 ( .A(n20875), .B(\stack[0][61] ), .Z(n21174) );
  NAND U21403 ( .A(n21176), .B(n21177), .Z(n4837) );
  NANDN U21404 ( .A(n6659), .B(n20866), .Z(n21177) );
  IV U21405 ( .A(\stack[1][62] ), .Z(n6659) );
  NANDN U21406 ( .A(n20866), .B(n21178), .Z(n21176) );
  NAND U21407 ( .A(n21179), .B(n21180), .Z(n21178) );
  NANDN U21408 ( .A(n4967), .B(\stack[2][62] ), .Z(n21180) );
  NANDN U21409 ( .A(n20875), .B(\stack[0][62] ), .Z(n21179) );
  NAND U21410 ( .A(n21181), .B(n21182), .Z(n4836) );
  NANDN U21411 ( .A(n6684), .B(n20866), .Z(n21182) );
  IV U21412 ( .A(\stack[1][63] ), .Z(n6684) );
  NANDN U21413 ( .A(n20866), .B(n21183), .Z(n21181) );
  NAND U21414 ( .A(n21184), .B(n21185), .Z(n21183) );
  NANDN U21415 ( .A(n4967), .B(\stack[2][63] ), .Z(n21185) );
  NANDN U21416 ( .A(n20875), .B(\stack[0][63] ), .Z(n21184) );
  NAND U21417 ( .A(n21186), .B(n21187), .Z(n4835) );
  NANDN U21418 ( .A(n21188), .B(\stack[2][0] ), .Z(n21187) );
  NANDN U21419 ( .A(n20866), .B(n21189), .Z(n21186) );
  NAND U21420 ( .A(n21190), .B(n21191), .Z(n21189) );
  NANDN U21421 ( .A(n4967), .B(\stack[3][0] ), .Z(n21191) );
  NANDN U21422 ( .A(n5169), .B(n4967), .Z(n21190) );
  IV U21423 ( .A(\stack[1][0] ), .Z(n5169) );
  NAND U21424 ( .A(n21192), .B(n21193), .Z(n4834) );
  NANDN U21425 ( .A(n21188), .B(\stack[2][1] ), .Z(n21193) );
  NANDN U21426 ( .A(n20866), .B(n21194), .Z(n21192) );
  NAND U21427 ( .A(n21195), .B(n21196), .Z(n21194) );
  NANDN U21428 ( .A(n4967), .B(\stack[3][1] ), .Z(n21196) );
  NANDN U21429 ( .A(n5195), .B(n4967), .Z(n21195) );
  IV U21430 ( .A(\stack[1][1] ), .Z(n5195) );
  NAND U21431 ( .A(n21197), .B(n21198), .Z(n4833) );
  NANDN U21432 ( .A(n21188), .B(\stack[2][2] ), .Z(n21198) );
  NANDN U21433 ( .A(n20866), .B(n21199), .Z(n21197) );
  NAND U21434 ( .A(n21200), .B(n21201), .Z(n21199) );
  NANDN U21435 ( .A(n4967), .B(\stack[3][2] ), .Z(n21201) );
  NANDN U21436 ( .A(n5219), .B(n4967), .Z(n21200) );
  IV U21437 ( .A(\stack[1][2] ), .Z(n5219) );
  NAND U21438 ( .A(n21202), .B(n21203), .Z(n4832) );
  NANDN U21439 ( .A(n21188), .B(\stack[2][3] ), .Z(n21203) );
  NANDN U21440 ( .A(n20866), .B(n21204), .Z(n21202) );
  NAND U21441 ( .A(n21205), .B(n21206), .Z(n21204) );
  NANDN U21442 ( .A(n4967), .B(\stack[3][3] ), .Z(n21206) );
  NANDN U21443 ( .A(n5243), .B(n4967), .Z(n21205) );
  IV U21444 ( .A(\stack[1][3] ), .Z(n5243) );
  NAND U21445 ( .A(n21207), .B(n21208), .Z(n4831) );
  NANDN U21446 ( .A(n21188), .B(\stack[2][4] ), .Z(n21208) );
  NANDN U21447 ( .A(n20866), .B(n21209), .Z(n21207) );
  NAND U21448 ( .A(n21210), .B(n21211), .Z(n21209) );
  NANDN U21449 ( .A(n4967), .B(\stack[3][4] ), .Z(n21211) );
  NANDN U21450 ( .A(n5267), .B(n4967), .Z(n21210) );
  IV U21451 ( .A(\stack[1][4] ), .Z(n5267) );
  NAND U21452 ( .A(n21212), .B(n21213), .Z(n4830) );
  NANDN U21453 ( .A(n21188), .B(\stack[2][5] ), .Z(n21213) );
  NANDN U21454 ( .A(n20866), .B(n21214), .Z(n21212) );
  NAND U21455 ( .A(n21215), .B(n21216), .Z(n21214) );
  NANDN U21456 ( .A(n4967), .B(\stack[3][5] ), .Z(n21216) );
  NANDN U21457 ( .A(n5292), .B(n4967), .Z(n21215) );
  IV U21458 ( .A(\stack[1][5] ), .Z(n5292) );
  NAND U21459 ( .A(n21217), .B(n21218), .Z(n4829) );
  NANDN U21460 ( .A(n21188), .B(\stack[2][6] ), .Z(n21218) );
  NANDN U21461 ( .A(n20866), .B(n21219), .Z(n21217) );
  NAND U21462 ( .A(n21220), .B(n21221), .Z(n21219) );
  NANDN U21463 ( .A(n4967), .B(\stack[3][6] ), .Z(n21221) );
  NANDN U21464 ( .A(n5316), .B(n4967), .Z(n21220) );
  IV U21465 ( .A(\stack[1][6] ), .Z(n5316) );
  NAND U21466 ( .A(n21222), .B(n21223), .Z(n4828) );
  NANDN U21467 ( .A(n21188), .B(\stack[2][7] ), .Z(n21223) );
  NANDN U21468 ( .A(n20866), .B(n21224), .Z(n21222) );
  NAND U21469 ( .A(n21225), .B(n21226), .Z(n21224) );
  NANDN U21470 ( .A(n4967), .B(\stack[3][7] ), .Z(n21226) );
  NANDN U21471 ( .A(n5340), .B(n4967), .Z(n21225) );
  IV U21472 ( .A(\stack[1][7] ), .Z(n5340) );
  NAND U21473 ( .A(n21227), .B(n21228), .Z(n4827) );
  NANDN U21474 ( .A(n21188), .B(\stack[2][8] ), .Z(n21228) );
  NANDN U21475 ( .A(n20866), .B(n21229), .Z(n21227) );
  NAND U21476 ( .A(n21230), .B(n21231), .Z(n21229) );
  NANDN U21477 ( .A(n4967), .B(\stack[3][8] ), .Z(n21231) );
  NANDN U21478 ( .A(n5364), .B(n4967), .Z(n21230) );
  IV U21479 ( .A(\stack[1][8] ), .Z(n5364) );
  NAND U21480 ( .A(n21232), .B(n21233), .Z(n4826) );
  NANDN U21481 ( .A(n21188), .B(\stack[2][9] ), .Z(n21233) );
  NANDN U21482 ( .A(n20866), .B(n21234), .Z(n21232) );
  NAND U21483 ( .A(n21235), .B(n21236), .Z(n21234) );
  NANDN U21484 ( .A(n4967), .B(\stack[3][9] ), .Z(n21236) );
  NANDN U21485 ( .A(n5387), .B(n4967), .Z(n21235) );
  IV U21486 ( .A(\stack[1][9] ), .Z(n5387) );
  NAND U21487 ( .A(n21237), .B(n21238), .Z(n4825) );
  NANDN U21488 ( .A(n21188), .B(\stack[2][10] ), .Z(n21238) );
  NANDN U21489 ( .A(n20866), .B(n21239), .Z(n21237) );
  NAND U21490 ( .A(n21240), .B(n21241), .Z(n21239) );
  NANDN U21491 ( .A(n4967), .B(\stack[3][10] ), .Z(n21241) );
  NANDN U21492 ( .A(n20875), .B(\stack[1][10] ), .Z(n21240) );
  NAND U21493 ( .A(n21242), .B(n21243), .Z(n4824) );
  NANDN U21494 ( .A(n21188), .B(\stack[2][11] ), .Z(n21243) );
  NANDN U21495 ( .A(n20866), .B(n21244), .Z(n21242) );
  NAND U21496 ( .A(n21245), .B(n21246), .Z(n21244) );
  NANDN U21497 ( .A(n4967), .B(\stack[3][11] ), .Z(n21246) );
  NANDN U21498 ( .A(n20875), .B(\stack[1][11] ), .Z(n21245) );
  NAND U21499 ( .A(n21247), .B(n21248), .Z(n4823) );
  NANDN U21500 ( .A(n21188), .B(\stack[2][12] ), .Z(n21248) );
  NANDN U21501 ( .A(n20866), .B(n21249), .Z(n21247) );
  NAND U21502 ( .A(n21250), .B(n21251), .Z(n21249) );
  NANDN U21503 ( .A(n4967), .B(\stack[3][12] ), .Z(n21251) );
  NANDN U21504 ( .A(n20875), .B(\stack[1][12] ), .Z(n21250) );
  NAND U21505 ( .A(n21252), .B(n21253), .Z(n4822) );
  NANDN U21506 ( .A(n21188), .B(\stack[2][13] ), .Z(n21253) );
  NANDN U21507 ( .A(n20866), .B(n21254), .Z(n21252) );
  NAND U21508 ( .A(n21255), .B(n21256), .Z(n21254) );
  NANDN U21509 ( .A(n4967), .B(\stack[3][13] ), .Z(n21256) );
  NANDN U21510 ( .A(n20875), .B(\stack[1][13] ), .Z(n21255) );
  NAND U21511 ( .A(n21257), .B(n21258), .Z(n4821) );
  NANDN U21512 ( .A(n21188), .B(\stack[2][14] ), .Z(n21258) );
  NANDN U21513 ( .A(n20866), .B(n21259), .Z(n21257) );
  NAND U21514 ( .A(n21260), .B(n21261), .Z(n21259) );
  NANDN U21515 ( .A(n4967), .B(\stack[3][14] ), .Z(n21261) );
  NANDN U21516 ( .A(n20875), .B(\stack[1][14] ), .Z(n21260) );
  NAND U21517 ( .A(n21262), .B(n21263), .Z(n4820) );
  NANDN U21518 ( .A(n21188), .B(\stack[2][15] ), .Z(n21263) );
  NANDN U21519 ( .A(n20866), .B(n21264), .Z(n21262) );
  NAND U21520 ( .A(n21265), .B(n21266), .Z(n21264) );
  NANDN U21521 ( .A(n4967), .B(\stack[3][15] ), .Z(n21266) );
  NANDN U21522 ( .A(n20875), .B(\stack[1][15] ), .Z(n21265) );
  NAND U21523 ( .A(n21267), .B(n21268), .Z(n4819) );
  NANDN U21524 ( .A(n21188), .B(\stack[2][16] ), .Z(n21268) );
  NANDN U21525 ( .A(n20866), .B(n21269), .Z(n21267) );
  NAND U21526 ( .A(n21270), .B(n21271), .Z(n21269) );
  NANDN U21527 ( .A(n4967), .B(\stack[3][16] ), .Z(n21271) );
  NANDN U21528 ( .A(n20875), .B(\stack[1][16] ), .Z(n21270) );
  NAND U21529 ( .A(n21272), .B(n21273), .Z(n4818) );
  NANDN U21530 ( .A(n21188), .B(\stack[2][17] ), .Z(n21273) );
  NANDN U21531 ( .A(n20866), .B(n21274), .Z(n21272) );
  NAND U21532 ( .A(n21275), .B(n21276), .Z(n21274) );
  NANDN U21533 ( .A(n4967), .B(\stack[3][17] ), .Z(n21276) );
  NANDN U21534 ( .A(n20875), .B(\stack[1][17] ), .Z(n21275) );
  NAND U21535 ( .A(n21277), .B(n21278), .Z(n4817) );
  NANDN U21536 ( .A(n21188), .B(\stack[2][18] ), .Z(n21278) );
  NANDN U21537 ( .A(n20866), .B(n21279), .Z(n21277) );
  NAND U21538 ( .A(n21280), .B(n21281), .Z(n21279) );
  NANDN U21539 ( .A(n4967), .B(\stack[3][18] ), .Z(n21281) );
  NANDN U21540 ( .A(n20875), .B(\stack[1][18] ), .Z(n21280) );
  NAND U21541 ( .A(n21282), .B(n21283), .Z(n4816) );
  NANDN U21542 ( .A(n21188), .B(\stack[2][19] ), .Z(n21283) );
  NANDN U21543 ( .A(n20866), .B(n21284), .Z(n21282) );
  NAND U21544 ( .A(n21285), .B(n21286), .Z(n21284) );
  NANDN U21545 ( .A(n4967), .B(\stack[3][19] ), .Z(n21286) );
  NANDN U21546 ( .A(n20875), .B(\stack[1][19] ), .Z(n21285) );
  NAND U21547 ( .A(n21287), .B(n21288), .Z(n4815) );
  NANDN U21548 ( .A(n21188), .B(\stack[2][20] ), .Z(n21288) );
  NANDN U21549 ( .A(n20866), .B(n21289), .Z(n21287) );
  NAND U21550 ( .A(n21290), .B(n21291), .Z(n21289) );
  NANDN U21551 ( .A(n4967), .B(\stack[3][20] ), .Z(n21291) );
  NANDN U21552 ( .A(n20875), .B(\stack[1][20] ), .Z(n21290) );
  NAND U21553 ( .A(n21292), .B(n21293), .Z(n4814) );
  NANDN U21554 ( .A(n21188), .B(\stack[2][21] ), .Z(n21293) );
  NANDN U21555 ( .A(n20866), .B(n21294), .Z(n21292) );
  NAND U21556 ( .A(n21295), .B(n21296), .Z(n21294) );
  NANDN U21557 ( .A(n4967), .B(\stack[3][21] ), .Z(n21296) );
  NANDN U21558 ( .A(n20875), .B(\stack[1][21] ), .Z(n21295) );
  NAND U21559 ( .A(n21297), .B(n21298), .Z(n4813) );
  NANDN U21560 ( .A(n21188), .B(\stack[2][22] ), .Z(n21298) );
  NANDN U21561 ( .A(n20866), .B(n21299), .Z(n21297) );
  NAND U21562 ( .A(n21300), .B(n21301), .Z(n21299) );
  NANDN U21563 ( .A(n4967), .B(\stack[3][22] ), .Z(n21301) );
  NANDN U21564 ( .A(n20875), .B(\stack[1][22] ), .Z(n21300) );
  NAND U21565 ( .A(n21302), .B(n21303), .Z(n4812) );
  NANDN U21566 ( .A(n21188), .B(\stack[2][23] ), .Z(n21303) );
  NANDN U21567 ( .A(n20866), .B(n21304), .Z(n21302) );
  NAND U21568 ( .A(n21305), .B(n21306), .Z(n21304) );
  NANDN U21569 ( .A(n4967), .B(\stack[3][23] ), .Z(n21306) );
  NANDN U21570 ( .A(n20875), .B(\stack[1][23] ), .Z(n21305) );
  NAND U21571 ( .A(n21307), .B(n21308), .Z(n4811) );
  NANDN U21572 ( .A(n21188), .B(\stack[2][24] ), .Z(n21308) );
  NANDN U21573 ( .A(n20866), .B(n21309), .Z(n21307) );
  NAND U21574 ( .A(n21310), .B(n21311), .Z(n21309) );
  NANDN U21575 ( .A(n4967), .B(\stack[3][24] ), .Z(n21311) );
  NANDN U21576 ( .A(n20875), .B(\stack[1][24] ), .Z(n21310) );
  NAND U21577 ( .A(n21312), .B(n21313), .Z(n4810) );
  NANDN U21578 ( .A(n21188), .B(\stack[2][25] ), .Z(n21313) );
  NANDN U21579 ( .A(n20866), .B(n21314), .Z(n21312) );
  NAND U21580 ( .A(n21315), .B(n21316), .Z(n21314) );
  NANDN U21581 ( .A(n4967), .B(\stack[3][25] ), .Z(n21316) );
  NANDN U21582 ( .A(n20875), .B(\stack[1][25] ), .Z(n21315) );
  NAND U21583 ( .A(n21317), .B(n21318), .Z(n4809) );
  NANDN U21584 ( .A(n21188), .B(\stack[2][26] ), .Z(n21318) );
  NANDN U21585 ( .A(n20866), .B(n21319), .Z(n21317) );
  NAND U21586 ( .A(n21320), .B(n21321), .Z(n21319) );
  NANDN U21587 ( .A(n4967), .B(\stack[3][26] ), .Z(n21321) );
  NANDN U21588 ( .A(n20875), .B(\stack[1][26] ), .Z(n21320) );
  NAND U21589 ( .A(n21322), .B(n21323), .Z(n4808) );
  NANDN U21590 ( .A(n21188), .B(\stack[2][27] ), .Z(n21323) );
  NANDN U21591 ( .A(n20866), .B(n21324), .Z(n21322) );
  NAND U21592 ( .A(n21325), .B(n21326), .Z(n21324) );
  NANDN U21593 ( .A(n4967), .B(\stack[3][27] ), .Z(n21326) );
  NANDN U21594 ( .A(n20875), .B(\stack[1][27] ), .Z(n21325) );
  NAND U21595 ( .A(n21327), .B(n21328), .Z(n4807) );
  NANDN U21596 ( .A(n21188), .B(\stack[2][28] ), .Z(n21328) );
  NANDN U21597 ( .A(n20866), .B(n21329), .Z(n21327) );
  NAND U21598 ( .A(n21330), .B(n21331), .Z(n21329) );
  NANDN U21599 ( .A(n4967), .B(\stack[3][28] ), .Z(n21331) );
  NANDN U21600 ( .A(n20875), .B(\stack[1][28] ), .Z(n21330) );
  NAND U21601 ( .A(n21332), .B(n21333), .Z(n4806) );
  NANDN U21602 ( .A(n21188), .B(\stack[2][29] ), .Z(n21333) );
  NANDN U21603 ( .A(n20866), .B(n21334), .Z(n21332) );
  NAND U21604 ( .A(n21335), .B(n21336), .Z(n21334) );
  NANDN U21605 ( .A(n4967), .B(\stack[3][29] ), .Z(n21336) );
  NANDN U21606 ( .A(n20875), .B(\stack[1][29] ), .Z(n21335) );
  NAND U21607 ( .A(n21337), .B(n21338), .Z(n4805) );
  NANDN U21608 ( .A(n21188), .B(\stack[2][30] ), .Z(n21338) );
  NANDN U21609 ( .A(n20866), .B(n21339), .Z(n21337) );
  NAND U21610 ( .A(n21340), .B(n21341), .Z(n21339) );
  NANDN U21611 ( .A(n4967), .B(\stack[3][30] ), .Z(n21341) );
  NANDN U21612 ( .A(n20875), .B(\stack[1][30] ), .Z(n21340) );
  NAND U21613 ( .A(n21342), .B(n21343), .Z(n4804) );
  NANDN U21614 ( .A(n21188), .B(\stack[2][31] ), .Z(n21343) );
  NANDN U21615 ( .A(n20866), .B(n21344), .Z(n21342) );
  NAND U21616 ( .A(n21345), .B(n21346), .Z(n21344) );
  NANDN U21617 ( .A(n4967), .B(\stack[3][31] ), .Z(n21346) );
  NANDN U21618 ( .A(n20875), .B(\stack[1][31] ), .Z(n21345) );
  NAND U21619 ( .A(n21347), .B(n21348), .Z(n4803) );
  NANDN U21620 ( .A(n21188), .B(\stack[2][32] ), .Z(n21348) );
  NANDN U21621 ( .A(n20866), .B(n21349), .Z(n21347) );
  NAND U21622 ( .A(n21350), .B(n21351), .Z(n21349) );
  NANDN U21623 ( .A(n4967), .B(\stack[3][32] ), .Z(n21351) );
  NANDN U21624 ( .A(n20875), .B(\stack[1][32] ), .Z(n21350) );
  NAND U21625 ( .A(n21352), .B(n21353), .Z(n4802) );
  NANDN U21626 ( .A(n21188), .B(\stack[2][33] ), .Z(n21353) );
  NANDN U21627 ( .A(n20866), .B(n21354), .Z(n21352) );
  NAND U21628 ( .A(n21355), .B(n21356), .Z(n21354) );
  NANDN U21629 ( .A(n4967), .B(\stack[3][33] ), .Z(n21356) );
  NANDN U21630 ( .A(n20875), .B(\stack[1][33] ), .Z(n21355) );
  NAND U21631 ( .A(n21357), .B(n21358), .Z(n4801) );
  NANDN U21632 ( .A(n21188), .B(\stack[2][34] ), .Z(n21358) );
  NANDN U21633 ( .A(n20866), .B(n21359), .Z(n21357) );
  NAND U21634 ( .A(n21360), .B(n21361), .Z(n21359) );
  NANDN U21635 ( .A(n4967), .B(\stack[3][34] ), .Z(n21361) );
  NANDN U21636 ( .A(n20875), .B(\stack[1][34] ), .Z(n21360) );
  NAND U21637 ( .A(n21362), .B(n21363), .Z(n4800) );
  NANDN U21638 ( .A(n21188), .B(\stack[2][35] ), .Z(n21363) );
  NANDN U21639 ( .A(n20866), .B(n21364), .Z(n21362) );
  NAND U21640 ( .A(n21365), .B(n21366), .Z(n21364) );
  NANDN U21641 ( .A(n4967), .B(\stack[3][35] ), .Z(n21366) );
  NANDN U21642 ( .A(n20875), .B(\stack[1][35] ), .Z(n21365) );
  NAND U21643 ( .A(n21367), .B(n21368), .Z(n4799) );
  NANDN U21644 ( .A(n21188), .B(\stack[2][36] ), .Z(n21368) );
  NANDN U21645 ( .A(n20866), .B(n21369), .Z(n21367) );
  NAND U21646 ( .A(n21370), .B(n21371), .Z(n21369) );
  NANDN U21647 ( .A(n4967), .B(\stack[3][36] ), .Z(n21371) );
  NANDN U21648 ( .A(n20875), .B(\stack[1][36] ), .Z(n21370) );
  NAND U21649 ( .A(n21372), .B(n21373), .Z(n4798) );
  NANDN U21650 ( .A(n21188), .B(\stack[2][37] ), .Z(n21373) );
  NANDN U21651 ( .A(n20866), .B(n21374), .Z(n21372) );
  NAND U21652 ( .A(n21375), .B(n21376), .Z(n21374) );
  NANDN U21653 ( .A(n4967), .B(\stack[3][37] ), .Z(n21376) );
  NANDN U21654 ( .A(n20875), .B(\stack[1][37] ), .Z(n21375) );
  NAND U21655 ( .A(n21377), .B(n21378), .Z(n4797) );
  NANDN U21656 ( .A(n21188), .B(\stack[2][38] ), .Z(n21378) );
  NANDN U21657 ( .A(n20866), .B(n21379), .Z(n21377) );
  NAND U21658 ( .A(n21380), .B(n21381), .Z(n21379) );
  NANDN U21659 ( .A(n4967), .B(\stack[3][38] ), .Z(n21381) );
  NANDN U21660 ( .A(n20875), .B(\stack[1][38] ), .Z(n21380) );
  NAND U21661 ( .A(n21382), .B(n21383), .Z(n4796) );
  NANDN U21662 ( .A(n21188), .B(\stack[2][39] ), .Z(n21383) );
  NANDN U21663 ( .A(n20866), .B(n21384), .Z(n21382) );
  NAND U21664 ( .A(n21385), .B(n21386), .Z(n21384) );
  NANDN U21665 ( .A(n4967), .B(\stack[3][39] ), .Z(n21386) );
  NANDN U21666 ( .A(n20875), .B(\stack[1][39] ), .Z(n21385) );
  NAND U21667 ( .A(n21387), .B(n21388), .Z(n4795) );
  NANDN U21668 ( .A(n21188), .B(\stack[2][40] ), .Z(n21388) );
  NANDN U21669 ( .A(n20866), .B(n21389), .Z(n21387) );
  NAND U21670 ( .A(n21390), .B(n21391), .Z(n21389) );
  NANDN U21671 ( .A(n4967), .B(\stack[3][40] ), .Z(n21391) );
  NANDN U21672 ( .A(n20875), .B(\stack[1][40] ), .Z(n21390) );
  NAND U21673 ( .A(n21392), .B(n21393), .Z(n4794) );
  NANDN U21674 ( .A(n21188), .B(\stack[2][41] ), .Z(n21393) );
  NANDN U21675 ( .A(n20866), .B(n21394), .Z(n21392) );
  NAND U21676 ( .A(n21395), .B(n21396), .Z(n21394) );
  NANDN U21677 ( .A(n4967), .B(\stack[3][41] ), .Z(n21396) );
  NANDN U21678 ( .A(n20875), .B(\stack[1][41] ), .Z(n21395) );
  NAND U21679 ( .A(n21397), .B(n21398), .Z(n4793) );
  NANDN U21680 ( .A(n21188), .B(\stack[2][42] ), .Z(n21398) );
  NANDN U21681 ( .A(n20866), .B(n21399), .Z(n21397) );
  NAND U21682 ( .A(n21400), .B(n21401), .Z(n21399) );
  NANDN U21683 ( .A(n4967), .B(\stack[3][42] ), .Z(n21401) );
  NANDN U21684 ( .A(n20875), .B(\stack[1][42] ), .Z(n21400) );
  NAND U21685 ( .A(n21402), .B(n21403), .Z(n4792) );
  NANDN U21686 ( .A(n21188), .B(\stack[2][43] ), .Z(n21403) );
  NANDN U21687 ( .A(n20866), .B(n21404), .Z(n21402) );
  NAND U21688 ( .A(n21405), .B(n21406), .Z(n21404) );
  NANDN U21689 ( .A(n4967), .B(\stack[3][43] ), .Z(n21406) );
  NANDN U21690 ( .A(n20875), .B(\stack[1][43] ), .Z(n21405) );
  NAND U21691 ( .A(n21407), .B(n21408), .Z(n4791) );
  NANDN U21692 ( .A(n21188), .B(\stack[2][44] ), .Z(n21408) );
  NANDN U21693 ( .A(n20866), .B(n21409), .Z(n21407) );
  NAND U21694 ( .A(n21410), .B(n21411), .Z(n21409) );
  NANDN U21695 ( .A(n4967), .B(\stack[3][44] ), .Z(n21411) );
  NANDN U21696 ( .A(n20875), .B(\stack[1][44] ), .Z(n21410) );
  NAND U21697 ( .A(n21412), .B(n21413), .Z(n4790) );
  NANDN U21698 ( .A(n21188), .B(\stack[2][45] ), .Z(n21413) );
  NANDN U21699 ( .A(n20866), .B(n21414), .Z(n21412) );
  NAND U21700 ( .A(n21415), .B(n21416), .Z(n21414) );
  NANDN U21701 ( .A(n4967), .B(\stack[3][45] ), .Z(n21416) );
  NANDN U21702 ( .A(n20875), .B(\stack[1][45] ), .Z(n21415) );
  NAND U21703 ( .A(n21417), .B(n21418), .Z(n4789) );
  NANDN U21704 ( .A(n21188), .B(\stack[2][46] ), .Z(n21418) );
  NANDN U21705 ( .A(n20866), .B(n21419), .Z(n21417) );
  NAND U21706 ( .A(n21420), .B(n21421), .Z(n21419) );
  NANDN U21707 ( .A(n4967), .B(\stack[3][46] ), .Z(n21421) );
  NANDN U21708 ( .A(n20875), .B(\stack[1][46] ), .Z(n21420) );
  NAND U21709 ( .A(n21422), .B(n21423), .Z(n4788) );
  NANDN U21710 ( .A(n21188), .B(\stack[2][47] ), .Z(n21423) );
  NANDN U21711 ( .A(n20866), .B(n21424), .Z(n21422) );
  NAND U21712 ( .A(n21425), .B(n21426), .Z(n21424) );
  NANDN U21713 ( .A(n4967), .B(\stack[3][47] ), .Z(n21426) );
  NANDN U21714 ( .A(n20875), .B(\stack[1][47] ), .Z(n21425) );
  NAND U21715 ( .A(n21427), .B(n21428), .Z(n4787) );
  NANDN U21716 ( .A(n21188), .B(\stack[2][48] ), .Z(n21428) );
  NANDN U21717 ( .A(n20866), .B(n21429), .Z(n21427) );
  NAND U21718 ( .A(n21430), .B(n21431), .Z(n21429) );
  NANDN U21719 ( .A(n4967), .B(\stack[3][48] ), .Z(n21431) );
  NANDN U21720 ( .A(n20875), .B(\stack[1][48] ), .Z(n21430) );
  NAND U21721 ( .A(n21432), .B(n21433), .Z(n4786) );
  NANDN U21722 ( .A(n21188), .B(\stack[2][49] ), .Z(n21433) );
  NANDN U21723 ( .A(n20866), .B(n21434), .Z(n21432) );
  NAND U21724 ( .A(n21435), .B(n21436), .Z(n21434) );
  NANDN U21725 ( .A(n4967), .B(\stack[3][49] ), .Z(n21436) );
  NANDN U21726 ( .A(n20875), .B(\stack[1][49] ), .Z(n21435) );
  NAND U21727 ( .A(n21437), .B(n21438), .Z(n4785) );
  NANDN U21728 ( .A(n21188), .B(\stack[2][50] ), .Z(n21438) );
  NANDN U21729 ( .A(n20866), .B(n21439), .Z(n21437) );
  NAND U21730 ( .A(n21440), .B(n21441), .Z(n21439) );
  NANDN U21731 ( .A(n4967), .B(\stack[3][50] ), .Z(n21441) );
  NANDN U21732 ( .A(n20875), .B(\stack[1][50] ), .Z(n21440) );
  NAND U21733 ( .A(n21442), .B(n21443), .Z(n4784) );
  NANDN U21734 ( .A(n21188), .B(\stack[2][51] ), .Z(n21443) );
  NANDN U21735 ( .A(n20866), .B(n21444), .Z(n21442) );
  NAND U21736 ( .A(n21445), .B(n21446), .Z(n21444) );
  NANDN U21737 ( .A(n4967), .B(\stack[3][51] ), .Z(n21446) );
  NANDN U21738 ( .A(n20875), .B(\stack[1][51] ), .Z(n21445) );
  NAND U21739 ( .A(n21447), .B(n21448), .Z(n4783) );
  NANDN U21740 ( .A(n21188), .B(\stack[2][52] ), .Z(n21448) );
  NANDN U21741 ( .A(n20866), .B(n21449), .Z(n21447) );
  NAND U21742 ( .A(n21450), .B(n21451), .Z(n21449) );
  NANDN U21743 ( .A(n4967), .B(\stack[3][52] ), .Z(n21451) );
  NANDN U21744 ( .A(n20875), .B(\stack[1][52] ), .Z(n21450) );
  NAND U21745 ( .A(n21452), .B(n21453), .Z(n4782) );
  NANDN U21746 ( .A(n21188), .B(\stack[2][53] ), .Z(n21453) );
  NANDN U21747 ( .A(n20866), .B(n21454), .Z(n21452) );
  NAND U21748 ( .A(n21455), .B(n21456), .Z(n21454) );
  NANDN U21749 ( .A(n4967), .B(\stack[3][53] ), .Z(n21456) );
  NANDN U21750 ( .A(n20875), .B(\stack[1][53] ), .Z(n21455) );
  NAND U21751 ( .A(n21457), .B(n21458), .Z(n4781) );
  NANDN U21752 ( .A(n21188), .B(\stack[2][54] ), .Z(n21458) );
  NANDN U21753 ( .A(n20866), .B(n21459), .Z(n21457) );
  NAND U21754 ( .A(n21460), .B(n21461), .Z(n21459) );
  NANDN U21755 ( .A(n4967), .B(\stack[3][54] ), .Z(n21461) );
  NANDN U21756 ( .A(n20875), .B(\stack[1][54] ), .Z(n21460) );
  NAND U21757 ( .A(n21462), .B(n21463), .Z(n4780) );
  NANDN U21758 ( .A(n21188), .B(\stack[2][55] ), .Z(n21463) );
  NANDN U21759 ( .A(n20866), .B(n21464), .Z(n21462) );
  NAND U21760 ( .A(n21465), .B(n21466), .Z(n21464) );
  NANDN U21761 ( .A(n4967), .B(\stack[3][55] ), .Z(n21466) );
  NANDN U21762 ( .A(n20875), .B(\stack[1][55] ), .Z(n21465) );
  NAND U21763 ( .A(n21467), .B(n21468), .Z(n4779) );
  NANDN U21764 ( .A(n21188), .B(\stack[2][56] ), .Z(n21468) );
  NANDN U21765 ( .A(n20866), .B(n21469), .Z(n21467) );
  NAND U21766 ( .A(n21470), .B(n21471), .Z(n21469) );
  NANDN U21767 ( .A(n4967), .B(\stack[3][56] ), .Z(n21471) );
  NANDN U21768 ( .A(n20875), .B(\stack[1][56] ), .Z(n21470) );
  NAND U21769 ( .A(n21472), .B(n21473), .Z(n4778) );
  NANDN U21770 ( .A(n21188), .B(\stack[2][57] ), .Z(n21473) );
  NANDN U21771 ( .A(n20866), .B(n21474), .Z(n21472) );
  NAND U21772 ( .A(n21475), .B(n21476), .Z(n21474) );
  NANDN U21773 ( .A(n4967), .B(\stack[3][57] ), .Z(n21476) );
  NANDN U21774 ( .A(n20875), .B(\stack[1][57] ), .Z(n21475) );
  NAND U21775 ( .A(n21477), .B(n21478), .Z(n4777) );
  NANDN U21776 ( .A(n21188), .B(\stack[2][58] ), .Z(n21478) );
  NANDN U21777 ( .A(n20866), .B(n21479), .Z(n21477) );
  NAND U21778 ( .A(n21480), .B(n21481), .Z(n21479) );
  NANDN U21779 ( .A(n4967), .B(\stack[3][58] ), .Z(n21481) );
  NANDN U21780 ( .A(n20875), .B(\stack[1][58] ), .Z(n21480) );
  NAND U21781 ( .A(n21482), .B(n21483), .Z(n4776) );
  NANDN U21782 ( .A(n21188), .B(\stack[2][59] ), .Z(n21483) );
  NANDN U21783 ( .A(n20866), .B(n21484), .Z(n21482) );
  NAND U21784 ( .A(n21485), .B(n21486), .Z(n21484) );
  NANDN U21785 ( .A(n4967), .B(\stack[3][59] ), .Z(n21486) );
  NANDN U21786 ( .A(n20875), .B(\stack[1][59] ), .Z(n21485) );
  NAND U21787 ( .A(n21487), .B(n21488), .Z(n4775) );
  NANDN U21788 ( .A(n21188), .B(\stack[2][60] ), .Z(n21488) );
  NANDN U21789 ( .A(n20866), .B(n21489), .Z(n21487) );
  NAND U21790 ( .A(n21490), .B(n21491), .Z(n21489) );
  NANDN U21791 ( .A(n4967), .B(\stack[3][60] ), .Z(n21491) );
  NANDN U21792 ( .A(n20875), .B(\stack[1][60] ), .Z(n21490) );
  NAND U21793 ( .A(n21492), .B(n21493), .Z(n4774) );
  NANDN U21794 ( .A(n21188), .B(\stack[2][61] ), .Z(n21493) );
  NANDN U21795 ( .A(n20866), .B(n21494), .Z(n21492) );
  NAND U21796 ( .A(n21495), .B(n21496), .Z(n21494) );
  NANDN U21797 ( .A(n4967), .B(\stack[3][61] ), .Z(n21496) );
  NANDN U21798 ( .A(n20875), .B(\stack[1][61] ), .Z(n21495) );
  NAND U21799 ( .A(n21497), .B(n21498), .Z(n4773) );
  NANDN U21800 ( .A(n21188), .B(\stack[2][62] ), .Z(n21498) );
  NANDN U21801 ( .A(n20866), .B(n21499), .Z(n21497) );
  NAND U21802 ( .A(n21500), .B(n21501), .Z(n21499) );
  NANDN U21803 ( .A(n4967), .B(\stack[3][62] ), .Z(n21501) );
  NANDN U21804 ( .A(n20875), .B(\stack[1][62] ), .Z(n21500) );
  NAND U21805 ( .A(n21502), .B(n21503), .Z(n4772) );
  NANDN U21806 ( .A(n21188), .B(\stack[2][63] ), .Z(n21503) );
  NANDN U21807 ( .A(n20866), .B(n21504), .Z(n21502) );
  NAND U21808 ( .A(n21505), .B(n21506), .Z(n21504) );
  NANDN U21809 ( .A(n4967), .B(\stack[3][63] ), .Z(n21506) );
  NANDN U21810 ( .A(n20875), .B(\stack[1][63] ), .Z(n21505) );
  NAND U21811 ( .A(n21507), .B(n21508), .Z(n4771) );
  NANDN U21812 ( .A(n21188), .B(\stack[3][0] ), .Z(n21508) );
  NANDN U21813 ( .A(n20866), .B(n21509), .Z(n21507) );
  NAND U21814 ( .A(n21510), .B(n21511), .Z(n21509) );
  NANDN U21815 ( .A(n4967), .B(\stack[4][0] ), .Z(n21511) );
  NANDN U21816 ( .A(n20875), .B(\stack[2][0] ), .Z(n21510) );
  NAND U21817 ( .A(n21512), .B(n21513), .Z(n4770) );
  NANDN U21818 ( .A(n21188), .B(\stack[3][1] ), .Z(n21513) );
  NANDN U21819 ( .A(n20866), .B(n21514), .Z(n21512) );
  NAND U21820 ( .A(n21515), .B(n21516), .Z(n21514) );
  NANDN U21821 ( .A(n4967), .B(\stack[4][1] ), .Z(n21516) );
  NANDN U21822 ( .A(n20875), .B(\stack[2][1] ), .Z(n21515) );
  NAND U21823 ( .A(n21517), .B(n21518), .Z(n4769) );
  NANDN U21824 ( .A(n21188), .B(\stack[3][2] ), .Z(n21518) );
  NANDN U21825 ( .A(n20866), .B(n21519), .Z(n21517) );
  NAND U21826 ( .A(n21520), .B(n21521), .Z(n21519) );
  NANDN U21827 ( .A(n4967), .B(\stack[4][2] ), .Z(n21521) );
  NANDN U21828 ( .A(n20875), .B(\stack[2][2] ), .Z(n21520) );
  NAND U21829 ( .A(n21522), .B(n21523), .Z(n4768) );
  NANDN U21830 ( .A(n21188), .B(\stack[3][3] ), .Z(n21523) );
  NANDN U21831 ( .A(n20866), .B(n21524), .Z(n21522) );
  NAND U21832 ( .A(n21525), .B(n21526), .Z(n21524) );
  NANDN U21833 ( .A(n4967), .B(\stack[4][3] ), .Z(n21526) );
  NANDN U21834 ( .A(n20875), .B(\stack[2][3] ), .Z(n21525) );
  NAND U21835 ( .A(n21527), .B(n21528), .Z(n4767) );
  NANDN U21836 ( .A(n21188), .B(\stack[3][4] ), .Z(n21528) );
  NANDN U21837 ( .A(n20866), .B(n21529), .Z(n21527) );
  NAND U21838 ( .A(n21530), .B(n21531), .Z(n21529) );
  NANDN U21839 ( .A(n4967), .B(\stack[4][4] ), .Z(n21531) );
  NANDN U21840 ( .A(n20875), .B(\stack[2][4] ), .Z(n21530) );
  NAND U21841 ( .A(n21532), .B(n21533), .Z(n4766) );
  NANDN U21842 ( .A(n21188), .B(\stack[3][5] ), .Z(n21533) );
  NANDN U21843 ( .A(n20866), .B(n21534), .Z(n21532) );
  NAND U21844 ( .A(n21535), .B(n21536), .Z(n21534) );
  NANDN U21845 ( .A(n4967), .B(\stack[4][5] ), .Z(n21536) );
  NANDN U21846 ( .A(n20875), .B(\stack[2][5] ), .Z(n21535) );
  NAND U21847 ( .A(n21537), .B(n21538), .Z(n4765) );
  NANDN U21848 ( .A(n21188), .B(\stack[3][6] ), .Z(n21538) );
  NANDN U21849 ( .A(n20866), .B(n21539), .Z(n21537) );
  NAND U21850 ( .A(n21540), .B(n21541), .Z(n21539) );
  NANDN U21851 ( .A(n4967), .B(\stack[4][6] ), .Z(n21541) );
  NANDN U21852 ( .A(n20875), .B(\stack[2][6] ), .Z(n21540) );
  NAND U21853 ( .A(n21542), .B(n21543), .Z(n4764) );
  NANDN U21854 ( .A(n21188), .B(\stack[3][7] ), .Z(n21543) );
  NANDN U21855 ( .A(n20866), .B(n21544), .Z(n21542) );
  NAND U21856 ( .A(n21545), .B(n21546), .Z(n21544) );
  NANDN U21857 ( .A(n4967), .B(\stack[4][7] ), .Z(n21546) );
  NANDN U21858 ( .A(n20875), .B(\stack[2][7] ), .Z(n21545) );
  NAND U21859 ( .A(n21547), .B(n21548), .Z(n4763) );
  NANDN U21860 ( .A(n21188), .B(\stack[3][8] ), .Z(n21548) );
  NANDN U21861 ( .A(n20866), .B(n21549), .Z(n21547) );
  NAND U21862 ( .A(n21550), .B(n21551), .Z(n21549) );
  NANDN U21863 ( .A(n4967), .B(\stack[4][8] ), .Z(n21551) );
  NANDN U21864 ( .A(n20875), .B(\stack[2][8] ), .Z(n21550) );
  NAND U21865 ( .A(n21552), .B(n21553), .Z(n4762) );
  NANDN U21866 ( .A(n21188), .B(\stack[3][9] ), .Z(n21553) );
  NANDN U21867 ( .A(n20866), .B(n21554), .Z(n21552) );
  NAND U21868 ( .A(n21555), .B(n21556), .Z(n21554) );
  NANDN U21869 ( .A(n4967), .B(\stack[4][9] ), .Z(n21556) );
  NANDN U21870 ( .A(n20875), .B(\stack[2][9] ), .Z(n21555) );
  NAND U21871 ( .A(n21557), .B(n21558), .Z(n4761) );
  NANDN U21872 ( .A(n21188), .B(\stack[3][10] ), .Z(n21558) );
  NANDN U21873 ( .A(n20866), .B(n21559), .Z(n21557) );
  NAND U21874 ( .A(n21560), .B(n21561), .Z(n21559) );
  NANDN U21875 ( .A(n4967), .B(\stack[4][10] ), .Z(n21561) );
  NANDN U21876 ( .A(n20875), .B(\stack[2][10] ), .Z(n21560) );
  NAND U21877 ( .A(n21562), .B(n21563), .Z(n4760) );
  NANDN U21878 ( .A(n21188), .B(\stack[3][11] ), .Z(n21563) );
  NANDN U21879 ( .A(n20866), .B(n21564), .Z(n21562) );
  NAND U21880 ( .A(n21565), .B(n21566), .Z(n21564) );
  NANDN U21881 ( .A(n4967), .B(\stack[4][11] ), .Z(n21566) );
  NANDN U21882 ( .A(n20875), .B(\stack[2][11] ), .Z(n21565) );
  NAND U21883 ( .A(n21567), .B(n21568), .Z(n4759) );
  NANDN U21884 ( .A(n21188), .B(\stack[3][12] ), .Z(n21568) );
  NANDN U21885 ( .A(n20866), .B(n21569), .Z(n21567) );
  NAND U21886 ( .A(n21570), .B(n21571), .Z(n21569) );
  NANDN U21887 ( .A(n4967), .B(\stack[4][12] ), .Z(n21571) );
  NANDN U21888 ( .A(n20875), .B(\stack[2][12] ), .Z(n21570) );
  NAND U21889 ( .A(n21572), .B(n21573), .Z(n4758) );
  NANDN U21890 ( .A(n21188), .B(\stack[3][13] ), .Z(n21573) );
  NANDN U21891 ( .A(n20866), .B(n21574), .Z(n21572) );
  NAND U21892 ( .A(n21575), .B(n21576), .Z(n21574) );
  NANDN U21893 ( .A(n4967), .B(\stack[4][13] ), .Z(n21576) );
  NANDN U21894 ( .A(n20875), .B(\stack[2][13] ), .Z(n21575) );
  NAND U21895 ( .A(n21577), .B(n21578), .Z(n4757) );
  NANDN U21896 ( .A(n21188), .B(\stack[3][14] ), .Z(n21578) );
  NANDN U21897 ( .A(n20866), .B(n21579), .Z(n21577) );
  NAND U21898 ( .A(n21580), .B(n21581), .Z(n21579) );
  NANDN U21899 ( .A(n4967), .B(\stack[4][14] ), .Z(n21581) );
  NANDN U21900 ( .A(n20875), .B(\stack[2][14] ), .Z(n21580) );
  NAND U21901 ( .A(n21582), .B(n21583), .Z(n4756) );
  NANDN U21902 ( .A(n21188), .B(\stack[3][15] ), .Z(n21583) );
  NANDN U21903 ( .A(n20866), .B(n21584), .Z(n21582) );
  NAND U21904 ( .A(n21585), .B(n21586), .Z(n21584) );
  NANDN U21905 ( .A(n4967), .B(\stack[4][15] ), .Z(n21586) );
  NANDN U21906 ( .A(n20875), .B(\stack[2][15] ), .Z(n21585) );
  NAND U21907 ( .A(n21587), .B(n21588), .Z(n4755) );
  NANDN U21908 ( .A(n21188), .B(\stack[3][16] ), .Z(n21588) );
  NANDN U21909 ( .A(n20866), .B(n21589), .Z(n21587) );
  NAND U21910 ( .A(n21590), .B(n21591), .Z(n21589) );
  NANDN U21911 ( .A(n4967), .B(\stack[4][16] ), .Z(n21591) );
  NANDN U21912 ( .A(n20875), .B(\stack[2][16] ), .Z(n21590) );
  NAND U21913 ( .A(n21592), .B(n21593), .Z(n4754) );
  NANDN U21914 ( .A(n21188), .B(\stack[3][17] ), .Z(n21593) );
  NANDN U21915 ( .A(n20866), .B(n21594), .Z(n21592) );
  NAND U21916 ( .A(n21595), .B(n21596), .Z(n21594) );
  NANDN U21917 ( .A(n4967), .B(\stack[4][17] ), .Z(n21596) );
  NANDN U21918 ( .A(n20875), .B(\stack[2][17] ), .Z(n21595) );
  NAND U21919 ( .A(n21597), .B(n21598), .Z(n4753) );
  NANDN U21920 ( .A(n21188), .B(\stack[3][18] ), .Z(n21598) );
  NANDN U21921 ( .A(n20866), .B(n21599), .Z(n21597) );
  NAND U21922 ( .A(n21600), .B(n21601), .Z(n21599) );
  NANDN U21923 ( .A(n4967), .B(\stack[4][18] ), .Z(n21601) );
  NANDN U21924 ( .A(n20875), .B(\stack[2][18] ), .Z(n21600) );
  NAND U21925 ( .A(n21602), .B(n21603), .Z(n4752) );
  NANDN U21926 ( .A(n21188), .B(\stack[3][19] ), .Z(n21603) );
  NANDN U21927 ( .A(n20866), .B(n21604), .Z(n21602) );
  NAND U21928 ( .A(n21605), .B(n21606), .Z(n21604) );
  NANDN U21929 ( .A(n4967), .B(\stack[4][19] ), .Z(n21606) );
  NANDN U21930 ( .A(n20875), .B(\stack[2][19] ), .Z(n21605) );
  NAND U21931 ( .A(n21607), .B(n21608), .Z(n4751) );
  NANDN U21932 ( .A(n21188), .B(\stack[3][20] ), .Z(n21608) );
  NANDN U21933 ( .A(n20866), .B(n21609), .Z(n21607) );
  NAND U21934 ( .A(n21610), .B(n21611), .Z(n21609) );
  NANDN U21935 ( .A(n4967), .B(\stack[4][20] ), .Z(n21611) );
  NANDN U21936 ( .A(n20875), .B(\stack[2][20] ), .Z(n21610) );
  NAND U21937 ( .A(n21612), .B(n21613), .Z(n4750) );
  NANDN U21938 ( .A(n21188), .B(\stack[3][21] ), .Z(n21613) );
  NANDN U21939 ( .A(n20866), .B(n21614), .Z(n21612) );
  NAND U21940 ( .A(n21615), .B(n21616), .Z(n21614) );
  NANDN U21941 ( .A(n4967), .B(\stack[4][21] ), .Z(n21616) );
  NANDN U21942 ( .A(n20875), .B(\stack[2][21] ), .Z(n21615) );
  NAND U21943 ( .A(n21617), .B(n21618), .Z(n4749) );
  NANDN U21944 ( .A(n21188), .B(\stack[3][22] ), .Z(n21618) );
  NANDN U21945 ( .A(n20866), .B(n21619), .Z(n21617) );
  NAND U21946 ( .A(n21620), .B(n21621), .Z(n21619) );
  NANDN U21947 ( .A(n4967), .B(\stack[4][22] ), .Z(n21621) );
  NANDN U21948 ( .A(n20875), .B(\stack[2][22] ), .Z(n21620) );
  NAND U21949 ( .A(n21622), .B(n21623), .Z(n4748) );
  NANDN U21950 ( .A(n21188), .B(\stack[3][23] ), .Z(n21623) );
  NANDN U21951 ( .A(n20866), .B(n21624), .Z(n21622) );
  NAND U21952 ( .A(n21625), .B(n21626), .Z(n21624) );
  NANDN U21953 ( .A(n4967), .B(\stack[4][23] ), .Z(n21626) );
  NANDN U21954 ( .A(n20875), .B(\stack[2][23] ), .Z(n21625) );
  NAND U21955 ( .A(n21627), .B(n21628), .Z(n4747) );
  NANDN U21956 ( .A(n21188), .B(\stack[3][24] ), .Z(n21628) );
  NANDN U21957 ( .A(n20866), .B(n21629), .Z(n21627) );
  NAND U21958 ( .A(n21630), .B(n21631), .Z(n21629) );
  NANDN U21959 ( .A(n4967), .B(\stack[4][24] ), .Z(n21631) );
  NANDN U21960 ( .A(n20875), .B(\stack[2][24] ), .Z(n21630) );
  NAND U21961 ( .A(n21632), .B(n21633), .Z(n4746) );
  NANDN U21962 ( .A(n21188), .B(\stack[3][25] ), .Z(n21633) );
  NANDN U21963 ( .A(n20866), .B(n21634), .Z(n21632) );
  NAND U21964 ( .A(n21635), .B(n21636), .Z(n21634) );
  NANDN U21965 ( .A(n4967), .B(\stack[4][25] ), .Z(n21636) );
  NANDN U21966 ( .A(n20875), .B(\stack[2][25] ), .Z(n21635) );
  NAND U21967 ( .A(n21637), .B(n21638), .Z(n4745) );
  NANDN U21968 ( .A(n21188), .B(\stack[3][26] ), .Z(n21638) );
  NANDN U21969 ( .A(n20866), .B(n21639), .Z(n21637) );
  NAND U21970 ( .A(n21640), .B(n21641), .Z(n21639) );
  NANDN U21971 ( .A(n4967), .B(\stack[4][26] ), .Z(n21641) );
  NANDN U21972 ( .A(n20875), .B(\stack[2][26] ), .Z(n21640) );
  NAND U21973 ( .A(n21642), .B(n21643), .Z(n4744) );
  NANDN U21974 ( .A(n21188), .B(\stack[3][27] ), .Z(n21643) );
  NANDN U21975 ( .A(n20866), .B(n21644), .Z(n21642) );
  NAND U21976 ( .A(n21645), .B(n21646), .Z(n21644) );
  NANDN U21977 ( .A(n4967), .B(\stack[4][27] ), .Z(n21646) );
  NANDN U21978 ( .A(n20875), .B(\stack[2][27] ), .Z(n21645) );
  NAND U21979 ( .A(n21647), .B(n21648), .Z(n4743) );
  NANDN U21980 ( .A(n21188), .B(\stack[3][28] ), .Z(n21648) );
  NANDN U21981 ( .A(n20866), .B(n21649), .Z(n21647) );
  NAND U21982 ( .A(n21650), .B(n21651), .Z(n21649) );
  NANDN U21983 ( .A(n4967), .B(\stack[4][28] ), .Z(n21651) );
  NANDN U21984 ( .A(n20875), .B(\stack[2][28] ), .Z(n21650) );
  NAND U21985 ( .A(n21652), .B(n21653), .Z(n4742) );
  NANDN U21986 ( .A(n21188), .B(\stack[3][29] ), .Z(n21653) );
  NANDN U21987 ( .A(n20866), .B(n21654), .Z(n21652) );
  NAND U21988 ( .A(n21655), .B(n21656), .Z(n21654) );
  NANDN U21989 ( .A(n4967), .B(\stack[4][29] ), .Z(n21656) );
  NANDN U21990 ( .A(n20875), .B(\stack[2][29] ), .Z(n21655) );
  NAND U21991 ( .A(n21657), .B(n21658), .Z(n4741) );
  NANDN U21992 ( .A(n21188), .B(\stack[3][30] ), .Z(n21658) );
  NANDN U21993 ( .A(n20866), .B(n21659), .Z(n21657) );
  NAND U21994 ( .A(n21660), .B(n21661), .Z(n21659) );
  NANDN U21995 ( .A(n4967), .B(\stack[4][30] ), .Z(n21661) );
  NANDN U21996 ( .A(n20875), .B(\stack[2][30] ), .Z(n21660) );
  NAND U21997 ( .A(n21662), .B(n21663), .Z(n4740) );
  NANDN U21998 ( .A(n21188), .B(\stack[3][31] ), .Z(n21663) );
  NANDN U21999 ( .A(n20866), .B(n21664), .Z(n21662) );
  NAND U22000 ( .A(n21665), .B(n21666), .Z(n21664) );
  NANDN U22001 ( .A(n4967), .B(\stack[4][31] ), .Z(n21666) );
  NANDN U22002 ( .A(n20875), .B(\stack[2][31] ), .Z(n21665) );
  NAND U22003 ( .A(n21667), .B(n21668), .Z(n4739) );
  NANDN U22004 ( .A(n21188), .B(\stack[3][32] ), .Z(n21668) );
  NANDN U22005 ( .A(n20866), .B(n21669), .Z(n21667) );
  NAND U22006 ( .A(n21670), .B(n21671), .Z(n21669) );
  NANDN U22007 ( .A(n4967), .B(\stack[4][32] ), .Z(n21671) );
  NANDN U22008 ( .A(n20875), .B(\stack[2][32] ), .Z(n21670) );
  NAND U22009 ( .A(n21672), .B(n21673), .Z(n4738) );
  NANDN U22010 ( .A(n21188), .B(\stack[3][33] ), .Z(n21673) );
  NANDN U22011 ( .A(n20866), .B(n21674), .Z(n21672) );
  NAND U22012 ( .A(n21675), .B(n21676), .Z(n21674) );
  NANDN U22013 ( .A(n4967), .B(\stack[4][33] ), .Z(n21676) );
  NANDN U22014 ( .A(n20875), .B(\stack[2][33] ), .Z(n21675) );
  NAND U22015 ( .A(n21677), .B(n21678), .Z(n4737) );
  NANDN U22016 ( .A(n21188), .B(\stack[3][34] ), .Z(n21678) );
  NANDN U22017 ( .A(n20866), .B(n21679), .Z(n21677) );
  NAND U22018 ( .A(n21680), .B(n21681), .Z(n21679) );
  NANDN U22019 ( .A(n4967), .B(\stack[4][34] ), .Z(n21681) );
  NANDN U22020 ( .A(n20875), .B(\stack[2][34] ), .Z(n21680) );
  NAND U22021 ( .A(n21682), .B(n21683), .Z(n4736) );
  NANDN U22022 ( .A(n21188), .B(\stack[3][35] ), .Z(n21683) );
  NANDN U22023 ( .A(n20866), .B(n21684), .Z(n21682) );
  NAND U22024 ( .A(n21685), .B(n21686), .Z(n21684) );
  NANDN U22025 ( .A(n4967), .B(\stack[4][35] ), .Z(n21686) );
  NANDN U22026 ( .A(n20875), .B(\stack[2][35] ), .Z(n21685) );
  NAND U22027 ( .A(n21687), .B(n21688), .Z(n4735) );
  NANDN U22028 ( .A(n21188), .B(\stack[3][36] ), .Z(n21688) );
  NANDN U22029 ( .A(n20866), .B(n21689), .Z(n21687) );
  NAND U22030 ( .A(n21690), .B(n21691), .Z(n21689) );
  NANDN U22031 ( .A(n4967), .B(\stack[4][36] ), .Z(n21691) );
  NANDN U22032 ( .A(n20875), .B(\stack[2][36] ), .Z(n21690) );
  NAND U22033 ( .A(n21692), .B(n21693), .Z(n4734) );
  NANDN U22034 ( .A(n21188), .B(\stack[3][37] ), .Z(n21693) );
  NANDN U22035 ( .A(n20866), .B(n21694), .Z(n21692) );
  NAND U22036 ( .A(n21695), .B(n21696), .Z(n21694) );
  NANDN U22037 ( .A(n4967), .B(\stack[4][37] ), .Z(n21696) );
  NANDN U22038 ( .A(n20875), .B(\stack[2][37] ), .Z(n21695) );
  NAND U22039 ( .A(n21697), .B(n21698), .Z(n4733) );
  NANDN U22040 ( .A(n21188), .B(\stack[3][38] ), .Z(n21698) );
  NANDN U22041 ( .A(n20866), .B(n21699), .Z(n21697) );
  NAND U22042 ( .A(n21700), .B(n21701), .Z(n21699) );
  NANDN U22043 ( .A(n4967), .B(\stack[4][38] ), .Z(n21701) );
  NANDN U22044 ( .A(n20875), .B(\stack[2][38] ), .Z(n21700) );
  NAND U22045 ( .A(n21702), .B(n21703), .Z(n4732) );
  NANDN U22046 ( .A(n21188), .B(\stack[3][39] ), .Z(n21703) );
  NANDN U22047 ( .A(n20866), .B(n21704), .Z(n21702) );
  NAND U22048 ( .A(n21705), .B(n21706), .Z(n21704) );
  NANDN U22049 ( .A(n4967), .B(\stack[4][39] ), .Z(n21706) );
  NANDN U22050 ( .A(n20875), .B(\stack[2][39] ), .Z(n21705) );
  NAND U22051 ( .A(n21707), .B(n21708), .Z(n4731) );
  NANDN U22052 ( .A(n21188), .B(\stack[3][40] ), .Z(n21708) );
  NANDN U22053 ( .A(n20866), .B(n21709), .Z(n21707) );
  NAND U22054 ( .A(n21710), .B(n21711), .Z(n21709) );
  NANDN U22055 ( .A(n4967), .B(\stack[4][40] ), .Z(n21711) );
  NANDN U22056 ( .A(n20875), .B(\stack[2][40] ), .Z(n21710) );
  NAND U22057 ( .A(n21712), .B(n21713), .Z(n4730) );
  NANDN U22058 ( .A(n21188), .B(\stack[3][41] ), .Z(n21713) );
  NANDN U22059 ( .A(n20866), .B(n21714), .Z(n21712) );
  NAND U22060 ( .A(n21715), .B(n21716), .Z(n21714) );
  NANDN U22061 ( .A(n4967), .B(\stack[4][41] ), .Z(n21716) );
  NANDN U22062 ( .A(n20875), .B(\stack[2][41] ), .Z(n21715) );
  NAND U22063 ( .A(n21717), .B(n21718), .Z(n4729) );
  NANDN U22064 ( .A(n21188), .B(\stack[3][42] ), .Z(n21718) );
  NANDN U22065 ( .A(n20866), .B(n21719), .Z(n21717) );
  NAND U22066 ( .A(n21720), .B(n21721), .Z(n21719) );
  NANDN U22067 ( .A(n4967), .B(\stack[4][42] ), .Z(n21721) );
  NANDN U22068 ( .A(n20875), .B(\stack[2][42] ), .Z(n21720) );
  NAND U22069 ( .A(n21722), .B(n21723), .Z(n4728) );
  NANDN U22070 ( .A(n21188), .B(\stack[3][43] ), .Z(n21723) );
  NANDN U22071 ( .A(n20866), .B(n21724), .Z(n21722) );
  NAND U22072 ( .A(n21725), .B(n21726), .Z(n21724) );
  NANDN U22073 ( .A(n4967), .B(\stack[4][43] ), .Z(n21726) );
  NANDN U22074 ( .A(n20875), .B(\stack[2][43] ), .Z(n21725) );
  NAND U22075 ( .A(n21727), .B(n21728), .Z(n4727) );
  NANDN U22076 ( .A(n21188), .B(\stack[3][44] ), .Z(n21728) );
  NANDN U22077 ( .A(n20866), .B(n21729), .Z(n21727) );
  NAND U22078 ( .A(n21730), .B(n21731), .Z(n21729) );
  NANDN U22079 ( .A(n4967), .B(\stack[4][44] ), .Z(n21731) );
  NANDN U22080 ( .A(n20875), .B(\stack[2][44] ), .Z(n21730) );
  NAND U22081 ( .A(n21732), .B(n21733), .Z(n4726) );
  NANDN U22082 ( .A(n21188), .B(\stack[3][45] ), .Z(n21733) );
  NANDN U22083 ( .A(n20866), .B(n21734), .Z(n21732) );
  NAND U22084 ( .A(n21735), .B(n21736), .Z(n21734) );
  NANDN U22085 ( .A(n4967), .B(\stack[4][45] ), .Z(n21736) );
  NANDN U22086 ( .A(n20875), .B(\stack[2][45] ), .Z(n21735) );
  NAND U22087 ( .A(n21737), .B(n21738), .Z(n4725) );
  NANDN U22088 ( .A(n21188), .B(\stack[3][46] ), .Z(n21738) );
  NANDN U22089 ( .A(n20866), .B(n21739), .Z(n21737) );
  NAND U22090 ( .A(n21740), .B(n21741), .Z(n21739) );
  NANDN U22091 ( .A(n4967), .B(\stack[4][46] ), .Z(n21741) );
  NANDN U22092 ( .A(n20875), .B(\stack[2][46] ), .Z(n21740) );
  NAND U22093 ( .A(n21742), .B(n21743), .Z(n4724) );
  NANDN U22094 ( .A(n21188), .B(\stack[3][47] ), .Z(n21743) );
  NANDN U22095 ( .A(n20866), .B(n21744), .Z(n21742) );
  NAND U22096 ( .A(n21745), .B(n21746), .Z(n21744) );
  NANDN U22097 ( .A(n4967), .B(\stack[4][47] ), .Z(n21746) );
  NANDN U22098 ( .A(n20875), .B(\stack[2][47] ), .Z(n21745) );
  NAND U22099 ( .A(n21747), .B(n21748), .Z(n4723) );
  NANDN U22100 ( .A(n21188), .B(\stack[3][48] ), .Z(n21748) );
  NANDN U22101 ( .A(n20866), .B(n21749), .Z(n21747) );
  NAND U22102 ( .A(n21750), .B(n21751), .Z(n21749) );
  NANDN U22103 ( .A(n4967), .B(\stack[4][48] ), .Z(n21751) );
  NANDN U22104 ( .A(n20875), .B(\stack[2][48] ), .Z(n21750) );
  NAND U22105 ( .A(n21752), .B(n21753), .Z(n4722) );
  NANDN U22106 ( .A(n21188), .B(\stack[3][49] ), .Z(n21753) );
  NANDN U22107 ( .A(n20866), .B(n21754), .Z(n21752) );
  NAND U22108 ( .A(n21755), .B(n21756), .Z(n21754) );
  NANDN U22109 ( .A(n4967), .B(\stack[4][49] ), .Z(n21756) );
  NANDN U22110 ( .A(n20875), .B(\stack[2][49] ), .Z(n21755) );
  NAND U22111 ( .A(n21757), .B(n21758), .Z(n4721) );
  NANDN U22112 ( .A(n21188), .B(\stack[3][50] ), .Z(n21758) );
  NANDN U22113 ( .A(n20866), .B(n21759), .Z(n21757) );
  NAND U22114 ( .A(n21760), .B(n21761), .Z(n21759) );
  NANDN U22115 ( .A(n4967), .B(\stack[4][50] ), .Z(n21761) );
  NANDN U22116 ( .A(n20875), .B(\stack[2][50] ), .Z(n21760) );
  NAND U22117 ( .A(n21762), .B(n21763), .Z(n4720) );
  NANDN U22118 ( .A(n21188), .B(\stack[3][51] ), .Z(n21763) );
  NANDN U22119 ( .A(n20866), .B(n21764), .Z(n21762) );
  NAND U22120 ( .A(n21765), .B(n21766), .Z(n21764) );
  NANDN U22121 ( .A(n4967), .B(\stack[4][51] ), .Z(n21766) );
  NANDN U22122 ( .A(n20875), .B(\stack[2][51] ), .Z(n21765) );
  NAND U22123 ( .A(n21767), .B(n21768), .Z(n4719) );
  NANDN U22124 ( .A(n21188), .B(\stack[3][52] ), .Z(n21768) );
  NANDN U22125 ( .A(n20866), .B(n21769), .Z(n21767) );
  NAND U22126 ( .A(n21770), .B(n21771), .Z(n21769) );
  NANDN U22127 ( .A(n4967), .B(\stack[4][52] ), .Z(n21771) );
  NANDN U22128 ( .A(n20875), .B(\stack[2][52] ), .Z(n21770) );
  NAND U22129 ( .A(n21772), .B(n21773), .Z(n4718) );
  NANDN U22130 ( .A(n21188), .B(\stack[3][53] ), .Z(n21773) );
  NANDN U22131 ( .A(n20866), .B(n21774), .Z(n21772) );
  NAND U22132 ( .A(n21775), .B(n21776), .Z(n21774) );
  NANDN U22133 ( .A(n4967), .B(\stack[4][53] ), .Z(n21776) );
  NANDN U22134 ( .A(n20875), .B(\stack[2][53] ), .Z(n21775) );
  NAND U22135 ( .A(n21777), .B(n21778), .Z(n4717) );
  NANDN U22136 ( .A(n21188), .B(\stack[3][54] ), .Z(n21778) );
  NANDN U22137 ( .A(n20866), .B(n21779), .Z(n21777) );
  NAND U22138 ( .A(n21780), .B(n21781), .Z(n21779) );
  NANDN U22139 ( .A(n4967), .B(\stack[4][54] ), .Z(n21781) );
  NANDN U22140 ( .A(n20875), .B(\stack[2][54] ), .Z(n21780) );
  NAND U22141 ( .A(n21782), .B(n21783), .Z(n4716) );
  NANDN U22142 ( .A(n21188), .B(\stack[3][55] ), .Z(n21783) );
  NANDN U22143 ( .A(n20866), .B(n21784), .Z(n21782) );
  NAND U22144 ( .A(n21785), .B(n21786), .Z(n21784) );
  NANDN U22145 ( .A(n4967), .B(\stack[4][55] ), .Z(n21786) );
  NANDN U22146 ( .A(n20875), .B(\stack[2][55] ), .Z(n21785) );
  NAND U22147 ( .A(n21787), .B(n21788), .Z(n4715) );
  NANDN U22148 ( .A(n21188), .B(\stack[3][56] ), .Z(n21788) );
  NANDN U22149 ( .A(n20866), .B(n21789), .Z(n21787) );
  NAND U22150 ( .A(n21790), .B(n21791), .Z(n21789) );
  NANDN U22151 ( .A(n4967), .B(\stack[4][56] ), .Z(n21791) );
  NANDN U22152 ( .A(n20875), .B(\stack[2][56] ), .Z(n21790) );
  NAND U22153 ( .A(n21792), .B(n21793), .Z(n4714) );
  NANDN U22154 ( .A(n21188), .B(\stack[3][57] ), .Z(n21793) );
  NANDN U22155 ( .A(n20866), .B(n21794), .Z(n21792) );
  NAND U22156 ( .A(n21795), .B(n21796), .Z(n21794) );
  NANDN U22157 ( .A(n4967), .B(\stack[4][57] ), .Z(n21796) );
  NANDN U22158 ( .A(n20875), .B(\stack[2][57] ), .Z(n21795) );
  NAND U22159 ( .A(n21797), .B(n21798), .Z(n4713) );
  NANDN U22160 ( .A(n21188), .B(\stack[3][58] ), .Z(n21798) );
  NANDN U22161 ( .A(n20866), .B(n21799), .Z(n21797) );
  NAND U22162 ( .A(n21800), .B(n21801), .Z(n21799) );
  NANDN U22163 ( .A(n4967), .B(\stack[4][58] ), .Z(n21801) );
  NANDN U22164 ( .A(n20875), .B(\stack[2][58] ), .Z(n21800) );
  NAND U22165 ( .A(n21802), .B(n21803), .Z(n4712) );
  NANDN U22166 ( .A(n21188), .B(\stack[3][59] ), .Z(n21803) );
  NANDN U22167 ( .A(n20866), .B(n21804), .Z(n21802) );
  NAND U22168 ( .A(n21805), .B(n21806), .Z(n21804) );
  NANDN U22169 ( .A(n4967), .B(\stack[4][59] ), .Z(n21806) );
  NANDN U22170 ( .A(n20875), .B(\stack[2][59] ), .Z(n21805) );
  NAND U22171 ( .A(n21807), .B(n21808), .Z(n4711) );
  NANDN U22172 ( .A(n21188), .B(\stack[3][60] ), .Z(n21808) );
  NANDN U22173 ( .A(n20866), .B(n21809), .Z(n21807) );
  NAND U22174 ( .A(n21810), .B(n21811), .Z(n21809) );
  NANDN U22175 ( .A(n4967), .B(\stack[4][60] ), .Z(n21811) );
  NANDN U22176 ( .A(n20875), .B(\stack[2][60] ), .Z(n21810) );
  NAND U22177 ( .A(n21812), .B(n21813), .Z(n4710) );
  NANDN U22178 ( .A(n21188), .B(\stack[3][61] ), .Z(n21813) );
  NANDN U22179 ( .A(n20866), .B(n21814), .Z(n21812) );
  NAND U22180 ( .A(n21815), .B(n21816), .Z(n21814) );
  NANDN U22181 ( .A(n4967), .B(\stack[4][61] ), .Z(n21816) );
  NANDN U22182 ( .A(n20875), .B(\stack[2][61] ), .Z(n21815) );
  NAND U22183 ( .A(n21817), .B(n21818), .Z(n4709) );
  NANDN U22184 ( .A(n21188), .B(\stack[3][62] ), .Z(n21818) );
  NANDN U22185 ( .A(n20866), .B(n21819), .Z(n21817) );
  NAND U22186 ( .A(n21820), .B(n21821), .Z(n21819) );
  NANDN U22187 ( .A(n4967), .B(\stack[4][62] ), .Z(n21821) );
  NANDN U22188 ( .A(n20875), .B(\stack[2][62] ), .Z(n21820) );
  NAND U22189 ( .A(n21822), .B(n21823), .Z(n4708) );
  NANDN U22190 ( .A(n21188), .B(\stack[3][63] ), .Z(n21823) );
  NANDN U22191 ( .A(n20866), .B(n21824), .Z(n21822) );
  NAND U22192 ( .A(n21825), .B(n21826), .Z(n21824) );
  NANDN U22193 ( .A(n4967), .B(\stack[4][63] ), .Z(n21826) );
  NANDN U22194 ( .A(n20875), .B(\stack[2][63] ), .Z(n21825) );
  NAND U22195 ( .A(n21827), .B(n21828), .Z(n4707) );
  NANDN U22196 ( .A(n21188), .B(\stack[4][0] ), .Z(n21828) );
  NANDN U22197 ( .A(n20866), .B(n21829), .Z(n21827) );
  NAND U22198 ( .A(n21830), .B(n21831), .Z(n21829) );
  NANDN U22199 ( .A(n4967), .B(\stack[5][0] ), .Z(n21831) );
  NANDN U22200 ( .A(n20875), .B(\stack[3][0] ), .Z(n21830) );
  NAND U22201 ( .A(n21832), .B(n21833), .Z(n4706) );
  NANDN U22202 ( .A(n21188), .B(\stack[4][1] ), .Z(n21833) );
  NANDN U22203 ( .A(n20866), .B(n21834), .Z(n21832) );
  NAND U22204 ( .A(n21835), .B(n21836), .Z(n21834) );
  NANDN U22205 ( .A(n4967), .B(\stack[5][1] ), .Z(n21836) );
  NANDN U22206 ( .A(n20875), .B(\stack[3][1] ), .Z(n21835) );
  NAND U22207 ( .A(n21837), .B(n21838), .Z(n4705) );
  NANDN U22208 ( .A(n21188), .B(\stack[4][2] ), .Z(n21838) );
  NANDN U22209 ( .A(n20866), .B(n21839), .Z(n21837) );
  NAND U22210 ( .A(n21840), .B(n21841), .Z(n21839) );
  NANDN U22211 ( .A(n4967), .B(\stack[5][2] ), .Z(n21841) );
  NANDN U22212 ( .A(n20875), .B(\stack[3][2] ), .Z(n21840) );
  NAND U22213 ( .A(n21842), .B(n21843), .Z(n4704) );
  NANDN U22214 ( .A(n21188), .B(\stack[4][3] ), .Z(n21843) );
  NANDN U22215 ( .A(n20866), .B(n21844), .Z(n21842) );
  NAND U22216 ( .A(n21845), .B(n21846), .Z(n21844) );
  NANDN U22217 ( .A(n4967), .B(\stack[5][3] ), .Z(n21846) );
  NANDN U22218 ( .A(n20875), .B(\stack[3][3] ), .Z(n21845) );
  NAND U22219 ( .A(n21847), .B(n21848), .Z(n4703) );
  NANDN U22220 ( .A(n21188), .B(\stack[4][4] ), .Z(n21848) );
  NANDN U22221 ( .A(n20866), .B(n21849), .Z(n21847) );
  NAND U22222 ( .A(n21850), .B(n21851), .Z(n21849) );
  NANDN U22223 ( .A(n4967), .B(\stack[5][4] ), .Z(n21851) );
  NANDN U22224 ( .A(n20875), .B(\stack[3][4] ), .Z(n21850) );
  NAND U22225 ( .A(n21852), .B(n21853), .Z(n4702) );
  NANDN U22226 ( .A(n21188), .B(\stack[4][5] ), .Z(n21853) );
  NANDN U22227 ( .A(n20866), .B(n21854), .Z(n21852) );
  NAND U22228 ( .A(n21855), .B(n21856), .Z(n21854) );
  NANDN U22229 ( .A(n4967), .B(\stack[5][5] ), .Z(n21856) );
  NANDN U22230 ( .A(n20875), .B(\stack[3][5] ), .Z(n21855) );
  NAND U22231 ( .A(n21857), .B(n21858), .Z(n4701) );
  NANDN U22232 ( .A(n21188), .B(\stack[4][6] ), .Z(n21858) );
  NANDN U22233 ( .A(n20866), .B(n21859), .Z(n21857) );
  NAND U22234 ( .A(n21860), .B(n21861), .Z(n21859) );
  NANDN U22235 ( .A(n4967), .B(\stack[5][6] ), .Z(n21861) );
  NANDN U22236 ( .A(n20875), .B(\stack[3][6] ), .Z(n21860) );
  NAND U22237 ( .A(n21862), .B(n21863), .Z(n4700) );
  NANDN U22238 ( .A(n21188), .B(\stack[4][7] ), .Z(n21863) );
  NANDN U22239 ( .A(n20866), .B(n21864), .Z(n21862) );
  NAND U22240 ( .A(n21865), .B(n21866), .Z(n21864) );
  NANDN U22241 ( .A(n4967), .B(\stack[5][7] ), .Z(n21866) );
  NANDN U22242 ( .A(n20875), .B(\stack[3][7] ), .Z(n21865) );
  NAND U22243 ( .A(n21867), .B(n21868), .Z(n4699) );
  NANDN U22244 ( .A(n21188), .B(\stack[4][8] ), .Z(n21868) );
  NANDN U22245 ( .A(n20866), .B(n21869), .Z(n21867) );
  NAND U22246 ( .A(n21870), .B(n21871), .Z(n21869) );
  NANDN U22247 ( .A(n4967), .B(\stack[5][8] ), .Z(n21871) );
  NANDN U22248 ( .A(n20875), .B(\stack[3][8] ), .Z(n21870) );
  NAND U22249 ( .A(n21872), .B(n21873), .Z(n4698) );
  NANDN U22250 ( .A(n21188), .B(\stack[4][9] ), .Z(n21873) );
  NANDN U22251 ( .A(n20866), .B(n21874), .Z(n21872) );
  NAND U22252 ( .A(n21875), .B(n21876), .Z(n21874) );
  NANDN U22253 ( .A(n4967), .B(\stack[5][9] ), .Z(n21876) );
  NANDN U22254 ( .A(n20875), .B(\stack[3][9] ), .Z(n21875) );
  NAND U22255 ( .A(n21877), .B(n21878), .Z(n4697) );
  NANDN U22256 ( .A(n21188), .B(\stack[4][10] ), .Z(n21878) );
  NANDN U22257 ( .A(n20866), .B(n21879), .Z(n21877) );
  NAND U22258 ( .A(n21880), .B(n21881), .Z(n21879) );
  NANDN U22259 ( .A(n4967), .B(\stack[5][10] ), .Z(n21881) );
  NANDN U22260 ( .A(n20875), .B(\stack[3][10] ), .Z(n21880) );
  NAND U22261 ( .A(n21882), .B(n21883), .Z(n4696) );
  NANDN U22262 ( .A(n21188), .B(\stack[4][11] ), .Z(n21883) );
  NANDN U22263 ( .A(n20866), .B(n21884), .Z(n21882) );
  NAND U22264 ( .A(n21885), .B(n21886), .Z(n21884) );
  NANDN U22265 ( .A(n4967), .B(\stack[5][11] ), .Z(n21886) );
  NANDN U22266 ( .A(n20875), .B(\stack[3][11] ), .Z(n21885) );
  NAND U22267 ( .A(n21887), .B(n21888), .Z(n4695) );
  NANDN U22268 ( .A(n21188), .B(\stack[4][12] ), .Z(n21888) );
  NANDN U22269 ( .A(n20866), .B(n21889), .Z(n21887) );
  NAND U22270 ( .A(n21890), .B(n21891), .Z(n21889) );
  NANDN U22271 ( .A(n4967), .B(\stack[5][12] ), .Z(n21891) );
  NANDN U22272 ( .A(n20875), .B(\stack[3][12] ), .Z(n21890) );
  NAND U22273 ( .A(n21892), .B(n21893), .Z(n4694) );
  NANDN U22274 ( .A(n21188), .B(\stack[4][13] ), .Z(n21893) );
  NANDN U22275 ( .A(n20866), .B(n21894), .Z(n21892) );
  NAND U22276 ( .A(n21895), .B(n21896), .Z(n21894) );
  NANDN U22277 ( .A(n4967), .B(\stack[5][13] ), .Z(n21896) );
  NANDN U22278 ( .A(n20875), .B(\stack[3][13] ), .Z(n21895) );
  NAND U22279 ( .A(n21897), .B(n21898), .Z(n4693) );
  NANDN U22280 ( .A(n21188), .B(\stack[4][14] ), .Z(n21898) );
  NANDN U22281 ( .A(n20866), .B(n21899), .Z(n21897) );
  NAND U22282 ( .A(n21900), .B(n21901), .Z(n21899) );
  NANDN U22283 ( .A(n4967), .B(\stack[5][14] ), .Z(n21901) );
  NANDN U22284 ( .A(n20875), .B(\stack[3][14] ), .Z(n21900) );
  NAND U22285 ( .A(n21902), .B(n21903), .Z(n4692) );
  NANDN U22286 ( .A(n21188), .B(\stack[4][15] ), .Z(n21903) );
  NANDN U22287 ( .A(n20866), .B(n21904), .Z(n21902) );
  NAND U22288 ( .A(n21905), .B(n21906), .Z(n21904) );
  NANDN U22289 ( .A(n4967), .B(\stack[5][15] ), .Z(n21906) );
  NANDN U22290 ( .A(n20875), .B(\stack[3][15] ), .Z(n21905) );
  NAND U22291 ( .A(n21907), .B(n21908), .Z(n4691) );
  NANDN U22292 ( .A(n21188), .B(\stack[4][16] ), .Z(n21908) );
  NANDN U22293 ( .A(n20866), .B(n21909), .Z(n21907) );
  NAND U22294 ( .A(n21910), .B(n21911), .Z(n21909) );
  NANDN U22295 ( .A(n4967), .B(\stack[5][16] ), .Z(n21911) );
  NANDN U22296 ( .A(n20875), .B(\stack[3][16] ), .Z(n21910) );
  NAND U22297 ( .A(n21912), .B(n21913), .Z(n4690) );
  NANDN U22298 ( .A(n21188), .B(\stack[4][17] ), .Z(n21913) );
  NANDN U22299 ( .A(n20866), .B(n21914), .Z(n21912) );
  NAND U22300 ( .A(n21915), .B(n21916), .Z(n21914) );
  NANDN U22301 ( .A(n4967), .B(\stack[5][17] ), .Z(n21916) );
  NANDN U22302 ( .A(n20875), .B(\stack[3][17] ), .Z(n21915) );
  NAND U22303 ( .A(n21917), .B(n21918), .Z(n4689) );
  NANDN U22304 ( .A(n21188), .B(\stack[4][18] ), .Z(n21918) );
  NANDN U22305 ( .A(n20866), .B(n21919), .Z(n21917) );
  NAND U22306 ( .A(n21920), .B(n21921), .Z(n21919) );
  NANDN U22307 ( .A(n4967), .B(\stack[5][18] ), .Z(n21921) );
  NANDN U22308 ( .A(n20875), .B(\stack[3][18] ), .Z(n21920) );
  NAND U22309 ( .A(n21922), .B(n21923), .Z(n4688) );
  NANDN U22310 ( .A(n21188), .B(\stack[4][19] ), .Z(n21923) );
  NANDN U22311 ( .A(n20866), .B(n21924), .Z(n21922) );
  NAND U22312 ( .A(n21925), .B(n21926), .Z(n21924) );
  NANDN U22313 ( .A(n4967), .B(\stack[5][19] ), .Z(n21926) );
  NANDN U22314 ( .A(n20875), .B(\stack[3][19] ), .Z(n21925) );
  NAND U22315 ( .A(n21927), .B(n21928), .Z(n4687) );
  NANDN U22316 ( .A(n21188), .B(\stack[4][20] ), .Z(n21928) );
  NANDN U22317 ( .A(n20866), .B(n21929), .Z(n21927) );
  NAND U22318 ( .A(n21930), .B(n21931), .Z(n21929) );
  NANDN U22319 ( .A(n4967), .B(\stack[5][20] ), .Z(n21931) );
  NANDN U22320 ( .A(n20875), .B(\stack[3][20] ), .Z(n21930) );
  NAND U22321 ( .A(n21932), .B(n21933), .Z(n4686) );
  NANDN U22322 ( .A(n21188), .B(\stack[4][21] ), .Z(n21933) );
  NANDN U22323 ( .A(n20866), .B(n21934), .Z(n21932) );
  NAND U22324 ( .A(n21935), .B(n21936), .Z(n21934) );
  NANDN U22325 ( .A(n4967), .B(\stack[5][21] ), .Z(n21936) );
  NANDN U22326 ( .A(n20875), .B(\stack[3][21] ), .Z(n21935) );
  NAND U22327 ( .A(n21937), .B(n21938), .Z(n4685) );
  NANDN U22328 ( .A(n21188), .B(\stack[4][22] ), .Z(n21938) );
  NANDN U22329 ( .A(n20866), .B(n21939), .Z(n21937) );
  NAND U22330 ( .A(n21940), .B(n21941), .Z(n21939) );
  NANDN U22331 ( .A(n4967), .B(\stack[5][22] ), .Z(n21941) );
  NANDN U22332 ( .A(n20875), .B(\stack[3][22] ), .Z(n21940) );
  NAND U22333 ( .A(n21942), .B(n21943), .Z(n4684) );
  NANDN U22334 ( .A(n21188), .B(\stack[4][23] ), .Z(n21943) );
  NANDN U22335 ( .A(n20866), .B(n21944), .Z(n21942) );
  NAND U22336 ( .A(n21945), .B(n21946), .Z(n21944) );
  NANDN U22337 ( .A(n4967), .B(\stack[5][23] ), .Z(n21946) );
  NANDN U22338 ( .A(n20875), .B(\stack[3][23] ), .Z(n21945) );
  NAND U22339 ( .A(n21947), .B(n21948), .Z(n4683) );
  NANDN U22340 ( .A(n21188), .B(\stack[4][24] ), .Z(n21948) );
  NANDN U22341 ( .A(n20866), .B(n21949), .Z(n21947) );
  NAND U22342 ( .A(n21950), .B(n21951), .Z(n21949) );
  NANDN U22343 ( .A(n4967), .B(\stack[5][24] ), .Z(n21951) );
  NANDN U22344 ( .A(n20875), .B(\stack[3][24] ), .Z(n21950) );
  NAND U22345 ( .A(n21952), .B(n21953), .Z(n4682) );
  NANDN U22346 ( .A(n21188), .B(\stack[4][25] ), .Z(n21953) );
  NANDN U22347 ( .A(n20866), .B(n21954), .Z(n21952) );
  NAND U22348 ( .A(n21955), .B(n21956), .Z(n21954) );
  NANDN U22349 ( .A(n4967), .B(\stack[5][25] ), .Z(n21956) );
  NANDN U22350 ( .A(n20875), .B(\stack[3][25] ), .Z(n21955) );
  NAND U22351 ( .A(n21957), .B(n21958), .Z(n4681) );
  NANDN U22352 ( .A(n21188), .B(\stack[4][26] ), .Z(n21958) );
  NANDN U22353 ( .A(n20866), .B(n21959), .Z(n21957) );
  NAND U22354 ( .A(n21960), .B(n21961), .Z(n21959) );
  NANDN U22355 ( .A(n4967), .B(\stack[5][26] ), .Z(n21961) );
  NANDN U22356 ( .A(n20875), .B(\stack[3][26] ), .Z(n21960) );
  NAND U22357 ( .A(n21962), .B(n21963), .Z(n4680) );
  NANDN U22358 ( .A(n21188), .B(\stack[4][27] ), .Z(n21963) );
  NANDN U22359 ( .A(n20866), .B(n21964), .Z(n21962) );
  NAND U22360 ( .A(n21965), .B(n21966), .Z(n21964) );
  NANDN U22361 ( .A(n4967), .B(\stack[5][27] ), .Z(n21966) );
  NANDN U22362 ( .A(n20875), .B(\stack[3][27] ), .Z(n21965) );
  NAND U22363 ( .A(n21967), .B(n21968), .Z(n4679) );
  NANDN U22364 ( .A(n21188), .B(\stack[4][28] ), .Z(n21968) );
  NANDN U22365 ( .A(n20866), .B(n21969), .Z(n21967) );
  NAND U22366 ( .A(n21970), .B(n21971), .Z(n21969) );
  NANDN U22367 ( .A(n4967), .B(\stack[5][28] ), .Z(n21971) );
  NANDN U22368 ( .A(n20875), .B(\stack[3][28] ), .Z(n21970) );
  NAND U22369 ( .A(n21972), .B(n21973), .Z(n4678) );
  NANDN U22370 ( .A(n21188), .B(\stack[4][29] ), .Z(n21973) );
  NANDN U22371 ( .A(n20866), .B(n21974), .Z(n21972) );
  NAND U22372 ( .A(n21975), .B(n21976), .Z(n21974) );
  NANDN U22373 ( .A(n4967), .B(\stack[5][29] ), .Z(n21976) );
  NANDN U22374 ( .A(n20875), .B(\stack[3][29] ), .Z(n21975) );
  NAND U22375 ( .A(n21977), .B(n21978), .Z(n4677) );
  NANDN U22376 ( .A(n21188), .B(\stack[4][30] ), .Z(n21978) );
  NANDN U22377 ( .A(n20866), .B(n21979), .Z(n21977) );
  NAND U22378 ( .A(n21980), .B(n21981), .Z(n21979) );
  NANDN U22379 ( .A(n4967), .B(\stack[5][30] ), .Z(n21981) );
  NANDN U22380 ( .A(n20875), .B(\stack[3][30] ), .Z(n21980) );
  NAND U22381 ( .A(n21982), .B(n21983), .Z(n4676) );
  NANDN U22382 ( .A(n21188), .B(\stack[4][31] ), .Z(n21983) );
  NANDN U22383 ( .A(n20866), .B(n21984), .Z(n21982) );
  NAND U22384 ( .A(n21985), .B(n21986), .Z(n21984) );
  NANDN U22385 ( .A(n4967), .B(\stack[5][31] ), .Z(n21986) );
  NANDN U22386 ( .A(n20875), .B(\stack[3][31] ), .Z(n21985) );
  NAND U22387 ( .A(n21987), .B(n21988), .Z(n4675) );
  NANDN U22388 ( .A(n21188), .B(\stack[4][32] ), .Z(n21988) );
  NANDN U22389 ( .A(n20866), .B(n21989), .Z(n21987) );
  NAND U22390 ( .A(n21990), .B(n21991), .Z(n21989) );
  NANDN U22391 ( .A(n4967), .B(\stack[5][32] ), .Z(n21991) );
  NANDN U22392 ( .A(n20875), .B(\stack[3][32] ), .Z(n21990) );
  NAND U22393 ( .A(n21992), .B(n21993), .Z(n4674) );
  NANDN U22394 ( .A(n21188), .B(\stack[4][33] ), .Z(n21993) );
  NANDN U22395 ( .A(n20866), .B(n21994), .Z(n21992) );
  NAND U22396 ( .A(n21995), .B(n21996), .Z(n21994) );
  NANDN U22397 ( .A(n4967), .B(\stack[5][33] ), .Z(n21996) );
  NANDN U22398 ( .A(n20875), .B(\stack[3][33] ), .Z(n21995) );
  NAND U22399 ( .A(n21997), .B(n21998), .Z(n4673) );
  NANDN U22400 ( .A(n21188), .B(\stack[4][34] ), .Z(n21998) );
  NANDN U22401 ( .A(n20866), .B(n21999), .Z(n21997) );
  NAND U22402 ( .A(n22000), .B(n22001), .Z(n21999) );
  NANDN U22403 ( .A(n4967), .B(\stack[5][34] ), .Z(n22001) );
  NANDN U22404 ( .A(n20875), .B(\stack[3][34] ), .Z(n22000) );
  NAND U22405 ( .A(n22002), .B(n22003), .Z(n4672) );
  NANDN U22406 ( .A(n21188), .B(\stack[4][35] ), .Z(n22003) );
  NANDN U22407 ( .A(n20866), .B(n22004), .Z(n22002) );
  NAND U22408 ( .A(n22005), .B(n22006), .Z(n22004) );
  NANDN U22409 ( .A(n4967), .B(\stack[5][35] ), .Z(n22006) );
  NANDN U22410 ( .A(n20875), .B(\stack[3][35] ), .Z(n22005) );
  NAND U22411 ( .A(n22007), .B(n22008), .Z(n4671) );
  NANDN U22412 ( .A(n21188), .B(\stack[4][36] ), .Z(n22008) );
  NANDN U22413 ( .A(n20866), .B(n22009), .Z(n22007) );
  NAND U22414 ( .A(n22010), .B(n22011), .Z(n22009) );
  NANDN U22415 ( .A(n4967), .B(\stack[5][36] ), .Z(n22011) );
  NANDN U22416 ( .A(n20875), .B(\stack[3][36] ), .Z(n22010) );
  NAND U22417 ( .A(n22012), .B(n22013), .Z(n4670) );
  NANDN U22418 ( .A(n21188), .B(\stack[4][37] ), .Z(n22013) );
  NANDN U22419 ( .A(n20866), .B(n22014), .Z(n22012) );
  NAND U22420 ( .A(n22015), .B(n22016), .Z(n22014) );
  NANDN U22421 ( .A(n4967), .B(\stack[5][37] ), .Z(n22016) );
  NANDN U22422 ( .A(n20875), .B(\stack[3][37] ), .Z(n22015) );
  NAND U22423 ( .A(n22017), .B(n22018), .Z(n4669) );
  NANDN U22424 ( .A(n21188), .B(\stack[4][38] ), .Z(n22018) );
  NANDN U22425 ( .A(n20866), .B(n22019), .Z(n22017) );
  NAND U22426 ( .A(n22020), .B(n22021), .Z(n22019) );
  NANDN U22427 ( .A(n4967), .B(\stack[5][38] ), .Z(n22021) );
  NANDN U22428 ( .A(n20875), .B(\stack[3][38] ), .Z(n22020) );
  NAND U22429 ( .A(n22022), .B(n22023), .Z(n4668) );
  NANDN U22430 ( .A(n21188), .B(\stack[4][39] ), .Z(n22023) );
  NANDN U22431 ( .A(n20866), .B(n22024), .Z(n22022) );
  NAND U22432 ( .A(n22025), .B(n22026), .Z(n22024) );
  NANDN U22433 ( .A(n4967), .B(\stack[5][39] ), .Z(n22026) );
  NANDN U22434 ( .A(n20875), .B(\stack[3][39] ), .Z(n22025) );
  NAND U22435 ( .A(n22027), .B(n22028), .Z(n4667) );
  NANDN U22436 ( .A(n21188), .B(\stack[4][40] ), .Z(n22028) );
  NANDN U22437 ( .A(n20866), .B(n22029), .Z(n22027) );
  NAND U22438 ( .A(n22030), .B(n22031), .Z(n22029) );
  NANDN U22439 ( .A(n4967), .B(\stack[5][40] ), .Z(n22031) );
  NANDN U22440 ( .A(n20875), .B(\stack[3][40] ), .Z(n22030) );
  NAND U22441 ( .A(n22032), .B(n22033), .Z(n4666) );
  NANDN U22442 ( .A(n21188), .B(\stack[4][41] ), .Z(n22033) );
  NANDN U22443 ( .A(n20866), .B(n22034), .Z(n22032) );
  NAND U22444 ( .A(n22035), .B(n22036), .Z(n22034) );
  NANDN U22445 ( .A(n4967), .B(\stack[5][41] ), .Z(n22036) );
  NANDN U22446 ( .A(n20875), .B(\stack[3][41] ), .Z(n22035) );
  NAND U22447 ( .A(n22037), .B(n22038), .Z(n4665) );
  NANDN U22448 ( .A(n21188), .B(\stack[4][42] ), .Z(n22038) );
  NANDN U22449 ( .A(n20866), .B(n22039), .Z(n22037) );
  NAND U22450 ( .A(n22040), .B(n22041), .Z(n22039) );
  NANDN U22451 ( .A(n4967), .B(\stack[5][42] ), .Z(n22041) );
  NANDN U22452 ( .A(n20875), .B(\stack[3][42] ), .Z(n22040) );
  NAND U22453 ( .A(n22042), .B(n22043), .Z(n4664) );
  NANDN U22454 ( .A(n21188), .B(\stack[4][43] ), .Z(n22043) );
  NANDN U22455 ( .A(n20866), .B(n22044), .Z(n22042) );
  NAND U22456 ( .A(n22045), .B(n22046), .Z(n22044) );
  NANDN U22457 ( .A(n4967), .B(\stack[5][43] ), .Z(n22046) );
  NANDN U22458 ( .A(n20875), .B(\stack[3][43] ), .Z(n22045) );
  NAND U22459 ( .A(n22047), .B(n22048), .Z(n4663) );
  NANDN U22460 ( .A(n21188), .B(\stack[4][44] ), .Z(n22048) );
  NANDN U22461 ( .A(n20866), .B(n22049), .Z(n22047) );
  NAND U22462 ( .A(n22050), .B(n22051), .Z(n22049) );
  NANDN U22463 ( .A(n4967), .B(\stack[5][44] ), .Z(n22051) );
  NANDN U22464 ( .A(n20875), .B(\stack[3][44] ), .Z(n22050) );
  NAND U22465 ( .A(n22052), .B(n22053), .Z(n4662) );
  NANDN U22466 ( .A(n21188), .B(\stack[4][45] ), .Z(n22053) );
  NANDN U22467 ( .A(n20866), .B(n22054), .Z(n22052) );
  NAND U22468 ( .A(n22055), .B(n22056), .Z(n22054) );
  NANDN U22469 ( .A(n4967), .B(\stack[5][45] ), .Z(n22056) );
  NANDN U22470 ( .A(n20875), .B(\stack[3][45] ), .Z(n22055) );
  NAND U22471 ( .A(n22057), .B(n22058), .Z(n4661) );
  NANDN U22472 ( .A(n21188), .B(\stack[4][46] ), .Z(n22058) );
  NANDN U22473 ( .A(n20866), .B(n22059), .Z(n22057) );
  NAND U22474 ( .A(n22060), .B(n22061), .Z(n22059) );
  NANDN U22475 ( .A(n4967), .B(\stack[5][46] ), .Z(n22061) );
  NANDN U22476 ( .A(n20875), .B(\stack[3][46] ), .Z(n22060) );
  NAND U22477 ( .A(n22062), .B(n22063), .Z(n4660) );
  NANDN U22478 ( .A(n21188), .B(\stack[4][47] ), .Z(n22063) );
  NANDN U22479 ( .A(n20866), .B(n22064), .Z(n22062) );
  NAND U22480 ( .A(n22065), .B(n22066), .Z(n22064) );
  NANDN U22481 ( .A(n4967), .B(\stack[5][47] ), .Z(n22066) );
  NANDN U22482 ( .A(n20875), .B(\stack[3][47] ), .Z(n22065) );
  NAND U22483 ( .A(n22067), .B(n22068), .Z(n4659) );
  NANDN U22484 ( .A(n21188), .B(\stack[4][48] ), .Z(n22068) );
  NANDN U22485 ( .A(n20866), .B(n22069), .Z(n22067) );
  NAND U22486 ( .A(n22070), .B(n22071), .Z(n22069) );
  NANDN U22487 ( .A(n4967), .B(\stack[5][48] ), .Z(n22071) );
  NANDN U22488 ( .A(n20875), .B(\stack[3][48] ), .Z(n22070) );
  NAND U22489 ( .A(n22072), .B(n22073), .Z(n4658) );
  NANDN U22490 ( .A(n21188), .B(\stack[4][49] ), .Z(n22073) );
  NANDN U22491 ( .A(n20866), .B(n22074), .Z(n22072) );
  NAND U22492 ( .A(n22075), .B(n22076), .Z(n22074) );
  NANDN U22493 ( .A(n4967), .B(\stack[5][49] ), .Z(n22076) );
  NANDN U22494 ( .A(n20875), .B(\stack[3][49] ), .Z(n22075) );
  NAND U22495 ( .A(n22077), .B(n22078), .Z(n4657) );
  NANDN U22496 ( .A(n21188), .B(\stack[4][50] ), .Z(n22078) );
  NANDN U22497 ( .A(n20866), .B(n22079), .Z(n22077) );
  NAND U22498 ( .A(n22080), .B(n22081), .Z(n22079) );
  NANDN U22499 ( .A(n4967), .B(\stack[5][50] ), .Z(n22081) );
  NANDN U22500 ( .A(n20875), .B(\stack[3][50] ), .Z(n22080) );
  NAND U22501 ( .A(n22082), .B(n22083), .Z(n4656) );
  NANDN U22502 ( .A(n21188), .B(\stack[4][51] ), .Z(n22083) );
  NANDN U22503 ( .A(n20866), .B(n22084), .Z(n22082) );
  NAND U22504 ( .A(n22085), .B(n22086), .Z(n22084) );
  NANDN U22505 ( .A(n4967), .B(\stack[5][51] ), .Z(n22086) );
  NANDN U22506 ( .A(n20875), .B(\stack[3][51] ), .Z(n22085) );
  NAND U22507 ( .A(n22087), .B(n22088), .Z(n4655) );
  NANDN U22508 ( .A(n21188), .B(\stack[4][52] ), .Z(n22088) );
  NANDN U22509 ( .A(n20866), .B(n22089), .Z(n22087) );
  NAND U22510 ( .A(n22090), .B(n22091), .Z(n22089) );
  NANDN U22511 ( .A(n4967), .B(\stack[5][52] ), .Z(n22091) );
  NANDN U22512 ( .A(n20875), .B(\stack[3][52] ), .Z(n22090) );
  NAND U22513 ( .A(n22092), .B(n22093), .Z(n4654) );
  NANDN U22514 ( .A(n21188), .B(\stack[4][53] ), .Z(n22093) );
  NANDN U22515 ( .A(n20866), .B(n22094), .Z(n22092) );
  NAND U22516 ( .A(n22095), .B(n22096), .Z(n22094) );
  NANDN U22517 ( .A(n4967), .B(\stack[5][53] ), .Z(n22096) );
  NANDN U22518 ( .A(n20875), .B(\stack[3][53] ), .Z(n22095) );
  NAND U22519 ( .A(n22097), .B(n22098), .Z(n4653) );
  NANDN U22520 ( .A(n21188), .B(\stack[4][54] ), .Z(n22098) );
  NANDN U22521 ( .A(n20866), .B(n22099), .Z(n22097) );
  NAND U22522 ( .A(n22100), .B(n22101), .Z(n22099) );
  NANDN U22523 ( .A(n4967), .B(\stack[5][54] ), .Z(n22101) );
  NANDN U22524 ( .A(n20875), .B(\stack[3][54] ), .Z(n22100) );
  NAND U22525 ( .A(n22102), .B(n22103), .Z(n4652) );
  NANDN U22526 ( .A(n21188), .B(\stack[4][55] ), .Z(n22103) );
  NANDN U22527 ( .A(n20866), .B(n22104), .Z(n22102) );
  NAND U22528 ( .A(n22105), .B(n22106), .Z(n22104) );
  NANDN U22529 ( .A(n4967), .B(\stack[5][55] ), .Z(n22106) );
  NANDN U22530 ( .A(n20875), .B(\stack[3][55] ), .Z(n22105) );
  NAND U22531 ( .A(n22107), .B(n22108), .Z(n4651) );
  NANDN U22532 ( .A(n21188), .B(\stack[4][56] ), .Z(n22108) );
  NANDN U22533 ( .A(n20866), .B(n22109), .Z(n22107) );
  NAND U22534 ( .A(n22110), .B(n22111), .Z(n22109) );
  NANDN U22535 ( .A(n4967), .B(\stack[5][56] ), .Z(n22111) );
  NANDN U22536 ( .A(n20875), .B(\stack[3][56] ), .Z(n22110) );
  NAND U22537 ( .A(n22112), .B(n22113), .Z(n4650) );
  NANDN U22538 ( .A(n21188), .B(\stack[4][57] ), .Z(n22113) );
  NANDN U22539 ( .A(n20866), .B(n22114), .Z(n22112) );
  NAND U22540 ( .A(n22115), .B(n22116), .Z(n22114) );
  NANDN U22541 ( .A(n4967), .B(\stack[5][57] ), .Z(n22116) );
  NANDN U22542 ( .A(n20875), .B(\stack[3][57] ), .Z(n22115) );
  NAND U22543 ( .A(n22117), .B(n22118), .Z(n4649) );
  NANDN U22544 ( .A(n21188), .B(\stack[4][58] ), .Z(n22118) );
  NANDN U22545 ( .A(n20866), .B(n22119), .Z(n22117) );
  NAND U22546 ( .A(n22120), .B(n22121), .Z(n22119) );
  NANDN U22547 ( .A(n4967), .B(\stack[5][58] ), .Z(n22121) );
  NANDN U22548 ( .A(n20875), .B(\stack[3][58] ), .Z(n22120) );
  NAND U22549 ( .A(n22122), .B(n22123), .Z(n4648) );
  NANDN U22550 ( .A(n21188), .B(\stack[4][59] ), .Z(n22123) );
  NANDN U22551 ( .A(n20866), .B(n22124), .Z(n22122) );
  NAND U22552 ( .A(n22125), .B(n22126), .Z(n22124) );
  NANDN U22553 ( .A(n4967), .B(\stack[5][59] ), .Z(n22126) );
  NANDN U22554 ( .A(n20875), .B(\stack[3][59] ), .Z(n22125) );
  NAND U22555 ( .A(n22127), .B(n22128), .Z(n4647) );
  NANDN U22556 ( .A(n21188), .B(\stack[4][60] ), .Z(n22128) );
  NANDN U22557 ( .A(n20866), .B(n22129), .Z(n22127) );
  NAND U22558 ( .A(n22130), .B(n22131), .Z(n22129) );
  NANDN U22559 ( .A(n4967), .B(\stack[5][60] ), .Z(n22131) );
  NANDN U22560 ( .A(n20875), .B(\stack[3][60] ), .Z(n22130) );
  NAND U22561 ( .A(n22132), .B(n22133), .Z(n4646) );
  NANDN U22562 ( .A(n21188), .B(\stack[4][61] ), .Z(n22133) );
  NANDN U22563 ( .A(n20866), .B(n22134), .Z(n22132) );
  NAND U22564 ( .A(n22135), .B(n22136), .Z(n22134) );
  NANDN U22565 ( .A(n4967), .B(\stack[5][61] ), .Z(n22136) );
  NANDN U22566 ( .A(n20875), .B(\stack[3][61] ), .Z(n22135) );
  NAND U22567 ( .A(n22137), .B(n22138), .Z(n4645) );
  NANDN U22568 ( .A(n21188), .B(\stack[4][62] ), .Z(n22138) );
  NANDN U22569 ( .A(n20866), .B(n22139), .Z(n22137) );
  NAND U22570 ( .A(n22140), .B(n22141), .Z(n22139) );
  NANDN U22571 ( .A(n4967), .B(\stack[5][62] ), .Z(n22141) );
  NANDN U22572 ( .A(n20875), .B(\stack[3][62] ), .Z(n22140) );
  NAND U22573 ( .A(n22142), .B(n22143), .Z(n4644) );
  NANDN U22574 ( .A(n21188), .B(\stack[4][63] ), .Z(n22143) );
  NANDN U22575 ( .A(n20866), .B(n22144), .Z(n22142) );
  NAND U22576 ( .A(n22145), .B(n22146), .Z(n22144) );
  NANDN U22577 ( .A(n4967), .B(\stack[5][63] ), .Z(n22146) );
  NANDN U22578 ( .A(n20875), .B(\stack[3][63] ), .Z(n22145) );
  NAND U22579 ( .A(n22147), .B(n22148), .Z(n4643) );
  NANDN U22580 ( .A(n21188), .B(\stack[5][0] ), .Z(n22148) );
  NANDN U22581 ( .A(n20866), .B(n22149), .Z(n22147) );
  NAND U22582 ( .A(n22150), .B(n22151), .Z(n22149) );
  NANDN U22583 ( .A(n4967), .B(\stack[6][0] ), .Z(n22151) );
  NANDN U22584 ( .A(n20875), .B(\stack[4][0] ), .Z(n22150) );
  NAND U22585 ( .A(n22152), .B(n22153), .Z(n4642) );
  NANDN U22586 ( .A(n21188), .B(\stack[5][1] ), .Z(n22153) );
  NANDN U22587 ( .A(n20866), .B(n22154), .Z(n22152) );
  NAND U22588 ( .A(n22155), .B(n22156), .Z(n22154) );
  NANDN U22589 ( .A(n4967), .B(\stack[6][1] ), .Z(n22156) );
  NANDN U22590 ( .A(n20875), .B(\stack[4][1] ), .Z(n22155) );
  NAND U22591 ( .A(n22157), .B(n22158), .Z(n4641) );
  NANDN U22592 ( .A(n21188), .B(\stack[5][2] ), .Z(n22158) );
  NANDN U22593 ( .A(n20866), .B(n22159), .Z(n22157) );
  NAND U22594 ( .A(n22160), .B(n22161), .Z(n22159) );
  NANDN U22595 ( .A(n4967), .B(\stack[6][2] ), .Z(n22161) );
  NANDN U22596 ( .A(n20875), .B(\stack[4][2] ), .Z(n22160) );
  NAND U22597 ( .A(n22162), .B(n22163), .Z(n4640) );
  NANDN U22598 ( .A(n21188), .B(\stack[5][3] ), .Z(n22163) );
  NANDN U22599 ( .A(n20866), .B(n22164), .Z(n22162) );
  NAND U22600 ( .A(n22165), .B(n22166), .Z(n22164) );
  NANDN U22601 ( .A(n4967), .B(\stack[6][3] ), .Z(n22166) );
  NANDN U22602 ( .A(n20875), .B(\stack[4][3] ), .Z(n22165) );
  NAND U22603 ( .A(n22167), .B(n22168), .Z(n4639) );
  NANDN U22604 ( .A(n21188), .B(\stack[5][4] ), .Z(n22168) );
  NANDN U22605 ( .A(n20866), .B(n22169), .Z(n22167) );
  NAND U22606 ( .A(n22170), .B(n22171), .Z(n22169) );
  NANDN U22607 ( .A(n4967), .B(\stack[6][4] ), .Z(n22171) );
  NANDN U22608 ( .A(n20875), .B(\stack[4][4] ), .Z(n22170) );
  NAND U22609 ( .A(n22172), .B(n22173), .Z(n4638) );
  NANDN U22610 ( .A(n21188), .B(\stack[5][5] ), .Z(n22173) );
  NANDN U22611 ( .A(n20866), .B(n22174), .Z(n22172) );
  NAND U22612 ( .A(n22175), .B(n22176), .Z(n22174) );
  NANDN U22613 ( .A(n4967), .B(\stack[6][5] ), .Z(n22176) );
  NANDN U22614 ( .A(n20875), .B(\stack[4][5] ), .Z(n22175) );
  NAND U22615 ( .A(n22177), .B(n22178), .Z(n4637) );
  NANDN U22616 ( .A(n21188), .B(\stack[5][6] ), .Z(n22178) );
  NANDN U22617 ( .A(n20866), .B(n22179), .Z(n22177) );
  NAND U22618 ( .A(n22180), .B(n22181), .Z(n22179) );
  NANDN U22619 ( .A(n4967), .B(\stack[6][6] ), .Z(n22181) );
  NANDN U22620 ( .A(n20875), .B(\stack[4][6] ), .Z(n22180) );
  NAND U22621 ( .A(n22182), .B(n22183), .Z(n4636) );
  NANDN U22622 ( .A(n21188), .B(\stack[5][7] ), .Z(n22183) );
  NANDN U22623 ( .A(n20866), .B(n22184), .Z(n22182) );
  NAND U22624 ( .A(n22185), .B(n22186), .Z(n22184) );
  NANDN U22625 ( .A(n4967), .B(\stack[6][7] ), .Z(n22186) );
  NANDN U22626 ( .A(n20875), .B(\stack[4][7] ), .Z(n22185) );
  NAND U22627 ( .A(n22187), .B(n22188), .Z(n4635) );
  NANDN U22628 ( .A(n21188), .B(\stack[5][8] ), .Z(n22188) );
  NANDN U22629 ( .A(n20866), .B(n22189), .Z(n22187) );
  NAND U22630 ( .A(n22190), .B(n22191), .Z(n22189) );
  NANDN U22631 ( .A(n4967), .B(\stack[6][8] ), .Z(n22191) );
  NANDN U22632 ( .A(n20875), .B(\stack[4][8] ), .Z(n22190) );
  NAND U22633 ( .A(n22192), .B(n22193), .Z(n4634) );
  NANDN U22634 ( .A(n21188), .B(\stack[5][9] ), .Z(n22193) );
  NANDN U22635 ( .A(n20866), .B(n22194), .Z(n22192) );
  NAND U22636 ( .A(n22195), .B(n22196), .Z(n22194) );
  NANDN U22637 ( .A(n4967), .B(\stack[6][9] ), .Z(n22196) );
  NANDN U22638 ( .A(n20875), .B(\stack[4][9] ), .Z(n22195) );
  NAND U22639 ( .A(n22197), .B(n22198), .Z(n4633) );
  NANDN U22640 ( .A(n21188), .B(\stack[5][10] ), .Z(n22198) );
  NANDN U22641 ( .A(n20866), .B(n22199), .Z(n22197) );
  NAND U22642 ( .A(n22200), .B(n22201), .Z(n22199) );
  NANDN U22643 ( .A(n4967), .B(\stack[6][10] ), .Z(n22201) );
  NANDN U22644 ( .A(n20875), .B(\stack[4][10] ), .Z(n22200) );
  NAND U22645 ( .A(n22202), .B(n22203), .Z(n4632) );
  NANDN U22646 ( .A(n21188), .B(\stack[5][11] ), .Z(n22203) );
  NANDN U22647 ( .A(n20866), .B(n22204), .Z(n22202) );
  NAND U22648 ( .A(n22205), .B(n22206), .Z(n22204) );
  NANDN U22649 ( .A(n4967), .B(\stack[6][11] ), .Z(n22206) );
  NANDN U22650 ( .A(n20875), .B(\stack[4][11] ), .Z(n22205) );
  NAND U22651 ( .A(n22207), .B(n22208), .Z(n4631) );
  NANDN U22652 ( .A(n21188), .B(\stack[5][12] ), .Z(n22208) );
  NANDN U22653 ( .A(n20866), .B(n22209), .Z(n22207) );
  NAND U22654 ( .A(n22210), .B(n22211), .Z(n22209) );
  NANDN U22655 ( .A(n4967), .B(\stack[6][12] ), .Z(n22211) );
  NANDN U22656 ( .A(n20875), .B(\stack[4][12] ), .Z(n22210) );
  NAND U22657 ( .A(n22212), .B(n22213), .Z(n4630) );
  NANDN U22658 ( .A(n21188), .B(\stack[5][13] ), .Z(n22213) );
  NANDN U22659 ( .A(n20866), .B(n22214), .Z(n22212) );
  NAND U22660 ( .A(n22215), .B(n22216), .Z(n22214) );
  NANDN U22661 ( .A(n4967), .B(\stack[6][13] ), .Z(n22216) );
  NANDN U22662 ( .A(n20875), .B(\stack[4][13] ), .Z(n22215) );
  NAND U22663 ( .A(n22217), .B(n22218), .Z(n4629) );
  NANDN U22664 ( .A(n21188), .B(\stack[5][14] ), .Z(n22218) );
  NANDN U22665 ( .A(n20866), .B(n22219), .Z(n22217) );
  NAND U22666 ( .A(n22220), .B(n22221), .Z(n22219) );
  NANDN U22667 ( .A(n4967), .B(\stack[6][14] ), .Z(n22221) );
  NANDN U22668 ( .A(n20875), .B(\stack[4][14] ), .Z(n22220) );
  NAND U22669 ( .A(n22222), .B(n22223), .Z(n4628) );
  NANDN U22670 ( .A(n21188), .B(\stack[5][15] ), .Z(n22223) );
  NANDN U22671 ( .A(n20866), .B(n22224), .Z(n22222) );
  NAND U22672 ( .A(n22225), .B(n22226), .Z(n22224) );
  NANDN U22673 ( .A(n4967), .B(\stack[6][15] ), .Z(n22226) );
  NANDN U22674 ( .A(n20875), .B(\stack[4][15] ), .Z(n22225) );
  NAND U22675 ( .A(n22227), .B(n22228), .Z(n4627) );
  NANDN U22676 ( .A(n21188), .B(\stack[5][16] ), .Z(n22228) );
  NANDN U22677 ( .A(n20866), .B(n22229), .Z(n22227) );
  NAND U22678 ( .A(n22230), .B(n22231), .Z(n22229) );
  NANDN U22679 ( .A(n4967), .B(\stack[6][16] ), .Z(n22231) );
  NANDN U22680 ( .A(n20875), .B(\stack[4][16] ), .Z(n22230) );
  NAND U22681 ( .A(n22232), .B(n22233), .Z(n4626) );
  NANDN U22682 ( .A(n21188), .B(\stack[5][17] ), .Z(n22233) );
  NANDN U22683 ( .A(n20866), .B(n22234), .Z(n22232) );
  NAND U22684 ( .A(n22235), .B(n22236), .Z(n22234) );
  NANDN U22685 ( .A(n4967), .B(\stack[6][17] ), .Z(n22236) );
  NANDN U22686 ( .A(n20875), .B(\stack[4][17] ), .Z(n22235) );
  NAND U22687 ( .A(n22237), .B(n22238), .Z(n4625) );
  NANDN U22688 ( .A(n21188), .B(\stack[5][18] ), .Z(n22238) );
  NANDN U22689 ( .A(n20866), .B(n22239), .Z(n22237) );
  NAND U22690 ( .A(n22240), .B(n22241), .Z(n22239) );
  NANDN U22691 ( .A(n4967), .B(\stack[6][18] ), .Z(n22241) );
  NANDN U22692 ( .A(n20875), .B(\stack[4][18] ), .Z(n22240) );
  NAND U22693 ( .A(n22242), .B(n22243), .Z(n4624) );
  NANDN U22694 ( .A(n21188), .B(\stack[5][19] ), .Z(n22243) );
  NANDN U22695 ( .A(n20866), .B(n22244), .Z(n22242) );
  NAND U22696 ( .A(n22245), .B(n22246), .Z(n22244) );
  NANDN U22697 ( .A(n4967), .B(\stack[6][19] ), .Z(n22246) );
  NANDN U22698 ( .A(n20875), .B(\stack[4][19] ), .Z(n22245) );
  NAND U22699 ( .A(n22247), .B(n22248), .Z(n4623) );
  NANDN U22700 ( .A(n21188), .B(\stack[5][20] ), .Z(n22248) );
  NANDN U22701 ( .A(n20866), .B(n22249), .Z(n22247) );
  NAND U22702 ( .A(n22250), .B(n22251), .Z(n22249) );
  NANDN U22703 ( .A(n4967), .B(\stack[6][20] ), .Z(n22251) );
  NANDN U22704 ( .A(n20875), .B(\stack[4][20] ), .Z(n22250) );
  NAND U22705 ( .A(n22252), .B(n22253), .Z(n4622) );
  NANDN U22706 ( .A(n21188), .B(\stack[5][21] ), .Z(n22253) );
  NANDN U22707 ( .A(n20866), .B(n22254), .Z(n22252) );
  NAND U22708 ( .A(n22255), .B(n22256), .Z(n22254) );
  NANDN U22709 ( .A(n4967), .B(\stack[6][21] ), .Z(n22256) );
  NANDN U22710 ( .A(n20875), .B(\stack[4][21] ), .Z(n22255) );
  NAND U22711 ( .A(n22257), .B(n22258), .Z(n4621) );
  NANDN U22712 ( .A(n21188), .B(\stack[5][22] ), .Z(n22258) );
  NANDN U22713 ( .A(n20866), .B(n22259), .Z(n22257) );
  NAND U22714 ( .A(n22260), .B(n22261), .Z(n22259) );
  NANDN U22715 ( .A(n4967), .B(\stack[6][22] ), .Z(n22261) );
  NANDN U22716 ( .A(n20875), .B(\stack[4][22] ), .Z(n22260) );
  NAND U22717 ( .A(n22262), .B(n22263), .Z(n4620) );
  NANDN U22718 ( .A(n21188), .B(\stack[5][23] ), .Z(n22263) );
  NANDN U22719 ( .A(n20866), .B(n22264), .Z(n22262) );
  NAND U22720 ( .A(n22265), .B(n22266), .Z(n22264) );
  NANDN U22721 ( .A(n4967), .B(\stack[6][23] ), .Z(n22266) );
  NANDN U22722 ( .A(n20875), .B(\stack[4][23] ), .Z(n22265) );
  NAND U22723 ( .A(n22267), .B(n22268), .Z(n4619) );
  NANDN U22724 ( .A(n21188), .B(\stack[5][24] ), .Z(n22268) );
  NANDN U22725 ( .A(n20866), .B(n22269), .Z(n22267) );
  NAND U22726 ( .A(n22270), .B(n22271), .Z(n22269) );
  NANDN U22727 ( .A(n4967), .B(\stack[6][24] ), .Z(n22271) );
  NANDN U22728 ( .A(n20875), .B(\stack[4][24] ), .Z(n22270) );
  NAND U22729 ( .A(n22272), .B(n22273), .Z(n4618) );
  NANDN U22730 ( .A(n21188), .B(\stack[5][25] ), .Z(n22273) );
  NANDN U22731 ( .A(n20866), .B(n22274), .Z(n22272) );
  NAND U22732 ( .A(n22275), .B(n22276), .Z(n22274) );
  NANDN U22733 ( .A(n4967), .B(\stack[6][25] ), .Z(n22276) );
  NANDN U22734 ( .A(n20875), .B(\stack[4][25] ), .Z(n22275) );
  NAND U22735 ( .A(n22277), .B(n22278), .Z(n4617) );
  NANDN U22736 ( .A(n21188), .B(\stack[5][26] ), .Z(n22278) );
  NANDN U22737 ( .A(n20866), .B(n22279), .Z(n22277) );
  NAND U22738 ( .A(n22280), .B(n22281), .Z(n22279) );
  NANDN U22739 ( .A(n4967), .B(\stack[6][26] ), .Z(n22281) );
  NANDN U22740 ( .A(n20875), .B(\stack[4][26] ), .Z(n22280) );
  NAND U22741 ( .A(n22282), .B(n22283), .Z(n4616) );
  NANDN U22742 ( .A(n21188), .B(\stack[5][27] ), .Z(n22283) );
  NANDN U22743 ( .A(n20866), .B(n22284), .Z(n22282) );
  NAND U22744 ( .A(n22285), .B(n22286), .Z(n22284) );
  NANDN U22745 ( .A(n4967), .B(\stack[6][27] ), .Z(n22286) );
  NANDN U22746 ( .A(n20875), .B(\stack[4][27] ), .Z(n22285) );
  NAND U22747 ( .A(n22287), .B(n22288), .Z(n4615) );
  NANDN U22748 ( .A(n21188), .B(\stack[5][28] ), .Z(n22288) );
  NANDN U22749 ( .A(n20866), .B(n22289), .Z(n22287) );
  NAND U22750 ( .A(n22290), .B(n22291), .Z(n22289) );
  NANDN U22751 ( .A(n4967), .B(\stack[6][28] ), .Z(n22291) );
  NANDN U22752 ( .A(n20875), .B(\stack[4][28] ), .Z(n22290) );
  NAND U22753 ( .A(n22292), .B(n22293), .Z(n4614) );
  NANDN U22754 ( .A(n21188), .B(\stack[5][29] ), .Z(n22293) );
  NANDN U22755 ( .A(n20866), .B(n22294), .Z(n22292) );
  NAND U22756 ( .A(n22295), .B(n22296), .Z(n22294) );
  NANDN U22757 ( .A(n4967), .B(\stack[6][29] ), .Z(n22296) );
  NANDN U22758 ( .A(n20875), .B(\stack[4][29] ), .Z(n22295) );
  NAND U22759 ( .A(n22297), .B(n22298), .Z(n4613) );
  NANDN U22760 ( .A(n21188), .B(\stack[5][30] ), .Z(n22298) );
  NANDN U22761 ( .A(n20866), .B(n22299), .Z(n22297) );
  NAND U22762 ( .A(n22300), .B(n22301), .Z(n22299) );
  NANDN U22763 ( .A(n4967), .B(\stack[6][30] ), .Z(n22301) );
  NANDN U22764 ( .A(n20875), .B(\stack[4][30] ), .Z(n22300) );
  NAND U22765 ( .A(n22302), .B(n22303), .Z(n4612) );
  NANDN U22766 ( .A(n21188), .B(\stack[5][31] ), .Z(n22303) );
  NANDN U22767 ( .A(n20866), .B(n22304), .Z(n22302) );
  NAND U22768 ( .A(n22305), .B(n22306), .Z(n22304) );
  NANDN U22769 ( .A(n4967), .B(\stack[6][31] ), .Z(n22306) );
  NANDN U22770 ( .A(n20875), .B(\stack[4][31] ), .Z(n22305) );
  NAND U22771 ( .A(n22307), .B(n22308), .Z(n4611) );
  NANDN U22772 ( .A(n21188), .B(\stack[5][32] ), .Z(n22308) );
  NANDN U22773 ( .A(n20866), .B(n22309), .Z(n22307) );
  NAND U22774 ( .A(n22310), .B(n22311), .Z(n22309) );
  NANDN U22775 ( .A(n4967), .B(\stack[6][32] ), .Z(n22311) );
  NANDN U22776 ( .A(n20875), .B(\stack[4][32] ), .Z(n22310) );
  NAND U22777 ( .A(n22312), .B(n22313), .Z(n4610) );
  NANDN U22778 ( .A(n21188), .B(\stack[5][33] ), .Z(n22313) );
  NANDN U22779 ( .A(n20866), .B(n22314), .Z(n22312) );
  NAND U22780 ( .A(n22315), .B(n22316), .Z(n22314) );
  NANDN U22781 ( .A(n4967), .B(\stack[6][33] ), .Z(n22316) );
  NANDN U22782 ( .A(n20875), .B(\stack[4][33] ), .Z(n22315) );
  NAND U22783 ( .A(n22317), .B(n22318), .Z(n4609) );
  NANDN U22784 ( .A(n21188), .B(\stack[5][34] ), .Z(n22318) );
  NANDN U22785 ( .A(n20866), .B(n22319), .Z(n22317) );
  NAND U22786 ( .A(n22320), .B(n22321), .Z(n22319) );
  NANDN U22787 ( .A(n4967), .B(\stack[6][34] ), .Z(n22321) );
  NANDN U22788 ( .A(n20875), .B(\stack[4][34] ), .Z(n22320) );
  NAND U22789 ( .A(n22322), .B(n22323), .Z(n4608) );
  NANDN U22790 ( .A(n21188), .B(\stack[5][35] ), .Z(n22323) );
  NANDN U22791 ( .A(n20866), .B(n22324), .Z(n22322) );
  NAND U22792 ( .A(n22325), .B(n22326), .Z(n22324) );
  NANDN U22793 ( .A(n4967), .B(\stack[6][35] ), .Z(n22326) );
  NANDN U22794 ( .A(n20875), .B(\stack[4][35] ), .Z(n22325) );
  NAND U22795 ( .A(n22327), .B(n22328), .Z(n4607) );
  NANDN U22796 ( .A(n21188), .B(\stack[5][36] ), .Z(n22328) );
  NANDN U22797 ( .A(n20866), .B(n22329), .Z(n22327) );
  NAND U22798 ( .A(n22330), .B(n22331), .Z(n22329) );
  NANDN U22799 ( .A(n4967), .B(\stack[6][36] ), .Z(n22331) );
  NANDN U22800 ( .A(n20875), .B(\stack[4][36] ), .Z(n22330) );
  NAND U22801 ( .A(n22332), .B(n22333), .Z(n4606) );
  NANDN U22802 ( .A(n21188), .B(\stack[5][37] ), .Z(n22333) );
  NANDN U22803 ( .A(n20866), .B(n22334), .Z(n22332) );
  NAND U22804 ( .A(n22335), .B(n22336), .Z(n22334) );
  NANDN U22805 ( .A(n4967), .B(\stack[6][37] ), .Z(n22336) );
  NANDN U22806 ( .A(n20875), .B(\stack[4][37] ), .Z(n22335) );
  NAND U22807 ( .A(n22337), .B(n22338), .Z(n4605) );
  NANDN U22808 ( .A(n21188), .B(\stack[5][38] ), .Z(n22338) );
  NANDN U22809 ( .A(n20866), .B(n22339), .Z(n22337) );
  NAND U22810 ( .A(n22340), .B(n22341), .Z(n22339) );
  NANDN U22811 ( .A(n4967), .B(\stack[6][38] ), .Z(n22341) );
  NANDN U22812 ( .A(n20875), .B(\stack[4][38] ), .Z(n22340) );
  NAND U22813 ( .A(n22342), .B(n22343), .Z(n4604) );
  NANDN U22814 ( .A(n21188), .B(\stack[5][39] ), .Z(n22343) );
  NANDN U22815 ( .A(n20866), .B(n22344), .Z(n22342) );
  NAND U22816 ( .A(n22345), .B(n22346), .Z(n22344) );
  NANDN U22817 ( .A(n4967), .B(\stack[6][39] ), .Z(n22346) );
  NANDN U22818 ( .A(n20875), .B(\stack[4][39] ), .Z(n22345) );
  NAND U22819 ( .A(n22347), .B(n22348), .Z(n4603) );
  NANDN U22820 ( .A(n21188), .B(\stack[5][40] ), .Z(n22348) );
  NANDN U22821 ( .A(n20866), .B(n22349), .Z(n22347) );
  NAND U22822 ( .A(n22350), .B(n22351), .Z(n22349) );
  NANDN U22823 ( .A(n4967), .B(\stack[6][40] ), .Z(n22351) );
  NANDN U22824 ( .A(n20875), .B(\stack[4][40] ), .Z(n22350) );
  NAND U22825 ( .A(n22352), .B(n22353), .Z(n4602) );
  NANDN U22826 ( .A(n21188), .B(\stack[5][41] ), .Z(n22353) );
  NANDN U22827 ( .A(n20866), .B(n22354), .Z(n22352) );
  NAND U22828 ( .A(n22355), .B(n22356), .Z(n22354) );
  NANDN U22829 ( .A(n4967), .B(\stack[6][41] ), .Z(n22356) );
  NANDN U22830 ( .A(n20875), .B(\stack[4][41] ), .Z(n22355) );
  NAND U22831 ( .A(n22357), .B(n22358), .Z(n4601) );
  NANDN U22832 ( .A(n21188), .B(\stack[5][42] ), .Z(n22358) );
  NANDN U22833 ( .A(n20866), .B(n22359), .Z(n22357) );
  NAND U22834 ( .A(n22360), .B(n22361), .Z(n22359) );
  NANDN U22835 ( .A(n4967), .B(\stack[6][42] ), .Z(n22361) );
  NANDN U22836 ( .A(n20875), .B(\stack[4][42] ), .Z(n22360) );
  NAND U22837 ( .A(n22362), .B(n22363), .Z(n4600) );
  NANDN U22838 ( .A(n21188), .B(\stack[5][43] ), .Z(n22363) );
  NANDN U22839 ( .A(n20866), .B(n22364), .Z(n22362) );
  NAND U22840 ( .A(n22365), .B(n22366), .Z(n22364) );
  NANDN U22841 ( .A(n4967), .B(\stack[6][43] ), .Z(n22366) );
  NANDN U22842 ( .A(n20875), .B(\stack[4][43] ), .Z(n22365) );
  NAND U22843 ( .A(n22367), .B(n22368), .Z(n4599) );
  NANDN U22844 ( .A(n21188), .B(\stack[5][44] ), .Z(n22368) );
  NANDN U22845 ( .A(n20866), .B(n22369), .Z(n22367) );
  NAND U22846 ( .A(n22370), .B(n22371), .Z(n22369) );
  NANDN U22847 ( .A(n4967), .B(\stack[6][44] ), .Z(n22371) );
  NANDN U22848 ( .A(n20875), .B(\stack[4][44] ), .Z(n22370) );
  NAND U22849 ( .A(n22372), .B(n22373), .Z(n4598) );
  NANDN U22850 ( .A(n21188), .B(\stack[5][45] ), .Z(n22373) );
  NANDN U22851 ( .A(n20866), .B(n22374), .Z(n22372) );
  NAND U22852 ( .A(n22375), .B(n22376), .Z(n22374) );
  NANDN U22853 ( .A(n4967), .B(\stack[6][45] ), .Z(n22376) );
  NANDN U22854 ( .A(n20875), .B(\stack[4][45] ), .Z(n22375) );
  NAND U22855 ( .A(n22377), .B(n22378), .Z(n4597) );
  NANDN U22856 ( .A(n21188), .B(\stack[5][46] ), .Z(n22378) );
  NANDN U22857 ( .A(n20866), .B(n22379), .Z(n22377) );
  NAND U22858 ( .A(n22380), .B(n22381), .Z(n22379) );
  NANDN U22859 ( .A(n4967), .B(\stack[6][46] ), .Z(n22381) );
  NANDN U22860 ( .A(n20875), .B(\stack[4][46] ), .Z(n22380) );
  NAND U22861 ( .A(n22382), .B(n22383), .Z(n4596) );
  NANDN U22862 ( .A(n21188), .B(\stack[5][47] ), .Z(n22383) );
  NANDN U22863 ( .A(n20866), .B(n22384), .Z(n22382) );
  NAND U22864 ( .A(n22385), .B(n22386), .Z(n22384) );
  NANDN U22865 ( .A(n4967), .B(\stack[6][47] ), .Z(n22386) );
  NANDN U22866 ( .A(n20875), .B(\stack[4][47] ), .Z(n22385) );
  NAND U22867 ( .A(n22387), .B(n22388), .Z(n4595) );
  NANDN U22868 ( .A(n21188), .B(\stack[5][48] ), .Z(n22388) );
  NANDN U22869 ( .A(n20866), .B(n22389), .Z(n22387) );
  NAND U22870 ( .A(n22390), .B(n22391), .Z(n22389) );
  NANDN U22871 ( .A(n4967), .B(\stack[6][48] ), .Z(n22391) );
  NANDN U22872 ( .A(n20875), .B(\stack[4][48] ), .Z(n22390) );
  NAND U22873 ( .A(n22392), .B(n22393), .Z(n4594) );
  NANDN U22874 ( .A(n21188), .B(\stack[5][49] ), .Z(n22393) );
  NANDN U22875 ( .A(n20866), .B(n22394), .Z(n22392) );
  NAND U22876 ( .A(n22395), .B(n22396), .Z(n22394) );
  NANDN U22877 ( .A(n4967), .B(\stack[6][49] ), .Z(n22396) );
  NANDN U22878 ( .A(n20875), .B(\stack[4][49] ), .Z(n22395) );
  NAND U22879 ( .A(n22397), .B(n22398), .Z(n4593) );
  NANDN U22880 ( .A(n21188), .B(\stack[5][50] ), .Z(n22398) );
  NANDN U22881 ( .A(n20866), .B(n22399), .Z(n22397) );
  NAND U22882 ( .A(n22400), .B(n22401), .Z(n22399) );
  NANDN U22883 ( .A(n4967), .B(\stack[6][50] ), .Z(n22401) );
  NANDN U22884 ( .A(n20875), .B(\stack[4][50] ), .Z(n22400) );
  NAND U22885 ( .A(n22402), .B(n22403), .Z(n4592) );
  NANDN U22886 ( .A(n21188), .B(\stack[5][51] ), .Z(n22403) );
  NANDN U22887 ( .A(n20866), .B(n22404), .Z(n22402) );
  NAND U22888 ( .A(n22405), .B(n22406), .Z(n22404) );
  NANDN U22889 ( .A(n4967), .B(\stack[6][51] ), .Z(n22406) );
  NANDN U22890 ( .A(n20875), .B(\stack[4][51] ), .Z(n22405) );
  NAND U22891 ( .A(n22407), .B(n22408), .Z(n4591) );
  NANDN U22892 ( .A(n21188), .B(\stack[5][52] ), .Z(n22408) );
  NANDN U22893 ( .A(n20866), .B(n22409), .Z(n22407) );
  NAND U22894 ( .A(n22410), .B(n22411), .Z(n22409) );
  NANDN U22895 ( .A(n4967), .B(\stack[6][52] ), .Z(n22411) );
  NANDN U22896 ( .A(n20875), .B(\stack[4][52] ), .Z(n22410) );
  NAND U22897 ( .A(n22412), .B(n22413), .Z(n4590) );
  NANDN U22898 ( .A(n21188), .B(\stack[5][53] ), .Z(n22413) );
  NANDN U22899 ( .A(n20866), .B(n22414), .Z(n22412) );
  NAND U22900 ( .A(n22415), .B(n22416), .Z(n22414) );
  NANDN U22901 ( .A(n4967), .B(\stack[6][53] ), .Z(n22416) );
  NANDN U22902 ( .A(n20875), .B(\stack[4][53] ), .Z(n22415) );
  NAND U22903 ( .A(n22417), .B(n22418), .Z(n4589) );
  NANDN U22904 ( .A(n21188), .B(\stack[5][54] ), .Z(n22418) );
  NANDN U22905 ( .A(n20866), .B(n22419), .Z(n22417) );
  NAND U22906 ( .A(n22420), .B(n22421), .Z(n22419) );
  NANDN U22907 ( .A(n4967), .B(\stack[6][54] ), .Z(n22421) );
  NANDN U22908 ( .A(n20875), .B(\stack[4][54] ), .Z(n22420) );
  NAND U22909 ( .A(n22422), .B(n22423), .Z(n4588) );
  NANDN U22910 ( .A(n21188), .B(\stack[5][55] ), .Z(n22423) );
  NANDN U22911 ( .A(n20866), .B(n22424), .Z(n22422) );
  NAND U22912 ( .A(n22425), .B(n22426), .Z(n22424) );
  NANDN U22913 ( .A(n4967), .B(\stack[6][55] ), .Z(n22426) );
  NANDN U22914 ( .A(n20875), .B(\stack[4][55] ), .Z(n22425) );
  NAND U22915 ( .A(n22427), .B(n22428), .Z(n4587) );
  NANDN U22916 ( .A(n21188), .B(\stack[5][56] ), .Z(n22428) );
  NANDN U22917 ( .A(n20866), .B(n22429), .Z(n22427) );
  NAND U22918 ( .A(n22430), .B(n22431), .Z(n22429) );
  NANDN U22919 ( .A(n4967), .B(\stack[6][56] ), .Z(n22431) );
  NANDN U22920 ( .A(n20875), .B(\stack[4][56] ), .Z(n22430) );
  NAND U22921 ( .A(n22432), .B(n22433), .Z(n4586) );
  NANDN U22922 ( .A(n21188), .B(\stack[5][57] ), .Z(n22433) );
  NANDN U22923 ( .A(n20866), .B(n22434), .Z(n22432) );
  NAND U22924 ( .A(n22435), .B(n22436), .Z(n22434) );
  NANDN U22925 ( .A(n4967), .B(\stack[6][57] ), .Z(n22436) );
  NANDN U22926 ( .A(n20875), .B(\stack[4][57] ), .Z(n22435) );
  NAND U22927 ( .A(n22437), .B(n22438), .Z(n4585) );
  NANDN U22928 ( .A(n21188), .B(\stack[5][58] ), .Z(n22438) );
  NANDN U22929 ( .A(n20866), .B(n22439), .Z(n22437) );
  NAND U22930 ( .A(n22440), .B(n22441), .Z(n22439) );
  NANDN U22931 ( .A(n4967), .B(\stack[6][58] ), .Z(n22441) );
  NANDN U22932 ( .A(n20875), .B(\stack[4][58] ), .Z(n22440) );
  NAND U22933 ( .A(n22442), .B(n22443), .Z(n4584) );
  NANDN U22934 ( .A(n21188), .B(\stack[5][59] ), .Z(n22443) );
  NANDN U22935 ( .A(n20866), .B(n22444), .Z(n22442) );
  NAND U22936 ( .A(n22445), .B(n22446), .Z(n22444) );
  NANDN U22937 ( .A(n4967), .B(\stack[6][59] ), .Z(n22446) );
  NANDN U22938 ( .A(n20875), .B(\stack[4][59] ), .Z(n22445) );
  NAND U22939 ( .A(n22447), .B(n22448), .Z(n4583) );
  NANDN U22940 ( .A(n21188), .B(\stack[5][60] ), .Z(n22448) );
  NANDN U22941 ( .A(n20866), .B(n22449), .Z(n22447) );
  NAND U22942 ( .A(n22450), .B(n22451), .Z(n22449) );
  NANDN U22943 ( .A(n4967), .B(\stack[6][60] ), .Z(n22451) );
  NANDN U22944 ( .A(n20875), .B(\stack[4][60] ), .Z(n22450) );
  NAND U22945 ( .A(n22452), .B(n22453), .Z(n4582) );
  NANDN U22946 ( .A(n21188), .B(\stack[5][61] ), .Z(n22453) );
  NANDN U22947 ( .A(n20866), .B(n22454), .Z(n22452) );
  NAND U22948 ( .A(n22455), .B(n22456), .Z(n22454) );
  NANDN U22949 ( .A(n4967), .B(\stack[6][61] ), .Z(n22456) );
  NANDN U22950 ( .A(n20875), .B(\stack[4][61] ), .Z(n22455) );
  NAND U22951 ( .A(n22457), .B(n22458), .Z(n4581) );
  NANDN U22952 ( .A(n21188), .B(\stack[5][62] ), .Z(n22458) );
  NANDN U22953 ( .A(n20866), .B(n22459), .Z(n22457) );
  NAND U22954 ( .A(n22460), .B(n22461), .Z(n22459) );
  NANDN U22955 ( .A(n4967), .B(\stack[6][62] ), .Z(n22461) );
  NANDN U22956 ( .A(n20875), .B(\stack[4][62] ), .Z(n22460) );
  NAND U22957 ( .A(n22462), .B(n22463), .Z(n4580) );
  NANDN U22958 ( .A(n21188), .B(\stack[5][63] ), .Z(n22463) );
  NANDN U22959 ( .A(n20866), .B(n22464), .Z(n22462) );
  NAND U22960 ( .A(n22465), .B(n22466), .Z(n22464) );
  NANDN U22961 ( .A(n4967), .B(\stack[6][63] ), .Z(n22466) );
  NANDN U22962 ( .A(n20875), .B(\stack[4][63] ), .Z(n22465) );
  NAND U22963 ( .A(n22467), .B(n22468), .Z(n4579) );
  NANDN U22964 ( .A(n21188), .B(\stack[6][0] ), .Z(n22468) );
  NANDN U22965 ( .A(n20866), .B(n22469), .Z(n22467) );
  NANDN U22966 ( .A(n22470), .B(n22471), .Z(n22469) );
  NANDN U22967 ( .A(n20875), .B(\stack[5][0] ), .Z(n22471) );
  NAND U22968 ( .A(n22472), .B(n22473), .Z(n4578) );
  NANDN U22969 ( .A(n21188), .B(\stack[6][1] ), .Z(n22473) );
  NANDN U22970 ( .A(n20866), .B(n22474), .Z(n22472) );
  NANDN U22971 ( .A(n22475), .B(n22476), .Z(n22474) );
  NANDN U22972 ( .A(n20875), .B(\stack[5][1] ), .Z(n22476) );
  NAND U22973 ( .A(n22477), .B(n22478), .Z(n4577) );
  NANDN U22974 ( .A(n21188), .B(\stack[6][2] ), .Z(n22478) );
  NANDN U22975 ( .A(n20866), .B(n22479), .Z(n22477) );
  NANDN U22976 ( .A(n22480), .B(n22481), .Z(n22479) );
  NANDN U22977 ( .A(n20875), .B(\stack[5][2] ), .Z(n22481) );
  NAND U22978 ( .A(n22482), .B(n22483), .Z(n4576) );
  NANDN U22979 ( .A(n21188), .B(\stack[6][3] ), .Z(n22483) );
  NANDN U22980 ( .A(n20866), .B(n22484), .Z(n22482) );
  NANDN U22981 ( .A(n22485), .B(n22486), .Z(n22484) );
  NANDN U22982 ( .A(n20875), .B(\stack[5][3] ), .Z(n22486) );
  NAND U22983 ( .A(n22487), .B(n22488), .Z(n4575) );
  NANDN U22984 ( .A(n21188), .B(\stack[6][4] ), .Z(n22488) );
  NANDN U22985 ( .A(n20866), .B(n22489), .Z(n22487) );
  NANDN U22986 ( .A(n22490), .B(n22491), .Z(n22489) );
  NANDN U22987 ( .A(n20875), .B(\stack[5][4] ), .Z(n22491) );
  NAND U22988 ( .A(n22492), .B(n22493), .Z(n4574) );
  NANDN U22989 ( .A(n21188), .B(\stack[6][5] ), .Z(n22493) );
  NANDN U22990 ( .A(n20866), .B(n22494), .Z(n22492) );
  NANDN U22991 ( .A(n22495), .B(n22496), .Z(n22494) );
  NANDN U22992 ( .A(n20875), .B(\stack[5][5] ), .Z(n22496) );
  NAND U22993 ( .A(n22497), .B(n22498), .Z(n4573) );
  NANDN U22994 ( .A(n21188), .B(\stack[6][6] ), .Z(n22498) );
  NANDN U22995 ( .A(n20866), .B(n22499), .Z(n22497) );
  NANDN U22996 ( .A(n22500), .B(n22501), .Z(n22499) );
  NANDN U22997 ( .A(n20875), .B(\stack[5][6] ), .Z(n22501) );
  NAND U22998 ( .A(n22502), .B(n22503), .Z(n4572) );
  NANDN U22999 ( .A(n21188), .B(\stack[6][7] ), .Z(n22503) );
  NANDN U23000 ( .A(n20866), .B(n22504), .Z(n22502) );
  NANDN U23001 ( .A(n22505), .B(n22506), .Z(n22504) );
  NANDN U23002 ( .A(n20875), .B(\stack[5][7] ), .Z(n22506) );
  NAND U23003 ( .A(n22507), .B(n22508), .Z(n4571) );
  NANDN U23004 ( .A(n21188), .B(\stack[6][8] ), .Z(n22508) );
  NANDN U23005 ( .A(n20866), .B(n22509), .Z(n22507) );
  NANDN U23006 ( .A(n22510), .B(n22511), .Z(n22509) );
  NANDN U23007 ( .A(n20875), .B(\stack[5][8] ), .Z(n22511) );
  NAND U23008 ( .A(n22512), .B(n22513), .Z(n4570) );
  NANDN U23009 ( .A(n21188), .B(\stack[6][9] ), .Z(n22513) );
  NANDN U23010 ( .A(n20866), .B(n22514), .Z(n22512) );
  NANDN U23011 ( .A(n22515), .B(n22516), .Z(n22514) );
  NANDN U23012 ( .A(n20875), .B(\stack[5][9] ), .Z(n22516) );
  NAND U23013 ( .A(n22517), .B(n22518), .Z(n4569) );
  NANDN U23014 ( .A(n21188), .B(\stack[6][10] ), .Z(n22518) );
  NANDN U23015 ( .A(n20866), .B(n22519), .Z(n22517) );
  NANDN U23016 ( .A(n22520), .B(n22521), .Z(n22519) );
  NANDN U23017 ( .A(n20875), .B(\stack[5][10] ), .Z(n22521) );
  NAND U23018 ( .A(n22522), .B(n22523), .Z(n4568) );
  NANDN U23019 ( .A(n21188), .B(\stack[6][11] ), .Z(n22523) );
  NANDN U23020 ( .A(n20866), .B(n22524), .Z(n22522) );
  NANDN U23021 ( .A(n22525), .B(n22526), .Z(n22524) );
  NANDN U23022 ( .A(n20875), .B(\stack[5][11] ), .Z(n22526) );
  NAND U23023 ( .A(n22527), .B(n22528), .Z(n4567) );
  NANDN U23024 ( .A(n21188), .B(\stack[6][12] ), .Z(n22528) );
  NANDN U23025 ( .A(n20866), .B(n22529), .Z(n22527) );
  NANDN U23026 ( .A(n22530), .B(n22531), .Z(n22529) );
  NANDN U23027 ( .A(n20875), .B(\stack[5][12] ), .Z(n22531) );
  NAND U23028 ( .A(n22532), .B(n22533), .Z(n4566) );
  NANDN U23029 ( .A(n21188), .B(\stack[6][13] ), .Z(n22533) );
  NANDN U23030 ( .A(n20866), .B(n22534), .Z(n22532) );
  NANDN U23031 ( .A(n22535), .B(n22536), .Z(n22534) );
  NANDN U23032 ( .A(n20875), .B(\stack[5][13] ), .Z(n22536) );
  NAND U23033 ( .A(n22537), .B(n22538), .Z(n4565) );
  NANDN U23034 ( .A(n21188), .B(\stack[6][14] ), .Z(n22538) );
  NANDN U23035 ( .A(n20866), .B(n22539), .Z(n22537) );
  NANDN U23036 ( .A(n22540), .B(n22541), .Z(n22539) );
  NANDN U23037 ( .A(n20875), .B(\stack[5][14] ), .Z(n22541) );
  NAND U23038 ( .A(n22542), .B(n22543), .Z(n4564) );
  NANDN U23039 ( .A(n21188), .B(\stack[6][15] ), .Z(n22543) );
  NANDN U23040 ( .A(n20866), .B(n22544), .Z(n22542) );
  NANDN U23041 ( .A(n22545), .B(n22546), .Z(n22544) );
  NANDN U23042 ( .A(n20875), .B(\stack[5][15] ), .Z(n22546) );
  NAND U23043 ( .A(n22547), .B(n22548), .Z(n4563) );
  NANDN U23044 ( .A(n21188), .B(\stack[6][16] ), .Z(n22548) );
  NANDN U23045 ( .A(n20866), .B(n22549), .Z(n22547) );
  NANDN U23046 ( .A(n22550), .B(n22551), .Z(n22549) );
  NANDN U23047 ( .A(n20875), .B(\stack[5][16] ), .Z(n22551) );
  NAND U23048 ( .A(n22552), .B(n22553), .Z(n4562) );
  NANDN U23049 ( .A(n21188), .B(\stack[6][17] ), .Z(n22553) );
  NANDN U23050 ( .A(n20866), .B(n22554), .Z(n22552) );
  NANDN U23051 ( .A(n22555), .B(n22556), .Z(n22554) );
  NANDN U23052 ( .A(n20875), .B(\stack[5][17] ), .Z(n22556) );
  NAND U23053 ( .A(n22557), .B(n22558), .Z(n4561) );
  NANDN U23054 ( .A(n21188), .B(\stack[6][18] ), .Z(n22558) );
  NANDN U23055 ( .A(n20866), .B(n22559), .Z(n22557) );
  NANDN U23056 ( .A(n22560), .B(n22561), .Z(n22559) );
  NANDN U23057 ( .A(n20875), .B(\stack[5][18] ), .Z(n22561) );
  NAND U23058 ( .A(n22562), .B(n22563), .Z(n4560) );
  NANDN U23059 ( .A(n21188), .B(\stack[6][19] ), .Z(n22563) );
  NANDN U23060 ( .A(n20866), .B(n22564), .Z(n22562) );
  NANDN U23061 ( .A(n22565), .B(n22566), .Z(n22564) );
  NANDN U23062 ( .A(n20875), .B(\stack[5][19] ), .Z(n22566) );
  NAND U23063 ( .A(n22567), .B(n22568), .Z(n4559) );
  NANDN U23064 ( .A(n21188), .B(\stack[6][20] ), .Z(n22568) );
  NANDN U23065 ( .A(n20866), .B(n22569), .Z(n22567) );
  NANDN U23066 ( .A(n22570), .B(n22571), .Z(n22569) );
  NANDN U23067 ( .A(n20875), .B(\stack[5][20] ), .Z(n22571) );
  NAND U23068 ( .A(n22572), .B(n22573), .Z(n4558) );
  NANDN U23069 ( .A(n21188), .B(\stack[6][21] ), .Z(n22573) );
  NANDN U23070 ( .A(n20866), .B(n22574), .Z(n22572) );
  NANDN U23071 ( .A(n22575), .B(n22576), .Z(n22574) );
  NANDN U23072 ( .A(n20875), .B(\stack[5][21] ), .Z(n22576) );
  NAND U23073 ( .A(n22577), .B(n22578), .Z(n4557) );
  NANDN U23074 ( .A(n21188), .B(\stack[6][22] ), .Z(n22578) );
  NANDN U23075 ( .A(n20866), .B(n22579), .Z(n22577) );
  NANDN U23076 ( .A(n22580), .B(n22581), .Z(n22579) );
  NANDN U23077 ( .A(n20875), .B(\stack[5][22] ), .Z(n22581) );
  NAND U23078 ( .A(n22582), .B(n22583), .Z(n4556) );
  NANDN U23079 ( .A(n21188), .B(\stack[6][23] ), .Z(n22583) );
  NANDN U23080 ( .A(n20866), .B(n22584), .Z(n22582) );
  NANDN U23081 ( .A(n22585), .B(n22586), .Z(n22584) );
  NANDN U23082 ( .A(n20875), .B(\stack[5][23] ), .Z(n22586) );
  NAND U23083 ( .A(n22587), .B(n22588), .Z(n4555) );
  NANDN U23084 ( .A(n21188), .B(\stack[6][24] ), .Z(n22588) );
  NANDN U23085 ( .A(n20866), .B(n22589), .Z(n22587) );
  NANDN U23086 ( .A(n22590), .B(n22591), .Z(n22589) );
  NANDN U23087 ( .A(n20875), .B(\stack[5][24] ), .Z(n22591) );
  NAND U23088 ( .A(n22592), .B(n22593), .Z(n4554) );
  NANDN U23089 ( .A(n21188), .B(\stack[6][25] ), .Z(n22593) );
  NANDN U23090 ( .A(n20866), .B(n22594), .Z(n22592) );
  NANDN U23091 ( .A(n22595), .B(n22596), .Z(n22594) );
  NANDN U23092 ( .A(n20875), .B(\stack[5][25] ), .Z(n22596) );
  NAND U23093 ( .A(n22597), .B(n22598), .Z(n4553) );
  NANDN U23094 ( .A(n21188), .B(\stack[6][26] ), .Z(n22598) );
  NANDN U23095 ( .A(n20866), .B(n22599), .Z(n22597) );
  NANDN U23096 ( .A(n22600), .B(n22601), .Z(n22599) );
  NANDN U23097 ( .A(n20875), .B(\stack[5][26] ), .Z(n22601) );
  NAND U23098 ( .A(n22602), .B(n22603), .Z(n4552) );
  NANDN U23099 ( .A(n21188), .B(\stack[6][27] ), .Z(n22603) );
  NANDN U23100 ( .A(n20866), .B(n22604), .Z(n22602) );
  NANDN U23101 ( .A(n22605), .B(n22606), .Z(n22604) );
  NANDN U23102 ( .A(n20875), .B(\stack[5][27] ), .Z(n22606) );
  NAND U23103 ( .A(n22607), .B(n22608), .Z(n4551) );
  NANDN U23104 ( .A(n21188), .B(\stack[6][28] ), .Z(n22608) );
  NANDN U23105 ( .A(n20866), .B(n22609), .Z(n22607) );
  NANDN U23106 ( .A(n22610), .B(n22611), .Z(n22609) );
  NANDN U23107 ( .A(n20875), .B(\stack[5][28] ), .Z(n22611) );
  NAND U23108 ( .A(n22612), .B(n22613), .Z(n4550) );
  NANDN U23109 ( .A(n21188), .B(\stack[6][29] ), .Z(n22613) );
  NANDN U23110 ( .A(n20866), .B(n22614), .Z(n22612) );
  NANDN U23111 ( .A(n22615), .B(n22616), .Z(n22614) );
  NANDN U23112 ( .A(n20875), .B(\stack[5][29] ), .Z(n22616) );
  NAND U23113 ( .A(n22617), .B(n22618), .Z(n4549) );
  NANDN U23114 ( .A(n21188), .B(\stack[6][30] ), .Z(n22618) );
  NANDN U23115 ( .A(n20866), .B(n22619), .Z(n22617) );
  NANDN U23116 ( .A(n22620), .B(n22621), .Z(n22619) );
  NANDN U23117 ( .A(n20875), .B(\stack[5][30] ), .Z(n22621) );
  NAND U23118 ( .A(n22622), .B(n22623), .Z(n4548) );
  NANDN U23119 ( .A(n21188), .B(\stack[6][31] ), .Z(n22623) );
  NANDN U23120 ( .A(n20866), .B(n22624), .Z(n22622) );
  NANDN U23121 ( .A(n22625), .B(n22626), .Z(n22624) );
  NANDN U23122 ( .A(n20875), .B(\stack[5][31] ), .Z(n22626) );
  NAND U23123 ( .A(n22627), .B(n22628), .Z(n4547) );
  NANDN U23124 ( .A(n21188), .B(\stack[6][32] ), .Z(n22628) );
  NANDN U23125 ( .A(n20866), .B(n22629), .Z(n22627) );
  NANDN U23126 ( .A(n22630), .B(n22631), .Z(n22629) );
  NANDN U23127 ( .A(n20875), .B(\stack[5][32] ), .Z(n22631) );
  NAND U23128 ( .A(n22632), .B(n22633), .Z(n4546) );
  NANDN U23129 ( .A(n21188), .B(\stack[6][33] ), .Z(n22633) );
  NANDN U23130 ( .A(n20866), .B(n22634), .Z(n22632) );
  NANDN U23131 ( .A(n22635), .B(n22636), .Z(n22634) );
  NANDN U23132 ( .A(n20875), .B(\stack[5][33] ), .Z(n22636) );
  NAND U23133 ( .A(n22637), .B(n22638), .Z(n4545) );
  NANDN U23134 ( .A(n21188), .B(\stack[6][34] ), .Z(n22638) );
  NANDN U23135 ( .A(n20866), .B(n22639), .Z(n22637) );
  NANDN U23136 ( .A(n22640), .B(n22641), .Z(n22639) );
  NANDN U23137 ( .A(n20875), .B(\stack[5][34] ), .Z(n22641) );
  NAND U23138 ( .A(n22642), .B(n22643), .Z(n4544) );
  NANDN U23139 ( .A(n21188), .B(\stack[6][35] ), .Z(n22643) );
  NANDN U23140 ( .A(n20866), .B(n22644), .Z(n22642) );
  NANDN U23141 ( .A(n22645), .B(n22646), .Z(n22644) );
  NANDN U23142 ( .A(n20875), .B(\stack[5][35] ), .Z(n22646) );
  NAND U23143 ( .A(n22647), .B(n22648), .Z(n4543) );
  NANDN U23144 ( .A(n21188), .B(\stack[6][36] ), .Z(n22648) );
  NANDN U23145 ( .A(n20866), .B(n22649), .Z(n22647) );
  NANDN U23146 ( .A(n22650), .B(n22651), .Z(n22649) );
  NANDN U23147 ( .A(n20875), .B(\stack[5][36] ), .Z(n22651) );
  NAND U23148 ( .A(n22652), .B(n22653), .Z(n4542) );
  NANDN U23149 ( .A(n21188), .B(\stack[6][37] ), .Z(n22653) );
  NANDN U23150 ( .A(n20866), .B(n22654), .Z(n22652) );
  NANDN U23151 ( .A(n22655), .B(n22656), .Z(n22654) );
  NANDN U23152 ( .A(n20875), .B(\stack[5][37] ), .Z(n22656) );
  NAND U23153 ( .A(n22657), .B(n22658), .Z(n4541) );
  NANDN U23154 ( .A(n21188), .B(\stack[6][38] ), .Z(n22658) );
  NANDN U23155 ( .A(n20866), .B(n22659), .Z(n22657) );
  NANDN U23156 ( .A(n22660), .B(n22661), .Z(n22659) );
  NANDN U23157 ( .A(n20875), .B(\stack[5][38] ), .Z(n22661) );
  NAND U23158 ( .A(n22662), .B(n22663), .Z(n4540) );
  NANDN U23159 ( .A(n21188), .B(\stack[6][39] ), .Z(n22663) );
  NANDN U23160 ( .A(n20866), .B(n22664), .Z(n22662) );
  NANDN U23161 ( .A(n22665), .B(n22666), .Z(n22664) );
  NANDN U23162 ( .A(n20875), .B(\stack[5][39] ), .Z(n22666) );
  NAND U23163 ( .A(n22667), .B(n22668), .Z(n4539) );
  NANDN U23164 ( .A(n21188), .B(\stack[6][40] ), .Z(n22668) );
  NANDN U23165 ( .A(n20866), .B(n22669), .Z(n22667) );
  NANDN U23166 ( .A(n22670), .B(n22671), .Z(n22669) );
  NANDN U23167 ( .A(n20875), .B(\stack[5][40] ), .Z(n22671) );
  NAND U23168 ( .A(n22672), .B(n22673), .Z(n4538) );
  NANDN U23169 ( .A(n21188), .B(\stack[6][41] ), .Z(n22673) );
  NANDN U23170 ( .A(n20866), .B(n22674), .Z(n22672) );
  NANDN U23171 ( .A(n22675), .B(n22676), .Z(n22674) );
  NANDN U23172 ( .A(n20875), .B(\stack[5][41] ), .Z(n22676) );
  NAND U23173 ( .A(n22677), .B(n22678), .Z(n4537) );
  NANDN U23174 ( .A(n21188), .B(\stack[6][42] ), .Z(n22678) );
  NANDN U23175 ( .A(n20866), .B(n22679), .Z(n22677) );
  NANDN U23176 ( .A(n22680), .B(n22681), .Z(n22679) );
  NANDN U23177 ( .A(n20875), .B(\stack[5][42] ), .Z(n22681) );
  NAND U23178 ( .A(n22682), .B(n22683), .Z(n4536) );
  NANDN U23179 ( .A(n21188), .B(\stack[6][43] ), .Z(n22683) );
  NANDN U23180 ( .A(n20866), .B(n22684), .Z(n22682) );
  NANDN U23181 ( .A(n22685), .B(n22686), .Z(n22684) );
  NANDN U23182 ( .A(n20875), .B(\stack[5][43] ), .Z(n22686) );
  NAND U23183 ( .A(n22687), .B(n22688), .Z(n4535) );
  NANDN U23184 ( .A(n21188), .B(\stack[6][44] ), .Z(n22688) );
  NANDN U23185 ( .A(n20866), .B(n22689), .Z(n22687) );
  NANDN U23186 ( .A(n22690), .B(n22691), .Z(n22689) );
  NANDN U23187 ( .A(n20875), .B(\stack[5][44] ), .Z(n22691) );
  NAND U23188 ( .A(n22692), .B(n22693), .Z(n4534) );
  NANDN U23189 ( .A(n21188), .B(\stack[6][45] ), .Z(n22693) );
  NANDN U23190 ( .A(n20866), .B(n22694), .Z(n22692) );
  NANDN U23191 ( .A(n22695), .B(n22696), .Z(n22694) );
  NANDN U23192 ( .A(n20875), .B(\stack[5][45] ), .Z(n22696) );
  NAND U23193 ( .A(n22697), .B(n22698), .Z(n4533) );
  NANDN U23194 ( .A(n21188), .B(\stack[6][46] ), .Z(n22698) );
  NANDN U23195 ( .A(n20866), .B(n22699), .Z(n22697) );
  NANDN U23196 ( .A(n22700), .B(n22701), .Z(n22699) );
  NANDN U23197 ( .A(n20875), .B(\stack[5][46] ), .Z(n22701) );
  NAND U23198 ( .A(n22702), .B(n22703), .Z(n4532) );
  NANDN U23199 ( .A(n21188), .B(\stack[6][47] ), .Z(n22703) );
  NANDN U23200 ( .A(n20866), .B(n22704), .Z(n22702) );
  NANDN U23201 ( .A(n22705), .B(n22706), .Z(n22704) );
  NANDN U23202 ( .A(n20875), .B(\stack[5][47] ), .Z(n22706) );
  NAND U23203 ( .A(n22707), .B(n22708), .Z(n4531) );
  NANDN U23204 ( .A(n21188), .B(\stack[6][48] ), .Z(n22708) );
  NANDN U23205 ( .A(n20866), .B(n22709), .Z(n22707) );
  NANDN U23206 ( .A(n22710), .B(n22711), .Z(n22709) );
  NANDN U23207 ( .A(n20875), .B(\stack[5][48] ), .Z(n22711) );
  NAND U23208 ( .A(n22712), .B(n22713), .Z(n4530) );
  NANDN U23209 ( .A(n21188), .B(\stack[6][49] ), .Z(n22713) );
  NANDN U23210 ( .A(n20866), .B(n22714), .Z(n22712) );
  NANDN U23211 ( .A(n22715), .B(n22716), .Z(n22714) );
  NANDN U23212 ( .A(n20875), .B(\stack[5][49] ), .Z(n22716) );
  NAND U23213 ( .A(n22717), .B(n22718), .Z(n4529) );
  NANDN U23214 ( .A(n21188), .B(\stack[6][50] ), .Z(n22718) );
  NANDN U23215 ( .A(n20866), .B(n22719), .Z(n22717) );
  NANDN U23216 ( .A(n22720), .B(n22721), .Z(n22719) );
  NANDN U23217 ( .A(n20875), .B(\stack[5][50] ), .Z(n22721) );
  NAND U23218 ( .A(n22722), .B(n22723), .Z(n4528) );
  NANDN U23219 ( .A(n21188), .B(\stack[6][51] ), .Z(n22723) );
  NANDN U23220 ( .A(n20866), .B(n22724), .Z(n22722) );
  NANDN U23221 ( .A(n22725), .B(n22726), .Z(n22724) );
  NANDN U23222 ( .A(n20875), .B(\stack[5][51] ), .Z(n22726) );
  NAND U23223 ( .A(n22727), .B(n22728), .Z(n4527) );
  NANDN U23224 ( .A(n21188), .B(\stack[6][52] ), .Z(n22728) );
  NANDN U23225 ( .A(n20866), .B(n22729), .Z(n22727) );
  NANDN U23226 ( .A(n22730), .B(n22731), .Z(n22729) );
  NANDN U23227 ( .A(n20875), .B(\stack[5][52] ), .Z(n22731) );
  NAND U23228 ( .A(n22732), .B(n22733), .Z(n4526) );
  NANDN U23229 ( .A(n21188), .B(\stack[6][53] ), .Z(n22733) );
  NANDN U23230 ( .A(n20866), .B(n22734), .Z(n22732) );
  NANDN U23231 ( .A(n22735), .B(n22736), .Z(n22734) );
  NANDN U23232 ( .A(n20875), .B(\stack[5][53] ), .Z(n22736) );
  NAND U23233 ( .A(n22737), .B(n22738), .Z(n4525) );
  NANDN U23234 ( .A(n21188), .B(\stack[6][54] ), .Z(n22738) );
  NANDN U23235 ( .A(n20866), .B(n22739), .Z(n22737) );
  NANDN U23236 ( .A(n22740), .B(n22741), .Z(n22739) );
  NANDN U23237 ( .A(n20875), .B(\stack[5][54] ), .Z(n22741) );
  NAND U23238 ( .A(n22742), .B(n22743), .Z(n4524) );
  NANDN U23239 ( .A(n21188), .B(\stack[6][55] ), .Z(n22743) );
  NANDN U23240 ( .A(n20866), .B(n22744), .Z(n22742) );
  NANDN U23241 ( .A(n22745), .B(n22746), .Z(n22744) );
  NANDN U23242 ( .A(n20875), .B(\stack[5][55] ), .Z(n22746) );
  NAND U23243 ( .A(n22747), .B(n22748), .Z(n4523) );
  NANDN U23244 ( .A(n21188), .B(\stack[6][56] ), .Z(n22748) );
  NANDN U23245 ( .A(n20866), .B(n22749), .Z(n22747) );
  NANDN U23246 ( .A(n22750), .B(n22751), .Z(n22749) );
  NANDN U23247 ( .A(n20875), .B(\stack[5][56] ), .Z(n22751) );
  NAND U23248 ( .A(n22752), .B(n22753), .Z(n4522) );
  NANDN U23249 ( .A(n21188), .B(\stack[6][57] ), .Z(n22753) );
  NANDN U23250 ( .A(n20866), .B(n22754), .Z(n22752) );
  NANDN U23251 ( .A(n22755), .B(n22756), .Z(n22754) );
  NANDN U23252 ( .A(n20875), .B(\stack[5][57] ), .Z(n22756) );
  NAND U23253 ( .A(n22757), .B(n22758), .Z(n4521) );
  NANDN U23254 ( .A(n21188), .B(\stack[6][58] ), .Z(n22758) );
  NANDN U23255 ( .A(n20866), .B(n22759), .Z(n22757) );
  NANDN U23256 ( .A(n22760), .B(n22761), .Z(n22759) );
  NANDN U23257 ( .A(n20875), .B(\stack[5][58] ), .Z(n22761) );
  NAND U23258 ( .A(n22762), .B(n22763), .Z(n4520) );
  NANDN U23259 ( .A(n21188), .B(\stack[6][59] ), .Z(n22763) );
  NANDN U23260 ( .A(n20866), .B(n22764), .Z(n22762) );
  NANDN U23261 ( .A(n22765), .B(n22766), .Z(n22764) );
  NANDN U23262 ( .A(n20875), .B(\stack[5][59] ), .Z(n22766) );
  NAND U23263 ( .A(n22767), .B(n22768), .Z(n4519) );
  NANDN U23264 ( .A(n21188), .B(\stack[6][60] ), .Z(n22768) );
  NANDN U23265 ( .A(n20866), .B(n22769), .Z(n22767) );
  NANDN U23266 ( .A(n22770), .B(n22771), .Z(n22769) );
  NANDN U23267 ( .A(n20875), .B(\stack[5][60] ), .Z(n22771) );
  NAND U23268 ( .A(n22772), .B(n22773), .Z(n4518) );
  NANDN U23269 ( .A(n21188), .B(\stack[6][61] ), .Z(n22773) );
  NANDN U23270 ( .A(n20866), .B(n22774), .Z(n22772) );
  NANDN U23271 ( .A(n22775), .B(n22776), .Z(n22774) );
  NANDN U23272 ( .A(n20875), .B(\stack[5][61] ), .Z(n22776) );
  NAND U23273 ( .A(n22777), .B(n22778), .Z(n4517) );
  NANDN U23274 ( .A(n21188), .B(\stack[6][62] ), .Z(n22778) );
  NANDN U23275 ( .A(n20866), .B(n22779), .Z(n22777) );
  NANDN U23276 ( .A(n22780), .B(n22781), .Z(n22779) );
  NANDN U23277 ( .A(n20875), .B(\stack[5][62] ), .Z(n22781) );
  NAND U23278 ( .A(n22782), .B(n22783), .Z(n4516) );
  NANDN U23279 ( .A(n21188), .B(\stack[6][63] ), .Z(n22783) );
  IV U23280 ( .A(n20866), .Z(n21188) );
  NANDN U23281 ( .A(n20866), .B(n22784), .Z(n22782) );
  NANDN U23282 ( .A(n22785), .B(n22786), .Z(n22784) );
  NANDN U23283 ( .A(n20875), .B(\stack[5][63] ), .Z(n22786) );
  NOR U23284 ( .A(n4967), .B(n6671), .Z(n20866) );
  NAND U23285 ( .A(n22787), .B(n22788), .Z(n6671) );
  NOR U23286 ( .A(n5168), .B(n20167), .Z(n22788) );
  ANDN U23287 ( .B(n20152), .A(n22789), .Z(n20167) );
  NOR U23288 ( .A(n20152), .B(n22789), .Z(n5168) );
  NANDN U23289 ( .A(opcode[2]), .B(opcode[1]), .Z(n22789) );
  ANDN U23290 ( .B(n20153), .A(n20166), .Z(n22787) );
  AND U23291 ( .A(n22790), .B(opcode[0]), .Z(n20166) );
  ANDN U23292 ( .B(n20156), .A(opcode[2]), .Z(n22790) );
  IV U23293 ( .A(opcode[1]), .Z(n20156) );
  NANDN U23294 ( .A(n20863), .B(opcode[1]), .Z(n20153) );
  IV U23295 ( .A(opcode[2]), .Z(n20863) );
  NANDN U23296 ( .A(n22475), .B(n22791), .Z(n4504) );
  NANDN U23297 ( .A(n20875), .B(\stack[6][1] ), .Z(n22791) );
  AND U23298 ( .A(\stack[7][1] ), .B(n20875), .Z(n22475) );
  NANDN U23299 ( .A(n22480), .B(n22792), .Z(n4495) );
  NANDN U23300 ( .A(n20875), .B(\stack[6][2] ), .Z(n22792) );
  AND U23301 ( .A(\stack[7][2] ), .B(n20875), .Z(n22480) );
  NANDN U23302 ( .A(n22485), .B(n22793), .Z(n4486) );
  NANDN U23303 ( .A(n20875), .B(\stack[6][3] ), .Z(n22793) );
  AND U23304 ( .A(\stack[7][3] ), .B(n20875), .Z(n22485) );
  NANDN U23305 ( .A(n22490), .B(n22794), .Z(n4477) );
  NANDN U23306 ( .A(n20875), .B(\stack[6][4] ), .Z(n22794) );
  AND U23307 ( .A(\stack[7][4] ), .B(n20875), .Z(n22490) );
  NANDN U23308 ( .A(n22495), .B(n22795), .Z(n4468) );
  NANDN U23309 ( .A(n20875), .B(\stack[6][5] ), .Z(n22795) );
  AND U23310 ( .A(\stack[7][5] ), .B(n20875), .Z(n22495) );
  NANDN U23311 ( .A(n22500), .B(n22796), .Z(n4459) );
  NANDN U23312 ( .A(n20875), .B(\stack[6][6] ), .Z(n22796) );
  AND U23313 ( .A(\stack[7][6] ), .B(n20875), .Z(n22500) );
  NANDN U23314 ( .A(n22505), .B(n22797), .Z(n4450) );
  NANDN U23315 ( .A(n20875), .B(\stack[6][7] ), .Z(n22797) );
  AND U23316 ( .A(\stack[7][7] ), .B(n20875), .Z(n22505) );
  NANDN U23317 ( .A(n22510), .B(n22798), .Z(n4441) );
  NANDN U23318 ( .A(n20875), .B(\stack[6][8] ), .Z(n22798) );
  AND U23319 ( .A(\stack[7][8] ), .B(n20875), .Z(n22510) );
  NANDN U23320 ( .A(n22515), .B(n22799), .Z(n4432) );
  NANDN U23321 ( .A(n20875), .B(\stack[6][9] ), .Z(n22799) );
  AND U23322 ( .A(\stack[7][9] ), .B(n20875), .Z(n22515) );
  NANDN U23323 ( .A(n22520), .B(n22800), .Z(n4423) );
  NANDN U23324 ( .A(n20875), .B(\stack[6][10] ), .Z(n22800) );
  AND U23325 ( .A(\stack[7][10] ), .B(n20875), .Z(n22520) );
  NANDN U23326 ( .A(n22525), .B(n22801), .Z(n4414) );
  NANDN U23327 ( .A(n20875), .B(\stack[6][11] ), .Z(n22801) );
  AND U23328 ( .A(\stack[7][11] ), .B(n20875), .Z(n22525) );
  NANDN U23329 ( .A(n22530), .B(n22802), .Z(n4405) );
  NANDN U23330 ( .A(n20875), .B(\stack[6][12] ), .Z(n22802) );
  AND U23331 ( .A(\stack[7][12] ), .B(n20875), .Z(n22530) );
  NANDN U23332 ( .A(n22535), .B(n22803), .Z(n4396) );
  NANDN U23333 ( .A(n20875), .B(\stack[6][13] ), .Z(n22803) );
  AND U23334 ( .A(\stack[7][13] ), .B(n20875), .Z(n22535) );
  NANDN U23335 ( .A(n22540), .B(n22804), .Z(n4387) );
  NANDN U23336 ( .A(n20875), .B(\stack[6][14] ), .Z(n22804) );
  AND U23337 ( .A(\stack[7][14] ), .B(n20875), .Z(n22540) );
  NANDN U23338 ( .A(n22545), .B(n22805), .Z(n4378) );
  NANDN U23339 ( .A(n20875), .B(\stack[6][15] ), .Z(n22805) );
  AND U23340 ( .A(\stack[7][15] ), .B(n20875), .Z(n22545) );
  NANDN U23341 ( .A(n22550), .B(n22806), .Z(n4369) );
  NANDN U23342 ( .A(n20875), .B(\stack[6][16] ), .Z(n22806) );
  AND U23343 ( .A(\stack[7][16] ), .B(n20875), .Z(n22550) );
  NANDN U23344 ( .A(n22555), .B(n22807), .Z(n4360) );
  NANDN U23345 ( .A(n20875), .B(\stack[6][17] ), .Z(n22807) );
  AND U23346 ( .A(\stack[7][17] ), .B(n20875), .Z(n22555) );
  NANDN U23347 ( .A(n22560), .B(n22808), .Z(n4351) );
  NANDN U23348 ( .A(n20875), .B(\stack[6][18] ), .Z(n22808) );
  AND U23349 ( .A(\stack[7][18] ), .B(n20875), .Z(n22560) );
  NANDN U23350 ( .A(n22565), .B(n22809), .Z(n4342) );
  NANDN U23351 ( .A(n20875), .B(\stack[6][19] ), .Z(n22809) );
  AND U23352 ( .A(\stack[7][19] ), .B(n20875), .Z(n22565) );
  NANDN U23353 ( .A(n22570), .B(n22810), .Z(n4333) );
  NANDN U23354 ( .A(n20875), .B(\stack[6][20] ), .Z(n22810) );
  AND U23355 ( .A(\stack[7][20] ), .B(n20875), .Z(n22570) );
  NANDN U23356 ( .A(n22575), .B(n22811), .Z(n4324) );
  NANDN U23357 ( .A(n20875), .B(\stack[6][21] ), .Z(n22811) );
  AND U23358 ( .A(\stack[7][21] ), .B(n20875), .Z(n22575) );
  NANDN U23359 ( .A(n22580), .B(n22812), .Z(n4315) );
  NANDN U23360 ( .A(n20875), .B(\stack[6][22] ), .Z(n22812) );
  AND U23361 ( .A(\stack[7][22] ), .B(n20875), .Z(n22580) );
  NANDN U23362 ( .A(n22585), .B(n22813), .Z(n4306) );
  NANDN U23363 ( .A(n20875), .B(\stack[6][23] ), .Z(n22813) );
  AND U23364 ( .A(\stack[7][23] ), .B(n20875), .Z(n22585) );
  NANDN U23365 ( .A(n22590), .B(n22814), .Z(n4297) );
  NANDN U23366 ( .A(n20875), .B(\stack[6][24] ), .Z(n22814) );
  AND U23367 ( .A(\stack[7][24] ), .B(n20875), .Z(n22590) );
  NANDN U23368 ( .A(n22595), .B(n22815), .Z(n4288) );
  NANDN U23369 ( .A(n20875), .B(\stack[6][25] ), .Z(n22815) );
  AND U23370 ( .A(\stack[7][25] ), .B(n20875), .Z(n22595) );
  NANDN U23371 ( .A(n22600), .B(n22816), .Z(n4279) );
  NANDN U23372 ( .A(n20875), .B(\stack[6][26] ), .Z(n22816) );
  AND U23373 ( .A(\stack[7][26] ), .B(n20875), .Z(n22600) );
  NANDN U23374 ( .A(n22605), .B(n22817), .Z(n4270) );
  NANDN U23375 ( .A(n20875), .B(\stack[6][27] ), .Z(n22817) );
  AND U23376 ( .A(\stack[7][27] ), .B(n20875), .Z(n22605) );
  NANDN U23377 ( .A(n22610), .B(n22818), .Z(n4261) );
  NANDN U23378 ( .A(n20875), .B(\stack[6][28] ), .Z(n22818) );
  AND U23379 ( .A(\stack[7][28] ), .B(n20875), .Z(n22610) );
  NANDN U23380 ( .A(n22615), .B(n22819), .Z(n4252) );
  NANDN U23381 ( .A(n20875), .B(\stack[6][29] ), .Z(n22819) );
  AND U23382 ( .A(\stack[7][29] ), .B(n20875), .Z(n22615) );
  NANDN U23383 ( .A(n22620), .B(n22820), .Z(n4243) );
  NANDN U23384 ( .A(n20875), .B(\stack[6][30] ), .Z(n22820) );
  AND U23385 ( .A(\stack[7][30] ), .B(n20875), .Z(n22620) );
  NANDN U23386 ( .A(n22625), .B(n22821), .Z(n4234) );
  NANDN U23387 ( .A(n20875), .B(\stack[6][31] ), .Z(n22821) );
  AND U23388 ( .A(\stack[7][31] ), .B(n20875), .Z(n22625) );
  NANDN U23389 ( .A(n22630), .B(n22822), .Z(n4225) );
  NANDN U23390 ( .A(n20875), .B(\stack[6][32] ), .Z(n22822) );
  AND U23391 ( .A(\stack[7][32] ), .B(n20875), .Z(n22630) );
  NANDN U23392 ( .A(n22635), .B(n22823), .Z(n4216) );
  NANDN U23393 ( .A(n20875), .B(\stack[6][33] ), .Z(n22823) );
  AND U23394 ( .A(\stack[7][33] ), .B(n20875), .Z(n22635) );
  NANDN U23395 ( .A(n22640), .B(n22824), .Z(n4207) );
  NANDN U23396 ( .A(n20875), .B(\stack[6][34] ), .Z(n22824) );
  AND U23397 ( .A(\stack[7][34] ), .B(n20875), .Z(n22640) );
  NANDN U23398 ( .A(n22645), .B(n22825), .Z(n4198) );
  NANDN U23399 ( .A(n20875), .B(\stack[6][35] ), .Z(n22825) );
  AND U23400 ( .A(\stack[7][35] ), .B(n20875), .Z(n22645) );
  NANDN U23401 ( .A(n22650), .B(n22826), .Z(n4189) );
  NANDN U23402 ( .A(n20875), .B(\stack[6][36] ), .Z(n22826) );
  AND U23403 ( .A(\stack[7][36] ), .B(n20875), .Z(n22650) );
  NANDN U23404 ( .A(n22655), .B(n22827), .Z(n4180) );
  NANDN U23405 ( .A(n20875), .B(\stack[6][37] ), .Z(n22827) );
  AND U23406 ( .A(\stack[7][37] ), .B(n20875), .Z(n22655) );
  NANDN U23407 ( .A(n22660), .B(n22828), .Z(n4171) );
  NANDN U23408 ( .A(n20875), .B(\stack[6][38] ), .Z(n22828) );
  AND U23409 ( .A(\stack[7][38] ), .B(n20875), .Z(n22660) );
  NANDN U23410 ( .A(n22665), .B(n22829), .Z(n4162) );
  NANDN U23411 ( .A(n20875), .B(\stack[6][39] ), .Z(n22829) );
  AND U23412 ( .A(\stack[7][39] ), .B(n20875), .Z(n22665) );
  NANDN U23413 ( .A(n22670), .B(n22830), .Z(n4153) );
  NANDN U23414 ( .A(n20875), .B(\stack[6][40] ), .Z(n22830) );
  AND U23415 ( .A(\stack[7][40] ), .B(n20875), .Z(n22670) );
  NANDN U23416 ( .A(n22675), .B(n22831), .Z(n4144) );
  NANDN U23417 ( .A(n20875), .B(\stack[6][41] ), .Z(n22831) );
  AND U23418 ( .A(\stack[7][41] ), .B(n20875), .Z(n22675) );
  NANDN U23419 ( .A(n22680), .B(n22832), .Z(n4135) );
  NANDN U23420 ( .A(n20875), .B(\stack[6][42] ), .Z(n22832) );
  AND U23421 ( .A(\stack[7][42] ), .B(n20875), .Z(n22680) );
  NANDN U23422 ( .A(n22685), .B(n22833), .Z(n4126) );
  NANDN U23423 ( .A(n20875), .B(\stack[6][43] ), .Z(n22833) );
  AND U23424 ( .A(\stack[7][43] ), .B(n20875), .Z(n22685) );
  NANDN U23425 ( .A(n22690), .B(n22834), .Z(n4117) );
  NANDN U23426 ( .A(n20875), .B(\stack[6][44] ), .Z(n22834) );
  AND U23427 ( .A(\stack[7][44] ), .B(n20875), .Z(n22690) );
  NANDN U23428 ( .A(n22695), .B(n22835), .Z(n4108) );
  NANDN U23429 ( .A(n20875), .B(\stack[6][45] ), .Z(n22835) );
  AND U23430 ( .A(\stack[7][45] ), .B(n20875), .Z(n22695) );
  NANDN U23431 ( .A(n22700), .B(n22836), .Z(n4099) );
  NANDN U23432 ( .A(n20875), .B(\stack[6][46] ), .Z(n22836) );
  AND U23433 ( .A(\stack[7][46] ), .B(n20875), .Z(n22700) );
  NANDN U23434 ( .A(n22705), .B(n22837), .Z(n4090) );
  NANDN U23435 ( .A(n20875), .B(\stack[6][47] ), .Z(n22837) );
  AND U23436 ( .A(\stack[7][47] ), .B(n20875), .Z(n22705) );
  NANDN U23437 ( .A(n22710), .B(n22838), .Z(n4081) );
  NANDN U23438 ( .A(n20875), .B(\stack[6][48] ), .Z(n22838) );
  AND U23439 ( .A(\stack[7][48] ), .B(n20875), .Z(n22710) );
  NANDN U23440 ( .A(n22715), .B(n22839), .Z(n4072) );
  NANDN U23441 ( .A(n20875), .B(\stack[6][49] ), .Z(n22839) );
  AND U23442 ( .A(\stack[7][49] ), .B(n20875), .Z(n22715) );
  NANDN U23443 ( .A(n22720), .B(n22840), .Z(n4063) );
  NANDN U23444 ( .A(n20875), .B(\stack[6][50] ), .Z(n22840) );
  AND U23445 ( .A(\stack[7][50] ), .B(n20875), .Z(n22720) );
  NANDN U23446 ( .A(n22725), .B(n22841), .Z(n4054) );
  NANDN U23447 ( .A(n20875), .B(\stack[6][51] ), .Z(n22841) );
  AND U23448 ( .A(\stack[7][51] ), .B(n20875), .Z(n22725) );
  NANDN U23449 ( .A(n22730), .B(n22842), .Z(n4045) );
  NANDN U23450 ( .A(n20875), .B(\stack[6][52] ), .Z(n22842) );
  AND U23451 ( .A(\stack[7][52] ), .B(n20875), .Z(n22730) );
  NANDN U23452 ( .A(n22735), .B(n22843), .Z(n4036) );
  NANDN U23453 ( .A(n20875), .B(\stack[6][53] ), .Z(n22843) );
  AND U23454 ( .A(\stack[7][53] ), .B(n20875), .Z(n22735) );
  NANDN U23455 ( .A(n22740), .B(n22844), .Z(n4027) );
  NANDN U23456 ( .A(n20875), .B(\stack[6][54] ), .Z(n22844) );
  AND U23457 ( .A(\stack[7][54] ), .B(n20875), .Z(n22740) );
  NANDN U23458 ( .A(n22745), .B(n22845), .Z(n4018) );
  NANDN U23459 ( .A(n20875), .B(\stack[6][55] ), .Z(n22845) );
  AND U23460 ( .A(\stack[7][55] ), .B(n20875), .Z(n22745) );
  NANDN U23461 ( .A(n22750), .B(n22846), .Z(n4009) );
  NANDN U23462 ( .A(n20875), .B(\stack[6][56] ), .Z(n22846) );
  AND U23463 ( .A(\stack[7][56] ), .B(n20875), .Z(n22750) );
  NANDN U23464 ( .A(n22755), .B(n22847), .Z(n4000) );
  NANDN U23465 ( .A(n20875), .B(\stack[6][57] ), .Z(n22847) );
  AND U23466 ( .A(\stack[7][57] ), .B(n20875), .Z(n22755) );
  NANDN U23467 ( .A(n22760), .B(n22848), .Z(n3991) );
  NANDN U23468 ( .A(n20875), .B(\stack[6][58] ), .Z(n22848) );
  AND U23469 ( .A(\stack[7][58] ), .B(n20875), .Z(n22760) );
  NANDN U23470 ( .A(n22765), .B(n22849), .Z(n3982) );
  NANDN U23471 ( .A(n20875), .B(\stack[6][59] ), .Z(n22849) );
  AND U23472 ( .A(\stack[7][59] ), .B(n20875), .Z(n22765) );
  NANDN U23473 ( .A(n22770), .B(n22850), .Z(n3973) );
  NANDN U23474 ( .A(n20875), .B(\stack[6][60] ), .Z(n22850) );
  AND U23475 ( .A(\stack[7][60] ), .B(n20875), .Z(n22770) );
  NANDN U23476 ( .A(n22775), .B(n22851), .Z(n3964) );
  NANDN U23477 ( .A(n20875), .B(\stack[6][61] ), .Z(n22851) );
  AND U23478 ( .A(\stack[7][61] ), .B(n20875), .Z(n22775) );
  NANDN U23479 ( .A(n22780), .B(n22852), .Z(n3955) );
  NANDN U23480 ( .A(n20875), .B(\stack[6][62] ), .Z(n22852) );
  AND U23481 ( .A(\stack[7][62] ), .B(n20875), .Z(n22780) );
  NANDN U23482 ( .A(n22785), .B(n22853), .Z(n3948) );
  NANDN U23483 ( .A(n20875), .B(\stack[6][63] ), .Z(n22853) );
  AND U23484 ( .A(\stack[7][63] ), .B(n20875), .Z(n22785) );
  NANDN U23485 ( .A(n22470), .B(n22854), .Z(n3941) );
  NANDN U23486 ( .A(n20875), .B(\stack[6][0] ), .Z(n22854) );
  AND U23487 ( .A(\stack[7][0] ), .B(n20875), .Z(n22470) );
  IV U23488 ( .A(n4967), .Z(n20875) );
  AND U23489 ( .A(n22855), .B(opcode[2]), .Z(n4967) );
  ANDN U23490 ( .B(n20152), .A(opcode[1]), .Z(n22855) );
  IV U23491 ( .A(opcode[0]), .Z(n20152) );
endmodule

