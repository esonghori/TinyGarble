
module sum_N1024_CC32 ( clk, rst, a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n5) );
  NAND U6 ( .A(a[0]), .B(b[0]), .Z(n3) );
  NAND U7 ( .A(n1), .B(carry_on), .Z(n2) );
  NAND U8 ( .A(n3), .B(n2), .Z(n4) );
  XOR U9 ( .A(n5), .B(n4), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n9) );
  NAND U11 ( .A(a[1]), .B(b[1]), .Z(n7) );
  NAND U12 ( .A(n5), .B(n4), .Z(n6) );
  NAND U13 ( .A(n7), .B(n6), .Z(n8) );
  XOR U14 ( .A(n9), .B(n8), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n13) );
  NAND U16 ( .A(a[2]), .B(b[2]), .Z(n11) );
  NAND U17 ( .A(n9), .B(n8), .Z(n10) );
  NAND U18 ( .A(n11), .B(n10), .Z(n12) );
  XOR U19 ( .A(n13), .B(n12), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n17) );
  NAND U21 ( .A(a[3]), .B(b[3]), .Z(n15) );
  NAND U22 ( .A(n13), .B(n12), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n16) );
  XOR U24 ( .A(n17), .B(n16), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n21) );
  NAND U26 ( .A(a[4]), .B(b[4]), .Z(n19) );
  NAND U27 ( .A(n17), .B(n16), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n20) );
  XOR U29 ( .A(n21), .B(n20), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n25) );
  NAND U31 ( .A(a[5]), .B(b[5]), .Z(n23) );
  NAND U32 ( .A(n21), .B(n20), .Z(n22) );
  NAND U33 ( .A(n23), .B(n22), .Z(n24) );
  XOR U34 ( .A(n25), .B(n24), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n29) );
  NAND U36 ( .A(a[6]), .B(b[6]), .Z(n27) );
  NAND U37 ( .A(n25), .B(n24), .Z(n26) );
  NAND U38 ( .A(n27), .B(n26), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n33) );
  NAND U41 ( .A(a[7]), .B(b[7]), .Z(n31) );
  NAND U42 ( .A(n29), .B(n28), .Z(n30) );
  NAND U43 ( .A(n31), .B(n30), .Z(n32) );
  XOR U44 ( .A(n33), .B(n32), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n37) );
  NAND U46 ( .A(a[8]), .B(b[8]), .Z(n35) );
  NAND U47 ( .A(n33), .B(n32), .Z(n34) );
  NAND U48 ( .A(n35), .B(n34), .Z(n36) );
  XOR U49 ( .A(n37), .B(n36), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n41) );
  NAND U51 ( .A(a[9]), .B(b[9]), .Z(n39) );
  NAND U52 ( .A(n37), .B(n36), .Z(n38) );
  NAND U53 ( .A(n39), .B(n38), .Z(n40) );
  XOR U54 ( .A(n41), .B(n40), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n45) );
  NAND U56 ( .A(a[10]), .B(b[10]), .Z(n43) );
  NAND U57 ( .A(n41), .B(n40), .Z(n42) );
  NAND U58 ( .A(n43), .B(n42), .Z(n44) );
  XOR U59 ( .A(n45), .B(n44), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n49) );
  NAND U61 ( .A(a[11]), .B(b[11]), .Z(n47) );
  NAND U62 ( .A(n45), .B(n44), .Z(n46) );
  NAND U63 ( .A(n47), .B(n46), .Z(n48) );
  XOR U64 ( .A(n49), .B(n48), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n53) );
  NAND U66 ( .A(a[12]), .B(b[12]), .Z(n51) );
  NAND U67 ( .A(n49), .B(n48), .Z(n50) );
  NAND U68 ( .A(n51), .B(n50), .Z(n52) );
  XOR U69 ( .A(n53), .B(n52), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n57) );
  NAND U71 ( .A(a[13]), .B(b[13]), .Z(n55) );
  NAND U72 ( .A(n53), .B(n52), .Z(n54) );
  NAND U73 ( .A(n55), .B(n54), .Z(n56) );
  XOR U74 ( .A(n57), .B(n56), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n61) );
  NAND U76 ( .A(a[14]), .B(b[14]), .Z(n59) );
  NAND U77 ( .A(n57), .B(n56), .Z(n58) );
  NAND U78 ( .A(n59), .B(n58), .Z(n60) );
  XOR U79 ( .A(n61), .B(n60), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n65) );
  NAND U81 ( .A(a[15]), .B(b[15]), .Z(n63) );
  NAND U82 ( .A(n61), .B(n60), .Z(n62) );
  NAND U83 ( .A(n63), .B(n62), .Z(n64) );
  XOR U84 ( .A(n65), .B(n64), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n69) );
  NAND U86 ( .A(a[16]), .B(b[16]), .Z(n67) );
  NAND U87 ( .A(n65), .B(n64), .Z(n66) );
  NAND U88 ( .A(n67), .B(n66), .Z(n68) );
  XOR U89 ( .A(n69), .B(n68), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n73) );
  NAND U91 ( .A(a[17]), .B(b[17]), .Z(n71) );
  NAND U92 ( .A(n69), .B(n68), .Z(n70) );
  NAND U93 ( .A(n71), .B(n70), .Z(n72) );
  XOR U94 ( .A(n73), .B(n72), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n77) );
  NAND U96 ( .A(a[18]), .B(b[18]), .Z(n75) );
  NAND U97 ( .A(n73), .B(n72), .Z(n74) );
  NAND U98 ( .A(n75), .B(n74), .Z(n76) );
  XOR U99 ( .A(n77), .B(n76), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n81) );
  NAND U101 ( .A(a[19]), .B(b[19]), .Z(n79) );
  NAND U102 ( .A(n77), .B(n76), .Z(n78) );
  NAND U103 ( .A(n79), .B(n78), .Z(n80) );
  XOR U104 ( .A(n81), .B(n80), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n85) );
  NAND U106 ( .A(a[20]), .B(b[20]), .Z(n83) );
  NAND U107 ( .A(n81), .B(n80), .Z(n82) );
  NAND U108 ( .A(n83), .B(n82), .Z(n84) );
  XOR U109 ( .A(n85), .B(n84), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n89) );
  NAND U111 ( .A(a[21]), .B(b[21]), .Z(n87) );
  NAND U112 ( .A(n85), .B(n84), .Z(n86) );
  NAND U113 ( .A(n87), .B(n86), .Z(n88) );
  XOR U114 ( .A(n89), .B(n88), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n93) );
  NAND U116 ( .A(a[22]), .B(b[22]), .Z(n91) );
  NAND U117 ( .A(n89), .B(n88), .Z(n90) );
  NAND U118 ( .A(n91), .B(n90), .Z(n92) );
  XOR U119 ( .A(n93), .B(n92), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n97) );
  NAND U121 ( .A(a[23]), .B(b[23]), .Z(n95) );
  NAND U122 ( .A(n93), .B(n92), .Z(n94) );
  NAND U123 ( .A(n95), .B(n94), .Z(n96) );
  XOR U124 ( .A(n97), .B(n96), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n101) );
  NAND U126 ( .A(a[24]), .B(b[24]), .Z(n99) );
  NAND U127 ( .A(n97), .B(n96), .Z(n98) );
  NAND U128 ( .A(n99), .B(n98), .Z(n100) );
  XOR U129 ( .A(n101), .B(n100), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n105) );
  NAND U131 ( .A(a[25]), .B(b[25]), .Z(n103) );
  NAND U132 ( .A(n101), .B(n100), .Z(n102) );
  NAND U133 ( .A(n103), .B(n102), .Z(n104) );
  XOR U134 ( .A(n105), .B(n104), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n109) );
  NAND U136 ( .A(a[26]), .B(b[26]), .Z(n107) );
  NAND U137 ( .A(n105), .B(n104), .Z(n106) );
  NAND U138 ( .A(n107), .B(n106), .Z(n108) );
  XOR U139 ( .A(n109), .B(n108), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n113) );
  NAND U141 ( .A(a[27]), .B(b[27]), .Z(n111) );
  NAND U142 ( .A(n109), .B(n108), .Z(n110) );
  NAND U143 ( .A(n111), .B(n110), .Z(n112) );
  XOR U144 ( .A(n113), .B(n112), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n117) );
  NAND U146 ( .A(a[28]), .B(b[28]), .Z(n115) );
  NAND U147 ( .A(n113), .B(n112), .Z(n114) );
  NAND U148 ( .A(n115), .B(n114), .Z(n116) );
  XOR U149 ( .A(n117), .B(n116), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n121) );
  NAND U151 ( .A(a[29]), .B(b[29]), .Z(n119) );
  NAND U152 ( .A(n117), .B(n116), .Z(n118) );
  NAND U153 ( .A(n119), .B(n118), .Z(n120) );
  XOR U154 ( .A(n121), .B(n120), .Z(c[30]) );
  NAND U155 ( .A(a[30]), .B(b[30]), .Z(n123) );
  NAND U156 ( .A(n121), .B(n120), .Z(n122) );
  AND U157 ( .A(n123), .B(n122), .Z(n125) );
  XOR U158 ( .A(a[31]), .B(b[31]), .Z(n124) );
  XNOR U159 ( .A(n125), .B(n124), .Z(c[31]) );
  NAND U160 ( .A(a[31]), .B(b[31]), .Z(n127) );
  NANDN U161 ( .A(n125), .B(n124), .Z(n126) );
  NAND U162 ( .A(n127), .B(n126), .Z(carry_on_d) );
endmodule

