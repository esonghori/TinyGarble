
module mult_N32_CC1 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [63:0] o;
  input clk, rst;
  wire   \mult_26/A2[31] , \mult_26/A2[32] , \mult_26/A2[33] ,
         \mult_26/A2[34] , \mult_26/A2[35] , \mult_26/A2[36] ,
         \mult_26/A2[37] , \mult_26/A2[38] , \mult_26/A2[39] ,
         \mult_26/A2[40] , \mult_26/A2[41] , \mult_26/A2[42] ,
         \mult_26/A2[43] , \mult_26/A2[44] , \mult_26/A2[45] ,
         \mult_26/A2[46] , \mult_26/A2[47] , \mult_26/A2[48] ,
         \mult_26/A2[49] , \mult_26/A2[50] , \mult_26/A2[51] ,
         \mult_26/A2[52] , \mult_26/A2[53] , \mult_26/A2[54] ,
         \mult_26/A2[55] , \mult_26/A2[56] , \mult_26/A2[57] ,
         \mult_26/A2[58] , \mult_26/A2[59] , \mult_26/A2[60] ,
         \mult_26/A2[61] , \mult_26/A1[31] , \mult_26/A1[32] ,
         \mult_26/A1[33] , \mult_26/A1[34] , \mult_26/A1[35] ,
         \mult_26/A1[36] , \mult_26/A1[37] , \mult_26/A1[38] ,
         \mult_26/A1[39] , \mult_26/A1[40] , \mult_26/A1[41] ,
         \mult_26/A1[42] , \mult_26/A1[43] , \mult_26/A1[44] ,
         \mult_26/A1[45] , \mult_26/A1[46] , \mult_26/A1[47] ,
         \mult_26/A1[48] , \mult_26/A1[49] , \mult_26/A1[50] ,
         \mult_26/A1[51] , \mult_26/A1[52] , \mult_26/A1[53] ,
         \mult_26/A1[54] , \mult_26/A1[55] , \mult_26/A1[56] ,
         \mult_26/A1[57] , \mult_26/A1[58] , \mult_26/A1[59] ,
         \mult_26/A1[60] , \mult_26/SUMB[16][1] , \mult_26/SUMB[16][2] ,
         \mult_26/SUMB[16][3] , \mult_26/SUMB[16][4] , \mult_26/SUMB[16][5] ,
         \mult_26/SUMB[16][6] , \mult_26/SUMB[16][7] , \mult_26/SUMB[16][8] ,
         \mult_26/SUMB[16][9] , \mult_26/SUMB[16][10] , \mult_26/SUMB[16][11] ,
         \mult_26/SUMB[16][12] , \mult_26/SUMB[16][13] ,
         \mult_26/SUMB[16][14] , \mult_26/SUMB[16][15] ,
         \mult_26/SUMB[16][16] , \mult_26/SUMB[16][17] ,
         \mult_26/SUMB[16][18] , \mult_26/SUMB[16][19] ,
         \mult_26/SUMB[16][20] , \mult_26/SUMB[16][21] ,
         \mult_26/SUMB[16][22] , \mult_26/SUMB[16][23] ,
         \mult_26/SUMB[16][24] , \mult_26/SUMB[16][25] ,
         \mult_26/SUMB[16][26] , \mult_26/SUMB[16][27] ,
         \mult_26/SUMB[16][28] , \mult_26/SUMB[16][29] ,
         \mult_26/SUMB[16][30] , \mult_26/SUMB[17][1] , \mult_26/SUMB[17][2] ,
         \mult_26/SUMB[17][3] , \mult_26/SUMB[17][4] , \mult_26/SUMB[17][5] ,
         \mult_26/SUMB[17][6] , \mult_26/SUMB[17][7] , \mult_26/SUMB[17][8] ,
         \mult_26/SUMB[17][9] , \mult_26/SUMB[17][10] , \mult_26/SUMB[17][11] ,
         \mult_26/SUMB[17][12] , \mult_26/SUMB[17][13] ,
         \mult_26/SUMB[17][14] , \mult_26/SUMB[17][15] ,
         \mult_26/SUMB[17][16] , \mult_26/SUMB[17][17] ,
         \mult_26/SUMB[17][18] , \mult_26/SUMB[17][19] ,
         \mult_26/SUMB[17][20] , \mult_26/SUMB[17][21] ,
         \mult_26/SUMB[17][22] , \mult_26/SUMB[17][23] ,
         \mult_26/SUMB[17][24] , \mult_26/SUMB[17][25] ,
         \mult_26/SUMB[17][26] , \mult_26/SUMB[17][27] ,
         \mult_26/SUMB[17][28] , \mult_26/SUMB[17][29] ,
         \mult_26/SUMB[17][30] , \mult_26/SUMB[18][1] , \mult_26/SUMB[18][2] ,
         \mult_26/SUMB[18][3] , \mult_26/SUMB[18][4] , \mult_26/SUMB[18][5] ,
         \mult_26/SUMB[18][6] , \mult_26/SUMB[18][7] , \mult_26/SUMB[18][8] ,
         \mult_26/SUMB[18][9] , \mult_26/SUMB[18][10] , \mult_26/SUMB[18][11] ,
         \mult_26/SUMB[18][12] , \mult_26/SUMB[18][13] ,
         \mult_26/SUMB[18][14] , \mult_26/SUMB[18][15] ,
         \mult_26/SUMB[18][16] , \mult_26/SUMB[18][17] ,
         \mult_26/SUMB[18][18] , \mult_26/SUMB[18][19] ,
         \mult_26/SUMB[18][20] , \mult_26/SUMB[18][21] ,
         \mult_26/SUMB[18][22] , \mult_26/SUMB[18][23] ,
         \mult_26/SUMB[18][24] , \mult_26/SUMB[18][25] ,
         \mult_26/SUMB[18][26] , \mult_26/SUMB[18][27] ,
         \mult_26/SUMB[18][28] , \mult_26/SUMB[18][29] ,
         \mult_26/SUMB[18][30] , \mult_26/SUMB[19][1] , \mult_26/SUMB[19][2] ,
         \mult_26/SUMB[19][3] , \mult_26/SUMB[19][4] , \mult_26/SUMB[19][5] ,
         \mult_26/SUMB[19][6] , \mult_26/SUMB[19][7] , \mult_26/SUMB[19][8] ,
         \mult_26/SUMB[19][9] , \mult_26/SUMB[19][10] , \mult_26/SUMB[19][11] ,
         \mult_26/SUMB[19][12] , \mult_26/SUMB[19][13] ,
         \mult_26/SUMB[19][14] , \mult_26/SUMB[19][15] ,
         \mult_26/SUMB[19][16] , \mult_26/SUMB[19][17] ,
         \mult_26/SUMB[19][18] , \mult_26/SUMB[19][19] ,
         \mult_26/SUMB[19][20] , \mult_26/SUMB[19][21] ,
         \mult_26/SUMB[19][22] , \mult_26/SUMB[19][23] ,
         \mult_26/SUMB[19][24] , \mult_26/SUMB[19][25] ,
         \mult_26/SUMB[19][26] , \mult_26/SUMB[19][27] ,
         \mult_26/SUMB[19][28] , \mult_26/SUMB[19][29] ,
         \mult_26/SUMB[19][30] , \mult_26/SUMB[20][1] , \mult_26/SUMB[20][2] ,
         \mult_26/SUMB[20][3] , \mult_26/SUMB[20][4] , \mult_26/SUMB[20][5] ,
         \mult_26/SUMB[20][6] , \mult_26/SUMB[20][7] , \mult_26/SUMB[20][8] ,
         \mult_26/SUMB[20][9] , \mult_26/SUMB[20][10] , \mult_26/SUMB[20][11] ,
         \mult_26/SUMB[20][12] , \mult_26/SUMB[20][13] ,
         \mult_26/SUMB[20][14] , \mult_26/SUMB[20][15] ,
         \mult_26/SUMB[20][16] , \mult_26/SUMB[20][17] ,
         \mult_26/SUMB[20][18] , \mult_26/SUMB[20][19] ,
         \mult_26/SUMB[20][20] , \mult_26/SUMB[20][21] ,
         \mult_26/SUMB[20][22] , \mult_26/SUMB[20][23] ,
         \mult_26/SUMB[20][24] , \mult_26/SUMB[20][25] ,
         \mult_26/SUMB[20][26] , \mult_26/SUMB[20][27] ,
         \mult_26/SUMB[20][28] , \mult_26/SUMB[20][29] ,
         \mult_26/SUMB[20][30] , \mult_26/SUMB[21][1] , \mult_26/SUMB[21][2] ,
         \mult_26/SUMB[21][3] , \mult_26/SUMB[21][4] , \mult_26/SUMB[21][5] ,
         \mult_26/SUMB[21][6] , \mult_26/SUMB[21][7] , \mult_26/SUMB[21][8] ,
         \mult_26/SUMB[21][9] , \mult_26/SUMB[21][10] , \mult_26/SUMB[21][11] ,
         \mult_26/SUMB[21][12] , \mult_26/SUMB[21][13] ,
         \mult_26/SUMB[21][14] , \mult_26/SUMB[21][15] ,
         \mult_26/SUMB[21][16] , \mult_26/SUMB[21][17] ,
         \mult_26/SUMB[21][18] , \mult_26/SUMB[21][19] ,
         \mult_26/SUMB[21][20] , \mult_26/SUMB[21][21] ,
         \mult_26/SUMB[21][22] , \mult_26/SUMB[21][23] ,
         \mult_26/SUMB[21][24] , \mult_26/SUMB[21][25] ,
         \mult_26/SUMB[21][26] , \mult_26/SUMB[21][27] ,
         \mult_26/SUMB[21][28] , \mult_26/SUMB[21][29] ,
         \mult_26/SUMB[21][30] , \mult_26/SUMB[22][1] , \mult_26/SUMB[22][2] ,
         \mult_26/SUMB[22][3] , \mult_26/SUMB[22][4] , \mult_26/SUMB[22][5] ,
         \mult_26/SUMB[22][6] , \mult_26/SUMB[22][7] , \mult_26/SUMB[22][8] ,
         \mult_26/SUMB[22][9] , \mult_26/SUMB[22][10] , \mult_26/SUMB[22][11] ,
         \mult_26/SUMB[22][12] , \mult_26/SUMB[22][13] ,
         \mult_26/SUMB[22][14] , \mult_26/SUMB[22][15] ,
         \mult_26/SUMB[22][16] , \mult_26/SUMB[22][17] ,
         \mult_26/SUMB[22][18] , \mult_26/SUMB[22][19] ,
         \mult_26/SUMB[22][20] , \mult_26/SUMB[22][21] ,
         \mult_26/SUMB[22][22] , \mult_26/SUMB[22][23] ,
         \mult_26/SUMB[22][24] , \mult_26/SUMB[22][25] ,
         \mult_26/SUMB[22][26] , \mult_26/SUMB[22][27] ,
         \mult_26/SUMB[22][28] , \mult_26/SUMB[22][29] ,
         \mult_26/SUMB[22][30] , \mult_26/SUMB[23][1] , \mult_26/SUMB[23][2] ,
         \mult_26/SUMB[23][3] , \mult_26/SUMB[23][4] , \mult_26/SUMB[23][5] ,
         \mult_26/SUMB[23][6] , \mult_26/SUMB[23][7] , \mult_26/SUMB[23][8] ,
         \mult_26/SUMB[23][9] , \mult_26/SUMB[23][10] , \mult_26/SUMB[23][11] ,
         \mult_26/SUMB[23][12] , \mult_26/SUMB[23][13] ,
         \mult_26/SUMB[23][14] , \mult_26/SUMB[23][15] ,
         \mult_26/SUMB[23][16] , \mult_26/SUMB[23][17] ,
         \mult_26/SUMB[23][18] , \mult_26/SUMB[23][19] ,
         \mult_26/SUMB[23][20] , \mult_26/SUMB[23][21] ,
         \mult_26/SUMB[23][22] , \mult_26/SUMB[23][23] ,
         \mult_26/SUMB[23][24] , \mult_26/SUMB[23][25] ,
         \mult_26/SUMB[23][26] , \mult_26/SUMB[23][27] ,
         \mult_26/SUMB[23][28] , \mult_26/SUMB[23][29] ,
         \mult_26/SUMB[23][30] , \mult_26/SUMB[24][1] , \mult_26/SUMB[24][2] ,
         \mult_26/SUMB[24][3] , \mult_26/SUMB[24][4] , \mult_26/SUMB[24][5] ,
         \mult_26/SUMB[24][6] , \mult_26/SUMB[24][7] , \mult_26/SUMB[24][8] ,
         \mult_26/SUMB[24][9] , \mult_26/SUMB[24][10] , \mult_26/SUMB[24][11] ,
         \mult_26/SUMB[24][12] , \mult_26/SUMB[24][13] ,
         \mult_26/SUMB[24][14] , \mult_26/SUMB[24][15] ,
         \mult_26/SUMB[24][16] , \mult_26/SUMB[24][17] ,
         \mult_26/SUMB[24][18] , \mult_26/SUMB[24][19] ,
         \mult_26/SUMB[24][20] , \mult_26/SUMB[24][21] ,
         \mult_26/SUMB[24][22] , \mult_26/SUMB[24][23] ,
         \mult_26/SUMB[24][24] , \mult_26/SUMB[24][25] ,
         \mult_26/SUMB[24][26] , \mult_26/SUMB[24][27] ,
         \mult_26/SUMB[24][28] , \mult_26/SUMB[24][29] ,
         \mult_26/SUMB[24][30] , \mult_26/SUMB[25][1] , \mult_26/SUMB[25][2] ,
         \mult_26/SUMB[25][3] , \mult_26/SUMB[25][4] , \mult_26/SUMB[25][5] ,
         \mult_26/SUMB[25][6] , \mult_26/SUMB[25][7] , \mult_26/SUMB[25][8] ,
         \mult_26/SUMB[25][9] , \mult_26/SUMB[25][10] , \mult_26/SUMB[25][11] ,
         \mult_26/SUMB[25][12] , \mult_26/SUMB[25][13] ,
         \mult_26/SUMB[25][14] , \mult_26/SUMB[25][15] ,
         \mult_26/SUMB[25][16] , \mult_26/SUMB[25][17] ,
         \mult_26/SUMB[25][18] , \mult_26/SUMB[25][19] ,
         \mult_26/SUMB[25][20] , \mult_26/SUMB[25][21] ,
         \mult_26/SUMB[25][22] , \mult_26/SUMB[25][23] ,
         \mult_26/SUMB[25][24] , \mult_26/SUMB[25][25] ,
         \mult_26/SUMB[25][26] , \mult_26/SUMB[25][27] ,
         \mult_26/SUMB[25][28] , \mult_26/SUMB[25][29] ,
         \mult_26/SUMB[25][30] , \mult_26/SUMB[26][1] , \mult_26/SUMB[26][2] ,
         \mult_26/SUMB[26][3] , \mult_26/SUMB[26][4] , \mult_26/SUMB[26][5] ,
         \mult_26/SUMB[26][6] , \mult_26/SUMB[26][7] , \mult_26/SUMB[26][8] ,
         \mult_26/SUMB[26][9] , \mult_26/SUMB[26][10] , \mult_26/SUMB[26][11] ,
         \mult_26/SUMB[26][12] , \mult_26/SUMB[26][13] ,
         \mult_26/SUMB[26][14] , \mult_26/SUMB[26][15] ,
         \mult_26/SUMB[26][16] , \mult_26/SUMB[26][17] ,
         \mult_26/SUMB[26][18] , \mult_26/SUMB[26][19] ,
         \mult_26/SUMB[26][20] , \mult_26/SUMB[26][21] ,
         \mult_26/SUMB[26][22] , \mult_26/SUMB[26][23] ,
         \mult_26/SUMB[26][24] , \mult_26/SUMB[26][25] ,
         \mult_26/SUMB[26][26] , \mult_26/SUMB[26][27] ,
         \mult_26/SUMB[26][28] , \mult_26/SUMB[26][29] ,
         \mult_26/SUMB[26][30] , \mult_26/SUMB[27][1] , \mult_26/SUMB[27][2] ,
         \mult_26/SUMB[27][3] , \mult_26/SUMB[27][4] , \mult_26/SUMB[27][5] ,
         \mult_26/SUMB[27][6] , \mult_26/SUMB[27][7] , \mult_26/SUMB[27][8] ,
         \mult_26/SUMB[27][9] , \mult_26/SUMB[27][10] , \mult_26/SUMB[27][11] ,
         \mult_26/SUMB[27][12] , \mult_26/SUMB[27][13] ,
         \mult_26/SUMB[27][14] , \mult_26/SUMB[27][15] ,
         \mult_26/SUMB[27][16] , \mult_26/SUMB[27][17] ,
         \mult_26/SUMB[27][18] , \mult_26/SUMB[27][19] ,
         \mult_26/SUMB[27][20] , \mult_26/SUMB[27][21] ,
         \mult_26/SUMB[27][22] , \mult_26/SUMB[27][23] ,
         \mult_26/SUMB[27][24] , \mult_26/SUMB[27][25] ,
         \mult_26/SUMB[27][26] , \mult_26/SUMB[27][27] ,
         \mult_26/SUMB[27][28] , \mult_26/SUMB[27][29] ,
         \mult_26/SUMB[27][30] , \mult_26/SUMB[28][1] , \mult_26/SUMB[28][2] ,
         \mult_26/SUMB[28][3] , \mult_26/SUMB[28][4] , \mult_26/SUMB[28][5] ,
         \mult_26/SUMB[28][6] , \mult_26/SUMB[28][7] , \mult_26/SUMB[28][8] ,
         \mult_26/SUMB[28][9] , \mult_26/SUMB[28][10] , \mult_26/SUMB[28][11] ,
         \mult_26/SUMB[28][12] , \mult_26/SUMB[28][13] ,
         \mult_26/SUMB[28][14] , \mult_26/SUMB[28][15] ,
         \mult_26/SUMB[28][16] , \mult_26/SUMB[28][17] ,
         \mult_26/SUMB[28][18] , \mult_26/SUMB[28][19] ,
         \mult_26/SUMB[28][20] , \mult_26/SUMB[28][21] ,
         \mult_26/SUMB[28][22] , \mult_26/SUMB[28][23] ,
         \mult_26/SUMB[28][24] , \mult_26/SUMB[28][25] ,
         \mult_26/SUMB[28][26] , \mult_26/SUMB[28][27] ,
         \mult_26/SUMB[28][28] , \mult_26/SUMB[28][29] ,
         \mult_26/SUMB[28][30] , \mult_26/SUMB[29][1] , \mult_26/SUMB[29][2] ,
         \mult_26/SUMB[29][3] , \mult_26/SUMB[29][4] , \mult_26/SUMB[29][5] ,
         \mult_26/SUMB[29][6] , \mult_26/SUMB[29][7] , \mult_26/SUMB[29][8] ,
         \mult_26/SUMB[29][9] , \mult_26/SUMB[29][10] , \mult_26/SUMB[29][11] ,
         \mult_26/SUMB[29][12] , \mult_26/SUMB[29][13] ,
         \mult_26/SUMB[29][14] , \mult_26/SUMB[29][15] ,
         \mult_26/SUMB[29][16] , \mult_26/SUMB[29][17] ,
         \mult_26/SUMB[29][18] , \mult_26/SUMB[29][19] ,
         \mult_26/SUMB[29][20] , \mult_26/SUMB[29][21] ,
         \mult_26/SUMB[29][22] , \mult_26/SUMB[29][23] ,
         \mult_26/SUMB[29][24] , \mult_26/SUMB[29][25] ,
         \mult_26/SUMB[29][26] , \mult_26/SUMB[29][27] ,
         \mult_26/SUMB[29][28] , \mult_26/SUMB[29][29] ,
         \mult_26/SUMB[29][30] , \mult_26/SUMB[30][1] , \mult_26/SUMB[30][2] ,
         \mult_26/SUMB[30][3] , \mult_26/SUMB[30][4] , \mult_26/SUMB[30][5] ,
         \mult_26/SUMB[30][6] , \mult_26/SUMB[30][7] , \mult_26/SUMB[30][8] ,
         \mult_26/SUMB[30][9] , \mult_26/SUMB[30][10] , \mult_26/SUMB[30][11] ,
         \mult_26/SUMB[30][12] , \mult_26/SUMB[30][13] ,
         \mult_26/SUMB[30][14] , \mult_26/SUMB[30][15] ,
         \mult_26/SUMB[30][16] , \mult_26/SUMB[30][17] ,
         \mult_26/SUMB[30][18] , \mult_26/SUMB[30][19] ,
         \mult_26/SUMB[30][20] , \mult_26/SUMB[30][21] ,
         \mult_26/SUMB[30][22] , \mult_26/SUMB[30][23] ,
         \mult_26/SUMB[30][24] , \mult_26/SUMB[30][25] ,
         \mult_26/SUMB[30][26] , \mult_26/SUMB[30][27] ,
         \mult_26/SUMB[30][28] , \mult_26/SUMB[30][29] ,
         \mult_26/SUMB[30][30] , \mult_26/SUMB[31][0] , \mult_26/SUMB[31][1] ,
         \mult_26/SUMB[31][2] , \mult_26/SUMB[31][3] , \mult_26/SUMB[31][4] ,
         \mult_26/SUMB[31][5] , \mult_26/SUMB[31][6] , \mult_26/SUMB[31][7] ,
         \mult_26/SUMB[31][8] , \mult_26/SUMB[31][9] , \mult_26/SUMB[31][10] ,
         \mult_26/SUMB[31][11] , \mult_26/SUMB[31][12] ,
         \mult_26/SUMB[31][13] , \mult_26/SUMB[31][14] ,
         \mult_26/SUMB[31][15] , \mult_26/SUMB[31][16] ,
         \mult_26/SUMB[31][17] , \mult_26/SUMB[31][18] ,
         \mult_26/SUMB[31][19] , \mult_26/SUMB[31][20] ,
         \mult_26/SUMB[31][21] , \mult_26/SUMB[31][22] ,
         \mult_26/SUMB[31][23] , \mult_26/SUMB[31][24] ,
         \mult_26/SUMB[31][25] , \mult_26/SUMB[31][26] ,
         \mult_26/SUMB[31][27] , \mult_26/SUMB[31][28] ,
         \mult_26/SUMB[31][29] , \mult_26/SUMB[31][30] ,
         \mult_26/CARRYB[16][0] , \mult_26/CARRYB[16][1] ,
         \mult_26/CARRYB[16][2] , \mult_26/CARRYB[16][3] ,
         \mult_26/CARRYB[16][4] , \mult_26/CARRYB[16][5] ,
         \mult_26/CARRYB[16][6] , \mult_26/CARRYB[16][7] ,
         \mult_26/CARRYB[16][8] , \mult_26/CARRYB[16][9] ,
         \mult_26/CARRYB[16][10] , \mult_26/CARRYB[16][11] ,
         \mult_26/CARRYB[16][12] , \mult_26/CARRYB[16][13] ,
         \mult_26/CARRYB[16][14] , \mult_26/CARRYB[16][15] ,
         \mult_26/CARRYB[16][16] , \mult_26/CARRYB[16][17] ,
         \mult_26/CARRYB[16][18] , \mult_26/CARRYB[16][19] ,
         \mult_26/CARRYB[16][20] , \mult_26/CARRYB[16][21] ,
         \mult_26/CARRYB[16][22] , \mult_26/CARRYB[16][23] ,
         \mult_26/CARRYB[16][24] , \mult_26/CARRYB[16][25] ,
         \mult_26/CARRYB[16][26] , \mult_26/CARRYB[16][27] ,
         \mult_26/CARRYB[16][28] , \mult_26/CARRYB[16][29] ,
         \mult_26/CARRYB[16][30] , \mult_26/CARRYB[17][0] ,
         \mult_26/CARRYB[17][1] , \mult_26/CARRYB[17][2] ,
         \mult_26/CARRYB[17][3] , \mult_26/CARRYB[17][4] ,
         \mult_26/CARRYB[17][5] , \mult_26/CARRYB[17][6] ,
         \mult_26/CARRYB[17][7] , \mult_26/CARRYB[17][8] ,
         \mult_26/CARRYB[17][9] , \mult_26/CARRYB[17][10] ,
         \mult_26/CARRYB[17][11] , \mult_26/CARRYB[17][12] ,
         \mult_26/CARRYB[17][13] , \mult_26/CARRYB[17][14] ,
         \mult_26/CARRYB[17][15] , \mult_26/CARRYB[17][16] ,
         \mult_26/CARRYB[17][17] , \mult_26/CARRYB[17][18] ,
         \mult_26/CARRYB[17][19] , \mult_26/CARRYB[17][20] ,
         \mult_26/CARRYB[17][21] , \mult_26/CARRYB[17][22] ,
         \mult_26/CARRYB[17][23] , \mult_26/CARRYB[17][24] ,
         \mult_26/CARRYB[17][25] , \mult_26/CARRYB[17][26] ,
         \mult_26/CARRYB[17][27] , \mult_26/CARRYB[17][28] ,
         \mult_26/CARRYB[17][29] , \mult_26/CARRYB[17][30] ,
         \mult_26/CARRYB[18][0] , \mult_26/CARRYB[18][1] ,
         \mult_26/CARRYB[18][2] , \mult_26/CARRYB[18][3] ,
         \mult_26/CARRYB[18][4] , \mult_26/CARRYB[18][5] ,
         \mult_26/CARRYB[18][6] , \mult_26/CARRYB[18][7] ,
         \mult_26/CARRYB[18][8] , \mult_26/CARRYB[18][9] ,
         \mult_26/CARRYB[18][10] , \mult_26/CARRYB[18][11] ,
         \mult_26/CARRYB[18][12] , \mult_26/CARRYB[18][13] ,
         \mult_26/CARRYB[18][14] , \mult_26/CARRYB[18][15] ,
         \mult_26/CARRYB[18][16] , \mult_26/CARRYB[18][17] ,
         \mult_26/CARRYB[18][18] , \mult_26/CARRYB[18][19] ,
         \mult_26/CARRYB[18][20] , \mult_26/CARRYB[18][21] ,
         \mult_26/CARRYB[18][22] , \mult_26/CARRYB[18][23] ,
         \mult_26/CARRYB[18][24] , \mult_26/CARRYB[18][25] ,
         \mult_26/CARRYB[18][26] , \mult_26/CARRYB[18][27] ,
         \mult_26/CARRYB[18][28] , \mult_26/CARRYB[18][29] ,
         \mult_26/CARRYB[18][30] , \mult_26/CARRYB[19][0] ,
         \mult_26/CARRYB[19][1] , \mult_26/CARRYB[19][2] ,
         \mult_26/CARRYB[19][3] , \mult_26/CARRYB[19][4] ,
         \mult_26/CARRYB[19][5] , \mult_26/CARRYB[19][6] ,
         \mult_26/CARRYB[19][7] , \mult_26/CARRYB[19][8] ,
         \mult_26/CARRYB[19][9] , \mult_26/CARRYB[19][10] ,
         \mult_26/CARRYB[19][11] , \mult_26/CARRYB[19][12] ,
         \mult_26/CARRYB[19][13] , \mult_26/CARRYB[19][14] ,
         \mult_26/CARRYB[19][15] , \mult_26/CARRYB[19][16] ,
         \mult_26/CARRYB[19][17] , \mult_26/CARRYB[19][18] ,
         \mult_26/CARRYB[19][19] , \mult_26/CARRYB[19][20] ,
         \mult_26/CARRYB[19][21] , \mult_26/CARRYB[19][22] ,
         \mult_26/CARRYB[19][23] , \mult_26/CARRYB[19][24] ,
         \mult_26/CARRYB[19][25] , \mult_26/CARRYB[19][26] ,
         \mult_26/CARRYB[19][27] , \mult_26/CARRYB[19][28] ,
         \mult_26/CARRYB[19][29] , \mult_26/CARRYB[19][30] ,
         \mult_26/CARRYB[20][0] , \mult_26/CARRYB[20][1] ,
         \mult_26/CARRYB[20][2] , \mult_26/CARRYB[20][3] ,
         \mult_26/CARRYB[20][4] , \mult_26/CARRYB[20][5] ,
         \mult_26/CARRYB[20][6] , \mult_26/CARRYB[20][7] ,
         \mult_26/CARRYB[20][8] , \mult_26/CARRYB[20][9] ,
         \mult_26/CARRYB[20][10] , \mult_26/CARRYB[20][11] ,
         \mult_26/CARRYB[20][12] , \mult_26/CARRYB[20][13] ,
         \mult_26/CARRYB[20][14] , \mult_26/CARRYB[20][15] ,
         \mult_26/CARRYB[20][16] , \mult_26/CARRYB[20][17] ,
         \mult_26/CARRYB[20][18] , \mult_26/CARRYB[20][19] ,
         \mult_26/CARRYB[20][20] , \mult_26/CARRYB[20][21] ,
         \mult_26/CARRYB[20][22] , \mult_26/CARRYB[20][23] ,
         \mult_26/CARRYB[20][24] , \mult_26/CARRYB[20][25] ,
         \mult_26/CARRYB[20][26] , \mult_26/CARRYB[20][27] ,
         \mult_26/CARRYB[20][28] , \mult_26/CARRYB[20][29] ,
         \mult_26/CARRYB[20][30] , \mult_26/CARRYB[21][0] ,
         \mult_26/CARRYB[21][1] , \mult_26/CARRYB[21][2] ,
         \mult_26/CARRYB[21][3] , \mult_26/CARRYB[21][4] ,
         \mult_26/CARRYB[21][5] , \mult_26/CARRYB[21][6] ,
         \mult_26/CARRYB[21][7] , \mult_26/CARRYB[21][8] ,
         \mult_26/CARRYB[21][9] , \mult_26/CARRYB[21][10] ,
         \mult_26/CARRYB[21][11] , \mult_26/CARRYB[21][12] ,
         \mult_26/CARRYB[21][13] , \mult_26/CARRYB[21][14] ,
         \mult_26/CARRYB[21][15] , \mult_26/CARRYB[21][16] ,
         \mult_26/CARRYB[21][17] , \mult_26/CARRYB[21][18] ,
         \mult_26/CARRYB[21][19] , \mult_26/CARRYB[21][20] ,
         \mult_26/CARRYB[21][21] , \mult_26/CARRYB[21][22] ,
         \mult_26/CARRYB[21][23] , \mult_26/CARRYB[21][24] ,
         \mult_26/CARRYB[21][25] , \mult_26/CARRYB[21][26] ,
         \mult_26/CARRYB[21][27] , \mult_26/CARRYB[21][28] ,
         \mult_26/CARRYB[21][29] , \mult_26/CARRYB[21][30] ,
         \mult_26/CARRYB[22][0] , \mult_26/CARRYB[22][1] ,
         \mult_26/CARRYB[22][2] , \mult_26/CARRYB[22][3] ,
         \mult_26/CARRYB[22][4] , \mult_26/CARRYB[22][5] ,
         \mult_26/CARRYB[22][6] , \mult_26/CARRYB[22][7] ,
         \mult_26/CARRYB[22][8] , \mult_26/CARRYB[22][9] ,
         \mult_26/CARRYB[22][10] , \mult_26/CARRYB[22][11] ,
         \mult_26/CARRYB[22][12] , \mult_26/CARRYB[22][13] ,
         \mult_26/CARRYB[22][14] , \mult_26/CARRYB[22][15] ,
         \mult_26/CARRYB[22][16] , \mult_26/CARRYB[22][17] ,
         \mult_26/CARRYB[22][18] , \mult_26/CARRYB[22][19] ,
         \mult_26/CARRYB[22][20] , \mult_26/CARRYB[22][21] ,
         \mult_26/CARRYB[22][22] , \mult_26/CARRYB[22][23] ,
         \mult_26/CARRYB[22][24] , \mult_26/CARRYB[22][25] ,
         \mult_26/CARRYB[22][26] , \mult_26/CARRYB[22][27] ,
         \mult_26/CARRYB[22][28] , \mult_26/CARRYB[22][29] ,
         \mult_26/CARRYB[22][30] , \mult_26/CARRYB[23][0] ,
         \mult_26/CARRYB[23][1] , \mult_26/CARRYB[23][2] ,
         \mult_26/CARRYB[23][3] , \mult_26/CARRYB[23][4] ,
         \mult_26/CARRYB[23][5] , \mult_26/CARRYB[23][6] ,
         \mult_26/CARRYB[23][7] , \mult_26/CARRYB[23][8] ,
         \mult_26/CARRYB[23][9] , \mult_26/CARRYB[23][10] ,
         \mult_26/CARRYB[23][11] , \mult_26/CARRYB[23][12] ,
         \mult_26/CARRYB[23][13] , \mult_26/CARRYB[23][14] ,
         \mult_26/CARRYB[23][15] , \mult_26/CARRYB[23][16] ,
         \mult_26/CARRYB[23][17] , \mult_26/CARRYB[23][18] ,
         \mult_26/CARRYB[23][19] , \mult_26/CARRYB[23][20] ,
         \mult_26/CARRYB[23][21] , \mult_26/CARRYB[23][22] ,
         \mult_26/CARRYB[23][23] , \mult_26/CARRYB[23][24] ,
         \mult_26/CARRYB[23][25] , \mult_26/CARRYB[23][26] ,
         \mult_26/CARRYB[23][27] , \mult_26/CARRYB[23][28] ,
         \mult_26/CARRYB[23][29] , \mult_26/CARRYB[23][30] ,
         \mult_26/CARRYB[24][0] , \mult_26/CARRYB[24][1] ,
         \mult_26/CARRYB[24][2] , \mult_26/CARRYB[24][3] ,
         \mult_26/CARRYB[24][4] , \mult_26/CARRYB[24][5] ,
         \mult_26/CARRYB[24][6] , \mult_26/CARRYB[24][7] ,
         \mult_26/CARRYB[24][8] , \mult_26/CARRYB[24][9] ,
         \mult_26/CARRYB[24][10] , \mult_26/CARRYB[24][11] ,
         \mult_26/CARRYB[24][12] , \mult_26/CARRYB[24][13] ,
         \mult_26/CARRYB[24][14] , \mult_26/CARRYB[24][15] ,
         \mult_26/CARRYB[24][16] , \mult_26/CARRYB[24][17] ,
         \mult_26/CARRYB[24][18] , \mult_26/CARRYB[24][19] ,
         \mult_26/CARRYB[24][20] , \mult_26/CARRYB[24][21] ,
         \mult_26/CARRYB[24][22] , \mult_26/CARRYB[24][23] ,
         \mult_26/CARRYB[24][24] , \mult_26/CARRYB[24][25] ,
         \mult_26/CARRYB[24][26] , \mult_26/CARRYB[24][27] ,
         \mult_26/CARRYB[24][28] , \mult_26/CARRYB[24][29] ,
         \mult_26/CARRYB[24][30] , \mult_26/CARRYB[25][0] ,
         \mult_26/CARRYB[25][1] , \mult_26/CARRYB[25][2] ,
         \mult_26/CARRYB[25][3] , \mult_26/CARRYB[25][4] ,
         \mult_26/CARRYB[25][5] , \mult_26/CARRYB[25][6] ,
         \mult_26/CARRYB[25][7] , \mult_26/CARRYB[25][8] ,
         \mult_26/CARRYB[25][9] , \mult_26/CARRYB[25][10] ,
         \mult_26/CARRYB[25][11] , \mult_26/CARRYB[25][12] ,
         \mult_26/CARRYB[25][13] , \mult_26/CARRYB[25][14] ,
         \mult_26/CARRYB[25][15] , \mult_26/CARRYB[25][16] ,
         \mult_26/CARRYB[25][17] , \mult_26/CARRYB[25][18] ,
         \mult_26/CARRYB[25][19] , \mult_26/CARRYB[25][20] ,
         \mult_26/CARRYB[25][21] , \mult_26/CARRYB[25][22] ,
         \mult_26/CARRYB[25][23] , \mult_26/CARRYB[25][24] ,
         \mult_26/CARRYB[25][25] , \mult_26/CARRYB[25][26] ,
         \mult_26/CARRYB[25][27] , \mult_26/CARRYB[25][28] ,
         \mult_26/CARRYB[25][29] , \mult_26/CARRYB[25][30] ,
         \mult_26/CARRYB[26][0] , \mult_26/CARRYB[26][1] ,
         \mult_26/CARRYB[26][2] , \mult_26/CARRYB[26][3] ,
         \mult_26/CARRYB[26][4] , \mult_26/CARRYB[26][5] ,
         \mult_26/CARRYB[26][6] , \mult_26/CARRYB[26][7] ,
         \mult_26/CARRYB[26][8] , \mult_26/CARRYB[26][9] ,
         \mult_26/CARRYB[26][10] , \mult_26/CARRYB[26][11] ,
         \mult_26/CARRYB[26][12] , \mult_26/CARRYB[26][13] ,
         \mult_26/CARRYB[26][14] , \mult_26/CARRYB[26][15] ,
         \mult_26/CARRYB[26][16] , \mult_26/CARRYB[26][17] ,
         \mult_26/CARRYB[26][18] , \mult_26/CARRYB[26][19] ,
         \mult_26/CARRYB[26][20] , \mult_26/CARRYB[26][21] ,
         \mult_26/CARRYB[26][22] , \mult_26/CARRYB[26][23] ,
         \mult_26/CARRYB[26][24] , \mult_26/CARRYB[26][25] ,
         \mult_26/CARRYB[26][26] , \mult_26/CARRYB[26][27] ,
         \mult_26/CARRYB[26][28] , \mult_26/CARRYB[26][29] ,
         \mult_26/CARRYB[26][30] , \mult_26/CARRYB[27][0] ,
         \mult_26/CARRYB[27][1] , \mult_26/CARRYB[27][2] ,
         \mult_26/CARRYB[27][3] , \mult_26/CARRYB[27][4] ,
         \mult_26/CARRYB[27][5] , \mult_26/CARRYB[27][6] ,
         \mult_26/CARRYB[27][7] , \mult_26/CARRYB[27][8] ,
         \mult_26/CARRYB[27][9] , \mult_26/CARRYB[27][10] ,
         \mult_26/CARRYB[27][11] , \mult_26/CARRYB[27][12] ,
         \mult_26/CARRYB[27][13] , \mult_26/CARRYB[27][14] ,
         \mult_26/CARRYB[27][15] , \mult_26/CARRYB[27][16] ,
         \mult_26/CARRYB[27][17] , \mult_26/CARRYB[27][18] ,
         \mult_26/CARRYB[27][19] , \mult_26/CARRYB[27][20] ,
         \mult_26/CARRYB[27][21] , \mult_26/CARRYB[27][22] ,
         \mult_26/CARRYB[27][23] , \mult_26/CARRYB[27][24] ,
         \mult_26/CARRYB[27][25] , \mult_26/CARRYB[27][26] ,
         \mult_26/CARRYB[27][27] , \mult_26/CARRYB[27][28] ,
         \mult_26/CARRYB[27][29] , \mult_26/CARRYB[27][30] ,
         \mult_26/CARRYB[28][0] , \mult_26/CARRYB[28][1] ,
         \mult_26/CARRYB[28][2] , \mult_26/CARRYB[28][3] ,
         \mult_26/CARRYB[28][4] , \mult_26/CARRYB[28][5] ,
         \mult_26/CARRYB[28][6] , \mult_26/CARRYB[28][7] ,
         \mult_26/CARRYB[28][8] , \mult_26/CARRYB[28][9] ,
         \mult_26/CARRYB[28][10] , \mult_26/CARRYB[28][11] ,
         \mult_26/CARRYB[28][12] , \mult_26/CARRYB[28][13] ,
         \mult_26/CARRYB[28][14] , \mult_26/CARRYB[28][15] ,
         \mult_26/CARRYB[28][16] , \mult_26/CARRYB[28][17] ,
         \mult_26/CARRYB[28][18] , \mult_26/CARRYB[28][19] ,
         \mult_26/CARRYB[28][20] , \mult_26/CARRYB[28][21] ,
         \mult_26/CARRYB[28][22] , \mult_26/CARRYB[28][23] ,
         \mult_26/CARRYB[28][24] , \mult_26/CARRYB[28][25] ,
         \mult_26/CARRYB[28][26] , \mult_26/CARRYB[28][27] ,
         \mult_26/CARRYB[28][28] , \mult_26/CARRYB[28][29] ,
         \mult_26/CARRYB[28][30] , \mult_26/CARRYB[29][0] ,
         \mult_26/CARRYB[29][1] , \mult_26/CARRYB[29][2] ,
         \mult_26/CARRYB[29][3] , \mult_26/CARRYB[29][4] ,
         \mult_26/CARRYB[29][5] , \mult_26/CARRYB[29][6] ,
         \mult_26/CARRYB[29][7] , \mult_26/CARRYB[29][8] ,
         \mult_26/CARRYB[29][9] , \mult_26/CARRYB[29][10] ,
         \mult_26/CARRYB[29][11] , \mult_26/CARRYB[29][12] ,
         \mult_26/CARRYB[29][13] , \mult_26/CARRYB[29][14] ,
         \mult_26/CARRYB[29][15] , \mult_26/CARRYB[29][16] ,
         \mult_26/CARRYB[29][17] , \mult_26/CARRYB[29][18] ,
         \mult_26/CARRYB[29][19] , \mult_26/CARRYB[29][20] ,
         \mult_26/CARRYB[29][21] , \mult_26/CARRYB[29][22] ,
         \mult_26/CARRYB[29][23] , \mult_26/CARRYB[29][24] ,
         \mult_26/CARRYB[29][25] , \mult_26/CARRYB[29][26] ,
         \mult_26/CARRYB[29][27] , \mult_26/CARRYB[29][28] ,
         \mult_26/CARRYB[29][29] , \mult_26/CARRYB[29][30] ,
         \mult_26/CARRYB[30][0] , \mult_26/CARRYB[30][1] ,
         \mult_26/CARRYB[30][2] , \mult_26/CARRYB[30][3] ,
         \mult_26/CARRYB[30][4] , \mult_26/CARRYB[30][5] ,
         \mult_26/CARRYB[30][6] , \mult_26/CARRYB[30][7] ,
         \mult_26/CARRYB[30][8] , \mult_26/CARRYB[30][9] ,
         \mult_26/CARRYB[30][10] , \mult_26/CARRYB[30][11] ,
         \mult_26/CARRYB[30][12] , \mult_26/CARRYB[30][13] ,
         \mult_26/CARRYB[30][14] , \mult_26/CARRYB[30][15] ,
         \mult_26/CARRYB[30][16] , \mult_26/CARRYB[30][17] ,
         \mult_26/CARRYB[30][18] , \mult_26/CARRYB[30][19] ,
         \mult_26/CARRYB[30][20] , \mult_26/CARRYB[30][21] ,
         \mult_26/CARRYB[30][22] , \mult_26/CARRYB[30][23] ,
         \mult_26/CARRYB[30][24] , \mult_26/CARRYB[30][25] ,
         \mult_26/CARRYB[30][26] , \mult_26/CARRYB[30][27] ,
         \mult_26/CARRYB[30][28] , \mult_26/CARRYB[30][29] ,
         \mult_26/CARRYB[30][30] , \mult_26/CARRYB[31][0] ,
         \mult_26/CARRYB[31][1] , \mult_26/CARRYB[31][2] ,
         \mult_26/CARRYB[31][3] , \mult_26/CARRYB[31][4] ,
         \mult_26/CARRYB[31][5] , \mult_26/CARRYB[31][6] ,
         \mult_26/CARRYB[31][7] , \mult_26/CARRYB[31][8] ,
         \mult_26/CARRYB[31][9] , \mult_26/CARRYB[31][10] ,
         \mult_26/CARRYB[31][11] , \mult_26/CARRYB[31][12] ,
         \mult_26/CARRYB[31][13] , \mult_26/CARRYB[31][14] ,
         \mult_26/CARRYB[31][15] , \mult_26/CARRYB[31][16] ,
         \mult_26/CARRYB[31][17] , \mult_26/CARRYB[31][18] ,
         \mult_26/CARRYB[31][19] , \mult_26/CARRYB[31][20] ,
         \mult_26/CARRYB[31][21] , \mult_26/CARRYB[31][22] ,
         \mult_26/CARRYB[31][23] , \mult_26/CARRYB[31][24] ,
         \mult_26/CARRYB[31][25] , \mult_26/CARRYB[31][26] ,
         \mult_26/CARRYB[31][27] , \mult_26/CARRYB[31][28] ,
         \mult_26/CARRYB[31][29] , \mult_26/CARRYB[31][30] ,
         \mult_26/SUMB[1][1] , \mult_26/SUMB[1][2] , \mult_26/SUMB[1][3] ,
         \mult_26/SUMB[1][4] , \mult_26/SUMB[1][5] , \mult_26/SUMB[1][6] ,
         \mult_26/SUMB[1][7] , \mult_26/SUMB[1][8] , \mult_26/SUMB[1][9] ,
         \mult_26/SUMB[1][10] , \mult_26/SUMB[1][11] , \mult_26/SUMB[1][12] ,
         \mult_26/SUMB[1][13] , \mult_26/SUMB[1][14] , \mult_26/SUMB[1][15] ,
         \mult_26/SUMB[1][16] , \mult_26/SUMB[1][17] , \mult_26/SUMB[1][18] ,
         \mult_26/SUMB[1][19] , \mult_26/SUMB[1][20] , \mult_26/SUMB[1][21] ,
         \mult_26/SUMB[1][22] , \mult_26/SUMB[1][23] , \mult_26/SUMB[1][24] ,
         \mult_26/SUMB[1][25] , \mult_26/SUMB[1][26] , \mult_26/SUMB[1][27] ,
         \mult_26/SUMB[1][28] , \mult_26/SUMB[1][29] , \mult_26/SUMB[1][30] ,
         \mult_26/SUMB[2][1] , \mult_26/SUMB[2][2] , \mult_26/SUMB[2][3] ,
         \mult_26/SUMB[2][4] , \mult_26/SUMB[2][5] , \mult_26/SUMB[2][6] ,
         \mult_26/SUMB[2][7] , \mult_26/SUMB[2][8] , \mult_26/SUMB[2][9] ,
         \mult_26/SUMB[2][10] , \mult_26/SUMB[2][11] , \mult_26/SUMB[2][12] ,
         \mult_26/SUMB[2][13] , \mult_26/SUMB[2][14] , \mult_26/SUMB[2][15] ,
         \mult_26/SUMB[2][16] , \mult_26/SUMB[2][17] , \mult_26/SUMB[2][18] ,
         \mult_26/SUMB[2][19] , \mult_26/SUMB[2][20] , \mult_26/SUMB[2][21] ,
         \mult_26/SUMB[2][22] , \mult_26/SUMB[2][23] , \mult_26/SUMB[2][24] ,
         \mult_26/SUMB[2][25] , \mult_26/SUMB[2][26] , \mult_26/SUMB[2][27] ,
         \mult_26/SUMB[2][28] , \mult_26/SUMB[2][29] , \mult_26/SUMB[2][30] ,
         \mult_26/SUMB[3][1] , \mult_26/SUMB[3][2] , \mult_26/SUMB[3][3] ,
         \mult_26/SUMB[3][4] , \mult_26/SUMB[3][5] , \mult_26/SUMB[3][6] ,
         \mult_26/SUMB[3][7] , \mult_26/SUMB[3][8] , \mult_26/SUMB[3][9] ,
         \mult_26/SUMB[3][10] , \mult_26/SUMB[3][11] , \mult_26/SUMB[3][12] ,
         \mult_26/SUMB[3][13] , \mult_26/SUMB[3][14] , \mult_26/SUMB[3][15] ,
         \mult_26/SUMB[3][16] , \mult_26/SUMB[3][17] , \mult_26/SUMB[3][18] ,
         \mult_26/SUMB[3][19] , \mult_26/SUMB[3][20] , \mult_26/SUMB[3][21] ,
         \mult_26/SUMB[3][22] , \mult_26/SUMB[3][23] , \mult_26/SUMB[3][24] ,
         \mult_26/SUMB[3][25] , \mult_26/SUMB[3][26] , \mult_26/SUMB[3][27] ,
         \mult_26/SUMB[3][28] , \mult_26/SUMB[3][29] , \mult_26/SUMB[3][30] ,
         \mult_26/SUMB[4][1] , \mult_26/SUMB[4][2] , \mult_26/SUMB[4][3] ,
         \mult_26/SUMB[4][4] , \mult_26/SUMB[4][5] , \mult_26/SUMB[4][6] ,
         \mult_26/SUMB[4][7] , \mult_26/SUMB[4][8] , \mult_26/SUMB[4][9] ,
         \mult_26/SUMB[4][10] , \mult_26/SUMB[4][11] , \mult_26/SUMB[4][12] ,
         \mult_26/SUMB[4][13] , \mult_26/SUMB[4][14] , \mult_26/SUMB[4][15] ,
         \mult_26/SUMB[4][16] , \mult_26/SUMB[4][17] , \mult_26/SUMB[4][18] ,
         \mult_26/SUMB[4][19] , \mult_26/SUMB[4][20] , \mult_26/SUMB[4][21] ,
         \mult_26/SUMB[4][22] , \mult_26/SUMB[4][23] , \mult_26/SUMB[4][24] ,
         \mult_26/SUMB[4][25] , \mult_26/SUMB[4][26] , \mult_26/SUMB[4][27] ,
         \mult_26/SUMB[4][28] , \mult_26/SUMB[4][29] , \mult_26/SUMB[4][30] ,
         \mult_26/SUMB[5][1] , \mult_26/SUMB[5][2] , \mult_26/SUMB[5][3] ,
         \mult_26/SUMB[5][4] , \mult_26/SUMB[5][5] , \mult_26/SUMB[5][6] ,
         \mult_26/SUMB[5][7] , \mult_26/SUMB[5][8] , \mult_26/SUMB[5][9] ,
         \mult_26/SUMB[5][10] , \mult_26/SUMB[5][11] , \mult_26/SUMB[5][12] ,
         \mult_26/SUMB[5][13] , \mult_26/SUMB[5][14] , \mult_26/SUMB[5][15] ,
         \mult_26/SUMB[5][16] , \mult_26/SUMB[5][17] , \mult_26/SUMB[5][18] ,
         \mult_26/SUMB[5][19] , \mult_26/SUMB[5][20] , \mult_26/SUMB[5][21] ,
         \mult_26/SUMB[5][22] , \mult_26/SUMB[5][23] , \mult_26/SUMB[5][24] ,
         \mult_26/SUMB[5][25] , \mult_26/SUMB[5][26] , \mult_26/SUMB[5][27] ,
         \mult_26/SUMB[5][28] , \mult_26/SUMB[5][29] , \mult_26/SUMB[5][30] ,
         \mult_26/SUMB[6][1] , \mult_26/SUMB[6][2] , \mult_26/SUMB[6][3] ,
         \mult_26/SUMB[6][4] , \mult_26/SUMB[6][5] , \mult_26/SUMB[6][6] ,
         \mult_26/SUMB[6][7] , \mult_26/SUMB[6][8] , \mult_26/SUMB[6][9] ,
         \mult_26/SUMB[6][10] , \mult_26/SUMB[6][11] , \mult_26/SUMB[6][12] ,
         \mult_26/SUMB[6][13] , \mult_26/SUMB[6][14] , \mult_26/SUMB[6][15] ,
         \mult_26/SUMB[6][16] , \mult_26/SUMB[6][17] , \mult_26/SUMB[6][18] ,
         \mult_26/SUMB[6][19] , \mult_26/SUMB[6][20] , \mult_26/SUMB[6][21] ,
         \mult_26/SUMB[6][22] , \mult_26/SUMB[6][23] , \mult_26/SUMB[6][24] ,
         \mult_26/SUMB[6][25] , \mult_26/SUMB[6][26] , \mult_26/SUMB[6][27] ,
         \mult_26/SUMB[6][28] , \mult_26/SUMB[6][29] , \mult_26/SUMB[6][30] ,
         \mult_26/SUMB[7][1] , \mult_26/SUMB[7][2] , \mult_26/SUMB[7][3] ,
         \mult_26/SUMB[7][4] , \mult_26/SUMB[7][5] , \mult_26/SUMB[7][6] ,
         \mult_26/SUMB[7][7] , \mult_26/SUMB[7][8] , \mult_26/SUMB[7][9] ,
         \mult_26/SUMB[7][10] , \mult_26/SUMB[7][11] , \mult_26/SUMB[7][12] ,
         \mult_26/SUMB[7][13] , \mult_26/SUMB[7][14] , \mult_26/SUMB[7][15] ,
         \mult_26/SUMB[7][16] , \mult_26/SUMB[7][17] , \mult_26/SUMB[7][18] ,
         \mult_26/SUMB[7][19] , \mult_26/SUMB[7][20] , \mult_26/SUMB[7][21] ,
         \mult_26/SUMB[7][22] , \mult_26/SUMB[7][23] , \mult_26/SUMB[7][24] ,
         \mult_26/SUMB[7][25] , \mult_26/SUMB[7][26] , \mult_26/SUMB[7][27] ,
         \mult_26/SUMB[7][28] , \mult_26/SUMB[7][29] , \mult_26/SUMB[7][30] ,
         \mult_26/SUMB[8][1] , \mult_26/SUMB[8][2] , \mult_26/SUMB[8][3] ,
         \mult_26/SUMB[8][4] , \mult_26/SUMB[8][5] , \mult_26/SUMB[8][6] ,
         \mult_26/SUMB[8][7] , \mult_26/SUMB[8][8] , \mult_26/SUMB[8][9] ,
         \mult_26/SUMB[8][10] , \mult_26/SUMB[8][11] , \mult_26/SUMB[8][12] ,
         \mult_26/SUMB[8][13] , \mult_26/SUMB[8][14] , \mult_26/SUMB[8][15] ,
         \mult_26/SUMB[8][16] , \mult_26/SUMB[8][17] , \mult_26/SUMB[8][18] ,
         \mult_26/SUMB[8][19] , \mult_26/SUMB[8][20] , \mult_26/SUMB[8][21] ,
         \mult_26/SUMB[8][22] , \mult_26/SUMB[8][23] , \mult_26/SUMB[8][24] ,
         \mult_26/SUMB[8][25] , \mult_26/SUMB[8][26] , \mult_26/SUMB[8][27] ,
         \mult_26/SUMB[8][28] , \mult_26/SUMB[8][29] , \mult_26/SUMB[8][30] ,
         \mult_26/SUMB[9][1] , \mult_26/SUMB[9][2] , \mult_26/SUMB[9][3] ,
         \mult_26/SUMB[9][4] , \mult_26/SUMB[9][5] , \mult_26/SUMB[9][6] ,
         \mult_26/SUMB[9][7] , \mult_26/SUMB[9][8] , \mult_26/SUMB[9][9] ,
         \mult_26/SUMB[9][10] , \mult_26/SUMB[9][11] , \mult_26/SUMB[9][12] ,
         \mult_26/SUMB[9][13] , \mult_26/SUMB[9][14] , \mult_26/SUMB[9][15] ,
         \mult_26/SUMB[9][16] , \mult_26/SUMB[9][17] , \mult_26/SUMB[9][18] ,
         \mult_26/SUMB[9][19] , \mult_26/SUMB[9][20] , \mult_26/SUMB[9][21] ,
         \mult_26/SUMB[9][22] , \mult_26/SUMB[9][23] , \mult_26/SUMB[9][24] ,
         \mult_26/SUMB[9][25] , \mult_26/SUMB[9][26] , \mult_26/SUMB[9][27] ,
         \mult_26/SUMB[9][28] , \mult_26/SUMB[9][29] , \mult_26/SUMB[9][30] ,
         \mult_26/SUMB[10][1] , \mult_26/SUMB[10][2] , \mult_26/SUMB[10][3] ,
         \mult_26/SUMB[10][4] , \mult_26/SUMB[10][5] , \mult_26/SUMB[10][6] ,
         \mult_26/SUMB[10][7] , \mult_26/SUMB[10][8] , \mult_26/SUMB[10][9] ,
         \mult_26/SUMB[10][10] , \mult_26/SUMB[10][11] ,
         \mult_26/SUMB[10][12] , \mult_26/SUMB[10][13] ,
         \mult_26/SUMB[10][14] , \mult_26/SUMB[10][15] ,
         \mult_26/SUMB[10][16] , \mult_26/SUMB[10][17] ,
         \mult_26/SUMB[10][18] , \mult_26/SUMB[10][19] ,
         \mult_26/SUMB[10][20] , \mult_26/SUMB[10][21] ,
         \mult_26/SUMB[10][22] , \mult_26/SUMB[10][23] ,
         \mult_26/SUMB[10][24] , \mult_26/SUMB[10][25] ,
         \mult_26/SUMB[10][26] , \mult_26/SUMB[10][27] ,
         \mult_26/SUMB[10][28] , \mult_26/SUMB[10][29] ,
         \mult_26/SUMB[10][30] , \mult_26/SUMB[11][1] , \mult_26/SUMB[11][2] ,
         \mult_26/SUMB[11][3] , \mult_26/SUMB[11][4] , \mult_26/SUMB[11][5] ,
         \mult_26/SUMB[11][6] , \mult_26/SUMB[11][7] , \mult_26/SUMB[11][8] ,
         \mult_26/SUMB[11][9] , \mult_26/SUMB[11][10] , \mult_26/SUMB[11][11] ,
         \mult_26/SUMB[11][12] , \mult_26/SUMB[11][13] ,
         \mult_26/SUMB[11][14] , \mult_26/SUMB[11][15] ,
         \mult_26/SUMB[11][16] , \mult_26/SUMB[11][17] ,
         \mult_26/SUMB[11][18] , \mult_26/SUMB[11][19] ,
         \mult_26/SUMB[11][20] , \mult_26/SUMB[11][21] ,
         \mult_26/SUMB[11][22] , \mult_26/SUMB[11][23] ,
         \mult_26/SUMB[11][24] , \mult_26/SUMB[11][25] ,
         \mult_26/SUMB[11][26] , \mult_26/SUMB[11][27] ,
         \mult_26/SUMB[11][28] , \mult_26/SUMB[11][29] ,
         \mult_26/SUMB[11][30] , \mult_26/SUMB[12][1] , \mult_26/SUMB[12][2] ,
         \mult_26/SUMB[12][3] , \mult_26/SUMB[12][4] , \mult_26/SUMB[12][5] ,
         \mult_26/SUMB[12][6] , \mult_26/SUMB[12][7] , \mult_26/SUMB[12][8] ,
         \mult_26/SUMB[12][9] , \mult_26/SUMB[12][10] , \mult_26/SUMB[12][11] ,
         \mult_26/SUMB[12][12] , \mult_26/SUMB[12][13] ,
         \mult_26/SUMB[12][14] , \mult_26/SUMB[12][15] ,
         \mult_26/SUMB[12][16] , \mult_26/SUMB[12][17] ,
         \mult_26/SUMB[12][18] , \mult_26/SUMB[12][19] ,
         \mult_26/SUMB[12][20] , \mult_26/SUMB[12][21] ,
         \mult_26/SUMB[12][22] , \mult_26/SUMB[12][23] ,
         \mult_26/SUMB[12][24] , \mult_26/SUMB[12][25] ,
         \mult_26/SUMB[12][26] , \mult_26/SUMB[12][27] ,
         \mult_26/SUMB[12][28] , \mult_26/SUMB[12][29] ,
         \mult_26/SUMB[12][30] , \mult_26/SUMB[13][1] , \mult_26/SUMB[13][2] ,
         \mult_26/SUMB[13][3] , \mult_26/SUMB[13][4] , \mult_26/SUMB[13][5] ,
         \mult_26/SUMB[13][6] , \mult_26/SUMB[13][7] , \mult_26/SUMB[13][8] ,
         \mult_26/SUMB[13][9] , \mult_26/SUMB[13][10] , \mult_26/SUMB[13][11] ,
         \mult_26/SUMB[13][12] , \mult_26/SUMB[13][13] ,
         \mult_26/SUMB[13][14] , \mult_26/SUMB[13][15] ,
         \mult_26/SUMB[13][16] , \mult_26/SUMB[13][17] ,
         \mult_26/SUMB[13][18] , \mult_26/SUMB[13][19] ,
         \mult_26/SUMB[13][20] , \mult_26/SUMB[13][21] ,
         \mult_26/SUMB[13][22] , \mult_26/SUMB[13][23] ,
         \mult_26/SUMB[13][24] , \mult_26/SUMB[13][25] ,
         \mult_26/SUMB[13][26] , \mult_26/SUMB[13][27] ,
         \mult_26/SUMB[13][28] , \mult_26/SUMB[13][29] ,
         \mult_26/SUMB[13][30] , \mult_26/SUMB[14][1] , \mult_26/SUMB[14][2] ,
         \mult_26/SUMB[14][3] , \mult_26/SUMB[14][4] , \mult_26/SUMB[14][5] ,
         \mult_26/SUMB[14][6] , \mult_26/SUMB[14][7] , \mult_26/SUMB[14][8] ,
         \mult_26/SUMB[14][9] , \mult_26/SUMB[14][10] , \mult_26/SUMB[14][11] ,
         \mult_26/SUMB[14][12] , \mult_26/SUMB[14][13] ,
         \mult_26/SUMB[14][14] , \mult_26/SUMB[14][15] ,
         \mult_26/SUMB[14][16] , \mult_26/SUMB[14][17] ,
         \mult_26/SUMB[14][18] , \mult_26/SUMB[14][19] ,
         \mult_26/SUMB[14][20] , \mult_26/SUMB[14][21] ,
         \mult_26/SUMB[14][22] , \mult_26/SUMB[14][23] ,
         \mult_26/SUMB[14][24] , \mult_26/SUMB[14][25] ,
         \mult_26/SUMB[14][26] , \mult_26/SUMB[14][27] ,
         \mult_26/SUMB[14][28] , \mult_26/SUMB[14][29] ,
         \mult_26/SUMB[14][30] , \mult_26/SUMB[15][1] , \mult_26/SUMB[15][2] ,
         \mult_26/SUMB[15][3] , \mult_26/SUMB[15][4] , \mult_26/SUMB[15][5] ,
         \mult_26/SUMB[15][6] , \mult_26/SUMB[15][7] , \mult_26/SUMB[15][8] ,
         \mult_26/SUMB[15][9] , \mult_26/SUMB[15][10] , \mult_26/SUMB[15][11] ,
         \mult_26/SUMB[15][12] , \mult_26/SUMB[15][13] ,
         \mult_26/SUMB[15][14] , \mult_26/SUMB[15][15] ,
         \mult_26/SUMB[15][16] , \mult_26/SUMB[15][17] ,
         \mult_26/SUMB[15][18] , \mult_26/SUMB[15][19] ,
         \mult_26/SUMB[15][20] , \mult_26/SUMB[15][21] ,
         \mult_26/SUMB[15][22] , \mult_26/SUMB[15][23] ,
         \mult_26/SUMB[15][24] , \mult_26/SUMB[15][25] ,
         \mult_26/SUMB[15][26] , \mult_26/SUMB[15][27] ,
         \mult_26/SUMB[15][28] , \mult_26/SUMB[15][29] ,
         \mult_26/SUMB[15][30] , \mult_26/CARRYB[1][0] ,
         \mult_26/CARRYB[1][1] , \mult_26/CARRYB[1][2] ,
         \mult_26/CARRYB[1][3] , \mult_26/CARRYB[1][4] ,
         \mult_26/CARRYB[1][5] , \mult_26/CARRYB[1][6] ,
         \mult_26/CARRYB[1][7] , \mult_26/CARRYB[1][8] ,
         \mult_26/CARRYB[1][9] , \mult_26/CARRYB[1][10] ,
         \mult_26/CARRYB[1][11] , \mult_26/CARRYB[1][12] ,
         \mult_26/CARRYB[1][13] , \mult_26/CARRYB[1][14] ,
         \mult_26/CARRYB[1][15] , \mult_26/CARRYB[1][16] ,
         \mult_26/CARRYB[1][17] , \mult_26/CARRYB[1][18] ,
         \mult_26/CARRYB[1][19] , \mult_26/CARRYB[1][20] ,
         \mult_26/CARRYB[1][21] , \mult_26/CARRYB[1][22] ,
         \mult_26/CARRYB[1][23] , \mult_26/CARRYB[1][24] ,
         \mult_26/CARRYB[1][25] , \mult_26/CARRYB[1][26] ,
         \mult_26/CARRYB[1][27] , \mult_26/CARRYB[1][28] ,
         \mult_26/CARRYB[1][29] , \mult_26/CARRYB[1][30] ,
         \mult_26/CARRYB[2][0] , \mult_26/CARRYB[2][1] ,
         \mult_26/CARRYB[2][2] , \mult_26/CARRYB[2][3] ,
         \mult_26/CARRYB[2][4] , \mult_26/CARRYB[2][5] ,
         \mult_26/CARRYB[2][6] , \mult_26/CARRYB[2][7] ,
         \mult_26/CARRYB[2][8] , \mult_26/CARRYB[2][9] ,
         \mult_26/CARRYB[2][10] , \mult_26/CARRYB[2][11] ,
         \mult_26/CARRYB[2][12] , \mult_26/CARRYB[2][13] ,
         \mult_26/CARRYB[2][14] , \mult_26/CARRYB[2][15] ,
         \mult_26/CARRYB[2][16] , \mult_26/CARRYB[2][17] ,
         \mult_26/CARRYB[2][18] , \mult_26/CARRYB[2][19] ,
         \mult_26/CARRYB[2][20] , \mult_26/CARRYB[2][21] ,
         \mult_26/CARRYB[2][22] , \mult_26/CARRYB[2][23] ,
         \mult_26/CARRYB[2][24] , \mult_26/CARRYB[2][25] ,
         \mult_26/CARRYB[2][26] , \mult_26/CARRYB[2][27] ,
         \mult_26/CARRYB[2][28] , \mult_26/CARRYB[2][29] ,
         \mult_26/CARRYB[2][30] , \mult_26/CARRYB[3][0] ,
         \mult_26/CARRYB[3][1] , \mult_26/CARRYB[3][2] ,
         \mult_26/CARRYB[3][3] , \mult_26/CARRYB[3][4] ,
         \mult_26/CARRYB[3][5] , \mult_26/CARRYB[3][6] ,
         \mult_26/CARRYB[3][7] , \mult_26/CARRYB[3][8] ,
         \mult_26/CARRYB[3][9] , \mult_26/CARRYB[3][10] ,
         \mult_26/CARRYB[3][11] , \mult_26/CARRYB[3][12] ,
         \mult_26/CARRYB[3][13] , \mult_26/CARRYB[3][14] ,
         \mult_26/CARRYB[3][15] , \mult_26/CARRYB[3][16] ,
         \mult_26/CARRYB[3][17] , \mult_26/CARRYB[3][18] ,
         \mult_26/CARRYB[3][19] , \mult_26/CARRYB[3][20] ,
         \mult_26/CARRYB[3][21] , \mult_26/CARRYB[3][22] ,
         \mult_26/CARRYB[3][23] , \mult_26/CARRYB[3][24] ,
         \mult_26/CARRYB[3][25] , \mult_26/CARRYB[3][26] ,
         \mult_26/CARRYB[3][27] , \mult_26/CARRYB[3][28] ,
         \mult_26/CARRYB[3][29] , \mult_26/CARRYB[3][30] ,
         \mult_26/CARRYB[4][0] , \mult_26/CARRYB[4][1] ,
         \mult_26/CARRYB[4][2] , \mult_26/CARRYB[4][3] ,
         \mult_26/CARRYB[4][4] , \mult_26/CARRYB[4][5] ,
         \mult_26/CARRYB[4][6] , \mult_26/CARRYB[4][7] ,
         \mult_26/CARRYB[4][8] , \mult_26/CARRYB[4][9] ,
         \mult_26/CARRYB[4][10] , \mult_26/CARRYB[4][11] ,
         \mult_26/CARRYB[4][12] , \mult_26/CARRYB[4][13] ,
         \mult_26/CARRYB[4][14] , \mult_26/CARRYB[4][15] ,
         \mult_26/CARRYB[4][16] , \mult_26/CARRYB[4][17] ,
         \mult_26/CARRYB[4][18] , \mult_26/CARRYB[4][19] ,
         \mult_26/CARRYB[4][20] , \mult_26/CARRYB[4][21] ,
         \mult_26/CARRYB[4][22] , \mult_26/CARRYB[4][23] ,
         \mult_26/CARRYB[4][24] , \mult_26/CARRYB[4][25] ,
         \mult_26/CARRYB[4][26] , \mult_26/CARRYB[4][27] ,
         \mult_26/CARRYB[4][28] , \mult_26/CARRYB[4][29] ,
         \mult_26/CARRYB[4][30] , \mult_26/CARRYB[5][0] ,
         \mult_26/CARRYB[5][1] , \mult_26/CARRYB[5][2] ,
         \mult_26/CARRYB[5][3] , \mult_26/CARRYB[5][4] ,
         \mult_26/CARRYB[5][5] , \mult_26/CARRYB[5][6] ,
         \mult_26/CARRYB[5][7] , \mult_26/CARRYB[5][8] ,
         \mult_26/CARRYB[5][9] , \mult_26/CARRYB[5][10] ,
         \mult_26/CARRYB[5][11] , \mult_26/CARRYB[5][12] ,
         \mult_26/CARRYB[5][13] , \mult_26/CARRYB[5][14] ,
         \mult_26/CARRYB[5][15] , \mult_26/CARRYB[5][16] ,
         \mult_26/CARRYB[5][17] , \mult_26/CARRYB[5][18] ,
         \mult_26/CARRYB[5][19] , \mult_26/CARRYB[5][20] ,
         \mult_26/CARRYB[5][21] , \mult_26/CARRYB[5][22] ,
         \mult_26/CARRYB[5][23] , \mult_26/CARRYB[5][24] ,
         \mult_26/CARRYB[5][25] , \mult_26/CARRYB[5][26] ,
         \mult_26/CARRYB[5][27] , \mult_26/CARRYB[5][28] ,
         \mult_26/CARRYB[5][29] , \mult_26/CARRYB[5][30] ,
         \mult_26/CARRYB[6][0] , \mult_26/CARRYB[6][1] ,
         \mult_26/CARRYB[6][2] , \mult_26/CARRYB[6][3] ,
         \mult_26/CARRYB[6][4] , \mult_26/CARRYB[6][5] ,
         \mult_26/CARRYB[6][6] , \mult_26/CARRYB[6][7] ,
         \mult_26/CARRYB[6][8] , \mult_26/CARRYB[6][9] ,
         \mult_26/CARRYB[6][10] , \mult_26/CARRYB[6][11] ,
         \mult_26/CARRYB[6][12] , \mult_26/CARRYB[6][13] ,
         \mult_26/CARRYB[6][14] , \mult_26/CARRYB[6][15] ,
         \mult_26/CARRYB[6][16] , \mult_26/CARRYB[6][17] ,
         \mult_26/CARRYB[6][18] , \mult_26/CARRYB[6][19] ,
         \mult_26/CARRYB[6][20] , \mult_26/CARRYB[6][21] ,
         \mult_26/CARRYB[6][22] , \mult_26/CARRYB[6][23] ,
         \mult_26/CARRYB[6][24] , \mult_26/CARRYB[6][25] ,
         \mult_26/CARRYB[6][26] , \mult_26/CARRYB[6][27] ,
         \mult_26/CARRYB[6][28] , \mult_26/CARRYB[6][29] ,
         \mult_26/CARRYB[6][30] , \mult_26/CARRYB[7][0] ,
         \mult_26/CARRYB[7][1] , \mult_26/CARRYB[7][2] ,
         \mult_26/CARRYB[7][3] , \mult_26/CARRYB[7][4] ,
         \mult_26/CARRYB[7][5] , \mult_26/CARRYB[7][6] ,
         \mult_26/CARRYB[7][7] , \mult_26/CARRYB[7][8] ,
         \mult_26/CARRYB[7][9] , \mult_26/CARRYB[7][10] ,
         \mult_26/CARRYB[7][11] , \mult_26/CARRYB[7][12] ,
         \mult_26/CARRYB[7][13] , \mult_26/CARRYB[7][14] ,
         \mult_26/CARRYB[7][15] , \mult_26/CARRYB[7][16] ,
         \mult_26/CARRYB[7][17] , \mult_26/CARRYB[7][18] ,
         \mult_26/CARRYB[7][19] , \mult_26/CARRYB[7][20] ,
         \mult_26/CARRYB[7][21] , \mult_26/CARRYB[7][22] ,
         \mult_26/CARRYB[7][23] , \mult_26/CARRYB[7][24] ,
         \mult_26/CARRYB[7][25] , \mult_26/CARRYB[7][26] ,
         \mult_26/CARRYB[7][27] , \mult_26/CARRYB[7][28] ,
         \mult_26/CARRYB[7][29] , \mult_26/CARRYB[7][30] ,
         \mult_26/CARRYB[8][0] , \mult_26/CARRYB[8][1] ,
         \mult_26/CARRYB[8][2] , \mult_26/CARRYB[8][3] ,
         \mult_26/CARRYB[8][4] , \mult_26/CARRYB[8][5] ,
         \mult_26/CARRYB[8][6] , \mult_26/CARRYB[8][7] ,
         \mult_26/CARRYB[8][8] , \mult_26/CARRYB[8][9] ,
         \mult_26/CARRYB[8][10] , \mult_26/CARRYB[8][11] ,
         \mult_26/CARRYB[8][12] , \mult_26/CARRYB[8][13] ,
         \mult_26/CARRYB[8][14] , \mult_26/CARRYB[8][15] ,
         \mult_26/CARRYB[8][16] , \mult_26/CARRYB[8][17] ,
         \mult_26/CARRYB[8][18] , \mult_26/CARRYB[8][19] ,
         \mult_26/CARRYB[8][20] , \mult_26/CARRYB[8][21] ,
         \mult_26/CARRYB[8][22] , \mult_26/CARRYB[8][23] ,
         \mult_26/CARRYB[8][24] , \mult_26/CARRYB[8][25] ,
         \mult_26/CARRYB[8][26] , \mult_26/CARRYB[8][27] ,
         \mult_26/CARRYB[8][28] , \mult_26/CARRYB[8][29] ,
         \mult_26/CARRYB[8][30] , \mult_26/CARRYB[9][0] ,
         \mult_26/CARRYB[9][1] , \mult_26/CARRYB[9][2] ,
         \mult_26/CARRYB[9][3] , \mult_26/CARRYB[9][4] ,
         \mult_26/CARRYB[9][5] , \mult_26/CARRYB[9][6] ,
         \mult_26/CARRYB[9][7] , \mult_26/CARRYB[9][8] ,
         \mult_26/CARRYB[9][9] , \mult_26/CARRYB[9][10] ,
         \mult_26/CARRYB[9][11] , \mult_26/CARRYB[9][12] ,
         \mult_26/CARRYB[9][13] , \mult_26/CARRYB[9][14] ,
         \mult_26/CARRYB[9][15] , \mult_26/CARRYB[9][16] ,
         \mult_26/CARRYB[9][17] , \mult_26/CARRYB[9][18] ,
         \mult_26/CARRYB[9][19] , \mult_26/CARRYB[9][20] ,
         \mult_26/CARRYB[9][21] , \mult_26/CARRYB[9][22] ,
         \mult_26/CARRYB[9][23] , \mult_26/CARRYB[9][24] ,
         \mult_26/CARRYB[9][25] , \mult_26/CARRYB[9][26] ,
         \mult_26/CARRYB[9][27] , \mult_26/CARRYB[9][28] ,
         \mult_26/CARRYB[9][29] , \mult_26/CARRYB[9][30] ,
         \mult_26/CARRYB[10][0] , \mult_26/CARRYB[10][1] ,
         \mult_26/CARRYB[10][2] , \mult_26/CARRYB[10][3] ,
         \mult_26/CARRYB[10][4] , \mult_26/CARRYB[10][5] ,
         \mult_26/CARRYB[10][6] , \mult_26/CARRYB[10][7] ,
         \mult_26/CARRYB[10][8] , \mult_26/CARRYB[10][9] ,
         \mult_26/CARRYB[10][10] , \mult_26/CARRYB[10][11] ,
         \mult_26/CARRYB[10][12] , \mult_26/CARRYB[10][13] ,
         \mult_26/CARRYB[10][14] , \mult_26/CARRYB[10][15] ,
         \mult_26/CARRYB[10][16] , \mult_26/CARRYB[10][17] ,
         \mult_26/CARRYB[10][18] , \mult_26/CARRYB[10][19] ,
         \mult_26/CARRYB[10][20] , \mult_26/CARRYB[10][21] ,
         \mult_26/CARRYB[10][22] , \mult_26/CARRYB[10][23] ,
         \mult_26/CARRYB[10][24] , \mult_26/CARRYB[10][25] ,
         \mult_26/CARRYB[10][26] , \mult_26/CARRYB[10][27] ,
         \mult_26/CARRYB[10][28] , \mult_26/CARRYB[10][29] ,
         \mult_26/CARRYB[10][30] , \mult_26/CARRYB[11][0] ,
         \mult_26/CARRYB[11][1] , \mult_26/CARRYB[11][2] ,
         \mult_26/CARRYB[11][3] , \mult_26/CARRYB[11][4] ,
         \mult_26/CARRYB[11][5] , \mult_26/CARRYB[11][6] ,
         \mult_26/CARRYB[11][7] , \mult_26/CARRYB[11][8] ,
         \mult_26/CARRYB[11][9] , \mult_26/CARRYB[11][10] ,
         \mult_26/CARRYB[11][11] , \mult_26/CARRYB[11][12] ,
         \mult_26/CARRYB[11][13] , \mult_26/CARRYB[11][14] ,
         \mult_26/CARRYB[11][15] , \mult_26/CARRYB[11][16] ,
         \mult_26/CARRYB[11][17] , \mult_26/CARRYB[11][18] ,
         \mult_26/CARRYB[11][19] , \mult_26/CARRYB[11][20] ,
         \mult_26/CARRYB[11][21] , \mult_26/CARRYB[11][22] ,
         \mult_26/CARRYB[11][23] , \mult_26/CARRYB[11][24] ,
         \mult_26/CARRYB[11][25] , \mult_26/CARRYB[11][26] ,
         \mult_26/CARRYB[11][27] , \mult_26/CARRYB[11][28] ,
         \mult_26/CARRYB[11][29] , \mult_26/CARRYB[11][30] ,
         \mult_26/CARRYB[12][0] , \mult_26/CARRYB[12][1] ,
         \mult_26/CARRYB[12][2] , \mult_26/CARRYB[12][3] ,
         \mult_26/CARRYB[12][4] , \mult_26/CARRYB[12][5] ,
         \mult_26/CARRYB[12][6] , \mult_26/CARRYB[12][7] ,
         \mult_26/CARRYB[12][8] , \mult_26/CARRYB[12][9] ,
         \mult_26/CARRYB[12][10] , \mult_26/CARRYB[12][11] ,
         \mult_26/CARRYB[12][12] , \mult_26/CARRYB[12][13] ,
         \mult_26/CARRYB[12][14] , \mult_26/CARRYB[12][15] ,
         \mult_26/CARRYB[12][16] , \mult_26/CARRYB[12][17] ,
         \mult_26/CARRYB[12][18] , \mult_26/CARRYB[12][19] ,
         \mult_26/CARRYB[12][20] , \mult_26/CARRYB[12][21] ,
         \mult_26/CARRYB[12][22] , \mult_26/CARRYB[12][23] ,
         \mult_26/CARRYB[12][24] , \mult_26/CARRYB[12][25] ,
         \mult_26/CARRYB[12][26] , \mult_26/CARRYB[12][27] ,
         \mult_26/CARRYB[12][28] , \mult_26/CARRYB[12][29] ,
         \mult_26/CARRYB[12][30] , \mult_26/CARRYB[13][0] ,
         \mult_26/CARRYB[13][1] , \mult_26/CARRYB[13][2] ,
         \mult_26/CARRYB[13][3] , \mult_26/CARRYB[13][4] ,
         \mult_26/CARRYB[13][5] , \mult_26/CARRYB[13][6] ,
         \mult_26/CARRYB[13][7] , \mult_26/CARRYB[13][8] ,
         \mult_26/CARRYB[13][9] , \mult_26/CARRYB[13][10] ,
         \mult_26/CARRYB[13][11] , \mult_26/CARRYB[13][12] ,
         \mult_26/CARRYB[13][13] , \mult_26/CARRYB[13][14] ,
         \mult_26/CARRYB[13][15] , \mult_26/CARRYB[13][16] ,
         \mult_26/CARRYB[13][17] , \mult_26/CARRYB[13][18] ,
         \mult_26/CARRYB[13][19] , \mult_26/CARRYB[13][20] ,
         \mult_26/CARRYB[13][21] , \mult_26/CARRYB[13][22] ,
         \mult_26/CARRYB[13][23] , \mult_26/CARRYB[13][24] ,
         \mult_26/CARRYB[13][25] , \mult_26/CARRYB[13][26] ,
         \mult_26/CARRYB[13][27] , \mult_26/CARRYB[13][28] ,
         \mult_26/CARRYB[13][29] , \mult_26/CARRYB[13][30] ,
         \mult_26/CARRYB[14][0] , \mult_26/CARRYB[14][1] ,
         \mult_26/CARRYB[14][2] , \mult_26/CARRYB[14][3] ,
         \mult_26/CARRYB[14][4] , \mult_26/CARRYB[14][5] ,
         \mult_26/CARRYB[14][6] , \mult_26/CARRYB[14][7] ,
         \mult_26/CARRYB[14][8] , \mult_26/CARRYB[14][9] ,
         \mult_26/CARRYB[14][10] , \mult_26/CARRYB[14][11] ,
         \mult_26/CARRYB[14][12] , \mult_26/CARRYB[14][13] ,
         \mult_26/CARRYB[14][14] , \mult_26/CARRYB[14][15] ,
         \mult_26/CARRYB[14][16] , \mult_26/CARRYB[14][17] ,
         \mult_26/CARRYB[14][18] , \mult_26/CARRYB[14][19] ,
         \mult_26/CARRYB[14][20] , \mult_26/CARRYB[14][21] ,
         \mult_26/CARRYB[14][22] , \mult_26/CARRYB[14][23] ,
         \mult_26/CARRYB[14][24] , \mult_26/CARRYB[14][25] ,
         \mult_26/CARRYB[14][26] , \mult_26/CARRYB[14][27] ,
         \mult_26/CARRYB[14][28] , \mult_26/CARRYB[14][29] ,
         \mult_26/CARRYB[14][30] , \mult_26/CARRYB[15][0] ,
         \mult_26/CARRYB[15][1] , \mult_26/CARRYB[15][2] ,
         \mult_26/CARRYB[15][3] , \mult_26/CARRYB[15][4] ,
         \mult_26/CARRYB[15][5] , \mult_26/CARRYB[15][6] ,
         \mult_26/CARRYB[15][7] , \mult_26/CARRYB[15][8] ,
         \mult_26/CARRYB[15][9] , \mult_26/CARRYB[15][10] ,
         \mult_26/CARRYB[15][11] , \mult_26/CARRYB[15][12] ,
         \mult_26/CARRYB[15][13] , \mult_26/CARRYB[15][14] ,
         \mult_26/CARRYB[15][15] , \mult_26/CARRYB[15][16] ,
         \mult_26/CARRYB[15][17] , \mult_26/CARRYB[15][18] ,
         \mult_26/CARRYB[15][19] , \mult_26/CARRYB[15][20] ,
         \mult_26/CARRYB[15][21] , \mult_26/CARRYB[15][22] ,
         \mult_26/CARRYB[15][23] , \mult_26/CARRYB[15][24] ,
         \mult_26/CARRYB[15][25] , \mult_26/CARRYB[15][26] ,
         \mult_26/CARRYB[15][27] , \mult_26/CARRYB[15][28] ,
         \mult_26/CARRYB[15][29] , \mult_26/CARRYB[15][30] ,
         \mult_26/ab[0][1] , \mult_26/ab[0][2] , \mult_26/ab[0][3] ,
         \mult_26/ab[0][4] , \mult_26/ab[0][5] , \mult_26/ab[0][6] ,
         \mult_26/ab[0][7] , \mult_26/ab[0][8] , \mult_26/ab[0][9] ,
         \mult_26/ab[0][10] , \mult_26/ab[0][11] , \mult_26/ab[0][12] ,
         \mult_26/ab[0][13] , \mult_26/ab[0][14] , \mult_26/ab[0][15] ,
         \mult_26/ab[0][16] , \mult_26/ab[0][17] , \mult_26/ab[0][18] ,
         \mult_26/ab[0][19] , \mult_26/ab[0][20] , \mult_26/ab[0][21] ,
         \mult_26/ab[0][22] , \mult_26/ab[0][23] , \mult_26/ab[0][24] ,
         \mult_26/ab[0][25] , \mult_26/ab[0][26] , \mult_26/ab[0][27] ,
         \mult_26/ab[0][28] , \mult_26/ab[0][29] , \mult_26/ab[0][30] ,
         \mult_26/ab[0][31] , \mult_26/ab[1][0] , \mult_26/ab[1][1] ,
         \mult_26/ab[1][2] , \mult_26/ab[1][3] , \mult_26/ab[1][4] ,
         \mult_26/ab[1][5] , \mult_26/ab[1][6] , \mult_26/ab[1][7] ,
         \mult_26/ab[1][8] , \mult_26/ab[1][9] , \mult_26/ab[1][10] ,
         \mult_26/ab[1][11] , \mult_26/ab[1][12] , \mult_26/ab[1][13] ,
         \mult_26/ab[1][14] , \mult_26/ab[1][15] , \mult_26/ab[1][16] ,
         \mult_26/ab[1][17] , \mult_26/ab[1][18] , \mult_26/ab[1][19] ,
         \mult_26/ab[1][20] , \mult_26/ab[1][21] , \mult_26/ab[1][22] ,
         \mult_26/ab[1][23] , \mult_26/ab[1][24] , \mult_26/ab[1][25] ,
         \mult_26/ab[1][26] , \mult_26/ab[1][27] , \mult_26/ab[1][28] ,
         \mult_26/ab[1][29] , \mult_26/ab[1][30] , \mult_26/ab[1][31] ,
         \mult_26/ab[2][0] , \mult_26/ab[2][1] , \mult_26/ab[2][2] ,
         \mult_26/ab[2][3] , \mult_26/ab[2][4] , \mult_26/ab[2][5] ,
         \mult_26/ab[2][6] , \mult_26/ab[2][7] , \mult_26/ab[2][8] ,
         \mult_26/ab[2][9] , \mult_26/ab[2][10] , \mult_26/ab[2][11] ,
         \mult_26/ab[2][12] , \mult_26/ab[2][13] , \mult_26/ab[2][14] ,
         \mult_26/ab[2][15] , \mult_26/ab[2][16] , \mult_26/ab[2][17] ,
         \mult_26/ab[2][18] , \mult_26/ab[2][19] , \mult_26/ab[2][20] ,
         \mult_26/ab[2][21] , \mult_26/ab[2][22] , \mult_26/ab[2][23] ,
         \mult_26/ab[2][24] , \mult_26/ab[2][25] , \mult_26/ab[2][26] ,
         \mult_26/ab[2][27] , \mult_26/ab[2][28] , \mult_26/ab[2][29] ,
         \mult_26/ab[2][30] , \mult_26/ab[2][31] , \mult_26/ab[3][0] ,
         \mult_26/ab[3][1] , \mult_26/ab[3][2] , \mult_26/ab[3][3] ,
         \mult_26/ab[3][4] , \mult_26/ab[3][5] , \mult_26/ab[3][6] ,
         \mult_26/ab[3][7] , \mult_26/ab[3][8] , \mult_26/ab[3][9] ,
         \mult_26/ab[3][10] , \mult_26/ab[3][11] , \mult_26/ab[3][12] ,
         \mult_26/ab[3][13] , \mult_26/ab[3][14] , \mult_26/ab[3][15] ,
         \mult_26/ab[3][16] , \mult_26/ab[3][17] , \mult_26/ab[3][18] ,
         \mult_26/ab[3][19] , \mult_26/ab[3][20] , \mult_26/ab[3][21] ,
         \mult_26/ab[3][22] , \mult_26/ab[3][23] , \mult_26/ab[3][24] ,
         \mult_26/ab[3][25] , \mult_26/ab[3][26] , \mult_26/ab[3][27] ,
         \mult_26/ab[3][28] , \mult_26/ab[3][29] , \mult_26/ab[3][30] ,
         \mult_26/ab[3][31] , \mult_26/ab[4][0] , \mult_26/ab[4][1] ,
         \mult_26/ab[4][2] , \mult_26/ab[4][3] , \mult_26/ab[4][4] ,
         \mult_26/ab[4][5] , \mult_26/ab[4][6] , \mult_26/ab[4][7] ,
         \mult_26/ab[4][8] , \mult_26/ab[4][9] , \mult_26/ab[4][10] ,
         \mult_26/ab[4][11] , \mult_26/ab[4][12] , \mult_26/ab[4][13] ,
         \mult_26/ab[4][14] , \mult_26/ab[4][15] , \mult_26/ab[4][16] ,
         \mult_26/ab[4][17] , \mult_26/ab[4][18] , \mult_26/ab[4][19] ,
         \mult_26/ab[4][20] , \mult_26/ab[4][21] , \mult_26/ab[4][22] ,
         \mult_26/ab[4][23] , \mult_26/ab[4][24] , \mult_26/ab[4][25] ,
         \mult_26/ab[4][26] , \mult_26/ab[4][27] , \mult_26/ab[4][28] ,
         \mult_26/ab[4][29] , \mult_26/ab[4][30] , \mult_26/ab[4][31] ,
         \mult_26/ab[5][0] , \mult_26/ab[5][1] , \mult_26/ab[5][2] ,
         \mult_26/ab[5][3] , \mult_26/ab[5][4] , \mult_26/ab[5][5] ,
         \mult_26/ab[5][6] , \mult_26/ab[5][7] , \mult_26/ab[5][8] ,
         \mult_26/ab[5][9] , \mult_26/ab[5][10] , \mult_26/ab[5][11] ,
         \mult_26/ab[5][12] , \mult_26/ab[5][13] , \mult_26/ab[5][14] ,
         \mult_26/ab[5][15] , \mult_26/ab[5][16] , \mult_26/ab[5][17] ,
         \mult_26/ab[5][18] , \mult_26/ab[5][19] , \mult_26/ab[5][20] ,
         \mult_26/ab[5][21] , \mult_26/ab[5][22] , \mult_26/ab[5][23] ,
         \mult_26/ab[5][24] , \mult_26/ab[5][25] , \mult_26/ab[5][26] ,
         \mult_26/ab[5][27] , \mult_26/ab[5][28] , \mult_26/ab[5][29] ,
         \mult_26/ab[5][30] , \mult_26/ab[5][31] , \mult_26/ab[6][0] ,
         \mult_26/ab[6][1] , \mult_26/ab[6][2] , \mult_26/ab[6][3] ,
         \mult_26/ab[6][4] , \mult_26/ab[6][5] , \mult_26/ab[6][6] ,
         \mult_26/ab[6][7] , \mult_26/ab[6][8] , \mult_26/ab[6][9] ,
         \mult_26/ab[6][10] , \mult_26/ab[6][11] , \mult_26/ab[6][12] ,
         \mult_26/ab[6][13] , \mult_26/ab[6][14] , \mult_26/ab[6][15] ,
         \mult_26/ab[6][16] , \mult_26/ab[6][17] , \mult_26/ab[6][18] ,
         \mult_26/ab[6][19] , \mult_26/ab[6][20] , \mult_26/ab[6][21] ,
         \mult_26/ab[6][22] , \mult_26/ab[6][23] , \mult_26/ab[6][24] ,
         \mult_26/ab[6][25] , \mult_26/ab[6][26] , \mult_26/ab[6][27] ,
         \mult_26/ab[6][28] , \mult_26/ab[6][29] , \mult_26/ab[6][30] ,
         \mult_26/ab[6][31] , \mult_26/ab[7][0] , \mult_26/ab[7][1] ,
         \mult_26/ab[7][2] , \mult_26/ab[7][3] , \mult_26/ab[7][4] ,
         \mult_26/ab[7][5] , \mult_26/ab[7][6] , \mult_26/ab[7][7] ,
         \mult_26/ab[7][8] , \mult_26/ab[7][9] , \mult_26/ab[7][10] ,
         \mult_26/ab[7][11] , \mult_26/ab[7][12] , \mult_26/ab[7][13] ,
         \mult_26/ab[7][14] , \mult_26/ab[7][15] , \mult_26/ab[7][16] ,
         \mult_26/ab[7][17] , \mult_26/ab[7][18] , \mult_26/ab[7][19] ,
         \mult_26/ab[7][20] , \mult_26/ab[7][21] , \mult_26/ab[7][22] ,
         \mult_26/ab[7][23] , \mult_26/ab[7][24] , \mult_26/ab[7][25] ,
         \mult_26/ab[7][26] , \mult_26/ab[7][27] , \mult_26/ab[7][28] ,
         \mult_26/ab[7][29] , \mult_26/ab[7][30] , \mult_26/ab[7][31] ,
         \mult_26/ab[8][0] , \mult_26/ab[8][1] , \mult_26/ab[8][2] ,
         \mult_26/ab[8][3] , \mult_26/ab[8][4] , \mult_26/ab[8][5] ,
         \mult_26/ab[8][6] , \mult_26/ab[8][7] , \mult_26/ab[8][8] ,
         \mult_26/ab[8][9] , \mult_26/ab[8][10] , \mult_26/ab[8][11] ,
         \mult_26/ab[8][12] , \mult_26/ab[8][13] , \mult_26/ab[8][14] ,
         \mult_26/ab[8][15] , \mult_26/ab[8][16] , \mult_26/ab[8][17] ,
         \mult_26/ab[8][18] , \mult_26/ab[8][19] , \mult_26/ab[8][20] ,
         \mult_26/ab[8][21] , \mult_26/ab[8][22] , \mult_26/ab[8][23] ,
         \mult_26/ab[8][24] , \mult_26/ab[8][25] , \mult_26/ab[8][26] ,
         \mult_26/ab[8][27] , \mult_26/ab[8][28] , \mult_26/ab[8][29] ,
         \mult_26/ab[8][30] , \mult_26/ab[8][31] , \mult_26/ab[9][0] ,
         \mult_26/ab[9][1] , \mult_26/ab[9][2] , \mult_26/ab[9][3] ,
         \mult_26/ab[9][4] , \mult_26/ab[9][5] , \mult_26/ab[9][6] ,
         \mult_26/ab[9][7] , \mult_26/ab[9][8] , \mult_26/ab[9][9] ,
         \mult_26/ab[9][10] , \mult_26/ab[9][11] , \mult_26/ab[9][12] ,
         \mult_26/ab[9][13] , \mult_26/ab[9][14] , \mult_26/ab[9][15] ,
         \mult_26/ab[9][16] , \mult_26/ab[9][17] , \mult_26/ab[9][18] ,
         \mult_26/ab[9][19] , \mult_26/ab[9][20] , \mult_26/ab[9][21] ,
         \mult_26/ab[9][22] , \mult_26/ab[9][23] , \mult_26/ab[9][24] ,
         \mult_26/ab[9][25] , \mult_26/ab[9][26] , \mult_26/ab[9][27] ,
         \mult_26/ab[9][28] , \mult_26/ab[9][29] , \mult_26/ab[9][30] ,
         \mult_26/ab[9][31] , \mult_26/ab[10][0] , \mult_26/ab[10][1] ,
         \mult_26/ab[10][2] , \mult_26/ab[10][3] , \mult_26/ab[10][4] ,
         \mult_26/ab[10][5] , \mult_26/ab[10][6] , \mult_26/ab[10][7] ,
         \mult_26/ab[10][8] , \mult_26/ab[10][9] , \mult_26/ab[10][10] ,
         \mult_26/ab[10][11] , \mult_26/ab[10][12] , \mult_26/ab[10][13] ,
         \mult_26/ab[10][14] , \mult_26/ab[10][15] , \mult_26/ab[10][16] ,
         \mult_26/ab[10][17] , \mult_26/ab[10][18] , \mult_26/ab[10][19] ,
         \mult_26/ab[10][20] , \mult_26/ab[10][21] , \mult_26/ab[10][22] ,
         \mult_26/ab[10][23] , \mult_26/ab[10][24] , \mult_26/ab[10][25] ,
         \mult_26/ab[10][26] , \mult_26/ab[10][27] , \mult_26/ab[10][28] ,
         \mult_26/ab[10][29] , \mult_26/ab[10][30] , \mult_26/ab[10][31] ,
         \mult_26/ab[11][0] , \mult_26/ab[11][1] , \mult_26/ab[11][2] ,
         \mult_26/ab[11][3] , \mult_26/ab[11][4] , \mult_26/ab[11][5] ,
         \mult_26/ab[11][6] , \mult_26/ab[11][7] , \mult_26/ab[11][8] ,
         \mult_26/ab[11][9] , \mult_26/ab[11][10] , \mult_26/ab[11][11] ,
         \mult_26/ab[11][12] , \mult_26/ab[11][13] , \mult_26/ab[11][14] ,
         \mult_26/ab[11][15] , \mult_26/ab[11][16] , \mult_26/ab[11][17] ,
         \mult_26/ab[11][18] , \mult_26/ab[11][19] , \mult_26/ab[11][20] ,
         \mult_26/ab[11][21] , \mult_26/ab[11][22] , \mult_26/ab[11][23] ,
         \mult_26/ab[11][24] , \mult_26/ab[11][25] , \mult_26/ab[11][26] ,
         \mult_26/ab[11][27] , \mult_26/ab[11][28] , \mult_26/ab[11][29] ,
         \mult_26/ab[11][30] , \mult_26/ab[11][31] , \mult_26/ab[12][0] ,
         \mult_26/ab[12][1] , \mult_26/ab[12][2] , \mult_26/ab[12][3] ,
         \mult_26/ab[12][4] , \mult_26/ab[12][5] , \mult_26/ab[12][6] ,
         \mult_26/ab[12][7] , \mult_26/ab[12][8] , \mult_26/ab[12][9] ,
         \mult_26/ab[12][10] , \mult_26/ab[12][11] , \mult_26/ab[12][12] ,
         \mult_26/ab[12][13] , \mult_26/ab[12][14] , \mult_26/ab[12][15] ,
         \mult_26/ab[12][16] , \mult_26/ab[12][17] , \mult_26/ab[12][18] ,
         \mult_26/ab[12][19] , \mult_26/ab[12][20] , \mult_26/ab[12][21] ,
         \mult_26/ab[12][22] , \mult_26/ab[12][23] , \mult_26/ab[12][24] ,
         \mult_26/ab[12][25] , \mult_26/ab[12][26] , \mult_26/ab[12][27] ,
         \mult_26/ab[12][28] , \mult_26/ab[12][29] , \mult_26/ab[12][30] ,
         \mult_26/ab[12][31] , \mult_26/ab[13][0] , \mult_26/ab[13][1] ,
         \mult_26/ab[13][2] , \mult_26/ab[13][3] , \mult_26/ab[13][4] ,
         \mult_26/ab[13][5] , \mult_26/ab[13][6] , \mult_26/ab[13][7] ,
         \mult_26/ab[13][8] , \mult_26/ab[13][9] , \mult_26/ab[13][10] ,
         \mult_26/ab[13][11] , \mult_26/ab[13][12] , \mult_26/ab[13][13] ,
         \mult_26/ab[13][14] , \mult_26/ab[13][15] , \mult_26/ab[13][16] ,
         \mult_26/ab[13][17] , \mult_26/ab[13][18] , \mult_26/ab[13][19] ,
         \mult_26/ab[13][20] , \mult_26/ab[13][21] , \mult_26/ab[13][22] ,
         \mult_26/ab[13][23] , \mult_26/ab[13][24] , \mult_26/ab[13][25] ,
         \mult_26/ab[13][26] , \mult_26/ab[13][27] , \mult_26/ab[13][28] ,
         \mult_26/ab[13][29] , \mult_26/ab[13][30] , \mult_26/ab[13][31] ,
         \mult_26/ab[14][0] , \mult_26/ab[14][1] , \mult_26/ab[14][2] ,
         \mult_26/ab[14][3] , \mult_26/ab[14][4] , \mult_26/ab[14][5] ,
         \mult_26/ab[14][6] , \mult_26/ab[14][7] , \mult_26/ab[14][8] ,
         \mult_26/ab[14][9] , \mult_26/ab[14][10] , \mult_26/ab[14][11] ,
         \mult_26/ab[14][12] , \mult_26/ab[14][13] , \mult_26/ab[14][14] ,
         \mult_26/ab[14][15] , \mult_26/ab[14][16] , \mult_26/ab[14][17] ,
         \mult_26/ab[14][18] , \mult_26/ab[14][19] , \mult_26/ab[14][20] ,
         \mult_26/ab[14][21] , \mult_26/ab[14][22] , \mult_26/ab[14][23] ,
         \mult_26/ab[14][24] , \mult_26/ab[14][25] , \mult_26/ab[14][26] ,
         \mult_26/ab[14][27] , \mult_26/ab[14][28] , \mult_26/ab[14][29] ,
         \mult_26/ab[14][30] , \mult_26/ab[14][31] , \mult_26/ab[15][0] ,
         \mult_26/ab[15][1] , \mult_26/ab[15][2] , \mult_26/ab[15][3] ,
         \mult_26/ab[15][4] , \mult_26/ab[15][5] , \mult_26/ab[15][6] ,
         \mult_26/ab[15][7] , \mult_26/ab[15][8] , \mult_26/ab[15][9] ,
         \mult_26/ab[15][10] , \mult_26/ab[15][11] , \mult_26/ab[15][12] ,
         \mult_26/ab[15][13] , \mult_26/ab[15][14] , \mult_26/ab[15][15] ,
         \mult_26/ab[15][16] , \mult_26/ab[15][17] , \mult_26/ab[15][18] ,
         \mult_26/ab[15][19] , \mult_26/ab[15][20] , \mult_26/ab[15][21] ,
         \mult_26/ab[15][22] , \mult_26/ab[15][23] , \mult_26/ab[15][24] ,
         \mult_26/ab[15][25] , \mult_26/ab[15][26] , \mult_26/ab[15][27] ,
         \mult_26/ab[15][28] , \mult_26/ab[15][29] , \mult_26/ab[15][30] ,
         \mult_26/ab[15][31] , \mult_26/ab[16][0] , \mult_26/ab[16][1] ,
         \mult_26/ab[16][2] , \mult_26/ab[16][3] , \mult_26/ab[16][4] ,
         \mult_26/ab[16][5] , \mult_26/ab[16][6] , \mult_26/ab[16][7] ,
         \mult_26/ab[16][8] , \mult_26/ab[16][9] , \mult_26/ab[16][10] ,
         \mult_26/ab[16][11] , \mult_26/ab[16][12] , \mult_26/ab[16][13] ,
         \mult_26/ab[16][14] , \mult_26/ab[16][15] , \mult_26/ab[16][16] ,
         \mult_26/ab[16][17] , \mult_26/ab[16][18] , \mult_26/ab[16][19] ,
         \mult_26/ab[16][20] , \mult_26/ab[16][21] , \mult_26/ab[16][22] ,
         \mult_26/ab[16][23] , \mult_26/ab[16][24] , \mult_26/ab[16][25] ,
         \mult_26/ab[16][26] , \mult_26/ab[16][27] , \mult_26/ab[16][28] ,
         \mult_26/ab[16][29] , \mult_26/ab[16][30] , \mult_26/ab[16][31] ,
         \mult_26/ab[17][0] , \mult_26/ab[17][1] , \mult_26/ab[17][2] ,
         \mult_26/ab[17][3] , \mult_26/ab[17][4] , \mult_26/ab[17][5] ,
         \mult_26/ab[17][6] , \mult_26/ab[17][7] , \mult_26/ab[17][8] ,
         \mult_26/ab[17][9] , \mult_26/ab[17][10] , \mult_26/ab[17][11] ,
         \mult_26/ab[17][12] , \mult_26/ab[17][13] , \mult_26/ab[17][14] ,
         \mult_26/ab[17][15] , \mult_26/ab[17][16] , \mult_26/ab[17][17] ,
         \mult_26/ab[17][18] , \mult_26/ab[17][19] , \mult_26/ab[17][20] ,
         \mult_26/ab[17][21] , \mult_26/ab[17][22] , \mult_26/ab[17][23] ,
         \mult_26/ab[17][24] , \mult_26/ab[17][25] , \mult_26/ab[17][26] ,
         \mult_26/ab[17][27] , \mult_26/ab[17][28] , \mult_26/ab[17][29] ,
         \mult_26/ab[17][30] , \mult_26/ab[17][31] , \mult_26/ab[18][0] ,
         \mult_26/ab[18][1] , \mult_26/ab[18][2] , \mult_26/ab[18][3] ,
         \mult_26/ab[18][4] , \mult_26/ab[18][5] , \mult_26/ab[18][6] ,
         \mult_26/ab[18][7] , \mult_26/ab[18][8] , \mult_26/ab[18][9] ,
         \mult_26/ab[18][10] , \mult_26/ab[18][11] , \mult_26/ab[18][12] ,
         \mult_26/ab[18][13] , \mult_26/ab[18][14] , \mult_26/ab[18][15] ,
         \mult_26/ab[18][16] , \mult_26/ab[18][17] , \mult_26/ab[18][18] ,
         \mult_26/ab[18][19] , \mult_26/ab[18][20] , \mult_26/ab[18][21] ,
         \mult_26/ab[18][22] , \mult_26/ab[18][23] , \mult_26/ab[18][24] ,
         \mult_26/ab[18][25] , \mult_26/ab[18][26] , \mult_26/ab[18][27] ,
         \mult_26/ab[18][28] , \mult_26/ab[18][29] , \mult_26/ab[18][30] ,
         \mult_26/ab[18][31] , \mult_26/ab[19][0] , \mult_26/ab[19][1] ,
         \mult_26/ab[19][2] , \mult_26/ab[19][3] , \mult_26/ab[19][4] ,
         \mult_26/ab[19][5] , \mult_26/ab[19][6] , \mult_26/ab[19][7] ,
         \mult_26/ab[19][8] , \mult_26/ab[19][9] , \mult_26/ab[19][10] ,
         \mult_26/ab[19][11] , \mult_26/ab[19][12] , \mult_26/ab[19][13] ,
         \mult_26/ab[19][14] , \mult_26/ab[19][15] , \mult_26/ab[19][16] ,
         \mult_26/ab[19][17] , \mult_26/ab[19][18] , \mult_26/ab[19][19] ,
         \mult_26/ab[19][20] , \mult_26/ab[19][21] , \mult_26/ab[19][22] ,
         \mult_26/ab[19][23] , \mult_26/ab[19][24] , \mult_26/ab[19][25] ,
         \mult_26/ab[19][26] , \mult_26/ab[19][27] , \mult_26/ab[19][28] ,
         \mult_26/ab[19][29] , \mult_26/ab[19][30] , \mult_26/ab[19][31] ,
         \mult_26/ab[20][0] , \mult_26/ab[20][1] , \mult_26/ab[20][2] ,
         \mult_26/ab[20][3] , \mult_26/ab[20][4] , \mult_26/ab[20][5] ,
         \mult_26/ab[20][6] , \mult_26/ab[20][7] , \mult_26/ab[20][8] ,
         \mult_26/ab[20][9] , \mult_26/ab[20][10] , \mult_26/ab[20][11] ,
         \mult_26/ab[20][12] , \mult_26/ab[20][13] , \mult_26/ab[20][14] ,
         \mult_26/ab[20][15] , \mult_26/ab[20][16] , \mult_26/ab[20][17] ,
         \mult_26/ab[20][18] , \mult_26/ab[20][19] , \mult_26/ab[20][20] ,
         \mult_26/ab[20][21] , \mult_26/ab[20][22] , \mult_26/ab[20][23] ,
         \mult_26/ab[20][24] , \mult_26/ab[20][25] , \mult_26/ab[20][26] ,
         \mult_26/ab[20][27] , \mult_26/ab[20][28] , \mult_26/ab[20][29] ,
         \mult_26/ab[20][30] , \mult_26/ab[20][31] , \mult_26/ab[21][0] ,
         \mult_26/ab[21][1] , \mult_26/ab[21][2] , \mult_26/ab[21][3] ,
         \mult_26/ab[21][4] , \mult_26/ab[21][5] , \mult_26/ab[21][6] ,
         \mult_26/ab[21][7] , \mult_26/ab[21][8] , \mult_26/ab[21][9] ,
         \mult_26/ab[21][10] , \mult_26/ab[21][11] , \mult_26/ab[21][12] ,
         \mult_26/ab[21][13] , \mult_26/ab[21][14] , \mult_26/ab[21][15] ,
         \mult_26/ab[21][16] , \mult_26/ab[21][17] , \mult_26/ab[21][18] ,
         \mult_26/ab[21][19] , \mult_26/ab[21][20] , \mult_26/ab[21][21] ,
         \mult_26/ab[21][22] , \mult_26/ab[21][23] , \mult_26/ab[21][24] ,
         \mult_26/ab[21][25] , \mult_26/ab[21][26] , \mult_26/ab[21][27] ,
         \mult_26/ab[21][28] , \mult_26/ab[21][29] , \mult_26/ab[21][30] ,
         \mult_26/ab[21][31] , \mult_26/ab[22][0] , \mult_26/ab[22][1] ,
         \mult_26/ab[22][2] , \mult_26/ab[22][3] , \mult_26/ab[22][4] ,
         \mult_26/ab[22][5] , \mult_26/ab[22][6] , \mult_26/ab[22][7] ,
         \mult_26/ab[22][8] , \mult_26/ab[22][9] , \mult_26/ab[22][10] ,
         \mult_26/ab[22][11] , \mult_26/ab[22][12] , \mult_26/ab[22][13] ,
         \mult_26/ab[22][14] , \mult_26/ab[22][15] , \mult_26/ab[22][16] ,
         \mult_26/ab[22][17] , \mult_26/ab[22][18] , \mult_26/ab[22][19] ,
         \mult_26/ab[22][20] , \mult_26/ab[22][21] , \mult_26/ab[22][22] ,
         \mult_26/ab[22][23] , \mult_26/ab[22][24] , \mult_26/ab[22][25] ,
         \mult_26/ab[22][26] , \mult_26/ab[22][27] , \mult_26/ab[22][28] ,
         \mult_26/ab[22][29] , \mult_26/ab[22][30] , \mult_26/ab[22][31] ,
         \mult_26/ab[23][0] , \mult_26/ab[23][1] , \mult_26/ab[23][2] ,
         \mult_26/ab[23][3] , \mult_26/ab[23][4] , \mult_26/ab[23][5] ,
         \mult_26/ab[23][6] , \mult_26/ab[23][7] , \mult_26/ab[23][8] ,
         \mult_26/ab[23][9] , \mult_26/ab[23][10] , \mult_26/ab[23][11] ,
         \mult_26/ab[23][12] , \mult_26/ab[23][13] , \mult_26/ab[23][14] ,
         \mult_26/ab[23][15] , \mult_26/ab[23][16] , \mult_26/ab[23][17] ,
         \mult_26/ab[23][18] , \mult_26/ab[23][19] , \mult_26/ab[23][20] ,
         \mult_26/ab[23][21] , \mult_26/ab[23][22] , \mult_26/ab[23][23] ,
         \mult_26/ab[23][24] , \mult_26/ab[23][25] , \mult_26/ab[23][26] ,
         \mult_26/ab[23][27] , \mult_26/ab[23][28] , \mult_26/ab[23][29] ,
         \mult_26/ab[23][30] , \mult_26/ab[23][31] , \mult_26/ab[24][0] ,
         \mult_26/ab[24][1] , \mult_26/ab[24][2] , \mult_26/ab[24][3] ,
         \mult_26/ab[24][4] , \mult_26/ab[24][5] , \mult_26/ab[24][6] ,
         \mult_26/ab[24][7] , \mult_26/ab[24][8] , \mult_26/ab[24][9] ,
         \mult_26/ab[24][10] , \mult_26/ab[24][11] , \mult_26/ab[24][12] ,
         \mult_26/ab[24][13] , \mult_26/ab[24][14] , \mult_26/ab[24][15] ,
         \mult_26/ab[24][16] , \mult_26/ab[24][17] , \mult_26/ab[24][18] ,
         \mult_26/ab[24][19] , \mult_26/ab[24][20] , \mult_26/ab[24][21] ,
         \mult_26/ab[24][22] , \mult_26/ab[24][23] , \mult_26/ab[24][24] ,
         \mult_26/ab[24][25] , \mult_26/ab[24][26] , \mult_26/ab[24][27] ,
         \mult_26/ab[24][28] , \mult_26/ab[24][29] , \mult_26/ab[24][30] ,
         \mult_26/ab[24][31] , \mult_26/ab[25][0] , \mult_26/ab[25][1] ,
         \mult_26/ab[25][2] , \mult_26/ab[25][3] , \mult_26/ab[25][4] ,
         \mult_26/ab[25][5] , \mult_26/ab[25][6] , \mult_26/ab[25][7] ,
         \mult_26/ab[25][8] , \mult_26/ab[25][9] , \mult_26/ab[25][10] ,
         \mult_26/ab[25][11] , \mult_26/ab[25][12] , \mult_26/ab[25][13] ,
         \mult_26/ab[25][14] , \mult_26/ab[25][15] , \mult_26/ab[25][16] ,
         \mult_26/ab[25][17] , \mult_26/ab[25][18] , \mult_26/ab[25][19] ,
         \mult_26/ab[25][20] , \mult_26/ab[25][21] , \mult_26/ab[25][22] ,
         \mult_26/ab[25][23] , \mult_26/ab[25][24] , \mult_26/ab[25][25] ,
         \mult_26/ab[25][26] , \mult_26/ab[25][27] , \mult_26/ab[25][28] ,
         \mult_26/ab[25][29] , \mult_26/ab[25][30] , \mult_26/ab[25][31] ,
         \mult_26/ab[26][0] , \mult_26/ab[26][1] , \mult_26/ab[26][2] ,
         \mult_26/ab[26][3] , \mult_26/ab[26][4] , \mult_26/ab[26][5] ,
         \mult_26/ab[26][6] , \mult_26/ab[26][7] , \mult_26/ab[26][8] ,
         \mult_26/ab[26][9] , \mult_26/ab[26][10] , \mult_26/ab[26][11] ,
         \mult_26/ab[26][12] , \mult_26/ab[26][13] , \mult_26/ab[26][14] ,
         \mult_26/ab[26][15] , \mult_26/ab[26][16] , \mult_26/ab[26][17] ,
         \mult_26/ab[26][18] , \mult_26/ab[26][19] , \mult_26/ab[26][20] ,
         \mult_26/ab[26][21] , \mult_26/ab[26][22] , \mult_26/ab[26][23] ,
         \mult_26/ab[26][24] , \mult_26/ab[26][25] , \mult_26/ab[26][26] ,
         \mult_26/ab[26][27] , \mult_26/ab[26][28] , \mult_26/ab[26][29] ,
         \mult_26/ab[26][30] , \mult_26/ab[26][31] , \mult_26/ab[27][0] ,
         \mult_26/ab[27][1] , \mult_26/ab[27][2] , \mult_26/ab[27][3] ,
         \mult_26/ab[27][4] , \mult_26/ab[27][5] , \mult_26/ab[27][6] ,
         \mult_26/ab[27][7] , \mult_26/ab[27][8] , \mult_26/ab[27][9] ,
         \mult_26/ab[27][10] , \mult_26/ab[27][11] , \mult_26/ab[27][12] ,
         \mult_26/ab[27][13] , \mult_26/ab[27][14] , \mult_26/ab[27][15] ,
         \mult_26/ab[27][16] , \mult_26/ab[27][17] , \mult_26/ab[27][18] ,
         \mult_26/ab[27][19] , \mult_26/ab[27][20] , \mult_26/ab[27][21] ,
         \mult_26/ab[27][22] , \mult_26/ab[27][23] , \mult_26/ab[27][24] ,
         \mult_26/ab[27][25] , \mult_26/ab[27][26] , \mult_26/ab[27][27] ,
         \mult_26/ab[27][28] , \mult_26/ab[27][29] , \mult_26/ab[27][30] ,
         \mult_26/ab[27][31] , \mult_26/ab[28][0] , \mult_26/ab[28][1] ,
         \mult_26/ab[28][2] , \mult_26/ab[28][3] , \mult_26/ab[28][4] ,
         \mult_26/ab[28][5] , \mult_26/ab[28][6] , \mult_26/ab[28][7] ,
         \mult_26/ab[28][8] , \mult_26/ab[28][9] , \mult_26/ab[28][10] ,
         \mult_26/ab[28][11] , \mult_26/ab[28][12] , \mult_26/ab[28][13] ,
         \mult_26/ab[28][14] , \mult_26/ab[28][15] , \mult_26/ab[28][16] ,
         \mult_26/ab[28][17] , \mult_26/ab[28][18] , \mult_26/ab[28][19] ,
         \mult_26/ab[28][20] , \mult_26/ab[28][21] , \mult_26/ab[28][22] ,
         \mult_26/ab[28][23] , \mult_26/ab[28][24] , \mult_26/ab[28][25] ,
         \mult_26/ab[28][26] , \mult_26/ab[28][27] , \mult_26/ab[28][28] ,
         \mult_26/ab[28][29] , \mult_26/ab[28][30] , \mult_26/ab[28][31] ,
         \mult_26/ab[29][0] , \mult_26/ab[29][1] , \mult_26/ab[29][2] ,
         \mult_26/ab[29][3] , \mult_26/ab[29][4] , \mult_26/ab[29][5] ,
         \mult_26/ab[29][6] , \mult_26/ab[29][7] , \mult_26/ab[29][8] ,
         \mult_26/ab[29][9] , \mult_26/ab[29][10] , \mult_26/ab[29][11] ,
         \mult_26/ab[29][12] , \mult_26/ab[29][13] , \mult_26/ab[29][14] ,
         \mult_26/ab[29][15] , \mult_26/ab[29][16] , \mult_26/ab[29][17] ,
         \mult_26/ab[29][18] , \mult_26/ab[29][19] , \mult_26/ab[29][20] ,
         \mult_26/ab[29][21] , \mult_26/ab[29][22] , \mult_26/ab[29][23] ,
         \mult_26/ab[29][24] , \mult_26/ab[29][25] , \mult_26/ab[29][26] ,
         \mult_26/ab[29][27] , \mult_26/ab[29][28] , \mult_26/ab[29][29] ,
         \mult_26/ab[29][30] , \mult_26/ab[29][31] , \mult_26/ab[30][0] ,
         \mult_26/ab[30][1] , \mult_26/ab[30][2] , \mult_26/ab[30][3] ,
         \mult_26/ab[30][4] , \mult_26/ab[30][5] , \mult_26/ab[30][6] ,
         \mult_26/ab[30][7] , \mult_26/ab[30][8] , \mult_26/ab[30][9] ,
         \mult_26/ab[30][10] , \mult_26/ab[30][11] , \mult_26/ab[30][12] ,
         \mult_26/ab[30][13] , \mult_26/ab[30][14] , \mult_26/ab[30][15] ,
         \mult_26/ab[30][16] , \mult_26/ab[30][17] , \mult_26/ab[30][18] ,
         \mult_26/ab[30][19] , \mult_26/ab[30][20] , \mult_26/ab[30][21] ,
         \mult_26/ab[30][22] , \mult_26/ab[30][23] , \mult_26/ab[30][24] ,
         \mult_26/ab[30][25] , \mult_26/ab[30][26] , \mult_26/ab[30][27] ,
         \mult_26/ab[30][28] , \mult_26/ab[30][29] , \mult_26/ab[30][30] ,
         \mult_26/ab[30][31] , \mult_26/ab[31][0] , \mult_26/ab[31][1] ,
         \mult_26/ab[31][2] , \mult_26/ab[31][3] , \mult_26/ab[31][4] ,
         \mult_26/ab[31][5] , \mult_26/ab[31][6] , \mult_26/ab[31][7] ,
         \mult_26/ab[31][8] , \mult_26/ab[31][9] , \mult_26/ab[31][10] ,
         \mult_26/ab[31][11] , \mult_26/ab[31][12] , \mult_26/ab[31][13] ,
         \mult_26/ab[31][14] , \mult_26/ab[31][15] , \mult_26/ab[31][16] ,
         \mult_26/ab[31][17] , \mult_26/ab[31][18] , \mult_26/ab[31][19] ,
         \mult_26/ab[31][20] , \mult_26/ab[31][21] , \mult_26/ab[31][22] ,
         \mult_26/ab[31][23] , \mult_26/ab[31][24] , \mult_26/ab[31][25] ,
         \mult_26/ab[31][26] , \mult_26/ab[31][27] , \mult_26/ab[31][28] ,
         \mult_26/ab[31][29] , \mult_26/ab[31][30] , \mult_26/ab[31][31] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186;
  assign o[31] = \mult_26/SUMB[31][0] ;

  FADDER \mult_26/S3_2_30  ( .CIN(\mult_26/ab[2][30] ), .IN0(
        \mult_26/CARRYB[1][30] ), .IN1(\mult_26/ab[1][31] ), .COUT(
        \mult_26/CARRYB[2][30] ), .SUM(\mult_26/SUMB[2][30] ) );
  FADDER \mult_26/S2_2_29  ( .CIN(\mult_26/ab[2][29] ), .IN0(
        \mult_26/CARRYB[1][29] ), .IN1(\mult_26/SUMB[1][30] ), .COUT(
        \mult_26/CARRYB[2][29] ), .SUM(\mult_26/SUMB[2][29] ) );
  FADDER \mult_26/S2_2_28  ( .CIN(\mult_26/ab[2][28] ), .IN0(
        \mult_26/CARRYB[1][28] ), .IN1(\mult_26/SUMB[1][29] ), .COUT(
        \mult_26/CARRYB[2][28] ), .SUM(\mult_26/SUMB[2][28] ) );
  FADDER \mult_26/S2_2_27  ( .CIN(\mult_26/ab[2][27] ), .IN0(
        \mult_26/CARRYB[1][27] ), .IN1(\mult_26/SUMB[1][28] ), .COUT(
        \mult_26/CARRYB[2][27] ), .SUM(\mult_26/SUMB[2][27] ) );
  FADDER \mult_26/S2_2_26  ( .CIN(\mult_26/ab[2][26] ), .IN0(
        \mult_26/CARRYB[1][26] ), .IN1(\mult_26/SUMB[1][27] ), .COUT(
        \mult_26/CARRYB[2][26] ), .SUM(\mult_26/SUMB[2][26] ) );
  FADDER \mult_26/S2_2_25  ( .CIN(\mult_26/ab[2][25] ), .IN0(
        \mult_26/CARRYB[1][25] ), .IN1(\mult_26/SUMB[1][26] ), .COUT(
        \mult_26/CARRYB[2][25] ), .SUM(\mult_26/SUMB[2][25] ) );
  FADDER \mult_26/S2_2_24  ( .CIN(\mult_26/ab[2][24] ), .IN0(
        \mult_26/CARRYB[1][24] ), .IN1(\mult_26/SUMB[1][25] ), .COUT(
        \mult_26/CARRYB[2][24] ), .SUM(\mult_26/SUMB[2][24] ) );
  FADDER \mult_26/S2_2_23  ( .CIN(\mult_26/ab[2][23] ), .IN0(
        \mult_26/CARRYB[1][23] ), .IN1(\mult_26/SUMB[1][24] ), .COUT(
        \mult_26/CARRYB[2][23] ), .SUM(\mult_26/SUMB[2][23] ) );
  FADDER \mult_26/S2_2_22  ( .CIN(\mult_26/ab[2][22] ), .IN0(
        \mult_26/CARRYB[1][22] ), .IN1(\mult_26/SUMB[1][23] ), .COUT(
        \mult_26/CARRYB[2][22] ), .SUM(\mult_26/SUMB[2][22] ) );
  FADDER \mult_26/S2_2_21  ( .CIN(\mult_26/ab[2][21] ), .IN0(
        \mult_26/CARRYB[1][21] ), .IN1(\mult_26/SUMB[1][22] ), .COUT(
        \mult_26/CARRYB[2][21] ), .SUM(\mult_26/SUMB[2][21] ) );
  FADDER \mult_26/S2_2_20  ( .CIN(\mult_26/ab[2][20] ), .IN0(
        \mult_26/CARRYB[1][20] ), .IN1(\mult_26/SUMB[1][21] ), .COUT(
        \mult_26/CARRYB[2][20] ), .SUM(\mult_26/SUMB[2][20] ) );
  FADDER \mult_26/S2_2_19  ( .CIN(\mult_26/ab[2][19] ), .IN0(
        \mult_26/CARRYB[1][19] ), .IN1(\mult_26/SUMB[1][20] ), .COUT(
        \mult_26/CARRYB[2][19] ), .SUM(\mult_26/SUMB[2][19] ) );
  FADDER \mult_26/S2_2_18  ( .CIN(\mult_26/ab[2][18] ), .IN0(
        \mult_26/CARRYB[1][18] ), .IN1(\mult_26/SUMB[1][19] ), .COUT(
        \mult_26/CARRYB[2][18] ), .SUM(\mult_26/SUMB[2][18] ) );
  FADDER \mult_26/S2_2_17  ( .CIN(\mult_26/ab[2][17] ), .IN0(
        \mult_26/CARRYB[1][17] ), .IN1(\mult_26/SUMB[1][18] ), .COUT(
        \mult_26/CARRYB[2][17] ), .SUM(\mult_26/SUMB[2][17] ) );
  FADDER \mult_26/S2_2_16  ( .CIN(\mult_26/ab[2][16] ), .IN0(
        \mult_26/CARRYB[1][16] ), .IN1(\mult_26/SUMB[1][17] ), .COUT(
        \mult_26/CARRYB[2][16] ), .SUM(\mult_26/SUMB[2][16] ) );
  FADDER \mult_26/S2_2_15  ( .CIN(\mult_26/ab[2][15] ), .IN0(
        \mult_26/CARRYB[1][15] ), .IN1(\mult_26/SUMB[1][16] ), .COUT(
        \mult_26/CARRYB[2][15] ), .SUM(\mult_26/SUMB[2][15] ) );
  FADDER \mult_26/S2_2_14  ( .CIN(\mult_26/ab[2][14] ), .IN0(
        \mult_26/CARRYB[1][14] ), .IN1(\mult_26/SUMB[1][15] ), .COUT(
        \mult_26/CARRYB[2][14] ), .SUM(\mult_26/SUMB[2][14] ) );
  FADDER \mult_26/S2_2_13  ( .CIN(\mult_26/ab[2][13] ), .IN0(
        \mult_26/CARRYB[1][13] ), .IN1(\mult_26/SUMB[1][14] ), .COUT(
        \mult_26/CARRYB[2][13] ), .SUM(\mult_26/SUMB[2][13] ) );
  FADDER \mult_26/S2_2_12  ( .CIN(\mult_26/ab[2][12] ), .IN0(
        \mult_26/CARRYB[1][12] ), .IN1(\mult_26/SUMB[1][13] ), .COUT(
        \mult_26/CARRYB[2][12] ), .SUM(\mult_26/SUMB[2][12] ) );
  FADDER \mult_26/S2_2_11  ( .CIN(\mult_26/ab[2][11] ), .IN0(
        \mult_26/CARRYB[1][11] ), .IN1(\mult_26/SUMB[1][12] ), .COUT(
        \mult_26/CARRYB[2][11] ), .SUM(\mult_26/SUMB[2][11] ) );
  FADDER \mult_26/S2_2_10  ( .CIN(\mult_26/ab[2][10] ), .IN0(
        \mult_26/CARRYB[1][10] ), .IN1(\mult_26/SUMB[1][11] ), .COUT(
        \mult_26/CARRYB[2][10] ), .SUM(\mult_26/SUMB[2][10] ) );
  FADDER \mult_26/S2_2_9  ( .CIN(\mult_26/ab[2][9] ), .IN0(
        \mult_26/CARRYB[1][9] ), .IN1(\mult_26/SUMB[1][10] ), .COUT(
        \mult_26/CARRYB[2][9] ), .SUM(\mult_26/SUMB[2][9] ) );
  FADDER \mult_26/S2_2_8  ( .CIN(\mult_26/ab[2][8] ), .IN0(
        \mult_26/CARRYB[1][8] ), .IN1(\mult_26/SUMB[1][9] ), .COUT(
        \mult_26/CARRYB[2][8] ), .SUM(\mult_26/SUMB[2][8] ) );
  FADDER \mult_26/S2_2_7  ( .CIN(\mult_26/ab[2][7] ), .IN0(
        \mult_26/CARRYB[1][7] ), .IN1(\mult_26/SUMB[1][8] ), .COUT(
        \mult_26/CARRYB[2][7] ), .SUM(\mult_26/SUMB[2][7] ) );
  FADDER \mult_26/S2_2_6  ( .CIN(\mult_26/ab[2][6] ), .IN0(
        \mult_26/CARRYB[1][6] ), .IN1(\mult_26/SUMB[1][7] ), .COUT(
        \mult_26/CARRYB[2][6] ), .SUM(\mult_26/SUMB[2][6] ) );
  FADDER \mult_26/S2_2_5  ( .CIN(\mult_26/ab[2][5] ), .IN0(
        \mult_26/CARRYB[1][5] ), .IN1(\mult_26/SUMB[1][6] ), .COUT(
        \mult_26/CARRYB[2][5] ), .SUM(\mult_26/SUMB[2][5] ) );
  FADDER \mult_26/S2_2_4  ( .CIN(\mult_26/ab[2][4] ), .IN0(
        \mult_26/CARRYB[1][4] ), .IN1(\mult_26/SUMB[1][5] ), .COUT(
        \mult_26/CARRYB[2][4] ), .SUM(\mult_26/SUMB[2][4] ) );
  FADDER \mult_26/S2_2_3  ( .CIN(\mult_26/ab[2][3] ), .IN0(
        \mult_26/CARRYB[1][3] ), .IN1(\mult_26/SUMB[1][4] ), .COUT(
        \mult_26/CARRYB[2][3] ), .SUM(\mult_26/SUMB[2][3] ) );
  FADDER \mult_26/S2_2_2  ( .CIN(\mult_26/ab[2][2] ), .IN0(
        \mult_26/CARRYB[1][2] ), .IN1(\mult_26/SUMB[1][3] ), .COUT(
        \mult_26/CARRYB[2][2] ), .SUM(\mult_26/SUMB[2][2] ) );
  FADDER \mult_26/S2_2_1  ( .CIN(\mult_26/ab[2][1] ), .IN0(
        \mult_26/CARRYB[1][1] ), .IN1(\mult_26/SUMB[1][2] ), .COUT(
        \mult_26/CARRYB[2][1] ), .SUM(\mult_26/SUMB[2][1] ) );
  FADDER \mult_26/S1_2_0  ( .CIN(\mult_26/ab[2][0] ), .IN0(
        \mult_26/CARRYB[1][0] ), .IN1(\mult_26/SUMB[1][1] ), .COUT(
        \mult_26/CARRYB[2][0] ), .SUM(o[2]) );
  FADDER \mult_26/S3_3_30  ( .CIN(\mult_26/ab[3][30] ), .IN0(
        \mult_26/CARRYB[2][30] ), .IN1(\mult_26/ab[2][31] ), .COUT(
        \mult_26/CARRYB[3][30] ), .SUM(\mult_26/SUMB[3][30] ) );
  FADDER \mult_26/S2_3_29  ( .CIN(\mult_26/ab[3][29] ), .IN0(
        \mult_26/CARRYB[2][29] ), .IN1(\mult_26/SUMB[2][30] ), .COUT(
        \mult_26/CARRYB[3][29] ), .SUM(\mult_26/SUMB[3][29] ) );
  FADDER \mult_26/S2_3_28  ( .CIN(\mult_26/ab[3][28] ), .IN0(
        \mult_26/CARRYB[2][28] ), .IN1(\mult_26/SUMB[2][29] ), .COUT(
        \mult_26/CARRYB[3][28] ), .SUM(\mult_26/SUMB[3][28] ) );
  FADDER \mult_26/S2_3_27  ( .CIN(\mult_26/ab[3][27] ), .IN0(
        \mult_26/CARRYB[2][27] ), .IN1(\mult_26/SUMB[2][28] ), .COUT(
        \mult_26/CARRYB[3][27] ), .SUM(\mult_26/SUMB[3][27] ) );
  FADDER \mult_26/S2_3_26  ( .CIN(\mult_26/ab[3][26] ), .IN0(
        \mult_26/CARRYB[2][26] ), .IN1(\mult_26/SUMB[2][27] ), .COUT(
        \mult_26/CARRYB[3][26] ), .SUM(\mult_26/SUMB[3][26] ) );
  FADDER \mult_26/S2_3_25  ( .CIN(\mult_26/ab[3][25] ), .IN0(
        \mult_26/CARRYB[2][25] ), .IN1(\mult_26/SUMB[2][26] ), .COUT(
        \mult_26/CARRYB[3][25] ), .SUM(\mult_26/SUMB[3][25] ) );
  FADDER \mult_26/S2_3_24  ( .CIN(\mult_26/ab[3][24] ), .IN0(
        \mult_26/CARRYB[2][24] ), .IN1(\mult_26/SUMB[2][25] ), .COUT(
        \mult_26/CARRYB[3][24] ), .SUM(\mult_26/SUMB[3][24] ) );
  FADDER \mult_26/S2_3_23  ( .CIN(\mult_26/ab[3][23] ), .IN0(
        \mult_26/CARRYB[2][23] ), .IN1(\mult_26/SUMB[2][24] ), .COUT(
        \mult_26/CARRYB[3][23] ), .SUM(\mult_26/SUMB[3][23] ) );
  FADDER \mult_26/S2_3_22  ( .CIN(\mult_26/ab[3][22] ), .IN0(
        \mult_26/CARRYB[2][22] ), .IN1(\mult_26/SUMB[2][23] ), .COUT(
        \mult_26/CARRYB[3][22] ), .SUM(\mult_26/SUMB[3][22] ) );
  FADDER \mult_26/S2_3_21  ( .CIN(\mult_26/ab[3][21] ), .IN0(
        \mult_26/CARRYB[2][21] ), .IN1(\mult_26/SUMB[2][22] ), .COUT(
        \mult_26/CARRYB[3][21] ), .SUM(\mult_26/SUMB[3][21] ) );
  FADDER \mult_26/S2_3_20  ( .CIN(\mult_26/ab[3][20] ), .IN0(
        \mult_26/CARRYB[2][20] ), .IN1(\mult_26/SUMB[2][21] ), .COUT(
        \mult_26/CARRYB[3][20] ), .SUM(\mult_26/SUMB[3][20] ) );
  FADDER \mult_26/S2_3_19  ( .CIN(\mult_26/ab[3][19] ), .IN0(
        \mult_26/CARRYB[2][19] ), .IN1(\mult_26/SUMB[2][20] ), .COUT(
        \mult_26/CARRYB[3][19] ), .SUM(\mult_26/SUMB[3][19] ) );
  FADDER \mult_26/S2_3_18  ( .CIN(\mult_26/ab[3][18] ), .IN0(
        \mult_26/CARRYB[2][18] ), .IN1(\mult_26/SUMB[2][19] ), .COUT(
        \mult_26/CARRYB[3][18] ), .SUM(\mult_26/SUMB[3][18] ) );
  FADDER \mult_26/S2_3_17  ( .CIN(\mult_26/ab[3][17] ), .IN0(
        \mult_26/CARRYB[2][17] ), .IN1(\mult_26/SUMB[2][18] ), .COUT(
        \mult_26/CARRYB[3][17] ), .SUM(\mult_26/SUMB[3][17] ) );
  FADDER \mult_26/S2_3_16  ( .CIN(\mult_26/ab[3][16] ), .IN0(
        \mult_26/CARRYB[2][16] ), .IN1(\mult_26/SUMB[2][17] ), .COUT(
        \mult_26/CARRYB[3][16] ), .SUM(\mult_26/SUMB[3][16] ) );
  FADDER \mult_26/S2_3_15  ( .CIN(\mult_26/ab[3][15] ), .IN0(
        \mult_26/CARRYB[2][15] ), .IN1(\mult_26/SUMB[2][16] ), .COUT(
        \mult_26/CARRYB[3][15] ), .SUM(\mult_26/SUMB[3][15] ) );
  FADDER \mult_26/S2_3_14  ( .CIN(\mult_26/ab[3][14] ), .IN0(
        \mult_26/CARRYB[2][14] ), .IN1(\mult_26/SUMB[2][15] ), .COUT(
        \mult_26/CARRYB[3][14] ), .SUM(\mult_26/SUMB[3][14] ) );
  FADDER \mult_26/S2_3_13  ( .CIN(\mult_26/ab[3][13] ), .IN0(
        \mult_26/CARRYB[2][13] ), .IN1(\mult_26/SUMB[2][14] ), .COUT(
        \mult_26/CARRYB[3][13] ), .SUM(\mult_26/SUMB[3][13] ) );
  FADDER \mult_26/S2_3_12  ( .CIN(\mult_26/ab[3][12] ), .IN0(
        \mult_26/CARRYB[2][12] ), .IN1(\mult_26/SUMB[2][13] ), .COUT(
        \mult_26/CARRYB[3][12] ), .SUM(\mult_26/SUMB[3][12] ) );
  FADDER \mult_26/S2_3_11  ( .CIN(\mult_26/ab[3][11] ), .IN0(
        \mult_26/CARRYB[2][11] ), .IN1(\mult_26/SUMB[2][12] ), .COUT(
        \mult_26/CARRYB[3][11] ), .SUM(\mult_26/SUMB[3][11] ) );
  FADDER \mult_26/S2_3_10  ( .CIN(\mult_26/ab[3][10] ), .IN0(
        \mult_26/CARRYB[2][10] ), .IN1(\mult_26/SUMB[2][11] ), .COUT(
        \mult_26/CARRYB[3][10] ), .SUM(\mult_26/SUMB[3][10] ) );
  FADDER \mult_26/S2_3_9  ( .CIN(\mult_26/ab[3][9] ), .IN0(
        \mult_26/CARRYB[2][9] ), .IN1(\mult_26/SUMB[2][10] ), .COUT(
        \mult_26/CARRYB[3][9] ), .SUM(\mult_26/SUMB[3][9] ) );
  FADDER \mult_26/S2_3_8  ( .CIN(\mult_26/ab[3][8] ), .IN0(
        \mult_26/CARRYB[2][8] ), .IN1(\mult_26/SUMB[2][9] ), .COUT(
        \mult_26/CARRYB[3][8] ), .SUM(\mult_26/SUMB[3][8] ) );
  FADDER \mult_26/S2_3_7  ( .CIN(\mult_26/ab[3][7] ), .IN0(
        \mult_26/CARRYB[2][7] ), .IN1(\mult_26/SUMB[2][8] ), .COUT(
        \mult_26/CARRYB[3][7] ), .SUM(\mult_26/SUMB[3][7] ) );
  FADDER \mult_26/S2_3_6  ( .CIN(\mult_26/ab[3][6] ), .IN0(
        \mult_26/CARRYB[2][6] ), .IN1(\mult_26/SUMB[2][7] ), .COUT(
        \mult_26/CARRYB[3][6] ), .SUM(\mult_26/SUMB[3][6] ) );
  FADDER \mult_26/S2_3_5  ( .CIN(\mult_26/ab[3][5] ), .IN0(
        \mult_26/CARRYB[2][5] ), .IN1(\mult_26/SUMB[2][6] ), .COUT(
        \mult_26/CARRYB[3][5] ), .SUM(\mult_26/SUMB[3][5] ) );
  FADDER \mult_26/S2_3_4  ( .CIN(\mult_26/ab[3][4] ), .IN0(
        \mult_26/CARRYB[2][4] ), .IN1(\mult_26/SUMB[2][5] ), .COUT(
        \mult_26/CARRYB[3][4] ), .SUM(\mult_26/SUMB[3][4] ) );
  FADDER \mult_26/S2_3_3  ( .CIN(\mult_26/ab[3][3] ), .IN0(
        \mult_26/CARRYB[2][3] ), .IN1(\mult_26/SUMB[2][4] ), .COUT(
        \mult_26/CARRYB[3][3] ), .SUM(\mult_26/SUMB[3][3] ) );
  FADDER \mult_26/S2_3_2  ( .CIN(\mult_26/ab[3][2] ), .IN0(
        \mult_26/CARRYB[2][2] ), .IN1(\mult_26/SUMB[2][3] ), .COUT(
        \mult_26/CARRYB[3][2] ), .SUM(\mult_26/SUMB[3][2] ) );
  FADDER \mult_26/S2_3_1  ( .CIN(\mult_26/ab[3][1] ), .IN0(
        \mult_26/CARRYB[2][1] ), .IN1(\mult_26/SUMB[2][2] ), .COUT(
        \mult_26/CARRYB[3][1] ), .SUM(\mult_26/SUMB[3][1] ) );
  FADDER \mult_26/S1_3_0  ( .CIN(\mult_26/ab[3][0] ), .IN0(
        \mult_26/CARRYB[2][0] ), .IN1(\mult_26/SUMB[2][1] ), .COUT(
        \mult_26/CARRYB[3][0] ), .SUM(o[3]) );
  FADDER \mult_26/S3_4_30  ( .CIN(\mult_26/ab[4][30] ), .IN0(
        \mult_26/CARRYB[3][30] ), .IN1(\mult_26/ab[3][31] ), .COUT(
        \mult_26/CARRYB[4][30] ), .SUM(\mult_26/SUMB[4][30] ) );
  FADDER \mult_26/S2_4_29  ( .CIN(\mult_26/ab[4][29] ), .IN0(
        \mult_26/CARRYB[3][29] ), .IN1(\mult_26/SUMB[3][30] ), .COUT(
        \mult_26/CARRYB[4][29] ), .SUM(\mult_26/SUMB[4][29] ) );
  FADDER \mult_26/S2_4_28  ( .CIN(\mult_26/ab[4][28] ), .IN0(
        \mult_26/CARRYB[3][28] ), .IN1(\mult_26/SUMB[3][29] ), .COUT(
        \mult_26/CARRYB[4][28] ), .SUM(\mult_26/SUMB[4][28] ) );
  FADDER \mult_26/S2_4_27  ( .CIN(\mult_26/ab[4][27] ), .IN0(
        \mult_26/CARRYB[3][27] ), .IN1(\mult_26/SUMB[3][28] ), .COUT(
        \mult_26/CARRYB[4][27] ), .SUM(\mult_26/SUMB[4][27] ) );
  FADDER \mult_26/S2_4_26  ( .CIN(\mult_26/ab[4][26] ), .IN0(
        \mult_26/CARRYB[3][26] ), .IN1(\mult_26/SUMB[3][27] ), .COUT(
        \mult_26/CARRYB[4][26] ), .SUM(\mult_26/SUMB[4][26] ) );
  FADDER \mult_26/S2_4_25  ( .CIN(\mult_26/ab[4][25] ), .IN0(
        \mult_26/CARRYB[3][25] ), .IN1(\mult_26/SUMB[3][26] ), .COUT(
        \mult_26/CARRYB[4][25] ), .SUM(\mult_26/SUMB[4][25] ) );
  FADDER \mult_26/S2_4_24  ( .CIN(\mult_26/ab[4][24] ), .IN0(
        \mult_26/CARRYB[3][24] ), .IN1(\mult_26/SUMB[3][25] ), .COUT(
        \mult_26/CARRYB[4][24] ), .SUM(\mult_26/SUMB[4][24] ) );
  FADDER \mult_26/S2_4_23  ( .CIN(\mult_26/ab[4][23] ), .IN0(
        \mult_26/CARRYB[3][23] ), .IN1(\mult_26/SUMB[3][24] ), .COUT(
        \mult_26/CARRYB[4][23] ), .SUM(\mult_26/SUMB[4][23] ) );
  FADDER \mult_26/S2_4_22  ( .CIN(\mult_26/ab[4][22] ), .IN0(
        \mult_26/CARRYB[3][22] ), .IN1(\mult_26/SUMB[3][23] ), .COUT(
        \mult_26/CARRYB[4][22] ), .SUM(\mult_26/SUMB[4][22] ) );
  FADDER \mult_26/S2_4_21  ( .CIN(\mult_26/ab[4][21] ), .IN0(
        \mult_26/CARRYB[3][21] ), .IN1(\mult_26/SUMB[3][22] ), .COUT(
        \mult_26/CARRYB[4][21] ), .SUM(\mult_26/SUMB[4][21] ) );
  FADDER \mult_26/S2_4_20  ( .CIN(\mult_26/ab[4][20] ), .IN0(
        \mult_26/CARRYB[3][20] ), .IN1(\mult_26/SUMB[3][21] ), .COUT(
        \mult_26/CARRYB[4][20] ), .SUM(\mult_26/SUMB[4][20] ) );
  FADDER \mult_26/S2_4_19  ( .CIN(\mult_26/ab[4][19] ), .IN0(
        \mult_26/CARRYB[3][19] ), .IN1(\mult_26/SUMB[3][20] ), .COUT(
        \mult_26/CARRYB[4][19] ), .SUM(\mult_26/SUMB[4][19] ) );
  FADDER \mult_26/S2_4_18  ( .CIN(\mult_26/ab[4][18] ), .IN0(
        \mult_26/CARRYB[3][18] ), .IN1(\mult_26/SUMB[3][19] ), .COUT(
        \mult_26/CARRYB[4][18] ), .SUM(\mult_26/SUMB[4][18] ) );
  FADDER \mult_26/S2_4_17  ( .CIN(\mult_26/ab[4][17] ), .IN0(
        \mult_26/CARRYB[3][17] ), .IN1(\mult_26/SUMB[3][18] ), .COUT(
        \mult_26/CARRYB[4][17] ), .SUM(\mult_26/SUMB[4][17] ) );
  FADDER \mult_26/S2_4_16  ( .CIN(\mult_26/ab[4][16] ), .IN0(
        \mult_26/CARRYB[3][16] ), .IN1(\mult_26/SUMB[3][17] ), .COUT(
        \mult_26/CARRYB[4][16] ), .SUM(\mult_26/SUMB[4][16] ) );
  FADDER \mult_26/S2_4_15  ( .CIN(\mult_26/ab[4][15] ), .IN0(
        \mult_26/CARRYB[3][15] ), .IN1(\mult_26/SUMB[3][16] ), .COUT(
        \mult_26/CARRYB[4][15] ), .SUM(\mult_26/SUMB[4][15] ) );
  FADDER \mult_26/S2_4_14  ( .CIN(\mult_26/ab[4][14] ), .IN0(
        \mult_26/CARRYB[3][14] ), .IN1(\mult_26/SUMB[3][15] ), .COUT(
        \mult_26/CARRYB[4][14] ), .SUM(\mult_26/SUMB[4][14] ) );
  FADDER \mult_26/S2_4_13  ( .CIN(\mult_26/ab[4][13] ), .IN0(
        \mult_26/CARRYB[3][13] ), .IN1(\mult_26/SUMB[3][14] ), .COUT(
        \mult_26/CARRYB[4][13] ), .SUM(\mult_26/SUMB[4][13] ) );
  FADDER \mult_26/S2_4_12  ( .CIN(\mult_26/ab[4][12] ), .IN0(
        \mult_26/CARRYB[3][12] ), .IN1(\mult_26/SUMB[3][13] ), .COUT(
        \mult_26/CARRYB[4][12] ), .SUM(\mult_26/SUMB[4][12] ) );
  FADDER \mult_26/S2_4_11  ( .CIN(\mult_26/ab[4][11] ), .IN0(
        \mult_26/CARRYB[3][11] ), .IN1(\mult_26/SUMB[3][12] ), .COUT(
        \mult_26/CARRYB[4][11] ), .SUM(\mult_26/SUMB[4][11] ) );
  FADDER \mult_26/S2_4_10  ( .CIN(\mult_26/ab[4][10] ), .IN0(
        \mult_26/CARRYB[3][10] ), .IN1(\mult_26/SUMB[3][11] ), .COUT(
        \mult_26/CARRYB[4][10] ), .SUM(\mult_26/SUMB[4][10] ) );
  FADDER \mult_26/S2_4_9  ( .CIN(\mult_26/ab[4][9] ), .IN0(
        \mult_26/CARRYB[3][9] ), .IN1(\mult_26/SUMB[3][10] ), .COUT(
        \mult_26/CARRYB[4][9] ), .SUM(\mult_26/SUMB[4][9] ) );
  FADDER \mult_26/S2_4_8  ( .CIN(\mult_26/ab[4][8] ), .IN0(
        \mult_26/CARRYB[3][8] ), .IN1(\mult_26/SUMB[3][9] ), .COUT(
        \mult_26/CARRYB[4][8] ), .SUM(\mult_26/SUMB[4][8] ) );
  FADDER \mult_26/S2_4_7  ( .CIN(\mult_26/ab[4][7] ), .IN0(
        \mult_26/CARRYB[3][7] ), .IN1(\mult_26/SUMB[3][8] ), .COUT(
        \mult_26/CARRYB[4][7] ), .SUM(\mult_26/SUMB[4][7] ) );
  FADDER \mult_26/S2_4_6  ( .CIN(\mult_26/ab[4][6] ), .IN0(
        \mult_26/CARRYB[3][6] ), .IN1(\mult_26/SUMB[3][7] ), .COUT(
        \mult_26/CARRYB[4][6] ), .SUM(\mult_26/SUMB[4][6] ) );
  FADDER \mult_26/S2_4_5  ( .CIN(\mult_26/ab[4][5] ), .IN0(
        \mult_26/CARRYB[3][5] ), .IN1(\mult_26/SUMB[3][6] ), .COUT(
        \mult_26/CARRYB[4][5] ), .SUM(\mult_26/SUMB[4][5] ) );
  FADDER \mult_26/S2_4_4  ( .CIN(\mult_26/ab[4][4] ), .IN0(
        \mult_26/CARRYB[3][4] ), .IN1(\mult_26/SUMB[3][5] ), .COUT(
        \mult_26/CARRYB[4][4] ), .SUM(\mult_26/SUMB[4][4] ) );
  FADDER \mult_26/S2_4_3  ( .CIN(\mult_26/ab[4][3] ), .IN0(
        \mult_26/CARRYB[3][3] ), .IN1(\mult_26/SUMB[3][4] ), .COUT(
        \mult_26/CARRYB[4][3] ), .SUM(\mult_26/SUMB[4][3] ) );
  FADDER \mult_26/S2_4_2  ( .CIN(\mult_26/ab[4][2] ), .IN0(
        \mult_26/CARRYB[3][2] ), .IN1(\mult_26/SUMB[3][3] ), .COUT(
        \mult_26/CARRYB[4][2] ), .SUM(\mult_26/SUMB[4][2] ) );
  FADDER \mult_26/S2_4_1  ( .CIN(\mult_26/ab[4][1] ), .IN0(
        \mult_26/CARRYB[3][1] ), .IN1(\mult_26/SUMB[3][2] ), .COUT(
        \mult_26/CARRYB[4][1] ), .SUM(\mult_26/SUMB[4][1] ) );
  FADDER \mult_26/S1_4_0  ( .CIN(\mult_26/ab[4][0] ), .IN0(
        \mult_26/CARRYB[3][0] ), .IN1(\mult_26/SUMB[3][1] ), .COUT(
        \mult_26/CARRYB[4][0] ), .SUM(o[4]) );
  FADDER \mult_26/S3_5_30  ( .CIN(\mult_26/ab[5][30] ), .IN0(
        \mult_26/CARRYB[4][30] ), .IN1(\mult_26/ab[4][31] ), .COUT(
        \mult_26/CARRYB[5][30] ), .SUM(\mult_26/SUMB[5][30] ) );
  FADDER \mult_26/S2_5_29  ( .CIN(\mult_26/ab[5][29] ), .IN0(
        \mult_26/CARRYB[4][29] ), .IN1(\mult_26/SUMB[4][30] ), .COUT(
        \mult_26/CARRYB[5][29] ), .SUM(\mult_26/SUMB[5][29] ) );
  FADDER \mult_26/S2_5_28  ( .CIN(\mult_26/ab[5][28] ), .IN0(
        \mult_26/CARRYB[4][28] ), .IN1(\mult_26/SUMB[4][29] ), .COUT(
        \mult_26/CARRYB[5][28] ), .SUM(\mult_26/SUMB[5][28] ) );
  FADDER \mult_26/S2_5_27  ( .CIN(\mult_26/ab[5][27] ), .IN0(
        \mult_26/CARRYB[4][27] ), .IN1(\mult_26/SUMB[4][28] ), .COUT(
        \mult_26/CARRYB[5][27] ), .SUM(\mult_26/SUMB[5][27] ) );
  FADDER \mult_26/S2_5_26  ( .CIN(\mult_26/ab[5][26] ), .IN0(
        \mult_26/CARRYB[4][26] ), .IN1(\mult_26/SUMB[4][27] ), .COUT(
        \mult_26/CARRYB[5][26] ), .SUM(\mult_26/SUMB[5][26] ) );
  FADDER \mult_26/S2_5_25  ( .CIN(\mult_26/ab[5][25] ), .IN0(
        \mult_26/CARRYB[4][25] ), .IN1(\mult_26/SUMB[4][26] ), .COUT(
        \mult_26/CARRYB[5][25] ), .SUM(\mult_26/SUMB[5][25] ) );
  FADDER \mult_26/S2_5_24  ( .CIN(\mult_26/ab[5][24] ), .IN0(
        \mult_26/CARRYB[4][24] ), .IN1(\mult_26/SUMB[4][25] ), .COUT(
        \mult_26/CARRYB[5][24] ), .SUM(\mult_26/SUMB[5][24] ) );
  FADDER \mult_26/S2_5_23  ( .CIN(\mult_26/ab[5][23] ), .IN0(
        \mult_26/CARRYB[4][23] ), .IN1(\mult_26/SUMB[4][24] ), .COUT(
        \mult_26/CARRYB[5][23] ), .SUM(\mult_26/SUMB[5][23] ) );
  FADDER \mult_26/S2_5_22  ( .CIN(\mult_26/ab[5][22] ), .IN0(
        \mult_26/CARRYB[4][22] ), .IN1(\mult_26/SUMB[4][23] ), .COUT(
        \mult_26/CARRYB[5][22] ), .SUM(\mult_26/SUMB[5][22] ) );
  FADDER \mult_26/S2_5_21  ( .CIN(\mult_26/ab[5][21] ), .IN0(
        \mult_26/CARRYB[4][21] ), .IN1(\mult_26/SUMB[4][22] ), .COUT(
        \mult_26/CARRYB[5][21] ), .SUM(\mult_26/SUMB[5][21] ) );
  FADDER \mult_26/S2_5_20  ( .CIN(\mult_26/ab[5][20] ), .IN0(
        \mult_26/CARRYB[4][20] ), .IN1(\mult_26/SUMB[4][21] ), .COUT(
        \mult_26/CARRYB[5][20] ), .SUM(\mult_26/SUMB[5][20] ) );
  FADDER \mult_26/S2_5_19  ( .CIN(\mult_26/ab[5][19] ), .IN0(
        \mult_26/CARRYB[4][19] ), .IN1(\mult_26/SUMB[4][20] ), .COUT(
        \mult_26/CARRYB[5][19] ), .SUM(\mult_26/SUMB[5][19] ) );
  FADDER \mult_26/S2_5_18  ( .CIN(\mult_26/ab[5][18] ), .IN0(
        \mult_26/CARRYB[4][18] ), .IN1(\mult_26/SUMB[4][19] ), .COUT(
        \mult_26/CARRYB[5][18] ), .SUM(\mult_26/SUMB[5][18] ) );
  FADDER \mult_26/S2_5_17  ( .CIN(\mult_26/ab[5][17] ), .IN0(
        \mult_26/CARRYB[4][17] ), .IN1(\mult_26/SUMB[4][18] ), .COUT(
        \mult_26/CARRYB[5][17] ), .SUM(\mult_26/SUMB[5][17] ) );
  FADDER \mult_26/S2_5_16  ( .CIN(\mult_26/ab[5][16] ), .IN0(
        \mult_26/CARRYB[4][16] ), .IN1(\mult_26/SUMB[4][17] ), .COUT(
        \mult_26/CARRYB[5][16] ), .SUM(\mult_26/SUMB[5][16] ) );
  FADDER \mult_26/S2_5_15  ( .CIN(\mult_26/ab[5][15] ), .IN0(
        \mult_26/CARRYB[4][15] ), .IN1(\mult_26/SUMB[4][16] ), .COUT(
        \mult_26/CARRYB[5][15] ), .SUM(\mult_26/SUMB[5][15] ) );
  FADDER \mult_26/S2_5_14  ( .CIN(\mult_26/ab[5][14] ), .IN0(
        \mult_26/CARRYB[4][14] ), .IN1(\mult_26/SUMB[4][15] ), .COUT(
        \mult_26/CARRYB[5][14] ), .SUM(\mult_26/SUMB[5][14] ) );
  FADDER \mult_26/S2_5_13  ( .CIN(\mult_26/ab[5][13] ), .IN0(
        \mult_26/CARRYB[4][13] ), .IN1(\mult_26/SUMB[4][14] ), .COUT(
        \mult_26/CARRYB[5][13] ), .SUM(\mult_26/SUMB[5][13] ) );
  FADDER \mult_26/S2_5_12  ( .CIN(\mult_26/ab[5][12] ), .IN0(
        \mult_26/CARRYB[4][12] ), .IN1(\mult_26/SUMB[4][13] ), .COUT(
        \mult_26/CARRYB[5][12] ), .SUM(\mult_26/SUMB[5][12] ) );
  FADDER \mult_26/S2_5_11  ( .CIN(\mult_26/ab[5][11] ), .IN0(
        \mult_26/CARRYB[4][11] ), .IN1(\mult_26/SUMB[4][12] ), .COUT(
        \mult_26/CARRYB[5][11] ), .SUM(\mult_26/SUMB[5][11] ) );
  FADDER \mult_26/S2_5_10  ( .CIN(\mult_26/ab[5][10] ), .IN0(
        \mult_26/CARRYB[4][10] ), .IN1(\mult_26/SUMB[4][11] ), .COUT(
        \mult_26/CARRYB[5][10] ), .SUM(\mult_26/SUMB[5][10] ) );
  FADDER \mult_26/S2_5_9  ( .CIN(\mult_26/ab[5][9] ), .IN0(
        \mult_26/CARRYB[4][9] ), .IN1(\mult_26/SUMB[4][10] ), .COUT(
        \mult_26/CARRYB[5][9] ), .SUM(\mult_26/SUMB[5][9] ) );
  FADDER \mult_26/S2_5_8  ( .CIN(\mult_26/ab[5][8] ), .IN0(
        \mult_26/CARRYB[4][8] ), .IN1(\mult_26/SUMB[4][9] ), .COUT(
        \mult_26/CARRYB[5][8] ), .SUM(\mult_26/SUMB[5][8] ) );
  FADDER \mult_26/S2_5_7  ( .CIN(\mult_26/ab[5][7] ), .IN0(
        \mult_26/CARRYB[4][7] ), .IN1(\mult_26/SUMB[4][8] ), .COUT(
        \mult_26/CARRYB[5][7] ), .SUM(\mult_26/SUMB[5][7] ) );
  FADDER \mult_26/S2_5_6  ( .CIN(\mult_26/ab[5][6] ), .IN0(
        \mult_26/CARRYB[4][6] ), .IN1(\mult_26/SUMB[4][7] ), .COUT(
        \mult_26/CARRYB[5][6] ), .SUM(\mult_26/SUMB[5][6] ) );
  FADDER \mult_26/S2_5_5  ( .CIN(\mult_26/ab[5][5] ), .IN0(
        \mult_26/CARRYB[4][5] ), .IN1(\mult_26/SUMB[4][6] ), .COUT(
        \mult_26/CARRYB[5][5] ), .SUM(\mult_26/SUMB[5][5] ) );
  FADDER \mult_26/S2_5_4  ( .CIN(\mult_26/ab[5][4] ), .IN0(
        \mult_26/CARRYB[4][4] ), .IN1(\mult_26/SUMB[4][5] ), .COUT(
        \mult_26/CARRYB[5][4] ), .SUM(\mult_26/SUMB[5][4] ) );
  FADDER \mult_26/S2_5_3  ( .CIN(\mult_26/ab[5][3] ), .IN0(
        \mult_26/CARRYB[4][3] ), .IN1(\mult_26/SUMB[4][4] ), .COUT(
        \mult_26/CARRYB[5][3] ), .SUM(\mult_26/SUMB[5][3] ) );
  FADDER \mult_26/S2_5_2  ( .CIN(\mult_26/ab[5][2] ), .IN0(
        \mult_26/CARRYB[4][2] ), .IN1(\mult_26/SUMB[4][3] ), .COUT(
        \mult_26/CARRYB[5][2] ), .SUM(\mult_26/SUMB[5][2] ) );
  FADDER \mult_26/S2_5_1  ( .CIN(\mult_26/ab[5][1] ), .IN0(
        \mult_26/CARRYB[4][1] ), .IN1(\mult_26/SUMB[4][2] ), .COUT(
        \mult_26/CARRYB[5][1] ), .SUM(\mult_26/SUMB[5][1] ) );
  FADDER \mult_26/S1_5_0  ( .CIN(\mult_26/ab[5][0] ), .IN0(
        \mult_26/CARRYB[4][0] ), .IN1(\mult_26/SUMB[4][1] ), .COUT(
        \mult_26/CARRYB[5][0] ), .SUM(o[5]) );
  FADDER \mult_26/S3_6_30  ( .CIN(\mult_26/ab[6][30] ), .IN0(
        \mult_26/CARRYB[5][30] ), .IN1(\mult_26/ab[5][31] ), .COUT(
        \mult_26/CARRYB[6][30] ), .SUM(\mult_26/SUMB[6][30] ) );
  FADDER \mult_26/S2_6_29  ( .CIN(\mult_26/ab[6][29] ), .IN0(
        \mult_26/CARRYB[5][29] ), .IN1(\mult_26/SUMB[5][30] ), .COUT(
        \mult_26/CARRYB[6][29] ), .SUM(\mult_26/SUMB[6][29] ) );
  FADDER \mult_26/S2_6_28  ( .CIN(\mult_26/ab[6][28] ), .IN0(
        \mult_26/CARRYB[5][28] ), .IN1(\mult_26/SUMB[5][29] ), .COUT(
        \mult_26/CARRYB[6][28] ), .SUM(\mult_26/SUMB[6][28] ) );
  FADDER \mult_26/S2_6_27  ( .CIN(\mult_26/ab[6][27] ), .IN0(
        \mult_26/CARRYB[5][27] ), .IN1(\mult_26/SUMB[5][28] ), .COUT(
        \mult_26/CARRYB[6][27] ), .SUM(\mult_26/SUMB[6][27] ) );
  FADDER \mult_26/S2_6_26  ( .CIN(\mult_26/ab[6][26] ), .IN0(
        \mult_26/CARRYB[5][26] ), .IN1(\mult_26/SUMB[5][27] ), .COUT(
        \mult_26/CARRYB[6][26] ), .SUM(\mult_26/SUMB[6][26] ) );
  FADDER \mult_26/S2_6_25  ( .CIN(\mult_26/ab[6][25] ), .IN0(
        \mult_26/CARRYB[5][25] ), .IN1(\mult_26/SUMB[5][26] ), .COUT(
        \mult_26/CARRYB[6][25] ), .SUM(\mult_26/SUMB[6][25] ) );
  FADDER \mult_26/S2_6_24  ( .CIN(\mult_26/ab[6][24] ), .IN0(
        \mult_26/CARRYB[5][24] ), .IN1(\mult_26/SUMB[5][25] ), .COUT(
        \mult_26/CARRYB[6][24] ), .SUM(\mult_26/SUMB[6][24] ) );
  FADDER \mult_26/S2_6_23  ( .CIN(\mult_26/ab[6][23] ), .IN0(
        \mult_26/CARRYB[5][23] ), .IN1(\mult_26/SUMB[5][24] ), .COUT(
        \mult_26/CARRYB[6][23] ), .SUM(\mult_26/SUMB[6][23] ) );
  FADDER \mult_26/S2_6_22  ( .CIN(\mult_26/ab[6][22] ), .IN0(
        \mult_26/CARRYB[5][22] ), .IN1(\mult_26/SUMB[5][23] ), .COUT(
        \mult_26/CARRYB[6][22] ), .SUM(\mult_26/SUMB[6][22] ) );
  FADDER \mult_26/S2_6_21  ( .CIN(\mult_26/ab[6][21] ), .IN0(
        \mult_26/CARRYB[5][21] ), .IN1(\mult_26/SUMB[5][22] ), .COUT(
        \mult_26/CARRYB[6][21] ), .SUM(\mult_26/SUMB[6][21] ) );
  FADDER \mult_26/S2_6_20  ( .CIN(\mult_26/ab[6][20] ), .IN0(
        \mult_26/CARRYB[5][20] ), .IN1(\mult_26/SUMB[5][21] ), .COUT(
        \mult_26/CARRYB[6][20] ), .SUM(\mult_26/SUMB[6][20] ) );
  FADDER \mult_26/S2_6_19  ( .CIN(\mult_26/ab[6][19] ), .IN0(
        \mult_26/CARRYB[5][19] ), .IN1(\mult_26/SUMB[5][20] ), .COUT(
        \mult_26/CARRYB[6][19] ), .SUM(\mult_26/SUMB[6][19] ) );
  FADDER \mult_26/S2_6_18  ( .CIN(\mult_26/ab[6][18] ), .IN0(
        \mult_26/CARRYB[5][18] ), .IN1(\mult_26/SUMB[5][19] ), .COUT(
        \mult_26/CARRYB[6][18] ), .SUM(\mult_26/SUMB[6][18] ) );
  FADDER \mult_26/S2_6_17  ( .CIN(\mult_26/ab[6][17] ), .IN0(
        \mult_26/CARRYB[5][17] ), .IN1(\mult_26/SUMB[5][18] ), .COUT(
        \mult_26/CARRYB[6][17] ), .SUM(\mult_26/SUMB[6][17] ) );
  FADDER \mult_26/S2_6_16  ( .CIN(\mult_26/ab[6][16] ), .IN0(
        \mult_26/CARRYB[5][16] ), .IN1(\mult_26/SUMB[5][17] ), .COUT(
        \mult_26/CARRYB[6][16] ), .SUM(\mult_26/SUMB[6][16] ) );
  FADDER \mult_26/S2_6_15  ( .CIN(\mult_26/ab[6][15] ), .IN0(
        \mult_26/CARRYB[5][15] ), .IN1(\mult_26/SUMB[5][16] ), .COUT(
        \mult_26/CARRYB[6][15] ), .SUM(\mult_26/SUMB[6][15] ) );
  FADDER \mult_26/S2_6_14  ( .CIN(\mult_26/ab[6][14] ), .IN0(
        \mult_26/CARRYB[5][14] ), .IN1(\mult_26/SUMB[5][15] ), .COUT(
        \mult_26/CARRYB[6][14] ), .SUM(\mult_26/SUMB[6][14] ) );
  FADDER \mult_26/S2_6_13  ( .CIN(\mult_26/ab[6][13] ), .IN0(
        \mult_26/CARRYB[5][13] ), .IN1(\mult_26/SUMB[5][14] ), .COUT(
        \mult_26/CARRYB[6][13] ), .SUM(\mult_26/SUMB[6][13] ) );
  FADDER \mult_26/S2_6_12  ( .CIN(\mult_26/ab[6][12] ), .IN0(
        \mult_26/CARRYB[5][12] ), .IN1(\mult_26/SUMB[5][13] ), .COUT(
        \mult_26/CARRYB[6][12] ), .SUM(\mult_26/SUMB[6][12] ) );
  FADDER \mult_26/S2_6_11  ( .CIN(\mult_26/ab[6][11] ), .IN0(
        \mult_26/CARRYB[5][11] ), .IN1(\mult_26/SUMB[5][12] ), .COUT(
        \mult_26/CARRYB[6][11] ), .SUM(\mult_26/SUMB[6][11] ) );
  FADDER \mult_26/S2_6_10  ( .CIN(\mult_26/ab[6][10] ), .IN0(
        \mult_26/CARRYB[5][10] ), .IN1(\mult_26/SUMB[5][11] ), .COUT(
        \mult_26/CARRYB[6][10] ), .SUM(\mult_26/SUMB[6][10] ) );
  FADDER \mult_26/S2_6_9  ( .CIN(\mult_26/ab[6][9] ), .IN0(
        \mult_26/CARRYB[5][9] ), .IN1(\mult_26/SUMB[5][10] ), .COUT(
        \mult_26/CARRYB[6][9] ), .SUM(\mult_26/SUMB[6][9] ) );
  FADDER \mult_26/S2_6_8  ( .CIN(\mult_26/ab[6][8] ), .IN0(
        \mult_26/CARRYB[5][8] ), .IN1(\mult_26/SUMB[5][9] ), .COUT(
        \mult_26/CARRYB[6][8] ), .SUM(\mult_26/SUMB[6][8] ) );
  FADDER \mult_26/S2_6_7  ( .CIN(\mult_26/ab[6][7] ), .IN0(
        \mult_26/CARRYB[5][7] ), .IN1(\mult_26/SUMB[5][8] ), .COUT(
        \mult_26/CARRYB[6][7] ), .SUM(\mult_26/SUMB[6][7] ) );
  FADDER \mult_26/S2_6_6  ( .CIN(\mult_26/ab[6][6] ), .IN0(
        \mult_26/CARRYB[5][6] ), .IN1(\mult_26/SUMB[5][7] ), .COUT(
        \mult_26/CARRYB[6][6] ), .SUM(\mult_26/SUMB[6][6] ) );
  FADDER \mult_26/S2_6_5  ( .CIN(\mult_26/ab[6][5] ), .IN0(
        \mult_26/CARRYB[5][5] ), .IN1(\mult_26/SUMB[5][6] ), .COUT(
        \mult_26/CARRYB[6][5] ), .SUM(\mult_26/SUMB[6][5] ) );
  FADDER \mult_26/S2_6_4  ( .CIN(\mult_26/ab[6][4] ), .IN0(
        \mult_26/CARRYB[5][4] ), .IN1(\mult_26/SUMB[5][5] ), .COUT(
        \mult_26/CARRYB[6][4] ), .SUM(\mult_26/SUMB[6][4] ) );
  FADDER \mult_26/S2_6_3  ( .CIN(\mult_26/ab[6][3] ), .IN0(
        \mult_26/CARRYB[5][3] ), .IN1(\mult_26/SUMB[5][4] ), .COUT(
        \mult_26/CARRYB[6][3] ), .SUM(\mult_26/SUMB[6][3] ) );
  FADDER \mult_26/S2_6_2  ( .CIN(\mult_26/ab[6][2] ), .IN0(
        \mult_26/CARRYB[5][2] ), .IN1(\mult_26/SUMB[5][3] ), .COUT(
        \mult_26/CARRYB[6][2] ), .SUM(\mult_26/SUMB[6][2] ) );
  FADDER \mult_26/S2_6_1  ( .CIN(\mult_26/ab[6][1] ), .IN0(
        \mult_26/CARRYB[5][1] ), .IN1(\mult_26/SUMB[5][2] ), .COUT(
        \mult_26/CARRYB[6][1] ), .SUM(\mult_26/SUMB[6][1] ) );
  FADDER \mult_26/S1_6_0  ( .CIN(\mult_26/ab[6][0] ), .IN0(
        \mult_26/CARRYB[5][0] ), .IN1(\mult_26/SUMB[5][1] ), .COUT(
        \mult_26/CARRYB[6][0] ), .SUM(o[6]) );
  FADDER \mult_26/S3_7_30  ( .CIN(\mult_26/ab[7][30] ), .IN0(
        \mult_26/CARRYB[6][30] ), .IN1(\mult_26/ab[6][31] ), .COUT(
        \mult_26/CARRYB[7][30] ), .SUM(\mult_26/SUMB[7][30] ) );
  FADDER \mult_26/S2_7_29  ( .CIN(\mult_26/ab[7][29] ), .IN0(
        \mult_26/CARRYB[6][29] ), .IN1(\mult_26/SUMB[6][30] ), .COUT(
        \mult_26/CARRYB[7][29] ), .SUM(\mult_26/SUMB[7][29] ) );
  FADDER \mult_26/S2_7_28  ( .CIN(\mult_26/ab[7][28] ), .IN0(
        \mult_26/CARRYB[6][28] ), .IN1(\mult_26/SUMB[6][29] ), .COUT(
        \mult_26/CARRYB[7][28] ), .SUM(\mult_26/SUMB[7][28] ) );
  FADDER \mult_26/S2_7_27  ( .CIN(\mult_26/ab[7][27] ), .IN0(
        \mult_26/CARRYB[6][27] ), .IN1(\mult_26/SUMB[6][28] ), .COUT(
        \mult_26/CARRYB[7][27] ), .SUM(\mult_26/SUMB[7][27] ) );
  FADDER \mult_26/S2_7_26  ( .CIN(\mult_26/ab[7][26] ), .IN0(
        \mult_26/CARRYB[6][26] ), .IN1(\mult_26/SUMB[6][27] ), .COUT(
        \mult_26/CARRYB[7][26] ), .SUM(\mult_26/SUMB[7][26] ) );
  FADDER \mult_26/S2_7_25  ( .CIN(\mult_26/ab[7][25] ), .IN0(
        \mult_26/CARRYB[6][25] ), .IN1(\mult_26/SUMB[6][26] ), .COUT(
        \mult_26/CARRYB[7][25] ), .SUM(\mult_26/SUMB[7][25] ) );
  FADDER \mult_26/S2_7_24  ( .CIN(\mult_26/ab[7][24] ), .IN0(
        \mult_26/CARRYB[6][24] ), .IN1(\mult_26/SUMB[6][25] ), .COUT(
        \mult_26/CARRYB[7][24] ), .SUM(\mult_26/SUMB[7][24] ) );
  FADDER \mult_26/S2_7_23  ( .CIN(\mult_26/ab[7][23] ), .IN0(
        \mult_26/CARRYB[6][23] ), .IN1(\mult_26/SUMB[6][24] ), .COUT(
        \mult_26/CARRYB[7][23] ), .SUM(\mult_26/SUMB[7][23] ) );
  FADDER \mult_26/S2_7_22  ( .CIN(\mult_26/ab[7][22] ), .IN0(
        \mult_26/CARRYB[6][22] ), .IN1(\mult_26/SUMB[6][23] ), .COUT(
        \mult_26/CARRYB[7][22] ), .SUM(\mult_26/SUMB[7][22] ) );
  FADDER \mult_26/S2_7_21  ( .CIN(\mult_26/ab[7][21] ), .IN0(
        \mult_26/CARRYB[6][21] ), .IN1(\mult_26/SUMB[6][22] ), .COUT(
        \mult_26/CARRYB[7][21] ), .SUM(\mult_26/SUMB[7][21] ) );
  FADDER \mult_26/S2_7_20  ( .CIN(\mult_26/ab[7][20] ), .IN0(
        \mult_26/CARRYB[6][20] ), .IN1(\mult_26/SUMB[6][21] ), .COUT(
        \mult_26/CARRYB[7][20] ), .SUM(\mult_26/SUMB[7][20] ) );
  FADDER \mult_26/S2_7_19  ( .CIN(\mult_26/ab[7][19] ), .IN0(
        \mult_26/CARRYB[6][19] ), .IN1(\mult_26/SUMB[6][20] ), .COUT(
        \mult_26/CARRYB[7][19] ), .SUM(\mult_26/SUMB[7][19] ) );
  FADDER \mult_26/S2_7_18  ( .CIN(\mult_26/ab[7][18] ), .IN0(
        \mult_26/CARRYB[6][18] ), .IN1(\mult_26/SUMB[6][19] ), .COUT(
        \mult_26/CARRYB[7][18] ), .SUM(\mult_26/SUMB[7][18] ) );
  FADDER \mult_26/S2_7_17  ( .CIN(\mult_26/ab[7][17] ), .IN0(
        \mult_26/CARRYB[6][17] ), .IN1(\mult_26/SUMB[6][18] ), .COUT(
        \mult_26/CARRYB[7][17] ), .SUM(\mult_26/SUMB[7][17] ) );
  FADDER \mult_26/S2_7_16  ( .CIN(\mult_26/ab[7][16] ), .IN0(
        \mult_26/CARRYB[6][16] ), .IN1(\mult_26/SUMB[6][17] ), .COUT(
        \mult_26/CARRYB[7][16] ), .SUM(\mult_26/SUMB[7][16] ) );
  FADDER \mult_26/S2_7_15  ( .CIN(\mult_26/ab[7][15] ), .IN0(
        \mult_26/CARRYB[6][15] ), .IN1(\mult_26/SUMB[6][16] ), .COUT(
        \mult_26/CARRYB[7][15] ), .SUM(\mult_26/SUMB[7][15] ) );
  FADDER \mult_26/S2_7_14  ( .CIN(\mult_26/ab[7][14] ), .IN0(
        \mult_26/CARRYB[6][14] ), .IN1(\mult_26/SUMB[6][15] ), .COUT(
        \mult_26/CARRYB[7][14] ), .SUM(\mult_26/SUMB[7][14] ) );
  FADDER \mult_26/S2_7_13  ( .CIN(\mult_26/ab[7][13] ), .IN0(
        \mult_26/CARRYB[6][13] ), .IN1(\mult_26/SUMB[6][14] ), .COUT(
        \mult_26/CARRYB[7][13] ), .SUM(\mult_26/SUMB[7][13] ) );
  FADDER \mult_26/S2_7_12  ( .CIN(\mult_26/ab[7][12] ), .IN0(
        \mult_26/CARRYB[6][12] ), .IN1(\mult_26/SUMB[6][13] ), .COUT(
        \mult_26/CARRYB[7][12] ), .SUM(\mult_26/SUMB[7][12] ) );
  FADDER \mult_26/S2_7_11  ( .CIN(\mult_26/ab[7][11] ), .IN0(
        \mult_26/CARRYB[6][11] ), .IN1(\mult_26/SUMB[6][12] ), .COUT(
        \mult_26/CARRYB[7][11] ), .SUM(\mult_26/SUMB[7][11] ) );
  FADDER \mult_26/S2_7_10  ( .CIN(\mult_26/ab[7][10] ), .IN0(
        \mult_26/CARRYB[6][10] ), .IN1(\mult_26/SUMB[6][11] ), .COUT(
        \mult_26/CARRYB[7][10] ), .SUM(\mult_26/SUMB[7][10] ) );
  FADDER \mult_26/S2_7_9  ( .CIN(\mult_26/ab[7][9] ), .IN0(
        \mult_26/CARRYB[6][9] ), .IN1(\mult_26/SUMB[6][10] ), .COUT(
        \mult_26/CARRYB[7][9] ), .SUM(\mult_26/SUMB[7][9] ) );
  FADDER \mult_26/S2_7_8  ( .CIN(\mult_26/ab[7][8] ), .IN0(
        \mult_26/CARRYB[6][8] ), .IN1(\mult_26/SUMB[6][9] ), .COUT(
        \mult_26/CARRYB[7][8] ), .SUM(\mult_26/SUMB[7][8] ) );
  FADDER \mult_26/S2_7_7  ( .CIN(\mult_26/ab[7][7] ), .IN0(
        \mult_26/CARRYB[6][7] ), .IN1(\mult_26/SUMB[6][8] ), .COUT(
        \mult_26/CARRYB[7][7] ), .SUM(\mult_26/SUMB[7][7] ) );
  FADDER \mult_26/S2_7_6  ( .CIN(\mult_26/ab[7][6] ), .IN0(
        \mult_26/CARRYB[6][6] ), .IN1(\mult_26/SUMB[6][7] ), .COUT(
        \mult_26/CARRYB[7][6] ), .SUM(\mult_26/SUMB[7][6] ) );
  FADDER \mult_26/S2_7_5  ( .CIN(\mult_26/ab[7][5] ), .IN0(
        \mult_26/CARRYB[6][5] ), .IN1(\mult_26/SUMB[6][6] ), .COUT(
        \mult_26/CARRYB[7][5] ), .SUM(\mult_26/SUMB[7][5] ) );
  FADDER \mult_26/S2_7_4  ( .CIN(\mult_26/ab[7][4] ), .IN0(
        \mult_26/CARRYB[6][4] ), .IN1(\mult_26/SUMB[6][5] ), .COUT(
        \mult_26/CARRYB[7][4] ), .SUM(\mult_26/SUMB[7][4] ) );
  FADDER \mult_26/S2_7_3  ( .CIN(\mult_26/ab[7][3] ), .IN0(
        \mult_26/CARRYB[6][3] ), .IN1(\mult_26/SUMB[6][4] ), .COUT(
        \mult_26/CARRYB[7][3] ), .SUM(\mult_26/SUMB[7][3] ) );
  FADDER \mult_26/S2_7_2  ( .CIN(\mult_26/ab[7][2] ), .IN0(
        \mult_26/CARRYB[6][2] ), .IN1(\mult_26/SUMB[6][3] ), .COUT(
        \mult_26/CARRYB[7][2] ), .SUM(\mult_26/SUMB[7][2] ) );
  FADDER \mult_26/S2_7_1  ( .CIN(\mult_26/ab[7][1] ), .IN0(
        \mult_26/CARRYB[6][1] ), .IN1(\mult_26/SUMB[6][2] ), .COUT(
        \mult_26/CARRYB[7][1] ), .SUM(\mult_26/SUMB[7][1] ) );
  FADDER \mult_26/S1_7_0  ( .CIN(\mult_26/ab[7][0] ), .IN0(
        \mult_26/CARRYB[6][0] ), .IN1(\mult_26/SUMB[6][1] ), .COUT(
        \mult_26/CARRYB[7][0] ), .SUM(o[7]) );
  FADDER \mult_26/S3_8_30  ( .CIN(\mult_26/ab[8][30] ), .IN0(
        \mult_26/CARRYB[7][30] ), .IN1(\mult_26/ab[7][31] ), .COUT(
        \mult_26/CARRYB[8][30] ), .SUM(\mult_26/SUMB[8][30] ) );
  FADDER \mult_26/S2_8_29  ( .CIN(\mult_26/ab[8][29] ), .IN0(
        \mult_26/CARRYB[7][29] ), .IN1(\mult_26/SUMB[7][30] ), .COUT(
        \mult_26/CARRYB[8][29] ), .SUM(\mult_26/SUMB[8][29] ) );
  FADDER \mult_26/S2_8_28  ( .CIN(\mult_26/ab[8][28] ), .IN0(
        \mult_26/CARRYB[7][28] ), .IN1(\mult_26/SUMB[7][29] ), .COUT(
        \mult_26/CARRYB[8][28] ), .SUM(\mult_26/SUMB[8][28] ) );
  FADDER \mult_26/S2_8_27  ( .CIN(\mult_26/ab[8][27] ), .IN0(
        \mult_26/CARRYB[7][27] ), .IN1(\mult_26/SUMB[7][28] ), .COUT(
        \mult_26/CARRYB[8][27] ), .SUM(\mult_26/SUMB[8][27] ) );
  FADDER \mult_26/S2_8_26  ( .CIN(\mult_26/ab[8][26] ), .IN0(
        \mult_26/CARRYB[7][26] ), .IN1(\mult_26/SUMB[7][27] ), .COUT(
        \mult_26/CARRYB[8][26] ), .SUM(\mult_26/SUMB[8][26] ) );
  FADDER \mult_26/S2_8_25  ( .CIN(\mult_26/ab[8][25] ), .IN0(
        \mult_26/CARRYB[7][25] ), .IN1(\mult_26/SUMB[7][26] ), .COUT(
        \mult_26/CARRYB[8][25] ), .SUM(\mult_26/SUMB[8][25] ) );
  FADDER \mult_26/S2_8_24  ( .CIN(\mult_26/ab[8][24] ), .IN0(
        \mult_26/CARRYB[7][24] ), .IN1(\mult_26/SUMB[7][25] ), .COUT(
        \mult_26/CARRYB[8][24] ), .SUM(\mult_26/SUMB[8][24] ) );
  FADDER \mult_26/S2_8_23  ( .CIN(\mult_26/ab[8][23] ), .IN0(
        \mult_26/CARRYB[7][23] ), .IN1(\mult_26/SUMB[7][24] ), .COUT(
        \mult_26/CARRYB[8][23] ), .SUM(\mult_26/SUMB[8][23] ) );
  FADDER \mult_26/S2_8_22  ( .CIN(\mult_26/ab[8][22] ), .IN0(
        \mult_26/CARRYB[7][22] ), .IN1(\mult_26/SUMB[7][23] ), .COUT(
        \mult_26/CARRYB[8][22] ), .SUM(\mult_26/SUMB[8][22] ) );
  FADDER \mult_26/S2_8_21  ( .CIN(\mult_26/ab[8][21] ), .IN0(
        \mult_26/CARRYB[7][21] ), .IN1(\mult_26/SUMB[7][22] ), .COUT(
        \mult_26/CARRYB[8][21] ), .SUM(\mult_26/SUMB[8][21] ) );
  FADDER \mult_26/S2_8_20  ( .CIN(\mult_26/ab[8][20] ), .IN0(
        \mult_26/CARRYB[7][20] ), .IN1(\mult_26/SUMB[7][21] ), .COUT(
        \mult_26/CARRYB[8][20] ), .SUM(\mult_26/SUMB[8][20] ) );
  FADDER \mult_26/S2_8_19  ( .CIN(\mult_26/ab[8][19] ), .IN0(
        \mult_26/CARRYB[7][19] ), .IN1(\mult_26/SUMB[7][20] ), .COUT(
        \mult_26/CARRYB[8][19] ), .SUM(\mult_26/SUMB[8][19] ) );
  FADDER \mult_26/S2_8_18  ( .CIN(\mult_26/ab[8][18] ), .IN0(
        \mult_26/CARRYB[7][18] ), .IN1(\mult_26/SUMB[7][19] ), .COUT(
        \mult_26/CARRYB[8][18] ), .SUM(\mult_26/SUMB[8][18] ) );
  FADDER \mult_26/S2_8_17  ( .CIN(\mult_26/ab[8][17] ), .IN0(
        \mult_26/CARRYB[7][17] ), .IN1(\mult_26/SUMB[7][18] ), .COUT(
        \mult_26/CARRYB[8][17] ), .SUM(\mult_26/SUMB[8][17] ) );
  FADDER \mult_26/S2_8_16  ( .CIN(\mult_26/ab[8][16] ), .IN0(
        \mult_26/CARRYB[7][16] ), .IN1(\mult_26/SUMB[7][17] ), .COUT(
        \mult_26/CARRYB[8][16] ), .SUM(\mult_26/SUMB[8][16] ) );
  FADDER \mult_26/S2_8_15  ( .CIN(\mult_26/ab[8][15] ), .IN0(
        \mult_26/CARRYB[7][15] ), .IN1(\mult_26/SUMB[7][16] ), .COUT(
        \mult_26/CARRYB[8][15] ), .SUM(\mult_26/SUMB[8][15] ) );
  FADDER \mult_26/S2_8_14  ( .CIN(\mult_26/ab[8][14] ), .IN0(
        \mult_26/CARRYB[7][14] ), .IN1(\mult_26/SUMB[7][15] ), .COUT(
        \mult_26/CARRYB[8][14] ), .SUM(\mult_26/SUMB[8][14] ) );
  FADDER \mult_26/S2_8_13  ( .CIN(\mult_26/ab[8][13] ), .IN0(
        \mult_26/CARRYB[7][13] ), .IN1(\mult_26/SUMB[7][14] ), .COUT(
        \mult_26/CARRYB[8][13] ), .SUM(\mult_26/SUMB[8][13] ) );
  FADDER \mult_26/S2_8_12  ( .CIN(\mult_26/ab[8][12] ), .IN0(
        \mult_26/CARRYB[7][12] ), .IN1(\mult_26/SUMB[7][13] ), .COUT(
        \mult_26/CARRYB[8][12] ), .SUM(\mult_26/SUMB[8][12] ) );
  FADDER \mult_26/S2_8_11  ( .CIN(\mult_26/ab[8][11] ), .IN0(
        \mult_26/CARRYB[7][11] ), .IN1(\mult_26/SUMB[7][12] ), .COUT(
        \mult_26/CARRYB[8][11] ), .SUM(\mult_26/SUMB[8][11] ) );
  FADDER \mult_26/S2_8_10  ( .CIN(\mult_26/ab[8][10] ), .IN0(
        \mult_26/CARRYB[7][10] ), .IN1(\mult_26/SUMB[7][11] ), .COUT(
        \mult_26/CARRYB[8][10] ), .SUM(\mult_26/SUMB[8][10] ) );
  FADDER \mult_26/S2_8_9  ( .CIN(\mult_26/ab[8][9] ), .IN0(
        \mult_26/CARRYB[7][9] ), .IN1(\mult_26/SUMB[7][10] ), .COUT(
        \mult_26/CARRYB[8][9] ), .SUM(\mult_26/SUMB[8][9] ) );
  FADDER \mult_26/S2_8_8  ( .CIN(\mult_26/ab[8][8] ), .IN0(
        \mult_26/CARRYB[7][8] ), .IN1(\mult_26/SUMB[7][9] ), .COUT(
        \mult_26/CARRYB[8][8] ), .SUM(\mult_26/SUMB[8][8] ) );
  FADDER \mult_26/S2_8_7  ( .CIN(\mult_26/ab[8][7] ), .IN0(
        \mult_26/CARRYB[7][7] ), .IN1(\mult_26/SUMB[7][8] ), .COUT(
        \mult_26/CARRYB[8][7] ), .SUM(\mult_26/SUMB[8][7] ) );
  FADDER \mult_26/S2_8_6  ( .CIN(\mult_26/ab[8][6] ), .IN0(
        \mult_26/CARRYB[7][6] ), .IN1(\mult_26/SUMB[7][7] ), .COUT(
        \mult_26/CARRYB[8][6] ), .SUM(\mult_26/SUMB[8][6] ) );
  FADDER \mult_26/S2_8_5  ( .CIN(\mult_26/ab[8][5] ), .IN0(
        \mult_26/CARRYB[7][5] ), .IN1(\mult_26/SUMB[7][6] ), .COUT(
        \mult_26/CARRYB[8][5] ), .SUM(\mult_26/SUMB[8][5] ) );
  FADDER \mult_26/S2_8_4  ( .CIN(\mult_26/ab[8][4] ), .IN0(
        \mult_26/CARRYB[7][4] ), .IN1(\mult_26/SUMB[7][5] ), .COUT(
        \mult_26/CARRYB[8][4] ), .SUM(\mult_26/SUMB[8][4] ) );
  FADDER \mult_26/S2_8_3  ( .CIN(\mult_26/ab[8][3] ), .IN0(
        \mult_26/CARRYB[7][3] ), .IN1(\mult_26/SUMB[7][4] ), .COUT(
        \mult_26/CARRYB[8][3] ), .SUM(\mult_26/SUMB[8][3] ) );
  FADDER \mult_26/S2_8_2  ( .CIN(\mult_26/ab[8][2] ), .IN0(
        \mult_26/CARRYB[7][2] ), .IN1(\mult_26/SUMB[7][3] ), .COUT(
        \mult_26/CARRYB[8][2] ), .SUM(\mult_26/SUMB[8][2] ) );
  FADDER \mult_26/S2_8_1  ( .CIN(\mult_26/ab[8][1] ), .IN0(
        \mult_26/CARRYB[7][1] ), .IN1(\mult_26/SUMB[7][2] ), .COUT(
        \mult_26/CARRYB[8][1] ), .SUM(\mult_26/SUMB[8][1] ) );
  FADDER \mult_26/S1_8_0  ( .CIN(\mult_26/ab[8][0] ), .IN0(
        \mult_26/CARRYB[7][0] ), .IN1(\mult_26/SUMB[7][1] ), .COUT(
        \mult_26/CARRYB[8][0] ), .SUM(o[8]) );
  FADDER \mult_26/S3_9_30  ( .CIN(\mult_26/ab[9][30] ), .IN0(
        \mult_26/CARRYB[8][30] ), .IN1(\mult_26/ab[8][31] ), .COUT(
        \mult_26/CARRYB[9][30] ), .SUM(\mult_26/SUMB[9][30] ) );
  FADDER \mult_26/S2_9_29  ( .CIN(\mult_26/ab[9][29] ), .IN0(
        \mult_26/CARRYB[8][29] ), .IN1(\mult_26/SUMB[8][30] ), .COUT(
        \mult_26/CARRYB[9][29] ), .SUM(\mult_26/SUMB[9][29] ) );
  FADDER \mult_26/S2_9_28  ( .CIN(\mult_26/ab[9][28] ), .IN0(
        \mult_26/CARRYB[8][28] ), .IN1(\mult_26/SUMB[8][29] ), .COUT(
        \mult_26/CARRYB[9][28] ), .SUM(\mult_26/SUMB[9][28] ) );
  FADDER \mult_26/S2_9_27  ( .CIN(\mult_26/ab[9][27] ), .IN0(
        \mult_26/CARRYB[8][27] ), .IN1(\mult_26/SUMB[8][28] ), .COUT(
        \mult_26/CARRYB[9][27] ), .SUM(\mult_26/SUMB[9][27] ) );
  FADDER \mult_26/S2_9_26  ( .CIN(\mult_26/ab[9][26] ), .IN0(
        \mult_26/CARRYB[8][26] ), .IN1(\mult_26/SUMB[8][27] ), .COUT(
        \mult_26/CARRYB[9][26] ), .SUM(\mult_26/SUMB[9][26] ) );
  FADDER \mult_26/S2_9_25  ( .CIN(\mult_26/ab[9][25] ), .IN0(
        \mult_26/CARRYB[8][25] ), .IN1(\mult_26/SUMB[8][26] ), .COUT(
        \mult_26/CARRYB[9][25] ), .SUM(\mult_26/SUMB[9][25] ) );
  FADDER \mult_26/S2_9_24  ( .CIN(\mult_26/ab[9][24] ), .IN0(
        \mult_26/CARRYB[8][24] ), .IN1(\mult_26/SUMB[8][25] ), .COUT(
        \mult_26/CARRYB[9][24] ), .SUM(\mult_26/SUMB[9][24] ) );
  FADDER \mult_26/S2_9_23  ( .CIN(\mult_26/ab[9][23] ), .IN0(
        \mult_26/CARRYB[8][23] ), .IN1(\mult_26/SUMB[8][24] ), .COUT(
        \mult_26/CARRYB[9][23] ), .SUM(\mult_26/SUMB[9][23] ) );
  FADDER \mult_26/S2_9_22  ( .CIN(\mult_26/ab[9][22] ), .IN0(
        \mult_26/CARRYB[8][22] ), .IN1(\mult_26/SUMB[8][23] ), .COUT(
        \mult_26/CARRYB[9][22] ), .SUM(\mult_26/SUMB[9][22] ) );
  FADDER \mult_26/S2_9_21  ( .CIN(\mult_26/ab[9][21] ), .IN0(
        \mult_26/CARRYB[8][21] ), .IN1(\mult_26/SUMB[8][22] ), .COUT(
        \mult_26/CARRYB[9][21] ), .SUM(\mult_26/SUMB[9][21] ) );
  FADDER \mult_26/S2_9_20  ( .CIN(\mult_26/ab[9][20] ), .IN0(
        \mult_26/CARRYB[8][20] ), .IN1(\mult_26/SUMB[8][21] ), .COUT(
        \mult_26/CARRYB[9][20] ), .SUM(\mult_26/SUMB[9][20] ) );
  FADDER \mult_26/S2_9_19  ( .CIN(\mult_26/ab[9][19] ), .IN0(
        \mult_26/CARRYB[8][19] ), .IN1(\mult_26/SUMB[8][20] ), .COUT(
        \mult_26/CARRYB[9][19] ), .SUM(\mult_26/SUMB[9][19] ) );
  FADDER \mult_26/S2_9_18  ( .CIN(\mult_26/ab[9][18] ), .IN0(
        \mult_26/CARRYB[8][18] ), .IN1(\mult_26/SUMB[8][19] ), .COUT(
        \mult_26/CARRYB[9][18] ), .SUM(\mult_26/SUMB[9][18] ) );
  FADDER \mult_26/S2_9_17  ( .CIN(\mult_26/ab[9][17] ), .IN0(
        \mult_26/CARRYB[8][17] ), .IN1(\mult_26/SUMB[8][18] ), .COUT(
        \mult_26/CARRYB[9][17] ), .SUM(\mult_26/SUMB[9][17] ) );
  FADDER \mult_26/S2_9_16  ( .CIN(\mult_26/ab[9][16] ), .IN0(
        \mult_26/CARRYB[8][16] ), .IN1(\mult_26/SUMB[8][17] ), .COUT(
        \mult_26/CARRYB[9][16] ), .SUM(\mult_26/SUMB[9][16] ) );
  FADDER \mult_26/S2_9_15  ( .CIN(\mult_26/ab[9][15] ), .IN0(
        \mult_26/CARRYB[8][15] ), .IN1(\mult_26/SUMB[8][16] ), .COUT(
        \mult_26/CARRYB[9][15] ), .SUM(\mult_26/SUMB[9][15] ) );
  FADDER \mult_26/S2_9_14  ( .CIN(\mult_26/ab[9][14] ), .IN0(
        \mult_26/CARRYB[8][14] ), .IN1(\mult_26/SUMB[8][15] ), .COUT(
        \mult_26/CARRYB[9][14] ), .SUM(\mult_26/SUMB[9][14] ) );
  FADDER \mult_26/S2_9_13  ( .CIN(\mult_26/ab[9][13] ), .IN0(
        \mult_26/CARRYB[8][13] ), .IN1(\mult_26/SUMB[8][14] ), .COUT(
        \mult_26/CARRYB[9][13] ), .SUM(\mult_26/SUMB[9][13] ) );
  FADDER \mult_26/S2_9_12  ( .CIN(\mult_26/ab[9][12] ), .IN0(
        \mult_26/CARRYB[8][12] ), .IN1(\mult_26/SUMB[8][13] ), .COUT(
        \mult_26/CARRYB[9][12] ), .SUM(\mult_26/SUMB[9][12] ) );
  FADDER \mult_26/S2_9_11  ( .CIN(\mult_26/ab[9][11] ), .IN0(
        \mult_26/CARRYB[8][11] ), .IN1(\mult_26/SUMB[8][12] ), .COUT(
        \mult_26/CARRYB[9][11] ), .SUM(\mult_26/SUMB[9][11] ) );
  FADDER \mult_26/S2_9_10  ( .CIN(\mult_26/ab[9][10] ), .IN0(
        \mult_26/CARRYB[8][10] ), .IN1(\mult_26/SUMB[8][11] ), .COUT(
        \mult_26/CARRYB[9][10] ), .SUM(\mult_26/SUMB[9][10] ) );
  FADDER \mult_26/S2_9_9  ( .CIN(\mult_26/ab[9][9] ), .IN0(
        \mult_26/CARRYB[8][9] ), .IN1(\mult_26/SUMB[8][10] ), .COUT(
        \mult_26/CARRYB[9][9] ), .SUM(\mult_26/SUMB[9][9] ) );
  FADDER \mult_26/S2_9_8  ( .CIN(\mult_26/ab[9][8] ), .IN0(
        \mult_26/CARRYB[8][8] ), .IN1(\mult_26/SUMB[8][9] ), .COUT(
        \mult_26/CARRYB[9][8] ), .SUM(\mult_26/SUMB[9][8] ) );
  FADDER \mult_26/S2_9_7  ( .CIN(\mult_26/ab[9][7] ), .IN0(
        \mult_26/CARRYB[8][7] ), .IN1(\mult_26/SUMB[8][8] ), .COUT(
        \mult_26/CARRYB[9][7] ), .SUM(\mult_26/SUMB[9][7] ) );
  FADDER \mult_26/S2_9_6  ( .CIN(\mult_26/ab[9][6] ), .IN0(
        \mult_26/CARRYB[8][6] ), .IN1(\mult_26/SUMB[8][7] ), .COUT(
        \mult_26/CARRYB[9][6] ), .SUM(\mult_26/SUMB[9][6] ) );
  FADDER \mult_26/S2_9_5  ( .CIN(\mult_26/ab[9][5] ), .IN0(
        \mult_26/CARRYB[8][5] ), .IN1(\mult_26/SUMB[8][6] ), .COUT(
        \mult_26/CARRYB[9][5] ), .SUM(\mult_26/SUMB[9][5] ) );
  FADDER \mult_26/S2_9_4  ( .CIN(\mult_26/ab[9][4] ), .IN0(
        \mult_26/CARRYB[8][4] ), .IN1(\mult_26/SUMB[8][5] ), .COUT(
        \mult_26/CARRYB[9][4] ), .SUM(\mult_26/SUMB[9][4] ) );
  FADDER \mult_26/S2_9_3  ( .CIN(\mult_26/ab[9][3] ), .IN0(
        \mult_26/CARRYB[8][3] ), .IN1(\mult_26/SUMB[8][4] ), .COUT(
        \mult_26/CARRYB[9][3] ), .SUM(\mult_26/SUMB[9][3] ) );
  FADDER \mult_26/S2_9_2  ( .CIN(\mult_26/ab[9][2] ), .IN0(
        \mult_26/CARRYB[8][2] ), .IN1(\mult_26/SUMB[8][3] ), .COUT(
        \mult_26/CARRYB[9][2] ), .SUM(\mult_26/SUMB[9][2] ) );
  FADDER \mult_26/S2_9_1  ( .CIN(\mult_26/ab[9][1] ), .IN0(
        \mult_26/CARRYB[8][1] ), .IN1(\mult_26/SUMB[8][2] ), .COUT(
        \mult_26/CARRYB[9][1] ), .SUM(\mult_26/SUMB[9][1] ) );
  FADDER \mult_26/S1_9_0  ( .CIN(\mult_26/ab[9][0] ), .IN0(
        \mult_26/CARRYB[8][0] ), .IN1(\mult_26/SUMB[8][1] ), .COUT(
        \mult_26/CARRYB[9][0] ), .SUM(o[9]) );
  FADDER \mult_26/S3_10_30  ( .CIN(\mult_26/ab[10][30] ), .IN0(
        \mult_26/CARRYB[9][30] ), .IN1(\mult_26/ab[9][31] ), .COUT(
        \mult_26/CARRYB[10][30] ), .SUM(\mult_26/SUMB[10][30] ) );
  FADDER \mult_26/S2_10_29  ( .CIN(\mult_26/ab[10][29] ), .IN0(
        \mult_26/CARRYB[9][29] ), .IN1(\mult_26/SUMB[9][30] ), .COUT(
        \mult_26/CARRYB[10][29] ), .SUM(\mult_26/SUMB[10][29] ) );
  FADDER \mult_26/S2_10_28  ( .CIN(\mult_26/ab[10][28] ), .IN0(
        \mult_26/CARRYB[9][28] ), .IN1(\mult_26/SUMB[9][29] ), .COUT(
        \mult_26/CARRYB[10][28] ), .SUM(\mult_26/SUMB[10][28] ) );
  FADDER \mult_26/S2_10_27  ( .CIN(\mult_26/ab[10][27] ), .IN0(
        \mult_26/CARRYB[9][27] ), .IN1(\mult_26/SUMB[9][28] ), .COUT(
        \mult_26/CARRYB[10][27] ), .SUM(\mult_26/SUMB[10][27] ) );
  FADDER \mult_26/S2_10_26  ( .CIN(\mult_26/ab[10][26] ), .IN0(
        \mult_26/CARRYB[9][26] ), .IN1(\mult_26/SUMB[9][27] ), .COUT(
        \mult_26/CARRYB[10][26] ), .SUM(\mult_26/SUMB[10][26] ) );
  FADDER \mult_26/S2_10_25  ( .CIN(\mult_26/ab[10][25] ), .IN0(
        \mult_26/CARRYB[9][25] ), .IN1(\mult_26/SUMB[9][26] ), .COUT(
        \mult_26/CARRYB[10][25] ), .SUM(\mult_26/SUMB[10][25] ) );
  FADDER \mult_26/S2_10_24  ( .CIN(\mult_26/ab[10][24] ), .IN0(
        \mult_26/CARRYB[9][24] ), .IN1(\mult_26/SUMB[9][25] ), .COUT(
        \mult_26/CARRYB[10][24] ), .SUM(\mult_26/SUMB[10][24] ) );
  FADDER \mult_26/S2_10_23  ( .CIN(\mult_26/ab[10][23] ), .IN0(
        \mult_26/CARRYB[9][23] ), .IN1(\mult_26/SUMB[9][24] ), .COUT(
        \mult_26/CARRYB[10][23] ), .SUM(\mult_26/SUMB[10][23] ) );
  FADDER \mult_26/S2_10_22  ( .CIN(\mult_26/ab[10][22] ), .IN0(
        \mult_26/CARRYB[9][22] ), .IN1(\mult_26/SUMB[9][23] ), .COUT(
        \mult_26/CARRYB[10][22] ), .SUM(\mult_26/SUMB[10][22] ) );
  FADDER \mult_26/S2_10_21  ( .CIN(\mult_26/ab[10][21] ), .IN0(
        \mult_26/CARRYB[9][21] ), .IN1(\mult_26/SUMB[9][22] ), .COUT(
        \mult_26/CARRYB[10][21] ), .SUM(\mult_26/SUMB[10][21] ) );
  FADDER \mult_26/S2_10_20  ( .CIN(\mult_26/ab[10][20] ), .IN0(
        \mult_26/CARRYB[9][20] ), .IN1(\mult_26/SUMB[9][21] ), .COUT(
        \mult_26/CARRYB[10][20] ), .SUM(\mult_26/SUMB[10][20] ) );
  FADDER \mult_26/S2_10_19  ( .CIN(\mult_26/ab[10][19] ), .IN0(
        \mult_26/CARRYB[9][19] ), .IN1(\mult_26/SUMB[9][20] ), .COUT(
        \mult_26/CARRYB[10][19] ), .SUM(\mult_26/SUMB[10][19] ) );
  FADDER \mult_26/S2_10_18  ( .CIN(\mult_26/ab[10][18] ), .IN0(
        \mult_26/CARRYB[9][18] ), .IN1(\mult_26/SUMB[9][19] ), .COUT(
        \mult_26/CARRYB[10][18] ), .SUM(\mult_26/SUMB[10][18] ) );
  FADDER \mult_26/S2_10_17  ( .CIN(\mult_26/ab[10][17] ), .IN0(
        \mult_26/CARRYB[9][17] ), .IN1(\mult_26/SUMB[9][18] ), .COUT(
        \mult_26/CARRYB[10][17] ), .SUM(\mult_26/SUMB[10][17] ) );
  FADDER \mult_26/S2_10_16  ( .CIN(\mult_26/ab[10][16] ), .IN0(
        \mult_26/CARRYB[9][16] ), .IN1(\mult_26/SUMB[9][17] ), .COUT(
        \mult_26/CARRYB[10][16] ), .SUM(\mult_26/SUMB[10][16] ) );
  FADDER \mult_26/S2_10_15  ( .CIN(\mult_26/ab[10][15] ), .IN0(
        \mult_26/CARRYB[9][15] ), .IN1(\mult_26/SUMB[9][16] ), .COUT(
        \mult_26/CARRYB[10][15] ), .SUM(\mult_26/SUMB[10][15] ) );
  FADDER \mult_26/S2_10_14  ( .CIN(\mult_26/ab[10][14] ), .IN0(
        \mult_26/CARRYB[9][14] ), .IN1(\mult_26/SUMB[9][15] ), .COUT(
        \mult_26/CARRYB[10][14] ), .SUM(\mult_26/SUMB[10][14] ) );
  FADDER \mult_26/S2_10_13  ( .CIN(\mult_26/ab[10][13] ), .IN0(
        \mult_26/CARRYB[9][13] ), .IN1(\mult_26/SUMB[9][14] ), .COUT(
        \mult_26/CARRYB[10][13] ), .SUM(\mult_26/SUMB[10][13] ) );
  FADDER \mult_26/S2_10_12  ( .CIN(\mult_26/ab[10][12] ), .IN0(
        \mult_26/CARRYB[9][12] ), .IN1(\mult_26/SUMB[9][13] ), .COUT(
        \mult_26/CARRYB[10][12] ), .SUM(\mult_26/SUMB[10][12] ) );
  FADDER \mult_26/S2_10_11  ( .CIN(\mult_26/ab[10][11] ), .IN0(
        \mult_26/CARRYB[9][11] ), .IN1(\mult_26/SUMB[9][12] ), .COUT(
        \mult_26/CARRYB[10][11] ), .SUM(\mult_26/SUMB[10][11] ) );
  FADDER \mult_26/S2_10_10  ( .CIN(\mult_26/ab[10][10] ), .IN0(
        \mult_26/CARRYB[9][10] ), .IN1(\mult_26/SUMB[9][11] ), .COUT(
        \mult_26/CARRYB[10][10] ), .SUM(\mult_26/SUMB[10][10] ) );
  FADDER \mult_26/S2_10_9  ( .CIN(\mult_26/ab[10][9] ), .IN0(
        \mult_26/CARRYB[9][9] ), .IN1(\mult_26/SUMB[9][10] ), .COUT(
        \mult_26/CARRYB[10][9] ), .SUM(\mult_26/SUMB[10][9] ) );
  FADDER \mult_26/S2_10_8  ( .CIN(\mult_26/ab[10][8] ), .IN0(
        \mult_26/CARRYB[9][8] ), .IN1(\mult_26/SUMB[9][9] ), .COUT(
        \mult_26/CARRYB[10][8] ), .SUM(\mult_26/SUMB[10][8] ) );
  FADDER \mult_26/S2_10_7  ( .CIN(\mult_26/ab[10][7] ), .IN0(
        \mult_26/CARRYB[9][7] ), .IN1(\mult_26/SUMB[9][8] ), .COUT(
        \mult_26/CARRYB[10][7] ), .SUM(\mult_26/SUMB[10][7] ) );
  FADDER \mult_26/S2_10_6  ( .CIN(\mult_26/ab[10][6] ), .IN0(
        \mult_26/CARRYB[9][6] ), .IN1(\mult_26/SUMB[9][7] ), .COUT(
        \mult_26/CARRYB[10][6] ), .SUM(\mult_26/SUMB[10][6] ) );
  FADDER \mult_26/S2_10_5  ( .CIN(\mult_26/ab[10][5] ), .IN0(
        \mult_26/CARRYB[9][5] ), .IN1(\mult_26/SUMB[9][6] ), .COUT(
        \mult_26/CARRYB[10][5] ), .SUM(\mult_26/SUMB[10][5] ) );
  FADDER \mult_26/S2_10_4  ( .CIN(\mult_26/ab[10][4] ), .IN0(
        \mult_26/CARRYB[9][4] ), .IN1(\mult_26/SUMB[9][5] ), .COUT(
        \mult_26/CARRYB[10][4] ), .SUM(\mult_26/SUMB[10][4] ) );
  FADDER \mult_26/S2_10_3  ( .CIN(\mult_26/ab[10][3] ), .IN0(
        \mult_26/CARRYB[9][3] ), .IN1(\mult_26/SUMB[9][4] ), .COUT(
        \mult_26/CARRYB[10][3] ), .SUM(\mult_26/SUMB[10][3] ) );
  FADDER \mult_26/S2_10_2  ( .CIN(\mult_26/ab[10][2] ), .IN0(
        \mult_26/CARRYB[9][2] ), .IN1(\mult_26/SUMB[9][3] ), .COUT(
        \mult_26/CARRYB[10][2] ), .SUM(\mult_26/SUMB[10][2] ) );
  FADDER \mult_26/S2_10_1  ( .CIN(\mult_26/ab[10][1] ), .IN0(
        \mult_26/CARRYB[9][1] ), .IN1(\mult_26/SUMB[9][2] ), .COUT(
        \mult_26/CARRYB[10][1] ), .SUM(\mult_26/SUMB[10][1] ) );
  FADDER \mult_26/S1_10_0  ( .CIN(\mult_26/ab[10][0] ), .IN0(
        \mult_26/CARRYB[9][0] ), .IN1(\mult_26/SUMB[9][1] ), .COUT(
        \mult_26/CARRYB[10][0] ), .SUM(o[10]) );
  FADDER \mult_26/S3_11_30  ( .CIN(\mult_26/ab[11][30] ), .IN0(
        \mult_26/CARRYB[10][30] ), .IN1(\mult_26/ab[10][31] ), .COUT(
        \mult_26/CARRYB[11][30] ), .SUM(\mult_26/SUMB[11][30] ) );
  FADDER \mult_26/S2_11_29  ( .CIN(\mult_26/ab[11][29] ), .IN0(
        \mult_26/CARRYB[10][29] ), .IN1(\mult_26/SUMB[10][30] ), .COUT(
        \mult_26/CARRYB[11][29] ), .SUM(\mult_26/SUMB[11][29] ) );
  FADDER \mult_26/S2_11_28  ( .CIN(\mult_26/ab[11][28] ), .IN0(
        \mult_26/CARRYB[10][28] ), .IN1(\mult_26/SUMB[10][29] ), .COUT(
        \mult_26/CARRYB[11][28] ), .SUM(\mult_26/SUMB[11][28] ) );
  FADDER \mult_26/S2_11_27  ( .CIN(\mult_26/ab[11][27] ), .IN0(
        \mult_26/CARRYB[10][27] ), .IN1(\mult_26/SUMB[10][28] ), .COUT(
        \mult_26/CARRYB[11][27] ), .SUM(\mult_26/SUMB[11][27] ) );
  FADDER \mult_26/S2_11_26  ( .CIN(\mult_26/ab[11][26] ), .IN0(
        \mult_26/CARRYB[10][26] ), .IN1(\mult_26/SUMB[10][27] ), .COUT(
        \mult_26/CARRYB[11][26] ), .SUM(\mult_26/SUMB[11][26] ) );
  FADDER \mult_26/S2_11_25  ( .CIN(\mult_26/ab[11][25] ), .IN0(
        \mult_26/CARRYB[10][25] ), .IN1(\mult_26/SUMB[10][26] ), .COUT(
        \mult_26/CARRYB[11][25] ), .SUM(\mult_26/SUMB[11][25] ) );
  FADDER \mult_26/S2_11_24  ( .CIN(\mult_26/ab[11][24] ), .IN0(
        \mult_26/CARRYB[10][24] ), .IN1(\mult_26/SUMB[10][25] ), .COUT(
        \mult_26/CARRYB[11][24] ), .SUM(\mult_26/SUMB[11][24] ) );
  FADDER \mult_26/S2_11_23  ( .CIN(\mult_26/ab[11][23] ), .IN0(
        \mult_26/CARRYB[10][23] ), .IN1(\mult_26/SUMB[10][24] ), .COUT(
        \mult_26/CARRYB[11][23] ), .SUM(\mult_26/SUMB[11][23] ) );
  FADDER \mult_26/S2_11_22  ( .CIN(\mult_26/ab[11][22] ), .IN0(
        \mult_26/CARRYB[10][22] ), .IN1(\mult_26/SUMB[10][23] ), .COUT(
        \mult_26/CARRYB[11][22] ), .SUM(\mult_26/SUMB[11][22] ) );
  FADDER \mult_26/S2_11_21  ( .CIN(\mult_26/ab[11][21] ), .IN0(
        \mult_26/CARRYB[10][21] ), .IN1(\mult_26/SUMB[10][22] ), .COUT(
        \mult_26/CARRYB[11][21] ), .SUM(\mult_26/SUMB[11][21] ) );
  FADDER \mult_26/S2_11_20  ( .CIN(\mult_26/ab[11][20] ), .IN0(
        \mult_26/CARRYB[10][20] ), .IN1(\mult_26/SUMB[10][21] ), .COUT(
        \mult_26/CARRYB[11][20] ), .SUM(\mult_26/SUMB[11][20] ) );
  FADDER \mult_26/S2_11_19  ( .CIN(\mult_26/ab[11][19] ), .IN0(
        \mult_26/CARRYB[10][19] ), .IN1(\mult_26/SUMB[10][20] ), .COUT(
        \mult_26/CARRYB[11][19] ), .SUM(\mult_26/SUMB[11][19] ) );
  FADDER \mult_26/S2_11_18  ( .CIN(\mult_26/ab[11][18] ), .IN0(
        \mult_26/CARRYB[10][18] ), .IN1(\mult_26/SUMB[10][19] ), .COUT(
        \mult_26/CARRYB[11][18] ), .SUM(\mult_26/SUMB[11][18] ) );
  FADDER \mult_26/S2_11_17  ( .CIN(\mult_26/ab[11][17] ), .IN0(
        \mult_26/CARRYB[10][17] ), .IN1(\mult_26/SUMB[10][18] ), .COUT(
        \mult_26/CARRYB[11][17] ), .SUM(\mult_26/SUMB[11][17] ) );
  FADDER \mult_26/S2_11_16  ( .CIN(\mult_26/ab[11][16] ), .IN0(
        \mult_26/CARRYB[10][16] ), .IN1(\mult_26/SUMB[10][17] ), .COUT(
        \mult_26/CARRYB[11][16] ), .SUM(\mult_26/SUMB[11][16] ) );
  FADDER \mult_26/S2_11_15  ( .CIN(\mult_26/ab[11][15] ), .IN0(
        \mult_26/CARRYB[10][15] ), .IN1(\mult_26/SUMB[10][16] ), .COUT(
        \mult_26/CARRYB[11][15] ), .SUM(\mult_26/SUMB[11][15] ) );
  FADDER \mult_26/S2_11_14  ( .CIN(\mult_26/ab[11][14] ), .IN0(
        \mult_26/CARRYB[10][14] ), .IN1(\mult_26/SUMB[10][15] ), .COUT(
        \mult_26/CARRYB[11][14] ), .SUM(\mult_26/SUMB[11][14] ) );
  FADDER \mult_26/S2_11_13  ( .CIN(\mult_26/ab[11][13] ), .IN0(
        \mult_26/CARRYB[10][13] ), .IN1(\mult_26/SUMB[10][14] ), .COUT(
        \mult_26/CARRYB[11][13] ), .SUM(\mult_26/SUMB[11][13] ) );
  FADDER \mult_26/S2_11_12  ( .CIN(\mult_26/ab[11][12] ), .IN0(
        \mult_26/CARRYB[10][12] ), .IN1(\mult_26/SUMB[10][13] ), .COUT(
        \mult_26/CARRYB[11][12] ), .SUM(\mult_26/SUMB[11][12] ) );
  FADDER \mult_26/S2_11_11  ( .CIN(\mult_26/ab[11][11] ), .IN0(
        \mult_26/CARRYB[10][11] ), .IN1(\mult_26/SUMB[10][12] ), .COUT(
        \mult_26/CARRYB[11][11] ), .SUM(\mult_26/SUMB[11][11] ) );
  FADDER \mult_26/S2_11_10  ( .CIN(\mult_26/ab[11][10] ), .IN0(
        \mult_26/CARRYB[10][10] ), .IN1(\mult_26/SUMB[10][11] ), .COUT(
        \mult_26/CARRYB[11][10] ), .SUM(\mult_26/SUMB[11][10] ) );
  FADDER \mult_26/S2_11_9  ( .CIN(\mult_26/ab[11][9] ), .IN0(
        \mult_26/CARRYB[10][9] ), .IN1(\mult_26/SUMB[10][10] ), .COUT(
        \mult_26/CARRYB[11][9] ), .SUM(\mult_26/SUMB[11][9] ) );
  FADDER \mult_26/S2_11_8  ( .CIN(\mult_26/ab[11][8] ), .IN0(
        \mult_26/CARRYB[10][8] ), .IN1(\mult_26/SUMB[10][9] ), .COUT(
        \mult_26/CARRYB[11][8] ), .SUM(\mult_26/SUMB[11][8] ) );
  FADDER \mult_26/S2_11_7  ( .CIN(\mult_26/ab[11][7] ), .IN0(
        \mult_26/CARRYB[10][7] ), .IN1(\mult_26/SUMB[10][8] ), .COUT(
        \mult_26/CARRYB[11][7] ), .SUM(\mult_26/SUMB[11][7] ) );
  FADDER \mult_26/S2_11_6  ( .CIN(\mult_26/ab[11][6] ), .IN0(
        \mult_26/CARRYB[10][6] ), .IN1(\mult_26/SUMB[10][7] ), .COUT(
        \mult_26/CARRYB[11][6] ), .SUM(\mult_26/SUMB[11][6] ) );
  FADDER \mult_26/S2_11_5  ( .CIN(\mult_26/ab[11][5] ), .IN0(
        \mult_26/CARRYB[10][5] ), .IN1(\mult_26/SUMB[10][6] ), .COUT(
        \mult_26/CARRYB[11][5] ), .SUM(\mult_26/SUMB[11][5] ) );
  FADDER \mult_26/S2_11_4  ( .CIN(\mult_26/ab[11][4] ), .IN0(
        \mult_26/CARRYB[10][4] ), .IN1(\mult_26/SUMB[10][5] ), .COUT(
        \mult_26/CARRYB[11][4] ), .SUM(\mult_26/SUMB[11][4] ) );
  FADDER \mult_26/S2_11_3  ( .CIN(\mult_26/ab[11][3] ), .IN0(
        \mult_26/CARRYB[10][3] ), .IN1(\mult_26/SUMB[10][4] ), .COUT(
        \mult_26/CARRYB[11][3] ), .SUM(\mult_26/SUMB[11][3] ) );
  FADDER \mult_26/S2_11_2  ( .CIN(\mult_26/ab[11][2] ), .IN0(
        \mult_26/CARRYB[10][2] ), .IN1(\mult_26/SUMB[10][3] ), .COUT(
        \mult_26/CARRYB[11][2] ), .SUM(\mult_26/SUMB[11][2] ) );
  FADDER \mult_26/S2_11_1  ( .CIN(\mult_26/ab[11][1] ), .IN0(
        \mult_26/CARRYB[10][1] ), .IN1(\mult_26/SUMB[10][2] ), .COUT(
        \mult_26/CARRYB[11][1] ), .SUM(\mult_26/SUMB[11][1] ) );
  FADDER \mult_26/S1_11_0  ( .CIN(\mult_26/ab[11][0] ), .IN0(
        \mult_26/CARRYB[10][0] ), .IN1(\mult_26/SUMB[10][1] ), .COUT(
        \mult_26/CARRYB[11][0] ), .SUM(o[11]) );
  FADDER \mult_26/S3_12_30  ( .CIN(\mult_26/ab[12][30] ), .IN0(
        \mult_26/CARRYB[11][30] ), .IN1(\mult_26/ab[11][31] ), .COUT(
        \mult_26/CARRYB[12][30] ), .SUM(\mult_26/SUMB[12][30] ) );
  FADDER \mult_26/S2_12_29  ( .CIN(\mult_26/ab[12][29] ), .IN0(
        \mult_26/CARRYB[11][29] ), .IN1(\mult_26/SUMB[11][30] ), .COUT(
        \mult_26/CARRYB[12][29] ), .SUM(\mult_26/SUMB[12][29] ) );
  FADDER \mult_26/S2_12_28  ( .CIN(\mult_26/ab[12][28] ), .IN0(
        \mult_26/CARRYB[11][28] ), .IN1(\mult_26/SUMB[11][29] ), .COUT(
        \mult_26/CARRYB[12][28] ), .SUM(\mult_26/SUMB[12][28] ) );
  FADDER \mult_26/S2_12_27  ( .CIN(\mult_26/ab[12][27] ), .IN0(
        \mult_26/CARRYB[11][27] ), .IN1(\mult_26/SUMB[11][28] ), .COUT(
        \mult_26/CARRYB[12][27] ), .SUM(\mult_26/SUMB[12][27] ) );
  FADDER \mult_26/S2_12_26  ( .CIN(\mult_26/ab[12][26] ), .IN0(
        \mult_26/CARRYB[11][26] ), .IN1(\mult_26/SUMB[11][27] ), .COUT(
        \mult_26/CARRYB[12][26] ), .SUM(\mult_26/SUMB[12][26] ) );
  FADDER \mult_26/S2_12_25  ( .CIN(\mult_26/ab[12][25] ), .IN0(
        \mult_26/CARRYB[11][25] ), .IN1(\mult_26/SUMB[11][26] ), .COUT(
        \mult_26/CARRYB[12][25] ), .SUM(\mult_26/SUMB[12][25] ) );
  FADDER \mult_26/S2_12_24  ( .CIN(\mult_26/ab[12][24] ), .IN0(
        \mult_26/CARRYB[11][24] ), .IN1(\mult_26/SUMB[11][25] ), .COUT(
        \mult_26/CARRYB[12][24] ), .SUM(\mult_26/SUMB[12][24] ) );
  FADDER \mult_26/S2_12_23  ( .CIN(\mult_26/ab[12][23] ), .IN0(
        \mult_26/CARRYB[11][23] ), .IN1(\mult_26/SUMB[11][24] ), .COUT(
        \mult_26/CARRYB[12][23] ), .SUM(\mult_26/SUMB[12][23] ) );
  FADDER \mult_26/S2_12_22  ( .CIN(\mult_26/ab[12][22] ), .IN0(
        \mult_26/CARRYB[11][22] ), .IN1(\mult_26/SUMB[11][23] ), .COUT(
        \mult_26/CARRYB[12][22] ), .SUM(\mult_26/SUMB[12][22] ) );
  FADDER \mult_26/S2_12_21  ( .CIN(\mult_26/ab[12][21] ), .IN0(
        \mult_26/CARRYB[11][21] ), .IN1(\mult_26/SUMB[11][22] ), .COUT(
        \mult_26/CARRYB[12][21] ), .SUM(\mult_26/SUMB[12][21] ) );
  FADDER \mult_26/S2_12_20  ( .CIN(\mult_26/ab[12][20] ), .IN0(
        \mult_26/CARRYB[11][20] ), .IN1(\mult_26/SUMB[11][21] ), .COUT(
        \mult_26/CARRYB[12][20] ), .SUM(\mult_26/SUMB[12][20] ) );
  FADDER \mult_26/S2_12_19  ( .CIN(\mult_26/ab[12][19] ), .IN0(
        \mult_26/CARRYB[11][19] ), .IN1(\mult_26/SUMB[11][20] ), .COUT(
        \mult_26/CARRYB[12][19] ), .SUM(\mult_26/SUMB[12][19] ) );
  FADDER \mult_26/S2_12_18  ( .CIN(\mult_26/ab[12][18] ), .IN0(
        \mult_26/CARRYB[11][18] ), .IN1(\mult_26/SUMB[11][19] ), .COUT(
        \mult_26/CARRYB[12][18] ), .SUM(\mult_26/SUMB[12][18] ) );
  FADDER \mult_26/S2_12_17  ( .CIN(\mult_26/ab[12][17] ), .IN0(
        \mult_26/CARRYB[11][17] ), .IN1(\mult_26/SUMB[11][18] ), .COUT(
        \mult_26/CARRYB[12][17] ), .SUM(\mult_26/SUMB[12][17] ) );
  FADDER \mult_26/S2_12_16  ( .CIN(\mult_26/ab[12][16] ), .IN0(
        \mult_26/CARRYB[11][16] ), .IN1(\mult_26/SUMB[11][17] ), .COUT(
        \mult_26/CARRYB[12][16] ), .SUM(\mult_26/SUMB[12][16] ) );
  FADDER \mult_26/S2_12_15  ( .CIN(\mult_26/ab[12][15] ), .IN0(
        \mult_26/CARRYB[11][15] ), .IN1(\mult_26/SUMB[11][16] ), .COUT(
        \mult_26/CARRYB[12][15] ), .SUM(\mult_26/SUMB[12][15] ) );
  FADDER \mult_26/S2_12_14  ( .CIN(\mult_26/ab[12][14] ), .IN0(
        \mult_26/CARRYB[11][14] ), .IN1(\mult_26/SUMB[11][15] ), .COUT(
        \mult_26/CARRYB[12][14] ), .SUM(\mult_26/SUMB[12][14] ) );
  FADDER \mult_26/S2_12_13  ( .CIN(\mult_26/ab[12][13] ), .IN0(
        \mult_26/CARRYB[11][13] ), .IN1(\mult_26/SUMB[11][14] ), .COUT(
        \mult_26/CARRYB[12][13] ), .SUM(\mult_26/SUMB[12][13] ) );
  FADDER \mult_26/S2_12_12  ( .CIN(\mult_26/ab[12][12] ), .IN0(
        \mult_26/CARRYB[11][12] ), .IN1(\mult_26/SUMB[11][13] ), .COUT(
        \mult_26/CARRYB[12][12] ), .SUM(\mult_26/SUMB[12][12] ) );
  FADDER \mult_26/S2_12_11  ( .CIN(\mult_26/ab[12][11] ), .IN0(
        \mult_26/CARRYB[11][11] ), .IN1(\mult_26/SUMB[11][12] ), .COUT(
        \mult_26/CARRYB[12][11] ), .SUM(\mult_26/SUMB[12][11] ) );
  FADDER \mult_26/S2_12_10  ( .CIN(\mult_26/ab[12][10] ), .IN0(
        \mult_26/CARRYB[11][10] ), .IN1(\mult_26/SUMB[11][11] ), .COUT(
        \mult_26/CARRYB[12][10] ), .SUM(\mult_26/SUMB[12][10] ) );
  FADDER \mult_26/S2_12_9  ( .CIN(\mult_26/ab[12][9] ), .IN0(
        \mult_26/CARRYB[11][9] ), .IN1(\mult_26/SUMB[11][10] ), .COUT(
        \mult_26/CARRYB[12][9] ), .SUM(\mult_26/SUMB[12][9] ) );
  FADDER \mult_26/S2_12_8  ( .CIN(\mult_26/ab[12][8] ), .IN0(
        \mult_26/CARRYB[11][8] ), .IN1(\mult_26/SUMB[11][9] ), .COUT(
        \mult_26/CARRYB[12][8] ), .SUM(\mult_26/SUMB[12][8] ) );
  FADDER \mult_26/S2_12_7  ( .CIN(\mult_26/ab[12][7] ), .IN0(
        \mult_26/CARRYB[11][7] ), .IN1(\mult_26/SUMB[11][8] ), .COUT(
        \mult_26/CARRYB[12][7] ), .SUM(\mult_26/SUMB[12][7] ) );
  FADDER \mult_26/S2_12_6  ( .CIN(\mult_26/ab[12][6] ), .IN0(
        \mult_26/CARRYB[11][6] ), .IN1(\mult_26/SUMB[11][7] ), .COUT(
        \mult_26/CARRYB[12][6] ), .SUM(\mult_26/SUMB[12][6] ) );
  FADDER \mult_26/S2_12_5  ( .CIN(\mult_26/ab[12][5] ), .IN0(
        \mult_26/CARRYB[11][5] ), .IN1(\mult_26/SUMB[11][6] ), .COUT(
        \mult_26/CARRYB[12][5] ), .SUM(\mult_26/SUMB[12][5] ) );
  FADDER \mult_26/S2_12_4  ( .CIN(\mult_26/ab[12][4] ), .IN0(
        \mult_26/CARRYB[11][4] ), .IN1(\mult_26/SUMB[11][5] ), .COUT(
        \mult_26/CARRYB[12][4] ), .SUM(\mult_26/SUMB[12][4] ) );
  FADDER \mult_26/S2_12_3  ( .CIN(\mult_26/ab[12][3] ), .IN0(
        \mult_26/CARRYB[11][3] ), .IN1(\mult_26/SUMB[11][4] ), .COUT(
        \mult_26/CARRYB[12][3] ), .SUM(\mult_26/SUMB[12][3] ) );
  FADDER \mult_26/S2_12_2  ( .CIN(\mult_26/ab[12][2] ), .IN0(
        \mult_26/CARRYB[11][2] ), .IN1(\mult_26/SUMB[11][3] ), .COUT(
        \mult_26/CARRYB[12][2] ), .SUM(\mult_26/SUMB[12][2] ) );
  FADDER \mult_26/S2_12_1  ( .CIN(\mult_26/ab[12][1] ), .IN0(
        \mult_26/CARRYB[11][1] ), .IN1(\mult_26/SUMB[11][2] ), .COUT(
        \mult_26/CARRYB[12][1] ), .SUM(\mult_26/SUMB[12][1] ) );
  FADDER \mult_26/S1_12_0  ( .CIN(\mult_26/ab[12][0] ), .IN0(
        \mult_26/CARRYB[11][0] ), .IN1(\mult_26/SUMB[11][1] ), .COUT(
        \mult_26/CARRYB[12][0] ), .SUM(o[12]) );
  FADDER \mult_26/S3_13_30  ( .CIN(\mult_26/ab[13][30] ), .IN0(
        \mult_26/CARRYB[12][30] ), .IN1(\mult_26/ab[12][31] ), .COUT(
        \mult_26/CARRYB[13][30] ), .SUM(\mult_26/SUMB[13][30] ) );
  FADDER \mult_26/S2_13_29  ( .CIN(\mult_26/ab[13][29] ), .IN0(
        \mult_26/CARRYB[12][29] ), .IN1(\mult_26/SUMB[12][30] ), .COUT(
        \mult_26/CARRYB[13][29] ), .SUM(\mult_26/SUMB[13][29] ) );
  FADDER \mult_26/S2_13_28  ( .CIN(\mult_26/ab[13][28] ), .IN0(
        \mult_26/CARRYB[12][28] ), .IN1(\mult_26/SUMB[12][29] ), .COUT(
        \mult_26/CARRYB[13][28] ), .SUM(\mult_26/SUMB[13][28] ) );
  FADDER \mult_26/S2_13_27  ( .CIN(\mult_26/ab[13][27] ), .IN0(
        \mult_26/CARRYB[12][27] ), .IN1(\mult_26/SUMB[12][28] ), .COUT(
        \mult_26/CARRYB[13][27] ), .SUM(\mult_26/SUMB[13][27] ) );
  FADDER \mult_26/S2_13_26  ( .CIN(\mult_26/ab[13][26] ), .IN0(
        \mult_26/CARRYB[12][26] ), .IN1(\mult_26/SUMB[12][27] ), .COUT(
        \mult_26/CARRYB[13][26] ), .SUM(\mult_26/SUMB[13][26] ) );
  FADDER \mult_26/S2_13_25  ( .CIN(\mult_26/ab[13][25] ), .IN0(
        \mult_26/CARRYB[12][25] ), .IN1(\mult_26/SUMB[12][26] ), .COUT(
        \mult_26/CARRYB[13][25] ), .SUM(\mult_26/SUMB[13][25] ) );
  FADDER \mult_26/S2_13_24  ( .CIN(\mult_26/ab[13][24] ), .IN0(
        \mult_26/CARRYB[12][24] ), .IN1(\mult_26/SUMB[12][25] ), .COUT(
        \mult_26/CARRYB[13][24] ), .SUM(\mult_26/SUMB[13][24] ) );
  FADDER \mult_26/S2_13_23  ( .CIN(\mult_26/ab[13][23] ), .IN0(
        \mult_26/CARRYB[12][23] ), .IN1(\mult_26/SUMB[12][24] ), .COUT(
        \mult_26/CARRYB[13][23] ), .SUM(\mult_26/SUMB[13][23] ) );
  FADDER \mult_26/S2_13_22  ( .CIN(\mult_26/ab[13][22] ), .IN0(
        \mult_26/CARRYB[12][22] ), .IN1(\mult_26/SUMB[12][23] ), .COUT(
        \mult_26/CARRYB[13][22] ), .SUM(\mult_26/SUMB[13][22] ) );
  FADDER \mult_26/S2_13_21  ( .CIN(\mult_26/ab[13][21] ), .IN0(
        \mult_26/CARRYB[12][21] ), .IN1(\mult_26/SUMB[12][22] ), .COUT(
        \mult_26/CARRYB[13][21] ), .SUM(\mult_26/SUMB[13][21] ) );
  FADDER \mult_26/S2_13_20  ( .CIN(\mult_26/ab[13][20] ), .IN0(
        \mult_26/CARRYB[12][20] ), .IN1(\mult_26/SUMB[12][21] ), .COUT(
        \mult_26/CARRYB[13][20] ), .SUM(\mult_26/SUMB[13][20] ) );
  FADDER \mult_26/S2_13_19  ( .CIN(\mult_26/ab[13][19] ), .IN0(
        \mult_26/CARRYB[12][19] ), .IN1(\mult_26/SUMB[12][20] ), .COUT(
        \mult_26/CARRYB[13][19] ), .SUM(\mult_26/SUMB[13][19] ) );
  FADDER \mult_26/S2_13_18  ( .CIN(\mult_26/ab[13][18] ), .IN0(
        \mult_26/CARRYB[12][18] ), .IN1(\mult_26/SUMB[12][19] ), .COUT(
        \mult_26/CARRYB[13][18] ), .SUM(\mult_26/SUMB[13][18] ) );
  FADDER \mult_26/S2_13_17  ( .CIN(\mult_26/ab[13][17] ), .IN0(
        \mult_26/CARRYB[12][17] ), .IN1(\mult_26/SUMB[12][18] ), .COUT(
        \mult_26/CARRYB[13][17] ), .SUM(\mult_26/SUMB[13][17] ) );
  FADDER \mult_26/S2_13_16  ( .CIN(\mult_26/ab[13][16] ), .IN0(
        \mult_26/CARRYB[12][16] ), .IN1(\mult_26/SUMB[12][17] ), .COUT(
        \mult_26/CARRYB[13][16] ), .SUM(\mult_26/SUMB[13][16] ) );
  FADDER \mult_26/S2_13_15  ( .CIN(\mult_26/ab[13][15] ), .IN0(
        \mult_26/CARRYB[12][15] ), .IN1(\mult_26/SUMB[12][16] ), .COUT(
        \mult_26/CARRYB[13][15] ), .SUM(\mult_26/SUMB[13][15] ) );
  FADDER \mult_26/S2_13_14  ( .CIN(\mult_26/ab[13][14] ), .IN0(
        \mult_26/CARRYB[12][14] ), .IN1(\mult_26/SUMB[12][15] ), .COUT(
        \mult_26/CARRYB[13][14] ), .SUM(\mult_26/SUMB[13][14] ) );
  FADDER \mult_26/S2_13_13  ( .CIN(\mult_26/ab[13][13] ), .IN0(
        \mult_26/CARRYB[12][13] ), .IN1(\mult_26/SUMB[12][14] ), .COUT(
        \mult_26/CARRYB[13][13] ), .SUM(\mult_26/SUMB[13][13] ) );
  FADDER \mult_26/S2_13_12  ( .CIN(\mult_26/ab[13][12] ), .IN0(
        \mult_26/CARRYB[12][12] ), .IN1(\mult_26/SUMB[12][13] ), .COUT(
        \mult_26/CARRYB[13][12] ), .SUM(\mult_26/SUMB[13][12] ) );
  FADDER \mult_26/S2_13_11  ( .CIN(\mult_26/ab[13][11] ), .IN0(
        \mult_26/CARRYB[12][11] ), .IN1(\mult_26/SUMB[12][12] ), .COUT(
        \mult_26/CARRYB[13][11] ), .SUM(\mult_26/SUMB[13][11] ) );
  FADDER \mult_26/S2_13_10  ( .CIN(\mult_26/ab[13][10] ), .IN0(
        \mult_26/CARRYB[12][10] ), .IN1(\mult_26/SUMB[12][11] ), .COUT(
        \mult_26/CARRYB[13][10] ), .SUM(\mult_26/SUMB[13][10] ) );
  FADDER \mult_26/S2_13_9  ( .CIN(\mult_26/ab[13][9] ), .IN0(
        \mult_26/CARRYB[12][9] ), .IN1(\mult_26/SUMB[12][10] ), .COUT(
        \mult_26/CARRYB[13][9] ), .SUM(\mult_26/SUMB[13][9] ) );
  FADDER \mult_26/S2_13_8  ( .CIN(\mult_26/ab[13][8] ), .IN0(
        \mult_26/CARRYB[12][8] ), .IN1(\mult_26/SUMB[12][9] ), .COUT(
        \mult_26/CARRYB[13][8] ), .SUM(\mult_26/SUMB[13][8] ) );
  FADDER \mult_26/S2_13_7  ( .CIN(\mult_26/ab[13][7] ), .IN0(
        \mult_26/CARRYB[12][7] ), .IN1(\mult_26/SUMB[12][8] ), .COUT(
        \mult_26/CARRYB[13][7] ), .SUM(\mult_26/SUMB[13][7] ) );
  FADDER \mult_26/S2_13_6  ( .CIN(\mult_26/ab[13][6] ), .IN0(
        \mult_26/CARRYB[12][6] ), .IN1(\mult_26/SUMB[12][7] ), .COUT(
        \mult_26/CARRYB[13][6] ), .SUM(\mult_26/SUMB[13][6] ) );
  FADDER \mult_26/S2_13_5  ( .CIN(\mult_26/ab[13][5] ), .IN0(
        \mult_26/CARRYB[12][5] ), .IN1(\mult_26/SUMB[12][6] ), .COUT(
        \mult_26/CARRYB[13][5] ), .SUM(\mult_26/SUMB[13][5] ) );
  FADDER \mult_26/S2_13_4  ( .CIN(\mult_26/ab[13][4] ), .IN0(
        \mult_26/CARRYB[12][4] ), .IN1(\mult_26/SUMB[12][5] ), .COUT(
        \mult_26/CARRYB[13][4] ), .SUM(\mult_26/SUMB[13][4] ) );
  FADDER \mult_26/S2_13_3  ( .CIN(\mult_26/ab[13][3] ), .IN0(
        \mult_26/CARRYB[12][3] ), .IN1(\mult_26/SUMB[12][4] ), .COUT(
        \mult_26/CARRYB[13][3] ), .SUM(\mult_26/SUMB[13][3] ) );
  FADDER \mult_26/S2_13_2  ( .CIN(\mult_26/ab[13][2] ), .IN0(
        \mult_26/CARRYB[12][2] ), .IN1(\mult_26/SUMB[12][3] ), .COUT(
        \mult_26/CARRYB[13][2] ), .SUM(\mult_26/SUMB[13][2] ) );
  FADDER \mult_26/S2_13_1  ( .CIN(\mult_26/ab[13][1] ), .IN0(
        \mult_26/CARRYB[12][1] ), .IN1(\mult_26/SUMB[12][2] ), .COUT(
        \mult_26/CARRYB[13][1] ), .SUM(\mult_26/SUMB[13][1] ) );
  FADDER \mult_26/S1_13_0  ( .CIN(\mult_26/ab[13][0] ), .IN0(
        \mult_26/CARRYB[12][0] ), .IN1(\mult_26/SUMB[12][1] ), .COUT(
        \mult_26/CARRYB[13][0] ), .SUM(o[13]) );
  FADDER \mult_26/S3_14_30  ( .CIN(\mult_26/ab[14][30] ), .IN0(
        \mult_26/CARRYB[13][30] ), .IN1(\mult_26/ab[13][31] ), .COUT(
        \mult_26/CARRYB[14][30] ), .SUM(\mult_26/SUMB[14][30] ) );
  FADDER \mult_26/S2_14_29  ( .CIN(\mult_26/ab[14][29] ), .IN0(
        \mult_26/CARRYB[13][29] ), .IN1(\mult_26/SUMB[13][30] ), .COUT(
        \mult_26/CARRYB[14][29] ), .SUM(\mult_26/SUMB[14][29] ) );
  FADDER \mult_26/S2_14_28  ( .CIN(\mult_26/ab[14][28] ), .IN0(
        \mult_26/CARRYB[13][28] ), .IN1(\mult_26/SUMB[13][29] ), .COUT(
        \mult_26/CARRYB[14][28] ), .SUM(\mult_26/SUMB[14][28] ) );
  FADDER \mult_26/S2_14_27  ( .CIN(\mult_26/ab[14][27] ), .IN0(
        \mult_26/CARRYB[13][27] ), .IN1(\mult_26/SUMB[13][28] ), .COUT(
        \mult_26/CARRYB[14][27] ), .SUM(\mult_26/SUMB[14][27] ) );
  FADDER \mult_26/S2_14_26  ( .CIN(\mult_26/ab[14][26] ), .IN0(
        \mult_26/CARRYB[13][26] ), .IN1(\mult_26/SUMB[13][27] ), .COUT(
        \mult_26/CARRYB[14][26] ), .SUM(\mult_26/SUMB[14][26] ) );
  FADDER \mult_26/S2_14_25  ( .CIN(\mult_26/ab[14][25] ), .IN0(
        \mult_26/CARRYB[13][25] ), .IN1(\mult_26/SUMB[13][26] ), .COUT(
        \mult_26/CARRYB[14][25] ), .SUM(\mult_26/SUMB[14][25] ) );
  FADDER \mult_26/S2_14_24  ( .CIN(\mult_26/ab[14][24] ), .IN0(
        \mult_26/CARRYB[13][24] ), .IN1(\mult_26/SUMB[13][25] ), .COUT(
        \mult_26/CARRYB[14][24] ), .SUM(\mult_26/SUMB[14][24] ) );
  FADDER \mult_26/S2_14_23  ( .CIN(\mult_26/ab[14][23] ), .IN0(
        \mult_26/CARRYB[13][23] ), .IN1(\mult_26/SUMB[13][24] ), .COUT(
        \mult_26/CARRYB[14][23] ), .SUM(\mult_26/SUMB[14][23] ) );
  FADDER \mult_26/S2_14_22  ( .CIN(\mult_26/ab[14][22] ), .IN0(
        \mult_26/CARRYB[13][22] ), .IN1(\mult_26/SUMB[13][23] ), .COUT(
        \mult_26/CARRYB[14][22] ), .SUM(\mult_26/SUMB[14][22] ) );
  FADDER \mult_26/S2_14_21  ( .CIN(\mult_26/ab[14][21] ), .IN0(
        \mult_26/CARRYB[13][21] ), .IN1(\mult_26/SUMB[13][22] ), .COUT(
        \mult_26/CARRYB[14][21] ), .SUM(\mult_26/SUMB[14][21] ) );
  FADDER \mult_26/S2_14_20  ( .CIN(\mult_26/ab[14][20] ), .IN0(
        \mult_26/CARRYB[13][20] ), .IN1(\mult_26/SUMB[13][21] ), .COUT(
        \mult_26/CARRYB[14][20] ), .SUM(\mult_26/SUMB[14][20] ) );
  FADDER \mult_26/S2_14_19  ( .CIN(\mult_26/ab[14][19] ), .IN0(
        \mult_26/CARRYB[13][19] ), .IN1(\mult_26/SUMB[13][20] ), .COUT(
        \mult_26/CARRYB[14][19] ), .SUM(\mult_26/SUMB[14][19] ) );
  FADDER \mult_26/S2_14_18  ( .CIN(\mult_26/ab[14][18] ), .IN0(
        \mult_26/CARRYB[13][18] ), .IN1(\mult_26/SUMB[13][19] ), .COUT(
        \mult_26/CARRYB[14][18] ), .SUM(\mult_26/SUMB[14][18] ) );
  FADDER \mult_26/S2_14_17  ( .CIN(\mult_26/ab[14][17] ), .IN0(
        \mult_26/CARRYB[13][17] ), .IN1(\mult_26/SUMB[13][18] ), .COUT(
        \mult_26/CARRYB[14][17] ), .SUM(\mult_26/SUMB[14][17] ) );
  FADDER \mult_26/S2_14_16  ( .CIN(\mult_26/ab[14][16] ), .IN0(
        \mult_26/CARRYB[13][16] ), .IN1(\mult_26/SUMB[13][17] ), .COUT(
        \mult_26/CARRYB[14][16] ), .SUM(\mult_26/SUMB[14][16] ) );
  FADDER \mult_26/S2_14_15  ( .CIN(\mult_26/ab[14][15] ), .IN0(
        \mult_26/CARRYB[13][15] ), .IN1(\mult_26/SUMB[13][16] ), .COUT(
        \mult_26/CARRYB[14][15] ), .SUM(\mult_26/SUMB[14][15] ) );
  FADDER \mult_26/S2_14_14  ( .CIN(\mult_26/ab[14][14] ), .IN0(
        \mult_26/CARRYB[13][14] ), .IN1(\mult_26/SUMB[13][15] ), .COUT(
        \mult_26/CARRYB[14][14] ), .SUM(\mult_26/SUMB[14][14] ) );
  FADDER \mult_26/S2_14_13  ( .CIN(\mult_26/ab[14][13] ), .IN0(
        \mult_26/CARRYB[13][13] ), .IN1(\mult_26/SUMB[13][14] ), .COUT(
        \mult_26/CARRYB[14][13] ), .SUM(\mult_26/SUMB[14][13] ) );
  FADDER \mult_26/S2_14_12  ( .CIN(\mult_26/ab[14][12] ), .IN0(
        \mult_26/CARRYB[13][12] ), .IN1(\mult_26/SUMB[13][13] ), .COUT(
        \mult_26/CARRYB[14][12] ), .SUM(\mult_26/SUMB[14][12] ) );
  FADDER \mult_26/S2_14_11  ( .CIN(\mult_26/ab[14][11] ), .IN0(
        \mult_26/CARRYB[13][11] ), .IN1(\mult_26/SUMB[13][12] ), .COUT(
        \mult_26/CARRYB[14][11] ), .SUM(\mult_26/SUMB[14][11] ) );
  FADDER \mult_26/S2_14_10  ( .CIN(\mult_26/ab[14][10] ), .IN0(
        \mult_26/CARRYB[13][10] ), .IN1(\mult_26/SUMB[13][11] ), .COUT(
        \mult_26/CARRYB[14][10] ), .SUM(\mult_26/SUMB[14][10] ) );
  FADDER \mult_26/S2_14_9  ( .CIN(\mult_26/ab[14][9] ), .IN0(
        \mult_26/CARRYB[13][9] ), .IN1(\mult_26/SUMB[13][10] ), .COUT(
        \mult_26/CARRYB[14][9] ), .SUM(\mult_26/SUMB[14][9] ) );
  FADDER \mult_26/S2_14_8  ( .CIN(\mult_26/ab[14][8] ), .IN0(
        \mult_26/CARRYB[13][8] ), .IN1(\mult_26/SUMB[13][9] ), .COUT(
        \mult_26/CARRYB[14][8] ), .SUM(\mult_26/SUMB[14][8] ) );
  FADDER \mult_26/S2_14_7  ( .CIN(\mult_26/ab[14][7] ), .IN0(
        \mult_26/CARRYB[13][7] ), .IN1(\mult_26/SUMB[13][8] ), .COUT(
        \mult_26/CARRYB[14][7] ), .SUM(\mult_26/SUMB[14][7] ) );
  FADDER \mult_26/S2_14_6  ( .CIN(\mult_26/ab[14][6] ), .IN0(
        \mult_26/CARRYB[13][6] ), .IN1(\mult_26/SUMB[13][7] ), .COUT(
        \mult_26/CARRYB[14][6] ), .SUM(\mult_26/SUMB[14][6] ) );
  FADDER \mult_26/S2_14_5  ( .CIN(\mult_26/ab[14][5] ), .IN0(
        \mult_26/CARRYB[13][5] ), .IN1(\mult_26/SUMB[13][6] ), .COUT(
        \mult_26/CARRYB[14][5] ), .SUM(\mult_26/SUMB[14][5] ) );
  FADDER \mult_26/S2_14_4  ( .CIN(\mult_26/ab[14][4] ), .IN0(
        \mult_26/CARRYB[13][4] ), .IN1(\mult_26/SUMB[13][5] ), .COUT(
        \mult_26/CARRYB[14][4] ), .SUM(\mult_26/SUMB[14][4] ) );
  FADDER \mult_26/S2_14_3  ( .CIN(\mult_26/ab[14][3] ), .IN0(
        \mult_26/CARRYB[13][3] ), .IN1(\mult_26/SUMB[13][4] ), .COUT(
        \mult_26/CARRYB[14][3] ), .SUM(\mult_26/SUMB[14][3] ) );
  FADDER \mult_26/S2_14_2  ( .CIN(\mult_26/ab[14][2] ), .IN0(
        \mult_26/CARRYB[13][2] ), .IN1(\mult_26/SUMB[13][3] ), .COUT(
        \mult_26/CARRYB[14][2] ), .SUM(\mult_26/SUMB[14][2] ) );
  FADDER \mult_26/S2_14_1  ( .CIN(\mult_26/ab[14][1] ), .IN0(
        \mult_26/CARRYB[13][1] ), .IN1(\mult_26/SUMB[13][2] ), .COUT(
        \mult_26/CARRYB[14][1] ), .SUM(\mult_26/SUMB[14][1] ) );
  FADDER \mult_26/S1_14_0  ( .CIN(\mult_26/ab[14][0] ), .IN0(
        \mult_26/CARRYB[13][0] ), .IN1(\mult_26/SUMB[13][1] ), .COUT(
        \mult_26/CARRYB[14][0] ), .SUM(o[14]) );
  FADDER \mult_26/S3_15_30  ( .CIN(\mult_26/ab[15][30] ), .IN0(
        \mult_26/CARRYB[14][30] ), .IN1(\mult_26/ab[14][31] ), .COUT(
        \mult_26/CARRYB[15][30] ), .SUM(\mult_26/SUMB[15][30] ) );
  FADDER \mult_26/S2_15_29  ( .CIN(\mult_26/ab[15][29] ), .IN0(
        \mult_26/CARRYB[14][29] ), .IN1(\mult_26/SUMB[14][30] ), .COUT(
        \mult_26/CARRYB[15][29] ), .SUM(\mult_26/SUMB[15][29] ) );
  FADDER \mult_26/S2_15_28  ( .CIN(\mult_26/ab[15][28] ), .IN0(
        \mult_26/CARRYB[14][28] ), .IN1(\mult_26/SUMB[14][29] ), .COUT(
        \mult_26/CARRYB[15][28] ), .SUM(\mult_26/SUMB[15][28] ) );
  FADDER \mult_26/S2_15_27  ( .CIN(\mult_26/ab[15][27] ), .IN0(
        \mult_26/CARRYB[14][27] ), .IN1(\mult_26/SUMB[14][28] ), .COUT(
        \mult_26/CARRYB[15][27] ), .SUM(\mult_26/SUMB[15][27] ) );
  FADDER \mult_26/S2_15_26  ( .CIN(\mult_26/ab[15][26] ), .IN0(
        \mult_26/CARRYB[14][26] ), .IN1(\mult_26/SUMB[14][27] ), .COUT(
        \mult_26/CARRYB[15][26] ), .SUM(\mult_26/SUMB[15][26] ) );
  FADDER \mult_26/S2_15_25  ( .CIN(\mult_26/ab[15][25] ), .IN0(
        \mult_26/CARRYB[14][25] ), .IN1(\mult_26/SUMB[14][26] ), .COUT(
        \mult_26/CARRYB[15][25] ), .SUM(\mult_26/SUMB[15][25] ) );
  FADDER \mult_26/S2_15_24  ( .CIN(\mult_26/ab[15][24] ), .IN0(
        \mult_26/CARRYB[14][24] ), .IN1(\mult_26/SUMB[14][25] ), .COUT(
        \mult_26/CARRYB[15][24] ), .SUM(\mult_26/SUMB[15][24] ) );
  FADDER \mult_26/S2_15_23  ( .CIN(\mult_26/ab[15][23] ), .IN0(
        \mult_26/CARRYB[14][23] ), .IN1(\mult_26/SUMB[14][24] ), .COUT(
        \mult_26/CARRYB[15][23] ), .SUM(\mult_26/SUMB[15][23] ) );
  FADDER \mult_26/S2_15_22  ( .CIN(\mult_26/ab[15][22] ), .IN0(
        \mult_26/CARRYB[14][22] ), .IN1(\mult_26/SUMB[14][23] ), .COUT(
        \mult_26/CARRYB[15][22] ), .SUM(\mult_26/SUMB[15][22] ) );
  FADDER \mult_26/S2_15_21  ( .CIN(\mult_26/ab[15][21] ), .IN0(
        \mult_26/CARRYB[14][21] ), .IN1(\mult_26/SUMB[14][22] ), .COUT(
        \mult_26/CARRYB[15][21] ), .SUM(\mult_26/SUMB[15][21] ) );
  FADDER \mult_26/S2_15_20  ( .CIN(\mult_26/ab[15][20] ), .IN0(
        \mult_26/CARRYB[14][20] ), .IN1(\mult_26/SUMB[14][21] ), .COUT(
        \mult_26/CARRYB[15][20] ), .SUM(\mult_26/SUMB[15][20] ) );
  FADDER \mult_26/S2_15_19  ( .CIN(\mult_26/ab[15][19] ), .IN0(
        \mult_26/CARRYB[14][19] ), .IN1(\mult_26/SUMB[14][20] ), .COUT(
        \mult_26/CARRYB[15][19] ), .SUM(\mult_26/SUMB[15][19] ) );
  FADDER \mult_26/S2_15_18  ( .CIN(\mult_26/ab[15][18] ), .IN0(
        \mult_26/CARRYB[14][18] ), .IN1(\mult_26/SUMB[14][19] ), .COUT(
        \mult_26/CARRYB[15][18] ), .SUM(\mult_26/SUMB[15][18] ) );
  FADDER \mult_26/S2_15_17  ( .CIN(\mult_26/ab[15][17] ), .IN0(
        \mult_26/CARRYB[14][17] ), .IN1(\mult_26/SUMB[14][18] ), .COUT(
        \mult_26/CARRYB[15][17] ), .SUM(\mult_26/SUMB[15][17] ) );
  FADDER \mult_26/S2_15_16  ( .CIN(\mult_26/ab[15][16] ), .IN0(
        \mult_26/CARRYB[14][16] ), .IN1(\mult_26/SUMB[14][17] ), .COUT(
        \mult_26/CARRYB[15][16] ), .SUM(\mult_26/SUMB[15][16] ) );
  FADDER \mult_26/S2_15_15  ( .CIN(\mult_26/ab[15][15] ), .IN0(
        \mult_26/CARRYB[14][15] ), .IN1(\mult_26/SUMB[14][16] ), .COUT(
        \mult_26/CARRYB[15][15] ), .SUM(\mult_26/SUMB[15][15] ) );
  FADDER \mult_26/S2_15_14  ( .CIN(\mult_26/ab[15][14] ), .IN0(
        \mult_26/CARRYB[14][14] ), .IN1(\mult_26/SUMB[14][15] ), .COUT(
        \mult_26/CARRYB[15][14] ), .SUM(\mult_26/SUMB[15][14] ) );
  FADDER \mult_26/S2_15_13  ( .CIN(\mult_26/ab[15][13] ), .IN0(
        \mult_26/CARRYB[14][13] ), .IN1(\mult_26/SUMB[14][14] ), .COUT(
        \mult_26/CARRYB[15][13] ), .SUM(\mult_26/SUMB[15][13] ) );
  FADDER \mult_26/S2_15_12  ( .CIN(\mult_26/ab[15][12] ), .IN0(
        \mult_26/CARRYB[14][12] ), .IN1(\mult_26/SUMB[14][13] ), .COUT(
        \mult_26/CARRYB[15][12] ), .SUM(\mult_26/SUMB[15][12] ) );
  FADDER \mult_26/S2_15_11  ( .CIN(\mult_26/ab[15][11] ), .IN0(
        \mult_26/CARRYB[14][11] ), .IN1(\mult_26/SUMB[14][12] ), .COUT(
        \mult_26/CARRYB[15][11] ), .SUM(\mult_26/SUMB[15][11] ) );
  FADDER \mult_26/S2_15_10  ( .CIN(\mult_26/ab[15][10] ), .IN0(
        \mult_26/CARRYB[14][10] ), .IN1(\mult_26/SUMB[14][11] ), .COUT(
        \mult_26/CARRYB[15][10] ), .SUM(\mult_26/SUMB[15][10] ) );
  FADDER \mult_26/S2_15_9  ( .CIN(\mult_26/ab[15][9] ), .IN0(
        \mult_26/CARRYB[14][9] ), .IN1(\mult_26/SUMB[14][10] ), .COUT(
        \mult_26/CARRYB[15][9] ), .SUM(\mult_26/SUMB[15][9] ) );
  FADDER \mult_26/S2_15_8  ( .CIN(\mult_26/ab[15][8] ), .IN0(
        \mult_26/CARRYB[14][8] ), .IN1(\mult_26/SUMB[14][9] ), .COUT(
        \mult_26/CARRYB[15][8] ), .SUM(\mult_26/SUMB[15][8] ) );
  FADDER \mult_26/S2_15_7  ( .CIN(\mult_26/ab[15][7] ), .IN0(
        \mult_26/CARRYB[14][7] ), .IN1(\mult_26/SUMB[14][8] ), .COUT(
        \mult_26/CARRYB[15][7] ), .SUM(\mult_26/SUMB[15][7] ) );
  FADDER \mult_26/S2_15_6  ( .CIN(\mult_26/ab[15][6] ), .IN0(
        \mult_26/CARRYB[14][6] ), .IN1(\mult_26/SUMB[14][7] ), .COUT(
        \mult_26/CARRYB[15][6] ), .SUM(\mult_26/SUMB[15][6] ) );
  FADDER \mult_26/S2_15_5  ( .CIN(\mult_26/ab[15][5] ), .IN0(
        \mult_26/CARRYB[14][5] ), .IN1(\mult_26/SUMB[14][6] ), .COUT(
        \mult_26/CARRYB[15][5] ), .SUM(\mult_26/SUMB[15][5] ) );
  FADDER \mult_26/S2_15_4  ( .CIN(\mult_26/ab[15][4] ), .IN0(
        \mult_26/CARRYB[14][4] ), .IN1(\mult_26/SUMB[14][5] ), .COUT(
        \mult_26/CARRYB[15][4] ), .SUM(\mult_26/SUMB[15][4] ) );
  FADDER \mult_26/S2_15_3  ( .CIN(\mult_26/ab[15][3] ), .IN0(
        \mult_26/CARRYB[14][3] ), .IN1(\mult_26/SUMB[14][4] ), .COUT(
        \mult_26/CARRYB[15][3] ), .SUM(\mult_26/SUMB[15][3] ) );
  FADDER \mult_26/S2_15_2  ( .CIN(\mult_26/ab[15][2] ), .IN0(
        \mult_26/CARRYB[14][2] ), .IN1(\mult_26/SUMB[14][3] ), .COUT(
        \mult_26/CARRYB[15][2] ), .SUM(\mult_26/SUMB[15][2] ) );
  FADDER \mult_26/S2_15_1  ( .CIN(\mult_26/ab[15][1] ), .IN0(
        \mult_26/CARRYB[14][1] ), .IN1(\mult_26/SUMB[14][2] ), .COUT(
        \mult_26/CARRYB[15][1] ), .SUM(\mult_26/SUMB[15][1] ) );
  FADDER \mult_26/S1_15_0  ( .CIN(\mult_26/ab[15][0] ), .IN0(
        \mult_26/CARRYB[14][0] ), .IN1(\mult_26/SUMB[14][1] ), .COUT(
        \mult_26/CARRYB[15][0] ), .SUM(o[15]) );
  FADDER \mult_26/S3_16_30  ( .CIN(\mult_26/ab[16][30] ), .IN0(
        \mult_26/CARRYB[15][30] ), .IN1(\mult_26/ab[15][31] ), .COUT(
        \mult_26/CARRYB[16][30] ), .SUM(\mult_26/SUMB[16][30] ) );
  FADDER \mult_26/S2_16_29  ( .CIN(\mult_26/ab[16][29] ), .IN0(
        \mult_26/CARRYB[15][29] ), .IN1(\mult_26/SUMB[15][30] ), .COUT(
        \mult_26/CARRYB[16][29] ), .SUM(\mult_26/SUMB[16][29] ) );
  FADDER \mult_26/S2_16_28  ( .CIN(\mult_26/ab[16][28] ), .IN0(
        \mult_26/CARRYB[15][28] ), .IN1(\mult_26/SUMB[15][29] ), .COUT(
        \mult_26/CARRYB[16][28] ), .SUM(\mult_26/SUMB[16][28] ) );
  FADDER \mult_26/S2_16_27  ( .CIN(\mult_26/ab[16][27] ), .IN0(
        \mult_26/CARRYB[15][27] ), .IN1(\mult_26/SUMB[15][28] ), .COUT(
        \mult_26/CARRYB[16][27] ), .SUM(\mult_26/SUMB[16][27] ) );
  FADDER \mult_26/S2_16_26  ( .CIN(\mult_26/ab[16][26] ), .IN0(
        \mult_26/CARRYB[15][26] ), .IN1(\mult_26/SUMB[15][27] ), .COUT(
        \mult_26/CARRYB[16][26] ), .SUM(\mult_26/SUMB[16][26] ) );
  FADDER \mult_26/S2_16_25  ( .CIN(\mult_26/ab[16][25] ), .IN0(
        \mult_26/CARRYB[15][25] ), .IN1(\mult_26/SUMB[15][26] ), .COUT(
        \mult_26/CARRYB[16][25] ), .SUM(\mult_26/SUMB[16][25] ) );
  FADDER \mult_26/S2_16_24  ( .CIN(\mult_26/ab[16][24] ), .IN0(
        \mult_26/CARRYB[15][24] ), .IN1(\mult_26/SUMB[15][25] ), .COUT(
        \mult_26/CARRYB[16][24] ), .SUM(\mult_26/SUMB[16][24] ) );
  FADDER \mult_26/S2_16_23  ( .CIN(\mult_26/ab[16][23] ), .IN0(
        \mult_26/CARRYB[15][23] ), .IN1(\mult_26/SUMB[15][24] ), .COUT(
        \mult_26/CARRYB[16][23] ), .SUM(\mult_26/SUMB[16][23] ) );
  FADDER \mult_26/S2_16_22  ( .CIN(\mult_26/ab[16][22] ), .IN0(
        \mult_26/CARRYB[15][22] ), .IN1(\mult_26/SUMB[15][23] ), .COUT(
        \mult_26/CARRYB[16][22] ), .SUM(\mult_26/SUMB[16][22] ) );
  FADDER \mult_26/S2_16_21  ( .CIN(\mult_26/ab[16][21] ), .IN0(
        \mult_26/CARRYB[15][21] ), .IN1(\mult_26/SUMB[15][22] ), .COUT(
        \mult_26/CARRYB[16][21] ), .SUM(\mult_26/SUMB[16][21] ) );
  FADDER \mult_26/S2_16_20  ( .CIN(\mult_26/ab[16][20] ), .IN0(
        \mult_26/CARRYB[15][20] ), .IN1(\mult_26/SUMB[15][21] ), .COUT(
        \mult_26/CARRYB[16][20] ), .SUM(\mult_26/SUMB[16][20] ) );
  FADDER \mult_26/S2_16_19  ( .CIN(\mult_26/ab[16][19] ), .IN0(
        \mult_26/CARRYB[15][19] ), .IN1(\mult_26/SUMB[15][20] ), .COUT(
        \mult_26/CARRYB[16][19] ), .SUM(\mult_26/SUMB[16][19] ) );
  FADDER \mult_26/S2_16_18  ( .CIN(\mult_26/ab[16][18] ), .IN0(
        \mult_26/CARRYB[15][18] ), .IN1(\mult_26/SUMB[15][19] ), .COUT(
        \mult_26/CARRYB[16][18] ), .SUM(\mult_26/SUMB[16][18] ) );
  FADDER \mult_26/S2_16_17  ( .CIN(\mult_26/ab[16][17] ), .IN0(
        \mult_26/CARRYB[15][17] ), .IN1(\mult_26/SUMB[15][18] ), .COUT(
        \mult_26/CARRYB[16][17] ), .SUM(\mult_26/SUMB[16][17] ) );
  FADDER \mult_26/S2_16_16  ( .CIN(\mult_26/ab[16][16] ), .IN0(
        \mult_26/CARRYB[15][16] ), .IN1(\mult_26/SUMB[15][17] ), .COUT(
        \mult_26/CARRYB[16][16] ), .SUM(\mult_26/SUMB[16][16] ) );
  FADDER \mult_26/S2_16_15  ( .CIN(\mult_26/ab[16][15] ), .IN0(
        \mult_26/CARRYB[15][15] ), .IN1(\mult_26/SUMB[15][16] ), .COUT(
        \mult_26/CARRYB[16][15] ), .SUM(\mult_26/SUMB[16][15] ) );
  FADDER \mult_26/S2_16_14  ( .CIN(\mult_26/ab[16][14] ), .IN0(
        \mult_26/CARRYB[15][14] ), .IN1(\mult_26/SUMB[15][15] ), .COUT(
        \mult_26/CARRYB[16][14] ), .SUM(\mult_26/SUMB[16][14] ) );
  FADDER \mult_26/S2_16_13  ( .CIN(\mult_26/ab[16][13] ), .IN0(
        \mult_26/CARRYB[15][13] ), .IN1(\mult_26/SUMB[15][14] ), .COUT(
        \mult_26/CARRYB[16][13] ), .SUM(\mult_26/SUMB[16][13] ) );
  FADDER \mult_26/S2_16_12  ( .CIN(\mult_26/ab[16][12] ), .IN0(
        \mult_26/CARRYB[15][12] ), .IN1(\mult_26/SUMB[15][13] ), .COUT(
        \mult_26/CARRYB[16][12] ), .SUM(\mult_26/SUMB[16][12] ) );
  FADDER \mult_26/S2_16_11  ( .CIN(\mult_26/ab[16][11] ), .IN0(
        \mult_26/CARRYB[15][11] ), .IN1(\mult_26/SUMB[15][12] ), .COUT(
        \mult_26/CARRYB[16][11] ), .SUM(\mult_26/SUMB[16][11] ) );
  FADDER \mult_26/S2_16_10  ( .CIN(\mult_26/ab[16][10] ), .IN0(
        \mult_26/CARRYB[15][10] ), .IN1(\mult_26/SUMB[15][11] ), .COUT(
        \mult_26/CARRYB[16][10] ), .SUM(\mult_26/SUMB[16][10] ) );
  FADDER \mult_26/S2_16_9  ( .CIN(\mult_26/ab[16][9] ), .IN0(
        \mult_26/CARRYB[15][9] ), .IN1(\mult_26/SUMB[15][10] ), .COUT(
        \mult_26/CARRYB[16][9] ), .SUM(\mult_26/SUMB[16][9] ) );
  FADDER \mult_26/S2_16_8  ( .CIN(\mult_26/ab[16][8] ), .IN0(
        \mult_26/CARRYB[15][8] ), .IN1(\mult_26/SUMB[15][9] ), .COUT(
        \mult_26/CARRYB[16][8] ), .SUM(\mult_26/SUMB[16][8] ) );
  FADDER \mult_26/S2_16_7  ( .CIN(\mult_26/ab[16][7] ), .IN0(
        \mult_26/CARRYB[15][7] ), .IN1(\mult_26/SUMB[15][8] ), .COUT(
        \mult_26/CARRYB[16][7] ), .SUM(\mult_26/SUMB[16][7] ) );
  FADDER \mult_26/S2_16_6  ( .CIN(\mult_26/ab[16][6] ), .IN0(
        \mult_26/CARRYB[15][6] ), .IN1(\mult_26/SUMB[15][7] ), .COUT(
        \mult_26/CARRYB[16][6] ), .SUM(\mult_26/SUMB[16][6] ) );
  FADDER \mult_26/S2_16_5  ( .CIN(\mult_26/ab[16][5] ), .IN0(
        \mult_26/CARRYB[15][5] ), .IN1(\mult_26/SUMB[15][6] ), .COUT(
        \mult_26/CARRYB[16][5] ), .SUM(\mult_26/SUMB[16][5] ) );
  FADDER \mult_26/S2_16_4  ( .CIN(\mult_26/ab[16][4] ), .IN0(
        \mult_26/CARRYB[15][4] ), .IN1(\mult_26/SUMB[15][5] ), .COUT(
        \mult_26/CARRYB[16][4] ), .SUM(\mult_26/SUMB[16][4] ) );
  FADDER \mult_26/S2_16_3  ( .CIN(\mult_26/ab[16][3] ), .IN0(
        \mult_26/CARRYB[15][3] ), .IN1(\mult_26/SUMB[15][4] ), .COUT(
        \mult_26/CARRYB[16][3] ), .SUM(\mult_26/SUMB[16][3] ) );
  FADDER \mult_26/S2_16_2  ( .CIN(\mult_26/ab[16][2] ), .IN0(
        \mult_26/CARRYB[15][2] ), .IN1(\mult_26/SUMB[15][3] ), .COUT(
        \mult_26/CARRYB[16][2] ), .SUM(\mult_26/SUMB[16][2] ) );
  FADDER \mult_26/S2_16_1  ( .CIN(\mult_26/ab[16][1] ), .IN0(
        \mult_26/CARRYB[15][1] ), .IN1(\mult_26/SUMB[15][2] ), .COUT(
        \mult_26/CARRYB[16][1] ), .SUM(\mult_26/SUMB[16][1] ) );
  FADDER \mult_26/S1_16_0  ( .CIN(\mult_26/ab[16][0] ), .IN0(
        \mult_26/CARRYB[15][0] ), .IN1(\mult_26/SUMB[15][1] ), .COUT(
        \mult_26/CARRYB[16][0] ), .SUM(o[16]) );
  FADDER \mult_26/S3_17_30  ( .CIN(\mult_26/ab[17][30] ), .IN0(
        \mult_26/CARRYB[16][30] ), .IN1(\mult_26/ab[16][31] ), .COUT(
        \mult_26/CARRYB[17][30] ), .SUM(\mult_26/SUMB[17][30] ) );
  FADDER \mult_26/S2_17_29  ( .CIN(\mult_26/ab[17][29] ), .IN0(
        \mult_26/CARRYB[16][29] ), .IN1(\mult_26/SUMB[16][30] ), .COUT(
        \mult_26/CARRYB[17][29] ), .SUM(\mult_26/SUMB[17][29] ) );
  FADDER \mult_26/S2_17_28  ( .CIN(\mult_26/ab[17][28] ), .IN0(
        \mult_26/CARRYB[16][28] ), .IN1(\mult_26/SUMB[16][29] ), .COUT(
        \mult_26/CARRYB[17][28] ), .SUM(\mult_26/SUMB[17][28] ) );
  FADDER \mult_26/S2_17_27  ( .CIN(\mult_26/ab[17][27] ), .IN0(
        \mult_26/CARRYB[16][27] ), .IN1(\mult_26/SUMB[16][28] ), .COUT(
        \mult_26/CARRYB[17][27] ), .SUM(\mult_26/SUMB[17][27] ) );
  FADDER \mult_26/S2_17_26  ( .CIN(\mult_26/ab[17][26] ), .IN0(
        \mult_26/CARRYB[16][26] ), .IN1(\mult_26/SUMB[16][27] ), .COUT(
        \mult_26/CARRYB[17][26] ), .SUM(\mult_26/SUMB[17][26] ) );
  FADDER \mult_26/S2_17_25  ( .CIN(\mult_26/ab[17][25] ), .IN0(
        \mult_26/CARRYB[16][25] ), .IN1(\mult_26/SUMB[16][26] ), .COUT(
        \mult_26/CARRYB[17][25] ), .SUM(\mult_26/SUMB[17][25] ) );
  FADDER \mult_26/S2_17_24  ( .CIN(\mult_26/ab[17][24] ), .IN0(
        \mult_26/CARRYB[16][24] ), .IN1(\mult_26/SUMB[16][25] ), .COUT(
        \mult_26/CARRYB[17][24] ), .SUM(\mult_26/SUMB[17][24] ) );
  FADDER \mult_26/S2_17_23  ( .CIN(\mult_26/ab[17][23] ), .IN0(
        \mult_26/CARRYB[16][23] ), .IN1(\mult_26/SUMB[16][24] ), .COUT(
        \mult_26/CARRYB[17][23] ), .SUM(\mult_26/SUMB[17][23] ) );
  FADDER \mult_26/S2_17_22  ( .CIN(\mult_26/ab[17][22] ), .IN0(
        \mult_26/CARRYB[16][22] ), .IN1(\mult_26/SUMB[16][23] ), .COUT(
        \mult_26/CARRYB[17][22] ), .SUM(\mult_26/SUMB[17][22] ) );
  FADDER \mult_26/S2_17_21  ( .CIN(\mult_26/ab[17][21] ), .IN0(
        \mult_26/CARRYB[16][21] ), .IN1(\mult_26/SUMB[16][22] ), .COUT(
        \mult_26/CARRYB[17][21] ), .SUM(\mult_26/SUMB[17][21] ) );
  FADDER \mult_26/S2_17_20  ( .CIN(\mult_26/ab[17][20] ), .IN0(
        \mult_26/CARRYB[16][20] ), .IN1(\mult_26/SUMB[16][21] ), .COUT(
        \mult_26/CARRYB[17][20] ), .SUM(\mult_26/SUMB[17][20] ) );
  FADDER \mult_26/S2_17_19  ( .CIN(\mult_26/ab[17][19] ), .IN0(
        \mult_26/CARRYB[16][19] ), .IN1(\mult_26/SUMB[16][20] ), .COUT(
        \mult_26/CARRYB[17][19] ), .SUM(\mult_26/SUMB[17][19] ) );
  FADDER \mult_26/S2_17_18  ( .CIN(\mult_26/ab[17][18] ), .IN0(
        \mult_26/CARRYB[16][18] ), .IN1(\mult_26/SUMB[16][19] ), .COUT(
        \mult_26/CARRYB[17][18] ), .SUM(\mult_26/SUMB[17][18] ) );
  FADDER \mult_26/S2_17_17  ( .CIN(\mult_26/ab[17][17] ), .IN0(
        \mult_26/CARRYB[16][17] ), .IN1(\mult_26/SUMB[16][18] ), .COUT(
        \mult_26/CARRYB[17][17] ), .SUM(\mult_26/SUMB[17][17] ) );
  FADDER \mult_26/S2_17_16  ( .CIN(\mult_26/ab[17][16] ), .IN0(
        \mult_26/CARRYB[16][16] ), .IN1(\mult_26/SUMB[16][17] ), .COUT(
        \mult_26/CARRYB[17][16] ), .SUM(\mult_26/SUMB[17][16] ) );
  FADDER \mult_26/S2_17_15  ( .CIN(\mult_26/ab[17][15] ), .IN0(
        \mult_26/CARRYB[16][15] ), .IN1(\mult_26/SUMB[16][16] ), .COUT(
        \mult_26/CARRYB[17][15] ), .SUM(\mult_26/SUMB[17][15] ) );
  FADDER \mult_26/S2_17_14  ( .CIN(\mult_26/ab[17][14] ), .IN0(
        \mult_26/CARRYB[16][14] ), .IN1(\mult_26/SUMB[16][15] ), .COUT(
        \mult_26/CARRYB[17][14] ), .SUM(\mult_26/SUMB[17][14] ) );
  FADDER \mult_26/S2_17_13  ( .CIN(\mult_26/ab[17][13] ), .IN0(
        \mult_26/CARRYB[16][13] ), .IN1(\mult_26/SUMB[16][14] ), .COUT(
        \mult_26/CARRYB[17][13] ), .SUM(\mult_26/SUMB[17][13] ) );
  FADDER \mult_26/S2_17_12  ( .CIN(\mult_26/ab[17][12] ), .IN0(
        \mult_26/CARRYB[16][12] ), .IN1(\mult_26/SUMB[16][13] ), .COUT(
        \mult_26/CARRYB[17][12] ), .SUM(\mult_26/SUMB[17][12] ) );
  FADDER \mult_26/S2_17_11  ( .CIN(\mult_26/ab[17][11] ), .IN0(
        \mult_26/CARRYB[16][11] ), .IN1(\mult_26/SUMB[16][12] ), .COUT(
        \mult_26/CARRYB[17][11] ), .SUM(\mult_26/SUMB[17][11] ) );
  FADDER \mult_26/S2_17_10  ( .CIN(\mult_26/ab[17][10] ), .IN0(
        \mult_26/CARRYB[16][10] ), .IN1(\mult_26/SUMB[16][11] ), .COUT(
        \mult_26/CARRYB[17][10] ), .SUM(\mult_26/SUMB[17][10] ) );
  FADDER \mult_26/S2_17_9  ( .CIN(\mult_26/ab[17][9] ), .IN0(
        \mult_26/CARRYB[16][9] ), .IN1(\mult_26/SUMB[16][10] ), .COUT(
        \mult_26/CARRYB[17][9] ), .SUM(\mult_26/SUMB[17][9] ) );
  FADDER \mult_26/S2_17_8  ( .CIN(\mult_26/ab[17][8] ), .IN0(
        \mult_26/CARRYB[16][8] ), .IN1(\mult_26/SUMB[16][9] ), .COUT(
        \mult_26/CARRYB[17][8] ), .SUM(\mult_26/SUMB[17][8] ) );
  FADDER \mult_26/S2_17_7  ( .CIN(\mult_26/ab[17][7] ), .IN0(
        \mult_26/CARRYB[16][7] ), .IN1(\mult_26/SUMB[16][8] ), .COUT(
        \mult_26/CARRYB[17][7] ), .SUM(\mult_26/SUMB[17][7] ) );
  FADDER \mult_26/S2_17_6  ( .CIN(\mult_26/ab[17][6] ), .IN0(
        \mult_26/CARRYB[16][6] ), .IN1(\mult_26/SUMB[16][7] ), .COUT(
        \mult_26/CARRYB[17][6] ), .SUM(\mult_26/SUMB[17][6] ) );
  FADDER \mult_26/S2_17_5  ( .CIN(\mult_26/ab[17][5] ), .IN0(
        \mult_26/CARRYB[16][5] ), .IN1(\mult_26/SUMB[16][6] ), .COUT(
        \mult_26/CARRYB[17][5] ), .SUM(\mult_26/SUMB[17][5] ) );
  FADDER \mult_26/S2_17_4  ( .CIN(\mult_26/ab[17][4] ), .IN0(
        \mult_26/CARRYB[16][4] ), .IN1(\mult_26/SUMB[16][5] ), .COUT(
        \mult_26/CARRYB[17][4] ), .SUM(\mult_26/SUMB[17][4] ) );
  FADDER \mult_26/S2_17_3  ( .CIN(\mult_26/ab[17][3] ), .IN0(
        \mult_26/CARRYB[16][3] ), .IN1(\mult_26/SUMB[16][4] ), .COUT(
        \mult_26/CARRYB[17][3] ), .SUM(\mult_26/SUMB[17][3] ) );
  FADDER \mult_26/S2_17_2  ( .CIN(\mult_26/ab[17][2] ), .IN0(
        \mult_26/CARRYB[16][2] ), .IN1(\mult_26/SUMB[16][3] ), .COUT(
        \mult_26/CARRYB[17][2] ), .SUM(\mult_26/SUMB[17][2] ) );
  FADDER \mult_26/S2_17_1  ( .CIN(\mult_26/ab[17][1] ), .IN0(
        \mult_26/CARRYB[16][1] ), .IN1(\mult_26/SUMB[16][2] ), .COUT(
        \mult_26/CARRYB[17][1] ), .SUM(\mult_26/SUMB[17][1] ) );
  FADDER \mult_26/S1_17_0  ( .CIN(\mult_26/ab[17][0] ), .IN0(
        \mult_26/CARRYB[16][0] ), .IN1(\mult_26/SUMB[16][1] ), .COUT(
        \mult_26/CARRYB[17][0] ), .SUM(o[17]) );
  FADDER \mult_26/S3_18_30  ( .CIN(\mult_26/ab[18][30] ), .IN0(
        \mult_26/CARRYB[17][30] ), .IN1(\mult_26/ab[17][31] ), .COUT(
        \mult_26/CARRYB[18][30] ), .SUM(\mult_26/SUMB[18][30] ) );
  FADDER \mult_26/S2_18_29  ( .CIN(\mult_26/ab[18][29] ), .IN0(
        \mult_26/CARRYB[17][29] ), .IN1(\mult_26/SUMB[17][30] ), .COUT(
        \mult_26/CARRYB[18][29] ), .SUM(\mult_26/SUMB[18][29] ) );
  FADDER \mult_26/S2_18_28  ( .CIN(\mult_26/ab[18][28] ), .IN0(
        \mult_26/CARRYB[17][28] ), .IN1(\mult_26/SUMB[17][29] ), .COUT(
        \mult_26/CARRYB[18][28] ), .SUM(\mult_26/SUMB[18][28] ) );
  FADDER \mult_26/S2_18_27  ( .CIN(\mult_26/ab[18][27] ), .IN0(
        \mult_26/CARRYB[17][27] ), .IN1(\mult_26/SUMB[17][28] ), .COUT(
        \mult_26/CARRYB[18][27] ), .SUM(\mult_26/SUMB[18][27] ) );
  FADDER \mult_26/S2_18_26  ( .CIN(\mult_26/ab[18][26] ), .IN0(
        \mult_26/CARRYB[17][26] ), .IN1(\mult_26/SUMB[17][27] ), .COUT(
        \mult_26/CARRYB[18][26] ), .SUM(\mult_26/SUMB[18][26] ) );
  FADDER \mult_26/S2_18_25  ( .CIN(\mult_26/ab[18][25] ), .IN0(
        \mult_26/CARRYB[17][25] ), .IN1(\mult_26/SUMB[17][26] ), .COUT(
        \mult_26/CARRYB[18][25] ), .SUM(\mult_26/SUMB[18][25] ) );
  FADDER \mult_26/S2_18_24  ( .CIN(\mult_26/ab[18][24] ), .IN0(
        \mult_26/CARRYB[17][24] ), .IN1(\mult_26/SUMB[17][25] ), .COUT(
        \mult_26/CARRYB[18][24] ), .SUM(\mult_26/SUMB[18][24] ) );
  FADDER \mult_26/S2_18_23  ( .CIN(\mult_26/ab[18][23] ), .IN0(
        \mult_26/CARRYB[17][23] ), .IN1(\mult_26/SUMB[17][24] ), .COUT(
        \mult_26/CARRYB[18][23] ), .SUM(\mult_26/SUMB[18][23] ) );
  FADDER \mult_26/S2_18_22  ( .CIN(\mult_26/ab[18][22] ), .IN0(
        \mult_26/CARRYB[17][22] ), .IN1(\mult_26/SUMB[17][23] ), .COUT(
        \mult_26/CARRYB[18][22] ), .SUM(\mult_26/SUMB[18][22] ) );
  FADDER \mult_26/S2_18_21  ( .CIN(\mult_26/ab[18][21] ), .IN0(
        \mult_26/CARRYB[17][21] ), .IN1(\mult_26/SUMB[17][22] ), .COUT(
        \mult_26/CARRYB[18][21] ), .SUM(\mult_26/SUMB[18][21] ) );
  FADDER \mult_26/S2_18_20  ( .CIN(\mult_26/ab[18][20] ), .IN0(
        \mult_26/CARRYB[17][20] ), .IN1(\mult_26/SUMB[17][21] ), .COUT(
        \mult_26/CARRYB[18][20] ), .SUM(\mult_26/SUMB[18][20] ) );
  FADDER \mult_26/S2_18_19  ( .CIN(\mult_26/ab[18][19] ), .IN0(
        \mult_26/CARRYB[17][19] ), .IN1(\mult_26/SUMB[17][20] ), .COUT(
        \mult_26/CARRYB[18][19] ), .SUM(\mult_26/SUMB[18][19] ) );
  FADDER \mult_26/S2_18_18  ( .CIN(\mult_26/ab[18][18] ), .IN0(
        \mult_26/CARRYB[17][18] ), .IN1(\mult_26/SUMB[17][19] ), .COUT(
        \mult_26/CARRYB[18][18] ), .SUM(\mult_26/SUMB[18][18] ) );
  FADDER \mult_26/S2_18_17  ( .CIN(\mult_26/ab[18][17] ), .IN0(
        \mult_26/CARRYB[17][17] ), .IN1(\mult_26/SUMB[17][18] ), .COUT(
        \mult_26/CARRYB[18][17] ), .SUM(\mult_26/SUMB[18][17] ) );
  FADDER \mult_26/S2_18_16  ( .CIN(\mult_26/ab[18][16] ), .IN0(
        \mult_26/CARRYB[17][16] ), .IN1(\mult_26/SUMB[17][17] ), .COUT(
        \mult_26/CARRYB[18][16] ), .SUM(\mult_26/SUMB[18][16] ) );
  FADDER \mult_26/S2_18_15  ( .CIN(\mult_26/ab[18][15] ), .IN0(
        \mult_26/CARRYB[17][15] ), .IN1(\mult_26/SUMB[17][16] ), .COUT(
        \mult_26/CARRYB[18][15] ), .SUM(\mult_26/SUMB[18][15] ) );
  FADDER \mult_26/S2_18_14  ( .CIN(\mult_26/ab[18][14] ), .IN0(
        \mult_26/CARRYB[17][14] ), .IN1(\mult_26/SUMB[17][15] ), .COUT(
        \mult_26/CARRYB[18][14] ), .SUM(\mult_26/SUMB[18][14] ) );
  FADDER \mult_26/S2_18_13  ( .CIN(\mult_26/ab[18][13] ), .IN0(
        \mult_26/CARRYB[17][13] ), .IN1(\mult_26/SUMB[17][14] ), .COUT(
        \mult_26/CARRYB[18][13] ), .SUM(\mult_26/SUMB[18][13] ) );
  FADDER \mult_26/S2_18_12  ( .CIN(\mult_26/ab[18][12] ), .IN0(
        \mult_26/CARRYB[17][12] ), .IN1(\mult_26/SUMB[17][13] ), .COUT(
        \mult_26/CARRYB[18][12] ), .SUM(\mult_26/SUMB[18][12] ) );
  FADDER \mult_26/S2_18_11  ( .CIN(\mult_26/ab[18][11] ), .IN0(
        \mult_26/CARRYB[17][11] ), .IN1(\mult_26/SUMB[17][12] ), .COUT(
        \mult_26/CARRYB[18][11] ), .SUM(\mult_26/SUMB[18][11] ) );
  FADDER \mult_26/S2_18_10  ( .CIN(\mult_26/ab[18][10] ), .IN0(
        \mult_26/CARRYB[17][10] ), .IN1(\mult_26/SUMB[17][11] ), .COUT(
        \mult_26/CARRYB[18][10] ), .SUM(\mult_26/SUMB[18][10] ) );
  FADDER \mult_26/S2_18_9  ( .CIN(\mult_26/ab[18][9] ), .IN0(
        \mult_26/CARRYB[17][9] ), .IN1(\mult_26/SUMB[17][10] ), .COUT(
        \mult_26/CARRYB[18][9] ), .SUM(\mult_26/SUMB[18][9] ) );
  FADDER \mult_26/S2_18_8  ( .CIN(\mult_26/ab[18][8] ), .IN0(
        \mult_26/CARRYB[17][8] ), .IN1(\mult_26/SUMB[17][9] ), .COUT(
        \mult_26/CARRYB[18][8] ), .SUM(\mult_26/SUMB[18][8] ) );
  FADDER \mult_26/S2_18_7  ( .CIN(\mult_26/ab[18][7] ), .IN0(
        \mult_26/CARRYB[17][7] ), .IN1(\mult_26/SUMB[17][8] ), .COUT(
        \mult_26/CARRYB[18][7] ), .SUM(\mult_26/SUMB[18][7] ) );
  FADDER \mult_26/S2_18_6  ( .CIN(\mult_26/ab[18][6] ), .IN0(
        \mult_26/CARRYB[17][6] ), .IN1(\mult_26/SUMB[17][7] ), .COUT(
        \mult_26/CARRYB[18][6] ), .SUM(\mult_26/SUMB[18][6] ) );
  FADDER \mult_26/S2_18_5  ( .CIN(\mult_26/ab[18][5] ), .IN0(
        \mult_26/CARRYB[17][5] ), .IN1(\mult_26/SUMB[17][6] ), .COUT(
        \mult_26/CARRYB[18][5] ), .SUM(\mult_26/SUMB[18][5] ) );
  FADDER \mult_26/S2_18_4  ( .CIN(\mult_26/ab[18][4] ), .IN0(
        \mult_26/CARRYB[17][4] ), .IN1(\mult_26/SUMB[17][5] ), .COUT(
        \mult_26/CARRYB[18][4] ), .SUM(\mult_26/SUMB[18][4] ) );
  FADDER \mult_26/S2_18_3  ( .CIN(\mult_26/ab[18][3] ), .IN0(
        \mult_26/CARRYB[17][3] ), .IN1(\mult_26/SUMB[17][4] ), .COUT(
        \mult_26/CARRYB[18][3] ), .SUM(\mult_26/SUMB[18][3] ) );
  FADDER \mult_26/S2_18_2  ( .CIN(\mult_26/ab[18][2] ), .IN0(
        \mult_26/CARRYB[17][2] ), .IN1(\mult_26/SUMB[17][3] ), .COUT(
        \mult_26/CARRYB[18][2] ), .SUM(\mult_26/SUMB[18][2] ) );
  FADDER \mult_26/S2_18_1  ( .CIN(\mult_26/ab[18][1] ), .IN0(
        \mult_26/CARRYB[17][1] ), .IN1(\mult_26/SUMB[17][2] ), .COUT(
        \mult_26/CARRYB[18][1] ), .SUM(\mult_26/SUMB[18][1] ) );
  FADDER \mult_26/S1_18_0  ( .CIN(\mult_26/ab[18][0] ), .IN0(
        \mult_26/CARRYB[17][0] ), .IN1(\mult_26/SUMB[17][1] ), .COUT(
        \mult_26/CARRYB[18][0] ), .SUM(o[18]) );
  FADDER \mult_26/S3_19_30  ( .CIN(\mult_26/ab[19][30] ), .IN0(
        \mult_26/CARRYB[18][30] ), .IN1(\mult_26/ab[18][31] ), .COUT(
        \mult_26/CARRYB[19][30] ), .SUM(\mult_26/SUMB[19][30] ) );
  FADDER \mult_26/S2_19_29  ( .CIN(\mult_26/ab[19][29] ), .IN0(
        \mult_26/CARRYB[18][29] ), .IN1(\mult_26/SUMB[18][30] ), .COUT(
        \mult_26/CARRYB[19][29] ), .SUM(\mult_26/SUMB[19][29] ) );
  FADDER \mult_26/S2_19_28  ( .CIN(\mult_26/ab[19][28] ), .IN0(
        \mult_26/CARRYB[18][28] ), .IN1(\mult_26/SUMB[18][29] ), .COUT(
        \mult_26/CARRYB[19][28] ), .SUM(\mult_26/SUMB[19][28] ) );
  FADDER \mult_26/S2_19_27  ( .CIN(\mult_26/ab[19][27] ), .IN0(
        \mult_26/CARRYB[18][27] ), .IN1(\mult_26/SUMB[18][28] ), .COUT(
        \mult_26/CARRYB[19][27] ), .SUM(\mult_26/SUMB[19][27] ) );
  FADDER \mult_26/S2_19_26  ( .CIN(\mult_26/ab[19][26] ), .IN0(
        \mult_26/CARRYB[18][26] ), .IN1(\mult_26/SUMB[18][27] ), .COUT(
        \mult_26/CARRYB[19][26] ), .SUM(\mult_26/SUMB[19][26] ) );
  FADDER \mult_26/S2_19_25  ( .CIN(\mult_26/ab[19][25] ), .IN0(
        \mult_26/CARRYB[18][25] ), .IN1(\mult_26/SUMB[18][26] ), .COUT(
        \mult_26/CARRYB[19][25] ), .SUM(\mult_26/SUMB[19][25] ) );
  FADDER \mult_26/S2_19_24  ( .CIN(\mult_26/ab[19][24] ), .IN0(
        \mult_26/CARRYB[18][24] ), .IN1(\mult_26/SUMB[18][25] ), .COUT(
        \mult_26/CARRYB[19][24] ), .SUM(\mult_26/SUMB[19][24] ) );
  FADDER \mult_26/S2_19_23  ( .CIN(\mult_26/ab[19][23] ), .IN0(
        \mult_26/CARRYB[18][23] ), .IN1(\mult_26/SUMB[18][24] ), .COUT(
        \mult_26/CARRYB[19][23] ), .SUM(\mult_26/SUMB[19][23] ) );
  FADDER \mult_26/S2_19_22  ( .CIN(\mult_26/ab[19][22] ), .IN0(
        \mult_26/CARRYB[18][22] ), .IN1(\mult_26/SUMB[18][23] ), .COUT(
        \mult_26/CARRYB[19][22] ), .SUM(\mult_26/SUMB[19][22] ) );
  FADDER \mult_26/S2_19_21  ( .CIN(\mult_26/ab[19][21] ), .IN0(
        \mult_26/CARRYB[18][21] ), .IN1(\mult_26/SUMB[18][22] ), .COUT(
        \mult_26/CARRYB[19][21] ), .SUM(\mult_26/SUMB[19][21] ) );
  FADDER \mult_26/S2_19_20  ( .CIN(\mult_26/ab[19][20] ), .IN0(
        \mult_26/CARRYB[18][20] ), .IN1(\mult_26/SUMB[18][21] ), .COUT(
        \mult_26/CARRYB[19][20] ), .SUM(\mult_26/SUMB[19][20] ) );
  FADDER \mult_26/S2_19_19  ( .CIN(\mult_26/ab[19][19] ), .IN0(
        \mult_26/CARRYB[18][19] ), .IN1(\mult_26/SUMB[18][20] ), .COUT(
        \mult_26/CARRYB[19][19] ), .SUM(\mult_26/SUMB[19][19] ) );
  FADDER \mult_26/S2_19_18  ( .CIN(\mult_26/ab[19][18] ), .IN0(
        \mult_26/CARRYB[18][18] ), .IN1(\mult_26/SUMB[18][19] ), .COUT(
        \mult_26/CARRYB[19][18] ), .SUM(\mult_26/SUMB[19][18] ) );
  FADDER \mult_26/S2_19_17  ( .CIN(\mult_26/ab[19][17] ), .IN0(
        \mult_26/CARRYB[18][17] ), .IN1(\mult_26/SUMB[18][18] ), .COUT(
        \mult_26/CARRYB[19][17] ), .SUM(\mult_26/SUMB[19][17] ) );
  FADDER \mult_26/S2_19_16  ( .CIN(\mult_26/ab[19][16] ), .IN0(
        \mult_26/CARRYB[18][16] ), .IN1(\mult_26/SUMB[18][17] ), .COUT(
        \mult_26/CARRYB[19][16] ), .SUM(\mult_26/SUMB[19][16] ) );
  FADDER \mult_26/S2_19_15  ( .CIN(\mult_26/ab[19][15] ), .IN0(
        \mult_26/CARRYB[18][15] ), .IN1(\mult_26/SUMB[18][16] ), .COUT(
        \mult_26/CARRYB[19][15] ), .SUM(\mult_26/SUMB[19][15] ) );
  FADDER \mult_26/S2_19_14  ( .CIN(\mult_26/ab[19][14] ), .IN0(
        \mult_26/CARRYB[18][14] ), .IN1(\mult_26/SUMB[18][15] ), .COUT(
        \mult_26/CARRYB[19][14] ), .SUM(\mult_26/SUMB[19][14] ) );
  FADDER \mult_26/S2_19_13  ( .CIN(\mult_26/ab[19][13] ), .IN0(
        \mult_26/CARRYB[18][13] ), .IN1(\mult_26/SUMB[18][14] ), .COUT(
        \mult_26/CARRYB[19][13] ), .SUM(\mult_26/SUMB[19][13] ) );
  FADDER \mult_26/S2_19_12  ( .CIN(\mult_26/ab[19][12] ), .IN0(
        \mult_26/CARRYB[18][12] ), .IN1(\mult_26/SUMB[18][13] ), .COUT(
        \mult_26/CARRYB[19][12] ), .SUM(\mult_26/SUMB[19][12] ) );
  FADDER \mult_26/S2_19_11  ( .CIN(\mult_26/ab[19][11] ), .IN0(
        \mult_26/CARRYB[18][11] ), .IN1(\mult_26/SUMB[18][12] ), .COUT(
        \mult_26/CARRYB[19][11] ), .SUM(\mult_26/SUMB[19][11] ) );
  FADDER \mult_26/S2_19_10  ( .CIN(\mult_26/ab[19][10] ), .IN0(
        \mult_26/CARRYB[18][10] ), .IN1(\mult_26/SUMB[18][11] ), .COUT(
        \mult_26/CARRYB[19][10] ), .SUM(\mult_26/SUMB[19][10] ) );
  FADDER \mult_26/S2_19_9  ( .CIN(\mult_26/ab[19][9] ), .IN0(
        \mult_26/CARRYB[18][9] ), .IN1(\mult_26/SUMB[18][10] ), .COUT(
        \mult_26/CARRYB[19][9] ), .SUM(\mult_26/SUMB[19][9] ) );
  FADDER \mult_26/S2_19_8  ( .CIN(\mult_26/ab[19][8] ), .IN0(
        \mult_26/CARRYB[18][8] ), .IN1(\mult_26/SUMB[18][9] ), .COUT(
        \mult_26/CARRYB[19][8] ), .SUM(\mult_26/SUMB[19][8] ) );
  FADDER \mult_26/S2_19_7  ( .CIN(\mult_26/ab[19][7] ), .IN0(
        \mult_26/CARRYB[18][7] ), .IN1(\mult_26/SUMB[18][8] ), .COUT(
        \mult_26/CARRYB[19][7] ), .SUM(\mult_26/SUMB[19][7] ) );
  FADDER \mult_26/S2_19_6  ( .CIN(\mult_26/ab[19][6] ), .IN0(
        \mult_26/CARRYB[18][6] ), .IN1(\mult_26/SUMB[18][7] ), .COUT(
        \mult_26/CARRYB[19][6] ), .SUM(\mult_26/SUMB[19][6] ) );
  FADDER \mult_26/S2_19_5  ( .CIN(\mult_26/ab[19][5] ), .IN0(
        \mult_26/CARRYB[18][5] ), .IN1(\mult_26/SUMB[18][6] ), .COUT(
        \mult_26/CARRYB[19][5] ), .SUM(\mult_26/SUMB[19][5] ) );
  FADDER \mult_26/S2_19_4  ( .CIN(\mult_26/ab[19][4] ), .IN0(
        \mult_26/CARRYB[18][4] ), .IN1(\mult_26/SUMB[18][5] ), .COUT(
        \mult_26/CARRYB[19][4] ), .SUM(\mult_26/SUMB[19][4] ) );
  FADDER \mult_26/S2_19_3  ( .CIN(\mult_26/ab[19][3] ), .IN0(
        \mult_26/CARRYB[18][3] ), .IN1(\mult_26/SUMB[18][4] ), .COUT(
        \mult_26/CARRYB[19][3] ), .SUM(\mult_26/SUMB[19][3] ) );
  FADDER \mult_26/S2_19_2  ( .CIN(\mult_26/ab[19][2] ), .IN0(
        \mult_26/CARRYB[18][2] ), .IN1(\mult_26/SUMB[18][3] ), .COUT(
        \mult_26/CARRYB[19][2] ), .SUM(\mult_26/SUMB[19][2] ) );
  FADDER \mult_26/S2_19_1  ( .CIN(\mult_26/ab[19][1] ), .IN0(
        \mult_26/CARRYB[18][1] ), .IN1(\mult_26/SUMB[18][2] ), .COUT(
        \mult_26/CARRYB[19][1] ), .SUM(\mult_26/SUMB[19][1] ) );
  FADDER \mult_26/S1_19_0  ( .CIN(\mult_26/ab[19][0] ), .IN0(
        \mult_26/CARRYB[18][0] ), .IN1(\mult_26/SUMB[18][1] ), .COUT(
        \mult_26/CARRYB[19][0] ), .SUM(o[19]) );
  FADDER \mult_26/S3_20_30  ( .CIN(\mult_26/ab[20][30] ), .IN0(
        \mult_26/CARRYB[19][30] ), .IN1(\mult_26/ab[19][31] ), .COUT(
        \mult_26/CARRYB[20][30] ), .SUM(\mult_26/SUMB[20][30] ) );
  FADDER \mult_26/S2_20_29  ( .CIN(\mult_26/ab[20][29] ), .IN0(
        \mult_26/CARRYB[19][29] ), .IN1(\mult_26/SUMB[19][30] ), .COUT(
        \mult_26/CARRYB[20][29] ), .SUM(\mult_26/SUMB[20][29] ) );
  FADDER \mult_26/S2_20_28  ( .CIN(\mult_26/ab[20][28] ), .IN0(
        \mult_26/CARRYB[19][28] ), .IN1(\mult_26/SUMB[19][29] ), .COUT(
        \mult_26/CARRYB[20][28] ), .SUM(\mult_26/SUMB[20][28] ) );
  FADDER \mult_26/S2_20_27  ( .CIN(\mult_26/ab[20][27] ), .IN0(
        \mult_26/CARRYB[19][27] ), .IN1(\mult_26/SUMB[19][28] ), .COUT(
        \mult_26/CARRYB[20][27] ), .SUM(\mult_26/SUMB[20][27] ) );
  FADDER \mult_26/S2_20_26  ( .CIN(\mult_26/ab[20][26] ), .IN0(
        \mult_26/CARRYB[19][26] ), .IN1(\mult_26/SUMB[19][27] ), .COUT(
        \mult_26/CARRYB[20][26] ), .SUM(\mult_26/SUMB[20][26] ) );
  FADDER \mult_26/S2_20_25  ( .CIN(\mult_26/ab[20][25] ), .IN0(
        \mult_26/CARRYB[19][25] ), .IN1(\mult_26/SUMB[19][26] ), .COUT(
        \mult_26/CARRYB[20][25] ), .SUM(\mult_26/SUMB[20][25] ) );
  FADDER \mult_26/S2_20_24  ( .CIN(\mult_26/ab[20][24] ), .IN0(
        \mult_26/CARRYB[19][24] ), .IN1(\mult_26/SUMB[19][25] ), .COUT(
        \mult_26/CARRYB[20][24] ), .SUM(\mult_26/SUMB[20][24] ) );
  FADDER \mult_26/S2_20_23  ( .CIN(\mult_26/ab[20][23] ), .IN0(
        \mult_26/CARRYB[19][23] ), .IN1(\mult_26/SUMB[19][24] ), .COUT(
        \mult_26/CARRYB[20][23] ), .SUM(\mult_26/SUMB[20][23] ) );
  FADDER \mult_26/S2_20_22  ( .CIN(\mult_26/ab[20][22] ), .IN0(
        \mult_26/CARRYB[19][22] ), .IN1(\mult_26/SUMB[19][23] ), .COUT(
        \mult_26/CARRYB[20][22] ), .SUM(\mult_26/SUMB[20][22] ) );
  FADDER \mult_26/S2_20_21  ( .CIN(\mult_26/ab[20][21] ), .IN0(
        \mult_26/CARRYB[19][21] ), .IN1(\mult_26/SUMB[19][22] ), .COUT(
        \mult_26/CARRYB[20][21] ), .SUM(\mult_26/SUMB[20][21] ) );
  FADDER \mult_26/S2_20_20  ( .CIN(\mult_26/ab[20][20] ), .IN0(
        \mult_26/CARRYB[19][20] ), .IN1(\mult_26/SUMB[19][21] ), .COUT(
        \mult_26/CARRYB[20][20] ), .SUM(\mult_26/SUMB[20][20] ) );
  FADDER \mult_26/S2_20_19  ( .CIN(\mult_26/ab[20][19] ), .IN0(
        \mult_26/CARRYB[19][19] ), .IN1(\mult_26/SUMB[19][20] ), .COUT(
        \mult_26/CARRYB[20][19] ), .SUM(\mult_26/SUMB[20][19] ) );
  FADDER \mult_26/S2_20_18  ( .CIN(\mult_26/ab[20][18] ), .IN0(
        \mult_26/CARRYB[19][18] ), .IN1(\mult_26/SUMB[19][19] ), .COUT(
        \mult_26/CARRYB[20][18] ), .SUM(\mult_26/SUMB[20][18] ) );
  FADDER \mult_26/S2_20_17  ( .CIN(\mult_26/ab[20][17] ), .IN0(
        \mult_26/CARRYB[19][17] ), .IN1(\mult_26/SUMB[19][18] ), .COUT(
        \mult_26/CARRYB[20][17] ), .SUM(\mult_26/SUMB[20][17] ) );
  FADDER \mult_26/S2_20_16  ( .CIN(\mult_26/ab[20][16] ), .IN0(
        \mult_26/CARRYB[19][16] ), .IN1(\mult_26/SUMB[19][17] ), .COUT(
        \mult_26/CARRYB[20][16] ), .SUM(\mult_26/SUMB[20][16] ) );
  FADDER \mult_26/S2_20_15  ( .CIN(\mult_26/ab[20][15] ), .IN0(
        \mult_26/CARRYB[19][15] ), .IN1(\mult_26/SUMB[19][16] ), .COUT(
        \mult_26/CARRYB[20][15] ), .SUM(\mult_26/SUMB[20][15] ) );
  FADDER \mult_26/S2_20_14  ( .CIN(\mult_26/ab[20][14] ), .IN0(
        \mult_26/CARRYB[19][14] ), .IN1(\mult_26/SUMB[19][15] ), .COUT(
        \mult_26/CARRYB[20][14] ), .SUM(\mult_26/SUMB[20][14] ) );
  FADDER \mult_26/S2_20_13  ( .CIN(\mult_26/ab[20][13] ), .IN0(
        \mult_26/CARRYB[19][13] ), .IN1(\mult_26/SUMB[19][14] ), .COUT(
        \mult_26/CARRYB[20][13] ), .SUM(\mult_26/SUMB[20][13] ) );
  FADDER \mult_26/S2_20_12  ( .CIN(\mult_26/ab[20][12] ), .IN0(
        \mult_26/CARRYB[19][12] ), .IN1(\mult_26/SUMB[19][13] ), .COUT(
        \mult_26/CARRYB[20][12] ), .SUM(\mult_26/SUMB[20][12] ) );
  FADDER \mult_26/S2_20_11  ( .CIN(\mult_26/ab[20][11] ), .IN0(
        \mult_26/CARRYB[19][11] ), .IN1(\mult_26/SUMB[19][12] ), .COUT(
        \mult_26/CARRYB[20][11] ), .SUM(\mult_26/SUMB[20][11] ) );
  FADDER \mult_26/S2_20_10  ( .CIN(\mult_26/ab[20][10] ), .IN0(
        \mult_26/CARRYB[19][10] ), .IN1(\mult_26/SUMB[19][11] ), .COUT(
        \mult_26/CARRYB[20][10] ), .SUM(\mult_26/SUMB[20][10] ) );
  FADDER \mult_26/S2_20_9  ( .CIN(\mult_26/ab[20][9] ), .IN0(
        \mult_26/CARRYB[19][9] ), .IN1(\mult_26/SUMB[19][10] ), .COUT(
        \mult_26/CARRYB[20][9] ), .SUM(\mult_26/SUMB[20][9] ) );
  FADDER \mult_26/S2_20_8  ( .CIN(\mult_26/ab[20][8] ), .IN0(
        \mult_26/CARRYB[19][8] ), .IN1(\mult_26/SUMB[19][9] ), .COUT(
        \mult_26/CARRYB[20][8] ), .SUM(\mult_26/SUMB[20][8] ) );
  FADDER \mult_26/S2_20_7  ( .CIN(\mult_26/ab[20][7] ), .IN0(
        \mult_26/CARRYB[19][7] ), .IN1(\mult_26/SUMB[19][8] ), .COUT(
        \mult_26/CARRYB[20][7] ), .SUM(\mult_26/SUMB[20][7] ) );
  FADDER \mult_26/S2_20_6  ( .CIN(\mult_26/ab[20][6] ), .IN0(
        \mult_26/CARRYB[19][6] ), .IN1(\mult_26/SUMB[19][7] ), .COUT(
        \mult_26/CARRYB[20][6] ), .SUM(\mult_26/SUMB[20][6] ) );
  FADDER \mult_26/S2_20_5  ( .CIN(\mult_26/ab[20][5] ), .IN0(
        \mult_26/CARRYB[19][5] ), .IN1(\mult_26/SUMB[19][6] ), .COUT(
        \mult_26/CARRYB[20][5] ), .SUM(\mult_26/SUMB[20][5] ) );
  FADDER \mult_26/S2_20_4  ( .CIN(\mult_26/ab[20][4] ), .IN0(
        \mult_26/CARRYB[19][4] ), .IN1(\mult_26/SUMB[19][5] ), .COUT(
        \mult_26/CARRYB[20][4] ), .SUM(\mult_26/SUMB[20][4] ) );
  FADDER \mult_26/S2_20_3  ( .CIN(\mult_26/ab[20][3] ), .IN0(
        \mult_26/CARRYB[19][3] ), .IN1(\mult_26/SUMB[19][4] ), .COUT(
        \mult_26/CARRYB[20][3] ), .SUM(\mult_26/SUMB[20][3] ) );
  FADDER \mult_26/S2_20_2  ( .CIN(\mult_26/ab[20][2] ), .IN0(
        \mult_26/CARRYB[19][2] ), .IN1(\mult_26/SUMB[19][3] ), .COUT(
        \mult_26/CARRYB[20][2] ), .SUM(\mult_26/SUMB[20][2] ) );
  FADDER \mult_26/S2_20_1  ( .CIN(\mult_26/ab[20][1] ), .IN0(
        \mult_26/CARRYB[19][1] ), .IN1(\mult_26/SUMB[19][2] ), .COUT(
        \mult_26/CARRYB[20][1] ), .SUM(\mult_26/SUMB[20][1] ) );
  FADDER \mult_26/S1_20_0  ( .CIN(\mult_26/ab[20][0] ), .IN0(
        \mult_26/CARRYB[19][0] ), .IN1(\mult_26/SUMB[19][1] ), .COUT(
        \mult_26/CARRYB[20][0] ), .SUM(o[20]) );
  FADDER \mult_26/S3_21_30  ( .CIN(\mult_26/ab[21][30] ), .IN0(
        \mult_26/CARRYB[20][30] ), .IN1(\mult_26/ab[20][31] ), .COUT(
        \mult_26/CARRYB[21][30] ), .SUM(\mult_26/SUMB[21][30] ) );
  FADDER \mult_26/S2_21_29  ( .CIN(\mult_26/ab[21][29] ), .IN0(
        \mult_26/CARRYB[20][29] ), .IN1(\mult_26/SUMB[20][30] ), .COUT(
        \mult_26/CARRYB[21][29] ), .SUM(\mult_26/SUMB[21][29] ) );
  FADDER \mult_26/S2_21_28  ( .CIN(\mult_26/ab[21][28] ), .IN0(
        \mult_26/CARRYB[20][28] ), .IN1(\mult_26/SUMB[20][29] ), .COUT(
        \mult_26/CARRYB[21][28] ), .SUM(\mult_26/SUMB[21][28] ) );
  FADDER \mult_26/S2_21_27  ( .CIN(\mult_26/ab[21][27] ), .IN0(
        \mult_26/CARRYB[20][27] ), .IN1(\mult_26/SUMB[20][28] ), .COUT(
        \mult_26/CARRYB[21][27] ), .SUM(\mult_26/SUMB[21][27] ) );
  FADDER \mult_26/S2_21_26  ( .CIN(\mult_26/ab[21][26] ), .IN0(
        \mult_26/CARRYB[20][26] ), .IN1(\mult_26/SUMB[20][27] ), .COUT(
        \mult_26/CARRYB[21][26] ), .SUM(\mult_26/SUMB[21][26] ) );
  FADDER \mult_26/S2_21_25  ( .CIN(\mult_26/ab[21][25] ), .IN0(
        \mult_26/CARRYB[20][25] ), .IN1(\mult_26/SUMB[20][26] ), .COUT(
        \mult_26/CARRYB[21][25] ), .SUM(\mult_26/SUMB[21][25] ) );
  FADDER \mult_26/S2_21_24  ( .CIN(\mult_26/ab[21][24] ), .IN0(
        \mult_26/CARRYB[20][24] ), .IN1(\mult_26/SUMB[20][25] ), .COUT(
        \mult_26/CARRYB[21][24] ), .SUM(\mult_26/SUMB[21][24] ) );
  FADDER \mult_26/S2_21_23  ( .CIN(\mult_26/ab[21][23] ), .IN0(
        \mult_26/CARRYB[20][23] ), .IN1(\mult_26/SUMB[20][24] ), .COUT(
        \mult_26/CARRYB[21][23] ), .SUM(\mult_26/SUMB[21][23] ) );
  FADDER \mult_26/S2_21_22  ( .CIN(\mult_26/ab[21][22] ), .IN0(
        \mult_26/CARRYB[20][22] ), .IN1(\mult_26/SUMB[20][23] ), .COUT(
        \mult_26/CARRYB[21][22] ), .SUM(\mult_26/SUMB[21][22] ) );
  FADDER \mult_26/S2_21_21  ( .CIN(\mult_26/ab[21][21] ), .IN0(
        \mult_26/CARRYB[20][21] ), .IN1(\mult_26/SUMB[20][22] ), .COUT(
        \mult_26/CARRYB[21][21] ), .SUM(\mult_26/SUMB[21][21] ) );
  FADDER \mult_26/S2_21_20  ( .CIN(\mult_26/ab[21][20] ), .IN0(
        \mult_26/CARRYB[20][20] ), .IN1(\mult_26/SUMB[20][21] ), .COUT(
        \mult_26/CARRYB[21][20] ), .SUM(\mult_26/SUMB[21][20] ) );
  FADDER \mult_26/S2_21_19  ( .CIN(\mult_26/ab[21][19] ), .IN0(
        \mult_26/CARRYB[20][19] ), .IN1(\mult_26/SUMB[20][20] ), .COUT(
        \mult_26/CARRYB[21][19] ), .SUM(\mult_26/SUMB[21][19] ) );
  FADDER \mult_26/S2_21_18  ( .CIN(\mult_26/ab[21][18] ), .IN0(
        \mult_26/CARRYB[20][18] ), .IN1(\mult_26/SUMB[20][19] ), .COUT(
        \mult_26/CARRYB[21][18] ), .SUM(\mult_26/SUMB[21][18] ) );
  FADDER \mult_26/S2_21_17  ( .CIN(\mult_26/ab[21][17] ), .IN0(
        \mult_26/CARRYB[20][17] ), .IN1(\mult_26/SUMB[20][18] ), .COUT(
        \mult_26/CARRYB[21][17] ), .SUM(\mult_26/SUMB[21][17] ) );
  FADDER \mult_26/S2_21_16  ( .CIN(\mult_26/ab[21][16] ), .IN0(
        \mult_26/CARRYB[20][16] ), .IN1(\mult_26/SUMB[20][17] ), .COUT(
        \mult_26/CARRYB[21][16] ), .SUM(\mult_26/SUMB[21][16] ) );
  FADDER \mult_26/S2_21_15  ( .CIN(\mult_26/ab[21][15] ), .IN0(
        \mult_26/CARRYB[20][15] ), .IN1(\mult_26/SUMB[20][16] ), .COUT(
        \mult_26/CARRYB[21][15] ), .SUM(\mult_26/SUMB[21][15] ) );
  FADDER \mult_26/S2_21_14  ( .CIN(\mult_26/ab[21][14] ), .IN0(
        \mult_26/CARRYB[20][14] ), .IN1(\mult_26/SUMB[20][15] ), .COUT(
        \mult_26/CARRYB[21][14] ), .SUM(\mult_26/SUMB[21][14] ) );
  FADDER \mult_26/S2_21_13  ( .CIN(\mult_26/ab[21][13] ), .IN0(
        \mult_26/CARRYB[20][13] ), .IN1(\mult_26/SUMB[20][14] ), .COUT(
        \mult_26/CARRYB[21][13] ), .SUM(\mult_26/SUMB[21][13] ) );
  FADDER \mult_26/S2_21_12  ( .CIN(\mult_26/ab[21][12] ), .IN0(
        \mult_26/CARRYB[20][12] ), .IN1(\mult_26/SUMB[20][13] ), .COUT(
        \mult_26/CARRYB[21][12] ), .SUM(\mult_26/SUMB[21][12] ) );
  FADDER \mult_26/S2_21_11  ( .CIN(\mult_26/ab[21][11] ), .IN0(
        \mult_26/CARRYB[20][11] ), .IN1(\mult_26/SUMB[20][12] ), .COUT(
        \mult_26/CARRYB[21][11] ), .SUM(\mult_26/SUMB[21][11] ) );
  FADDER \mult_26/S2_21_10  ( .CIN(\mult_26/ab[21][10] ), .IN0(
        \mult_26/CARRYB[20][10] ), .IN1(\mult_26/SUMB[20][11] ), .COUT(
        \mult_26/CARRYB[21][10] ), .SUM(\mult_26/SUMB[21][10] ) );
  FADDER \mult_26/S2_21_9  ( .CIN(\mult_26/ab[21][9] ), .IN0(
        \mult_26/CARRYB[20][9] ), .IN1(\mult_26/SUMB[20][10] ), .COUT(
        \mult_26/CARRYB[21][9] ), .SUM(\mult_26/SUMB[21][9] ) );
  FADDER \mult_26/S2_21_8  ( .CIN(\mult_26/ab[21][8] ), .IN0(
        \mult_26/CARRYB[20][8] ), .IN1(\mult_26/SUMB[20][9] ), .COUT(
        \mult_26/CARRYB[21][8] ), .SUM(\mult_26/SUMB[21][8] ) );
  FADDER \mult_26/S2_21_7  ( .CIN(\mult_26/ab[21][7] ), .IN0(
        \mult_26/CARRYB[20][7] ), .IN1(\mult_26/SUMB[20][8] ), .COUT(
        \mult_26/CARRYB[21][7] ), .SUM(\mult_26/SUMB[21][7] ) );
  FADDER \mult_26/S2_21_6  ( .CIN(\mult_26/ab[21][6] ), .IN0(
        \mult_26/CARRYB[20][6] ), .IN1(\mult_26/SUMB[20][7] ), .COUT(
        \mult_26/CARRYB[21][6] ), .SUM(\mult_26/SUMB[21][6] ) );
  FADDER \mult_26/S2_21_5  ( .CIN(\mult_26/ab[21][5] ), .IN0(
        \mult_26/CARRYB[20][5] ), .IN1(\mult_26/SUMB[20][6] ), .COUT(
        \mult_26/CARRYB[21][5] ), .SUM(\mult_26/SUMB[21][5] ) );
  FADDER \mult_26/S2_21_4  ( .CIN(\mult_26/ab[21][4] ), .IN0(
        \mult_26/CARRYB[20][4] ), .IN1(\mult_26/SUMB[20][5] ), .COUT(
        \mult_26/CARRYB[21][4] ), .SUM(\mult_26/SUMB[21][4] ) );
  FADDER \mult_26/S2_21_3  ( .CIN(\mult_26/ab[21][3] ), .IN0(
        \mult_26/CARRYB[20][3] ), .IN1(\mult_26/SUMB[20][4] ), .COUT(
        \mult_26/CARRYB[21][3] ), .SUM(\mult_26/SUMB[21][3] ) );
  FADDER \mult_26/S2_21_2  ( .CIN(\mult_26/ab[21][2] ), .IN0(
        \mult_26/CARRYB[20][2] ), .IN1(\mult_26/SUMB[20][3] ), .COUT(
        \mult_26/CARRYB[21][2] ), .SUM(\mult_26/SUMB[21][2] ) );
  FADDER \mult_26/S2_21_1  ( .CIN(\mult_26/ab[21][1] ), .IN0(
        \mult_26/CARRYB[20][1] ), .IN1(\mult_26/SUMB[20][2] ), .COUT(
        \mult_26/CARRYB[21][1] ), .SUM(\mult_26/SUMB[21][1] ) );
  FADDER \mult_26/S1_21_0  ( .CIN(\mult_26/ab[21][0] ), .IN0(
        \mult_26/CARRYB[20][0] ), .IN1(\mult_26/SUMB[20][1] ), .COUT(
        \mult_26/CARRYB[21][0] ), .SUM(o[21]) );
  FADDER \mult_26/S3_22_30  ( .CIN(\mult_26/ab[22][30] ), .IN0(
        \mult_26/CARRYB[21][30] ), .IN1(\mult_26/ab[21][31] ), .COUT(
        \mult_26/CARRYB[22][30] ), .SUM(\mult_26/SUMB[22][30] ) );
  FADDER \mult_26/S2_22_29  ( .CIN(\mult_26/ab[22][29] ), .IN0(
        \mult_26/CARRYB[21][29] ), .IN1(\mult_26/SUMB[21][30] ), .COUT(
        \mult_26/CARRYB[22][29] ), .SUM(\mult_26/SUMB[22][29] ) );
  FADDER \mult_26/S2_22_28  ( .CIN(\mult_26/ab[22][28] ), .IN0(
        \mult_26/CARRYB[21][28] ), .IN1(\mult_26/SUMB[21][29] ), .COUT(
        \mult_26/CARRYB[22][28] ), .SUM(\mult_26/SUMB[22][28] ) );
  FADDER \mult_26/S2_22_27  ( .CIN(\mult_26/ab[22][27] ), .IN0(
        \mult_26/CARRYB[21][27] ), .IN1(\mult_26/SUMB[21][28] ), .COUT(
        \mult_26/CARRYB[22][27] ), .SUM(\mult_26/SUMB[22][27] ) );
  FADDER \mult_26/S2_22_26  ( .CIN(\mult_26/ab[22][26] ), .IN0(
        \mult_26/CARRYB[21][26] ), .IN1(\mult_26/SUMB[21][27] ), .COUT(
        \mult_26/CARRYB[22][26] ), .SUM(\mult_26/SUMB[22][26] ) );
  FADDER \mult_26/S2_22_25  ( .CIN(\mult_26/ab[22][25] ), .IN0(
        \mult_26/CARRYB[21][25] ), .IN1(\mult_26/SUMB[21][26] ), .COUT(
        \mult_26/CARRYB[22][25] ), .SUM(\mult_26/SUMB[22][25] ) );
  FADDER \mult_26/S2_22_24  ( .CIN(\mult_26/ab[22][24] ), .IN0(
        \mult_26/CARRYB[21][24] ), .IN1(\mult_26/SUMB[21][25] ), .COUT(
        \mult_26/CARRYB[22][24] ), .SUM(\mult_26/SUMB[22][24] ) );
  FADDER \mult_26/S2_22_23  ( .CIN(\mult_26/ab[22][23] ), .IN0(
        \mult_26/CARRYB[21][23] ), .IN1(\mult_26/SUMB[21][24] ), .COUT(
        \mult_26/CARRYB[22][23] ), .SUM(\mult_26/SUMB[22][23] ) );
  FADDER \mult_26/S2_22_22  ( .CIN(\mult_26/ab[22][22] ), .IN0(
        \mult_26/CARRYB[21][22] ), .IN1(\mult_26/SUMB[21][23] ), .COUT(
        \mult_26/CARRYB[22][22] ), .SUM(\mult_26/SUMB[22][22] ) );
  FADDER \mult_26/S2_22_21  ( .CIN(\mult_26/ab[22][21] ), .IN0(
        \mult_26/CARRYB[21][21] ), .IN1(\mult_26/SUMB[21][22] ), .COUT(
        \mult_26/CARRYB[22][21] ), .SUM(\mult_26/SUMB[22][21] ) );
  FADDER \mult_26/S2_22_20  ( .CIN(\mult_26/ab[22][20] ), .IN0(
        \mult_26/CARRYB[21][20] ), .IN1(\mult_26/SUMB[21][21] ), .COUT(
        \mult_26/CARRYB[22][20] ), .SUM(\mult_26/SUMB[22][20] ) );
  FADDER \mult_26/S2_22_19  ( .CIN(\mult_26/ab[22][19] ), .IN0(
        \mult_26/CARRYB[21][19] ), .IN1(\mult_26/SUMB[21][20] ), .COUT(
        \mult_26/CARRYB[22][19] ), .SUM(\mult_26/SUMB[22][19] ) );
  FADDER \mult_26/S2_22_18  ( .CIN(\mult_26/ab[22][18] ), .IN0(
        \mult_26/CARRYB[21][18] ), .IN1(\mult_26/SUMB[21][19] ), .COUT(
        \mult_26/CARRYB[22][18] ), .SUM(\mult_26/SUMB[22][18] ) );
  FADDER \mult_26/S2_22_17  ( .CIN(\mult_26/ab[22][17] ), .IN0(
        \mult_26/CARRYB[21][17] ), .IN1(\mult_26/SUMB[21][18] ), .COUT(
        \mult_26/CARRYB[22][17] ), .SUM(\mult_26/SUMB[22][17] ) );
  FADDER \mult_26/S2_22_16  ( .CIN(\mult_26/ab[22][16] ), .IN0(
        \mult_26/CARRYB[21][16] ), .IN1(\mult_26/SUMB[21][17] ), .COUT(
        \mult_26/CARRYB[22][16] ), .SUM(\mult_26/SUMB[22][16] ) );
  FADDER \mult_26/S2_22_15  ( .CIN(\mult_26/ab[22][15] ), .IN0(
        \mult_26/CARRYB[21][15] ), .IN1(\mult_26/SUMB[21][16] ), .COUT(
        \mult_26/CARRYB[22][15] ), .SUM(\mult_26/SUMB[22][15] ) );
  FADDER \mult_26/S2_22_14  ( .CIN(\mult_26/ab[22][14] ), .IN0(
        \mult_26/CARRYB[21][14] ), .IN1(\mult_26/SUMB[21][15] ), .COUT(
        \mult_26/CARRYB[22][14] ), .SUM(\mult_26/SUMB[22][14] ) );
  FADDER \mult_26/S2_22_13  ( .CIN(\mult_26/ab[22][13] ), .IN0(
        \mult_26/CARRYB[21][13] ), .IN1(\mult_26/SUMB[21][14] ), .COUT(
        \mult_26/CARRYB[22][13] ), .SUM(\mult_26/SUMB[22][13] ) );
  FADDER \mult_26/S2_22_12  ( .CIN(\mult_26/ab[22][12] ), .IN0(
        \mult_26/CARRYB[21][12] ), .IN1(\mult_26/SUMB[21][13] ), .COUT(
        \mult_26/CARRYB[22][12] ), .SUM(\mult_26/SUMB[22][12] ) );
  FADDER \mult_26/S2_22_11  ( .CIN(\mult_26/ab[22][11] ), .IN0(
        \mult_26/CARRYB[21][11] ), .IN1(\mult_26/SUMB[21][12] ), .COUT(
        \mult_26/CARRYB[22][11] ), .SUM(\mult_26/SUMB[22][11] ) );
  FADDER \mult_26/S2_22_10  ( .CIN(\mult_26/ab[22][10] ), .IN0(
        \mult_26/CARRYB[21][10] ), .IN1(\mult_26/SUMB[21][11] ), .COUT(
        \mult_26/CARRYB[22][10] ), .SUM(\mult_26/SUMB[22][10] ) );
  FADDER \mult_26/S2_22_9  ( .CIN(\mult_26/ab[22][9] ), .IN0(
        \mult_26/CARRYB[21][9] ), .IN1(\mult_26/SUMB[21][10] ), .COUT(
        \mult_26/CARRYB[22][9] ), .SUM(\mult_26/SUMB[22][9] ) );
  FADDER \mult_26/S2_22_8  ( .CIN(\mult_26/ab[22][8] ), .IN0(
        \mult_26/CARRYB[21][8] ), .IN1(\mult_26/SUMB[21][9] ), .COUT(
        \mult_26/CARRYB[22][8] ), .SUM(\mult_26/SUMB[22][8] ) );
  FADDER \mult_26/S2_22_7  ( .CIN(\mult_26/ab[22][7] ), .IN0(
        \mult_26/CARRYB[21][7] ), .IN1(\mult_26/SUMB[21][8] ), .COUT(
        \mult_26/CARRYB[22][7] ), .SUM(\mult_26/SUMB[22][7] ) );
  FADDER \mult_26/S2_22_6  ( .CIN(\mult_26/ab[22][6] ), .IN0(
        \mult_26/CARRYB[21][6] ), .IN1(\mult_26/SUMB[21][7] ), .COUT(
        \mult_26/CARRYB[22][6] ), .SUM(\mult_26/SUMB[22][6] ) );
  FADDER \mult_26/S2_22_5  ( .CIN(\mult_26/ab[22][5] ), .IN0(
        \mult_26/CARRYB[21][5] ), .IN1(\mult_26/SUMB[21][6] ), .COUT(
        \mult_26/CARRYB[22][5] ), .SUM(\mult_26/SUMB[22][5] ) );
  FADDER \mult_26/S2_22_4  ( .CIN(\mult_26/ab[22][4] ), .IN0(
        \mult_26/CARRYB[21][4] ), .IN1(\mult_26/SUMB[21][5] ), .COUT(
        \mult_26/CARRYB[22][4] ), .SUM(\mult_26/SUMB[22][4] ) );
  FADDER \mult_26/S2_22_3  ( .CIN(\mult_26/ab[22][3] ), .IN0(
        \mult_26/CARRYB[21][3] ), .IN1(\mult_26/SUMB[21][4] ), .COUT(
        \mult_26/CARRYB[22][3] ), .SUM(\mult_26/SUMB[22][3] ) );
  FADDER \mult_26/S2_22_2  ( .CIN(\mult_26/ab[22][2] ), .IN0(
        \mult_26/CARRYB[21][2] ), .IN1(\mult_26/SUMB[21][3] ), .COUT(
        \mult_26/CARRYB[22][2] ), .SUM(\mult_26/SUMB[22][2] ) );
  FADDER \mult_26/S2_22_1  ( .CIN(\mult_26/ab[22][1] ), .IN0(
        \mult_26/CARRYB[21][1] ), .IN1(\mult_26/SUMB[21][2] ), .COUT(
        \mult_26/CARRYB[22][1] ), .SUM(\mult_26/SUMB[22][1] ) );
  FADDER \mult_26/S1_22_0  ( .CIN(\mult_26/ab[22][0] ), .IN0(
        \mult_26/CARRYB[21][0] ), .IN1(\mult_26/SUMB[21][1] ), .COUT(
        \mult_26/CARRYB[22][0] ), .SUM(o[22]) );
  FADDER \mult_26/S3_23_30  ( .CIN(\mult_26/ab[23][30] ), .IN0(
        \mult_26/CARRYB[22][30] ), .IN1(\mult_26/ab[22][31] ), .COUT(
        \mult_26/CARRYB[23][30] ), .SUM(\mult_26/SUMB[23][30] ) );
  FADDER \mult_26/S2_23_29  ( .CIN(\mult_26/ab[23][29] ), .IN0(
        \mult_26/CARRYB[22][29] ), .IN1(\mult_26/SUMB[22][30] ), .COUT(
        \mult_26/CARRYB[23][29] ), .SUM(\mult_26/SUMB[23][29] ) );
  FADDER \mult_26/S2_23_28  ( .CIN(\mult_26/ab[23][28] ), .IN0(
        \mult_26/CARRYB[22][28] ), .IN1(\mult_26/SUMB[22][29] ), .COUT(
        \mult_26/CARRYB[23][28] ), .SUM(\mult_26/SUMB[23][28] ) );
  FADDER \mult_26/S2_23_27  ( .CIN(\mult_26/ab[23][27] ), .IN0(
        \mult_26/CARRYB[22][27] ), .IN1(\mult_26/SUMB[22][28] ), .COUT(
        \mult_26/CARRYB[23][27] ), .SUM(\mult_26/SUMB[23][27] ) );
  FADDER \mult_26/S2_23_26  ( .CIN(\mult_26/ab[23][26] ), .IN0(
        \mult_26/CARRYB[22][26] ), .IN1(\mult_26/SUMB[22][27] ), .COUT(
        \mult_26/CARRYB[23][26] ), .SUM(\mult_26/SUMB[23][26] ) );
  FADDER \mult_26/S2_23_25  ( .CIN(\mult_26/ab[23][25] ), .IN0(
        \mult_26/CARRYB[22][25] ), .IN1(\mult_26/SUMB[22][26] ), .COUT(
        \mult_26/CARRYB[23][25] ), .SUM(\mult_26/SUMB[23][25] ) );
  FADDER \mult_26/S2_23_24  ( .CIN(\mult_26/ab[23][24] ), .IN0(
        \mult_26/CARRYB[22][24] ), .IN1(\mult_26/SUMB[22][25] ), .COUT(
        \mult_26/CARRYB[23][24] ), .SUM(\mult_26/SUMB[23][24] ) );
  FADDER \mult_26/S2_23_23  ( .CIN(\mult_26/ab[23][23] ), .IN0(
        \mult_26/CARRYB[22][23] ), .IN1(\mult_26/SUMB[22][24] ), .COUT(
        \mult_26/CARRYB[23][23] ), .SUM(\mult_26/SUMB[23][23] ) );
  FADDER \mult_26/S2_23_22  ( .CIN(\mult_26/ab[23][22] ), .IN0(
        \mult_26/CARRYB[22][22] ), .IN1(\mult_26/SUMB[22][23] ), .COUT(
        \mult_26/CARRYB[23][22] ), .SUM(\mult_26/SUMB[23][22] ) );
  FADDER \mult_26/S2_23_21  ( .CIN(\mult_26/ab[23][21] ), .IN0(
        \mult_26/CARRYB[22][21] ), .IN1(\mult_26/SUMB[22][22] ), .COUT(
        \mult_26/CARRYB[23][21] ), .SUM(\mult_26/SUMB[23][21] ) );
  FADDER \mult_26/S2_23_20  ( .CIN(\mult_26/ab[23][20] ), .IN0(
        \mult_26/CARRYB[22][20] ), .IN1(\mult_26/SUMB[22][21] ), .COUT(
        \mult_26/CARRYB[23][20] ), .SUM(\mult_26/SUMB[23][20] ) );
  FADDER \mult_26/S2_23_19  ( .CIN(\mult_26/ab[23][19] ), .IN0(
        \mult_26/CARRYB[22][19] ), .IN1(\mult_26/SUMB[22][20] ), .COUT(
        \mult_26/CARRYB[23][19] ), .SUM(\mult_26/SUMB[23][19] ) );
  FADDER \mult_26/S2_23_18  ( .CIN(\mult_26/ab[23][18] ), .IN0(
        \mult_26/CARRYB[22][18] ), .IN1(\mult_26/SUMB[22][19] ), .COUT(
        \mult_26/CARRYB[23][18] ), .SUM(\mult_26/SUMB[23][18] ) );
  FADDER \mult_26/S2_23_17  ( .CIN(\mult_26/ab[23][17] ), .IN0(
        \mult_26/CARRYB[22][17] ), .IN1(\mult_26/SUMB[22][18] ), .COUT(
        \mult_26/CARRYB[23][17] ), .SUM(\mult_26/SUMB[23][17] ) );
  FADDER \mult_26/S2_23_16  ( .CIN(\mult_26/ab[23][16] ), .IN0(
        \mult_26/CARRYB[22][16] ), .IN1(\mult_26/SUMB[22][17] ), .COUT(
        \mult_26/CARRYB[23][16] ), .SUM(\mult_26/SUMB[23][16] ) );
  FADDER \mult_26/S2_23_15  ( .CIN(\mult_26/ab[23][15] ), .IN0(
        \mult_26/CARRYB[22][15] ), .IN1(\mult_26/SUMB[22][16] ), .COUT(
        \mult_26/CARRYB[23][15] ), .SUM(\mult_26/SUMB[23][15] ) );
  FADDER \mult_26/S2_23_14  ( .CIN(\mult_26/ab[23][14] ), .IN0(
        \mult_26/CARRYB[22][14] ), .IN1(\mult_26/SUMB[22][15] ), .COUT(
        \mult_26/CARRYB[23][14] ), .SUM(\mult_26/SUMB[23][14] ) );
  FADDER \mult_26/S2_23_13  ( .CIN(\mult_26/ab[23][13] ), .IN0(
        \mult_26/CARRYB[22][13] ), .IN1(\mult_26/SUMB[22][14] ), .COUT(
        \mult_26/CARRYB[23][13] ), .SUM(\mult_26/SUMB[23][13] ) );
  FADDER \mult_26/S2_23_12  ( .CIN(\mult_26/ab[23][12] ), .IN0(
        \mult_26/CARRYB[22][12] ), .IN1(\mult_26/SUMB[22][13] ), .COUT(
        \mult_26/CARRYB[23][12] ), .SUM(\mult_26/SUMB[23][12] ) );
  FADDER \mult_26/S2_23_11  ( .CIN(\mult_26/ab[23][11] ), .IN0(
        \mult_26/CARRYB[22][11] ), .IN1(\mult_26/SUMB[22][12] ), .COUT(
        \mult_26/CARRYB[23][11] ), .SUM(\mult_26/SUMB[23][11] ) );
  FADDER \mult_26/S2_23_10  ( .CIN(\mult_26/ab[23][10] ), .IN0(
        \mult_26/CARRYB[22][10] ), .IN1(\mult_26/SUMB[22][11] ), .COUT(
        \mult_26/CARRYB[23][10] ), .SUM(\mult_26/SUMB[23][10] ) );
  FADDER \mult_26/S2_23_9  ( .CIN(\mult_26/ab[23][9] ), .IN0(
        \mult_26/CARRYB[22][9] ), .IN1(\mult_26/SUMB[22][10] ), .COUT(
        \mult_26/CARRYB[23][9] ), .SUM(\mult_26/SUMB[23][9] ) );
  FADDER \mult_26/S2_23_8  ( .CIN(\mult_26/ab[23][8] ), .IN0(
        \mult_26/CARRYB[22][8] ), .IN1(\mult_26/SUMB[22][9] ), .COUT(
        \mult_26/CARRYB[23][8] ), .SUM(\mult_26/SUMB[23][8] ) );
  FADDER \mult_26/S2_23_7  ( .CIN(\mult_26/ab[23][7] ), .IN0(
        \mult_26/CARRYB[22][7] ), .IN1(\mult_26/SUMB[22][8] ), .COUT(
        \mult_26/CARRYB[23][7] ), .SUM(\mult_26/SUMB[23][7] ) );
  FADDER \mult_26/S2_23_6  ( .CIN(\mult_26/ab[23][6] ), .IN0(
        \mult_26/CARRYB[22][6] ), .IN1(\mult_26/SUMB[22][7] ), .COUT(
        \mult_26/CARRYB[23][6] ), .SUM(\mult_26/SUMB[23][6] ) );
  FADDER \mult_26/S2_23_5  ( .CIN(\mult_26/ab[23][5] ), .IN0(
        \mult_26/CARRYB[22][5] ), .IN1(\mult_26/SUMB[22][6] ), .COUT(
        \mult_26/CARRYB[23][5] ), .SUM(\mult_26/SUMB[23][5] ) );
  FADDER \mult_26/S2_23_4  ( .CIN(\mult_26/ab[23][4] ), .IN0(
        \mult_26/CARRYB[22][4] ), .IN1(\mult_26/SUMB[22][5] ), .COUT(
        \mult_26/CARRYB[23][4] ), .SUM(\mult_26/SUMB[23][4] ) );
  FADDER \mult_26/S2_23_3  ( .CIN(\mult_26/ab[23][3] ), .IN0(
        \mult_26/CARRYB[22][3] ), .IN1(\mult_26/SUMB[22][4] ), .COUT(
        \mult_26/CARRYB[23][3] ), .SUM(\mult_26/SUMB[23][3] ) );
  FADDER \mult_26/S2_23_2  ( .CIN(\mult_26/ab[23][2] ), .IN0(
        \mult_26/CARRYB[22][2] ), .IN1(\mult_26/SUMB[22][3] ), .COUT(
        \mult_26/CARRYB[23][2] ), .SUM(\mult_26/SUMB[23][2] ) );
  FADDER \mult_26/S2_23_1  ( .CIN(\mult_26/ab[23][1] ), .IN0(
        \mult_26/CARRYB[22][1] ), .IN1(\mult_26/SUMB[22][2] ), .COUT(
        \mult_26/CARRYB[23][1] ), .SUM(\mult_26/SUMB[23][1] ) );
  FADDER \mult_26/S1_23_0  ( .CIN(\mult_26/ab[23][0] ), .IN0(
        \mult_26/CARRYB[22][0] ), .IN1(\mult_26/SUMB[22][1] ), .COUT(
        \mult_26/CARRYB[23][0] ), .SUM(o[23]) );
  FADDER \mult_26/S3_24_30  ( .CIN(\mult_26/ab[24][30] ), .IN0(
        \mult_26/CARRYB[23][30] ), .IN1(\mult_26/ab[23][31] ), .COUT(
        \mult_26/CARRYB[24][30] ), .SUM(\mult_26/SUMB[24][30] ) );
  FADDER \mult_26/S2_24_29  ( .CIN(\mult_26/ab[24][29] ), .IN0(
        \mult_26/CARRYB[23][29] ), .IN1(\mult_26/SUMB[23][30] ), .COUT(
        \mult_26/CARRYB[24][29] ), .SUM(\mult_26/SUMB[24][29] ) );
  FADDER \mult_26/S2_24_28  ( .CIN(\mult_26/ab[24][28] ), .IN0(
        \mult_26/CARRYB[23][28] ), .IN1(\mult_26/SUMB[23][29] ), .COUT(
        \mult_26/CARRYB[24][28] ), .SUM(\mult_26/SUMB[24][28] ) );
  FADDER \mult_26/S2_24_27  ( .CIN(\mult_26/ab[24][27] ), .IN0(
        \mult_26/CARRYB[23][27] ), .IN1(\mult_26/SUMB[23][28] ), .COUT(
        \mult_26/CARRYB[24][27] ), .SUM(\mult_26/SUMB[24][27] ) );
  FADDER \mult_26/S2_24_26  ( .CIN(\mult_26/ab[24][26] ), .IN0(
        \mult_26/CARRYB[23][26] ), .IN1(\mult_26/SUMB[23][27] ), .COUT(
        \mult_26/CARRYB[24][26] ), .SUM(\mult_26/SUMB[24][26] ) );
  FADDER \mult_26/S2_24_25  ( .CIN(\mult_26/ab[24][25] ), .IN0(
        \mult_26/CARRYB[23][25] ), .IN1(\mult_26/SUMB[23][26] ), .COUT(
        \mult_26/CARRYB[24][25] ), .SUM(\mult_26/SUMB[24][25] ) );
  FADDER \mult_26/S2_24_24  ( .CIN(\mult_26/ab[24][24] ), .IN0(
        \mult_26/CARRYB[23][24] ), .IN1(\mult_26/SUMB[23][25] ), .COUT(
        \mult_26/CARRYB[24][24] ), .SUM(\mult_26/SUMB[24][24] ) );
  FADDER \mult_26/S2_24_23  ( .CIN(\mult_26/ab[24][23] ), .IN0(
        \mult_26/CARRYB[23][23] ), .IN1(\mult_26/SUMB[23][24] ), .COUT(
        \mult_26/CARRYB[24][23] ), .SUM(\mult_26/SUMB[24][23] ) );
  FADDER \mult_26/S2_24_22  ( .CIN(\mult_26/ab[24][22] ), .IN0(
        \mult_26/CARRYB[23][22] ), .IN1(\mult_26/SUMB[23][23] ), .COUT(
        \mult_26/CARRYB[24][22] ), .SUM(\mult_26/SUMB[24][22] ) );
  FADDER \mult_26/S2_24_21  ( .CIN(\mult_26/ab[24][21] ), .IN0(
        \mult_26/CARRYB[23][21] ), .IN1(\mult_26/SUMB[23][22] ), .COUT(
        \mult_26/CARRYB[24][21] ), .SUM(\mult_26/SUMB[24][21] ) );
  FADDER \mult_26/S2_24_20  ( .CIN(\mult_26/ab[24][20] ), .IN0(
        \mult_26/CARRYB[23][20] ), .IN1(\mult_26/SUMB[23][21] ), .COUT(
        \mult_26/CARRYB[24][20] ), .SUM(\mult_26/SUMB[24][20] ) );
  FADDER \mult_26/S2_24_19  ( .CIN(\mult_26/ab[24][19] ), .IN0(
        \mult_26/CARRYB[23][19] ), .IN1(\mult_26/SUMB[23][20] ), .COUT(
        \mult_26/CARRYB[24][19] ), .SUM(\mult_26/SUMB[24][19] ) );
  FADDER \mult_26/S2_24_18  ( .CIN(\mult_26/ab[24][18] ), .IN0(
        \mult_26/CARRYB[23][18] ), .IN1(\mult_26/SUMB[23][19] ), .COUT(
        \mult_26/CARRYB[24][18] ), .SUM(\mult_26/SUMB[24][18] ) );
  FADDER \mult_26/S2_24_17  ( .CIN(\mult_26/ab[24][17] ), .IN0(
        \mult_26/CARRYB[23][17] ), .IN1(\mult_26/SUMB[23][18] ), .COUT(
        \mult_26/CARRYB[24][17] ), .SUM(\mult_26/SUMB[24][17] ) );
  FADDER \mult_26/S2_24_16  ( .CIN(\mult_26/ab[24][16] ), .IN0(
        \mult_26/CARRYB[23][16] ), .IN1(\mult_26/SUMB[23][17] ), .COUT(
        \mult_26/CARRYB[24][16] ), .SUM(\mult_26/SUMB[24][16] ) );
  FADDER \mult_26/S2_24_15  ( .CIN(\mult_26/ab[24][15] ), .IN0(
        \mult_26/CARRYB[23][15] ), .IN1(\mult_26/SUMB[23][16] ), .COUT(
        \mult_26/CARRYB[24][15] ), .SUM(\mult_26/SUMB[24][15] ) );
  FADDER \mult_26/S2_24_14  ( .CIN(\mult_26/ab[24][14] ), .IN0(
        \mult_26/CARRYB[23][14] ), .IN1(\mult_26/SUMB[23][15] ), .COUT(
        \mult_26/CARRYB[24][14] ), .SUM(\mult_26/SUMB[24][14] ) );
  FADDER \mult_26/S2_24_13  ( .CIN(\mult_26/ab[24][13] ), .IN0(
        \mult_26/CARRYB[23][13] ), .IN1(\mult_26/SUMB[23][14] ), .COUT(
        \mult_26/CARRYB[24][13] ), .SUM(\mult_26/SUMB[24][13] ) );
  FADDER \mult_26/S2_24_12  ( .CIN(\mult_26/ab[24][12] ), .IN0(
        \mult_26/CARRYB[23][12] ), .IN1(\mult_26/SUMB[23][13] ), .COUT(
        \mult_26/CARRYB[24][12] ), .SUM(\mult_26/SUMB[24][12] ) );
  FADDER \mult_26/S2_24_11  ( .CIN(\mult_26/ab[24][11] ), .IN0(
        \mult_26/CARRYB[23][11] ), .IN1(\mult_26/SUMB[23][12] ), .COUT(
        \mult_26/CARRYB[24][11] ), .SUM(\mult_26/SUMB[24][11] ) );
  FADDER \mult_26/S2_24_10  ( .CIN(\mult_26/ab[24][10] ), .IN0(
        \mult_26/CARRYB[23][10] ), .IN1(\mult_26/SUMB[23][11] ), .COUT(
        \mult_26/CARRYB[24][10] ), .SUM(\mult_26/SUMB[24][10] ) );
  FADDER \mult_26/S2_24_9  ( .CIN(\mult_26/ab[24][9] ), .IN0(
        \mult_26/CARRYB[23][9] ), .IN1(\mult_26/SUMB[23][10] ), .COUT(
        \mult_26/CARRYB[24][9] ), .SUM(\mult_26/SUMB[24][9] ) );
  FADDER \mult_26/S2_24_8  ( .CIN(\mult_26/ab[24][8] ), .IN0(
        \mult_26/CARRYB[23][8] ), .IN1(\mult_26/SUMB[23][9] ), .COUT(
        \mult_26/CARRYB[24][8] ), .SUM(\mult_26/SUMB[24][8] ) );
  FADDER \mult_26/S2_24_7  ( .CIN(\mult_26/ab[24][7] ), .IN0(
        \mult_26/CARRYB[23][7] ), .IN1(\mult_26/SUMB[23][8] ), .COUT(
        \mult_26/CARRYB[24][7] ), .SUM(\mult_26/SUMB[24][7] ) );
  FADDER \mult_26/S2_24_6  ( .CIN(\mult_26/ab[24][6] ), .IN0(
        \mult_26/CARRYB[23][6] ), .IN1(\mult_26/SUMB[23][7] ), .COUT(
        \mult_26/CARRYB[24][6] ), .SUM(\mult_26/SUMB[24][6] ) );
  FADDER \mult_26/S2_24_5  ( .CIN(\mult_26/ab[24][5] ), .IN0(
        \mult_26/CARRYB[23][5] ), .IN1(\mult_26/SUMB[23][6] ), .COUT(
        \mult_26/CARRYB[24][5] ), .SUM(\mult_26/SUMB[24][5] ) );
  FADDER \mult_26/S2_24_4  ( .CIN(\mult_26/ab[24][4] ), .IN0(
        \mult_26/CARRYB[23][4] ), .IN1(\mult_26/SUMB[23][5] ), .COUT(
        \mult_26/CARRYB[24][4] ), .SUM(\mult_26/SUMB[24][4] ) );
  FADDER \mult_26/S2_24_3  ( .CIN(\mult_26/ab[24][3] ), .IN0(
        \mult_26/CARRYB[23][3] ), .IN1(\mult_26/SUMB[23][4] ), .COUT(
        \mult_26/CARRYB[24][3] ), .SUM(\mult_26/SUMB[24][3] ) );
  FADDER \mult_26/S2_24_2  ( .CIN(\mult_26/ab[24][2] ), .IN0(
        \mult_26/CARRYB[23][2] ), .IN1(\mult_26/SUMB[23][3] ), .COUT(
        \mult_26/CARRYB[24][2] ), .SUM(\mult_26/SUMB[24][2] ) );
  FADDER \mult_26/S2_24_1  ( .CIN(\mult_26/ab[24][1] ), .IN0(
        \mult_26/CARRYB[23][1] ), .IN1(\mult_26/SUMB[23][2] ), .COUT(
        \mult_26/CARRYB[24][1] ), .SUM(\mult_26/SUMB[24][1] ) );
  FADDER \mult_26/S1_24_0  ( .CIN(\mult_26/ab[24][0] ), .IN0(
        \mult_26/CARRYB[23][0] ), .IN1(\mult_26/SUMB[23][1] ), .COUT(
        \mult_26/CARRYB[24][0] ), .SUM(o[24]) );
  FADDER \mult_26/S3_25_30  ( .CIN(\mult_26/ab[25][30] ), .IN0(
        \mult_26/CARRYB[24][30] ), .IN1(\mult_26/ab[24][31] ), .COUT(
        \mult_26/CARRYB[25][30] ), .SUM(\mult_26/SUMB[25][30] ) );
  FADDER \mult_26/S2_25_29  ( .CIN(\mult_26/ab[25][29] ), .IN0(
        \mult_26/CARRYB[24][29] ), .IN1(\mult_26/SUMB[24][30] ), .COUT(
        \mult_26/CARRYB[25][29] ), .SUM(\mult_26/SUMB[25][29] ) );
  FADDER \mult_26/S2_25_28  ( .CIN(\mult_26/ab[25][28] ), .IN0(
        \mult_26/CARRYB[24][28] ), .IN1(\mult_26/SUMB[24][29] ), .COUT(
        \mult_26/CARRYB[25][28] ), .SUM(\mult_26/SUMB[25][28] ) );
  FADDER \mult_26/S2_25_27  ( .CIN(\mult_26/ab[25][27] ), .IN0(
        \mult_26/CARRYB[24][27] ), .IN1(\mult_26/SUMB[24][28] ), .COUT(
        \mult_26/CARRYB[25][27] ), .SUM(\mult_26/SUMB[25][27] ) );
  FADDER \mult_26/S2_25_26  ( .CIN(\mult_26/ab[25][26] ), .IN0(
        \mult_26/CARRYB[24][26] ), .IN1(\mult_26/SUMB[24][27] ), .COUT(
        \mult_26/CARRYB[25][26] ), .SUM(\mult_26/SUMB[25][26] ) );
  FADDER \mult_26/S2_25_25  ( .CIN(\mult_26/ab[25][25] ), .IN0(
        \mult_26/CARRYB[24][25] ), .IN1(\mult_26/SUMB[24][26] ), .COUT(
        \mult_26/CARRYB[25][25] ), .SUM(\mult_26/SUMB[25][25] ) );
  FADDER \mult_26/S2_25_24  ( .CIN(\mult_26/ab[25][24] ), .IN0(
        \mult_26/CARRYB[24][24] ), .IN1(\mult_26/SUMB[24][25] ), .COUT(
        \mult_26/CARRYB[25][24] ), .SUM(\mult_26/SUMB[25][24] ) );
  FADDER \mult_26/S2_25_23  ( .CIN(\mult_26/ab[25][23] ), .IN0(
        \mult_26/CARRYB[24][23] ), .IN1(\mult_26/SUMB[24][24] ), .COUT(
        \mult_26/CARRYB[25][23] ), .SUM(\mult_26/SUMB[25][23] ) );
  FADDER \mult_26/S2_25_22  ( .CIN(\mult_26/ab[25][22] ), .IN0(
        \mult_26/CARRYB[24][22] ), .IN1(\mult_26/SUMB[24][23] ), .COUT(
        \mult_26/CARRYB[25][22] ), .SUM(\mult_26/SUMB[25][22] ) );
  FADDER \mult_26/S2_25_21  ( .CIN(\mult_26/ab[25][21] ), .IN0(
        \mult_26/CARRYB[24][21] ), .IN1(\mult_26/SUMB[24][22] ), .COUT(
        \mult_26/CARRYB[25][21] ), .SUM(\mult_26/SUMB[25][21] ) );
  FADDER \mult_26/S2_25_20  ( .CIN(\mult_26/ab[25][20] ), .IN0(
        \mult_26/CARRYB[24][20] ), .IN1(\mult_26/SUMB[24][21] ), .COUT(
        \mult_26/CARRYB[25][20] ), .SUM(\mult_26/SUMB[25][20] ) );
  FADDER \mult_26/S2_25_19  ( .CIN(\mult_26/ab[25][19] ), .IN0(
        \mult_26/CARRYB[24][19] ), .IN1(\mult_26/SUMB[24][20] ), .COUT(
        \mult_26/CARRYB[25][19] ), .SUM(\mult_26/SUMB[25][19] ) );
  FADDER \mult_26/S2_25_18  ( .CIN(\mult_26/ab[25][18] ), .IN0(
        \mult_26/CARRYB[24][18] ), .IN1(\mult_26/SUMB[24][19] ), .COUT(
        \mult_26/CARRYB[25][18] ), .SUM(\mult_26/SUMB[25][18] ) );
  FADDER \mult_26/S2_25_17  ( .CIN(\mult_26/ab[25][17] ), .IN0(
        \mult_26/CARRYB[24][17] ), .IN1(\mult_26/SUMB[24][18] ), .COUT(
        \mult_26/CARRYB[25][17] ), .SUM(\mult_26/SUMB[25][17] ) );
  FADDER \mult_26/S2_25_16  ( .CIN(\mult_26/ab[25][16] ), .IN0(
        \mult_26/CARRYB[24][16] ), .IN1(\mult_26/SUMB[24][17] ), .COUT(
        \mult_26/CARRYB[25][16] ), .SUM(\mult_26/SUMB[25][16] ) );
  FADDER \mult_26/S2_25_15  ( .CIN(\mult_26/ab[25][15] ), .IN0(
        \mult_26/CARRYB[24][15] ), .IN1(\mult_26/SUMB[24][16] ), .COUT(
        \mult_26/CARRYB[25][15] ), .SUM(\mult_26/SUMB[25][15] ) );
  FADDER \mult_26/S2_25_14  ( .CIN(\mult_26/ab[25][14] ), .IN0(
        \mult_26/CARRYB[24][14] ), .IN1(\mult_26/SUMB[24][15] ), .COUT(
        \mult_26/CARRYB[25][14] ), .SUM(\mult_26/SUMB[25][14] ) );
  FADDER \mult_26/S2_25_13  ( .CIN(\mult_26/ab[25][13] ), .IN0(
        \mult_26/CARRYB[24][13] ), .IN1(\mult_26/SUMB[24][14] ), .COUT(
        \mult_26/CARRYB[25][13] ), .SUM(\mult_26/SUMB[25][13] ) );
  FADDER \mult_26/S2_25_12  ( .CIN(\mult_26/ab[25][12] ), .IN0(
        \mult_26/CARRYB[24][12] ), .IN1(\mult_26/SUMB[24][13] ), .COUT(
        \mult_26/CARRYB[25][12] ), .SUM(\mult_26/SUMB[25][12] ) );
  FADDER \mult_26/S2_25_11  ( .CIN(\mult_26/ab[25][11] ), .IN0(
        \mult_26/CARRYB[24][11] ), .IN1(\mult_26/SUMB[24][12] ), .COUT(
        \mult_26/CARRYB[25][11] ), .SUM(\mult_26/SUMB[25][11] ) );
  FADDER \mult_26/S2_25_10  ( .CIN(\mult_26/ab[25][10] ), .IN0(
        \mult_26/CARRYB[24][10] ), .IN1(\mult_26/SUMB[24][11] ), .COUT(
        \mult_26/CARRYB[25][10] ), .SUM(\mult_26/SUMB[25][10] ) );
  FADDER \mult_26/S2_25_9  ( .CIN(\mult_26/ab[25][9] ), .IN0(
        \mult_26/CARRYB[24][9] ), .IN1(\mult_26/SUMB[24][10] ), .COUT(
        \mult_26/CARRYB[25][9] ), .SUM(\mult_26/SUMB[25][9] ) );
  FADDER \mult_26/S2_25_8  ( .CIN(\mult_26/ab[25][8] ), .IN0(
        \mult_26/CARRYB[24][8] ), .IN1(\mult_26/SUMB[24][9] ), .COUT(
        \mult_26/CARRYB[25][8] ), .SUM(\mult_26/SUMB[25][8] ) );
  FADDER \mult_26/S2_25_7  ( .CIN(\mult_26/ab[25][7] ), .IN0(
        \mult_26/CARRYB[24][7] ), .IN1(\mult_26/SUMB[24][8] ), .COUT(
        \mult_26/CARRYB[25][7] ), .SUM(\mult_26/SUMB[25][7] ) );
  FADDER \mult_26/S2_25_6  ( .CIN(\mult_26/ab[25][6] ), .IN0(
        \mult_26/CARRYB[24][6] ), .IN1(\mult_26/SUMB[24][7] ), .COUT(
        \mult_26/CARRYB[25][6] ), .SUM(\mult_26/SUMB[25][6] ) );
  FADDER \mult_26/S2_25_5  ( .CIN(\mult_26/ab[25][5] ), .IN0(
        \mult_26/CARRYB[24][5] ), .IN1(\mult_26/SUMB[24][6] ), .COUT(
        \mult_26/CARRYB[25][5] ), .SUM(\mult_26/SUMB[25][5] ) );
  FADDER \mult_26/S2_25_4  ( .CIN(\mult_26/ab[25][4] ), .IN0(
        \mult_26/CARRYB[24][4] ), .IN1(\mult_26/SUMB[24][5] ), .COUT(
        \mult_26/CARRYB[25][4] ), .SUM(\mult_26/SUMB[25][4] ) );
  FADDER \mult_26/S2_25_3  ( .CIN(\mult_26/ab[25][3] ), .IN0(
        \mult_26/CARRYB[24][3] ), .IN1(\mult_26/SUMB[24][4] ), .COUT(
        \mult_26/CARRYB[25][3] ), .SUM(\mult_26/SUMB[25][3] ) );
  FADDER \mult_26/S2_25_2  ( .CIN(\mult_26/ab[25][2] ), .IN0(
        \mult_26/CARRYB[24][2] ), .IN1(\mult_26/SUMB[24][3] ), .COUT(
        \mult_26/CARRYB[25][2] ), .SUM(\mult_26/SUMB[25][2] ) );
  FADDER \mult_26/S2_25_1  ( .CIN(\mult_26/ab[25][1] ), .IN0(
        \mult_26/CARRYB[24][1] ), .IN1(\mult_26/SUMB[24][2] ), .COUT(
        \mult_26/CARRYB[25][1] ), .SUM(\mult_26/SUMB[25][1] ) );
  FADDER \mult_26/S1_25_0  ( .CIN(\mult_26/ab[25][0] ), .IN0(
        \mult_26/CARRYB[24][0] ), .IN1(\mult_26/SUMB[24][1] ), .COUT(
        \mult_26/CARRYB[25][0] ), .SUM(o[25]) );
  FADDER \mult_26/S3_26_30  ( .CIN(\mult_26/ab[26][30] ), .IN0(
        \mult_26/CARRYB[25][30] ), .IN1(\mult_26/ab[25][31] ), .COUT(
        \mult_26/CARRYB[26][30] ), .SUM(\mult_26/SUMB[26][30] ) );
  FADDER \mult_26/S2_26_29  ( .CIN(\mult_26/ab[26][29] ), .IN0(
        \mult_26/CARRYB[25][29] ), .IN1(\mult_26/SUMB[25][30] ), .COUT(
        \mult_26/CARRYB[26][29] ), .SUM(\mult_26/SUMB[26][29] ) );
  FADDER \mult_26/S2_26_28  ( .CIN(\mult_26/ab[26][28] ), .IN0(
        \mult_26/CARRYB[25][28] ), .IN1(\mult_26/SUMB[25][29] ), .COUT(
        \mult_26/CARRYB[26][28] ), .SUM(\mult_26/SUMB[26][28] ) );
  FADDER \mult_26/S2_26_27  ( .CIN(\mult_26/ab[26][27] ), .IN0(
        \mult_26/CARRYB[25][27] ), .IN1(\mult_26/SUMB[25][28] ), .COUT(
        \mult_26/CARRYB[26][27] ), .SUM(\mult_26/SUMB[26][27] ) );
  FADDER \mult_26/S2_26_26  ( .CIN(\mult_26/ab[26][26] ), .IN0(
        \mult_26/CARRYB[25][26] ), .IN1(\mult_26/SUMB[25][27] ), .COUT(
        \mult_26/CARRYB[26][26] ), .SUM(\mult_26/SUMB[26][26] ) );
  FADDER \mult_26/S2_26_25  ( .CIN(\mult_26/ab[26][25] ), .IN0(
        \mult_26/CARRYB[25][25] ), .IN1(\mult_26/SUMB[25][26] ), .COUT(
        \mult_26/CARRYB[26][25] ), .SUM(\mult_26/SUMB[26][25] ) );
  FADDER \mult_26/S2_26_24  ( .CIN(\mult_26/ab[26][24] ), .IN0(
        \mult_26/CARRYB[25][24] ), .IN1(\mult_26/SUMB[25][25] ), .COUT(
        \mult_26/CARRYB[26][24] ), .SUM(\mult_26/SUMB[26][24] ) );
  FADDER \mult_26/S2_26_23  ( .CIN(\mult_26/ab[26][23] ), .IN0(
        \mult_26/CARRYB[25][23] ), .IN1(\mult_26/SUMB[25][24] ), .COUT(
        \mult_26/CARRYB[26][23] ), .SUM(\mult_26/SUMB[26][23] ) );
  FADDER \mult_26/S2_26_22  ( .CIN(\mult_26/ab[26][22] ), .IN0(
        \mult_26/CARRYB[25][22] ), .IN1(\mult_26/SUMB[25][23] ), .COUT(
        \mult_26/CARRYB[26][22] ), .SUM(\mult_26/SUMB[26][22] ) );
  FADDER \mult_26/S2_26_21  ( .CIN(\mult_26/ab[26][21] ), .IN0(
        \mult_26/CARRYB[25][21] ), .IN1(\mult_26/SUMB[25][22] ), .COUT(
        \mult_26/CARRYB[26][21] ), .SUM(\mult_26/SUMB[26][21] ) );
  FADDER \mult_26/S2_26_20  ( .CIN(\mult_26/ab[26][20] ), .IN0(
        \mult_26/CARRYB[25][20] ), .IN1(\mult_26/SUMB[25][21] ), .COUT(
        \mult_26/CARRYB[26][20] ), .SUM(\mult_26/SUMB[26][20] ) );
  FADDER \mult_26/S2_26_19  ( .CIN(\mult_26/ab[26][19] ), .IN0(
        \mult_26/CARRYB[25][19] ), .IN1(\mult_26/SUMB[25][20] ), .COUT(
        \mult_26/CARRYB[26][19] ), .SUM(\mult_26/SUMB[26][19] ) );
  FADDER \mult_26/S2_26_18  ( .CIN(\mult_26/ab[26][18] ), .IN0(
        \mult_26/CARRYB[25][18] ), .IN1(\mult_26/SUMB[25][19] ), .COUT(
        \mult_26/CARRYB[26][18] ), .SUM(\mult_26/SUMB[26][18] ) );
  FADDER \mult_26/S2_26_17  ( .CIN(\mult_26/ab[26][17] ), .IN0(
        \mult_26/CARRYB[25][17] ), .IN1(\mult_26/SUMB[25][18] ), .COUT(
        \mult_26/CARRYB[26][17] ), .SUM(\mult_26/SUMB[26][17] ) );
  FADDER \mult_26/S2_26_16  ( .CIN(\mult_26/ab[26][16] ), .IN0(
        \mult_26/CARRYB[25][16] ), .IN1(\mult_26/SUMB[25][17] ), .COUT(
        \mult_26/CARRYB[26][16] ), .SUM(\mult_26/SUMB[26][16] ) );
  FADDER \mult_26/S2_26_15  ( .CIN(\mult_26/ab[26][15] ), .IN0(
        \mult_26/CARRYB[25][15] ), .IN1(\mult_26/SUMB[25][16] ), .COUT(
        \mult_26/CARRYB[26][15] ), .SUM(\mult_26/SUMB[26][15] ) );
  FADDER \mult_26/S2_26_14  ( .CIN(\mult_26/ab[26][14] ), .IN0(
        \mult_26/CARRYB[25][14] ), .IN1(\mult_26/SUMB[25][15] ), .COUT(
        \mult_26/CARRYB[26][14] ), .SUM(\mult_26/SUMB[26][14] ) );
  FADDER \mult_26/S2_26_13  ( .CIN(\mult_26/ab[26][13] ), .IN0(
        \mult_26/CARRYB[25][13] ), .IN1(\mult_26/SUMB[25][14] ), .COUT(
        \mult_26/CARRYB[26][13] ), .SUM(\mult_26/SUMB[26][13] ) );
  FADDER \mult_26/S2_26_12  ( .CIN(\mult_26/ab[26][12] ), .IN0(
        \mult_26/CARRYB[25][12] ), .IN1(\mult_26/SUMB[25][13] ), .COUT(
        \mult_26/CARRYB[26][12] ), .SUM(\mult_26/SUMB[26][12] ) );
  FADDER \mult_26/S2_26_11  ( .CIN(\mult_26/ab[26][11] ), .IN0(
        \mult_26/CARRYB[25][11] ), .IN1(\mult_26/SUMB[25][12] ), .COUT(
        \mult_26/CARRYB[26][11] ), .SUM(\mult_26/SUMB[26][11] ) );
  FADDER \mult_26/S2_26_10  ( .CIN(\mult_26/ab[26][10] ), .IN0(
        \mult_26/CARRYB[25][10] ), .IN1(\mult_26/SUMB[25][11] ), .COUT(
        \mult_26/CARRYB[26][10] ), .SUM(\mult_26/SUMB[26][10] ) );
  FADDER \mult_26/S2_26_9  ( .CIN(\mult_26/ab[26][9] ), .IN0(
        \mult_26/CARRYB[25][9] ), .IN1(\mult_26/SUMB[25][10] ), .COUT(
        \mult_26/CARRYB[26][9] ), .SUM(\mult_26/SUMB[26][9] ) );
  FADDER \mult_26/S2_26_8  ( .CIN(\mult_26/ab[26][8] ), .IN0(
        \mult_26/CARRYB[25][8] ), .IN1(\mult_26/SUMB[25][9] ), .COUT(
        \mult_26/CARRYB[26][8] ), .SUM(\mult_26/SUMB[26][8] ) );
  FADDER \mult_26/S2_26_7  ( .CIN(\mult_26/ab[26][7] ), .IN0(
        \mult_26/CARRYB[25][7] ), .IN1(\mult_26/SUMB[25][8] ), .COUT(
        \mult_26/CARRYB[26][7] ), .SUM(\mult_26/SUMB[26][7] ) );
  FADDER \mult_26/S2_26_6  ( .CIN(\mult_26/ab[26][6] ), .IN0(
        \mult_26/CARRYB[25][6] ), .IN1(\mult_26/SUMB[25][7] ), .COUT(
        \mult_26/CARRYB[26][6] ), .SUM(\mult_26/SUMB[26][6] ) );
  FADDER \mult_26/S2_26_5  ( .CIN(\mult_26/ab[26][5] ), .IN0(
        \mult_26/CARRYB[25][5] ), .IN1(\mult_26/SUMB[25][6] ), .COUT(
        \mult_26/CARRYB[26][5] ), .SUM(\mult_26/SUMB[26][5] ) );
  FADDER \mult_26/S2_26_4  ( .CIN(\mult_26/ab[26][4] ), .IN0(
        \mult_26/CARRYB[25][4] ), .IN1(\mult_26/SUMB[25][5] ), .COUT(
        \mult_26/CARRYB[26][4] ), .SUM(\mult_26/SUMB[26][4] ) );
  FADDER \mult_26/S2_26_3  ( .CIN(\mult_26/ab[26][3] ), .IN0(
        \mult_26/CARRYB[25][3] ), .IN1(\mult_26/SUMB[25][4] ), .COUT(
        \mult_26/CARRYB[26][3] ), .SUM(\mult_26/SUMB[26][3] ) );
  FADDER \mult_26/S2_26_2  ( .CIN(\mult_26/ab[26][2] ), .IN0(
        \mult_26/CARRYB[25][2] ), .IN1(\mult_26/SUMB[25][3] ), .COUT(
        \mult_26/CARRYB[26][2] ), .SUM(\mult_26/SUMB[26][2] ) );
  FADDER \mult_26/S2_26_1  ( .CIN(\mult_26/ab[26][1] ), .IN0(
        \mult_26/CARRYB[25][1] ), .IN1(\mult_26/SUMB[25][2] ), .COUT(
        \mult_26/CARRYB[26][1] ), .SUM(\mult_26/SUMB[26][1] ) );
  FADDER \mult_26/S1_26_0  ( .CIN(\mult_26/ab[26][0] ), .IN0(
        \mult_26/CARRYB[25][0] ), .IN1(\mult_26/SUMB[25][1] ), .COUT(
        \mult_26/CARRYB[26][0] ), .SUM(o[26]) );
  FADDER \mult_26/S3_27_30  ( .CIN(\mult_26/ab[27][30] ), .IN0(
        \mult_26/CARRYB[26][30] ), .IN1(\mult_26/ab[26][31] ), .COUT(
        \mult_26/CARRYB[27][30] ), .SUM(\mult_26/SUMB[27][30] ) );
  FADDER \mult_26/S2_27_29  ( .CIN(\mult_26/ab[27][29] ), .IN0(
        \mult_26/CARRYB[26][29] ), .IN1(\mult_26/SUMB[26][30] ), .COUT(
        \mult_26/CARRYB[27][29] ), .SUM(\mult_26/SUMB[27][29] ) );
  FADDER \mult_26/S2_27_28  ( .CIN(\mult_26/ab[27][28] ), .IN0(
        \mult_26/CARRYB[26][28] ), .IN1(\mult_26/SUMB[26][29] ), .COUT(
        \mult_26/CARRYB[27][28] ), .SUM(\mult_26/SUMB[27][28] ) );
  FADDER \mult_26/S2_27_27  ( .CIN(\mult_26/ab[27][27] ), .IN0(
        \mult_26/CARRYB[26][27] ), .IN1(\mult_26/SUMB[26][28] ), .COUT(
        \mult_26/CARRYB[27][27] ), .SUM(\mult_26/SUMB[27][27] ) );
  FADDER \mult_26/S2_27_26  ( .CIN(\mult_26/ab[27][26] ), .IN0(
        \mult_26/CARRYB[26][26] ), .IN1(\mult_26/SUMB[26][27] ), .COUT(
        \mult_26/CARRYB[27][26] ), .SUM(\mult_26/SUMB[27][26] ) );
  FADDER \mult_26/S2_27_25  ( .CIN(\mult_26/ab[27][25] ), .IN0(
        \mult_26/CARRYB[26][25] ), .IN1(\mult_26/SUMB[26][26] ), .COUT(
        \mult_26/CARRYB[27][25] ), .SUM(\mult_26/SUMB[27][25] ) );
  FADDER \mult_26/S2_27_24  ( .CIN(\mult_26/ab[27][24] ), .IN0(
        \mult_26/CARRYB[26][24] ), .IN1(\mult_26/SUMB[26][25] ), .COUT(
        \mult_26/CARRYB[27][24] ), .SUM(\mult_26/SUMB[27][24] ) );
  FADDER \mult_26/S2_27_23  ( .CIN(\mult_26/ab[27][23] ), .IN0(
        \mult_26/CARRYB[26][23] ), .IN1(\mult_26/SUMB[26][24] ), .COUT(
        \mult_26/CARRYB[27][23] ), .SUM(\mult_26/SUMB[27][23] ) );
  FADDER \mult_26/S2_27_22  ( .CIN(\mult_26/ab[27][22] ), .IN0(
        \mult_26/CARRYB[26][22] ), .IN1(\mult_26/SUMB[26][23] ), .COUT(
        \mult_26/CARRYB[27][22] ), .SUM(\mult_26/SUMB[27][22] ) );
  FADDER \mult_26/S2_27_21  ( .CIN(\mult_26/ab[27][21] ), .IN0(
        \mult_26/CARRYB[26][21] ), .IN1(\mult_26/SUMB[26][22] ), .COUT(
        \mult_26/CARRYB[27][21] ), .SUM(\mult_26/SUMB[27][21] ) );
  FADDER \mult_26/S2_27_20  ( .CIN(\mult_26/ab[27][20] ), .IN0(
        \mult_26/CARRYB[26][20] ), .IN1(\mult_26/SUMB[26][21] ), .COUT(
        \mult_26/CARRYB[27][20] ), .SUM(\mult_26/SUMB[27][20] ) );
  FADDER \mult_26/S2_27_19  ( .CIN(\mult_26/ab[27][19] ), .IN0(
        \mult_26/CARRYB[26][19] ), .IN1(\mult_26/SUMB[26][20] ), .COUT(
        \mult_26/CARRYB[27][19] ), .SUM(\mult_26/SUMB[27][19] ) );
  FADDER \mult_26/S2_27_18  ( .CIN(\mult_26/ab[27][18] ), .IN0(
        \mult_26/CARRYB[26][18] ), .IN1(\mult_26/SUMB[26][19] ), .COUT(
        \mult_26/CARRYB[27][18] ), .SUM(\mult_26/SUMB[27][18] ) );
  FADDER \mult_26/S2_27_17  ( .CIN(\mult_26/ab[27][17] ), .IN0(
        \mult_26/CARRYB[26][17] ), .IN1(\mult_26/SUMB[26][18] ), .COUT(
        \mult_26/CARRYB[27][17] ), .SUM(\mult_26/SUMB[27][17] ) );
  FADDER \mult_26/S2_27_16  ( .CIN(\mult_26/ab[27][16] ), .IN0(
        \mult_26/CARRYB[26][16] ), .IN1(\mult_26/SUMB[26][17] ), .COUT(
        \mult_26/CARRYB[27][16] ), .SUM(\mult_26/SUMB[27][16] ) );
  FADDER \mult_26/S2_27_15  ( .CIN(\mult_26/ab[27][15] ), .IN0(
        \mult_26/CARRYB[26][15] ), .IN1(\mult_26/SUMB[26][16] ), .COUT(
        \mult_26/CARRYB[27][15] ), .SUM(\mult_26/SUMB[27][15] ) );
  FADDER \mult_26/S2_27_14  ( .CIN(\mult_26/ab[27][14] ), .IN0(
        \mult_26/CARRYB[26][14] ), .IN1(\mult_26/SUMB[26][15] ), .COUT(
        \mult_26/CARRYB[27][14] ), .SUM(\mult_26/SUMB[27][14] ) );
  FADDER \mult_26/S2_27_13  ( .CIN(\mult_26/ab[27][13] ), .IN0(
        \mult_26/CARRYB[26][13] ), .IN1(\mult_26/SUMB[26][14] ), .COUT(
        \mult_26/CARRYB[27][13] ), .SUM(\mult_26/SUMB[27][13] ) );
  FADDER \mult_26/S2_27_12  ( .CIN(\mult_26/ab[27][12] ), .IN0(
        \mult_26/CARRYB[26][12] ), .IN1(\mult_26/SUMB[26][13] ), .COUT(
        \mult_26/CARRYB[27][12] ), .SUM(\mult_26/SUMB[27][12] ) );
  FADDER \mult_26/S2_27_11  ( .CIN(\mult_26/ab[27][11] ), .IN0(
        \mult_26/CARRYB[26][11] ), .IN1(\mult_26/SUMB[26][12] ), .COUT(
        \mult_26/CARRYB[27][11] ), .SUM(\mult_26/SUMB[27][11] ) );
  FADDER \mult_26/S2_27_10  ( .CIN(\mult_26/ab[27][10] ), .IN0(
        \mult_26/CARRYB[26][10] ), .IN1(\mult_26/SUMB[26][11] ), .COUT(
        \mult_26/CARRYB[27][10] ), .SUM(\mult_26/SUMB[27][10] ) );
  FADDER \mult_26/S2_27_9  ( .CIN(\mult_26/ab[27][9] ), .IN0(
        \mult_26/CARRYB[26][9] ), .IN1(\mult_26/SUMB[26][10] ), .COUT(
        \mult_26/CARRYB[27][9] ), .SUM(\mult_26/SUMB[27][9] ) );
  FADDER \mult_26/S2_27_8  ( .CIN(\mult_26/ab[27][8] ), .IN0(
        \mult_26/CARRYB[26][8] ), .IN1(\mult_26/SUMB[26][9] ), .COUT(
        \mult_26/CARRYB[27][8] ), .SUM(\mult_26/SUMB[27][8] ) );
  FADDER \mult_26/S2_27_7  ( .CIN(\mult_26/ab[27][7] ), .IN0(
        \mult_26/CARRYB[26][7] ), .IN1(\mult_26/SUMB[26][8] ), .COUT(
        \mult_26/CARRYB[27][7] ), .SUM(\mult_26/SUMB[27][7] ) );
  FADDER \mult_26/S2_27_6  ( .CIN(\mult_26/ab[27][6] ), .IN0(
        \mult_26/CARRYB[26][6] ), .IN1(\mult_26/SUMB[26][7] ), .COUT(
        \mult_26/CARRYB[27][6] ), .SUM(\mult_26/SUMB[27][6] ) );
  FADDER \mult_26/S2_27_5  ( .CIN(\mult_26/ab[27][5] ), .IN0(
        \mult_26/CARRYB[26][5] ), .IN1(\mult_26/SUMB[26][6] ), .COUT(
        \mult_26/CARRYB[27][5] ), .SUM(\mult_26/SUMB[27][5] ) );
  FADDER \mult_26/S2_27_4  ( .CIN(\mult_26/ab[27][4] ), .IN0(
        \mult_26/CARRYB[26][4] ), .IN1(\mult_26/SUMB[26][5] ), .COUT(
        \mult_26/CARRYB[27][4] ), .SUM(\mult_26/SUMB[27][4] ) );
  FADDER \mult_26/S2_27_3  ( .CIN(\mult_26/ab[27][3] ), .IN0(
        \mult_26/CARRYB[26][3] ), .IN1(\mult_26/SUMB[26][4] ), .COUT(
        \mult_26/CARRYB[27][3] ), .SUM(\mult_26/SUMB[27][3] ) );
  FADDER \mult_26/S2_27_2  ( .CIN(\mult_26/ab[27][2] ), .IN0(
        \mult_26/CARRYB[26][2] ), .IN1(\mult_26/SUMB[26][3] ), .COUT(
        \mult_26/CARRYB[27][2] ), .SUM(\mult_26/SUMB[27][2] ) );
  FADDER \mult_26/S2_27_1  ( .CIN(\mult_26/ab[27][1] ), .IN0(
        \mult_26/CARRYB[26][1] ), .IN1(\mult_26/SUMB[26][2] ), .COUT(
        \mult_26/CARRYB[27][1] ), .SUM(\mult_26/SUMB[27][1] ) );
  FADDER \mult_26/S1_27_0  ( .CIN(\mult_26/ab[27][0] ), .IN0(
        \mult_26/CARRYB[26][0] ), .IN1(\mult_26/SUMB[26][1] ), .COUT(
        \mult_26/CARRYB[27][0] ), .SUM(o[27]) );
  FADDER \mult_26/S3_28_30  ( .CIN(\mult_26/ab[28][30] ), .IN0(
        \mult_26/CARRYB[27][30] ), .IN1(\mult_26/ab[27][31] ), .COUT(
        \mult_26/CARRYB[28][30] ), .SUM(\mult_26/SUMB[28][30] ) );
  FADDER \mult_26/S2_28_29  ( .CIN(\mult_26/ab[28][29] ), .IN0(
        \mult_26/CARRYB[27][29] ), .IN1(\mult_26/SUMB[27][30] ), .COUT(
        \mult_26/CARRYB[28][29] ), .SUM(\mult_26/SUMB[28][29] ) );
  FADDER \mult_26/S2_28_28  ( .CIN(\mult_26/ab[28][28] ), .IN0(
        \mult_26/CARRYB[27][28] ), .IN1(\mult_26/SUMB[27][29] ), .COUT(
        \mult_26/CARRYB[28][28] ), .SUM(\mult_26/SUMB[28][28] ) );
  FADDER \mult_26/S2_28_27  ( .CIN(\mult_26/ab[28][27] ), .IN0(
        \mult_26/CARRYB[27][27] ), .IN1(\mult_26/SUMB[27][28] ), .COUT(
        \mult_26/CARRYB[28][27] ), .SUM(\mult_26/SUMB[28][27] ) );
  FADDER \mult_26/S2_28_26  ( .CIN(\mult_26/ab[28][26] ), .IN0(
        \mult_26/CARRYB[27][26] ), .IN1(\mult_26/SUMB[27][27] ), .COUT(
        \mult_26/CARRYB[28][26] ), .SUM(\mult_26/SUMB[28][26] ) );
  FADDER \mult_26/S2_28_25  ( .CIN(\mult_26/ab[28][25] ), .IN0(
        \mult_26/CARRYB[27][25] ), .IN1(\mult_26/SUMB[27][26] ), .COUT(
        \mult_26/CARRYB[28][25] ), .SUM(\mult_26/SUMB[28][25] ) );
  FADDER \mult_26/S2_28_24  ( .CIN(\mult_26/ab[28][24] ), .IN0(
        \mult_26/CARRYB[27][24] ), .IN1(\mult_26/SUMB[27][25] ), .COUT(
        \mult_26/CARRYB[28][24] ), .SUM(\mult_26/SUMB[28][24] ) );
  FADDER \mult_26/S2_28_23  ( .CIN(\mult_26/ab[28][23] ), .IN0(
        \mult_26/CARRYB[27][23] ), .IN1(\mult_26/SUMB[27][24] ), .COUT(
        \mult_26/CARRYB[28][23] ), .SUM(\mult_26/SUMB[28][23] ) );
  FADDER \mult_26/S2_28_22  ( .CIN(\mult_26/ab[28][22] ), .IN0(
        \mult_26/CARRYB[27][22] ), .IN1(\mult_26/SUMB[27][23] ), .COUT(
        \mult_26/CARRYB[28][22] ), .SUM(\mult_26/SUMB[28][22] ) );
  FADDER \mult_26/S2_28_21  ( .CIN(\mult_26/ab[28][21] ), .IN0(
        \mult_26/CARRYB[27][21] ), .IN1(\mult_26/SUMB[27][22] ), .COUT(
        \mult_26/CARRYB[28][21] ), .SUM(\mult_26/SUMB[28][21] ) );
  FADDER \mult_26/S2_28_20  ( .CIN(\mult_26/ab[28][20] ), .IN0(
        \mult_26/CARRYB[27][20] ), .IN1(\mult_26/SUMB[27][21] ), .COUT(
        \mult_26/CARRYB[28][20] ), .SUM(\mult_26/SUMB[28][20] ) );
  FADDER \mult_26/S2_28_19  ( .CIN(\mult_26/ab[28][19] ), .IN0(
        \mult_26/CARRYB[27][19] ), .IN1(\mult_26/SUMB[27][20] ), .COUT(
        \mult_26/CARRYB[28][19] ), .SUM(\mult_26/SUMB[28][19] ) );
  FADDER \mult_26/S2_28_18  ( .CIN(\mult_26/ab[28][18] ), .IN0(
        \mult_26/CARRYB[27][18] ), .IN1(\mult_26/SUMB[27][19] ), .COUT(
        \mult_26/CARRYB[28][18] ), .SUM(\mult_26/SUMB[28][18] ) );
  FADDER \mult_26/S2_28_17  ( .CIN(\mult_26/ab[28][17] ), .IN0(
        \mult_26/CARRYB[27][17] ), .IN1(\mult_26/SUMB[27][18] ), .COUT(
        \mult_26/CARRYB[28][17] ), .SUM(\mult_26/SUMB[28][17] ) );
  FADDER \mult_26/S2_28_16  ( .CIN(\mult_26/ab[28][16] ), .IN0(
        \mult_26/CARRYB[27][16] ), .IN1(\mult_26/SUMB[27][17] ), .COUT(
        \mult_26/CARRYB[28][16] ), .SUM(\mult_26/SUMB[28][16] ) );
  FADDER \mult_26/S2_28_15  ( .CIN(\mult_26/ab[28][15] ), .IN0(
        \mult_26/CARRYB[27][15] ), .IN1(\mult_26/SUMB[27][16] ), .COUT(
        \mult_26/CARRYB[28][15] ), .SUM(\mult_26/SUMB[28][15] ) );
  FADDER \mult_26/S2_28_14  ( .CIN(\mult_26/ab[28][14] ), .IN0(
        \mult_26/CARRYB[27][14] ), .IN1(\mult_26/SUMB[27][15] ), .COUT(
        \mult_26/CARRYB[28][14] ), .SUM(\mult_26/SUMB[28][14] ) );
  FADDER \mult_26/S2_28_13  ( .CIN(\mult_26/ab[28][13] ), .IN0(
        \mult_26/CARRYB[27][13] ), .IN1(\mult_26/SUMB[27][14] ), .COUT(
        \mult_26/CARRYB[28][13] ), .SUM(\mult_26/SUMB[28][13] ) );
  FADDER \mult_26/S2_28_12  ( .CIN(\mult_26/ab[28][12] ), .IN0(
        \mult_26/CARRYB[27][12] ), .IN1(\mult_26/SUMB[27][13] ), .COUT(
        \mult_26/CARRYB[28][12] ), .SUM(\mult_26/SUMB[28][12] ) );
  FADDER \mult_26/S2_28_11  ( .CIN(\mult_26/ab[28][11] ), .IN0(
        \mult_26/CARRYB[27][11] ), .IN1(\mult_26/SUMB[27][12] ), .COUT(
        \mult_26/CARRYB[28][11] ), .SUM(\mult_26/SUMB[28][11] ) );
  FADDER \mult_26/S2_28_10  ( .CIN(\mult_26/ab[28][10] ), .IN0(
        \mult_26/CARRYB[27][10] ), .IN1(\mult_26/SUMB[27][11] ), .COUT(
        \mult_26/CARRYB[28][10] ), .SUM(\mult_26/SUMB[28][10] ) );
  FADDER \mult_26/S2_28_9  ( .CIN(\mult_26/ab[28][9] ), .IN0(
        \mult_26/CARRYB[27][9] ), .IN1(\mult_26/SUMB[27][10] ), .COUT(
        \mult_26/CARRYB[28][9] ), .SUM(\mult_26/SUMB[28][9] ) );
  FADDER \mult_26/S2_28_8  ( .CIN(\mult_26/ab[28][8] ), .IN0(
        \mult_26/CARRYB[27][8] ), .IN1(\mult_26/SUMB[27][9] ), .COUT(
        \mult_26/CARRYB[28][8] ), .SUM(\mult_26/SUMB[28][8] ) );
  FADDER \mult_26/S2_28_7  ( .CIN(\mult_26/ab[28][7] ), .IN0(
        \mult_26/CARRYB[27][7] ), .IN1(\mult_26/SUMB[27][8] ), .COUT(
        \mult_26/CARRYB[28][7] ), .SUM(\mult_26/SUMB[28][7] ) );
  FADDER \mult_26/S2_28_6  ( .CIN(\mult_26/ab[28][6] ), .IN0(
        \mult_26/CARRYB[27][6] ), .IN1(\mult_26/SUMB[27][7] ), .COUT(
        \mult_26/CARRYB[28][6] ), .SUM(\mult_26/SUMB[28][6] ) );
  FADDER \mult_26/S2_28_5  ( .CIN(\mult_26/ab[28][5] ), .IN0(
        \mult_26/CARRYB[27][5] ), .IN1(\mult_26/SUMB[27][6] ), .COUT(
        \mult_26/CARRYB[28][5] ), .SUM(\mult_26/SUMB[28][5] ) );
  FADDER \mult_26/S2_28_4  ( .CIN(\mult_26/ab[28][4] ), .IN0(
        \mult_26/CARRYB[27][4] ), .IN1(\mult_26/SUMB[27][5] ), .COUT(
        \mult_26/CARRYB[28][4] ), .SUM(\mult_26/SUMB[28][4] ) );
  FADDER \mult_26/S2_28_3  ( .CIN(\mult_26/ab[28][3] ), .IN0(
        \mult_26/CARRYB[27][3] ), .IN1(\mult_26/SUMB[27][4] ), .COUT(
        \mult_26/CARRYB[28][3] ), .SUM(\mult_26/SUMB[28][3] ) );
  FADDER \mult_26/S2_28_2  ( .CIN(\mult_26/ab[28][2] ), .IN0(
        \mult_26/CARRYB[27][2] ), .IN1(\mult_26/SUMB[27][3] ), .COUT(
        \mult_26/CARRYB[28][2] ), .SUM(\mult_26/SUMB[28][2] ) );
  FADDER \mult_26/S2_28_1  ( .CIN(\mult_26/ab[28][1] ), .IN0(
        \mult_26/CARRYB[27][1] ), .IN1(\mult_26/SUMB[27][2] ), .COUT(
        \mult_26/CARRYB[28][1] ), .SUM(\mult_26/SUMB[28][1] ) );
  FADDER \mult_26/S1_28_0  ( .CIN(\mult_26/ab[28][0] ), .IN0(
        \mult_26/CARRYB[27][0] ), .IN1(\mult_26/SUMB[27][1] ), .COUT(
        \mult_26/CARRYB[28][0] ), .SUM(o[28]) );
  FADDER \mult_26/S3_29_30  ( .CIN(\mult_26/ab[29][30] ), .IN0(
        \mult_26/CARRYB[28][30] ), .IN1(\mult_26/ab[28][31] ), .COUT(
        \mult_26/CARRYB[29][30] ), .SUM(\mult_26/SUMB[29][30] ) );
  FADDER \mult_26/S2_29_29  ( .CIN(\mult_26/ab[29][29] ), .IN0(
        \mult_26/CARRYB[28][29] ), .IN1(\mult_26/SUMB[28][30] ), .COUT(
        \mult_26/CARRYB[29][29] ), .SUM(\mult_26/SUMB[29][29] ) );
  FADDER \mult_26/S2_29_28  ( .CIN(\mult_26/ab[29][28] ), .IN0(
        \mult_26/CARRYB[28][28] ), .IN1(\mult_26/SUMB[28][29] ), .COUT(
        \mult_26/CARRYB[29][28] ), .SUM(\mult_26/SUMB[29][28] ) );
  FADDER \mult_26/S2_29_27  ( .CIN(\mult_26/ab[29][27] ), .IN0(
        \mult_26/CARRYB[28][27] ), .IN1(\mult_26/SUMB[28][28] ), .COUT(
        \mult_26/CARRYB[29][27] ), .SUM(\mult_26/SUMB[29][27] ) );
  FADDER \mult_26/S2_29_26  ( .CIN(\mult_26/ab[29][26] ), .IN0(
        \mult_26/CARRYB[28][26] ), .IN1(\mult_26/SUMB[28][27] ), .COUT(
        \mult_26/CARRYB[29][26] ), .SUM(\mult_26/SUMB[29][26] ) );
  FADDER \mult_26/S2_29_25  ( .CIN(\mult_26/ab[29][25] ), .IN0(
        \mult_26/CARRYB[28][25] ), .IN1(\mult_26/SUMB[28][26] ), .COUT(
        \mult_26/CARRYB[29][25] ), .SUM(\mult_26/SUMB[29][25] ) );
  FADDER \mult_26/S2_29_24  ( .CIN(\mult_26/ab[29][24] ), .IN0(
        \mult_26/CARRYB[28][24] ), .IN1(\mult_26/SUMB[28][25] ), .COUT(
        \mult_26/CARRYB[29][24] ), .SUM(\mult_26/SUMB[29][24] ) );
  FADDER \mult_26/S2_29_23  ( .CIN(\mult_26/ab[29][23] ), .IN0(
        \mult_26/CARRYB[28][23] ), .IN1(\mult_26/SUMB[28][24] ), .COUT(
        \mult_26/CARRYB[29][23] ), .SUM(\mult_26/SUMB[29][23] ) );
  FADDER \mult_26/S2_29_22  ( .CIN(\mult_26/ab[29][22] ), .IN0(
        \mult_26/CARRYB[28][22] ), .IN1(\mult_26/SUMB[28][23] ), .COUT(
        \mult_26/CARRYB[29][22] ), .SUM(\mult_26/SUMB[29][22] ) );
  FADDER \mult_26/S2_29_21  ( .CIN(\mult_26/ab[29][21] ), .IN0(
        \mult_26/CARRYB[28][21] ), .IN1(\mult_26/SUMB[28][22] ), .COUT(
        \mult_26/CARRYB[29][21] ), .SUM(\mult_26/SUMB[29][21] ) );
  FADDER \mult_26/S2_29_20  ( .CIN(\mult_26/ab[29][20] ), .IN0(
        \mult_26/CARRYB[28][20] ), .IN1(\mult_26/SUMB[28][21] ), .COUT(
        \mult_26/CARRYB[29][20] ), .SUM(\mult_26/SUMB[29][20] ) );
  FADDER \mult_26/S2_29_19  ( .CIN(\mult_26/ab[29][19] ), .IN0(
        \mult_26/CARRYB[28][19] ), .IN1(\mult_26/SUMB[28][20] ), .COUT(
        \mult_26/CARRYB[29][19] ), .SUM(\mult_26/SUMB[29][19] ) );
  FADDER \mult_26/S2_29_18  ( .CIN(\mult_26/ab[29][18] ), .IN0(
        \mult_26/CARRYB[28][18] ), .IN1(\mult_26/SUMB[28][19] ), .COUT(
        \mult_26/CARRYB[29][18] ), .SUM(\mult_26/SUMB[29][18] ) );
  FADDER \mult_26/S2_29_17  ( .CIN(\mult_26/ab[29][17] ), .IN0(
        \mult_26/CARRYB[28][17] ), .IN1(\mult_26/SUMB[28][18] ), .COUT(
        \mult_26/CARRYB[29][17] ), .SUM(\mult_26/SUMB[29][17] ) );
  FADDER \mult_26/S2_29_16  ( .CIN(\mult_26/ab[29][16] ), .IN0(
        \mult_26/CARRYB[28][16] ), .IN1(\mult_26/SUMB[28][17] ), .COUT(
        \mult_26/CARRYB[29][16] ), .SUM(\mult_26/SUMB[29][16] ) );
  FADDER \mult_26/S2_29_15  ( .CIN(\mult_26/ab[29][15] ), .IN0(
        \mult_26/CARRYB[28][15] ), .IN1(\mult_26/SUMB[28][16] ), .COUT(
        \mult_26/CARRYB[29][15] ), .SUM(\mult_26/SUMB[29][15] ) );
  FADDER \mult_26/S2_29_14  ( .CIN(\mult_26/ab[29][14] ), .IN0(
        \mult_26/CARRYB[28][14] ), .IN1(\mult_26/SUMB[28][15] ), .COUT(
        \mult_26/CARRYB[29][14] ), .SUM(\mult_26/SUMB[29][14] ) );
  FADDER \mult_26/S2_29_13  ( .CIN(\mult_26/ab[29][13] ), .IN0(
        \mult_26/CARRYB[28][13] ), .IN1(\mult_26/SUMB[28][14] ), .COUT(
        \mult_26/CARRYB[29][13] ), .SUM(\mult_26/SUMB[29][13] ) );
  FADDER \mult_26/S2_29_12  ( .CIN(\mult_26/ab[29][12] ), .IN0(
        \mult_26/CARRYB[28][12] ), .IN1(\mult_26/SUMB[28][13] ), .COUT(
        \mult_26/CARRYB[29][12] ), .SUM(\mult_26/SUMB[29][12] ) );
  FADDER \mult_26/S2_29_11  ( .CIN(\mult_26/ab[29][11] ), .IN0(
        \mult_26/CARRYB[28][11] ), .IN1(\mult_26/SUMB[28][12] ), .COUT(
        \mult_26/CARRYB[29][11] ), .SUM(\mult_26/SUMB[29][11] ) );
  FADDER \mult_26/S2_29_10  ( .CIN(\mult_26/ab[29][10] ), .IN0(
        \mult_26/CARRYB[28][10] ), .IN1(\mult_26/SUMB[28][11] ), .COUT(
        \mult_26/CARRYB[29][10] ), .SUM(\mult_26/SUMB[29][10] ) );
  FADDER \mult_26/S2_29_9  ( .CIN(\mult_26/ab[29][9] ), .IN0(
        \mult_26/CARRYB[28][9] ), .IN1(\mult_26/SUMB[28][10] ), .COUT(
        \mult_26/CARRYB[29][9] ), .SUM(\mult_26/SUMB[29][9] ) );
  FADDER \mult_26/S2_29_8  ( .CIN(\mult_26/ab[29][8] ), .IN0(
        \mult_26/CARRYB[28][8] ), .IN1(\mult_26/SUMB[28][9] ), .COUT(
        \mult_26/CARRYB[29][8] ), .SUM(\mult_26/SUMB[29][8] ) );
  FADDER \mult_26/S2_29_7  ( .CIN(\mult_26/ab[29][7] ), .IN0(
        \mult_26/CARRYB[28][7] ), .IN1(\mult_26/SUMB[28][8] ), .COUT(
        \mult_26/CARRYB[29][7] ), .SUM(\mult_26/SUMB[29][7] ) );
  FADDER \mult_26/S2_29_6  ( .CIN(\mult_26/ab[29][6] ), .IN0(
        \mult_26/CARRYB[28][6] ), .IN1(\mult_26/SUMB[28][7] ), .COUT(
        \mult_26/CARRYB[29][6] ), .SUM(\mult_26/SUMB[29][6] ) );
  FADDER \mult_26/S2_29_5  ( .CIN(\mult_26/ab[29][5] ), .IN0(
        \mult_26/CARRYB[28][5] ), .IN1(\mult_26/SUMB[28][6] ), .COUT(
        \mult_26/CARRYB[29][5] ), .SUM(\mult_26/SUMB[29][5] ) );
  FADDER \mult_26/S2_29_4  ( .CIN(\mult_26/ab[29][4] ), .IN0(
        \mult_26/CARRYB[28][4] ), .IN1(\mult_26/SUMB[28][5] ), .COUT(
        \mult_26/CARRYB[29][4] ), .SUM(\mult_26/SUMB[29][4] ) );
  FADDER \mult_26/S2_29_3  ( .CIN(\mult_26/ab[29][3] ), .IN0(
        \mult_26/CARRYB[28][3] ), .IN1(\mult_26/SUMB[28][4] ), .COUT(
        \mult_26/CARRYB[29][3] ), .SUM(\mult_26/SUMB[29][3] ) );
  FADDER \mult_26/S2_29_2  ( .CIN(\mult_26/ab[29][2] ), .IN0(
        \mult_26/CARRYB[28][2] ), .IN1(\mult_26/SUMB[28][3] ), .COUT(
        \mult_26/CARRYB[29][2] ), .SUM(\mult_26/SUMB[29][2] ) );
  FADDER \mult_26/S2_29_1  ( .CIN(\mult_26/ab[29][1] ), .IN0(
        \mult_26/CARRYB[28][1] ), .IN1(\mult_26/SUMB[28][2] ), .COUT(
        \mult_26/CARRYB[29][1] ), .SUM(\mult_26/SUMB[29][1] ) );
  FADDER \mult_26/S1_29_0  ( .CIN(\mult_26/ab[29][0] ), .IN0(
        \mult_26/CARRYB[28][0] ), .IN1(\mult_26/SUMB[28][1] ), .COUT(
        \mult_26/CARRYB[29][0] ), .SUM(o[29]) );
  FADDER \mult_26/S3_30_30  ( .CIN(\mult_26/ab[30][30] ), .IN0(
        \mult_26/CARRYB[29][30] ), .IN1(\mult_26/ab[29][31] ), .COUT(
        \mult_26/CARRYB[30][30] ), .SUM(\mult_26/SUMB[30][30] ) );
  FADDER \mult_26/S2_30_29  ( .CIN(\mult_26/ab[30][29] ), .IN0(
        \mult_26/CARRYB[29][29] ), .IN1(\mult_26/SUMB[29][30] ), .COUT(
        \mult_26/CARRYB[30][29] ), .SUM(\mult_26/SUMB[30][29] ) );
  FADDER \mult_26/S2_30_28  ( .CIN(\mult_26/ab[30][28] ), .IN0(
        \mult_26/CARRYB[29][28] ), .IN1(\mult_26/SUMB[29][29] ), .COUT(
        \mult_26/CARRYB[30][28] ), .SUM(\mult_26/SUMB[30][28] ) );
  FADDER \mult_26/S2_30_27  ( .CIN(\mult_26/ab[30][27] ), .IN0(
        \mult_26/CARRYB[29][27] ), .IN1(\mult_26/SUMB[29][28] ), .COUT(
        \mult_26/CARRYB[30][27] ), .SUM(\mult_26/SUMB[30][27] ) );
  FADDER \mult_26/S2_30_26  ( .CIN(\mult_26/ab[30][26] ), .IN0(
        \mult_26/CARRYB[29][26] ), .IN1(\mult_26/SUMB[29][27] ), .COUT(
        \mult_26/CARRYB[30][26] ), .SUM(\mult_26/SUMB[30][26] ) );
  FADDER \mult_26/S2_30_25  ( .CIN(\mult_26/ab[30][25] ), .IN0(
        \mult_26/CARRYB[29][25] ), .IN1(\mult_26/SUMB[29][26] ), .COUT(
        \mult_26/CARRYB[30][25] ), .SUM(\mult_26/SUMB[30][25] ) );
  FADDER \mult_26/S2_30_24  ( .CIN(\mult_26/ab[30][24] ), .IN0(
        \mult_26/CARRYB[29][24] ), .IN1(\mult_26/SUMB[29][25] ), .COUT(
        \mult_26/CARRYB[30][24] ), .SUM(\mult_26/SUMB[30][24] ) );
  FADDER \mult_26/S2_30_23  ( .CIN(\mult_26/ab[30][23] ), .IN0(
        \mult_26/CARRYB[29][23] ), .IN1(\mult_26/SUMB[29][24] ), .COUT(
        \mult_26/CARRYB[30][23] ), .SUM(\mult_26/SUMB[30][23] ) );
  FADDER \mult_26/S2_30_22  ( .CIN(\mult_26/ab[30][22] ), .IN0(
        \mult_26/CARRYB[29][22] ), .IN1(\mult_26/SUMB[29][23] ), .COUT(
        \mult_26/CARRYB[30][22] ), .SUM(\mult_26/SUMB[30][22] ) );
  FADDER \mult_26/S2_30_21  ( .CIN(\mult_26/ab[30][21] ), .IN0(
        \mult_26/CARRYB[29][21] ), .IN1(\mult_26/SUMB[29][22] ), .COUT(
        \mult_26/CARRYB[30][21] ), .SUM(\mult_26/SUMB[30][21] ) );
  FADDER \mult_26/S2_30_20  ( .CIN(\mult_26/ab[30][20] ), .IN0(
        \mult_26/CARRYB[29][20] ), .IN1(\mult_26/SUMB[29][21] ), .COUT(
        \mult_26/CARRYB[30][20] ), .SUM(\mult_26/SUMB[30][20] ) );
  FADDER \mult_26/S2_30_19  ( .CIN(\mult_26/ab[30][19] ), .IN0(
        \mult_26/CARRYB[29][19] ), .IN1(\mult_26/SUMB[29][20] ), .COUT(
        \mult_26/CARRYB[30][19] ), .SUM(\mult_26/SUMB[30][19] ) );
  FADDER \mult_26/S2_30_18  ( .CIN(\mult_26/ab[30][18] ), .IN0(
        \mult_26/CARRYB[29][18] ), .IN1(\mult_26/SUMB[29][19] ), .COUT(
        \mult_26/CARRYB[30][18] ), .SUM(\mult_26/SUMB[30][18] ) );
  FADDER \mult_26/S2_30_17  ( .CIN(\mult_26/ab[30][17] ), .IN0(
        \mult_26/CARRYB[29][17] ), .IN1(\mult_26/SUMB[29][18] ), .COUT(
        \mult_26/CARRYB[30][17] ), .SUM(\mult_26/SUMB[30][17] ) );
  FADDER \mult_26/S2_30_16  ( .CIN(\mult_26/ab[30][16] ), .IN0(
        \mult_26/CARRYB[29][16] ), .IN1(\mult_26/SUMB[29][17] ), .COUT(
        \mult_26/CARRYB[30][16] ), .SUM(\mult_26/SUMB[30][16] ) );
  FADDER \mult_26/S2_30_15  ( .CIN(\mult_26/ab[30][15] ), .IN0(
        \mult_26/CARRYB[29][15] ), .IN1(\mult_26/SUMB[29][16] ), .COUT(
        \mult_26/CARRYB[30][15] ), .SUM(\mult_26/SUMB[30][15] ) );
  FADDER \mult_26/S2_30_14  ( .CIN(\mult_26/ab[30][14] ), .IN0(
        \mult_26/CARRYB[29][14] ), .IN1(\mult_26/SUMB[29][15] ), .COUT(
        \mult_26/CARRYB[30][14] ), .SUM(\mult_26/SUMB[30][14] ) );
  FADDER \mult_26/S2_30_13  ( .CIN(\mult_26/ab[30][13] ), .IN0(
        \mult_26/CARRYB[29][13] ), .IN1(\mult_26/SUMB[29][14] ), .COUT(
        \mult_26/CARRYB[30][13] ), .SUM(\mult_26/SUMB[30][13] ) );
  FADDER \mult_26/S2_30_12  ( .CIN(\mult_26/ab[30][12] ), .IN0(
        \mult_26/CARRYB[29][12] ), .IN1(\mult_26/SUMB[29][13] ), .COUT(
        \mult_26/CARRYB[30][12] ), .SUM(\mult_26/SUMB[30][12] ) );
  FADDER \mult_26/S2_30_11  ( .CIN(\mult_26/ab[30][11] ), .IN0(
        \mult_26/CARRYB[29][11] ), .IN1(\mult_26/SUMB[29][12] ), .COUT(
        \mult_26/CARRYB[30][11] ), .SUM(\mult_26/SUMB[30][11] ) );
  FADDER \mult_26/S2_30_10  ( .CIN(\mult_26/ab[30][10] ), .IN0(
        \mult_26/CARRYB[29][10] ), .IN1(\mult_26/SUMB[29][11] ), .COUT(
        \mult_26/CARRYB[30][10] ), .SUM(\mult_26/SUMB[30][10] ) );
  FADDER \mult_26/S2_30_9  ( .CIN(\mult_26/ab[30][9] ), .IN0(
        \mult_26/CARRYB[29][9] ), .IN1(\mult_26/SUMB[29][10] ), .COUT(
        \mult_26/CARRYB[30][9] ), .SUM(\mult_26/SUMB[30][9] ) );
  FADDER \mult_26/S2_30_8  ( .CIN(\mult_26/ab[30][8] ), .IN0(
        \mult_26/CARRYB[29][8] ), .IN1(\mult_26/SUMB[29][9] ), .COUT(
        \mult_26/CARRYB[30][8] ), .SUM(\mult_26/SUMB[30][8] ) );
  FADDER \mult_26/S2_30_7  ( .CIN(\mult_26/ab[30][7] ), .IN0(
        \mult_26/CARRYB[29][7] ), .IN1(\mult_26/SUMB[29][8] ), .COUT(
        \mult_26/CARRYB[30][7] ), .SUM(\mult_26/SUMB[30][7] ) );
  FADDER \mult_26/S2_30_6  ( .CIN(\mult_26/ab[30][6] ), .IN0(
        \mult_26/CARRYB[29][6] ), .IN1(\mult_26/SUMB[29][7] ), .COUT(
        \mult_26/CARRYB[30][6] ), .SUM(\mult_26/SUMB[30][6] ) );
  FADDER \mult_26/S2_30_5  ( .CIN(\mult_26/ab[30][5] ), .IN0(
        \mult_26/CARRYB[29][5] ), .IN1(\mult_26/SUMB[29][6] ), .COUT(
        \mult_26/CARRYB[30][5] ), .SUM(\mult_26/SUMB[30][5] ) );
  FADDER \mult_26/S2_30_4  ( .CIN(\mult_26/ab[30][4] ), .IN0(
        \mult_26/CARRYB[29][4] ), .IN1(\mult_26/SUMB[29][5] ), .COUT(
        \mult_26/CARRYB[30][4] ), .SUM(\mult_26/SUMB[30][4] ) );
  FADDER \mult_26/S2_30_3  ( .CIN(\mult_26/ab[30][3] ), .IN0(
        \mult_26/CARRYB[29][3] ), .IN1(\mult_26/SUMB[29][4] ), .COUT(
        \mult_26/CARRYB[30][3] ), .SUM(\mult_26/SUMB[30][3] ) );
  FADDER \mult_26/S2_30_2  ( .CIN(\mult_26/ab[30][2] ), .IN0(
        \mult_26/CARRYB[29][2] ), .IN1(\mult_26/SUMB[29][3] ), .COUT(
        \mult_26/CARRYB[30][2] ), .SUM(\mult_26/SUMB[30][2] ) );
  FADDER \mult_26/S2_30_1  ( .CIN(\mult_26/ab[30][1] ), .IN0(
        \mult_26/CARRYB[29][1] ), .IN1(\mult_26/SUMB[29][2] ), .COUT(
        \mult_26/CARRYB[30][1] ), .SUM(\mult_26/SUMB[30][1] ) );
  FADDER \mult_26/S1_30_0  ( .CIN(\mult_26/ab[30][0] ), .IN0(
        \mult_26/CARRYB[29][0] ), .IN1(\mult_26/SUMB[29][1] ), .COUT(
        \mult_26/CARRYB[30][0] ), .SUM(o[30]) );
  FADDER \mult_26/S5_30  ( .CIN(\mult_26/ab[31][30] ), .IN0(
        \mult_26/CARRYB[30][30] ), .IN1(\mult_26/ab[30][31] ), .COUT(
        \mult_26/CARRYB[31][30] ), .SUM(\mult_26/SUMB[31][30] ) );
  FADDER \mult_26/S4_29  ( .CIN(\mult_26/ab[31][29] ), .IN0(
        \mult_26/CARRYB[30][29] ), .IN1(\mult_26/SUMB[30][30] ), .COUT(
        \mult_26/CARRYB[31][29] ), .SUM(\mult_26/SUMB[31][29] ) );
  FADDER \mult_26/S4_28  ( .CIN(\mult_26/ab[31][28] ), .IN0(
        \mult_26/CARRYB[30][28] ), .IN1(\mult_26/SUMB[30][29] ), .COUT(
        \mult_26/CARRYB[31][28] ), .SUM(\mult_26/SUMB[31][28] ) );
  FADDER \mult_26/S4_27  ( .CIN(\mult_26/ab[31][27] ), .IN0(
        \mult_26/CARRYB[30][27] ), .IN1(\mult_26/SUMB[30][28] ), .COUT(
        \mult_26/CARRYB[31][27] ), .SUM(\mult_26/SUMB[31][27] ) );
  FADDER \mult_26/S4_26  ( .CIN(\mult_26/ab[31][26] ), .IN0(
        \mult_26/CARRYB[30][26] ), .IN1(\mult_26/SUMB[30][27] ), .COUT(
        \mult_26/CARRYB[31][26] ), .SUM(\mult_26/SUMB[31][26] ) );
  FADDER \mult_26/S4_25  ( .CIN(\mult_26/ab[31][25] ), .IN0(
        \mult_26/CARRYB[30][25] ), .IN1(\mult_26/SUMB[30][26] ), .COUT(
        \mult_26/CARRYB[31][25] ), .SUM(\mult_26/SUMB[31][25] ) );
  FADDER \mult_26/S4_24  ( .CIN(\mult_26/ab[31][24] ), .IN0(
        \mult_26/CARRYB[30][24] ), .IN1(\mult_26/SUMB[30][25] ), .COUT(
        \mult_26/CARRYB[31][24] ), .SUM(\mult_26/SUMB[31][24] ) );
  FADDER \mult_26/S4_23  ( .CIN(\mult_26/ab[31][23] ), .IN0(
        \mult_26/CARRYB[30][23] ), .IN1(\mult_26/SUMB[30][24] ), .COUT(
        \mult_26/CARRYB[31][23] ), .SUM(\mult_26/SUMB[31][23] ) );
  FADDER \mult_26/S4_22  ( .CIN(\mult_26/ab[31][22] ), .IN0(
        \mult_26/CARRYB[30][22] ), .IN1(\mult_26/SUMB[30][23] ), .COUT(
        \mult_26/CARRYB[31][22] ), .SUM(\mult_26/SUMB[31][22] ) );
  FADDER \mult_26/S4_21  ( .CIN(\mult_26/ab[31][21] ), .IN0(
        \mult_26/CARRYB[30][21] ), .IN1(\mult_26/SUMB[30][22] ), .COUT(
        \mult_26/CARRYB[31][21] ), .SUM(\mult_26/SUMB[31][21] ) );
  FADDER \mult_26/S4_20  ( .CIN(\mult_26/ab[31][20] ), .IN0(
        \mult_26/CARRYB[30][20] ), .IN1(\mult_26/SUMB[30][21] ), .COUT(
        \mult_26/CARRYB[31][20] ), .SUM(\mult_26/SUMB[31][20] ) );
  FADDER \mult_26/S4_19  ( .CIN(\mult_26/ab[31][19] ), .IN0(
        \mult_26/CARRYB[30][19] ), .IN1(\mult_26/SUMB[30][20] ), .COUT(
        \mult_26/CARRYB[31][19] ), .SUM(\mult_26/SUMB[31][19] ) );
  FADDER \mult_26/S4_18  ( .CIN(\mult_26/ab[31][18] ), .IN0(
        \mult_26/CARRYB[30][18] ), .IN1(\mult_26/SUMB[30][19] ), .COUT(
        \mult_26/CARRYB[31][18] ), .SUM(\mult_26/SUMB[31][18] ) );
  FADDER \mult_26/S4_17  ( .CIN(\mult_26/ab[31][17] ), .IN0(
        \mult_26/CARRYB[30][17] ), .IN1(\mult_26/SUMB[30][18] ), .COUT(
        \mult_26/CARRYB[31][17] ), .SUM(\mult_26/SUMB[31][17] ) );
  FADDER \mult_26/S4_16  ( .CIN(\mult_26/ab[31][16] ), .IN0(
        \mult_26/CARRYB[30][16] ), .IN1(\mult_26/SUMB[30][17] ), .COUT(
        \mult_26/CARRYB[31][16] ), .SUM(\mult_26/SUMB[31][16] ) );
  FADDER \mult_26/S4_15  ( .CIN(\mult_26/ab[31][15] ), .IN0(
        \mult_26/CARRYB[30][15] ), .IN1(\mult_26/SUMB[30][16] ), .COUT(
        \mult_26/CARRYB[31][15] ), .SUM(\mult_26/SUMB[31][15] ) );
  FADDER \mult_26/S4_14  ( .CIN(\mult_26/ab[31][14] ), .IN0(
        \mult_26/CARRYB[30][14] ), .IN1(\mult_26/SUMB[30][15] ), .COUT(
        \mult_26/CARRYB[31][14] ), .SUM(\mult_26/SUMB[31][14] ) );
  FADDER \mult_26/S4_13  ( .CIN(\mult_26/ab[31][13] ), .IN0(
        \mult_26/CARRYB[30][13] ), .IN1(\mult_26/SUMB[30][14] ), .COUT(
        \mult_26/CARRYB[31][13] ), .SUM(\mult_26/SUMB[31][13] ) );
  FADDER \mult_26/S4_12  ( .CIN(\mult_26/ab[31][12] ), .IN0(
        \mult_26/CARRYB[30][12] ), .IN1(\mult_26/SUMB[30][13] ), .COUT(
        \mult_26/CARRYB[31][12] ), .SUM(\mult_26/SUMB[31][12] ) );
  FADDER \mult_26/S4_11  ( .CIN(\mult_26/ab[31][11] ), .IN0(
        \mult_26/CARRYB[30][11] ), .IN1(\mult_26/SUMB[30][12] ), .COUT(
        \mult_26/CARRYB[31][11] ), .SUM(\mult_26/SUMB[31][11] ) );
  FADDER \mult_26/S4_10  ( .CIN(\mult_26/ab[31][10] ), .IN0(
        \mult_26/CARRYB[30][10] ), .IN1(\mult_26/SUMB[30][11] ), .COUT(
        \mult_26/CARRYB[31][10] ), .SUM(\mult_26/SUMB[31][10] ) );
  FADDER \mult_26/S4_9  ( .CIN(\mult_26/ab[31][9] ), .IN0(
        \mult_26/CARRYB[30][9] ), .IN1(\mult_26/SUMB[30][10] ), .COUT(
        \mult_26/CARRYB[31][9] ), .SUM(\mult_26/SUMB[31][9] ) );
  FADDER \mult_26/S4_8  ( .CIN(\mult_26/ab[31][8] ), .IN0(
        \mult_26/CARRYB[30][8] ), .IN1(\mult_26/SUMB[30][9] ), .COUT(
        \mult_26/CARRYB[31][8] ), .SUM(\mult_26/SUMB[31][8] ) );
  FADDER \mult_26/S4_7  ( .CIN(\mult_26/ab[31][7] ), .IN0(
        \mult_26/CARRYB[30][7] ), .IN1(\mult_26/SUMB[30][8] ), .COUT(
        \mult_26/CARRYB[31][7] ), .SUM(\mult_26/SUMB[31][7] ) );
  FADDER \mult_26/S4_6  ( .CIN(\mult_26/ab[31][6] ), .IN0(
        \mult_26/CARRYB[30][6] ), .IN1(\mult_26/SUMB[30][7] ), .COUT(
        \mult_26/CARRYB[31][6] ), .SUM(\mult_26/SUMB[31][6] ) );
  FADDER \mult_26/S4_5  ( .CIN(\mult_26/ab[31][5] ), .IN0(
        \mult_26/CARRYB[30][5] ), .IN1(\mult_26/SUMB[30][6] ), .COUT(
        \mult_26/CARRYB[31][5] ), .SUM(\mult_26/SUMB[31][5] ) );
  FADDER \mult_26/S4_4  ( .CIN(\mult_26/ab[31][4] ), .IN0(
        \mult_26/CARRYB[30][4] ), .IN1(\mult_26/SUMB[30][5] ), .COUT(
        \mult_26/CARRYB[31][4] ), .SUM(\mult_26/SUMB[31][4] ) );
  FADDER \mult_26/S4_3  ( .CIN(\mult_26/ab[31][3] ), .IN0(
        \mult_26/CARRYB[30][3] ), .IN1(\mult_26/SUMB[30][4] ), .COUT(
        \mult_26/CARRYB[31][3] ), .SUM(\mult_26/SUMB[31][3] ) );
  FADDER \mult_26/S4_2  ( .CIN(\mult_26/ab[31][2] ), .IN0(
        \mult_26/CARRYB[30][2] ), .IN1(\mult_26/SUMB[30][3] ), .COUT(
        \mult_26/CARRYB[31][2] ), .SUM(\mult_26/SUMB[31][2] ) );
  FADDER \mult_26/S4_1  ( .CIN(\mult_26/ab[31][1] ), .IN0(
        \mult_26/CARRYB[30][1] ), .IN1(\mult_26/SUMB[30][2] ), .COUT(
        \mult_26/CARRYB[31][1] ), .SUM(\mult_26/SUMB[31][1] ) );
  FADDER \mult_26/S4_0  ( .CIN(\mult_26/ab[31][0] ), .IN0(
        \mult_26/CARRYB[30][0] ), .IN1(\mult_26/SUMB[30][1] ), .COUT(
        \mult_26/CARRYB[31][0] ), .SUM(\mult_26/SUMB[31][0] ) );
  XNOR U2 ( .A(\mult_26/A2[33] ), .B(\mult_26/A1[33] ), .Z(n184) );
  XNOR U3 ( .A(\mult_26/A2[37] ), .B(\mult_26/A1[37] ), .Z(n157) );
  XNOR U4 ( .A(\mult_26/A2[41] ), .B(\mult_26/A1[41] ), .Z(n130) );
  XNOR U5 ( .A(\mult_26/A1[45] ), .B(\mult_26/A2[45] ), .Z(n102) );
  XOR U6 ( .A(\mult_26/A2[31] ), .B(\mult_26/A1[31] ), .Z(o[33]) );
  XNOR U7 ( .A(\mult_26/A2[34] ), .B(\mult_26/A1[34] ), .Z(n181) );
  XNOR U8 ( .A(\mult_26/A2[38] ), .B(\mult_26/A1[38] ), .Z(n154) );
  XNOR U9 ( .A(\mult_26/A2[42] ), .B(\mult_26/A1[42] ), .Z(n127) );
  XNOR U10 ( .A(\mult_26/A1[47] ), .B(\mult_26/A2[47] ), .Z(n95) );
  XNOR U11 ( .A(\mult_26/A2[49] ), .B(\mult_26/A1[49] ), .Z(n62) );
  XNOR U12 ( .A(\mult_26/A2[51] ), .B(\mult_26/A1[51] ), .Z(n52) );
  XNOR U13 ( .A(\mult_26/A2[53] ), .B(\mult_26/A1[53] ), .Z(n42) );
  XNOR U14 ( .A(\mult_26/A2[55] ), .B(\mult_26/A1[55] ), .Z(n32) );
  XNOR U15 ( .A(\mult_26/A2[57] ), .B(\mult_26/A1[57] ), .Z(n22) );
  XNOR U16 ( .A(\mult_26/A2[59] ), .B(\mult_26/A1[59] ), .Z(n12) );
  XOR U17 ( .A(\mult_26/A1[32] ), .B(\mult_26/A2[32] ), .Z(n186) );
  XNOR U18 ( .A(\mult_26/A2[35] ), .B(\mult_26/A1[35] ), .Z(n177) );
  XNOR U19 ( .A(\mult_26/A1[36] ), .B(\mult_26/A2[36] ), .Z(n159) );
  XNOR U20 ( .A(\mult_26/A2[39] ), .B(\mult_26/A1[39] ), .Z(n150) );
  XNOR U21 ( .A(\mult_26/A2[40] ), .B(\mult_26/A1[40] ), .Z(n132) );
  XNOR U22 ( .A(\mult_26/A2[43] ), .B(\mult_26/A1[43] ), .Z(n123) );
  XNOR U23 ( .A(\mult_26/A1[44] ), .B(\mult_26/A2[44] ), .Z(n105) );
  XNOR U24 ( .A(\mult_26/A1[46] ), .B(\mult_26/A2[46] ), .Z(n99) );
  XNOR U25 ( .A(\mult_26/A2[48] ), .B(\mult_26/A1[48] ), .Z(n67) );
  XNOR U26 ( .A(\mult_26/A2[50] ), .B(\mult_26/A1[50] ), .Z(n57) );
  XNOR U27 ( .A(\mult_26/A2[52] ), .B(\mult_26/A1[52] ), .Z(n47) );
  XNOR U28 ( .A(\mult_26/A2[54] ), .B(\mult_26/A1[54] ), .Z(n37) );
  XNOR U29 ( .A(\mult_26/A2[56] ), .B(\mult_26/A1[56] ), .Z(n27) );
  XNOR U30 ( .A(\mult_26/A2[58] ), .B(\mult_26/A1[58] ), .Z(n17) );
  XNOR U31 ( .A(\mult_26/A2[60] ), .B(\mult_26/A1[60] ), .Z(n7) );
  AND U32 ( .A(\mult_26/CARRYB[31][0] ), .B(\mult_26/SUMB[31][1] ), .Z(
        \mult_26/A2[31] ) );
  XOR U33 ( .A(\mult_26/SUMB[31][1] ), .B(\mult_26/CARRYB[31][0] ), .Z(o[32])
         );
  AND U34 ( .A(\mult_26/SUMB[31][2] ), .B(\mult_26/CARRYB[31][1] ), .Z(
        \mult_26/A2[32] ) );
  XOR U35 ( .A(\mult_26/SUMB[31][2] ), .B(\mult_26/CARRYB[31][1] ), .Z(
        \mult_26/A1[31] ) );
  AND U36 ( .A(\mult_26/SUMB[31][3] ), .B(\mult_26/CARRYB[31][2] ), .Z(
        \mult_26/A2[33] ) );
  XOR U37 ( .A(\mult_26/SUMB[31][3] ), .B(\mult_26/CARRYB[31][2] ), .Z(
        \mult_26/A1[32] ) );
  AND U38 ( .A(\mult_26/SUMB[31][4] ), .B(\mult_26/CARRYB[31][3] ), .Z(
        \mult_26/A2[34] ) );
  XOR U39 ( .A(\mult_26/SUMB[31][4] ), .B(\mult_26/CARRYB[31][3] ), .Z(
        \mult_26/A1[33] ) );
  AND U40 ( .A(\mult_26/SUMB[31][5] ), .B(\mult_26/CARRYB[31][4] ), .Z(
        \mult_26/A2[35] ) );
  XOR U41 ( .A(\mult_26/SUMB[31][5] ), .B(\mult_26/CARRYB[31][4] ), .Z(
        \mult_26/A1[34] ) );
  AND U42 ( .A(\mult_26/SUMB[31][6] ), .B(\mult_26/CARRYB[31][5] ), .Z(
        \mult_26/A2[36] ) );
  XOR U43 ( .A(\mult_26/SUMB[31][6] ), .B(\mult_26/CARRYB[31][5] ), .Z(
        \mult_26/A1[35] ) );
  AND U44 ( .A(\mult_26/SUMB[31][7] ), .B(\mult_26/CARRYB[31][6] ), .Z(
        \mult_26/A2[37] ) );
  XOR U45 ( .A(\mult_26/SUMB[31][7] ), .B(\mult_26/CARRYB[31][6] ), .Z(
        \mult_26/A1[36] ) );
  AND U46 ( .A(\mult_26/SUMB[31][8] ), .B(\mult_26/CARRYB[31][7] ), .Z(
        \mult_26/A2[38] ) );
  XOR U47 ( .A(\mult_26/SUMB[31][8] ), .B(\mult_26/CARRYB[31][7] ), .Z(
        \mult_26/A1[37] ) );
  AND U48 ( .A(\mult_26/SUMB[31][9] ), .B(\mult_26/CARRYB[31][8] ), .Z(
        \mult_26/A2[39] ) );
  XOR U49 ( .A(\mult_26/SUMB[31][9] ), .B(\mult_26/CARRYB[31][8] ), .Z(
        \mult_26/A1[38] ) );
  AND U50 ( .A(\mult_26/SUMB[31][10] ), .B(\mult_26/CARRYB[31][9] ), .Z(
        \mult_26/A2[40] ) );
  XOR U51 ( .A(\mult_26/SUMB[31][10] ), .B(\mult_26/CARRYB[31][9] ), .Z(
        \mult_26/A1[39] ) );
  AND U52 ( .A(\mult_26/SUMB[31][11] ), .B(\mult_26/CARRYB[31][10] ), .Z(
        \mult_26/A2[41] ) );
  XOR U53 ( .A(\mult_26/SUMB[31][11] ), .B(\mult_26/CARRYB[31][10] ), .Z(
        \mult_26/A1[40] ) );
  AND U54 ( .A(\mult_26/SUMB[31][12] ), .B(\mult_26/CARRYB[31][11] ), .Z(
        \mult_26/A2[42] ) );
  XOR U55 ( .A(\mult_26/SUMB[31][12] ), .B(\mult_26/CARRYB[31][11] ), .Z(
        \mult_26/A1[41] ) );
  AND U56 ( .A(\mult_26/SUMB[31][13] ), .B(\mult_26/CARRYB[31][12] ), .Z(
        \mult_26/A2[43] ) );
  XOR U57 ( .A(\mult_26/SUMB[31][13] ), .B(\mult_26/CARRYB[31][12] ), .Z(
        \mult_26/A1[42] ) );
  AND U58 ( .A(\mult_26/SUMB[31][14] ), .B(\mult_26/CARRYB[31][13] ), .Z(
        \mult_26/A2[44] ) );
  XOR U59 ( .A(\mult_26/SUMB[31][14] ), .B(\mult_26/CARRYB[31][13] ), .Z(
        \mult_26/A1[43] ) );
  AND U60 ( .A(\mult_26/SUMB[31][15] ), .B(\mult_26/CARRYB[31][14] ), .Z(
        \mult_26/A2[45] ) );
  XOR U61 ( .A(\mult_26/SUMB[31][15] ), .B(\mult_26/CARRYB[31][14] ), .Z(
        \mult_26/A1[44] ) );
  AND U62 ( .A(\mult_26/SUMB[31][16] ), .B(\mult_26/CARRYB[31][15] ), .Z(
        \mult_26/A2[46] ) );
  XOR U63 ( .A(\mult_26/SUMB[31][16] ), .B(\mult_26/CARRYB[31][15] ), .Z(
        \mult_26/A1[45] ) );
  AND U64 ( .A(\mult_26/SUMB[31][17] ), .B(\mult_26/CARRYB[31][16] ), .Z(
        \mult_26/A2[47] ) );
  XOR U65 ( .A(\mult_26/SUMB[31][17] ), .B(\mult_26/CARRYB[31][16] ), .Z(
        \mult_26/A1[46] ) );
  AND U66 ( .A(\mult_26/SUMB[31][18] ), .B(\mult_26/CARRYB[31][17] ), .Z(
        \mult_26/A2[48] ) );
  XOR U67 ( .A(\mult_26/SUMB[31][18] ), .B(\mult_26/CARRYB[31][17] ), .Z(
        \mult_26/A1[47] ) );
  AND U68 ( .A(\mult_26/SUMB[31][19] ), .B(\mult_26/CARRYB[31][18] ), .Z(
        \mult_26/A2[49] ) );
  XOR U69 ( .A(\mult_26/SUMB[31][19] ), .B(\mult_26/CARRYB[31][18] ), .Z(
        \mult_26/A1[48] ) );
  AND U70 ( .A(\mult_26/SUMB[31][20] ), .B(\mult_26/CARRYB[31][19] ), .Z(
        \mult_26/A2[50] ) );
  XOR U71 ( .A(\mult_26/SUMB[31][20] ), .B(\mult_26/CARRYB[31][19] ), .Z(
        \mult_26/A1[49] ) );
  AND U72 ( .A(\mult_26/SUMB[31][21] ), .B(\mult_26/CARRYB[31][20] ), .Z(
        \mult_26/A2[51] ) );
  XOR U73 ( .A(\mult_26/SUMB[31][21] ), .B(\mult_26/CARRYB[31][20] ), .Z(
        \mult_26/A1[50] ) );
  AND U74 ( .A(\mult_26/SUMB[31][22] ), .B(\mult_26/CARRYB[31][21] ), .Z(
        \mult_26/A2[52] ) );
  XOR U75 ( .A(\mult_26/SUMB[31][22] ), .B(\mult_26/CARRYB[31][21] ), .Z(
        \mult_26/A1[51] ) );
  AND U76 ( .A(\mult_26/SUMB[31][23] ), .B(\mult_26/CARRYB[31][22] ), .Z(
        \mult_26/A2[53] ) );
  XOR U77 ( .A(\mult_26/SUMB[31][23] ), .B(\mult_26/CARRYB[31][22] ), .Z(
        \mult_26/A1[52] ) );
  AND U78 ( .A(\mult_26/SUMB[31][24] ), .B(\mult_26/CARRYB[31][23] ), .Z(
        \mult_26/A2[54] ) );
  XOR U79 ( .A(\mult_26/SUMB[31][24] ), .B(\mult_26/CARRYB[31][23] ), .Z(
        \mult_26/A1[53] ) );
  AND U80 ( .A(\mult_26/SUMB[31][25] ), .B(\mult_26/CARRYB[31][24] ), .Z(
        \mult_26/A2[55] ) );
  XOR U81 ( .A(\mult_26/SUMB[31][25] ), .B(\mult_26/CARRYB[31][24] ), .Z(
        \mult_26/A1[54] ) );
  AND U82 ( .A(\mult_26/SUMB[31][26] ), .B(\mult_26/CARRYB[31][25] ), .Z(
        \mult_26/A2[56] ) );
  XOR U83 ( .A(\mult_26/SUMB[31][26] ), .B(\mult_26/CARRYB[31][25] ), .Z(
        \mult_26/A1[55] ) );
  AND U84 ( .A(\mult_26/SUMB[31][27] ), .B(\mult_26/CARRYB[31][26] ), .Z(
        \mult_26/A2[57] ) );
  XOR U85 ( .A(\mult_26/SUMB[31][27] ), .B(\mult_26/CARRYB[31][26] ), .Z(
        \mult_26/A1[56] ) );
  AND U86 ( .A(\mult_26/SUMB[31][28] ), .B(\mult_26/CARRYB[31][27] ), .Z(
        \mult_26/A2[58] ) );
  XOR U87 ( .A(\mult_26/SUMB[31][28] ), .B(\mult_26/CARRYB[31][27] ), .Z(
        \mult_26/A1[57] ) );
  AND U88 ( .A(\mult_26/SUMB[31][29] ), .B(\mult_26/CARRYB[31][28] ), .Z(
        \mult_26/A2[59] ) );
  XOR U89 ( .A(\mult_26/SUMB[31][29] ), .B(\mult_26/CARRYB[31][28] ), .Z(
        \mult_26/A1[58] ) );
  AND U90 ( .A(\mult_26/SUMB[31][30] ), .B(\mult_26/CARRYB[31][29] ), .Z(
        \mult_26/A2[60] ) );
  XOR U91 ( .A(\mult_26/SUMB[31][30] ), .B(\mult_26/CARRYB[31][29] ), .Z(
        \mult_26/A1[59] ) );
  AND U92 ( .A(\mult_26/ab[31][31] ), .B(\mult_26/CARRYB[31][30] ), .Z(
        \mult_26/A2[61] ) );
  XOR U93 ( .A(\mult_26/ab[31][31] ), .B(\mult_26/CARRYB[31][30] ), .Z(
        \mult_26/A1[60] ) );
  AND U94 ( .A(\mult_26/ab[1][0] ), .B(\mult_26/ab[0][1] ), .Z(
        \mult_26/CARRYB[1][0] ) );
  XOR U95 ( .A(\mult_26/ab[0][1] ), .B(\mult_26/ab[1][0] ), .Z(o[1]) );
  AND U96 ( .A(\mult_26/ab[1][1] ), .B(\mult_26/ab[0][2] ), .Z(
        \mult_26/CARRYB[1][1] ) );
  XOR U97 ( .A(\mult_26/ab[0][2] ), .B(\mult_26/ab[1][1] ), .Z(
        \mult_26/SUMB[1][1] ) );
  AND U98 ( .A(\mult_26/ab[1][2] ), .B(\mult_26/ab[0][3] ), .Z(
        \mult_26/CARRYB[1][2] ) );
  XOR U99 ( .A(\mult_26/ab[0][3] ), .B(\mult_26/ab[1][2] ), .Z(
        \mult_26/SUMB[1][2] ) );
  AND U100 ( .A(\mult_26/ab[1][3] ), .B(\mult_26/ab[0][4] ), .Z(
        \mult_26/CARRYB[1][3] ) );
  XOR U101 ( .A(\mult_26/ab[0][4] ), .B(\mult_26/ab[1][3] ), .Z(
        \mult_26/SUMB[1][3] ) );
  AND U102 ( .A(\mult_26/ab[1][4] ), .B(\mult_26/ab[0][5] ), .Z(
        \mult_26/CARRYB[1][4] ) );
  XOR U103 ( .A(\mult_26/ab[0][5] ), .B(\mult_26/ab[1][4] ), .Z(
        \mult_26/SUMB[1][4] ) );
  AND U104 ( .A(\mult_26/ab[1][5] ), .B(\mult_26/ab[0][6] ), .Z(
        \mult_26/CARRYB[1][5] ) );
  XOR U105 ( .A(\mult_26/ab[0][6] ), .B(\mult_26/ab[1][5] ), .Z(
        \mult_26/SUMB[1][5] ) );
  AND U106 ( .A(\mult_26/ab[1][6] ), .B(\mult_26/ab[0][7] ), .Z(
        \mult_26/CARRYB[1][6] ) );
  XOR U107 ( .A(\mult_26/ab[0][7] ), .B(\mult_26/ab[1][6] ), .Z(
        \mult_26/SUMB[1][6] ) );
  AND U108 ( .A(\mult_26/ab[1][7] ), .B(\mult_26/ab[0][8] ), .Z(
        \mult_26/CARRYB[1][7] ) );
  XOR U109 ( .A(\mult_26/ab[0][8] ), .B(\mult_26/ab[1][7] ), .Z(
        \mult_26/SUMB[1][7] ) );
  AND U110 ( .A(\mult_26/ab[1][8] ), .B(\mult_26/ab[0][9] ), .Z(
        \mult_26/CARRYB[1][8] ) );
  XOR U111 ( .A(\mult_26/ab[0][9] ), .B(\mult_26/ab[1][8] ), .Z(
        \mult_26/SUMB[1][8] ) );
  AND U112 ( .A(\mult_26/ab[1][9] ), .B(\mult_26/ab[0][10] ), .Z(
        \mult_26/CARRYB[1][9] ) );
  XOR U113 ( .A(\mult_26/ab[0][10] ), .B(\mult_26/ab[1][9] ), .Z(
        \mult_26/SUMB[1][9] ) );
  AND U114 ( .A(\mult_26/ab[1][10] ), .B(\mult_26/ab[0][11] ), .Z(
        \mult_26/CARRYB[1][10] ) );
  XOR U115 ( .A(\mult_26/ab[0][11] ), .B(\mult_26/ab[1][10] ), .Z(
        \mult_26/SUMB[1][10] ) );
  AND U116 ( .A(\mult_26/ab[1][11] ), .B(\mult_26/ab[0][12] ), .Z(
        \mult_26/CARRYB[1][11] ) );
  XOR U117 ( .A(\mult_26/ab[0][12] ), .B(\mult_26/ab[1][11] ), .Z(
        \mult_26/SUMB[1][11] ) );
  AND U118 ( .A(\mult_26/ab[1][12] ), .B(\mult_26/ab[0][13] ), .Z(
        \mult_26/CARRYB[1][12] ) );
  XOR U119 ( .A(\mult_26/ab[0][13] ), .B(\mult_26/ab[1][12] ), .Z(
        \mult_26/SUMB[1][12] ) );
  AND U120 ( .A(\mult_26/ab[1][13] ), .B(\mult_26/ab[0][14] ), .Z(
        \mult_26/CARRYB[1][13] ) );
  XOR U121 ( .A(\mult_26/ab[0][14] ), .B(\mult_26/ab[1][13] ), .Z(
        \mult_26/SUMB[1][13] ) );
  AND U122 ( .A(\mult_26/ab[1][14] ), .B(\mult_26/ab[0][15] ), .Z(
        \mult_26/CARRYB[1][14] ) );
  XOR U123 ( .A(\mult_26/ab[0][15] ), .B(\mult_26/ab[1][14] ), .Z(
        \mult_26/SUMB[1][14] ) );
  AND U124 ( .A(\mult_26/ab[1][15] ), .B(\mult_26/ab[0][16] ), .Z(
        \mult_26/CARRYB[1][15] ) );
  XOR U125 ( .A(\mult_26/ab[0][16] ), .B(\mult_26/ab[1][15] ), .Z(
        \mult_26/SUMB[1][15] ) );
  AND U126 ( .A(\mult_26/ab[1][16] ), .B(\mult_26/ab[0][17] ), .Z(
        \mult_26/CARRYB[1][16] ) );
  XOR U127 ( .A(\mult_26/ab[0][17] ), .B(\mult_26/ab[1][16] ), .Z(
        \mult_26/SUMB[1][16] ) );
  AND U128 ( .A(\mult_26/ab[1][17] ), .B(\mult_26/ab[0][18] ), .Z(
        \mult_26/CARRYB[1][17] ) );
  XOR U129 ( .A(\mult_26/ab[0][18] ), .B(\mult_26/ab[1][17] ), .Z(
        \mult_26/SUMB[1][17] ) );
  AND U130 ( .A(\mult_26/ab[1][18] ), .B(\mult_26/ab[0][19] ), .Z(
        \mult_26/CARRYB[1][18] ) );
  XOR U131 ( .A(\mult_26/ab[0][19] ), .B(\mult_26/ab[1][18] ), .Z(
        \mult_26/SUMB[1][18] ) );
  AND U132 ( .A(\mult_26/ab[1][19] ), .B(\mult_26/ab[0][20] ), .Z(
        \mult_26/CARRYB[1][19] ) );
  XOR U133 ( .A(\mult_26/ab[0][20] ), .B(\mult_26/ab[1][19] ), .Z(
        \mult_26/SUMB[1][19] ) );
  AND U134 ( .A(\mult_26/ab[1][20] ), .B(\mult_26/ab[0][21] ), .Z(
        \mult_26/CARRYB[1][20] ) );
  XOR U135 ( .A(\mult_26/ab[0][21] ), .B(\mult_26/ab[1][20] ), .Z(
        \mult_26/SUMB[1][20] ) );
  AND U136 ( .A(\mult_26/ab[1][21] ), .B(\mult_26/ab[0][22] ), .Z(
        \mult_26/CARRYB[1][21] ) );
  XOR U137 ( .A(\mult_26/ab[0][22] ), .B(\mult_26/ab[1][21] ), .Z(
        \mult_26/SUMB[1][21] ) );
  AND U138 ( .A(\mult_26/ab[1][22] ), .B(\mult_26/ab[0][23] ), .Z(
        \mult_26/CARRYB[1][22] ) );
  XOR U139 ( .A(\mult_26/ab[0][23] ), .B(\mult_26/ab[1][22] ), .Z(
        \mult_26/SUMB[1][22] ) );
  AND U140 ( .A(\mult_26/ab[1][23] ), .B(\mult_26/ab[0][24] ), .Z(
        \mult_26/CARRYB[1][23] ) );
  XOR U141 ( .A(\mult_26/ab[0][24] ), .B(\mult_26/ab[1][23] ), .Z(
        \mult_26/SUMB[1][23] ) );
  AND U142 ( .A(\mult_26/ab[1][24] ), .B(\mult_26/ab[0][25] ), .Z(
        \mult_26/CARRYB[1][24] ) );
  XOR U143 ( .A(\mult_26/ab[0][25] ), .B(\mult_26/ab[1][24] ), .Z(
        \mult_26/SUMB[1][24] ) );
  AND U144 ( .A(\mult_26/ab[1][25] ), .B(\mult_26/ab[0][26] ), .Z(
        \mult_26/CARRYB[1][25] ) );
  XOR U145 ( .A(\mult_26/ab[0][26] ), .B(\mult_26/ab[1][25] ), .Z(
        \mult_26/SUMB[1][25] ) );
  AND U146 ( .A(\mult_26/ab[1][26] ), .B(\mult_26/ab[0][27] ), .Z(
        \mult_26/CARRYB[1][26] ) );
  XOR U147 ( .A(\mult_26/ab[0][27] ), .B(\mult_26/ab[1][26] ), .Z(
        \mult_26/SUMB[1][26] ) );
  AND U148 ( .A(\mult_26/ab[1][27] ), .B(\mult_26/ab[0][28] ), .Z(
        \mult_26/CARRYB[1][27] ) );
  XOR U149 ( .A(\mult_26/ab[0][28] ), .B(\mult_26/ab[1][27] ), .Z(
        \mult_26/SUMB[1][27] ) );
  AND U150 ( .A(\mult_26/ab[1][28] ), .B(\mult_26/ab[0][29] ), .Z(
        \mult_26/CARRYB[1][28] ) );
  XOR U151 ( .A(\mult_26/ab[0][29] ), .B(\mult_26/ab[1][28] ), .Z(
        \mult_26/SUMB[1][28] ) );
  AND U152 ( .A(\mult_26/ab[1][29] ), .B(\mult_26/ab[0][30] ), .Z(
        \mult_26/CARRYB[1][29] ) );
  XOR U153 ( .A(\mult_26/ab[0][30] ), .B(\mult_26/ab[1][29] ), .Z(
        \mult_26/SUMB[1][29] ) );
  AND U154 ( .A(\mult_26/ab[1][30] ), .B(\mult_26/ab[0][31] ), .Z(
        \mult_26/CARRYB[1][30] ) );
  XOR U155 ( .A(\mult_26/ab[0][31] ), .B(\mult_26/ab[1][30] ), .Z(
        \mult_26/SUMB[1][30] ) );
  XOR U156 ( .A(n2), .B(\mult_26/A2[61] ), .Z(o[63]) );
  NANDN U157 ( .B(n3), .A(n4), .Z(n2) );
  NAND U158 ( .A(n5), .B(n6), .Z(n4) );
  XNOR U159 ( .A(n7), .B(n5), .Z(o[62]) );
  NANDN U160 ( .B(n8), .A(n9), .Z(n5) );
  NAND U161 ( .A(n10), .B(n11), .Z(n9) );
  OR U162 ( .A(\mult_26/A2[60] ), .B(\mult_26/A1[60] ), .Z(n6) );
  AND U163 ( .A(\mult_26/A2[60] ), .B(\mult_26/A1[60] ), .Z(n3) );
  XNOR U164 ( .A(n12), .B(n10), .Z(o[61]) );
  NANDN U165 ( .B(n13), .A(n14), .Z(n10) );
  NAND U166 ( .A(n15), .B(n16), .Z(n14) );
  OR U167 ( .A(\mult_26/A2[59] ), .B(\mult_26/A1[59] ), .Z(n11) );
  AND U168 ( .A(\mult_26/A2[59] ), .B(\mult_26/A1[59] ), .Z(n8) );
  XNOR U169 ( .A(n17), .B(n15), .Z(o[60]) );
  NANDN U170 ( .B(n18), .A(n19), .Z(n15) );
  NAND U171 ( .A(n20), .B(n21), .Z(n19) );
  OR U172 ( .A(\mult_26/A2[58] ), .B(\mult_26/A1[58] ), .Z(n16) );
  AND U173 ( .A(\mult_26/A2[58] ), .B(\mult_26/A1[58] ), .Z(n13) );
  XNOR U174 ( .A(n22), .B(n20), .Z(o[59]) );
  NANDN U175 ( .B(n23), .A(n24), .Z(n20) );
  NAND U176 ( .A(n25), .B(n26), .Z(n24) );
  OR U177 ( .A(\mult_26/A2[57] ), .B(\mult_26/A1[57] ), .Z(n21) );
  AND U178 ( .A(\mult_26/A2[57] ), .B(\mult_26/A1[57] ), .Z(n18) );
  XNOR U179 ( .A(n27), .B(n25), .Z(o[58]) );
  NANDN U180 ( .B(n28), .A(n29), .Z(n25) );
  NAND U181 ( .A(n30), .B(n31), .Z(n29) );
  OR U182 ( .A(\mult_26/A2[56] ), .B(\mult_26/A1[56] ), .Z(n26) );
  AND U183 ( .A(\mult_26/A2[56] ), .B(\mult_26/A1[56] ), .Z(n23) );
  XNOR U184 ( .A(n32), .B(n30), .Z(o[57]) );
  NANDN U185 ( .B(n33), .A(n34), .Z(n30) );
  NAND U186 ( .A(n35), .B(n36), .Z(n34) );
  OR U187 ( .A(\mult_26/A2[55] ), .B(\mult_26/A1[55] ), .Z(n31) );
  AND U188 ( .A(\mult_26/A2[55] ), .B(\mult_26/A1[55] ), .Z(n28) );
  XNOR U189 ( .A(n37), .B(n35), .Z(o[56]) );
  NANDN U190 ( .B(n38), .A(n39), .Z(n35) );
  NAND U191 ( .A(n40), .B(n41), .Z(n39) );
  OR U192 ( .A(\mult_26/A2[54] ), .B(\mult_26/A1[54] ), .Z(n36) );
  AND U193 ( .A(\mult_26/A2[54] ), .B(\mult_26/A1[54] ), .Z(n33) );
  XNOR U194 ( .A(n42), .B(n40), .Z(o[55]) );
  NANDN U195 ( .B(n43), .A(n44), .Z(n40) );
  NAND U196 ( .A(n45), .B(n46), .Z(n44) );
  OR U197 ( .A(\mult_26/A2[53] ), .B(\mult_26/A1[53] ), .Z(n41) );
  AND U198 ( .A(\mult_26/A2[53] ), .B(\mult_26/A1[53] ), .Z(n38) );
  XNOR U199 ( .A(n47), .B(n45), .Z(o[54]) );
  NANDN U200 ( .B(n48), .A(n49), .Z(n45) );
  NAND U201 ( .A(n50), .B(n51), .Z(n49) );
  OR U202 ( .A(\mult_26/A2[52] ), .B(\mult_26/A1[52] ), .Z(n46) );
  AND U203 ( .A(\mult_26/A2[52] ), .B(\mult_26/A1[52] ), .Z(n43) );
  XNOR U204 ( .A(n52), .B(n50), .Z(o[53]) );
  NANDN U205 ( .B(n53), .A(n54), .Z(n50) );
  NAND U206 ( .A(n55), .B(n56), .Z(n54) );
  OR U207 ( .A(\mult_26/A2[51] ), .B(\mult_26/A1[51] ), .Z(n51) );
  AND U208 ( .A(\mult_26/A2[51] ), .B(\mult_26/A1[51] ), .Z(n48) );
  XNOR U209 ( .A(n57), .B(n55), .Z(o[52]) );
  NANDN U210 ( .B(n58), .A(n59), .Z(n55) );
  NAND U211 ( .A(n60), .B(n61), .Z(n59) );
  OR U212 ( .A(\mult_26/A2[50] ), .B(\mult_26/A1[50] ), .Z(n56) );
  AND U213 ( .A(\mult_26/A2[50] ), .B(\mult_26/A1[50] ), .Z(n53) );
  XNOR U214 ( .A(n62), .B(n60), .Z(o[51]) );
  NANDN U215 ( .B(n63), .A(n64), .Z(n60) );
  NAND U216 ( .A(n65), .B(n66), .Z(n64) );
  OR U217 ( .A(\mult_26/A2[49] ), .B(\mult_26/A1[49] ), .Z(n61) );
  AND U218 ( .A(\mult_26/A2[49] ), .B(\mult_26/A1[49] ), .Z(n58) );
  XNOR U219 ( .A(n67), .B(n65), .Z(o[50]) );
  NANDN U220 ( .B(n68), .A(n69), .Z(n65) );
  NANDN U221 ( .B(n70), .A(n71), .Z(n69) );
  NANDN U222 ( .B(n72), .A(n73), .Z(n71) );
  NANDN U223 ( .B(n74), .A(n75), .Z(n73) );
  NANDN U224 ( .B(n76), .A(n77), .Z(n75) );
  NANDN U225 ( .B(n78), .A(n79), .Z(n77) );
  NANDN U226 ( .B(n80), .A(n81), .Z(n79) );
  NANDN U227 ( .B(n82), .A(n83), .Z(n81) );
  NANDN U228 ( .B(n84), .A(n85), .Z(n83) );
  NANDN U229 ( .B(n86), .A(n87), .Z(n85) );
  NANDN U230 ( .B(n88), .A(n89), .Z(n87) );
  AND U231 ( .A(n90), .B(n91), .Z(n89) );
  NAND U232 ( .A(n92), .B(n93), .Z(n91) );
  NAND U233 ( .A(n94), .B(n92), .Z(n90) );
  OR U234 ( .A(\mult_26/A2[48] ), .B(\mult_26/A1[48] ), .Z(n66) );
  AND U235 ( .A(\mult_26/A2[48] ), .B(\mult_26/A1[48] ), .Z(n63) );
  XOR U236 ( .A(n95), .B(n96), .Z(o[49]) );
  ANDN U237 ( .A(n97), .B(n72), .Z(n96) );
  NANDN U238 ( .B(n74), .A(n98), .Z(n97) );
  AND U239 ( .A(\mult_26/A2[47] ), .B(\mult_26/A1[47] ), .Z(n68) );
  NOR U240 ( .A(\mult_26/A1[47] ), .B(\mult_26/A2[47] ), .Z(n70) );
  XNOR U241 ( .A(n99), .B(n98), .Z(o[48]) );
  NANDN U242 ( .B(n76), .A(n100), .Z(n98) );
  NANDN U243 ( .B(n78), .A(n101), .Z(n100) );
  AND U244 ( .A(\mult_26/A2[46] ), .B(\mult_26/A1[46] ), .Z(n72) );
  NOR U245 ( .A(\mult_26/A1[46] ), .B(\mult_26/A2[46] ), .Z(n74) );
  XNOR U246 ( .A(n102), .B(n101), .Z(o[47]) );
  NANDN U247 ( .B(n80), .A(n103), .Z(n101) );
  NANDN U248 ( .B(n82), .A(n104), .Z(n103) );
  AND U249 ( .A(\mult_26/A2[45] ), .B(\mult_26/A1[45] ), .Z(n76) );
  NOR U250 ( .A(\mult_26/A1[45] ), .B(\mult_26/A2[45] ), .Z(n78) );
  XNOR U251 ( .A(n105), .B(n104), .Z(o[46]) );
  NANDN U252 ( .B(n84), .A(n106), .Z(n104) );
  NANDN U253 ( .B(n86), .A(n107), .Z(n106) );
  NAND U254 ( .A(n108), .B(n109), .Z(n86) );
  AND U255 ( .A(n110), .B(n111), .Z(n109) );
  ANDN U256 ( .A(n112), .B(n113), .Z(n108) );
  NANDN U257 ( .B(n114), .A(n115), .Z(n84) );
  NAND U258 ( .A(n116), .B(n112), .Z(n115) );
  NANDN U259 ( .B(n117), .A(n118), .Z(n116) );
  NAND U260 ( .A(n119), .B(n111), .Z(n118) );
  NANDN U261 ( .B(n120), .A(n121), .Z(n119) );
  NAND U262 ( .A(n110), .B(n122), .Z(n121) );
  AND U263 ( .A(\mult_26/A2[44] ), .B(\mult_26/A1[44] ), .Z(n80) );
  NOR U264 ( .A(\mult_26/A1[44] ), .B(\mult_26/A2[44] ), .Z(n82) );
  XOR U265 ( .A(n123), .B(n124), .Z(o[45]) );
  ANDN U266 ( .A(n125), .B(n117), .Z(n124) );
  NAND U267 ( .A(n126), .B(n111), .Z(n125) );
  OR U268 ( .A(\mult_26/A2[43] ), .B(\mult_26/A1[43] ), .Z(n112) );
  AND U269 ( .A(\mult_26/A2[43] ), .B(\mult_26/A1[43] ), .Z(n114) );
  XNOR U270 ( .A(n127), .B(n126), .Z(o[44]) );
  NANDN U271 ( .B(n120), .A(n128), .Z(n126) );
  NAND U272 ( .A(n129), .B(n110), .Z(n128) );
  OR U273 ( .A(\mult_26/A2[42] ), .B(\mult_26/A1[42] ), .Z(n111) );
  AND U274 ( .A(\mult_26/A2[42] ), .B(\mult_26/A1[42] ), .Z(n117) );
  XNOR U275 ( .A(n130), .B(n129), .Z(o[43]) );
  NANDN U276 ( .B(n122), .A(n131), .Z(n129) );
  NANDN U277 ( .B(n113), .A(n107), .Z(n131) );
  OR U278 ( .A(\mult_26/A2[41] ), .B(\mult_26/A1[41] ), .Z(n110) );
  AND U279 ( .A(\mult_26/A2[41] ), .B(\mult_26/A1[41] ), .Z(n120) );
  XNOR U280 ( .A(n132), .B(n107), .Z(o[42]) );
  NANDN U281 ( .B(n88), .A(n133), .Z(n107) );
  NANDN U282 ( .B(n134), .A(n92), .Z(n133) );
  AND U283 ( .A(n135), .B(n136), .Z(n92) );
  AND U284 ( .A(n137), .B(n138), .Z(n136) );
  ANDN U285 ( .A(n139), .B(n140), .Z(n135) );
  NANDN U286 ( .B(n141), .A(n142), .Z(n88) );
  NAND U287 ( .A(n143), .B(n139), .Z(n142) );
  NANDN U288 ( .B(n144), .A(n145), .Z(n143) );
  NAND U289 ( .A(n146), .B(n138), .Z(n145) );
  NANDN U290 ( .B(n147), .A(n148), .Z(n146) );
  NAND U291 ( .A(n137), .B(n149), .Z(n148) );
  AND U292 ( .A(\mult_26/A2[40] ), .B(\mult_26/A1[40] ), .Z(n122) );
  NOR U293 ( .A(\mult_26/A2[40] ), .B(\mult_26/A1[40] ), .Z(n113) );
  XOR U294 ( .A(n150), .B(n151), .Z(o[41]) );
  ANDN U295 ( .A(n152), .B(n144), .Z(n151) );
  NAND U296 ( .A(n153), .B(n138), .Z(n152) );
  OR U297 ( .A(\mult_26/A2[39] ), .B(\mult_26/A1[39] ), .Z(n139) );
  AND U298 ( .A(\mult_26/A2[39] ), .B(\mult_26/A1[39] ), .Z(n141) );
  XNOR U299 ( .A(n154), .B(n153), .Z(o[40]) );
  NANDN U300 ( .B(n147), .A(n155), .Z(n153) );
  NAND U301 ( .A(n156), .B(n137), .Z(n155) );
  OR U302 ( .A(\mult_26/A2[38] ), .B(\mult_26/A1[38] ), .Z(n138) );
  AND U303 ( .A(\mult_26/A2[38] ), .B(\mult_26/A1[38] ), .Z(n144) );
  XNOR U304 ( .A(n157), .B(n156), .Z(o[39]) );
  NANDN U305 ( .B(n149), .A(n158), .Z(n156) );
  OR U306 ( .A(n134), .B(n140), .Z(n158) );
  OR U307 ( .A(\mult_26/A2[37] ), .B(\mult_26/A1[37] ), .Z(n137) );
  AND U308 ( .A(\mult_26/A2[37] ), .B(\mult_26/A1[37] ), .Z(n147) );
  XOR U309 ( .A(n159), .B(n134), .Z(o[38]) );
  NOR U310 ( .A(n94), .B(n93), .Z(n134) );
  AND U311 ( .A(n160), .B(n161), .Z(n93) );
  AND U312 ( .A(n162), .B(n163), .Z(n161) );
  AND U313 ( .A(n164), .B(n165), .Z(n163) );
  ANDN U314 ( .A(n166), .B(n167), .Z(n160) );
  NANDN U315 ( .B(n168), .A(n169), .Z(n94) );
  NAND U316 ( .A(n170), .B(n162), .Z(n169) );
  NANDN U317 ( .B(n171), .A(n172), .Z(n170) );
  NAND U318 ( .A(n173), .B(n165), .Z(n172) );
  NANDN U319 ( .B(n174), .A(n175), .Z(n173) );
  NANDN U320 ( .B(n167), .A(n176), .Z(n175) );
  AND U321 ( .A(\mult_26/A2[36] ), .B(\mult_26/A1[36] ), .Z(n149) );
  NOR U322 ( .A(\mult_26/A1[36] ), .B(\mult_26/A2[36] ), .Z(n140) );
  XOR U323 ( .A(n177), .B(n178), .Z(o[37]) );
  ANDN U324 ( .A(n179), .B(n171), .Z(n178) );
  NAND U325 ( .A(n180), .B(n165), .Z(n179) );
  OR U326 ( .A(\mult_26/A2[35] ), .B(\mult_26/A1[35] ), .Z(n162) );
  AND U327 ( .A(\mult_26/A2[35] ), .B(\mult_26/A1[35] ), .Z(n168) );
  XNOR U328 ( .A(n181), .B(n180), .Z(o[36]) );
  NANDN U329 ( .B(n174), .A(n182), .Z(n180) );
  NANDN U330 ( .B(n167), .A(n183), .Z(n182) );
  OR U331 ( .A(\mult_26/A1[34] ), .B(\mult_26/A2[34] ), .Z(n165) );
  AND U332 ( .A(\mult_26/A2[34] ), .B(\mult_26/A1[34] ), .Z(n171) );
  XNOR U333 ( .A(n184), .B(n183), .Z(o[35]) );
  NANDN U334 ( .B(n176), .A(n185), .Z(n183) );
  NAND U335 ( .A(n164), .B(n166), .Z(n185) );
  NOR U336 ( .A(\mult_26/A1[33] ), .B(\mult_26/A2[33] ), .Z(n167) );
  AND U337 ( .A(\mult_26/A2[33] ), .B(\mult_26/A1[33] ), .Z(n174) );
  XOR U338 ( .A(n166), .B(n186), .Z(o[34]) );
  AND U339 ( .A(\mult_26/A2[32] ), .B(\mult_26/A1[32] ), .Z(n176) );
  OR U340 ( .A(\mult_26/A1[32] ), .B(\mult_26/A2[32] ), .Z(n164) );
  AND U341 ( .A(\mult_26/A2[31] ), .B(\mult_26/A1[31] ), .Z(n166) );
  AND U342 ( .A(e_input[0]), .B(g_input[0]), .Z(o[0]) );
  AND U343 ( .A(e_input[9]), .B(g_input[9]), .Z(\mult_26/ab[9][9] ) );
  AND U344 ( .A(g_input[9]), .B(e_input[8]), .Z(\mult_26/ab[9][8] ) );
  AND U345 ( .A(g_input[9]), .B(e_input[7]), .Z(\mult_26/ab[9][7] ) );
  AND U346 ( .A(g_input[9]), .B(e_input[6]), .Z(\mult_26/ab[9][6] ) );
  AND U347 ( .A(g_input[9]), .B(e_input[5]), .Z(\mult_26/ab[9][5] ) );
  AND U348 ( .A(g_input[9]), .B(e_input[4]), .Z(\mult_26/ab[9][4] ) );
  AND U349 ( .A(g_input[9]), .B(e_input[3]), .Z(\mult_26/ab[9][3] ) );
  AND U350 ( .A(g_input[9]), .B(e_input[31]), .Z(\mult_26/ab[9][31] ) );
  AND U351 ( .A(g_input[9]), .B(e_input[30]), .Z(\mult_26/ab[9][30] ) );
  AND U352 ( .A(g_input[9]), .B(e_input[2]), .Z(\mult_26/ab[9][2] ) );
  AND U353 ( .A(g_input[9]), .B(e_input[29]), .Z(\mult_26/ab[9][29] ) );
  AND U354 ( .A(g_input[9]), .B(e_input[28]), .Z(\mult_26/ab[9][28] ) );
  AND U355 ( .A(g_input[9]), .B(e_input[27]), .Z(\mult_26/ab[9][27] ) );
  AND U356 ( .A(g_input[9]), .B(e_input[26]), .Z(\mult_26/ab[9][26] ) );
  AND U357 ( .A(g_input[9]), .B(e_input[25]), .Z(\mult_26/ab[9][25] ) );
  AND U358 ( .A(g_input[9]), .B(e_input[24]), .Z(\mult_26/ab[9][24] ) );
  AND U359 ( .A(g_input[9]), .B(e_input[23]), .Z(\mult_26/ab[9][23] ) );
  AND U360 ( .A(g_input[9]), .B(e_input[22]), .Z(\mult_26/ab[9][22] ) );
  AND U361 ( .A(g_input[9]), .B(e_input[21]), .Z(\mult_26/ab[9][21] ) );
  AND U362 ( .A(g_input[9]), .B(e_input[20]), .Z(\mult_26/ab[9][20] ) );
  AND U363 ( .A(g_input[9]), .B(e_input[1]), .Z(\mult_26/ab[9][1] ) );
  AND U364 ( .A(g_input[9]), .B(e_input[19]), .Z(\mult_26/ab[9][19] ) );
  AND U365 ( .A(g_input[9]), .B(e_input[18]), .Z(\mult_26/ab[9][18] ) );
  AND U366 ( .A(g_input[9]), .B(e_input[17]), .Z(\mult_26/ab[9][17] ) );
  AND U367 ( .A(g_input[9]), .B(e_input[16]), .Z(\mult_26/ab[9][16] ) );
  AND U368 ( .A(g_input[9]), .B(e_input[15]), .Z(\mult_26/ab[9][15] ) );
  AND U369 ( .A(g_input[9]), .B(e_input[14]), .Z(\mult_26/ab[9][14] ) );
  AND U370 ( .A(g_input[9]), .B(e_input[13]), .Z(\mult_26/ab[9][13] ) );
  AND U371 ( .A(g_input[9]), .B(e_input[12]), .Z(\mult_26/ab[9][12] ) );
  AND U372 ( .A(g_input[9]), .B(e_input[11]), .Z(\mult_26/ab[9][11] ) );
  AND U373 ( .A(g_input[9]), .B(e_input[10]), .Z(\mult_26/ab[9][10] ) );
  AND U374 ( .A(e_input[0]), .B(g_input[9]), .Z(\mult_26/ab[9][0] ) );
  AND U375 ( .A(e_input[9]), .B(g_input[8]), .Z(\mult_26/ab[8][9] ) );
  AND U376 ( .A(e_input[8]), .B(g_input[8]), .Z(\mult_26/ab[8][8] ) );
  AND U377 ( .A(e_input[7]), .B(g_input[8]), .Z(\mult_26/ab[8][7] ) );
  AND U378 ( .A(e_input[6]), .B(g_input[8]), .Z(\mult_26/ab[8][6] ) );
  AND U379 ( .A(e_input[5]), .B(g_input[8]), .Z(\mult_26/ab[8][5] ) );
  AND U380 ( .A(e_input[4]), .B(g_input[8]), .Z(\mult_26/ab[8][4] ) );
  AND U381 ( .A(e_input[3]), .B(g_input[8]), .Z(\mult_26/ab[8][3] ) );
  AND U382 ( .A(e_input[31]), .B(g_input[8]), .Z(\mult_26/ab[8][31] ) );
  AND U383 ( .A(e_input[30]), .B(g_input[8]), .Z(\mult_26/ab[8][30] ) );
  AND U384 ( .A(e_input[2]), .B(g_input[8]), .Z(\mult_26/ab[8][2] ) );
  AND U385 ( .A(e_input[29]), .B(g_input[8]), .Z(\mult_26/ab[8][29] ) );
  AND U386 ( .A(e_input[28]), .B(g_input[8]), .Z(\mult_26/ab[8][28] ) );
  AND U387 ( .A(e_input[27]), .B(g_input[8]), .Z(\mult_26/ab[8][27] ) );
  AND U388 ( .A(e_input[26]), .B(g_input[8]), .Z(\mult_26/ab[8][26] ) );
  AND U389 ( .A(e_input[25]), .B(g_input[8]), .Z(\mult_26/ab[8][25] ) );
  AND U390 ( .A(e_input[24]), .B(g_input[8]), .Z(\mult_26/ab[8][24] ) );
  AND U391 ( .A(e_input[23]), .B(g_input[8]), .Z(\mult_26/ab[8][23] ) );
  AND U392 ( .A(e_input[22]), .B(g_input[8]), .Z(\mult_26/ab[8][22] ) );
  AND U393 ( .A(e_input[21]), .B(g_input[8]), .Z(\mult_26/ab[8][21] ) );
  AND U394 ( .A(e_input[20]), .B(g_input[8]), .Z(\mult_26/ab[8][20] ) );
  AND U395 ( .A(e_input[1]), .B(g_input[8]), .Z(\mult_26/ab[8][1] ) );
  AND U396 ( .A(e_input[19]), .B(g_input[8]), .Z(\mult_26/ab[8][19] ) );
  AND U397 ( .A(e_input[18]), .B(g_input[8]), .Z(\mult_26/ab[8][18] ) );
  AND U398 ( .A(e_input[17]), .B(g_input[8]), .Z(\mult_26/ab[8][17] ) );
  AND U399 ( .A(e_input[16]), .B(g_input[8]), .Z(\mult_26/ab[8][16] ) );
  AND U400 ( .A(e_input[15]), .B(g_input[8]), .Z(\mult_26/ab[8][15] ) );
  AND U401 ( .A(e_input[14]), .B(g_input[8]), .Z(\mult_26/ab[8][14] ) );
  AND U402 ( .A(e_input[13]), .B(g_input[8]), .Z(\mult_26/ab[8][13] ) );
  AND U403 ( .A(e_input[12]), .B(g_input[8]), .Z(\mult_26/ab[8][12] ) );
  AND U404 ( .A(e_input[11]), .B(g_input[8]), .Z(\mult_26/ab[8][11] ) );
  AND U405 ( .A(e_input[10]), .B(g_input[8]), .Z(\mult_26/ab[8][10] ) );
  AND U406 ( .A(g_input[8]), .B(e_input[0]), .Z(\mult_26/ab[8][0] ) );
  AND U407 ( .A(e_input[9]), .B(g_input[7]), .Z(\mult_26/ab[7][9] ) );
  AND U408 ( .A(e_input[8]), .B(g_input[7]), .Z(\mult_26/ab[7][8] ) );
  AND U409 ( .A(e_input[7]), .B(g_input[7]), .Z(\mult_26/ab[7][7] ) );
  AND U410 ( .A(e_input[6]), .B(g_input[7]), .Z(\mult_26/ab[7][6] ) );
  AND U411 ( .A(e_input[5]), .B(g_input[7]), .Z(\mult_26/ab[7][5] ) );
  AND U412 ( .A(e_input[4]), .B(g_input[7]), .Z(\mult_26/ab[7][4] ) );
  AND U413 ( .A(e_input[3]), .B(g_input[7]), .Z(\mult_26/ab[7][3] ) );
  AND U414 ( .A(e_input[31]), .B(g_input[7]), .Z(\mult_26/ab[7][31] ) );
  AND U415 ( .A(e_input[30]), .B(g_input[7]), .Z(\mult_26/ab[7][30] ) );
  AND U416 ( .A(e_input[2]), .B(g_input[7]), .Z(\mult_26/ab[7][2] ) );
  AND U417 ( .A(e_input[29]), .B(g_input[7]), .Z(\mult_26/ab[7][29] ) );
  AND U418 ( .A(e_input[28]), .B(g_input[7]), .Z(\mult_26/ab[7][28] ) );
  AND U419 ( .A(e_input[27]), .B(g_input[7]), .Z(\mult_26/ab[7][27] ) );
  AND U420 ( .A(e_input[26]), .B(g_input[7]), .Z(\mult_26/ab[7][26] ) );
  AND U421 ( .A(e_input[25]), .B(g_input[7]), .Z(\mult_26/ab[7][25] ) );
  AND U422 ( .A(e_input[24]), .B(g_input[7]), .Z(\mult_26/ab[7][24] ) );
  AND U423 ( .A(e_input[23]), .B(g_input[7]), .Z(\mult_26/ab[7][23] ) );
  AND U424 ( .A(e_input[22]), .B(g_input[7]), .Z(\mult_26/ab[7][22] ) );
  AND U425 ( .A(e_input[21]), .B(g_input[7]), .Z(\mult_26/ab[7][21] ) );
  AND U426 ( .A(e_input[20]), .B(g_input[7]), .Z(\mult_26/ab[7][20] ) );
  AND U427 ( .A(e_input[1]), .B(g_input[7]), .Z(\mult_26/ab[7][1] ) );
  AND U428 ( .A(e_input[19]), .B(g_input[7]), .Z(\mult_26/ab[7][19] ) );
  AND U429 ( .A(e_input[18]), .B(g_input[7]), .Z(\mult_26/ab[7][18] ) );
  AND U430 ( .A(e_input[17]), .B(g_input[7]), .Z(\mult_26/ab[7][17] ) );
  AND U431 ( .A(e_input[16]), .B(g_input[7]), .Z(\mult_26/ab[7][16] ) );
  AND U432 ( .A(e_input[15]), .B(g_input[7]), .Z(\mult_26/ab[7][15] ) );
  AND U433 ( .A(e_input[14]), .B(g_input[7]), .Z(\mult_26/ab[7][14] ) );
  AND U434 ( .A(e_input[13]), .B(g_input[7]), .Z(\mult_26/ab[7][13] ) );
  AND U435 ( .A(e_input[12]), .B(g_input[7]), .Z(\mult_26/ab[7][12] ) );
  AND U436 ( .A(e_input[11]), .B(g_input[7]), .Z(\mult_26/ab[7][11] ) );
  AND U437 ( .A(e_input[10]), .B(g_input[7]), .Z(\mult_26/ab[7][10] ) );
  AND U438 ( .A(g_input[7]), .B(e_input[0]), .Z(\mult_26/ab[7][0] ) );
  AND U439 ( .A(e_input[9]), .B(g_input[6]), .Z(\mult_26/ab[6][9] ) );
  AND U440 ( .A(e_input[8]), .B(g_input[6]), .Z(\mult_26/ab[6][8] ) );
  AND U441 ( .A(e_input[7]), .B(g_input[6]), .Z(\mult_26/ab[6][7] ) );
  AND U442 ( .A(e_input[6]), .B(g_input[6]), .Z(\mult_26/ab[6][6] ) );
  AND U443 ( .A(e_input[5]), .B(g_input[6]), .Z(\mult_26/ab[6][5] ) );
  AND U444 ( .A(e_input[4]), .B(g_input[6]), .Z(\mult_26/ab[6][4] ) );
  AND U445 ( .A(e_input[3]), .B(g_input[6]), .Z(\mult_26/ab[6][3] ) );
  AND U446 ( .A(e_input[31]), .B(g_input[6]), .Z(\mult_26/ab[6][31] ) );
  AND U447 ( .A(e_input[30]), .B(g_input[6]), .Z(\mult_26/ab[6][30] ) );
  AND U448 ( .A(e_input[2]), .B(g_input[6]), .Z(\mult_26/ab[6][2] ) );
  AND U449 ( .A(e_input[29]), .B(g_input[6]), .Z(\mult_26/ab[6][29] ) );
  AND U450 ( .A(e_input[28]), .B(g_input[6]), .Z(\mult_26/ab[6][28] ) );
  AND U451 ( .A(e_input[27]), .B(g_input[6]), .Z(\mult_26/ab[6][27] ) );
  AND U452 ( .A(e_input[26]), .B(g_input[6]), .Z(\mult_26/ab[6][26] ) );
  AND U453 ( .A(e_input[25]), .B(g_input[6]), .Z(\mult_26/ab[6][25] ) );
  AND U454 ( .A(e_input[24]), .B(g_input[6]), .Z(\mult_26/ab[6][24] ) );
  AND U455 ( .A(e_input[23]), .B(g_input[6]), .Z(\mult_26/ab[6][23] ) );
  AND U456 ( .A(e_input[22]), .B(g_input[6]), .Z(\mult_26/ab[6][22] ) );
  AND U457 ( .A(e_input[21]), .B(g_input[6]), .Z(\mult_26/ab[6][21] ) );
  AND U458 ( .A(e_input[20]), .B(g_input[6]), .Z(\mult_26/ab[6][20] ) );
  AND U459 ( .A(e_input[1]), .B(g_input[6]), .Z(\mult_26/ab[6][1] ) );
  AND U460 ( .A(e_input[19]), .B(g_input[6]), .Z(\mult_26/ab[6][19] ) );
  AND U461 ( .A(e_input[18]), .B(g_input[6]), .Z(\mult_26/ab[6][18] ) );
  AND U462 ( .A(e_input[17]), .B(g_input[6]), .Z(\mult_26/ab[6][17] ) );
  AND U463 ( .A(e_input[16]), .B(g_input[6]), .Z(\mult_26/ab[6][16] ) );
  AND U464 ( .A(e_input[15]), .B(g_input[6]), .Z(\mult_26/ab[6][15] ) );
  AND U465 ( .A(e_input[14]), .B(g_input[6]), .Z(\mult_26/ab[6][14] ) );
  AND U466 ( .A(e_input[13]), .B(g_input[6]), .Z(\mult_26/ab[6][13] ) );
  AND U467 ( .A(e_input[12]), .B(g_input[6]), .Z(\mult_26/ab[6][12] ) );
  AND U468 ( .A(e_input[11]), .B(g_input[6]), .Z(\mult_26/ab[6][11] ) );
  AND U469 ( .A(e_input[10]), .B(g_input[6]), .Z(\mult_26/ab[6][10] ) );
  AND U470 ( .A(g_input[6]), .B(e_input[0]), .Z(\mult_26/ab[6][0] ) );
  AND U471 ( .A(e_input[9]), .B(g_input[5]), .Z(\mult_26/ab[5][9] ) );
  AND U472 ( .A(e_input[8]), .B(g_input[5]), .Z(\mult_26/ab[5][8] ) );
  AND U473 ( .A(e_input[7]), .B(g_input[5]), .Z(\mult_26/ab[5][7] ) );
  AND U474 ( .A(e_input[6]), .B(g_input[5]), .Z(\mult_26/ab[5][6] ) );
  AND U475 ( .A(e_input[5]), .B(g_input[5]), .Z(\mult_26/ab[5][5] ) );
  AND U476 ( .A(e_input[4]), .B(g_input[5]), .Z(\mult_26/ab[5][4] ) );
  AND U477 ( .A(e_input[3]), .B(g_input[5]), .Z(\mult_26/ab[5][3] ) );
  AND U478 ( .A(e_input[31]), .B(g_input[5]), .Z(\mult_26/ab[5][31] ) );
  AND U479 ( .A(e_input[30]), .B(g_input[5]), .Z(\mult_26/ab[5][30] ) );
  AND U480 ( .A(e_input[2]), .B(g_input[5]), .Z(\mult_26/ab[5][2] ) );
  AND U481 ( .A(e_input[29]), .B(g_input[5]), .Z(\mult_26/ab[5][29] ) );
  AND U482 ( .A(e_input[28]), .B(g_input[5]), .Z(\mult_26/ab[5][28] ) );
  AND U483 ( .A(e_input[27]), .B(g_input[5]), .Z(\mult_26/ab[5][27] ) );
  AND U484 ( .A(e_input[26]), .B(g_input[5]), .Z(\mult_26/ab[5][26] ) );
  AND U485 ( .A(e_input[25]), .B(g_input[5]), .Z(\mult_26/ab[5][25] ) );
  AND U486 ( .A(e_input[24]), .B(g_input[5]), .Z(\mult_26/ab[5][24] ) );
  AND U487 ( .A(e_input[23]), .B(g_input[5]), .Z(\mult_26/ab[5][23] ) );
  AND U488 ( .A(e_input[22]), .B(g_input[5]), .Z(\mult_26/ab[5][22] ) );
  AND U489 ( .A(e_input[21]), .B(g_input[5]), .Z(\mult_26/ab[5][21] ) );
  AND U490 ( .A(e_input[20]), .B(g_input[5]), .Z(\mult_26/ab[5][20] ) );
  AND U491 ( .A(e_input[1]), .B(g_input[5]), .Z(\mult_26/ab[5][1] ) );
  AND U492 ( .A(e_input[19]), .B(g_input[5]), .Z(\mult_26/ab[5][19] ) );
  AND U493 ( .A(e_input[18]), .B(g_input[5]), .Z(\mult_26/ab[5][18] ) );
  AND U494 ( .A(e_input[17]), .B(g_input[5]), .Z(\mult_26/ab[5][17] ) );
  AND U495 ( .A(e_input[16]), .B(g_input[5]), .Z(\mult_26/ab[5][16] ) );
  AND U496 ( .A(e_input[15]), .B(g_input[5]), .Z(\mult_26/ab[5][15] ) );
  AND U497 ( .A(e_input[14]), .B(g_input[5]), .Z(\mult_26/ab[5][14] ) );
  AND U498 ( .A(e_input[13]), .B(g_input[5]), .Z(\mult_26/ab[5][13] ) );
  AND U499 ( .A(e_input[12]), .B(g_input[5]), .Z(\mult_26/ab[5][12] ) );
  AND U500 ( .A(e_input[11]), .B(g_input[5]), .Z(\mult_26/ab[5][11] ) );
  AND U501 ( .A(e_input[10]), .B(g_input[5]), .Z(\mult_26/ab[5][10] ) );
  AND U502 ( .A(g_input[5]), .B(e_input[0]), .Z(\mult_26/ab[5][0] ) );
  AND U503 ( .A(e_input[9]), .B(g_input[4]), .Z(\mult_26/ab[4][9] ) );
  AND U504 ( .A(e_input[8]), .B(g_input[4]), .Z(\mult_26/ab[4][8] ) );
  AND U505 ( .A(e_input[7]), .B(g_input[4]), .Z(\mult_26/ab[4][7] ) );
  AND U506 ( .A(e_input[6]), .B(g_input[4]), .Z(\mult_26/ab[4][6] ) );
  AND U507 ( .A(e_input[5]), .B(g_input[4]), .Z(\mult_26/ab[4][5] ) );
  AND U508 ( .A(e_input[4]), .B(g_input[4]), .Z(\mult_26/ab[4][4] ) );
  AND U509 ( .A(e_input[3]), .B(g_input[4]), .Z(\mult_26/ab[4][3] ) );
  AND U510 ( .A(e_input[31]), .B(g_input[4]), .Z(\mult_26/ab[4][31] ) );
  AND U511 ( .A(e_input[30]), .B(g_input[4]), .Z(\mult_26/ab[4][30] ) );
  AND U512 ( .A(e_input[2]), .B(g_input[4]), .Z(\mult_26/ab[4][2] ) );
  AND U513 ( .A(e_input[29]), .B(g_input[4]), .Z(\mult_26/ab[4][29] ) );
  AND U514 ( .A(e_input[28]), .B(g_input[4]), .Z(\mult_26/ab[4][28] ) );
  AND U515 ( .A(e_input[27]), .B(g_input[4]), .Z(\mult_26/ab[4][27] ) );
  AND U516 ( .A(e_input[26]), .B(g_input[4]), .Z(\mult_26/ab[4][26] ) );
  AND U517 ( .A(e_input[25]), .B(g_input[4]), .Z(\mult_26/ab[4][25] ) );
  AND U518 ( .A(e_input[24]), .B(g_input[4]), .Z(\mult_26/ab[4][24] ) );
  AND U519 ( .A(e_input[23]), .B(g_input[4]), .Z(\mult_26/ab[4][23] ) );
  AND U520 ( .A(e_input[22]), .B(g_input[4]), .Z(\mult_26/ab[4][22] ) );
  AND U521 ( .A(e_input[21]), .B(g_input[4]), .Z(\mult_26/ab[4][21] ) );
  AND U522 ( .A(e_input[20]), .B(g_input[4]), .Z(\mult_26/ab[4][20] ) );
  AND U523 ( .A(e_input[1]), .B(g_input[4]), .Z(\mult_26/ab[4][1] ) );
  AND U524 ( .A(e_input[19]), .B(g_input[4]), .Z(\mult_26/ab[4][19] ) );
  AND U525 ( .A(e_input[18]), .B(g_input[4]), .Z(\mult_26/ab[4][18] ) );
  AND U526 ( .A(e_input[17]), .B(g_input[4]), .Z(\mult_26/ab[4][17] ) );
  AND U527 ( .A(e_input[16]), .B(g_input[4]), .Z(\mult_26/ab[4][16] ) );
  AND U528 ( .A(e_input[15]), .B(g_input[4]), .Z(\mult_26/ab[4][15] ) );
  AND U529 ( .A(e_input[14]), .B(g_input[4]), .Z(\mult_26/ab[4][14] ) );
  AND U530 ( .A(e_input[13]), .B(g_input[4]), .Z(\mult_26/ab[4][13] ) );
  AND U531 ( .A(e_input[12]), .B(g_input[4]), .Z(\mult_26/ab[4][12] ) );
  AND U532 ( .A(e_input[11]), .B(g_input[4]), .Z(\mult_26/ab[4][11] ) );
  AND U533 ( .A(e_input[10]), .B(g_input[4]), .Z(\mult_26/ab[4][10] ) );
  AND U534 ( .A(g_input[4]), .B(e_input[0]), .Z(\mult_26/ab[4][0] ) );
  AND U535 ( .A(e_input[9]), .B(g_input[3]), .Z(\mult_26/ab[3][9] ) );
  AND U536 ( .A(e_input[8]), .B(g_input[3]), .Z(\mult_26/ab[3][8] ) );
  AND U537 ( .A(e_input[7]), .B(g_input[3]), .Z(\mult_26/ab[3][7] ) );
  AND U538 ( .A(e_input[6]), .B(g_input[3]), .Z(\mult_26/ab[3][6] ) );
  AND U539 ( .A(e_input[5]), .B(g_input[3]), .Z(\mult_26/ab[3][5] ) );
  AND U540 ( .A(e_input[4]), .B(g_input[3]), .Z(\mult_26/ab[3][4] ) );
  AND U541 ( .A(e_input[3]), .B(g_input[3]), .Z(\mult_26/ab[3][3] ) );
  AND U542 ( .A(e_input[31]), .B(g_input[3]), .Z(\mult_26/ab[3][31] ) );
  AND U543 ( .A(e_input[30]), .B(g_input[3]), .Z(\mult_26/ab[3][30] ) );
  AND U544 ( .A(e_input[2]), .B(g_input[3]), .Z(\mult_26/ab[3][2] ) );
  AND U545 ( .A(e_input[29]), .B(g_input[3]), .Z(\mult_26/ab[3][29] ) );
  AND U546 ( .A(e_input[28]), .B(g_input[3]), .Z(\mult_26/ab[3][28] ) );
  AND U547 ( .A(e_input[27]), .B(g_input[3]), .Z(\mult_26/ab[3][27] ) );
  AND U548 ( .A(e_input[26]), .B(g_input[3]), .Z(\mult_26/ab[3][26] ) );
  AND U549 ( .A(e_input[25]), .B(g_input[3]), .Z(\mult_26/ab[3][25] ) );
  AND U550 ( .A(e_input[24]), .B(g_input[3]), .Z(\mult_26/ab[3][24] ) );
  AND U551 ( .A(e_input[23]), .B(g_input[3]), .Z(\mult_26/ab[3][23] ) );
  AND U552 ( .A(e_input[22]), .B(g_input[3]), .Z(\mult_26/ab[3][22] ) );
  AND U553 ( .A(e_input[21]), .B(g_input[3]), .Z(\mult_26/ab[3][21] ) );
  AND U554 ( .A(e_input[20]), .B(g_input[3]), .Z(\mult_26/ab[3][20] ) );
  AND U555 ( .A(e_input[1]), .B(g_input[3]), .Z(\mult_26/ab[3][1] ) );
  AND U556 ( .A(e_input[19]), .B(g_input[3]), .Z(\mult_26/ab[3][19] ) );
  AND U557 ( .A(e_input[18]), .B(g_input[3]), .Z(\mult_26/ab[3][18] ) );
  AND U558 ( .A(e_input[17]), .B(g_input[3]), .Z(\mult_26/ab[3][17] ) );
  AND U559 ( .A(e_input[16]), .B(g_input[3]), .Z(\mult_26/ab[3][16] ) );
  AND U560 ( .A(e_input[15]), .B(g_input[3]), .Z(\mult_26/ab[3][15] ) );
  AND U561 ( .A(e_input[14]), .B(g_input[3]), .Z(\mult_26/ab[3][14] ) );
  AND U562 ( .A(e_input[13]), .B(g_input[3]), .Z(\mult_26/ab[3][13] ) );
  AND U563 ( .A(e_input[12]), .B(g_input[3]), .Z(\mult_26/ab[3][12] ) );
  AND U564 ( .A(e_input[11]), .B(g_input[3]), .Z(\mult_26/ab[3][11] ) );
  AND U565 ( .A(e_input[10]), .B(g_input[3]), .Z(\mult_26/ab[3][10] ) );
  AND U566 ( .A(g_input[3]), .B(e_input[0]), .Z(\mult_26/ab[3][0] ) );
  AND U567 ( .A(e_input[9]), .B(g_input[31]), .Z(\mult_26/ab[31][9] ) );
  AND U568 ( .A(e_input[8]), .B(g_input[31]), .Z(\mult_26/ab[31][8] ) );
  AND U569 ( .A(e_input[7]), .B(g_input[31]), .Z(\mult_26/ab[31][7] ) );
  AND U570 ( .A(e_input[6]), .B(g_input[31]), .Z(\mult_26/ab[31][6] ) );
  AND U571 ( .A(e_input[5]), .B(g_input[31]), .Z(\mult_26/ab[31][5] ) );
  AND U572 ( .A(e_input[4]), .B(g_input[31]), .Z(\mult_26/ab[31][4] ) );
  AND U573 ( .A(e_input[3]), .B(g_input[31]), .Z(\mult_26/ab[31][3] ) );
  AND U574 ( .A(e_input[31]), .B(g_input[31]), .Z(\mult_26/ab[31][31] ) );
  AND U575 ( .A(e_input[30]), .B(g_input[31]), .Z(\mult_26/ab[31][30] ) );
  AND U576 ( .A(e_input[2]), .B(g_input[31]), .Z(\mult_26/ab[31][2] ) );
  AND U577 ( .A(e_input[29]), .B(g_input[31]), .Z(\mult_26/ab[31][29] ) );
  AND U578 ( .A(e_input[28]), .B(g_input[31]), .Z(\mult_26/ab[31][28] ) );
  AND U579 ( .A(e_input[27]), .B(g_input[31]), .Z(\mult_26/ab[31][27] ) );
  AND U580 ( .A(e_input[26]), .B(g_input[31]), .Z(\mult_26/ab[31][26] ) );
  AND U581 ( .A(e_input[25]), .B(g_input[31]), .Z(\mult_26/ab[31][25] ) );
  AND U582 ( .A(e_input[24]), .B(g_input[31]), .Z(\mult_26/ab[31][24] ) );
  AND U583 ( .A(e_input[23]), .B(g_input[31]), .Z(\mult_26/ab[31][23] ) );
  AND U584 ( .A(e_input[22]), .B(g_input[31]), .Z(\mult_26/ab[31][22] ) );
  AND U585 ( .A(e_input[21]), .B(g_input[31]), .Z(\mult_26/ab[31][21] ) );
  AND U586 ( .A(e_input[20]), .B(g_input[31]), .Z(\mult_26/ab[31][20] ) );
  AND U587 ( .A(e_input[1]), .B(g_input[31]), .Z(\mult_26/ab[31][1] ) );
  AND U588 ( .A(e_input[19]), .B(g_input[31]), .Z(\mult_26/ab[31][19] ) );
  AND U589 ( .A(e_input[18]), .B(g_input[31]), .Z(\mult_26/ab[31][18] ) );
  AND U590 ( .A(e_input[17]), .B(g_input[31]), .Z(\mult_26/ab[31][17] ) );
  AND U591 ( .A(e_input[16]), .B(g_input[31]), .Z(\mult_26/ab[31][16] ) );
  AND U592 ( .A(e_input[15]), .B(g_input[31]), .Z(\mult_26/ab[31][15] ) );
  AND U593 ( .A(e_input[14]), .B(g_input[31]), .Z(\mult_26/ab[31][14] ) );
  AND U594 ( .A(e_input[13]), .B(g_input[31]), .Z(\mult_26/ab[31][13] ) );
  AND U595 ( .A(e_input[12]), .B(g_input[31]), .Z(\mult_26/ab[31][12] ) );
  AND U596 ( .A(e_input[11]), .B(g_input[31]), .Z(\mult_26/ab[31][11] ) );
  AND U597 ( .A(e_input[10]), .B(g_input[31]), .Z(\mult_26/ab[31][10] ) );
  AND U598 ( .A(g_input[31]), .B(e_input[0]), .Z(\mult_26/ab[31][0] ) );
  AND U599 ( .A(e_input[9]), .B(g_input[30]), .Z(\mult_26/ab[30][9] ) );
  AND U600 ( .A(e_input[8]), .B(g_input[30]), .Z(\mult_26/ab[30][8] ) );
  AND U601 ( .A(e_input[7]), .B(g_input[30]), .Z(\mult_26/ab[30][7] ) );
  AND U602 ( .A(e_input[6]), .B(g_input[30]), .Z(\mult_26/ab[30][6] ) );
  AND U603 ( .A(e_input[5]), .B(g_input[30]), .Z(\mult_26/ab[30][5] ) );
  AND U604 ( .A(e_input[4]), .B(g_input[30]), .Z(\mult_26/ab[30][4] ) );
  AND U605 ( .A(e_input[3]), .B(g_input[30]), .Z(\mult_26/ab[30][3] ) );
  AND U606 ( .A(e_input[31]), .B(g_input[30]), .Z(\mult_26/ab[30][31] ) );
  AND U607 ( .A(e_input[30]), .B(g_input[30]), .Z(\mult_26/ab[30][30] ) );
  AND U608 ( .A(e_input[2]), .B(g_input[30]), .Z(\mult_26/ab[30][2] ) );
  AND U609 ( .A(e_input[29]), .B(g_input[30]), .Z(\mult_26/ab[30][29] ) );
  AND U610 ( .A(e_input[28]), .B(g_input[30]), .Z(\mult_26/ab[30][28] ) );
  AND U611 ( .A(e_input[27]), .B(g_input[30]), .Z(\mult_26/ab[30][27] ) );
  AND U612 ( .A(e_input[26]), .B(g_input[30]), .Z(\mult_26/ab[30][26] ) );
  AND U613 ( .A(e_input[25]), .B(g_input[30]), .Z(\mult_26/ab[30][25] ) );
  AND U614 ( .A(e_input[24]), .B(g_input[30]), .Z(\mult_26/ab[30][24] ) );
  AND U615 ( .A(e_input[23]), .B(g_input[30]), .Z(\mult_26/ab[30][23] ) );
  AND U616 ( .A(e_input[22]), .B(g_input[30]), .Z(\mult_26/ab[30][22] ) );
  AND U617 ( .A(e_input[21]), .B(g_input[30]), .Z(\mult_26/ab[30][21] ) );
  AND U618 ( .A(e_input[20]), .B(g_input[30]), .Z(\mult_26/ab[30][20] ) );
  AND U619 ( .A(e_input[1]), .B(g_input[30]), .Z(\mult_26/ab[30][1] ) );
  AND U620 ( .A(e_input[19]), .B(g_input[30]), .Z(\mult_26/ab[30][19] ) );
  AND U621 ( .A(e_input[18]), .B(g_input[30]), .Z(\mult_26/ab[30][18] ) );
  AND U622 ( .A(e_input[17]), .B(g_input[30]), .Z(\mult_26/ab[30][17] ) );
  AND U623 ( .A(e_input[16]), .B(g_input[30]), .Z(\mult_26/ab[30][16] ) );
  AND U624 ( .A(e_input[15]), .B(g_input[30]), .Z(\mult_26/ab[30][15] ) );
  AND U625 ( .A(e_input[14]), .B(g_input[30]), .Z(\mult_26/ab[30][14] ) );
  AND U626 ( .A(e_input[13]), .B(g_input[30]), .Z(\mult_26/ab[30][13] ) );
  AND U627 ( .A(e_input[12]), .B(g_input[30]), .Z(\mult_26/ab[30][12] ) );
  AND U628 ( .A(e_input[11]), .B(g_input[30]), .Z(\mult_26/ab[30][11] ) );
  AND U629 ( .A(e_input[10]), .B(g_input[30]), .Z(\mult_26/ab[30][10] ) );
  AND U630 ( .A(g_input[30]), .B(e_input[0]), .Z(\mult_26/ab[30][0] ) );
  AND U631 ( .A(e_input[9]), .B(g_input[2]), .Z(\mult_26/ab[2][9] ) );
  AND U632 ( .A(e_input[8]), .B(g_input[2]), .Z(\mult_26/ab[2][8] ) );
  AND U633 ( .A(e_input[7]), .B(g_input[2]), .Z(\mult_26/ab[2][7] ) );
  AND U634 ( .A(e_input[6]), .B(g_input[2]), .Z(\mult_26/ab[2][6] ) );
  AND U635 ( .A(e_input[5]), .B(g_input[2]), .Z(\mult_26/ab[2][5] ) );
  AND U636 ( .A(e_input[4]), .B(g_input[2]), .Z(\mult_26/ab[2][4] ) );
  AND U637 ( .A(e_input[3]), .B(g_input[2]), .Z(\mult_26/ab[2][3] ) );
  AND U638 ( .A(e_input[31]), .B(g_input[2]), .Z(\mult_26/ab[2][31] ) );
  AND U639 ( .A(e_input[30]), .B(g_input[2]), .Z(\mult_26/ab[2][30] ) );
  AND U640 ( .A(e_input[2]), .B(g_input[2]), .Z(\mult_26/ab[2][2] ) );
  AND U641 ( .A(e_input[29]), .B(g_input[2]), .Z(\mult_26/ab[2][29] ) );
  AND U642 ( .A(e_input[28]), .B(g_input[2]), .Z(\mult_26/ab[2][28] ) );
  AND U643 ( .A(e_input[27]), .B(g_input[2]), .Z(\mult_26/ab[2][27] ) );
  AND U644 ( .A(e_input[26]), .B(g_input[2]), .Z(\mult_26/ab[2][26] ) );
  AND U645 ( .A(e_input[25]), .B(g_input[2]), .Z(\mult_26/ab[2][25] ) );
  AND U646 ( .A(e_input[24]), .B(g_input[2]), .Z(\mult_26/ab[2][24] ) );
  AND U647 ( .A(e_input[23]), .B(g_input[2]), .Z(\mult_26/ab[2][23] ) );
  AND U648 ( .A(e_input[22]), .B(g_input[2]), .Z(\mult_26/ab[2][22] ) );
  AND U649 ( .A(e_input[21]), .B(g_input[2]), .Z(\mult_26/ab[2][21] ) );
  AND U650 ( .A(e_input[20]), .B(g_input[2]), .Z(\mult_26/ab[2][20] ) );
  AND U651 ( .A(e_input[1]), .B(g_input[2]), .Z(\mult_26/ab[2][1] ) );
  AND U652 ( .A(e_input[19]), .B(g_input[2]), .Z(\mult_26/ab[2][19] ) );
  AND U653 ( .A(e_input[18]), .B(g_input[2]), .Z(\mult_26/ab[2][18] ) );
  AND U654 ( .A(e_input[17]), .B(g_input[2]), .Z(\mult_26/ab[2][17] ) );
  AND U655 ( .A(e_input[16]), .B(g_input[2]), .Z(\mult_26/ab[2][16] ) );
  AND U656 ( .A(e_input[15]), .B(g_input[2]), .Z(\mult_26/ab[2][15] ) );
  AND U657 ( .A(e_input[14]), .B(g_input[2]), .Z(\mult_26/ab[2][14] ) );
  AND U658 ( .A(e_input[13]), .B(g_input[2]), .Z(\mult_26/ab[2][13] ) );
  AND U659 ( .A(e_input[12]), .B(g_input[2]), .Z(\mult_26/ab[2][12] ) );
  AND U660 ( .A(e_input[11]), .B(g_input[2]), .Z(\mult_26/ab[2][11] ) );
  AND U661 ( .A(e_input[10]), .B(g_input[2]), .Z(\mult_26/ab[2][10] ) );
  AND U662 ( .A(g_input[2]), .B(e_input[0]), .Z(\mult_26/ab[2][0] ) );
  AND U663 ( .A(e_input[9]), .B(g_input[29]), .Z(\mult_26/ab[29][9] ) );
  AND U664 ( .A(e_input[8]), .B(g_input[29]), .Z(\mult_26/ab[29][8] ) );
  AND U665 ( .A(e_input[7]), .B(g_input[29]), .Z(\mult_26/ab[29][7] ) );
  AND U666 ( .A(e_input[6]), .B(g_input[29]), .Z(\mult_26/ab[29][6] ) );
  AND U667 ( .A(e_input[5]), .B(g_input[29]), .Z(\mult_26/ab[29][5] ) );
  AND U668 ( .A(e_input[4]), .B(g_input[29]), .Z(\mult_26/ab[29][4] ) );
  AND U669 ( .A(e_input[3]), .B(g_input[29]), .Z(\mult_26/ab[29][3] ) );
  AND U670 ( .A(e_input[31]), .B(g_input[29]), .Z(\mult_26/ab[29][31] ) );
  AND U671 ( .A(e_input[30]), .B(g_input[29]), .Z(\mult_26/ab[29][30] ) );
  AND U672 ( .A(e_input[2]), .B(g_input[29]), .Z(\mult_26/ab[29][2] ) );
  AND U673 ( .A(e_input[29]), .B(g_input[29]), .Z(\mult_26/ab[29][29] ) );
  AND U674 ( .A(e_input[28]), .B(g_input[29]), .Z(\mult_26/ab[29][28] ) );
  AND U675 ( .A(e_input[27]), .B(g_input[29]), .Z(\mult_26/ab[29][27] ) );
  AND U676 ( .A(e_input[26]), .B(g_input[29]), .Z(\mult_26/ab[29][26] ) );
  AND U677 ( .A(e_input[25]), .B(g_input[29]), .Z(\mult_26/ab[29][25] ) );
  AND U678 ( .A(e_input[24]), .B(g_input[29]), .Z(\mult_26/ab[29][24] ) );
  AND U679 ( .A(e_input[23]), .B(g_input[29]), .Z(\mult_26/ab[29][23] ) );
  AND U680 ( .A(e_input[22]), .B(g_input[29]), .Z(\mult_26/ab[29][22] ) );
  AND U681 ( .A(e_input[21]), .B(g_input[29]), .Z(\mult_26/ab[29][21] ) );
  AND U682 ( .A(e_input[20]), .B(g_input[29]), .Z(\mult_26/ab[29][20] ) );
  AND U683 ( .A(e_input[1]), .B(g_input[29]), .Z(\mult_26/ab[29][1] ) );
  AND U684 ( .A(e_input[19]), .B(g_input[29]), .Z(\mult_26/ab[29][19] ) );
  AND U685 ( .A(e_input[18]), .B(g_input[29]), .Z(\mult_26/ab[29][18] ) );
  AND U686 ( .A(e_input[17]), .B(g_input[29]), .Z(\mult_26/ab[29][17] ) );
  AND U687 ( .A(e_input[16]), .B(g_input[29]), .Z(\mult_26/ab[29][16] ) );
  AND U688 ( .A(e_input[15]), .B(g_input[29]), .Z(\mult_26/ab[29][15] ) );
  AND U689 ( .A(e_input[14]), .B(g_input[29]), .Z(\mult_26/ab[29][14] ) );
  AND U690 ( .A(e_input[13]), .B(g_input[29]), .Z(\mult_26/ab[29][13] ) );
  AND U691 ( .A(e_input[12]), .B(g_input[29]), .Z(\mult_26/ab[29][12] ) );
  AND U692 ( .A(e_input[11]), .B(g_input[29]), .Z(\mult_26/ab[29][11] ) );
  AND U693 ( .A(e_input[10]), .B(g_input[29]), .Z(\mult_26/ab[29][10] ) );
  AND U694 ( .A(g_input[29]), .B(e_input[0]), .Z(\mult_26/ab[29][0] ) );
  AND U695 ( .A(e_input[9]), .B(g_input[28]), .Z(\mult_26/ab[28][9] ) );
  AND U696 ( .A(e_input[8]), .B(g_input[28]), .Z(\mult_26/ab[28][8] ) );
  AND U697 ( .A(e_input[7]), .B(g_input[28]), .Z(\mult_26/ab[28][7] ) );
  AND U698 ( .A(e_input[6]), .B(g_input[28]), .Z(\mult_26/ab[28][6] ) );
  AND U699 ( .A(e_input[5]), .B(g_input[28]), .Z(\mult_26/ab[28][5] ) );
  AND U700 ( .A(e_input[4]), .B(g_input[28]), .Z(\mult_26/ab[28][4] ) );
  AND U701 ( .A(e_input[3]), .B(g_input[28]), .Z(\mult_26/ab[28][3] ) );
  AND U702 ( .A(e_input[31]), .B(g_input[28]), .Z(\mult_26/ab[28][31] ) );
  AND U703 ( .A(e_input[30]), .B(g_input[28]), .Z(\mult_26/ab[28][30] ) );
  AND U704 ( .A(e_input[2]), .B(g_input[28]), .Z(\mult_26/ab[28][2] ) );
  AND U705 ( .A(e_input[29]), .B(g_input[28]), .Z(\mult_26/ab[28][29] ) );
  AND U706 ( .A(e_input[28]), .B(g_input[28]), .Z(\mult_26/ab[28][28] ) );
  AND U707 ( .A(e_input[27]), .B(g_input[28]), .Z(\mult_26/ab[28][27] ) );
  AND U708 ( .A(e_input[26]), .B(g_input[28]), .Z(\mult_26/ab[28][26] ) );
  AND U709 ( .A(e_input[25]), .B(g_input[28]), .Z(\mult_26/ab[28][25] ) );
  AND U710 ( .A(e_input[24]), .B(g_input[28]), .Z(\mult_26/ab[28][24] ) );
  AND U711 ( .A(e_input[23]), .B(g_input[28]), .Z(\mult_26/ab[28][23] ) );
  AND U712 ( .A(e_input[22]), .B(g_input[28]), .Z(\mult_26/ab[28][22] ) );
  AND U713 ( .A(e_input[21]), .B(g_input[28]), .Z(\mult_26/ab[28][21] ) );
  AND U714 ( .A(e_input[20]), .B(g_input[28]), .Z(\mult_26/ab[28][20] ) );
  AND U715 ( .A(e_input[1]), .B(g_input[28]), .Z(\mult_26/ab[28][1] ) );
  AND U716 ( .A(e_input[19]), .B(g_input[28]), .Z(\mult_26/ab[28][19] ) );
  AND U717 ( .A(e_input[18]), .B(g_input[28]), .Z(\mult_26/ab[28][18] ) );
  AND U718 ( .A(e_input[17]), .B(g_input[28]), .Z(\mult_26/ab[28][17] ) );
  AND U719 ( .A(e_input[16]), .B(g_input[28]), .Z(\mult_26/ab[28][16] ) );
  AND U720 ( .A(e_input[15]), .B(g_input[28]), .Z(\mult_26/ab[28][15] ) );
  AND U721 ( .A(e_input[14]), .B(g_input[28]), .Z(\mult_26/ab[28][14] ) );
  AND U722 ( .A(e_input[13]), .B(g_input[28]), .Z(\mult_26/ab[28][13] ) );
  AND U723 ( .A(e_input[12]), .B(g_input[28]), .Z(\mult_26/ab[28][12] ) );
  AND U724 ( .A(e_input[11]), .B(g_input[28]), .Z(\mult_26/ab[28][11] ) );
  AND U725 ( .A(e_input[10]), .B(g_input[28]), .Z(\mult_26/ab[28][10] ) );
  AND U726 ( .A(g_input[28]), .B(e_input[0]), .Z(\mult_26/ab[28][0] ) );
  AND U727 ( .A(e_input[9]), .B(g_input[27]), .Z(\mult_26/ab[27][9] ) );
  AND U728 ( .A(e_input[8]), .B(g_input[27]), .Z(\mult_26/ab[27][8] ) );
  AND U729 ( .A(e_input[7]), .B(g_input[27]), .Z(\mult_26/ab[27][7] ) );
  AND U730 ( .A(e_input[6]), .B(g_input[27]), .Z(\mult_26/ab[27][6] ) );
  AND U731 ( .A(e_input[5]), .B(g_input[27]), .Z(\mult_26/ab[27][5] ) );
  AND U732 ( .A(e_input[4]), .B(g_input[27]), .Z(\mult_26/ab[27][4] ) );
  AND U733 ( .A(e_input[3]), .B(g_input[27]), .Z(\mult_26/ab[27][3] ) );
  AND U734 ( .A(e_input[31]), .B(g_input[27]), .Z(\mult_26/ab[27][31] ) );
  AND U735 ( .A(e_input[30]), .B(g_input[27]), .Z(\mult_26/ab[27][30] ) );
  AND U736 ( .A(e_input[2]), .B(g_input[27]), .Z(\mult_26/ab[27][2] ) );
  AND U737 ( .A(e_input[29]), .B(g_input[27]), .Z(\mult_26/ab[27][29] ) );
  AND U738 ( .A(e_input[28]), .B(g_input[27]), .Z(\mult_26/ab[27][28] ) );
  AND U739 ( .A(e_input[27]), .B(g_input[27]), .Z(\mult_26/ab[27][27] ) );
  AND U740 ( .A(e_input[26]), .B(g_input[27]), .Z(\mult_26/ab[27][26] ) );
  AND U741 ( .A(e_input[25]), .B(g_input[27]), .Z(\mult_26/ab[27][25] ) );
  AND U742 ( .A(e_input[24]), .B(g_input[27]), .Z(\mult_26/ab[27][24] ) );
  AND U743 ( .A(e_input[23]), .B(g_input[27]), .Z(\mult_26/ab[27][23] ) );
  AND U744 ( .A(e_input[22]), .B(g_input[27]), .Z(\mult_26/ab[27][22] ) );
  AND U745 ( .A(e_input[21]), .B(g_input[27]), .Z(\mult_26/ab[27][21] ) );
  AND U746 ( .A(e_input[20]), .B(g_input[27]), .Z(\mult_26/ab[27][20] ) );
  AND U747 ( .A(e_input[1]), .B(g_input[27]), .Z(\mult_26/ab[27][1] ) );
  AND U748 ( .A(e_input[19]), .B(g_input[27]), .Z(\mult_26/ab[27][19] ) );
  AND U749 ( .A(e_input[18]), .B(g_input[27]), .Z(\mult_26/ab[27][18] ) );
  AND U750 ( .A(e_input[17]), .B(g_input[27]), .Z(\mult_26/ab[27][17] ) );
  AND U751 ( .A(e_input[16]), .B(g_input[27]), .Z(\mult_26/ab[27][16] ) );
  AND U752 ( .A(e_input[15]), .B(g_input[27]), .Z(\mult_26/ab[27][15] ) );
  AND U753 ( .A(e_input[14]), .B(g_input[27]), .Z(\mult_26/ab[27][14] ) );
  AND U754 ( .A(e_input[13]), .B(g_input[27]), .Z(\mult_26/ab[27][13] ) );
  AND U755 ( .A(e_input[12]), .B(g_input[27]), .Z(\mult_26/ab[27][12] ) );
  AND U756 ( .A(e_input[11]), .B(g_input[27]), .Z(\mult_26/ab[27][11] ) );
  AND U757 ( .A(e_input[10]), .B(g_input[27]), .Z(\mult_26/ab[27][10] ) );
  AND U758 ( .A(g_input[27]), .B(e_input[0]), .Z(\mult_26/ab[27][0] ) );
  AND U759 ( .A(e_input[9]), .B(g_input[26]), .Z(\mult_26/ab[26][9] ) );
  AND U760 ( .A(e_input[8]), .B(g_input[26]), .Z(\mult_26/ab[26][8] ) );
  AND U761 ( .A(e_input[7]), .B(g_input[26]), .Z(\mult_26/ab[26][7] ) );
  AND U762 ( .A(e_input[6]), .B(g_input[26]), .Z(\mult_26/ab[26][6] ) );
  AND U763 ( .A(e_input[5]), .B(g_input[26]), .Z(\mult_26/ab[26][5] ) );
  AND U764 ( .A(e_input[4]), .B(g_input[26]), .Z(\mult_26/ab[26][4] ) );
  AND U765 ( .A(e_input[3]), .B(g_input[26]), .Z(\mult_26/ab[26][3] ) );
  AND U766 ( .A(e_input[31]), .B(g_input[26]), .Z(\mult_26/ab[26][31] ) );
  AND U767 ( .A(e_input[30]), .B(g_input[26]), .Z(\mult_26/ab[26][30] ) );
  AND U768 ( .A(e_input[2]), .B(g_input[26]), .Z(\mult_26/ab[26][2] ) );
  AND U769 ( .A(e_input[29]), .B(g_input[26]), .Z(\mult_26/ab[26][29] ) );
  AND U770 ( .A(e_input[28]), .B(g_input[26]), .Z(\mult_26/ab[26][28] ) );
  AND U771 ( .A(e_input[27]), .B(g_input[26]), .Z(\mult_26/ab[26][27] ) );
  AND U772 ( .A(e_input[26]), .B(g_input[26]), .Z(\mult_26/ab[26][26] ) );
  AND U773 ( .A(e_input[25]), .B(g_input[26]), .Z(\mult_26/ab[26][25] ) );
  AND U774 ( .A(e_input[24]), .B(g_input[26]), .Z(\mult_26/ab[26][24] ) );
  AND U775 ( .A(e_input[23]), .B(g_input[26]), .Z(\mult_26/ab[26][23] ) );
  AND U776 ( .A(e_input[22]), .B(g_input[26]), .Z(\mult_26/ab[26][22] ) );
  AND U777 ( .A(e_input[21]), .B(g_input[26]), .Z(\mult_26/ab[26][21] ) );
  AND U778 ( .A(e_input[20]), .B(g_input[26]), .Z(\mult_26/ab[26][20] ) );
  AND U779 ( .A(e_input[1]), .B(g_input[26]), .Z(\mult_26/ab[26][1] ) );
  AND U780 ( .A(e_input[19]), .B(g_input[26]), .Z(\mult_26/ab[26][19] ) );
  AND U781 ( .A(e_input[18]), .B(g_input[26]), .Z(\mult_26/ab[26][18] ) );
  AND U782 ( .A(e_input[17]), .B(g_input[26]), .Z(\mult_26/ab[26][17] ) );
  AND U783 ( .A(e_input[16]), .B(g_input[26]), .Z(\mult_26/ab[26][16] ) );
  AND U784 ( .A(e_input[15]), .B(g_input[26]), .Z(\mult_26/ab[26][15] ) );
  AND U785 ( .A(e_input[14]), .B(g_input[26]), .Z(\mult_26/ab[26][14] ) );
  AND U786 ( .A(e_input[13]), .B(g_input[26]), .Z(\mult_26/ab[26][13] ) );
  AND U787 ( .A(e_input[12]), .B(g_input[26]), .Z(\mult_26/ab[26][12] ) );
  AND U788 ( .A(e_input[11]), .B(g_input[26]), .Z(\mult_26/ab[26][11] ) );
  AND U789 ( .A(e_input[10]), .B(g_input[26]), .Z(\mult_26/ab[26][10] ) );
  AND U790 ( .A(g_input[26]), .B(e_input[0]), .Z(\mult_26/ab[26][0] ) );
  AND U791 ( .A(e_input[9]), .B(g_input[25]), .Z(\mult_26/ab[25][9] ) );
  AND U792 ( .A(e_input[8]), .B(g_input[25]), .Z(\mult_26/ab[25][8] ) );
  AND U793 ( .A(e_input[7]), .B(g_input[25]), .Z(\mult_26/ab[25][7] ) );
  AND U794 ( .A(e_input[6]), .B(g_input[25]), .Z(\mult_26/ab[25][6] ) );
  AND U795 ( .A(e_input[5]), .B(g_input[25]), .Z(\mult_26/ab[25][5] ) );
  AND U796 ( .A(e_input[4]), .B(g_input[25]), .Z(\mult_26/ab[25][4] ) );
  AND U797 ( .A(e_input[3]), .B(g_input[25]), .Z(\mult_26/ab[25][3] ) );
  AND U798 ( .A(e_input[31]), .B(g_input[25]), .Z(\mult_26/ab[25][31] ) );
  AND U799 ( .A(e_input[30]), .B(g_input[25]), .Z(\mult_26/ab[25][30] ) );
  AND U800 ( .A(e_input[2]), .B(g_input[25]), .Z(\mult_26/ab[25][2] ) );
  AND U801 ( .A(e_input[29]), .B(g_input[25]), .Z(\mult_26/ab[25][29] ) );
  AND U802 ( .A(e_input[28]), .B(g_input[25]), .Z(\mult_26/ab[25][28] ) );
  AND U803 ( .A(e_input[27]), .B(g_input[25]), .Z(\mult_26/ab[25][27] ) );
  AND U804 ( .A(e_input[26]), .B(g_input[25]), .Z(\mult_26/ab[25][26] ) );
  AND U805 ( .A(e_input[25]), .B(g_input[25]), .Z(\mult_26/ab[25][25] ) );
  AND U806 ( .A(e_input[24]), .B(g_input[25]), .Z(\mult_26/ab[25][24] ) );
  AND U807 ( .A(e_input[23]), .B(g_input[25]), .Z(\mult_26/ab[25][23] ) );
  AND U808 ( .A(e_input[22]), .B(g_input[25]), .Z(\mult_26/ab[25][22] ) );
  AND U809 ( .A(e_input[21]), .B(g_input[25]), .Z(\mult_26/ab[25][21] ) );
  AND U810 ( .A(e_input[20]), .B(g_input[25]), .Z(\mult_26/ab[25][20] ) );
  AND U811 ( .A(e_input[1]), .B(g_input[25]), .Z(\mult_26/ab[25][1] ) );
  AND U812 ( .A(e_input[19]), .B(g_input[25]), .Z(\mult_26/ab[25][19] ) );
  AND U813 ( .A(e_input[18]), .B(g_input[25]), .Z(\mult_26/ab[25][18] ) );
  AND U814 ( .A(e_input[17]), .B(g_input[25]), .Z(\mult_26/ab[25][17] ) );
  AND U815 ( .A(e_input[16]), .B(g_input[25]), .Z(\mult_26/ab[25][16] ) );
  AND U816 ( .A(e_input[15]), .B(g_input[25]), .Z(\mult_26/ab[25][15] ) );
  AND U817 ( .A(e_input[14]), .B(g_input[25]), .Z(\mult_26/ab[25][14] ) );
  AND U818 ( .A(e_input[13]), .B(g_input[25]), .Z(\mult_26/ab[25][13] ) );
  AND U819 ( .A(e_input[12]), .B(g_input[25]), .Z(\mult_26/ab[25][12] ) );
  AND U820 ( .A(e_input[11]), .B(g_input[25]), .Z(\mult_26/ab[25][11] ) );
  AND U821 ( .A(e_input[10]), .B(g_input[25]), .Z(\mult_26/ab[25][10] ) );
  AND U822 ( .A(g_input[25]), .B(e_input[0]), .Z(\mult_26/ab[25][0] ) );
  AND U823 ( .A(e_input[9]), .B(g_input[24]), .Z(\mult_26/ab[24][9] ) );
  AND U824 ( .A(e_input[8]), .B(g_input[24]), .Z(\mult_26/ab[24][8] ) );
  AND U825 ( .A(e_input[7]), .B(g_input[24]), .Z(\mult_26/ab[24][7] ) );
  AND U826 ( .A(e_input[6]), .B(g_input[24]), .Z(\mult_26/ab[24][6] ) );
  AND U827 ( .A(e_input[5]), .B(g_input[24]), .Z(\mult_26/ab[24][5] ) );
  AND U828 ( .A(e_input[4]), .B(g_input[24]), .Z(\mult_26/ab[24][4] ) );
  AND U829 ( .A(e_input[3]), .B(g_input[24]), .Z(\mult_26/ab[24][3] ) );
  AND U830 ( .A(e_input[31]), .B(g_input[24]), .Z(\mult_26/ab[24][31] ) );
  AND U831 ( .A(e_input[30]), .B(g_input[24]), .Z(\mult_26/ab[24][30] ) );
  AND U832 ( .A(e_input[2]), .B(g_input[24]), .Z(\mult_26/ab[24][2] ) );
  AND U833 ( .A(e_input[29]), .B(g_input[24]), .Z(\mult_26/ab[24][29] ) );
  AND U834 ( .A(e_input[28]), .B(g_input[24]), .Z(\mult_26/ab[24][28] ) );
  AND U835 ( .A(e_input[27]), .B(g_input[24]), .Z(\mult_26/ab[24][27] ) );
  AND U836 ( .A(e_input[26]), .B(g_input[24]), .Z(\mult_26/ab[24][26] ) );
  AND U837 ( .A(e_input[25]), .B(g_input[24]), .Z(\mult_26/ab[24][25] ) );
  AND U838 ( .A(e_input[24]), .B(g_input[24]), .Z(\mult_26/ab[24][24] ) );
  AND U839 ( .A(e_input[23]), .B(g_input[24]), .Z(\mult_26/ab[24][23] ) );
  AND U840 ( .A(e_input[22]), .B(g_input[24]), .Z(\mult_26/ab[24][22] ) );
  AND U841 ( .A(e_input[21]), .B(g_input[24]), .Z(\mult_26/ab[24][21] ) );
  AND U842 ( .A(e_input[20]), .B(g_input[24]), .Z(\mult_26/ab[24][20] ) );
  AND U843 ( .A(e_input[1]), .B(g_input[24]), .Z(\mult_26/ab[24][1] ) );
  AND U844 ( .A(e_input[19]), .B(g_input[24]), .Z(\mult_26/ab[24][19] ) );
  AND U845 ( .A(e_input[18]), .B(g_input[24]), .Z(\mult_26/ab[24][18] ) );
  AND U846 ( .A(e_input[17]), .B(g_input[24]), .Z(\mult_26/ab[24][17] ) );
  AND U847 ( .A(e_input[16]), .B(g_input[24]), .Z(\mult_26/ab[24][16] ) );
  AND U848 ( .A(e_input[15]), .B(g_input[24]), .Z(\mult_26/ab[24][15] ) );
  AND U849 ( .A(e_input[14]), .B(g_input[24]), .Z(\mult_26/ab[24][14] ) );
  AND U850 ( .A(e_input[13]), .B(g_input[24]), .Z(\mult_26/ab[24][13] ) );
  AND U851 ( .A(e_input[12]), .B(g_input[24]), .Z(\mult_26/ab[24][12] ) );
  AND U852 ( .A(e_input[11]), .B(g_input[24]), .Z(\mult_26/ab[24][11] ) );
  AND U853 ( .A(e_input[10]), .B(g_input[24]), .Z(\mult_26/ab[24][10] ) );
  AND U854 ( .A(g_input[24]), .B(e_input[0]), .Z(\mult_26/ab[24][0] ) );
  AND U855 ( .A(e_input[9]), .B(g_input[23]), .Z(\mult_26/ab[23][9] ) );
  AND U856 ( .A(e_input[8]), .B(g_input[23]), .Z(\mult_26/ab[23][8] ) );
  AND U857 ( .A(e_input[7]), .B(g_input[23]), .Z(\mult_26/ab[23][7] ) );
  AND U858 ( .A(e_input[6]), .B(g_input[23]), .Z(\mult_26/ab[23][6] ) );
  AND U859 ( .A(e_input[5]), .B(g_input[23]), .Z(\mult_26/ab[23][5] ) );
  AND U860 ( .A(e_input[4]), .B(g_input[23]), .Z(\mult_26/ab[23][4] ) );
  AND U861 ( .A(e_input[3]), .B(g_input[23]), .Z(\mult_26/ab[23][3] ) );
  AND U862 ( .A(e_input[31]), .B(g_input[23]), .Z(\mult_26/ab[23][31] ) );
  AND U863 ( .A(e_input[30]), .B(g_input[23]), .Z(\mult_26/ab[23][30] ) );
  AND U864 ( .A(e_input[2]), .B(g_input[23]), .Z(\mult_26/ab[23][2] ) );
  AND U865 ( .A(e_input[29]), .B(g_input[23]), .Z(\mult_26/ab[23][29] ) );
  AND U866 ( .A(e_input[28]), .B(g_input[23]), .Z(\mult_26/ab[23][28] ) );
  AND U867 ( .A(e_input[27]), .B(g_input[23]), .Z(\mult_26/ab[23][27] ) );
  AND U868 ( .A(e_input[26]), .B(g_input[23]), .Z(\mult_26/ab[23][26] ) );
  AND U869 ( .A(e_input[25]), .B(g_input[23]), .Z(\mult_26/ab[23][25] ) );
  AND U870 ( .A(e_input[24]), .B(g_input[23]), .Z(\mult_26/ab[23][24] ) );
  AND U871 ( .A(e_input[23]), .B(g_input[23]), .Z(\mult_26/ab[23][23] ) );
  AND U872 ( .A(e_input[22]), .B(g_input[23]), .Z(\mult_26/ab[23][22] ) );
  AND U873 ( .A(e_input[21]), .B(g_input[23]), .Z(\mult_26/ab[23][21] ) );
  AND U874 ( .A(e_input[20]), .B(g_input[23]), .Z(\mult_26/ab[23][20] ) );
  AND U875 ( .A(e_input[1]), .B(g_input[23]), .Z(\mult_26/ab[23][1] ) );
  AND U876 ( .A(e_input[19]), .B(g_input[23]), .Z(\mult_26/ab[23][19] ) );
  AND U877 ( .A(e_input[18]), .B(g_input[23]), .Z(\mult_26/ab[23][18] ) );
  AND U878 ( .A(e_input[17]), .B(g_input[23]), .Z(\mult_26/ab[23][17] ) );
  AND U879 ( .A(e_input[16]), .B(g_input[23]), .Z(\mult_26/ab[23][16] ) );
  AND U880 ( .A(e_input[15]), .B(g_input[23]), .Z(\mult_26/ab[23][15] ) );
  AND U881 ( .A(e_input[14]), .B(g_input[23]), .Z(\mult_26/ab[23][14] ) );
  AND U882 ( .A(e_input[13]), .B(g_input[23]), .Z(\mult_26/ab[23][13] ) );
  AND U883 ( .A(e_input[12]), .B(g_input[23]), .Z(\mult_26/ab[23][12] ) );
  AND U884 ( .A(e_input[11]), .B(g_input[23]), .Z(\mult_26/ab[23][11] ) );
  AND U885 ( .A(e_input[10]), .B(g_input[23]), .Z(\mult_26/ab[23][10] ) );
  AND U886 ( .A(g_input[23]), .B(e_input[0]), .Z(\mult_26/ab[23][0] ) );
  AND U887 ( .A(e_input[9]), .B(g_input[22]), .Z(\mult_26/ab[22][9] ) );
  AND U888 ( .A(e_input[8]), .B(g_input[22]), .Z(\mult_26/ab[22][8] ) );
  AND U889 ( .A(e_input[7]), .B(g_input[22]), .Z(\mult_26/ab[22][7] ) );
  AND U890 ( .A(e_input[6]), .B(g_input[22]), .Z(\mult_26/ab[22][6] ) );
  AND U891 ( .A(e_input[5]), .B(g_input[22]), .Z(\mult_26/ab[22][5] ) );
  AND U892 ( .A(e_input[4]), .B(g_input[22]), .Z(\mult_26/ab[22][4] ) );
  AND U893 ( .A(e_input[3]), .B(g_input[22]), .Z(\mult_26/ab[22][3] ) );
  AND U894 ( .A(e_input[31]), .B(g_input[22]), .Z(\mult_26/ab[22][31] ) );
  AND U895 ( .A(e_input[30]), .B(g_input[22]), .Z(\mult_26/ab[22][30] ) );
  AND U896 ( .A(e_input[2]), .B(g_input[22]), .Z(\mult_26/ab[22][2] ) );
  AND U897 ( .A(e_input[29]), .B(g_input[22]), .Z(\mult_26/ab[22][29] ) );
  AND U898 ( .A(e_input[28]), .B(g_input[22]), .Z(\mult_26/ab[22][28] ) );
  AND U899 ( .A(e_input[27]), .B(g_input[22]), .Z(\mult_26/ab[22][27] ) );
  AND U900 ( .A(e_input[26]), .B(g_input[22]), .Z(\mult_26/ab[22][26] ) );
  AND U901 ( .A(e_input[25]), .B(g_input[22]), .Z(\mult_26/ab[22][25] ) );
  AND U902 ( .A(e_input[24]), .B(g_input[22]), .Z(\mult_26/ab[22][24] ) );
  AND U903 ( .A(e_input[23]), .B(g_input[22]), .Z(\mult_26/ab[22][23] ) );
  AND U904 ( .A(e_input[22]), .B(g_input[22]), .Z(\mult_26/ab[22][22] ) );
  AND U905 ( .A(e_input[21]), .B(g_input[22]), .Z(\mult_26/ab[22][21] ) );
  AND U906 ( .A(e_input[20]), .B(g_input[22]), .Z(\mult_26/ab[22][20] ) );
  AND U907 ( .A(e_input[1]), .B(g_input[22]), .Z(\mult_26/ab[22][1] ) );
  AND U908 ( .A(e_input[19]), .B(g_input[22]), .Z(\mult_26/ab[22][19] ) );
  AND U909 ( .A(e_input[18]), .B(g_input[22]), .Z(\mult_26/ab[22][18] ) );
  AND U910 ( .A(e_input[17]), .B(g_input[22]), .Z(\mult_26/ab[22][17] ) );
  AND U911 ( .A(e_input[16]), .B(g_input[22]), .Z(\mult_26/ab[22][16] ) );
  AND U912 ( .A(e_input[15]), .B(g_input[22]), .Z(\mult_26/ab[22][15] ) );
  AND U913 ( .A(e_input[14]), .B(g_input[22]), .Z(\mult_26/ab[22][14] ) );
  AND U914 ( .A(e_input[13]), .B(g_input[22]), .Z(\mult_26/ab[22][13] ) );
  AND U915 ( .A(e_input[12]), .B(g_input[22]), .Z(\mult_26/ab[22][12] ) );
  AND U916 ( .A(e_input[11]), .B(g_input[22]), .Z(\mult_26/ab[22][11] ) );
  AND U917 ( .A(e_input[10]), .B(g_input[22]), .Z(\mult_26/ab[22][10] ) );
  AND U918 ( .A(g_input[22]), .B(e_input[0]), .Z(\mult_26/ab[22][0] ) );
  AND U919 ( .A(e_input[9]), .B(g_input[21]), .Z(\mult_26/ab[21][9] ) );
  AND U920 ( .A(e_input[8]), .B(g_input[21]), .Z(\mult_26/ab[21][8] ) );
  AND U921 ( .A(e_input[7]), .B(g_input[21]), .Z(\mult_26/ab[21][7] ) );
  AND U922 ( .A(e_input[6]), .B(g_input[21]), .Z(\mult_26/ab[21][6] ) );
  AND U923 ( .A(e_input[5]), .B(g_input[21]), .Z(\mult_26/ab[21][5] ) );
  AND U924 ( .A(e_input[4]), .B(g_input[21]), .Z(\mult_26/ab[21][4] ) );
  AND U925 ( .A(e_input[3]), .B(g_input[21]), .Z(\mult_26/ab[21][3] ) );
  AND U926 ( .A(e_input[31]), .B(g_input[21]), .Z(\mult_26/ab[21][31] ) );
  AND U927 ( .A(e_input[30]), .B(g_input[21]), .Z(\mult_26/ab[21][30] ) );
  AND U928 ( .A(e_input[2]), .B(g_input[21]), .Z(\mult_26/ab[21][2] ) );
  AND U929 ( .A(e_input[29]), .B(g_input[21]), .Z(\mult_26/ab[21][29] ) );
  AND U930 ( .A(e_input[28]), .B(g_input[21]), .Z(\mult_26/ab[21][28] ) );
  AND U931 ( .A(e_input[27]), .B(g_input[21]), .Z(\mult_26/ab[21][27] ) );
  AND U932 ( .A(e_input[26]), .B(g_input[21]), .Z(\mult_26/ab[21][26] ) );
  AND U933 ( .A(e_input[25]), .B(g_input[21]), .Z(\mult_26/ab[21][25] ) );
  AND U934 ( .A(e_input[24]), .B(g_input[21]), .Z(\mult_26/ab[21][24] ) );
  AND U935 ( .A(e_input[23]), .B(g_input[21]), .Z(\mult_26/ab[21][23] ) );
  AND U936 ( .A(e_input[22]), .B(g_input[21]), .Z(\mult_26/ab[21][22] ) );
  AND U937 ( .A(e_input[21]), .B(g_input[21]), .Z(\mult_26/ab[21][21] ) );
  AND U938 ( .A(e_input[20]), .B(g_input[21]), .Z(\mult_26/ab[21][20] ) );
  AND U939 ( .A(e_input[1]), .B(g_input[21]), .Z(\mult_26/ab[21][1] ) );
  AND U940 ( .A(e_input[19]), .B(g_input[21]), .Z(\mult_26/ab[21][19] ) );
  AND U941 ( .A(e_input[18]), .B(g_input[21]), .Z(\mult_26/ab[21][18] ) );
  AND U942 ( .A(e_input[17]), .B(g_input[21]), .Z(\mult_26/ab[21][17] ) );
  AND U943 ( .A(e_input[16]), .B(g_input[21]), .Z(\mult_26/ab[21][16] ) );
  AND U944 ( .A(e_input[15]), .B(g_input[21]), .Z(\mult_26/ab[21][15] ) );
  AND U945 ( .A(e_input[14]), .B(g_input[21]), .Z(\mult_26/ab[21][14] ) );
  AND U946 ( .A(e_input[13]), .B(g_input[21]), .Z(\mult_26/ab[21][13] ) );
  AND U947 ( .A(e_input[12]), .B(g_input[21]), .Z(\mult_26/ab[21][12] ) );
  AND U948 ( .A(e_input[11]), .B(g_input[21]), .Z(\mult_26/ab[21][11] ) );
  AND U949 ( .A(e_input[10]), .B(g_input[21]), .Z(\mult_26/ab[21][10] ) );
  AND U950 ( .A(g_input[21]), .B(e_input[0]), .Z(\mult_26/ab[21][0] ) );
  AND U951 ( .A(e_input[9]), .B(g_input[20]), .Z(\mult_26/ab[20][9] ) );
  AND U952 ( .A(e_input[8]), .B(g_input[20]), .Z(\mult_26/ab[20][8] ) );
  AND U953 ( .A(e_input[7]), .B(g_input[20]), .Z(\mult_26/ab[20][7] ) );
  AND U954 ( .A(e_input[6]), .B(g_input[20]), .Z(\mult_26/ab[20][6] ) );
  AND U955 ( .A(e_input[5]), .B(g_input[20]), .Z(\mult_26/ab[20][5] ) );
  AND U956 ( .A(e_input[4]), .B(g_input[20]), .Z(\mult_26/ab[20][4] ) );
  AND U957 ( .A(e_input[3]), .B(g_input[20]), .Z(\mult_26/ab[20][3] ) );
  AND U958 ( .A(e_input[31]), .B(g_input[20]), .Z(\mult_26/ab[20][31] ) );
  AND U959 ( .A(e_input[30]), .B(g_input[20]), .Z(\mult_26/ab[20][30] ) );
  AND U960 ( .A(e_input[2]), .B(g_input[20]), .Z(\mult_26/ab[20][2] ) );
  AND U961 ( .A(e_input[29]), .B(g_input[20]), .Z(\mult_26/ab[20][29] ) );
  AND U962 ( .A(e_input[28]), .B(g_input[20]), .Z(\mult_26/ab[20][28] ) );
  AND U963 ( .A(e_input[27]), .B(g_input[20]), .Z(\mult_26/ab[20][27] ) );
  AND U964 ( .A(e_input[26]), .B(g_input[20]), .Z(\mult_26/ab[20][26] ) );
  AND U965 ( .A(e_input[25]), .B(g_input[20]), .Z(\mult_26/ab[20][25] ) );
  AND U966 ( .A(e_input[24]), .B(g_input[20]), .Z(\mult_26/ab[20][24] ) );
  AND U967 ( .A(e_input[23]), .B(g_input[20]), .Z(\mult_26/ab[20][23] ) );
  AND U968 ( .A(e_input[22]), .B(g_input[20]), .Z(\mult_26/ab[20][22] ) );
  AND U969 ( .A(e_input[21]), .B(g_input[20]), .Z(\mult_26/ab[20][21] ) );
  AND U970 ( .A(e_input[20]), .B(g_input[20]), .Z(\mult_26/ab[20][20] ) );
  AND U971 ( .A(e_input[1]), .B(g_input[20]), .Z(\mult_26/ab[20][1] ) );
  AND U972 ( .A(e_input[19]), .B(g_input[20]), .Z(\mult_26/ab[20][19] ) );
  AND U973 ( .A(e_input[18]), .B(g_input[20]), .Z(\mult_26/ab[20][18] ) );
  AND U974 ( .A(e_input[17]), .B(g_input[20]), .Z(\mult_26/ab[20][17] ) );
  AND U975 ( .A(e_input[16]), .B(g_input[20]), .Z(\mult_26/ab[20][16] ) );
  AND U976 ( .A(e_input[15]), .B(g_input[20]), .Z(\mult_26/ab[20][15] ) );
  AND U977 ( .A(e_input[14]), .B(g_input[20]), .Z(\mult_26/ab[20][14] ) );
  AND U978 ( .A(e_input[13]), .B(g_input[20]), .Z(\mult_26/ab[20][13] ) );
  AND U979 ( .A(e_input[12]), .B(g_input[20]), .Z(\mult_26/ab[20][12] ) );
  AND U980 ( .A(e_input[11]), .B(g_input[20]), .Z(\mult_26/ab[20][11] ) );
  AND U981 ( .A(e_input[10]), .B(g_input[20]), .Z(\mult_26/ab[20][10] ) );
  AND U982 ( .A(g_input[20]), .B(e_input[0]), .Z(\mult_26/ab[20][0] ) );
  AND U983 ( .A(e_input[9]), .B(g_input[1]), .Z(\mult_26/ab[1][9] ) );
  AND U984 ( .A(e_input[8]), .B(g_input[1]), .Z(\mult_26/ab[1][8] ) );
  AND U985 ( .A(e_input[7]), .B(g_input[1]), .Z(\mult_26/ab[1][7] ) );
  AND U986 ( .A(e_input[6]), .B(g_input[1]), .Z(\mult_26/ab[1][6] ) );
  AND U987 ( .A(e_input[5]), .B(g_input[1]), .Z(\mult_26/ab[1][5] ) );
  AND U988 ( .A(e_input[4]), .B(g_input[1]), .Z(\mult_26/ab[1][4] ) );
  AND U989 ( .A(e_input[3]), .B(g_input[1]), .Z(\mult_26/ab[1][3] ) );
  AND U990 ( .A(e_input[31]), .B(g_input[1]), .Z(\mult_26/ab[1][31] ) );
  AND U991 ( .A(e_input[30]), .B(g_input[1]), .Z(\mult_26/ab[1][30] ) );
  AND U992 ( .A(e_input[2]), .B(g_input[1]), .Z(\mult_26/ab[1][2] ) );
  AND U993 ( .A(e_input[29]), .B(g_input[1]), .Z(\mult_26/ab[1][29] ) );
  AND U994 ( .A(e_input[28]), .B(g_input[1]), .Z(\mult_26/ab[1][28] ) );
  AND U995 ( .A(e_input[27]), .B(g_input[1]), .Z(\mult_26/ab[1][27] ) );
  AND U996 ( .A(e_input[26]), .B(g_input[1]), .Z(\mult_26/ab[1][26] ) );
  AND U997 ( .A(e_input[25]), .B(g_input[1]), .Z(\mult_26/ab[1][25] ) );
  AND U998 ( .A(e_input[24]), .B(g_input[1]), .Z(\mult_26/ab[1][24] ) );
  AND U999 ( .A(e_input[23]), .B(g_input[1]), .Z(\mult_26/ab[1][23] ) );
  AND U1000 ( .A(e_input[22]), .B(g_input[1]), .Z(\mult_26/ab[1][22] ) );
  AND U1001 ( .A(e_input[21]), .B(g_input[1]), .Z(\mult_26/ab[1][21] ) );
  AND U1002 ( .A(e_input[20]), .B(g_input[1]), .Z(\mult_26/ab[1][20] ) );
  AND U1003 ( .A(e_input[1]), .B(g_input[1]), .Z(\mult_26/ab[1][1] ) );
  AND U1004 ( .A(e_input[19]), .B(g_input[1]), .Z(\mult_26/ab[1][19] ) );
  AND U1005 ( .A(e_input[18]), .B(g_input[1]), .Z(\mult_26/ab[1][18] ) );
  AND U1006 ( .A(e_input[17]), .B(g_input[1]), .Z(\mult_26/ab[1][17] ) );
  AND U1007 ( .A(e_input[16]), .B(g_input[1]), .Z(\mult_26/ab[1][16] ) );
  AND U1008 ( .A(e_input[15]), .B(g_input[1]), .Z(\mult_26/ab[1][15] ) );
  AND U1009 ( .A(e_input[14]), .B(g_input[1]), .Z(\mult_26/ab[1][14] ) );
  AND U1010 ( .A(e_input[13]), .B(g_input[1]), .Z(\mult_26/ab[1][13] ) );
  AND U1011 ( .A(e_input[12]), .B(g_input[1]), .Z(\mult_26/ab[1][12] ) );
  AND U1012 ( .A(e_input[11]), .B(g_input[1]), .Z(\mult_26/ab[1][11] ) );
  AND U1013 ( .A(e_input[10]), .B(g_input[1]), .Z(\mult_26/ab[1][10] ) );
  AND U1014 ( .A(g_input[1]), .B(e_input[0]), .Z(\mult_26/ab[1][0] ) );
  AND U1015 ( .A(e_input[9]), .B(g_input[19]), .Z(\mult_26/ab[19][9] ) );
  AND U1016 ( .A(e_input[8]), .B(g_input[19]), .Z(\mult_26/ab[19][8] ) );
  AND U1017 ( .A(e_input[7]), .B(g_input[19]), .Z(\mult_26/ab[19][7] ) );
  AND U1018 ( .A(e_input[6]), .B(g_input[19]), .Z(\mult_26/ab[19][6] ) );
  AND U1019 ( .A(e_input[5]), .B(g_input[19]), .Z(\mult_26/ab[19][5] ) );
  AND U1020 ( .A(e_input[4]), .B(g_input[19]), .Z(\mult_26/ab[19][4] ) );
  AND U1021 ( .A(e_input[3]), .B(g_input[19]), .Z(\mult_26/ab[19][3] ) );
  AND U1022 ( .A(e_input[31]), .B(g_input[19]), .Z(\mult_26/ab[19][31] ) );
  AND U1023 ( .A(e_input[30]), .B(g_input[19]), .Z(\mult_26/ab[19][30] ) );
  AND U1024 ( .A(e_input[2]), .B(g_input[19]), .Z(\mult_26/ab[19][2] ) );
  AND U1025 ( .A(e_input[29]), .B(g_input[19]), .Z(\mult_26/ab[19][29] ) );
  AND U1026 ( .A(e_input[28]), .B(g_input[19]), .Z(\mult_26/ab[19][28] ) );
  AND U1027 ( .A(e_input[27]), .B(g_input[19]), .Z(\mult_26/ab[19][27] ) );
  AND U1028 ( .A(e_input[26]), .B(g_input[19]), .Z(\mult_26/ab[19][26] ) );
  AND U1029 ( .A(e_input[25]), .B(g_input[19]), .Z(\mult_26/ab[19][25] ) );
  AND U1030 ( .A(e_input[24]), .B(g_input[19]), .Z(\mult_26/ab[19][24] ) );
  AND U1031 ( .A(e_input[23]), .B(g_input[19]), .Z(\mult_26/ab[19][23] ) );
  AND U1032 ( .A(e_input[22]), .B(g_input[19]), .Z(\mult_26/ab[19][22] ) );
  AND U1033 ( .A(e_input[21]), .B(g_input[19]), .Z(\mult_26/ab[19][21] ) );
  AND U1034 ( .A(e_input[20]), .B(g_input[19]), .Z(\mult_26/ab[19][20] ) );
  AND U1035 ( .A(e_input[1]), .B(g_input[19]), .Z(\mult_26/ab[19][1] ) );
  AND U1036 ( .A(e_input[19]), .B(g_input[19]), .Z(\mult_26/ab[19][19] ) );
  AND U1037 ( .A(e_input[18]), .B(g_input[19]), .Z(\mult_26/ab[19][18] ) );
  AND U1038 ( .A(e_input[17]), .B(g_input[19]), .Z(\mult_26/ab[19][17] ) );
  AND U1039 ( .A(e_input[16]), .B(g_input[19]), .Z(\mult_26/ab[19][16] ) );
  AND U1040 ( .A(e_input[15]), .B(g_input[19]), .Z(\mult_26/ab[19][15] ) );
  AND U1041 ( .A(e_input[14]), .B(g_input[19]), .Z(\mult_26/ab[19][14] ) );
  AND U1042 ( .A(e_input[13]), .B(g_input[19]), .Z(\mult_26/ab[19][13] ) );
  AND U1043 ( .A(e_input[12]), .B(g_input[19]), .Z(\mult_26/ab[19][12] ) );
  AND U1044 ( .A(e_input[11]), .B(g_input[19]), .Z(\mult_26/ab[19][11] ) );
  AND U1045 ( .A(e_input[10]), .B(g_input[19]), .Z(\mult_26/ab[19][10] ) );
  AND U1046 ( .A(g_input[19]), .B(e_input[0]), .Z(\mult_26/ab[19][0] ) );
  AND U1047 ( .A(e_input[9]), .B(g_input[18]), .Z(\mult_26/ab[18][9] ) );
  AND U1048 ( .A(e_input[8]), .B(g_input[18]), .Z(\mult_26/ab[18][8] ) );
  AND U1049 ( .A(e_input[7]), .B(g_input[18]), .Z(\mult_26/ab[18][7] ) );
  AND U1050 ( .A(e_input[6]), .B(g_input[18]), .Z(\mult_26/ab[18][6] ) );
  AND U1051 ( .A(e_input[5]), .B(g_input[18]), .Z(\mult_26/ab[18][5] ) );
  AND U1052 ( .A(e_input[4]), .B(g_input[18]), .Z(\mult_26/ab[18][4] ) );
  AND U1053 ( .A(e_input[3]), .B(g_input[18]), .Z(\mult_26/ab[18][3] ) );
  AND U1054 ( .A(e_input[31]), .B(g_input[18]), .Z(\mult_26/ab[18][31] ) );
  AND U1055 ( .A(e_input[30]), .B(g_input[18]), .Z(\mult_26/ab[18][30] ) );
  AND U1056 ( .A(e_input[2]), .B(g_input[18]), .Z(\mult_26/ab[18][2] ) );
  AND U1057 ( .A(e_input[29]), .B(g_input[18]), .Z(\mult_26/ab[18][29] ) );
  AND U1058 ( .A(e_input[28]), .B(g_input[18]), .Z(\mult_26/ab[18][28] ) );
  AND U1059 ( .A(e_input[27]), .B(g_input[18]), .Z(\mult_26/ab[18][27] ) );
  AND U1060 ( .A(e_input[26]), .B(g_input[18]), .Z(\mult_26/ab[18][26] ) );
  AND U1061 ( .A(e_input[25]), .B(g_input[18]), .Z(\mult_26/ab[18][25] ) );
  AND U1062 ( .A(e_input[24]), .B(g_input[18]), .Z(\mult_26/ab[18][24] ) );
  AND U1063 ( .A(e_input[23]), .B(g_input[18]), .Z(\mult_26/ab[18][23] ) );
  AND U1064 ( .A(e_input[22]), .B(g_input[18]), .Z(\mult_26/ab[18][22] ) );
  AND U1065 ( .A(e_input[21]), .B(g_input[18]), .Z(\mult_26/ab[18][21] ) );
  AND U1066 ( .A(e_input[20]), .B(g_input[18]), .Z(\mult_26/ab[18][20] ) );
  AND U1067 ( .A(e_input[1]), .B(g_input[18]), .Z(\mult_26/ab[18][1] ) );
  AND U1068 ( .A(e_input[19]), .B(g_input[18]), .Z(\mult_26/ab[18][19] ) );
  AND U1069 ( .A(e_input[18]), .B(g_input[18]), .Z(\mult_26/ab[18][18] ) );
  AND U1070 ( .A(e_input[17]), .B(g_input[18]), .Z(\mult_26/ab[18][17] ) );
  AND U1071 ( .A(e_input[16]), .B(g_input[18]), .Z(\mult_26/ab[18][16] ) );
  AND U1072 ( .A(e_input[15]), .B(g_input[18]), .Z(\mult_26/ab[18][15] ) );
  AND U1073 ( .A(e_input[14]), .B(g_input[18]), .Z(\mult_26/ab[18][14] ) );
  AND U1074 ( .A(e_input[13]), .B(g_input[18]), .Z(\mult_26/ab[18][13] ) );
  AND U1075 ( .A(e_input[12]), .B(g_input[18]), .Z(\mult_26/ab[18][12] ) );
  AND U1076 ( .A(e_input[11]), .B(g_input[18]), .Z(\mult_26/ab[18][11] ) );
  AND U1077 ( .A(e_input[10]), .B(g_input[18]), .Z(\mult_26/ab[18][10] ) );
  AND U1078 ( .A(g_input[18]), .B(e_input[0]), .Z(\mult_26/ab[18][0] ) );
  AND U1079 ( .A(e_input[9]), .B(g_input[17]), .Z(\mult_26/ab[17][9] ) );
  AND U1080 ( .A(e_input[8]), .B(g_input[17]), .Z(\mult_26/ab[17][8] ) );
  AND U1081 ( .A(e_input[7]), .B(g_input[17]), .Z(\mult_26/ab[17][7] ) );
  AND U1082 ( .A(e_input[6]), .B(g_input[17]), .Z(\mult_26/ab[17][6] ) );
  AND U1083 ( .A(e_input[5]), .B(g_input[17]), .Z(\mult_26/ab[17][5] ) );
  AND U1084 ( .A(e_input[4]), .B(g_input[17]), .Z(\mult_26/ab[17][4] ) );
  AND U1085 ( .A(e_input[3]), .B(g_input[17]), .Z(\mult_26/ab[17][3] ) );
  AND U1086 ( .A(e_input[31]), .B(g_input[17]), .Z(\mult_26/ab[17][31] ) );
  AND U1087 ( .A(e_input[30]), .B(g_input[17]), .Z(\mult_26/ab[17][30] ) );
  AND U1088 ( .A(e_input[2]), .B(g_input[17]), .Z(\mult_26/ab[17][2] ) );
  AND U1089 ( .A(e_input[29]), .B(g_input[17]), .Z(\mult_26/ab[17][29] ) );
  AND U1090 ( .A(e_input[28]), .B(g_input[17]), .Z(\mult_26/ab[17][28] ) );
  AND U1091 ( .A(e_input[27]), .B(g_input[17]), .Z(\mult_26/ab[17][27] ) );
  AND U1092 ( .A(e_input[26]), .B(g_input[17]), .Z(\mult_26/ab[17][26] ) );
  AND U1093 ( .A(e_input[25]), .B(g_input[17]), .Z(\mult_26/ab[17][25] ) );
  AND U1094 ( .A(e_input[24]), .B(g_input[17]), .Z(\mult_26/ab[17][24] ) );
  AND U1095 ( .A(e_input[23]), .B(g_input[17]), .Z(\mult_26/ab[17][23] ) );
  AND U1096 ( .A(e_input[22]), .B(g_input[17]), .Z(\mult_26/ab[17][22] ) );
  AND U1097 ( .A(e_input[21]), .B(g_input[17]), .Z(\mult_26/ab[17][21] ) );
  AND U1098 ( .A(e_input[20]), .B(g_input[17]), .Z(\mult_26/ab[17][20] ) );
  AND U1099 ( .A(e_input[1]), .B(g_input[17]), .Z(\mult_26/ab[17][1] ) );
  AND U1100 ( .A(e_input[19]), .B(g_input[17]), .Z(\mult_26/ab[17][19] ) );
  AND U1101 ( .A(e_input[18]), .B(g_input[17]), .Z(\mult_26/ab[17][18] ) );
  AND U1102 ( .A(e_input[17]), .B(g_input[17]), .Z(\mult_26/ab[17][17] ) );
  AND U1103 ( .A(e_input[16]), .B(g_input[17]), .Z(\mult_26/ab[17][16] ) );
  AND U1104 ( .A(e_input[15]), .B(g_input[17]), .Z(\mult_26/ab[17][15] ) );
  AND U1105 ( .A(e_input[14]), .B(g_input[17]), .Z(\mult_26/ab[17][14] ) );
  AND U1106 ( .A(e_input[13]), .B(g_input[17]), .Z(\mult_26/ab[17][13] ) );
  AND U1107 ( .A(e_input[12]), .B(g_input[17]), .Z(\mult_26/ab[17][12] ) );
  AND U1108 ( .A(e_input[11]), .B(g_input[17]), .Z(\mult_26/ab[17][11] ) );
  AND U1109 ( .A(e_input[10]), .B(g_input[17]), .Z(\mult_26/ab[17][10] ) );
  AND U1110 ( .A(g_input[17]), .B(e_input[0]), .Z(\mult_26/ab[17][0] ) );
  AND U1111 ( .A(e_input[9]), .B(g_input[16]), .Z(\mult_26/ab[16][9] ) );
  AND U1112 ( .A(e_input[8]), .B(g_input[16]), .Z(\mult_26/ab[16][8] ) );
  AND U1113 ( .A(e_input[7]), .B(g_input[16]), .Z(\mult_26/ab[16][7] ) );
  AND U1114 ( .A(e_input[6]), .B(g_input[16]), .Z(\mult_26/ab[16][6] ) );
  AND U1115 ( .A(e_input[5]), .B(g_input[16]), .Z(\mult_26/ab[16][5] ) );
  AND U1116 ( .A(e_input[4]), .B(g_input[16]), .Z(\mult_26/ab[16][4] ) );
  AND U1117 ( .A(e_input[3]), .B(g_input[16]), .Z(\mult_26/ab[16][3] ) );
  AND U1118 ( .A(e_input[31]), .B(g_input[16]), .Z(\mult_26/ab[16][31] ) );
  AND U1119 ( .A(e_input[30]), .B(g_input[16]), .Z(\mult_26/ab[16][30] ) );
  AND U1120 ( .A(e_input[2]), .B(g_input[16]), .Z(\mult_26/ab[16][2] ) );
  AND U1121 ( .A(e_input[29]), .B(g_input[16]), .Z(\mult_26/ab[16][29] ) );
  AND U1122 ( .A(e_input[28]), .B(g_input[16]), .Z(\mult_26/ab[16][28] ) );
  AND U1123 ( .A(e_input[27]), .B(g_input[16]), .Z(\mult_26/ab[16][27] ) );
  AND U1124 ( .A(e_input[26]), .B(g_input[16]), .Z(\mult_26/ab[16][26] ) );
  AND U1125 ( .A(e_input[25]), .B(g_input[16]), .Z(\mult_26/ab[16][25] ) );
  AND U1126 ( .A(e_input[24]), .B(g_input[16]), .Z(\mult_26/ab[16][24] ) );
  AND U1127 ( .A(e_input[23]), .B(g_input[16]), .Z(\mult_26/ab[16][23] ) );
  AND U1128 ( .A(e_input[22]), .B(g_input[16]), .Z(\mult_26/ab[16][22] ) );
  AND U1129 ( .A(e_input[21]), .B(g_input[16]), .Z(\mult_26/ab[16][21] ) );
  AND U1130 ( .A(e_input[20]), .B(g_input[16]), .Z(\mult_26/ab[16][20] ) );
  AND U1131 ( .A(e_input[1]), .B(g_input[16]), .Z(\mult_26/ab[16][1] ) );
  AND U1132 ( .A(e_input[19]), .B(g_input[16]), .Z(\mult_26/ab[16][19] ) );
  AND U1133 ( .A(e_input[18]), .B(g_input[16]), .Z(\mult_26/ab[16][18] ) );
  AND U1134 ( .A(e_input[17]), .B(g_input[16]), .Z(\mult_26/ab[16][17] ) );
  AND U1135 ( .A(e_input[16]), .B(g_input[16]), .Z(\mult_26/ab[16][16] ) );
  AND U1136 ( .A(e_input[15]), .B(g_input[16]), .Z(\mult_26/ab[16][15] ) );
  AND U1137 ( .A(e_input[14]), .B(g_input[16]), .Z(\mult_26/ab[16][14] ) );
  AND U1138 ( .A(e_input[13]), .B(g_input[16]), .Z(\mult_26/ab[16][13] ) );
  AND U1139 ( .A(e_input[12]), .B(g_input[16]), .Z(\mult_26/ab[16][12] ) );
  AND U1140 ( .A(e_input[11]), .B(g_input[16]), .Z(\mult_26/ab[16][11] ) );
  AND U1141 ( .A(e_input[10]), .B(g_input[16]), .Z(\mult_26/ab[16][10] ) );
  AND U1142 ( .A(g_input[16]), .B(e_input[0]), .Z(\mult_26/ab[16][0] ) );
  AND U1143 ( .A(e_input[9]), .B(g_input[15]), .Z(\mult_26/ab[15][9] ) );
  AND U1144 ( .A(e_input[8]), .B(g_input[15]), .Z(\mult_26/ab[15][8] ) );
  AND U1145 ( .A(e_input[7]), .B(g_input[15]), .Z(\mult_26/ab[15][7] ) );
  AND U1146 ( .A(e_input[6]), .B(g_input[15]), .Z(\mult_26/ab[15][6] ) );
  AND U1147 ( .A(e_input[5]), .B(g_input[15]), .Z(\mult_26/ab[15][5] ) );
  AND U1148 ( .A(e_input[4]), .B(g_input[15]), .Z(\mult_26/ab[15][4] ) );
  AND U1149 ( .A(e_input[3]), .B(g_input[15]), .Z(\mult_26/ab[15][3] ) );
  AND U1150 ( .A(e_input[31]), .B(g_input[15]), .Z(\mult_26/ab[15][31] ) );
  AND U1151 ( .A(e_input[30]), .B(g_input[15]), .Z(\mult_26/ab[15][30] ) );
  AND U1152 ( .A(e_input[2]), .B(g_input[15]), .Z(\mult_26/ab[15][2] ) );
  AND U1153 ( .A(e_input[29]), .B(g_input[15]), .Z(\mult_26/ab[15][29] ) );
  AND U1154 ( .A(e_input[28]), .B(g_input[15]), .Z(\mult_26/ab[15][28] ) );
  AND U1155 ( .A(e_input[27]), .B(g_input[15]), .Z(\mult_26/ab[15][27] ) );
  AND U1156 ( .A(e_input[26]), .B(g_input[15]), .Z(\mult_26/ab[15][26] ) );
  AND U1157 ( .A(e_input[25]), .B(g_input[15]), .Z(\mult_26/ab[15][25] ) );
  AND U1158 ( .A(e_input[24]), .B(g_input[15]), .Z(\mult_26/ab[15][24] ) );
  AND U1159 ( .A(e_input[23]), .B(g_input[15]), .Z(\mult_26/ab[15][23] ) );
  AND U1160 ( .A(e_input[22]), .B(g_input[15]), .Z(\mult_26/ab[15][22] ) );
  AND U1161 ( .A(e_input[21]), .B(g_input[15]), .Z(\mult_26/ab[15][21] ) );
  AND U1162 ( .A(e_input[20]), .B(g_input[15]), .Z(\mult_26/ab[15][20] ) );
  AND U1163 ( .A(e_input[1]), .B(g_input[15]), .Z(\mult_26/ab[15][1] ) );
  AND U1164 ( .A(e_input[19]), .B(g_input[15]), .Z(\mult_26/ab[15][19] ) );
  AND U1165 ( .A(e_input[18]), .B(g_input[15]), .Z(\mult_26/ab[15][18] ) );
  AND U1166 ( .A(e_input[17]), .B(g_input[15]), .Z(\mult_26/ab[15][17] ) );
  AND U1167 ( .A(e_input[16]), .B(g_input[15]), .Z(\mult_26/ab[15][16] ) );
  AND U1168 ( .A(e_input[15]), .B(g_input[15]), .Z(\mult_26/ab[15][15] ) );
  AND U1169 ( .A(e_input[14]), .B(g_input[15]), .Z(\mult_26/ab[15][14] ) );
  AND U1170 ( .A(e_input[13]), .B(g_input[15]), .Z(\mult_26/ab[15][13] ) );
  AND U1171 ( .A(e_input[12]), .B(g_input[15]), .Z(\mult_26/ab[15][12] ) );
  AND U1172 ( .A(e_input[11]), .B(g_input[15]), .Z(\mult_26/ab[15][11] ) );
  AND U1173 ( .A(e_input[10]), .B(g_input[15]), .Z(\mult_26/ab[15][10] ) );
  AND U1174 ( .A(g_input[15]), .B(e_input[0]), .Z(\mult_26/ab[15][0] ) );
  AND U1175 ( .A(e_input[9]), .B(g_input[14]), .Z(\mult_26/ab[14][9] ) );
  AND U1176 ( .A(e_input[8]), .B(g_input[14]), .Z(\mult_26/ab[14][8] ) );
  AND U1177 ( .A(e_input[7]), .B(g_input[14]), .Z(\mult_26/ab[14][7] ) );
  AND U1178 ( .A(e_input[6]), .B(g_input[14]), .Z(\mult_26/ab[14][6] ) );
  AND U1179 ( .A(e_input[5]), .B(g_input[14]), .Z(\mult_26/ab[14][5] ) );
  AND U1180 ( .A(e_input[4]), .B(g_input[14]), .Z(\mult_26/ab[14][4] ) );
  AND U1181 ( .A(e_input[3]), .B(g_input[14]), .Z(\mult_26/ab[14][3] ) );
  AND U1182 ( .A(e_input[31]), .B(g_input[14]), .Z(\mult_26/ab[14][31] ) );
  AND U1183 ( .A(e_input[30]), .B(g_input[14]), .Z(\mult_26/ab[14][30] ) );
  AND U1184 ( .A(e_input[2]), .B(g_input[14]), .Z(\mult_26/ab[14][2] ) );
  AND U1185 ( .A(e_input[29]), .B(g_input[14]), .Z(\mult_26/ab[14][29] ) );
  AND U1186 ( .A(e_input[28]), .B(g_input[14]), .Z(\mult_26/ab[14][28] ) );
  AND U1187 ( .A(e_input[27]), .B(g_input[14]), .Z(\mult_26/ab[14][27] ) );
  AND U1188 ( .A(e_input[26]), .B(g_input[14]), .Z(\mult_26/ab[14][26] ) );
  AND U1189 ( .A(e_input[25]), .B(g_input[14]), .Z(\mult_26/ab[14][25] ) );
  AND U1190 ( .A(e_input[24]), .B(g_input[14]), .Z(\mult_26/ab[14][24] ) );
  AND U1191 ( .A(e_input[23]), .B(g_input[14]), .Z(\mult_26/ab[14][23] ) );
  AND U1192 ( .A(e_input[22]), .B(g_input[14]), .Z(\mult_26/ab[14][22] ) );
  AND U1193 ( .A(e_input[21]), .B(g_input[14]), .Z(\mult_26/ab[14][21] ) );
  AND U1194 ( .A(e_input[20]), .B(g_input[14]), .Z(\mult_26/ab[14][20] ) );
  AND U1195 ( .A(e_input[1]), .B(g_input[14]), .Z(\mult_26/ab[14][1] ) );
  AND U1196 ( .A(e_input[19]), .B(g_input[14]), .Z(\mult_26/ab[14][19] ) );
  AND U1197 ( .A(e_input[18]), .B(g_input[14]), .Z(\mult_26/ab[14][18] ) );
  AND U1198 ( .A(e_input[17]), .B(g_input[14]), .Z(\mult_26/ab[14][17] ) );
  AND U1199 ( .A(e_input[16]), .B(g_input[14]), .Z(\mult_26/ab[14][16] ) );
  AND U1200 ( .A(e_input[15]), .B(g_input[14]), .Z(\mult_26/ab[14][15] ) );
  AND U1201 ( .A(e_input[14]), .B(g_input[14]), .Z(\mult_26/ab[14][14] ) );
  AND U1202 ( .A(e_input[13]), .B(g_input[14]), .Z(\mult_26/ab[14][13] ) );
  AND U1203 ( .A(e_input[12]), .B(g_input[14]), .Z(\mult_26/ab[14][12] ) );
  AND U1204 ( .A(e_input[11]), .B(g_input[14]), .Z(\mult_26/ab[14][11] ) );
  AND U1205 ( .A(e_input[10]), .B(g_input[14]), .Z(\mult_26/ab[14][10] ) );
  AND U1206 ( .A(g_input[14]), .B(e_input[0]), .Z(\mult_26/ab[14][0] ) );
  AND U1207 ( .A(e_input[9]), .B(g_input[13]), .Z(\mult_26/ab[13][9] ) );
  AND U1208 ( .A(e_input[8]), .B(g_input[13]), .Z(\mult_26/ab[13][8] ) );
  AND U1209 ( .A(e_input[7]), .B(g_input[13]), .Z(\mult_26/ab[13][7] ) );
  AND U1210 ( .A(e_input[6]), .B(g_input[13]), .Z(\mult_26/ab[13][6] ) );
  AND U1211 ( .A(e_input[5]), .B(g_input[13]), .Z(\mult_26/ab[13][5] ) );
  AND U1212 ( .A(e_input[4]), .B(g_input[13]), .Z(\mult_26/ab[13][4] ) );
  AND U1213 ( .A(e_input[3]), .B(g_input[13]), .Z(\mult_26/ab[13][3] ) );
  AND U1214 ( .A(e_input[31]), .B(g_input[13]), .Z(\mult_26/ab[13][31] ) );
  AND U1215 ( .A(e_input[30]), .B(g_input[13]), .Z(\mult_26/ab[13][30] ) );
  AND U1216 ( .A(e_input[2]), .B(g_input[13]), .Z(\mult_26/ab[13][2] ) );
  AND U1217 ( .A(e_input[29]), .B(g_input[13]), .Z(\mult_26/ab[13][29] ) );
  AND U1218 ( .A(e_input[28]), .B(g_input[13]), .Z(\mult_26/ab[13][28] ) );
  AND U1219 ( .A(e_input[27]), .B(g_input[13]), .Z(\mult_26/ab[13][27] ) );
  AND U1220 ( .A(e_input[26]), .B(g_input[13]), .Z(\mult_26/ab[13][26] ) );
  AND U1221 ( .A(e_input[25]), .B(g_input[13]), .Z(\mult_26/ab[13][25] ) );
  AND U1222 ( .A(e_input[24]), .B(g_input[13]), .Z(\mult_26/ab[13][24] ) );
  AND U1223 ( .A(e_input[23]), .B(g_input[13]), .Z(\mult_26/ab[13][23] ) );
  AND U1224 ( .A(e_input[22]), .B(g_input[13]), .Z(\mult_26/ab[13][22] ) );
  AND U1225 ( .A(e_input[21]), .B(g_input[13]), .Z(\mult_26/ab[13][21] ) );
  AND U1226 ( .A(e_input[20]), .B(g_input[13]), .Z(\mult_26/ab[13][20] ) );
  AND U1227 ( .A(e_input[1]), .B(g_input[13]), .Z(\mult_26/ab[13][1] ) );
  AND U1228 ( .A(e_input[19]), .B(g_input[13]), .Z(\mult_26/ab[13][19] ) );
  AND U1229 ( .A(e_input[18]), .B(g_input[13]), .Z(\mult_26/ab[13][18] ) );
  AND U1230 ( .A(e_input[17]), .B(g_input[13]), .Z(\mult_26/ab[13][17] ) );
  AND U1231 ( .A(e_input[16]), .B(g_input[13]), .Z(\mult_26/ab[13][16] ) );
  AND U1232 ( .A(e_input[15]), .B(g_input[13]), .Z(\mult_26/ab[13][15] ) );
  AND U1233 ( .A(e_input[14]), .B(g_input[13]), .Z(\mult_26/ab[13][14] ) );
  AND U1234 ( .A(e_input[13]), .B(g_input[13]), .Z(\mult_26/ab[13][13] ) );
  AND U1235 ( .A(e_input[12]), .B(g_input[13]), .Z(\mult_26/ab[13][12] ) );
  AND U1236 ( .A(e_input[11]), .B(g_input[13]), .Z(\mult_26/ab[13][11] ) );
  AND U1237 ( .A(e_input[10]), .B(g_input[13]), .Z(\mult_26/ab[13][10] ) );
  AND U1238 ( .A(g_input[13]), .B(e_input[0]), .Z(\mult_26/ab[13][0] ) );
  AND U1239 ( .A(e_input[9]), .B(g_input[12]), .Z(\mult_26/ab[12][9] ) );
  AND U1240 ( .A(e_input[8]), .B(g_input[12]), .Z(\mult_26/ab[12][8] ) );
  AND U1241 ( .A(e_input[7]), .B(g_input[12]), .Z(\mult_26/ab[12][7] ) );
  AND U1242 ( .A(e_input[6]), .B(g_input[12]), .Z(\mult_26/ab[12][6] ) );
  AND U1243 ( .A(e_input[5]), .B(g_input[12]), .Z(\mult_26/ab[12][5] ) );
  AND U1244 ( .A(e_input[4]), .B(g_input[12]), .Z(\mult_26/ab[12][4] ) );
  AND U1245 ( .A(e_input[3]), .B(g_input[12]), .Z(\mult_26/ab[12][3] ) );
  AND U1246 ( .A(e_input[31]), .B(g_input[12]), .Z(\mult_26/ab[12][31] ) );
  AND U1247 ( .A(e_input[30]), .B(g_input[12]), .Z(\mult_26/ab[12][30] ) );
  AND U1248 ( .A(e_input[2]), .B(g_input[12]), .Z(\mult_26/ab[12][2] ) );
  AND U1249 ( .A(e_input[29]), .B(g_input[12]), .Z(\mult_26/ab[12][29] ) );
  AND U1250 ( .A(e_input[28]), .B(g_input[12]), .Z(\mult_26/ab[12][28] ) );
  AND U1251 ( .A(e_input[27]), .B(g_input[12]), .Z(\mult_26/ab[12][27] ) );
  AND U1252 ( .A(e_input[26]), .B(g_input[12]), .Z(\mult_26/ab[12][26] ) );
  AND U1253 ( .A(e_input[25]), .B(g_input[12]), .Z(\mult_26/ab[12][25] ) );
  AND U1254 ( .A(e_input[24]), .B(g_input[12]), .Z(\mult_26/ab[12][24] ) );
  AND U1255 ( .A(e_input[23]), .B(g_input[12]), .Z(\mult_26/ab[12][23] ) );
  AND U1256 ( .A(e_input[22]), .B(g_input[12]), .Z(\mult_26/ab[12][22] ) );
  AND U1257 ( .A(e_input[21]), .B(g_input[12]), .Z(\mult_26/ab[12][21] ) );
  AND U1258 ( .A(e_input[20]), .B(g_input[12]), .Z(\mult_26/ab[12][20] ) );
  AND U1259 ( .A(e_input[1]), .B(g_input[12]), .Z(\mult_26/ab[12][1] ) );
  AND U1260 ( .A(e_input[19]), .B(g_input[12]), .Z(\mult_26/ab[12][19] ) );
  AND U1261 ( .A(e_input[18]), .B(g_input[12]), .Z(\mult_26/ab[12][18] ) );
  AND U1262 ( .A(e_input[17]), .B(g_input[12]), .Z(\mult_26/ab[12][17] ) );
  AND U1263 ( .A(e_input[16]), .B(g_input[12]), .Z(\mult_26/ab[12][16] ) );
  AND U1264 ( .A(e_input[15]), .B(g_input[12]), .Z(\mult_26/ab[12][15] ) );
  AND U1265 ( .A(e_input[14]), .B(g_input[12]), .Z(\mult_26/ab[12][14] ) );
  AND U1266 ( .A(e_input[13]), .B(g_input[12]), .Z(\mult_26/ab[12][13] ) );
  AND U1267 ( .A(e_input[12]), .B(g_input[12]), .Z(\mult_26/ab[12][12] ) );
  AND U1268 ( .A(e_input[11]), .B(g_input[12]), .Z(\mult_26/ab[12][11] ) );
  AND U1269 ( .A(e_input[10]), .B(g_input[12]), .Z(\mult_26/ab[12][10] ) );
  AND U1270 ( .A(g_input[12]), .B(e_input[0]), .Z(\mult_26/ab[12][0] ) );
  AND U1271 ( .A(e_input[9]), .B(g_input[11]), .Z(\mult_26/ab[11][9] ) );
  AND U1272 ( .A(e_input[8]), .B(g_input[11]), .Z(\mult_26/ab[11][8] ) );
  AND U1273 ( .A(e_input[7]), .B(g_input[11]), .Z(\mult_26/ab[11][7] ) );
  AND U1274 ( .A(e_input[6]), .B(g_input[11]), .Z(\mult_26/ab[11][6] ) );
  AND U1275 ( .A(e_input[5]), .B(g_input[11]), .Z(\mult_26/ab[11][5] ) );
  AND U1276 ( .A(e_input[4]), .B(g_input[11]), .Z(\mult_26/ab[11][4] ) );
  AND U1277 ( .A(e_input[3]), .B(g_input[11]), .Z(\mult_26/ab[11][3] ) );
  AND U1278 ( .A(e_input[31]), .B(g_input[11]), .Z(\mult_26/ab[11][31] ) );
  AND U1279 ( .A(e_input[30]), .B(g_input[11]), .Z(\mult_26/ab[11][30] ) );
  AND U1280 ( .A(e_input[2]), .B(g_input[11]), .Z(\mult_26/ab[11][2] ) );
  AND U1281 ( .A(e_input[29]), .B(g_input[11]), .Z(\mult_26/ab[11][29] ) );
  AND U1282 ( .A(e_input[28]), .B(g_input[11]), .Z(\mult_26/ab[11][28] ) );
  AND U1283 ( .A(e_input[27]), .B(g_input[11]), .Z(\mult_26/ab[11][27] ) );
  AND U1284 ( .A(e_input[26]), .B(g_input[11]), .Z(\mult_26/ab[11][26] ) );
  AND U1285 ( .A(e_input[25]), .B(g_input[11]), .Z(\mult_26/ab[11][25] ) );
  AND U1286 ( .A(e_input[24]), .B(g_input[11]), .Z(\mult_26/ab[11][24] ) );
  AND U1287 ( .A(e_input[23]), .B(g_input[11]), .Z(\mult_26/ab[11][23] ) );
  AND U1288 ( .A(e_input[22]), .B(g_input[11]), .Z(\mult_26/ab[11][22] ) );
  AND U1289 ( .A(e_input[21]), .B(g_input[11]), .Z(\mult_26/ab[11][21] ) );
  AND U1290 ( .A(e_input[20]), .B(g_input[11]), .Z(\mult_26/ab[11][20] ) );
  AND U1291 ( .A(e_input[1]), .B(g_input[11]), .Z(\mult_26/ab[11][1] ) );
  AND U1292 ( .A(e_input[19]), .B(g_input[11]), .Z(\mult_26/ab[11][19] ) );
  AND U1293 ( .A(e_input[18]), .B(g_input[11]), .Z(\mult_26/ab[11][18] ) );
  AND U1294 ( .A(e_input[17]), .B(g_input[11]), .Z(\mult_26/ab[11][17] ) );
  AND U1295 ( .A(e_input[16]), .B(g_input[11]), .Z(\mult_26/ab[11][16] ) );
  AND U1296 ( .A(e_input[15]), .B(g_input[11]), .Z(\mult_26/ab[11][15] ) );
  AND U1297 ( .A(e_input[14]), .B(g_input[11]), .Z(\mult_26/ab[11][14] ) );
  AND U1298 ( .A(e_input[13]), .B(g_input[11]), .Z(\mult_26/ab[11][13] ) );
  AND U1299 ( .A(e_input[12]), .B(g_input[11]), .Z(\mult_26/ab[11][12] ) );
  AND U1300 ( .A(e_input[11]), .B(g_input[11]), .Z(\mult_26/ab[11][11] ) );
  AND U1301 ( .A(e_input[10]), .B(g_input[11]), .Z(\mult_26/ab[11][10] ) );
  AND U1302 ( .A(g_input[11]), .B(e_input[0]), .Z(\mult_26/ab[11][0] ) );
  AND U1303 ( .A(e_input[9]), .B(g_input[10]), .Z(\mult_26/ab[10][9] ) );
  AND U1304 ( .A(e_input[8]), .B(g_input[10]), .Z(\mult_26/ab[10][8] ) );
  AND U1305 ( .A(e_input[7]), .B(g_input[10]), .Z(\mult_26/ab[10][7] ) );
  AND U1306 ( .A(e_input[6]), .B(g_input[10]), .Z(\mult_26/ab[10][6] ) );
  AND U1307 ( .A(e_input[5]), .B(g_input[10]), .Z(\mult_26/ab[10][5] ) );
  AND U1308 ( .A(e_input[4]), .B(g_input[10]), .Z(\mult_26/ab[10][4] ) );
  AND U1309 ( .A(e_input[3]), .B(g_input[10]), .Z(\mult_26/ab[10][3] ) );
  AND U1310 ( .A(e_input[31]), .B(g_input[10]), .Z(\mult_26/ab[10][31] ) );
  AND U1311 ( .A(e_input[30]), .B(g_input[10]), .Z(\mult_26/ab[10][30] ) );
  AND U1312 ( .A(e_input[2]), .B(g_input[10]), .Z(\mult_26/ab[10][2] ) );
  AND U1313 ( .A(e_input[29]), .B(g_input[10]), .Z(\mult_26/ab[10][29] ) );
  AND U1314 ( .A(e_input[28]), .B(g_input[10]), .Z(\mult_26/ab[10][28] ) );
  AND U1315 ( .A(e_input[27]), .B(g_input[10]), .Z(\mult_26/ab[10][27] ) );
  AND U1316 ( .A(e_input[26]), .B(g_input[10]), .Z(\mult_26/ab[10][26] ) );
  AND U1317 ( .A(e_input[25]), .B(g_input[10]), .Z(\mult_26/ab[10][25] ) );
  AND U1318 ( .A(e_input[24]), .B(g_input[10]), .Z(\mult_26/ab[10][24] ) );
  AND U1319 ( .A(e_input[23]), .B(g_input[10]), .Z(\mult_26/ab[10][23] ) );
  AND U1320 ( .A(e_input[22]), .B(g_input[10]), .Z(\mult_26/ab[10][22] ) );
  AND U1321 ( .A(e_input[21]), .B(g_input[10]), .Z(\mult_26/ab[10][21] ) );
  AND U1322 ( .A(e_input[20]), .B(g_input[10]), .Z(\mult_26/ab[10][20] ) );
  AND U1323 ( .A(e_input[1]), .B(g_input[10]), .Z(\mult_26/ab[10][1] ) );
  AND U1324 ( .A(e_input[19]), .B(g_input[10]), .Z(\mult_26/ab[10][19] ) );
  AND U1325 ( .A(e_input[18]), .B(g_input[10]), .Z(\mult_26/ab[10][18] ) );
  AND U1326 ( .A(e_input[17]), .B(g_input[10]), .Z(\mult_26/ab[10][17] ) );
  AND U1327 ( .A(e_input[16]), .B(g_input[10]), .Z(\mult_26/ab[10][16] ) );
  AND U1328 ( .A(e_input[15]), .B(g_input[10]), .Z(\mult_26/ab[10][15] ) );
  AND U1329 ( .A(e_input[14]), .B(g_input[10]), .Z(\mult_26/ab[10][14] ) );
  AND U1330 ( .A(e_input[13]), .B(g_input[10]), .Z(\mult_26/ab[10][13] ) );
  AND U1331 ( .A(e_input[12]), .B(g_input[10]), .Z(\mult_26/ab[10][12] ) );
  AND U1332 ( .A(e_input[11]), .B(g_input[10]), .Z(\mult_26/ab[10][11] ) );
  AND U1333 ( .A(e_input[10]), .B(g_input[10]), .Z(\mult_26/ab[10][10] ) );
  AND U1334 ( .A(g_input[10]), .B(e_input[0]), .Z(\mult_26/ab[10][0] ) );
  AND U1335 ( .A(g_input[0]), .B(e_input[9]), .Z(\mult_26/ab[0][9] ) );
  AND U1336 ( .A(g_input[0]), .B(e_input[8]), .Z(\mult_26/ab[0][8] ) );
  AND U1337 ( .A(g_input[0]), .B(e_input[7]), .Z(\mult_26/ab[0][7] ) );
  AND U1338 ( .A(g_input[0]), .B(e_input[6]), .Z(\mult_26/ab[0][6] ) );
  AND U1339 ( .A(g_input[0]), .B(e_input[5]), .Z(\mult_26/ab[0][5] ) );
  AND U1340 ( .A(g_input[0]), .B(e_input[4]), .Z(\mult_26/ab[0][4] ) );
  AND U1341 ( .A(g_input[0]), .B(e_input[3]), .Z(\mult_26/ab[0][3] ) );
  AND U1342 ( .A(g_input[0]), .B(e_input[31]), .Z(\mult_26/ab[0][31] ) );
  AND U1343 ( .A(g_input[0]), .B(e_input[30]), .Z(\mult_26/ab[0][30] ) );
  AND U1344 ( .A(g_input[0]), .B(e_input[2]), .Z(\mult_26/ab[0][2] ) );
  AND U1345 ( .A(g_input[0]), .B(e_input[29]), .Z(\mult_26/ab[0][29] ) );
  AND U1346 ( .A(g_input[0]), .B(e_input[28]), .Z(\mult_26/ab[0][28] ) );
  AND U1347 ( .A(g_input[0]), .B(e_input[27]), .Z(\mult_26/ab[0][27] ) );
  AND U1348 ( .A(g_input[0]), .B(e_input[26]), .Z(\mult_26/ab[0][26] ) );
  AND U1349 ( .A(g_input[0]), .B(e_input[25]), .Z(\mult_26/ab[0][25] ) );
  AND U1350 ( .A(g_input[0]), .B(e_input[24]), .Z(\mult_26/ab[0][24] ) );
  AND U1351 ( .A(g_input[0]), .B(e_input[23]), .Z(\mult_26/ab[0][23] ) );
  AND U1352 ( .A(g_input[0]), .B(e_input[22]), .Z(\mult_26/ab[0][22] ) );
  AND U1353 ( .A(g_input[0]), .B(e_input[21]), .Z(\mult_26/ab[0][21] ) );
  AND U1354 ( .A(g_input[0]), .B(e_input[20]), .Z(\mult_26/ab[0][20] ) );
  AND U1355 ( .A(g_input[0]), .B(e_input[1]), .Z(\mult_26/ab[0][1] ) );
  AND U1356 ( .A(g_input[0]), .B(e_input[19]), .Z(\mult_26/ab[0][19] ) );
  AND U1357 ( .A(g_input[0]), .B(e_input[18]), .Z(\mult_26/ab[0][18] ) );
  AND U1358 ( .A(g_input[0]), .B(e_input[17]), .Z(\mult_26/ab[0][17] ) );
  AND U1359 ( .A(g_input[0]), .B(e_input[16]), .Z(\mult_26/ab[0][16] ) );
  AND U1360 ( .A(g_input[0]), .B(e_input[15]), .Z(\mult_26/ab[0][15] ) );
  AND U1361 ( .A(g_input[0]), .B(e_input[14]), .Z(\mult_26/ab[0][14] ) );
  AND U1362 ( .A(g_input[0]), .B(e_input[13]), .Z(\mult_26/ab[0][13] ) );
  AND U1363 ( .A(g_input[0]), .B(e_input[12]), .Z(\mult_26/ab[0][12] ) );
  AND U1364 ( .A(g_input[0]), .B(e_input[11]), .Z(\mult_26/ab[0][11] ) );
  AND U1365 ( .A(g_input[0]), .B(e_input[10]), .Z(\mult_26/ab[0][10] ) );
endmodule

