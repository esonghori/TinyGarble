
module mult_N128_CC4 ( clk, rst, a, b, c );
  input [127:0] a;
  input [31:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329;
  wire   [127:32] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U35 ( .A(n5993), .B(n6156), .Z(n6002) );
  XNOR U36 ( .A(n8165), .B(n8256), .Z(n8174) );
  XNOR U37 ( .A(n848), .B(n938), .Z(n852) );
  XNOR U38 ( .A(n6003), .B(n6155), .Z(n6007) );
  XNOR U39 ( .A(n5842), .B(n5976), .Z(n5846) );
  XNOR U40 ( .A(n6194), .B(n6328), .Z(n6198) );
  XNOR U41 ( .A(n6546), .B(n6680), .Z(n6550) );
  XNOR U42 ( .A(n6033), .B(n6149), .Z(n6037) );
  XNOR U43 ( .A(n6385), .B(n6501), .Z(n6389) );
  XNOR U44 ( .A(n6737), .B(n6853), .Z(n6741) );
  XNOR U45 ( .A(n7089), .B(n7205), .Z(n7093) );
  XNOR U46 ( .A(n1379), .B(n1482), .Z(n1383) );
  XNOR U47 ( .A(n1740), .B(n1843), .Z(n1744) );
  XNOR U48 ( .A(n5872), .B(n5970), .Z(n5876) );
  XNOR U49 ( .A(n6224), .B(n6322), .Z(n6228) );
  XNOR U50 ( .A(n6576), .B(n6674), .Z(n6580) );
  XNOR U51 ( .A(n6928), .B(n7026), .Z(n6932) );
  XNOR U52 ( .A(n7280), .B(n7378), .Z(n7284) );
  XNOR U53 ( .A(n7632), .B(n7730), .Z(n7636) );
  XNOR U54 ( .A(n6063), .B(n6143), .Z(n6067) );
  XNOR U55 ( .A(n6415), .B(n6495), .Z(n6419) );
  XNOR U56 ( .A(n6767), .B(n6847), .Z(n6771) );
  XNOR U57 ( .A(n7119), .B(n7199), .Z(n7123) );
  XNOR U58 ( .A(n7471), .B(n7551), .Z(n7475) );
  XNOR U59 ( .A(n7823), .B(n7903), .Z(n7827) );
  XNOR U60 ( .A(n8175), .B(n8255), .Z(n8179) );
  XNOR U61 ( .A(n1038), .B(n1117), .Z(n1042) );
  XNOR U62 ( .A(n5902), .B(n5964), .Z(n5906) );
  XNOR U63 ( .A(n6254), .B(n6316), .Z(n6258) );
  XNOR U64 ( .A(n6606), .B(n6668), .Z(n6610) );
  XNOR U65 ( .A(n6958), .B(n7020), .Z(n6962) );
  XNOR U66 ( .A(n7310), .B(n7372), .Z(n7314) );
  XNOR U67 ( .A(n7662), .B(n7724), .Z(n7666) );
  XNOR U68 ( .A(n8014), .B(n8076), .Z(n8018) );
  XNOR U69 ( .A(n8366), .B(n8428), .Z(n8370) );
  XNOR U70 ( .A(n8718), .B(n8780), .Z(n8722) );
  XNOR U71 ( .A(n692), .B(n753), .Z(n696) );
  XNOR U72 ( .A(n6093), .B(n6137), .Z(n6097) );
  XNOR U73 ( .A(n6445), .B(n6489), .Z(n6449) );
  XNOR U74 ( .A(n6797), .B(n6841), .Z(n6801) );
  XNOR U75 ( .A(n7149), .B(n7193), .Z(n7153) );
  XNOR U76 ( .A(n7501), .B(n7545), .Z(n7505) );
  XNOR U77 ( .A(n7853), .B(n7897), .Z(n7857) );
  XNOR U78 ( .A(n8205), .B(n8249), .Z(n8209) );
  XNOR U79 ( .A(n8557), .B(n8601), .Z(n8561) );
  XNOR U80 ( .A(n8909), .B(n8953), .Z(n8913) );
  XNOR U81 ( .A(n9261), .B(n9305), .Z(n9265) );
  XNOR U82 ( .A(n6108), .B(n6134), .Z(n6112) );
  XNOR U83 ( .A(n6460), .B(n6486), .Z(n6464) );
  XNOR U84 ( .A(n6812), .B(n6838), .Z(n6816) );
  XNOR U85 ( .A(n7164), .B(n7190), .Z(n7168) );
  XNOR U86 ( .A(n7516), .B(n7542), .Z(n7520) );
  XNOR U87 ( .A(n7868), .B(n7894), .Z(n7872) );
  XNOR U88 ( .A(n8220), .B(n8246), .Z(n8224) );
  XNOR U89 ( .A(n8572), .B(n8598), .Z(n8576) );
  XNOR U90 ( .A(n8924), .B(n8950), .Z(n8928) );
  XNOR U91 ( .A(n9276), .B(n9302), .Z(n9280) );
  XNOR U92 ( .A(n9628), .B(n9654), .Z(n9632) );
  XNOR U93 ( .A(n9975), .B(n10006), .Z(n9984) );
  ANDN U94 ( .B(n4344), .A(n4345), .Z(n4164) );
  XNOR U95 ( .A(n1684), .B(n1854), .Z(n1689) );
  XNOR U96 ( .A(n15887), .B(n16051), .Z(n15892) );
  XNOR U97 ( .A(n6527), .B(n6685), .Z(n6531) );
  XNOR U98 ( .A(n7055), .B(n7213), .Z(n7059) );
  XNOR U99 ( .A(n5827), .B(n5979), .Z(n5831) );
  XNOR U100 ( .A(n6174), .B(n6331), .Z(n6183) );
  XNOR U101 ( .A(n11144), .B(n11296), .Z(n11148) );
  XNOR U102 ( .A(n11497), .B(n11649), .Z(n11501) );
  XNOR U103 ( .A(n15018), .B(n15170), .Z(n15022) );
  XNOR U104 ( .A(n16448), .B(n16600), .Z(n16452) );
  XNOR U105 ( .A(n16802), .B(n16954), .Z(n16806) );
  XNOR U106 ( .A(n15903), .B(n16048), .Z(n15907) );
  XNOR U107 ( .A(n1705), .B(n1850), .Z(n1709) );
  XNOR U108 ( .A(n6018), .B(n6152), .Z(n6022) );
  XNOR U109 ( .A(n6370), .B(n6504), .Z(n6374) );
  XNOR U110 ( .A(n6717), .B(n6856), .Z(n6726) );
  XNOR U111 ( .A(n7779), .B(n7913), .Z(n7783) );
  XNOR U112 ( .A(n10982), .B(n11116), .Z(n10986) );
  XNOR U113 ( .A(n11336), .B(n11470), .Z(n11340) );
  XNOR U114 ( .A(n11688), .B(n11822), .Z(n11692) );
  XNOR U115 ( .A(n12040), .B(n12174), .Z(n12044) );
  XNOR U116 ( .A(n15033), .B(n15167), .Z(n15037) );
  XNOR U117 ( .A(n16463), .B(n16597), .Z(n16467) );
  XNOR U118 ( .A(n16817), .B(n16951), .Z(n16821) );
  XNOR U119 ( .A(n7432), .B(n7560), .Z(n7436) );
  XNOR U120 ( .A(n15918), .B(n16045), .Z(n15922) );
  XNOR U121 ( .A(n1720), .B(n1847), .Z(n1724) );
  XNOR U122 ( .A(n5857), .B(n5973), .Z(n5861) );
  XNOR U123 ( .A(n6209), .B(n6325), .Z(n6213) );
  XNOR U124 ( .A(n6561), .B(n6677), .Z(n6565) );
  XNOR U125 ( .A(n6913), .B(n7029), .Z(n6917) );
  XNOR U126 ( .A(n7260), .B(n7381), .Z(n7269) );
  XNOR U127 ( .A(n11174), .B(n11290), .Z(n11178) );
  XNOR U128 ( .A(n11527), .B(n11643), .Z(n11531) );
  XNOR U129 ( .A(n11879), .B(n11995), .Z(n11883) );
  XNOR U130 ( .A(n12231), .B(n12347), .Z(n12235) );
  XNOR U131 ( .A(n12583), .B(n12699), .Z(n12587) );
  XNOR U132 ( .A(n15048), .B(n15164), .Z(n15052) );
  XNOR U133 ( .A(n16478), .B(n16594), .Z(n16482) );
  XNOR U134 ( .A(n16832), .B(n16948), .Z(n16836) );
  XNOR U135 ( .A(n15933), .B(n16042), .Z(n15937) );
  XNOR U136 ( .A(n1545), .B(n1665), .Z(n1549) );
  XNOR U137 ( .A(n8156), .B(n8260), .Z(n8160) );
  XNOR U138 ( .A(n6048), .B(n6146), .Z(n6052) );
  XNOR U139 ( .A(n6400), .B(n6498), .Z(n6404) );
  XNOR U140 ( .A(n6752), .B(n6850), .Z(n6756) );
  XNOR U141 ( .A(n7104), .B(n7202), .Z(n7108) );
  XNOR U142 ( .A(n7456), .B(n7554), .Z(n7460) );
  XNOR U143 ( .A(n7803), .B(n7906), .Z(n7812) );
  XNOR U144 ( .A(n9217), .B(n9315), .Z(n9221) );
  XNOR U145 ( .A(n11012), .B(n11110), .Z(n11016) );
  XNOR U146 ( .A(n11366), .B(n11464), .Z(n11370) );
  XNOR U147 ( .A(n11718), .B(n11816), .Z(n11722) );
  XNOR U148 ( .A(n12070), .B(n12168), .Z(n12074) );
  XNOR U149 ( .A(n12422), .B(n12520), .Z(n12426) );
  XNOR U150 ( .A(n12774), .B(n12872), .Z(n12778) );
  XNOR U151 ( .A(n13126), .B(n13224), .Z(n13130) );
  XNOR U152 ( .A(n15063), .B(n15161), .Z(n15067) );
  XNOR U153 ( .A(n16493), .B(n16591), .Z(n16497) );
  XNOR U154 ( .A(n16847), .B(n16945), .Z(n16851) );
  XNOR U155 ( .A(n1199), .B(n1301), .Z(n1203) );
  XNOR U156 ( .A(n15948), .B(n16039), .Z(n15952) );
  XNOR U157 ( .A(n823), .B(n943), .Z(n827) );
  XNOR U158 ( .A(n1560), .B(n1662), .Z(n1564) );
  XNOR U159 ( .A(n1394), .B(n1479), .Z(n1398) );
  XNOR U160 ( .A(n5887), .B(n5967), .Z(n5891) );
  XNOR U161 ( .A(n6239), .B(n6319), .Z(n6243) );
  XNOR U162 ( .A(n6591), .B(n6671), .Z(n6595) );
  XNOR U163 ( .A(n6943), .B(n7023), .Z(n6947) );
  XNOR U164 ( .A(n7295), .B(n7375), .Z(n7299) );
  XNOR U165 ( .A(n7647), .B(n7727), .Z(n7651) );
  XNOR U166 ( .A(n7999), .B(n8079), .Z(n8003) );
  XNOR U167 ( .A(n8346), .B(n8431), .Z(n8355) );
  XNOR U168 ( .A(n11204), .B(n11284), .Z(n11208) );
  XNOR U169 ( .A(n11557), .B(n11637), .Z(n11561) );
  XNOR U170 ( .A(n11909), .B(n11989), .Z(n11913) );
  XNOR U171 ( .A(n12261), .B(n12341), .Z(n12265) );
  XNOR U172 ( .A(n12613), .B(n12693), .Z(n12617) );
  XNOR U173 ( .A(n12965), .B(n13045), .Z(n12969) );
  XNOR U174 ( .A(n13317), .B(n13397), .Z(n13321) );
  XNOR U175 ( .A(n13669), .B(n13749), .Z(n13673) );
  XNOR U176 ( .A(n16508), .B(n16588), .Z(n16512) );
  XNOR U177 ( .A(n16862), .B(n16942), .Z(n16866) );
  XNOR U178 ( .A(n1219), .B(n1297), .Z(n1223) );
  XNOR U179 ( .A(n9413), .B(n9487), .Z(n9417) );
  XNOR U180 ( .A(n15963), .B(n16036), .Z(n15967) );
  XNOR U181 ( .A(n667), .B(n758), .Z(n671) );
  XNOR U182 ( .A(n1048), .B(n1115), .Z(n1052) );
  XNOR U183 ( .A(n3214), .B(n3280), .Z(n3218) );
  XNOR U184 ( .A(n3574), .B(n3640), .Z(n3578) );
  XNOR U185 ( .A(n6078), .B(n6140), .Z(n6082) );
  XNOR U186 ( .A(n6430), .B(n6492), .Z(n6434) );
  XNOR U187 ( .A(n6782), .B(n6844), .Z(n6786) );
  XNOR U188 ( .A(n7134), .B(n7196), .Z(n7138) );
  XNOR U189 ( .A(n7486), .B(n7548), .Z(n7490) );
  XNOR U190 ( .A(n7838), .B(n7900), .Z(n7842) );
  XNOR U191 ( .A(n8190), .B(n8252), .Z(n8194) );
  XNOR U192 ( .A(n8542), .B(n8604), .Z(n8546) );
  XNOR U193 ( .A(n8889), .B(n8956), .Z(n8898) );
  XNOR U194 ( .A(n11042), .B(n11104), .Z(n11046) );
  XNOR U195 ( .A(n11396), .B(n11458), .Z(n11400) );
  XNOR U196 ( .A(n11748), .B(n11810), .Z(n11752) );
  XNOR U197 ( .A(n12100), .B(n12162), .Z(n12104) );
  XNOR U198 ( .A(n12452), .B(n12514), .Z(n12456) );
  XNOR U199 ( .A(n12804), .B(n12866), .Z(n12808) );
  XNOR U200 ( .A(n13156), .B(n13218), .Z(n13160) );
  XNOR U201 ( .A(n13508), .B(n13570), .Z(n13512) );
  XNOR U202 ( .A(n13860), .B(n13922), .Z(n13864) );
  XNOR U203 ( .A(n14212), .B(n14274), .Z(n14216) );
  XNOR U204 ( .A(n16523), .B(n16585), .Z(n16527) );
  XNOR U205 ( .A(n16877), .B(n16939), .Z(n16881) );
  XNOR U206 ( .A(n15978), .B(n16033), .Z(n15982) );
  XNOR U207 ( .A(n873), .B(n933), .Z(n877) );
  XNOR U208 ( .A(n4304), .B(n4358), .Z(n4308) );
  XNOR U209 ( .A(n10137), .B(n10187), .Z(n10141) );
  XNOR U210 ( .A(n5917), .B(n5961), .Z(n5921) );
  XNOR U211 ( .A(n6269), .B(n6313), .Z(n6273) );
  XNOR U212 ( .A(n6621), .B(n6665), .Z(n6625) );
  XNOR U213 ( .A(n6973), .B(n7017), .Z(n6977) );
  XNOR U214 ( .A(n7325), .B(n7369), .Z(n7329) );
  XNOR U215 ( .A(n7677), .B(n7721), .Z(n7681) );
  XNOR U216 ( .A(n8029), .B(n8073), .Z(n8033) );
  XNOR U217 ( .A(n8381), .B(n8425), .Z(n8385) );
  XNOR U218 ( .A(n8733), .B(n8777), .Z(n8737) );
  XNOR U219 ( .A(n9085), .B(n9129), .Z(n9089) );
  XNOR U220 ( .A(n9432), .B(n9481), .Z(n9441) );
  XNOR U221 ( .A(n9966), .B(n10010), .Z(n9970) );
  XNOR U222 ( .A(n11234), .B(n11278), .Z(n11238) );
  XNOR U223 ( .A(n11587), .B(n11631), .Z(n11591) );
  XNOR U224 ( .A(n11939), .B(n11983), .Z(n11943) );
  XNOR U225 ( .A(n12291), .B(n12335), .Z(n12295) );
  XNOR U226 ( .A(n12643), .B(n12687), .Z(n12647) );
  XNOR U227 ( .A(n12995), .B(n13039), .Z(n12999) );
  XNOR U228 ( .A(n13347), .B(n13391), .Z(n13351) );
  XNOR U229 ( .A(n13699), .B(n13743), .Z(n13703) );
  XNOR U230 ( .A(n14051), .B(n14095), .Z(n14055) );
  XNOR U231 ( .A(n14403), .B(n14447), .Z(n14407) );
  XNOR U232 ( .A(n14755), .B(n14799), .Z(n14759) );
  XNOR U233 ( .A(n16538), .B(n16582), .Z(n16542) );
  XNOR U234 ( .A(n16892), .B(n16936), .Z(n16896) );
  XNOR U235 ( .A(n15817), .B(n15855), .Z(n15821) );
  XNOR U236 ( .A(n3059), .B(n3095), .Z(n3063) );
  XNOR U237 ( .A(n3419), .B(n3455), .Z(n3423) );
  XNOR U238 ( .A(n3779), .B(n3815), .Z(n3783) );
  XNOR U239 ( .A(n4319), .B(n4355), .Z(n4323) );
  XNOR U240 ( .A(n10504), .B(n10536), .Z(n10508) );
  XNOR U241 ( .A(n5932), .B(n5958), .Z(n5936) );
  XNOR U242 ( .A(n6284), .B(n6310), .Z(n6288) );
  XNOR U243 ( .A(n6636), .B(n6662), .Z(n6640) );
  XNOR U244 ( .A(n6988), .B(n7014), .Z(n6992) );
  XNOR U245 ( .A(n7340), .B(n7366), .Z(n7344) );
  XNOR U246 ( .A(n7692), .B(n7718), .Z(n7696) );
  XNOR U247 ( .A(n8044), .B(n8070), .Z(n8048) );
  XNOR U248 ( .A(n8396), .B(n8422), .Z(n8400) );
  XNOR U249 ( .A(n8748), .B(n8774), .Z(n8752) );
  XNOR U250 ( .A(n9100), .B(n9126), .Z(n9104) );
  XNOR U251 ( .A(n9452), .B(n9478), .Z(n9456) );
  XNOR U252 ( .A(n9804), .B(n9830), .Z(n9808) );
  XNOR U253 ( .A(n11072), .B(n11098), .Z(n11076) );
  XNOR U254 ( .A(n11426), .B(n11452), .Z(n11430) );
  XNOR U255 ( .A(n11778), .B(n11804), .Z(n11782) );
  XNOR U256 ( .A(n12130), .B(n12156), .Z(n12134) );
  XNOR U257 ( .A(n12482), .B(n12508), .Z(n12486) );
  XNOR U258 ( .A(n12834), .B(n12860), .Z(n12838) );
  XNOR U259 ( .A(n13186), .B(n13212), .Z(n13190) );
  XNOR U260 ( .A(n13538), .B(n13564), .Z(n13542) );
  XNOR U261 ( .A(n13890), .B(n13916), .Z(n13894) );
  XNOR U262 ( .A(n14242), .B(n14268), .Z(n14246) );
  XNOR U263 ( .A(n14594), .B(n14620), .Z(n14598) );
  XNOR U264 ( .A(n14946), .B(n14972), .Z(n14950) );
  XNOR U265 ( .A(n15298), .B(n15324), .Z(n15302) );
  XNOR U266 ( .A(n16553), .B(n16579), .Z(n16557) );
  XNOR U267 ( .A(n16907), .B(n16933), .Z(n16911) );
  XNOR U268 ( .A(n5584), .B(n5603), .Z(n5588) );
  XNOR U269 ( .A(n10156), .B(n10181), .Z(n10165) );
  ANDN U270 ( .B(n3624), .A(n3625), .Z(n3444) );
  ANDN U271 ( .B(n4524), .A(n4525), .Z(n4344) );
  XNOR U272 ( .A(n4028), .B(n4197), .Z(n4033) );
  XNOR U273 ( .A(n6697), .B(n6862), .Z(n6702) );
  XNOR U274 ( .A(n7401), .B(n7566), .Z(n7406) );
  XNOR U275 ( .A(n9513), .B(n9678), .Z(n9518) );
  XNOR U276 ( .A(n15183), .B(n15348), .Z(n15188) );
  XNOR U277 ( .A(n15535), .B(n15700), .Z(n15540) );
  XNOR U278 ( .A(n2051), .B(n2214), .Z(n2055) );
  XNOR U279 ( .A(n4394), .B(n4556), .Z(n4398) );
  XNOR U280 ( .A(n7759), .B(n7917), .Z(n7763) );
  XNOR U281 ( .A(n8111), .B(n8269), .Z(n8115) );
  XNOR U282 ( .A(n9871), .B(n10029), .Z(n9875) );
  XNOR U283 ( .A(n13077), .B(n13235), .Z(n13081) );
  XNOR U284 ( .A(n13429), .B(n13587), .Z(n13433) );
  XNOR U285 ( .A(n18026), .B(n18184), .Z(n18030) );
  XNOR U286 ( .A(n17690), .B(n17848), .Z(n17694) );
  XNOR U287 ( .A(n17330), .B(n17486), .Z(n17324) );
  XNOR U288 ( .A(n1876), .B(n2032), .Z(n1880) );
  XNOR U289 ( .A(n2598), .B(n2754), .Z(n2602) );
  XNOR U290 ( .A(n2959), .B(n3115), .Z(n2963) );
  XNOR U291 ( .A(n3319), .B(n3475), .Z(n3323) );
  XNOR U292 ( .A(n3679), .B(n3835), .Z(n3683) );
  XNOR U293 ( .A(n4759), .B(n4915), .Z(n4763) );
  XNOR U294 ( .A(n5656), .B(n5477), .Z(n5479) );
  XNOR U295 ( .A(n8468), .B(n8620), .Z(n8472) );
  XNOR U296 ( .A(n8820), .B(n8972), .Z(n8824) );
  XNOR U297 ( .A(n9172), .B(n9324), .Z(n9176) );
  XNOR U298 ( .A(n10228), .B(n10380), .Z(n10232) );
  XNOR U299 ( .A(n10580), .B(n10734), .Z(n10584) );
  XNOR U300 ( .A(n10967), .B(n11119), .Z(n10971) );
  XNOR U301 ( .A(n11321), .B(n11473), .Z(n11325) );
  XNOR U302 ( .A(n11855), .B(n11676), .Z(n11678) );
  XNOR U303 ( .A(n11854), .B(n12002), .Z(n11849) );
  XNOR U304 ( .A(n12202), .B(n12354), .Z(n12206) );
  XNOR U305 ( .A(n12554), .B(n12706), .Z(n12558) );
  XNOR U306 ( .A(n12906), .B(n13058), .Z(n12910) );
  XNOR U307 ( .A(n13962), .B(n14114), .Z(n13966) );
  XNOR U308 ( .A(n14314), .B(n14466), .Z(n14318) );
  XNOR U309 ( .A(n14666), .B(n14818), .Z(n14670) );
  XNOR U310 ( .A(n16073), .B(n16224), .Z(n16077) );
  XNOR U311 ( .A(n16625), .B(n16777), .Z(n16629) );
  XNOR U312 ( .A(n16978), .B(n17130), .Z(n16982) );
  XNOR U313 ( .A(n4044), .B(n4194), .Z(n4048) );
  XNOR U314 ( .A(n5832), .B(n5978), .Z(n5836) );
  XNOR U315 ( .A(n6184), .B(n6330), .Z(n6188) );
  XNOR U316 ( .A(n6889), .B(n7035), .Z(n6893) );
  XNOR U317 ( .A(n7417), .B(n7563), .Z(n7421) );
  XNOR U318 ( .A(n9529), .B(n9675), .Z(n9533) );
  XNOR U319 ( .A(n15199), .B(n15345), .Z(n15203) );
  XNOR U320 ( .A(n15551), .B(n15697), .Z(n15555) );
  XNOR U321 ( .A(n1515), .B(n1671), .Z(n1519) );
  XNOR U322 ( .A(n2427), .B(n2572), .Z(n2431) );
  XNOR U323 ( .A(n4409), .B(n4553), .Z(n4413) );
  XNOR U324 ( .A(n8126), .B(n8266), .Z(n8130) );
  XNOR U325 ( .A(n9886), .B(n10026), .Z(n9890) );
  XNOR U326 ( .A(n13444), .B(n13584), .Z(n13448) );
  XNOR U327 ( .A(n13796), .B(n13936), .Z(n13800) );
  XNOR U328 ( .A(n18353), .B(n18493), .Z(n18357) );
  XNOR U329 ( .A(n18041), .B(n18181), .Z(n18045) );
  XNOR U330 ( .A(n17705), .B(n17845), .Z(n17709) );
  XNOR U331 ( .A(n17340), .B(n17483), .Z(n17344) );
  XNOR U332 ( .A(n1891), .B(n2029), .Z(n1895) );
  XNOR U333 ( .A(n2252), .B(n2390), .Z(n2256) );
  XNOR U334 ( .A(n2974), .B(n3112), .Z(n2978) );
  XNOR U335 ( .A(n3334), .B(n3472), .Z(n3338) );
  XNOR U336 ( .A(n3694), .B(n3832), .Z(n3698) );
  XNOR U337 ( .A(n4774), .B(n4912), .Z(n4778) );
  XNOR U338 ( .A(n5671), .B(n5492), .Z(n5494) );
  XNOR U339 ( .A(n8483), .B(n8617), .Z(n8487) );
  XNOR U340 ( .A(n8835), .B(n8969), .Z(n8839) );
  XNOR U341 ( .A(n9187), .B(n9321), .Z(n9191) );
  XNOR U342 ( .A(n10243), .B(n10377), .Z(n10247) );
  XNOR U343 ( .A(n10595), .B(n10731), .Z(n10599) );
  XNOR U344 ( .A(n11159), .B(n11293), .Z(n11163) );
  XNOR U345 ( .A(n11512), .B(n11646), .Z(n11516) );
  XNOR U346 ( .A(n11864), .B(n11998), .Z(n11868) );
  XNOR U347 ( .A(n12211), .B(n12350), .Z(n12220) );
  XNOR U348 ( .A(n12569), .B(n12703), .Z(n12577) );
  XNOR U349 ( .A(n12921), .B(n13055), .Z(n12925) );
  XNOR U350 ( .A(n13273), .B(n13407), .Z(n13277) );
  XNOR U351 ( .A(n14329), .B(n14463), .Z(n14333) );
  XNOR U352 ( .A(n14681), .B(n14815), .Z(n14685) );
  XNOR U353 ( .A(n16088), .B(n16221), .Z(n16092) );
  XNOR U354 ( .A(n16640), .B(n16774), .Z(n16644) );
  XNOR U355 ( .A(n16993), .B(n17127), .Z(n16997) );
  XNOR U356 ( .A(n1715), .B(n1848), .Z(n1719) );
  XNOR U357 ( .A(n4059), .B(n4191), .Z(n4063) );
  XNOR U358 ( .A(n5847), .B(n5975), .Z(n5851) );
  XNOR U359 ( .A(n6199), .B(n6327), .Z(n6203) );
  XNOR U360 ( .A(n6551), .B(n6679), .Z(n6555) );
  XNOR U361 ( .A(n6898), .B(n7031), .Z(n6907) );
  XNOR U362 ( .A(n7608), .B(n7736), .Z(n7612) );
  XNOR U363 ( .A(n7960), .B(n8088), .Z(n7964) );
  XNOR U364 ( .A(n9544), .B(n9672), .Z(n9548) );
  XNOR U365 ( .A(n15214), .B(n15342), .Z(n15218) );
  XNOR U366 ( .A(n15566), .B(n15694), .Z(n15570) );
  XNOR U367 ( .A(n1339), .B(n1490), .Z(n1343) );
  XNOR U368 ( .A(n2803), .B(n2930), .Z(n2807) );
  XNOR U369 ( .A(n4424), .B(n4550), .Z(n4428) );
  XNOR U370 ( .A(n8317), .B(n8439), .Z(n8321) );
  XNOR U371 ( .A(n9901), .B(n10023), .Z(n9905) );
  XNOR U372 ( .A(n13811), .B(n13933), .Z(n13815) );
  XNOR U373 ( .A(n14163), .B(n14285), .Z(n14167) );
  XNOR U374 ( .A(n18920), .B(n19042), .Z(n18924) );
  XNOR U375 ( .A(n18656), .B(n18778), .Z(n18660) );
  XNOR U376 ( .A(n18368), .B(n18490), .Z(n18372) );
  XNOR U377 ( .A(n18056), .B(n18178), .Z(n18060) );
  XNOR U378 ( .A(n17720), .B(n17842), .Z(n17724) );
  XNOR U379 ( .A(n17355), .B(n17480), .Z(n17359) );
  XNOR U380 ( .A(n2267), .B(n2387), .Z(n2271) );
  XNOR U381 ( .A(n2628), .B(n2748), .Z(n2632) );
  XNOR U382 ( .A(n3349), .B(n3469), .Z(n3353) );
  XNOR U383 ( .A(n3709), .B(n3829), .Z(n3713) );
  XNOR U384 ( .A(n4789), .B(n4909), .Z(n4793) );
  XNOR U385 ( .A(n5686), .B(n5507), .Z(n5509) );
  XNOR U386 ( .A(n5863), .B(n5683), .Z(n5685) );
  XNOR U387 ( .A(n8850), .B(n8966), .Z(n8854) );
  XNOR U388 ( .A(n9202), .B(n9318), .Z(n9206) );
  XNOR U389 ( .A(n10258), .B(n10374), .Z(n10262) );
  XNOR U390 ( .A(n10610), .B(n10728), .Z(n10614) );
  XNOR U391 ( .A(n10997), .B(n11113), .Z(n11001) );
  XNOR U392 ( .A(n11351), .B(n11467), .Z(n11355) );
  XNOR U393 ( .A(n11703), .B(n11819), .Z(n11707) );
  XNOR U394 ( .A(n12055), .B(n12171), .Z(n12059) );
  XNOR U395 ( .A(n12407), .B(n12523), .Z(n12411) );
  XNOR U396 ( .A(n12941), .B(n12762), .Z(n12764) );
  XNOR U397 ( .A(n12940), .B(n13052), .Z(n12935) );
  XNOR U398 ( .A(n13288), .B(n13404), .Z(n13292) );
  XNOR U399 ( .A(n13640), .B(n13756), .Z(n13644) );
  XNOR U400 ( .A(n14696), .B(n14812), .Z(n14700) );
  XNOR U401 ( .A(n16103), .B(n16218), .Z(n16107) );
  XNOR U402 ( .A(n16655), .B(n16771), .Z(n16659) );
  XNOR U403 ( .A(n17008), .B(n17124), .Z(n17012) );
  XNOR U404 ( .A(n1730), .B(n1845), .Z(n1734) );
  XNOR U405 ( .A(n4074), .B(n4188), .Z(n4078) );
  XNOR U406 ( .A(n6038), .B(n6148), .Z(n6042) );
  XNOR U407 ( .A(n6390), .B(n6500), .Z(n6394) );
  XNOR U408 ( .A(n6742), .B(n6852), .Z(n6746) );
  XNOR U409 ( .A(n7094), .B(n7204), .Z(n7098) );
  XNOR U410 ( .A(n7441), .B(n7556), .Z(n7450) );
  XNOR U411 ( .A(n7975), .B(n8085), .Z(n7979) );
  XNOR U412 ( .A(n9559), .B(n9669), .Z(n9563) );
  XNOR U413 ( .A(n15229), .B(n15339), .Z(n15233) );
  XNOR U414 ( .A(n15581), .B(n15691), .Z(n15585) );
  XNOR U415 ( .A(n1354), .B(n1487), .Z(n1358) );
  XNOR U416 ( .A(n973), .B(n1130), .Z(n977) );
  XNOR U417 ( .A(n2096), .B(n2205), .Z(n2100) );
  XNOR U418 ( .A(n3179), .B(n3287), .Z(n3183) );
  XNOR U419 ( .A(n4439), .B(n4547), .Z(n4443) );
  XNOR U420 ( .A(n8332), .B(n8436), .Z(n8336) );
  XNOR U421 ( .A(n8684), .B(n8788), .Z(n8688) );
  XNOR U422 ( .A(n9916), .B(n10020), .Z(n9920) );
  XNOR U423 ( .A(n14178), .B(n14282), .Z(n14182) );
  XNOR U424 ( .A(n14530), .B(n14634), .Z(n14534) );
  XNOR U425 ( .A(n19175), .B(n19279), .Z(n19179) );
  XNOR U426 ( .A(n18935), .B(n19039), .Z(n18939) );
  XNOR U427 ( .A(n18671), .B(n18775), .Z(n18675) );
  XNOR U428 ( .A(n18383), .B(n18487), .Z(n18387) );
  XNOR U429 ( .A(n18071), .B(n18175), .Z(n18075) );
  XNOR U430 ( .A(n17735), .B(n17839), .Z(n17739) );
  XNOR U431 ( .A(n17370), .B(n17477), .Z(n17374) );
  XNOR U432 ( .A(n1194), .B(n1302), .Z(n1198) );
  XNOR U433 ( .A(n2643), .B(n2745), .Z(n2647) );
  XNOR U434 ( .A(n3004), .B(n3106), .Z(n3008) );
  XNOR U435 ( .A(n3724), .B(n3826), .Z(n3728) );
  XNOR U436 ( .A(n4804), .B(n4906), .Z(n4808) );
  XNOR U437 ( .A(n5701), .B(n5522), .Z(n5524) );
  XNOR U438 ( .A(n5878), .B(n5698), .Z(n5700) );
  XNOR U439 ( .A(n10273), .B(n10371), .Z(n10277) );
  XNOR U440 ( .A(n10625), .B(n10725), .Z(n10629) );
  XNOR U441 ( .A(n11189), .B(n11287), .Z(n11193) );
  XNOR U442 ( .A(n11542), .B(n11640), .Z(n11546) );
  XNOR U443 ( .A(n11894), .B(n11992), .Z(n11898) );
  XNOR U444 ( .A(n12246), .B(n12344), .Z(n12250) );
  XNOR U445 ( .A(n12598), .B(n12696), .Z(n12602) );
  XNOR U446 ( .A(n12950), .B(n13048), .Z(n12954) );
  XNOR U447 ( .A(n13297), .B(n13400), .Z(n13306) );
  XNOR U448 ( .A(n13655), .B(n13753), .Z(n13663) );
  XNOR U449 ( .A(n14007), .B(n14105), .Z(n14011) );
  XNOR U450 ( .A(n16118), .B(n16215), .Z(n16122) );
  XNOR U451 ( .A(n16670), .B(n16768), .Z(n16674) );
  XNOR U452 ( .A(n17023), .B(n17121), .Z(n17027) );
  XNOR U453 ( .A(n4089), .B(n4185), .Z(n4093) );
  XNOR U454 ( .A(n6053), .B(n6145), .Z(n6057) );
  XNOR U455 ( .A(n6405), .B(n6497), .Z(n6409) );
  XNOR U456 ( .A(n6757), .B(n6849), .Z(n6761) );
  XNOR U457 ( .A(n7109), .B(n7201), .Z(n7113) );
  XNOR U458 ( .A(n7461), .B(n7553), .Z(n7465) );
  XNOR U459 ( .A(n7813), .B(n7905), .Z(n7817) );
  XNOR U460 ( .A(n9222), .B(n9314), .Z(n9226) );
  XNOR U461 ( .A(n9574), .B(n9666), .Z(n9578) );
  XNOR U462 ( .A(n15244), .B(n15336), .Z(n15248) );
  XNOR U463 ( .A(n15596), .B(n15688), .Z(n15600) );
  XNOR U464 ( .A(n1179), .B(n1305), .Z(n1183) );
  XNOR U465 ( .A(n798), .B(n948), .Z(n802) );
  XNOR U466 ( .A(n1750), .B(n1841), .Z(n1754) );
  XNOR U467 ( .A(n2111), .B(n2202), .Z(n2115) );
  XNOR U468 ( .A(n2472), .B(n2563), .Z(n2476) );
  XNOR U469 ( .A(n3554), .B(n3644), .Z(n3558) );
  XNOR U470 ( .A(n4454), .B(n4544), .Z(n4458) );
  XNOR U471 ( .A(n8699), .B(n8785), .Z(n8703) );
  XNOR U472 ( .A(n9051), .B(n9137), .Z(n9055) );
  XNOR U473 ( .A(n9931), .B(n10017), .Z(n9935) );
  XNOR U474 ( .A(n14545), .B(n14631), .Z(n14549) );
  XNOR U475 ( .A(n14897), .B(n14983), .Z(n14901) );
  XNOR U476 ( .A(n19598), .B(n19684), .Z(n19602) );
  XNOR U477 ( .A(n19406), .B(n19492), .Z(n19410) );
  XNOR U478 ( .A(n19190), .B(n19276), .Z(n19194) );
  XNOR U479 ( .A(n18950), .B(n19036), .Z(n18954) );
  XNOR U480 ( .A(n18686), .B(n18772), .Z(n18690) );
  XNOR U481 ( .A(n18398), .B(n18484), .Z(n18402) );
  XNOR U482 ( .A(n18086), .B(n18172), .Z(n18090) );
  XNOR U483 ( .A(n17750), .B(n17836), .Z(n17754) );
  XNOR U484 ( .A(n17385), .B(n17474), .Z(n17389) );
  XNOR U485 ( .A(n1209), .B(n1299), .Z(n1213) );
  XNOR U486 ( .A(n1033), .B(n1118), .Z(n1037) );
  XNOR U487 ( .A(n1575), .B(n1659), .Z(n1579) );
  XNOR U488 ( .A(n3019), .B(n3103), .Z(n3023) );
  XNOR U489 ( .A(n3379), .B(n3463), .Z(n3383) );
  XNOR U490 ( .A(n4819), .B(n4903), .Z(n4823) );
  XNOR U491 ( .A(n5716), .B(n5537), .Z(n5539) );
  XNOR U492 ( .A(n8532), .B(n8608), .Z(n8527) );
  XNOR U493 ( .A(n10288), .B(n10368), .Z(n10292) );
  XNOR U494 ( .A(n10640), .B(n10722), .Z(n10644) );
  XNOR U495 ( .A(n11027), .B(n11107), .Z(n11031) );
  XNOR U496 ( .A(n11381), .B(n11461), .Z(n11385) );
  XNOR U497 ( .A(n11733), .B(n11813), .Z(n11737) );
  XNOR U498 ( .A(n12085), .B(n12165), .Z(n12089) );
  XNOR U499 ( .A(n12437), .B(n12517), .Z(n12441) );
  XNOR U500 ( .A(n12789), .B(n12869), .Z(n12793) );
  XNOR U501 ( .A(n13141), .B(n13221), .Z(n13145) );
  XNOR U502 ( .A(n13493), .B(n13573), .Z(n13497) );
  XNOR U503 ( .A(n14027), .B(n13848), .Z(n13850) );
  XNOR U504 ( .A(n14026), .B(n14102), .Z(n14021) );
  XNOR U505 ( .A(n14374), .B(n14454), .Z(n14378) );
  XNOR U506 ( .A(n16133), .B(n16212), .Z(n16137) );
  XNOR U507 ( .A(n16685), .B(n16765), .Z(n16689) );
  XNOR U508 ( .A(n17038), .B(n17118), .Z(n17042) );
  XNOR U509 ( .A(n833), .B(n941), .Z(n837) );
  XNOR U510 ( .A(n4104), .B(n4182), .Z(n4108) );
  XNOR U511 ( .A(n5892), .B(n5966), .Z(n5896) );
  XNOR U512 ( .A(n6244), .B(n6318), .Z(n6248) );
  XNOR U513 ( .A(n6596), .B(n6670), .Z(n6600) );
  XNOR U514 ( .A(n6948), .B(n7022), .Z(n6952) );
  XNOR U515 ( .A(n7300), .B(n7374), .Z(n7304) );
  XNOR U516 ( .A(n7652), .B(n7726), .Z(n7656) );
  XNOR U517 ( .A(n8004), .B(n8078), .Z(n8008) );
  XNOR U518 ( .A(n8356), .B(n8430), .Z(n8360) );
  XNOR U519 ( .A(n9589), .B(n9663), .Z(n9593) );
  XNOR U520 ( .A(n15611), .B(n15685), .Z(n15615) );
  XNOR U521 ( .A(n622), .B(n767), .Z(n626) );
  XNOR U522 ( .A(n2126), .B(n2199), .Z(n2130) );
  XNOR U523 ( .A(n2487), .B(n2560), .Z(n2491) );
  XNOR U524 ( .A(n2848), .B(n2921), .Z(n2852) );
  XNOR U525 ( .A(n3929), .B(n4001), .Z(n3933) );
  XNOR U526 ( .A(n4469), .B(n4541), .Z(n4473) );
  XNOR U527 ( .A(n9066), .B(n9134), .Z(n9074) );
  XNOR U528 ( .A(n9946), .B(n10014), .Z(n9950) );
  XNOR U529 ( .A(n14912), .B(n14980), .Z(n14916) );
  XNOR U530 ( .A(n15440), .B(n15508), .Z(n15444) );
  XNOR U531 ( .A(n19781), .B(n19849), .Z(n19785) );
  XNOR U532 ( .A(n19613), .B(n19681), .Z(n19617) );
  XNOR U533 ( .A(n19421), .B(n19489), .Z(n19425) );
  XNOR U534 ( .A(n19205), .B(n19273), .Z(n19209) );
  XNOR U535 ( .A(n18965), .B(n19033), .Z(n18969) );
  XNOR U536 ( .A(n18701), .B(n18769), .Z(n18705) );
  XNOR U537 ( .A(n18413), .B(n18481), .Z(n18417) );
  XNOR U538 ( .A(n18101), .B(n18169), .Z(n18105) );
  XNOR U539 ( .A(n17765), .B(n17833), .Z(n17769) );
  XNOR U540 ( .A(n17400), .B(n17471), .Z(n17404) );
  XNOR U541 ( .A(n672), .B(n757), .Z(n676) );
  XNOR U542 ( .A(n1409), .B(n1476), .Z(n1413) );
  XNOR U543 ( .A(n1770), .B(n1837), .Z(n1774) );
  XNOR U544 ( .A(n4834), .B(n4900), .Z(n4838) );
  XNOR U545 ( .A(n5731), .B(n5552), .Z(n5554) );
  XNOR U546 ( .A(n5908), .B(n5728), .Z(n5730) );
  XNOR U547 ( .A(n10303), .B(n10365), .Z(n10307) );
  XNOR U548 ( .A(n10655), .B(n10719), .Z(n10659) );
  XNOR U549 ( .A(n11219), .B(n11281), .Z(n11223) );
  XNOR U550 ( .A(n11572), .B(n11634), .Z(n11576) );
  XNOR U551 ( .A(n11924), .B(n11986), .Z(n11928) );
  XNOR U552 ( .A(n12276), .B(n12338), .Z(n12280) );
  XNOR U553 ( .A(n12628), .B(n12690), .Z(n12632) );
  XNOR U554 ( .A(n12980), .B(n13042), .Z(n12984) );
  XNOR U555 ( .A(n13332), .B(n13394), .Z(n13336) );
  XNOR U556 ( .A(n13684), .B(n13746), .Z(n13688) );
  XNOR U557 ( .A(n14036), .B(n14098), .Z(n14040) );
  XNOR U558 ( .A(n14383), .B(n14450), .Z(n14392) );
  XNOR U559 ( .A(n14741), .B(n14803), .Z(n14749) );
  XNOR U560 ( .A(n16148), .B(n16209), .Z(n16152) );
  XNOR U561 ( .A(n16700), .B(n16762), .Z(n16704) );
  XNOR U562 ( .A(n17053), .B(n17115), .Z(n17057) );
  XNOR U563 ( .A(n868), .B(n934), .Z(n872) );
  XNOR U564 ( .A(n6083), .B(n6139), .Z(n6087) );
  XNOR U565 ( .A(n6435), .B(n6491), .Z(n6439) );
  XNOR U566 ( .A(n6787), .B(n6843), .Z(n6791) );
  XNOR U567 ( .A(n7139), .B(n7195), .Z(n7143) );
  XNOR U568 ( .A(n7491), .B(n7547), .Z(n7495) );
  XNOR U569 ( .A(n7843), .B(n7899), .Z(n7847) );
  XNOR U570 ( .A(n8195), .B(n8251), .Z(n8199) );
  XNOR U571 ( .A(n8547), .B(n8603), .Z(n8551) );
  XNOR U572 ( .A(n8899), .B(n8955), .Z(n8903) );
  XNOR U573 ( .A(n2502), .B(n2557), .Z(n2506) );
  XNOR U574 ( .A(n2863), .B(n2918), .Z(n2867) );
  XNOR U575 ( .A(n3224), .B(n3278), .Z(n3228) );
  XNOR U576 ( .A(n3764), .B(n3818), .Z(n3768) );
  XNOR U577 ( .A(n4124), .B(n4178), .Z(n4128) );
  XNOR U578 ( .A(n4484), .B(n4538), .Z(n4488) );
  XNOR U579 ( .A(n15279), .B(n15329), .Z(n15283) );
  XNOR U580 ( .A(n20060), .B(n20110), .Z(n20064) );
  XNOR U581 ( .A(n19940), .B(n19990), .Z(n19944) );
  XNOR U582 ( .A(n19796), .B(n19846), .Z(n19800) );
  XNOR U583 ( .A(n19628), .B(n19678), .Z(n19632) );
  XNOR U584 ( .A(n19436), .B(n19486), .Z(n19440) );
  XNOR U585 ( .A(n19220), .B(n19270), .Z(n19224) );
  XNOR U586 ( .A(n18980), .B(n19030), .Z(n18984) );
  XNOR U587 ( .A(n18716), .B(n18766), .Z(n18720) );
  XNOR U588 ( .A(n18428), .B(n18478), .Z(n18432) );
  XNOR U589 ( .A(n18116), .B(n18166), .Z(n18120) );
  XNOR U590 ( .A(n17780), .B(n17830), .Z(n17784) );
  XNOR U591 ( .A(n17415), .B(n17468), .Z(n17419) );
  XNOR U592 ( .A(n522), .B(n570), .Z(n526) );
  XNOR U593 ( .A(n883), .B(n931), .Z(n887) );
  XNOR U594 ( .A(n1244), .B(n1292), .Z(n1248) );
  XNOR U595 ( .A(n1605), .B(n1653), .Z(n1609) );
  XNOR U596 ( .A(n1966), .B(n2014), .Z(n1970) );
  XNOR U597 ( .A(n2327), .B(n2375), .Z(n2331) );
  XNOR U598 ( .A(n4849), .B(n4897), .Z(n4853) );
  XNOR U599 ( .A(n5746), .B(n5567), .Z(n5569) );
  XNOR U600 ( .A(n5923), .B(n5743), .Z(n5745) );
  XNOR U601 ( .A(n10142), .B(n10186), .Z(n10146) );
  XNOR U602 ( .A(n10670), .B(n10716), .Z(n10674) );
  XNOR U603 ( .A(n11057), .B(n11101), .Z(n11061) );
  XNOR U604 ( .A(n11411), .B(n11455), .Z(n11415) );
  XNOR U605 ( .A(n11763), .B(n11807), .Z(n11767) );
  XNOR U606 ( .A(n12115), .B(n12159), .Z(n12119) );
  XNOR U607 ( .A(n12467), .B(n12511), .Z(n12471) );
  XNOR U608 ( .A(n12819), .B(n12863), .Z(n12823) );
  XNOR U609 ( .A(n13171), .B(n13215), .Z(n13175) );
  XNOR U610 ( .A(n13523), .B(n13567), .Z(n13527) );
  XNOR U611 ( .A(n13875), .B(n13919), .Z(n13879) );
  XNOR U612 ( .A(n14227), .B(n14271), .Z(n14231) );
  XNOR U613 ( .A(n14579), .B(n14623), .Z(n14583) );
  XNOR U614 ( .A(n15113), .B(n14934), .Z(n14936) );
  XNOR U615 ( .A(n15112), .B(n15152), .Z(n15107) );
  XNOR U616 ( .A(n16163), .B(n16206), .Z(n16167) );
  XNOR U617 ( .A(n16715), .B(n16759), .Z(n16719) );
  XNOR U618 ( .A(n17068), .B(n17112), .Z(n17072) );
  XNOR U619 ( .A(n6098), .B(n6136), .Z(n6102) );
  XNOR U620 ( .A(n6450), .B(n6488), .Z(n6454) );
  XNOR U621 ( .A(n6802), .B(n6840), .Z(n6806) );
  XNOR U622 ( .A(n7154), .B(n7192), .Z(n7158) );
  XNOR U623 ( .A(n7506), .B(n7544), .Z(n7510) );
  XNOR U624 ( .A(n7858), .B(n7896), .Z(n7862) );
  XNOR U625 ( .A(n8210), .B(n8248), .Z(n8214) );
  XNOR U626 ( .A(n8562), .B(n8600), .Z(n8566) );
  XNOR U627 ( .A(n8914), .B(n8952), .Z(n8918) );
  XNOR U628 ( .A(n9266), .B(n9304), .Z(n9270) );
  XNOR U629 ( .A(n9613), .B(n9656), .Z(n9622) );
  XNOR U630 ( .A(n15993), .B(n16030), .Z(n15997) );
  XNOR U631 ( .A(n2878), .B(n2915), .Z(n2882) );
  XNOR U632 ( .A(n3239), .B(n3275), .Z(n3243) );
  XNOR U633 ( .A(n3599), .B(n3635), .Z(n3603) );
  XNOR U634 ( .A(n3959), .B(n3995), .Z(n3963) );
  XNOR U635 ( .A(n15646), .B(n15678), .Z(n15654) );
  XNOR U636 ( .A(n20171), .B(n20203), .Z(n20175) );
  XNOR U637 ( .A(n20075), .B(n20107), .Z(n20079) );
  XNOR U638 ( .A(n19955), .B(n19987), .Z(n19959) );
  XNOR U639 ( .A(n19811), .B(n19843), .Z(n19815) );
  XNOR U640 ( .A(n19643), .B(n19675), .Z(n19647) );
  XNOR U641 ( .A(n19451), .B(n19483), .Z(n19455) );
  XNOR U642 ( .A(n19235), .B(n19267), .Z(n19239) );
  XNOR U643 ( .A(n18995), .B(n19027), .Z(n18999) );
  XNOR U644 ( .A(n18731), .B(n18763), .Z(n18735) );
  XNOR U645 ( .A(n18443), .B(n18475), .Z(n18447) );
  XNOR U646 ( .A(n18131), .B(n18163), .Z(n18135) );
  XNOR U647 ( .A(n17795), .B(n17827), .Z(n17799) );
  XNOR U648 ( .A(n17430), .B(n17465), .Z(n17434) );
  XNOR U649 ( .A(n537), .B(n567), .Z(n541) );
  XNOR U650 ( .A(n898), .B(n928), .Z(n902) );
  XNOR U651 ( .A(n1259), .B(n1289), .Z(n1263) );
  XNOR U652 ( .A(n1620), .B(n1650), .Z(n1624) );
  XNOR U653 ( .A(n1981), .B(n2011), .Z(n1985) );
  XNOR U654 ( .A(n2342), .B(n2372), .Z(n2346) );
  XNOR U655 ( .A(n2703), .B(n2733), .Z(n2707) );
  XNOR U656 ( .A(n4504), .B(n4534), .Z(n4508) );
  XNOR U657 ( .A(n4864), .B(n4894), .Z(n4868) );
  XNOR U658 ( .A(n5938), .B(n5758), .Z(n5760) );
  XNOR U659 ( .A(n10509), .B(n10535), .Z(n10513) );
  XNOR U660 ( .A(n11249), .B(n11275), .Z(n11253) );
  XNOR U661 ( .A(n11602), .B(n11628), .Z(n11606) );
  XNOR U662 ( .A(n11954), .B(n11980), .Z(n11958) );
  XNOR U663 ( .A(n12306), .B(n12332), .Z(n12310) );
  XNOR U664 ( .A(n12658), .B(n12684), .Z(n12662) );
  XNOR U665 ( .A(n13010), .B(n13036), .Z(n13014) );
  XNOR U666 ( .A(n13362), .B(n13388), .Z(n13366) );
  XNOR U667 ( .A(n13714), .B(n13740), .Z(n13718) );
  XNOR U668 ( .A(n14066), .B(n14092), .Z(n14070) );
  XNOR U669 ( .A(n14418), .B(n14444), .Z(n14422) );
  XNOR U670 ( .A(n14770), .B(n14796), .Z(n14774) );
  XNOR U671 ( .A(n15122), .B(n15148), .Z(n15126) );
  XNOR U672 ( .A(n15469), .B(n15500), .Z(n15478) );
  XNOR U673 ( .A(n16730), .B(n16756), .Z(n16734) );
  XNOR U674 ( .A(n17083), .B(n17109), .Z(n17087) );
  XNOR U675 ( .A(n5943), .B(n5763), .Z(n5765) );
  XNOR U676 ( .A(n6113), .B(n6133), .Z(n6117) );
  XNOR U677 ( .A(n6465), .B(n6485), .Z(n6469) );
  XNOR U678 ( .A(n6817), .B(n6837), .Z(n6821) );
  XNOR U679 ( .A(n7169), .B(n7189), .Z(n7173) );
  XNOR U680 ( .A(n7521), .B(n7541), .Z(n7525) );
  XNOR U681 ( .A(n7873), .B(n7893), .Z(n7877) );
  XNOR U682 ( .A(n8225), .B(n8245), .Z(n8229) );
  XNOR U683 ( .A(n8577), .B(n8597), .Z(n8581) );
  XNOR U684 ( .A(n8929), .B(n8949), .Z(n8933) );
  XNOR U685 ( .A(n9281), .B(n9301), .Z(n9285) );
  XNOR U686 ( .A(n9633), .B(n9653), .Z(n9637) );
  XNOR U687 ( .A(n9985), .B(n10005), .Z(n9989) );
  XNOR U688 ( .A(n10342), .B(n10358), .Z(n10337) );
  ANDN U689 ( .B(n3084), .A(n3085), .Z(n2904) );
  ANDN U690 ( .B(n3804), .A(n3805), .Z(n3624) );
  ANDN U691 ( .B(n4704), .A(n4705), .Z(n4524) );
  XNOR U692 ( .A(n2226), .B(n2395), .Z(n2231) );
  XNOR U693 ( .A(n2587), .B(n2756), .Z(n2592) );
  XNOR U694 ( .A(n2948), .B(n3117), .Z(n2953) );
  XNOR U695 ( .A(n3308), .B(n3477), .Z(n3313) );
  XNOR U696 ( .A(n3668), .B(n3837), .Z(n3673) );
  XNOR U697 ( .A(n4748), .B(n4917), .Z(n4753) );
  XNOR U698 ( .A(n5646), .B(n5467), .Z(n5469) );
  XNOR U699 ( .A(n5823), .B(n5643), .Z(n5645) );
  XNOR U700 ( .A(n13423), .B(n13588), .Z(n13428) );
  XNOR U701 ( .A(n13775), .B(n13940), .Z(n13780) );
  XNOR U702 ( .A(n14127), .B(n14292), .Z(n14132) );
  XNOR U703 ( .A(n14479), .B(n14644), .Z(n14484) );
  XNOR U704 ( .A(n14831), .B(n14996), .Z(n14836) );
  XNOR U705 ( .A(n1690), .B(n1853), .Z(n1694) );
  XNOR U706 ( .A(n4034), .B(n4196), .Z(n4038) );
  XNOR U707 ( .A(n8287), .B(n8445), .Z(n8291) );
  XNOR U708 ( .A(n8639), .B(n8797), .Z(n8643) );
  XNOR U709 ( .A(n8991), .B(n9149), .Z(n8995) );
  XNOR U710 ( .A(n13253), .B(n13411), .Z(n13257) );
  XNOR U711 ( .A(n15365), .B(n15523), .Z(n15369) );
  XNOR U712 ( .A(n17861), .B(n18019), .Z(n17865) );
  XNOR U713 ( .A(n17510), .B(n17668), .Z(n17514) );
  XNOR U714 ( .A(n2056), .B(n2213), .Z(n2060) );
  XNOR U715 ( .A(n4399), .B(n4555), .Z(n4403) );
  XNOR U716 ( .A(n5833), .B(n5653), .Z(n5655) );
  XNOR U717 ( .A(n6532), .B(n6684), .Z(n6540) );
  XNOR U718 ( .A(n6884), .B(n7036), .Z(n6888) );
  XNOR U719 ( .A(n7236), .B(n7388), .Z(n7240) );
  XNOR U720 ( .A(n7764), .B(n7916), .Z(n7768) );
  XNOR U721 ( .A(n8116), .B(n8268), .Z(n8120) );
  XNOR U722 ( .A(n9348), .B(n9500), .Z(n9352) );
  XNOR U723 ( .A(n9700), .B(n9852), .Z(n9704) );
  XNOR U724 ( .A(n10052), .B(n10204), .Z(n10056) );
  XNOR U725 ( .A(n10404), .B(n10556), .Z(n10408) );
  XNOR U726 ( .A(n10758), .B(n10939), .Z(n10762) );
  XNOR U727 ( .A(n11150), .B(n10970), .Z(n10972) );
  XNOR U728 ( .A(n11327), .B(n11147), .Z(n11149) );
  XNOR U729 ( .A(n11503), .B(n11324), .Z(n11326) );
  XNOR U730 ( .A(n11679), .B(n11500), .Z(n11502) );
  XNOR U731 ( .A(n11668), .B(n11825), .Z(n11677) );
  XNOR U732 ( .A(n12026), .B(n12178), .Z(n12034) );
  XNOR U733 ( .A(n12378), .B(n12530), .Z(n12382) );
  XNOR U734 ( .A(n12730), .B(n12882), .Z(n12734) );
  XNOR U735 ( .A(n13082), .B(n13234), .Z(n13086) );
  XNOR U736 ( .A(n15722), .B(n15874), .Z(n15726) );
  XNOR U737 ( .A(n16248), .B(n16420), .Z(n16252) );
  XNOR U738 ( .A(n16631), .B(n16451), .Z(n16453) );
  XNOR U739 ( .A(n16808), .B(n16628), .Z(n16630) );
  XNOR U740 ( .A(n16984), .B(n16805), .Z(n16807) );
  XNOR U741 ( .A(n17160), .B(n16981), .Z(n16983) );
  XNOR U742 ( .A(n17149), .B(n17301), .Z(n17158) );
  XNOR U743 ( .A(n2603), .B(n2753), .Z(n2607) );
  XNOR U744 ( .A(n2964), .B(n3114), .Z(n2968) );
  XNOR U745 ( .A(n3324), .B(n3474), .Z(n3328) );
  XNOR U746 ( .A(n3684), .B(n3834), .Z(n3688) );
  XNOR U747 ( .A(n4764), .B(n4914), .Z(n4768) );
  XNOR U748 ( .A(n5661), .B(n5482), .Z(n5484) );
  XNOR U749 ( .A(n5838), .B(n5658), .Z(n5660) );
  XNOR U750 ( .A(n6008), .B(n6154), .Z(n6012) );
  XNOR U751 ( .A(n6355), .B(n6506), .Z(n6364) );
  XNOR U752 ( .A(n7593), .B(n7739), .Z(n7597) );
  XNOR U753 ( .A(n13791), .B(n13937), .Z(n13795) );
  XNOR U754 ( .A(n14143), .B(n14289), .Z(n14147) );
  XNOR U755 ( .A(n14495), .B(n14641), .Z(n14499) );
  XNOR U756 ( .A(n14847), .B(n14993), .Z(n14851) );
  XNOR U757 ( .A(n1886), .B(n2030), .Z(n1890) );
  XNOR U758 ( .A(n4049), .B(n4193), .Z(n4053) );
  XNOR U759 ( .A(n8654), .B(n8794), .Z(n8658) );
  XNOR U760 ( .A(n9006), .B(n9146), .Z(n9010) );
  XNOR U761 ( .A(n13620), .B(n13760), .Z(n13624) );
  XNOR U762 ( .A(n15380), .B(n15520), .Z(n15384) );
  XNOR U763 ( .A(n18500), .B(n18640), .Z(n18504) );
  XNOR U764 ( .A(n18200), .B(n18340), .Z(n18204) );
  XNOR U765 ( .A(n17876), .B(n18016), .Z(n17880) );
  XNOR U766 ( .A(n17525), .B(n17665), .Z(n17529) );
  XNOR U767 ( .A(n1520), .B(n1670), .Z(n1524) );
  XNOR U768 ( .A(n2432), .B(n2571), .Z(n2436) );
  XNOR U769 ( .A(n4414), .B(n4552), .Z(n4418) );
  XNOR U770 ( .A(n5848), .B(n5668), .Z(n5670) );
  XNOR U771 ( .A(n7251), .B(n7385), .Z(n7255) );
  XNOR U772 ( .A(n8131), .B(n8265), .Z(n8135) );
  XNOR U773 ( .A(n9363), .B(n9497), .Z(n9367) );
  XNOR U774 ( .A(n9715), .B(n9849), .Z(n9719) );
  XNOR U775 ( .A(n10067), .B(n10201), .Z(n10071) );
  XNOR U776 ( .A(n10419), .B(n10553), .Z(n10423) );
  XNOR U777 ( .A(n10773), .B(n10933), .Z(n10777) );
  XNOR U778 ( .A(n11165), .B(n10985), .Z(n10987) );
  XNOR U779 ( .A(n11342), .B(n11162), .Z(n11164) );
  XNOR U780 ( .A(n11518), .B(n11339), .Z(n11341) );
  XNOR U781 ( .A(n11694), .B(n11515), .Z(n11517) );
  XNOR U782 ( .A(n11870), .B(n11691), .Z(n11693) );
  XNOR U783 ( .A(n12046), .B(n11867), .Z(n11869) );
  XNOR U784 ( .A(n12222), .B(n12043), .Z(n12045) );
  XNOR U785 ( .A(n12398), .B(n12219), .Z(n12221) );
  XNOR U786 ( .A(n12397), .B(n12527), .Z(n12392) );
  XNOR U787 ( .A(n12745), .B(n12879), .Z(n12749) );
  XNOR U788 ( .A(n13097), .B(n13231), .Z(n13101) );
  XNOR U789 ( .A(n13449), .B(n13583), .Z(n13453) );
  XNOR U790 ( .A(n15737), .B(n15871), .Z(n15741) );
  XNOR U791 ( .A(n16263), .B(n16414), .Z(n16267) );
  XNOR U792 ( .A(n16646), .B(n16466), .Z(n16468) );
  XNOR U793 ( .A(n16823), .B(n16643), .Z(n16645) );
  XNOR U794 ( .A(n16999), .B(n16820), .Z(n16822) );
  XNOR U795 ( .A(n17175), .B(n16996), .Z(n16998) );
  XNOR U796 ( .A(n17169), .B(n17298), .Z(n17173) );
  XNOR U797 ( .A(n2979), .B(n3111), .Z(n2983) );
  XNOR U798 ( .A(n3339), .B(n3471), .Z(n3343) );
  XNOR U799 ( .A(n3699), .B(n3831), .Z(n3703) );
  XNOR U800 ( .A(n4779), .B(n4911), .Z(n4783) );
  XNOR U801 ( .A(n5676), .B(n5497), .Z(n5499) );
  XNOR U802 ( .A(n5853), .B(n5673), .Z(n5675) );
  XNOR U803 ( .A(n6023), .B(n6151), .Z(n6027) );
  XNOR U804 ( .A(n6375), .B(n6503), .Z(n6379) );
  XNOR U805 ( .A(n6727), .B(n6855), .Z(n6731) );
  XNOR U806 ( .A(n7084), .B(n7208), .Z(n7079) );
  XNOR U807 ( .A(n8488), .B(n8616), .Z(n8492) );
  XNOR U808 ( .A(n14158), .B(n14286), .Z(n14162) );
  XNOR U809 ( .A(n14510), .B(n14638), .Z(n14514) );
  XNOR U810 ( .A(n14862), .B(n14990), .Z(n14866) );
  XNOR U811 ( .A(n1901), .B(n2027), .Z(n1905) );
  XNOR U812 ( .A(n2262), .B(n2388), .Z(n2266) );
  XNOR U813 ( .A(n4064), .B(n4190), .Z(n4068) );
  XNOR U814 ( .A(n7965), .B(n8087), .Z(n7969) );
  XNOR U815 ( .A(n9021), .B(n9143), .Z(n9025) );
  XNOR U816 ( .A(n13987), .B(n14109), .Z(n13991) );
  XNOR U817 ( .A(n15395), .B(n15517), .Z(n15399) );
  XNOR U818 ( .A(n18791), .B(n18913), .Z(n18795) );
  XNOR U819 ( .A(n18515), .B(n18637), .Z(n18519) );
  XNOR U820 ( .A(n18215), .B(n18337), .Z(n18219) );
  XNOR U821 ( .A(n17891), .B(n18013), .Z(n17895) );
  XNOR U822 ( .A(n17540), .B(n17662), .Z(n17544) );
  XNOR U823 ( .A(n1535), .B(n1667), .Z(n1539) );
  XNOR U824 ( .A(n1154), .B(n1310), .Z(n1158) );
  XNOR U825 ( .A(n2808), .B(n2929), .Z(n2812) );
  XNOR U826 ( .A(n4429), .B(n4549), .Z(n4433) );
  XNOR U827 ( .A(n7794), .B(n7910), .Z(n7798) );
  XNOR U828 ( .A(n8322), .B(n8438), .Z(n8326) );
  XNOR U829 ( .A(n9378), .B(n9494), .Z(n9382) );
  XNOR U830 ( .A(n9730), .B(n9846), .Z(n9734) );
  XNOR U831 ( .A(n10082), .B(n10198), .Z(n10086) );
  XNOR U832 ( .A(n10434), .B(n10550), .Z(n10438) );
  XNOR U833 ( .A(n10788), .B(n10927), .Z(n10792) );
  XNOR U834 ( .A(n11180), .B(n11000), .Z(n11002) );
  XNOR U835 ( .A(n11357), .B(n11177), .Z(n11179) );
  XNOR U836 ( .A(n11533), .B(n11354), .Z(n11356) );
  XNOR U837 ( .A(n11709), .B(n11530), .Z(n11532) );
  XNOR U838 ( .A(n11885), .B(n11706), .Z(n11708) );
  XNOR U839 ( .A(n12061), .B(n11882), .Z(n11884) );
  XNOR U840 ( .A(n12237), .B(n12058), .Z(n12060) );
  XNOR U841 ( .A(n12413), .B(n12234), .Z(n12236) );
  XNOR U842 ( .A(n12589), .B(n12410), .Z(n12412) );
  XNOR U843 ( .A(n12765), .B(n12586), .Z(n12588) );
  XNOR U844 ( .A(n12754), .B(n12875), .Z(n12763) );
  XNOR U845 ( .A(n13112), .B(n13228), .Z(n13120) );
  XNOR U846 ( .A(n13464), .B(n13580), .Z(n13468) );
  XNOR U847 ( .A(n13816), .B(n13932), .Z(n13820) );
  XNOR U848 ( .A(n15752), .B(n15868), .Z(n15756) );
  XNOR U849 ( .A(n16278), .B(n16408), .Z(n16282) );
  XNOR U850 ( .A(n16661), .B(n16481), .Z(n16483) );
  XNOR U851 ( .A(n16838), .B(n16658), .Z(n16660) );
  XNOR U852 ( .A(n17014), .B(n16835), .Z(n16837) );
  XNOR U853 ( .A(n17190), .B(n17011), .Z(n17013) );
  XNOR U854 ( .A(n17184), .B(n17295), .Z(n17188) );
  XNOR U855 ( .A(n3354), .B(n3468), .Z(n3358) );
  XNOR U856 ( .A(n3714), .B(n3828), .Z(n3718) );
  XNOR U857 ( .A(n4794), .B(n4908), .Z(n4798) );
  XNOR U858 ( .A(n5691), .B(n5512), .Z(n5514) );
  XNOR U859 ( .A(n5868), .B(n5688), .Z(n5690) );
  XNOR U860 ( .A(n5862), .B(n5972), .Z(n5866) );
  XNOR U861 ( .A(n6214), .B(n6324), .Z(n6218) );
  XNOR U862 ( .A(n6566), .B(n6676), .Z(n6570) );
  XNOR U863 ( .A(n6918), .B(n7028), .Z(n6922) );
  XNOR U864 ( .A(n7270), .B(n7380), .Z(n7274) );
  XNOR U865 ( .A(n7627), .B(n7733), .Z(n7622) );
  XNOR U866 ( .A(n8855), .B(n8965), .Z(n8859) );
  XNOR U867 ( .A(n14525), .B(n14635), .Z(n14529) );
  XNOR U868 ( .A(n14877), .B(n14987), .Z(n14881) );
  XNOR U869 ( .A(n1916), .B(n2024), .Z(n1920) );
  XNOR U870 ( .A(n2277), .B(n2385), .Z(n2281) );
  XNOR U871 ( .A(n2638), .B(n2746), .Z(n2642) );
  XNOR U872 ( .A(n4079), .B(n4187), .Z(n4083) );
  XNOR U873 ( .A(n14354), .B(n14458), .Z(n14358) );
  XNOR U874 ( .A(n15410), .B(n15514), .Z(n15414) );
  XNOR U875 ( .A(n19286), .B(n19390), .Z(n19290) );
  XNOR U876 ( .A(n19058), .B(n19162), .Z(n19062) );
  XNOR U877 ( .A(n18806), .B(n18910), .Z(n18810) );
  XNOR U878 ( .A(n18530), .B(n18634), .Z(n18534) );
  XNOR U879 ( .A(n18230), .B(n18334), .Z(n18234) );
  XNOR U880 ( .A(n17906), .B(n18010), .Z(n17910) );
  XNOR U881 ( .A(n17555), .B(n17659), .Z(n17559) );
  XNOR U882 ( .A(n1359), .B(n1486), .Z(n1363) );
  XNOR U883 ( .A(n978), .B(n1129), .Z(n982) );
  XNOR U884 ( .A(n3184), .B(n3286), .Z(n3188) );
  XNOR U885 ( .A(n4444), .B(n4546), .Z(n4448) );
  XNOR U886 ( .A(n8337), .B(n8435), .Z(n8341) );
  XNOR U887 ( .A(n8689), .B(n8787), .Z(n8693) );
  XNOR U888 ( .A(n9393), .B(n9491), .Z(n9397) );
  XNOR U889 ( .A(n9745), .B(n9843), .Z(n9749) );
  XNOR U890 ( .A(n10097), .B(n10195), .Z(n10101) );
  XNOR U891 ( .A(n10449), .B(n10547), .Z(n10453) );
  XNOR U892 ( .A(n10803), .B(n10921), .Z(n10807) );
  XNOR U893 ( .A(n11195), .B(n11015), .Z(n11017) );
  XNOR U894 ( .A(n11372), .B(n11192), .Z(n11194) );
  XNOR U895 ( .A(n11548), .B(n11369), .Z(n11371) );
  XNOR U896 ( .A(n11724), .B(n11545), .Z(n11547) );
  XNOR U897 ( .A(n11900), .B(n11721), .Z(n11723) );
  XNOR U898 ( .A(n12076), .B(n11897), .Z(n11899) );
  XNOR U899 ( .A(n12252), .B(n12073), .Z(n12075) );
  XNOR U900 ( .A(n12428), .B(n12249), .Z(n12251) );
  XNOR U901 ( .A(n12604), .B(n12425), .Z(n12427) );
  XNOR U902 ( .A(n12780), .B(n12601), .Z(n12603) );
  XNOR U903 ( .A(n12956), .B(n12777), .Z(n12779) );
  XNOR U904 ( .A(n13132), .B(n12953), .Z(n12955) );
  XNOR U905 ( .A(n13308), .B(n13129), .Z(n13131) );
  XNOR U906 ( .A(n13484), .B(n13305), .Z(n13307) );
  XNOR U907 ( .A(n13483), .B(n13577), .Z(n13478) );
  XNOR U908 ( .A(n13831), .B(n13929), .Z(n13835) );
  XNOR U909 ( .A(n14183), .B(n14281), .Z(n14187) );
  XNOR U910 ( .A(n15767), .B(n15865), .Z(n15771) );
  XNOR U911 ( .A(n16293), .B(n16402), .Z(n16297) );
  XNOR U912 ( .A(n16676), .B(n16496), .Z(n16498) );
  XNOR U913 ( .A(n16853), .B(n16673), .Z(n16675) );
  XNOR U914 ( .A(n17029), .B(n16850), .Z(n16852) );
  XNOR U915 ( .A(n17205), .B(n17026), .Z(n17028) );
  XNOR U916 ( .A(n17199), .B(n17292), .Z(n17203) );
  XNOR U917 ( .A(n1008), .B(n1123), .Z(n1012) );
  XNOR U918 ( .A(n1555), .B(n1663), .Z(n1559) );
  XNOR U919 ( .A(n3729), .B(n3825), .Z(n3733) );
  XNOR U920 ( .A(n4809), .B(n4905), .Z(n4813) );
  XNOR U921 ( .A(n5706), .B(n5527), .Z(n5529) );
  XNOR U922 ( .A(n5883), .B(n5703), .Z(n5705) );
  XNOR U923 ( .A(n5877), .B(n5969), .Z(n5881) );
  XNOR U924 ( .A(n6229), .B(n6321), .Z(n6233) );
  XNOR U925 ( .A(n6581), .B(n6673), .Z(n6585) );
  XNOR U926 ( .A(n6933), .B(n7025), .Z(n6937) );
  XNOR U927 ( .A(n7285), .B(n7377), .Z(n7289) );
  XNOR U928 ( .A(n7637), .B(n7729), .Z(n7641) );
  XNOR U929 ( .A(n7984), .B(n8081), .Z(n7993) );
  XNOR U930 ( .A(n14892), .B(n14984), .Z(n14896) );
  XNOR U931 ( .A(n1389), .B(n1480), .Z(n1393) );
  XNOR U932 ( .A(n1931), .B(n2021), .Z(n1935) );
  XNOR U933 ( .A(n2292), .B(n2382), .Z(n2296) );
  XNOR U934 ( .A(n2653), .B(n2743), .Z(n2657) );
  XNOR U935 ( .A(n3014), .B(n3104), .Z(n3018) );
  XNOR U936 ( .A(n4094), .B(n4184), .Z(n4098) );
  XNOR U937 ( .A(n14721), .B(n14807), .Z(n14725) );
  XNOR U938 ( .A(n15425), .B(n15511), .Z(n15429) );
  XNOR U939 ( .A(n19505), .B(n19591), .Z(n19509) );
  XNOR U940 ( .A(n19301), .B(n19387), .Z(n19305) );
  XNOR U941 ( .A(n19073), .B(n19159), .Z(n19077) );
  XNOR U942 ( .A(n18821), .B(n18907), .Z(n18825) );
  XNOR U943 ( .A(n18545), .B(n18631), .Z(n18549) );
  XNOR U944 ( .A(n18245), .B(n18331), .Z(n18249) );
  XNOR U945 ( .A(n17921), .B(n18007), .Z(n17925) );
  XNOR U946 ( .A(n17570), .B(n17656), .Z(n17574) );
  XNOR U947 ( .A(n993), .B(n1126), .Z(n997) );
  XNOR U948 ( .A(n612), .B(n769), .Z(n616) );
  XNOR U949 ( .A(n1755), .B(n1840), .Z(n1759) );
  XNOR U950 ( .A(n3559), .B(n3643), .Z(n3563) );
  XNOR U951 ( .A(n4459), .B(n4543), .Z(n4463) );
  XNOR U952 ( .A(n5893), .B(n5713), .Z(n5715) );
  XNOR U953 ( .A(n8880), .B(n8960), .Z(n8884) );
  XNOR U954 ( .A(n9232), .B(n9312), .Z(n9236) );
  XNOR U955 ( .A(n9760), .B(n9840), .Z(n9764) );
  XNOR U956 ( .A(n10112), .B(n10192), .Z(n10116) );
  XNOR U957 ( .A(n10464), .B(n10544), .Z(n10468) );
  XNOR U958 ( .A(n10818), .B(n10915), .Z(n10822) );
  XNOR U959 ( .A(n11210), .B(n11030), .Z(n11032) );
  XNOR U960 ( .A(n11387), .B(n11207), .Z(n11209) );
  XNOR U961 ( .A(n11563), .B(n11384), .Z(n11386) );
  XNOR U962 ( .A(n11739), .B(n11560), .Z(n11562) );
  XNOR U963 ( .A(n11915), .B(n11736), .Z(n11738) );
  XNOR U964 ( .A(n12091), .B(n11912), .Z(n11914) );
  XNOR U965 ( .A(n12267), .B(n12088), .Z(n12090) );
  XNOR U966 ( .A(n12443), .B(n12264), .Z(n12266) );
  XNOR U967 ( .A(n12619), .B(n12440), .Z(n12442) );
  XNOR U968 ( .A(n12795), .B(n12616), .Z(n12618) );
  XNOR U969 ( .A(n12971), .B(n12792), .Z(n12794) );
  XNOR U970 ( .A(n13147), .B(n12968), .Z(n12970) );
  XNOR U971 ( .A(n13323), .B(n13144), .Z(n13146) );
  XNOR U972 ( .A(n13499), .B(n13320), .Z(n13322) );
  XNOR U973 ( .A(n13675), .B(n13496), .Z(n13498) );
  XNOR U974 ( .A(n13851), .B(n13672), .Z(n13674) );
  XNOR U975 ( .A(n13840), .B(n13925), .Z(n13849) );
  XNOR U976 ( .A(n14198), .B(n14278), .Z(n14206) );
  XNOR U977 ( .A(n14550), .B(n14630), .Z(n14554) );
  XNOR U978 ( .A(n15782), .B(n15862), .Z(n15786) );
  XNOR U979 ( .A(n16308), .B(n16396), .Z(n16312) );
  XNOR U980 ( .A(n16691), .B(n16511), .Z(n16513) );
  XNOR U981 ( .A(n16868), .B(n16688), .Z(n16690) );
  XNOR U982 ( .A(n17044), .B(n16865), .Z(n16867) );
  XNOR U983 ( .A(n17220), .B(n17041), .Z(n17043) );
  XNOR U984 ( .A(n17214), .B(n17289), .Z(n17218) );
  XNOR U985 ( .A(n1214), .B(n1298), .Z(n1218) );
  XNOR U986 ( .A(n452), .B(n584), .Z(n456) );
  XNOR U987 ( .A(n662), .B(n759), .Z(n666) );
  XNOR U988 ( .A(n4824), .B(n4902), .Z(n4828) );
  XNOR U989 ( .A(n5721), .B(n5542), .Z(n5544) );
  XNOR U990 ( .A(n5898), .B(n5718), .Z(n5720) );
  XNOR U991 ( .A(n6068), .B(n6142), .Z(n6072) );
  XNOR U992 ( .A(n6420), .B(n6494), .Z(n6424) );
  XNOR U993 ( .A(n6772), .B(n6846), .Z(n6776) );
  XNOR U994 ( .A(n7124), .B(n7198), .Z(n7128) );
  XNOR U995 ( .A(n7476), .B(n7550), .Z(n7480) );
  XNOR U996 ( .A(n7828), .B(n7902), .Z(n7832) );
  XNOR U997 ( .A(n8180), .B(n8254), .Z(n8184) );
  XNOR U998 ( .A(n8527), .B(n8606), .Z(n8536) );
  XNOR U999 ( .A(n15259), .B(n15333), .Z(n15263) );
  XNOR U1000 ( .A(n647), .B(n762), .Z(n651) );
  XNOR U1001 ( .A(n2307), .B(n2379), .Z(n2311) );
  XNOR U1002 ( .A(n2668), .B(n2740), .Z(n2672) );
  XNOR U1003 ( .A(n3029), .B(n3101), .Z(n3033) );
  XNOR U1004 ( .A(n3389), .B(n3461), .Z(n3393) );
  XNOR U1005 ( .A(n4109), .B(n4181), .Z(n4113) );
  XNOR U1006 ( .A(n15088), .B(n15156), .Z(n15092) );
  XNOR U1007 ( .A(n19856), .B(n19924), .Z(n19860) );
  XNOR U1008 ( .A(n19700), .B(n19768), .Z(n19704) );
  XNOR U1009 ( .A(n19520), .B(n19588), .Z(n19524) );
  XNOR U1010 ( .A(n19316), .B(n19384), .Z(n19320) );
  XNOR U1011 ( .A(n19088), .B(n19156), .Z(n19092) );
  XNOR U1012 ( .A(n18836), .B(n18904), .Z(n18840) );
  XNOR U1013 ( .A(n18560), .B(n18628), .Z(n18564) );
  XNOR U1014 ( .A(n18260), .B(n18328), .Z(n18264) );
  XNOR U1015 ( .A(n17936), .B(n18004), .Z(n17940) );
  XNOR U1016 ( .A(n17585), .B(n17653), .Z(n17589) );
  XNOR U1017 ( .A(n627), .B(n766), .Z(n631) );
  XNOR U1018 ( .A(n1229), .B(n1295), .Z(n1233) );
  XNOR U1019 ( .A(n1590), .B(n1656), .Z(n1594) );
  XNOR U1020 ( .A(n1951), .B(n2017), .Z(n1955) );
  XNOR U1021 ( .A(n3754), .B(n3820), .Z(n3758) );
  XNOR U1022 ( .A(n4474), .B(n4540), .Z(n4478) );
  XNOR U1023 ( .A(n9247), .B(n9309), .Z(n9255) );
  XNOR U1024 ( .A(n9775), .B(n9837), .Z(n9779) );
  XNOR U1025 ( .A(n10127), .B(n10189), .Z(n10131) );
  XNOR U1026 ( .A(n10479), .B(n10541), .Z(n10483) );
  XNOR U1027 ( .A(n10833), .B(n10909), .Z(n10837) );
  XNOR U1028 ( .A(n11225), .B(n11045), .Z(n11047) );
  XNOR U1029 ( .A(n11402), .B(n11222), .Z(n11224) );
  XNOR U1030 ( .A(n11578), .B(n11399), .Z(n11401) );
  XNOR U1031 ( .A(n11754), .B(n11575), .Z(n11577) );
  XNOR U1032 ( .A(n11930), .B(n11751), .Z(n11753) );
  XNOR U1033 ( .A(n12106), .B(n11927), .Z(n11929) );
  XNOR U1034 ( .A(n12282), .B(n12103), .Z(n12105) );
  XNOR U1035 ( .A(n12458), .B(n12279), .Z(n12281) );
  XNOR U1036 ( .A(n12634), .B(n12455), .Z(n12457) );
  XNOR U1037 ( .A(n12810), .B(n12631), .Z(n12633) );
  XNOR U1038 ( .A(n12986), .B(n12807), .Z(n12809) );
  XNOR U1039 ( .A(n13162), .B(n12983), .Z(n12985) );
  XNOR U1040 ( .A(n13338), .B(n13159), .Z(n13161) );
  XNOR U1041 ( .A(n13514), .B(n13335), .Z(n13337) );
  XNOR U1042 ( .A(n13690), .B(n13511), .Z(n13513) );
  XNOR U1043 ( .A(n13866), .B(n13687), .Z(n13689) );
  XNOR U1044 ( .A(n14042), .B(n13863), .Z(n13865) );
  XNOR U1045 ( .A(n14218), .B(n14039), .Z(n14041) );
  XNOR U1046 ( .A(n14394), .B(n14215), .Z(n14217) );
  XNOR U1047 ( .A(n14570), .B(n14391), .Z(n14393) );
  XNOR U1048 ( .A(n14569), .B(n14627), .Z(n14564) );
  XNOR U1049 ( .A(n14917), .B(n14979), .Z(n14921) );
  XNOR U1050 ( .A(n15797), .B(n15859), .Z(n15801) );
  XNOR U1051 ( .A(n16323), .B(n16390), .Z(n16327) );
  XNOR U1052 ( .A(n16706), .B(n16526), .Z(n16528) );
  XNOR U1053 ( .A(n16883), .B(n16703), .Z(n16705) );
  XNOR U1054 ( .A(n17059), .B(n16880), .Z(n16882) );
  XNOR U1055 ( .A(n17235), .B(n17056), .Z(n17058) );
  XNOR U1056 ( .A(n17229), .B(n17286), .Z(n17233) );
  XNOR U1057 ( .A(n677), .B(n756), .Z(n681) );
  XNOR U1058 ( .A(n4839), .B(n4899), .Z(n4843) );
  XNOR U1059 ( .A(n5736), .B(n5557), .Z(n5559) );
  XNOR U1060 ( .A(n5913), .B(n5733), .Z(n5735) );
  XNOR U1061 ( .A(n5907), .B(n5963), .Z(n5911) );
  XNOR U1062 ( .A(n6259), .B(n6315), .Z(n6263) );
  XNOR U1063 ( .A(n6611), .B(n6667), .Z(n6615) );
  XNOR U1064 ( .A(n6963), .B(n7019), .Z(n6967) );
  XNOR U1065 ( .A(n7315), .B(n7371), .Z(n7319) );
  XNOR U1066 ( .A(n7667), .B(n7723), .Z(n7671) );
  XNOR U1067 ( .A(n8019), .B(n8075), .Z(n8023) );
  XNOR U1068 ( .A(n8371), .B(n8427), .Z(n8375) );
  XNOR U1069 ( .A(n8723), .B(n8779), .Z(n8727) );
  XNOR U1070 ( .A(n9070), .B(n9131), .Z(n9079) );
  XNOR U1071 ( .A(n9604), .B(n9660), .Z(n9608) );
  XNOR U1072 ( .A(n15626), .B(n15682), .Z(n15630) );
  XNOR U1073 ( .A(n2683), .B(n2737), .Z(n2687) );
  XNOR U1074 ( .A(n3044), .B(n3098), .Z(n3048) );
  XNOR U1075 ( .A(n3404), .B(n3458), .Z(n3408) );
  XNOR U1076 ( .A(n15455), .B(n15505), .Z(n15459) );
  XNOR U1077 ( .A(n20003), .B(n20053), .Z(n20007) );
  XNOR U1078 ( .A(n19871), .B(n19921), .Z(n19875) );
  XNOR U1079 ( .A(n19715), .B(n19765), .Z(n19719) );
  XNOR U1080 ( .A(n19535), .B(n19585), .Z(n19539) );
  XNOR U1081 ( .A(n19331), .B(n19381), .Z(n19335) );
  XNOR U1082 ( .A(n19103), .B(n19153), .Z(n19107) );
  XNOR U1083 ( .A(n18851), .B(n18901), .Z(n18855) );
  XNOR U1084 ( .A(n18575), .B(n18625), .Z(n18579) );
  XNOR U1085 ( .A(n18275), .B(n18325), .Z(n18279) );
  XNOR U1086 ( .A(n17951), .B(n18001), .Z(n17955) );
  XNOR U1087 ( .A(n17600), .B(n17650), .Z(n17604) );
  XNOR U1088 ( .A(n702), .B(n751), .Z(n706) );
  XNOR U1089 ( .A(n1063), .B(n1112), .Z(n1067) );
  XNOR U1090 ( .A(n1424), .B(n1473), .Z(n1428) );
  XNOR U1091 ( .A(n1785), .B(n1834), .Z(n1789) );
  XNOR U1092 ( .A(n2146), .B(n2195), .Z(n2150) );
  XNOR U1093 ( .A(n2507), .B(n2556), .Z(n2511) );
  XNOR U1094 ( .A(n3769), .B(n3817), .Z(n3773) );
  XNOR U1095 ( .A(n4129), .B(n4177), .Z(n4133) );
  XNOR U1096 ( .A(n4489), .B(n4537), .Z(n4493) );
  XNOR U1097 ( .A(n10494), .B(n10538), .Z(n10498) );
  XNOR U1098 ( .A(n10848), .B(n10903), .Z(n10852) );
  XNOR U1099 ( .A(n11240), .B(n11060), .Z(n11062) );
  XNOR U1100 ( .A(n11417), .B(n11237), .Z(n11239) );
  XNOR U1101 ( .A(n11593), .B(n11414), .Z(n11416) );
  XNOR U1102 ( .A(n11769), .B(n11590), .Z(n11592) );
  XNOR U1103 ( .A(n11945), .B(n11766), .Z(n11768) );
  XNOR U1104 ( .A(n12121), .B(n11942), .Z(n11944) );
  XNOR U1105 ( .A(n12297), .B(n12118), .Z(n12120) );
  XNOR U1106 ( .A(n12473), .B(n12294), .Z(n12296) );
  XNOR U1107 ( .A(n12649), .B(n12470), .Z(n12472) );
  XNOR U1108 ( .A(n12825), .B(n12646), .Z(n12648) );
  XNOR U1109 ( .A(n13001), .B(n12822), .Z(n12824) );
  XNOR U1110 ( .A(n13177), .B(n12998), .Z(n13000) );
  XNOR U1111 ( .A(n13353), .B(n13174), .Z(n13176) );
  XNOR U1112 ( .A(n13529), .B(n13350), .Z(n13352) );
  XNOR U1113 ( .A(n13705), .B(n13526), .Z(n13528) );
  XNOR U1114 ( .A(n13881), .B(n13702), .Z(n13704) );
  XNOR U1115 ( .A(n14057), .B(n13878), .Z(n13880) );
  XNOR U1116 ( .A(n14233), .B(n14054), .Z(n14056) );
  XNOR U1117 ( .A(n14409), .B(n14230), .Z(n14232) );
  XNOR U1118 ( .A(n14585), .B(n14406), .Z(n14408) );
  XNOR U1119 ( .A(n14761), .B(n14582), .Z(n14584) );
  XNOR U1120 ( .A(n14937), .B(n14758), .Z(n14760) );
  XNOR U1121 ( .A(n14926), .B(n14975), .Z(n14935) );
  XNOR U1122 ( .A(n15284), .B(n15328), .Z(n15292) );
  XNOR U1123 ( .A(n16338), .B(n16384), .Z(n16342) );
  XNOR U1124 ( .A(n16721), .B(n16541), .Z(n16543) );
  XNOR U1125 ( .A(n16898), .B(n16718), .Z(n16720) );
  XNOR U1126 ( .A(n17074), .B(n16895), .Z(n16897) );
  XNOR U1127 ( .A(n17250), .B(n17071), .Z(n17073) );
  XNOR U1128 ( .A(n17244), .B(n17283), .Z(n17248) );
  XNOR U1129 ( .A(n4854), .B(n4896), .Z(n4858) );
  XNOR U1130 ( .A(n5751), .B(n5572), .Z(n5574) );
  XNOR U1131 ( .A(n5928), .B(n5748), .Z(n5750) );
  XNOR U1132 ( .A(n5922), .B(n5960), .Z(n5926) );
  XNOR U1133 ( .A(n6274), .B(n6312), .Z(n6278) );
  XNOR U1134 ( .A(n6626), .B(n6664), .Z(n6630) );
  XNOR U1135 ( .A(n6978), .B(n7016), .Z(n6982) );
  XNOR U1136 ( .A(n7330), .B(n7368), .Z(n7334) );
  XNOR U1137 ( .A(n7682), .B(n7720), .Z(n7686) );
  XNOR U1138 ( .A(n8034), .B(n8072), .Z(n8038) );
  XNOR U1139 ( .A(n8386), .B(n8424), .Z(n8390) );
  XNOR U1140 ( .A(n8738), .B(n8776), .Z(n8742) );
  XNOR U1141 ( .A(n9090), .B(n9128), .Z(n9094) );
  XNOR U1142 ( .A(n9442), .B(n9480), .Z(n9446) );
  XNOR U1143 ( .A(n9799), .B(n9833), .Z(n9794) );
  XNOR U1144 ( .A(n10147), .B(n10185), .Z(n10151) );
  XNOR U1145 ( .A(n15998), .B(n16029), .Z(n16002) );
  XNOR U1146 ( .A(n20210), .B(n20242), .Z(n20214) );
  XNOR U1147 ( .A(n20126), .B(n20158), .Z(n20130) );
  XNOR U1148 ( .A(n20018), .B(n20050), .Z(n20022) );
  XNOR U1149 ( .A(n19886), .B(n19918), .Z(n19890) );
  XNOR U1150 ( .A(n19730), .B(n19762), .Z(n19734) );
  XNOR U1151 ( .A(n19550), .B(n19582), .Z(n19554) );
  XNOR U1152 ( .A(n19346), .B(n19378), .Z(n19350) );
  XNOR U1153 ( .A(n19118), .B(n19150), .Z(n19122) );
  XNOR U1154 ( .A(n18866), .B(n18898), .Z(n18870) );
  XNOR U1155 ( .A(n18590), .B(n18622), .Z(n18594) );
  XNOR U1156 ( .A(n18290), .B(n18322), .Z(n18294) );
  XNOR U1157 ( .A(n17966), .B(n17998), .Z(n17970) );
  XNOR U1158 ( .A(n17615), .B(n17647), .Z(n17619) );
  XNOR U1159 ( .A(n717), .B(n748), .Z(n721) );
  XNOR U1160 ( .A(n1078), .B(n1109), .Z(n1082) );
  XNOR U1161 ( .A(n1439), .B(n1470), .Z(n1443) );
  XNOR U1162 ( .A(n1800), .B(n1831), .Z(n1804) );
  XNOR U1163 ( .A(n2161), .B(n2192), .Z(n2165) );
  XNOR U1164 ( .A(n2522), .B(n2553), .Z(n2526) );
  XNOR U1165 ( .A(n2883), .B(n2914), .Z(n2887) );
  XNOR U1166 ( .A(n3244), .B(n3274), .Z(n3248) );
  XNOR U1167 ( .A(n3604), .B(n3634), .Z(n3608) );
  XNOR U1168 ( .A(n3964), .B(n3994), .Z(n3968) );
  XNOR U1169 ( .A(n4324), .B(n4354), .Z(n4328) );
  XNOR U1170 ( .A(n4684), .B(n4714), .Z(n4688) );
  XNOR U1171 ( .A(n10863), .B(n10897), .Z(n10867) );
  XNOR U1172 ( .A(n11255), .B(n11075), .Z(n11077) );
  XNOR U1173 ( .A(n11432), .B(n11252), .Z(n11254) );
  XNOR U1174 ( .A(n11608), .B(n11429), .Z(n11431) );
  XNOR U1175 ( .A(n11784), .B(n11605), .Z(n11607) );
  XNOR U1176 ( .A(n11960), .B(n11781), .Z(n11783) );
  XNOR U1177 ( .A(n12136), .B(n11957), .Z(n11959) );
  XNOR U1178 ( .A(n12312), .B(n12133), .Z(n12135) );
  XNOR U1179 ( .A(n12488), .B(n12309), .Z(n12311) );
  XNOR U1180 ( .A(n12664), .B(n12485), .Z(n12487) );
  XNOR U1181 ( .A(n12840), .B(n12661), .Z(n12663) );
  XNOR U1182 ( .A(n13016), .B(n12837), .Z(n12839) );
  XNOR U1183 ( .A(n13192), .B(n13013), .Z(n13015) );
  XNOR U1184 ( .A(n13368), .B(n13189), .Z(n13191) );
  XNOR U1185 ( .A(n13544), .B(n13365), .Z(n13367) );
  XNOR U1186 ( .A(n13720), .B(n13541), .Z(n13543) );
  XNOR U1187 ( .A(n13896), .B(n13717), .Z(n13719) );
  XNOR U1188 ( .A(n14072), .B(n13893), .Z(n13895) );
  XNOR U1189 ( .A(n14248), .B(n14069), .Z(n14071) );
  XNOR U1190 ( .A(n14424), .B(n14245), .Z(n14247) );
  XNOR U1191 ( .A(n14600), .B(n14421), .Z(n14423) );
  XNOR U1192 ( .A(n14776), .B(n14597), .Z(n14599) );
  XNOR U1193 ( .A(n14952), .B(n14773), .Z(n14775) );
  XNOR U1194 ( .A(n15128), .B(n14949), .Z(n14951) );
  XNOR U1195 ( .A(n15304), .B(n15125), .Z(n15127) );
  XNOR U1196 ( .A(n15480), .B(n15301), .Z(n15303) );
  XNOR U1197 ( .A(n15656), .B(n15477), .Z(n15479) );
  XNOR U1198 ( .A(n15655), .B(n15677), .Z(n15650) );
  XNOR U1199 ( .A(n16353), .B(n16378), .Z(n16357) );
  XNOR U1200 ( .A(n16736), .B(n16556), .Z(n16558) );
  XNOR U1201 ( .A(n16913), .B(n16733), .Z(n16735) );
  XNOR U1202 ( .A(n17089), .B(n16910), .Z(n16912) );
  XNOR U1203 ( .A(n17265), .B(n17086), .Z(n17088) );
  XNOR U1204 ( .A(n17259), .B(n17280), .Z(n17263) );
  XNOR U1205 ( .A(n5049), .B(n5402), .Z(n5053) );
  XNOR U1206 ( .A(n5766), .B(n5587), .Z(n5589) );
  XNOR U1207 ( .A(n5760), .B(n5780), .Z(n5764) );
  XNOR U1208 ( .A(n5937), .B(n5957), .Z(n5941) );
  XNOR U1209 ( .A(n6289), .B(n6309), .Z(n6293) );
  XNOR U1210 ( .A(n6641), .B(n6661), .Z(n6645) );
  XNOR U1211 ( .A(n6993), .B(n7013), .Z(n6997) );
  XNOR U1212 ( .A(n7345), .B(n7365), .Z(n7349) );
  XNOR U1213 ( .A(n7697), .B(n7717), .Z(n7701) );
  XNOR U1214 ( .A(n8049), .B(n8069), .Z(n8053) );
  XNOR U1215 ( .A(n8401), .B(n8421), .Z(n8405) );
  XNOR U1216 ( .A(n8753), .B(n8773), .Z(n8757) );
  XNOR U1217 ( .A(n9105), .B(n9125), .Z(n9109) );
  XNOR U1218 ( .A(n9457), .B(n9477), .Z(n9461) );
  XNOR U1219 ( .A(n9809), .B(n9829), .Z(n9813) );
  XNOR U1220 ( .A(n10343), .B(n10164), .Z(n10166) );
  XNOR U1221 ( .A(n10514), .B(n10534), .Z(n10522) );
  ANDN U1222 ( .B(n3444), .A(n3445), .Z(n3264) );
  ANDN U1223 ( .B(n4164), .A(n4165), .Z(n3984) );
  ANDN U1224 ( .B(n4884), .A(n4885), .Z(n4704) );
  XNOR U1225 ( .A(n17680), .B(n17850), .Z(n17684) );
  XNOR U1226 ( .A(n17315), .B(n17488), .Z(n17320) );
  XNOR U1227 ( .A(n4928), .B(n5450), .Z(n4933) );
  XNOR U1228 ( .A(n5463), .B(n5627), .Z(n5468) );
  XNOR U1229 ( .A(n5639), .B(n5804), .Z(n5644) );
  XNOR U1230 ( .A(n5999), .B(n5820), .Z(n5821) );
  XNOR U1231 ( .A(n7049), .B(n7214), .Z(n7054) );
  XNOR U1232 ( .A(n7577), .B(n7742), .Z(n7582) );
  XNOR U1233 ( .A(n7929), .B(n8094), .Z(n7934) );
  XNOR U1234 ( .A(n8457), .B(n8622), .Z(n8462) );
  XNOR U1235 ( .A(n8809), .B(n8974), .Z(n8814) );
  XNOR U1236 ( .A(n9161), .B(n9326), .Z(n9166) );
  XNOR U1237 ( .A(n10217), .B(n10382), .Z(n10222) );
  XNOR U1238 ( .A(n10569), .B(n10736), .Z(n10574) );
  XNOR U1239 ( .A(n10956), .B(n11121), .Z(n10961) );
  XNOR U1240 ( .A(n11133), .B(n11298), .Z(n11138) );
  XNOR U1241 ( .A(n11491), .B(n11652), .Z(n11487) );
  XNOR U1242 ( .A(n11839), .B(n12004), .Z(n11844) );
  XNOR U1243 ( .A(n12191), .B(n12356), .Z(n12196) );
  XNOR U1244 ( .A(n12543), .B(n12708), .Z(n12548) );
  XNOR U1245 ( .A(n15711), .B(n15876), .Z(n15716) );
  XNOR U1246 ( .A(n16062), .B(n16226), .Z(n16067) );
  XNOR U1247 ( .A(n16437), .B(n16602), .Z(n16442) );
  XNOR U1248 ( .A(n16614), .B(n16779), .Z(n16619) );
  XNOR U1249 ( .A(n16972), .B(n17133), .Z(n16968) );
  XNOR U1250 ( .A(n2412), .B(n2575), .Z(n2416) );
  XNOR U1251 ( .A(n2773), .B(n2936), .Z(n2777) );
  XNOR U1252 ( .A(n3134), .B(n3296), .Z(n3138) );
  XNOR U1253 ( .A(n3494), .B(n3656), .Z(n3498) );
  XNOR U1254 ( .A(n3854), .B(n4016), .Z(n3858) );
  XNOR U1255 ( .A(n4214), .B(n4376), .Z(n4218) );
  XNOR U1256 ( .A(n7407), .B(n7565), .Z(n7411) );
  XNOR U1257 ( .A(n9519), .B(n9677), .Z(n9523) );
  XNOR U1258 ( .A(n13605), .B(n13763), .Z(n13609) );
  XNOR U1259 ( .A(n13957), .B(n14115), .Z(n13961) );
  XNOR U1260 ( .A(n14309), .B(n14467), .Z(n14313) );
  XNOR U1261 ( .A(n14661), .B(n14819), .Z(n14665) );
  XNOR U1262 ( .A(n15013), .B(n15171), .Z(n15017) );
  XNOR U1263 ( .A(n1504), .B(n1673), .Z(n1509) );
  XNOR U1264 ( .A(n2237), .B(n2393), .Z(n2241) );
  XNOR U1265 ( .A(n4579), .B(n4735), .Z(n4583) );
  XNOR U1266 ( .A(n6360), .B(n6508), .Z(n6355) );
  XNOR U1267 ( .A(n6708), .B(n6860), .Z(n6712) );
  XNOR U1268 ( .A(n9876), .B(n10028), .Z(n9880) );
  XNOR U1269 ( .A(n13258), .B(n13410), .Z(n13262) );
  XNOR U1270 ( .A(n15370), .B(n15522), .Z(n15374) );
  XNOR U1271 ( .A(n18031), .B(n18183), .Z(n18035) );
  XNOR U1272 ( .A(n17695), .B(n17847), .Z(n17699) );
  XNOR U1273 ( .A(n17325), .B(n17485), .Z(n17334) );
  XNOR U1274 ( .A(n1700), .B(n1851), .Z(n1704) );
  XNOR U1275 ( .A(n4944), .B(n5444), .Z(n4948) );
  XNOR U1276 ( .A(n5479), .B(n5624), .Z(n5483) );
  XNOR U1277 ( .A(n5655), .B(n5801), .Z(n5659) );
  XNOR U1278 ( .A(n6014), .B(n5835), .Z(n5837) );
  XNOR U1279 ( .A(n6190), .B(n6011), .Z(n6013) );
  XNOR U1280 ( .A(n6366), .B(n6187), .Z(n6189) );
  XNOR U1281 ( .A(n6542), .B(n6363), .Z(n6365) );
  XNOR U1282 ( .A(n7065), .B(n7211), .Z(n7069) );
  XNOR U1283 ( .A(n7945), .B(n8091), .Z(n7949) );
  XNOR U1284 ( .A(n8473), .B(n8619), .Z(n8477) );
  XNOR U1285 ( .A(n8825), .B(n8971), .Z(n8829) );
  XNOR U1286 ( .A(n9177), .B(n9323), .Z(n9181) );
  XNOR U1287 ( .A(n10233), .B(n10379), .Z(n10237) );
  XNOR U1288 ( .A(n10585), .B(n10733), .Z(n10589) );
  XNOR U1289 ( .A(n10972), .B(n11118), .Z(n10976) );
  XNOR U1290 ( .A(n11332), .B(n11152), .Z(n11154) );
  XNOR U1291 ( .A(n11508), .B(n11329), .Z(n11331) );
  XNOR U1292 ( .A(n11684), .B(n11505), .Z(n11507) );
  XNOR U1293 ( .A(n11860), .B(n11681), .Z(n11683) );
  XNOR U1294 ( .A(n11849), .B(n12000), .Z(n11858) );
  XNOR U1295 ( .A(n12207), .B(n12353), .Z(n12215) );
  XNOR U1296 ( .A(n12559), .B(n12705), .Z(n12563) );
  XNOR U1297 ( .A(n12911), .B(n13057), .Z(n12915) );
  XNOR U1298 ( .A(n15727), .B(n15873), .Z(n15731) );
  XNOR U1299 ( .A(n16078), .B(n16223), .Z(n16082) );
  XNOR U1300 ( .A(n16453), .B(n16599), .Z(n16457) );
  XNOR U1301 ( .A(n16630), .B(n16776), .Z(n16634) );
  XNOR U1302 ( .A(n16807), .B(n16953), .Z(n16811) );
  XNOR U1303 ( .A(n16983), .B(n17129), .Z(n16987) );
  XNOR U1304 ( .A(n2066), .B(n2211), .Z(n2070) );
  XNOR U1305 ( .A(n2788), .B(n2933), .Z(n2792) );
  XNOR U1306 ( .A(n3149), .B(n3293), .Z(n3153) );
  XNOR U1307 ( .A(n3509), .B(n3653), .Z(n3513) );
  XNOR U1308 ( .A(n3869), .B(n4013), .Z(n3873) );
  XNOR U1309 ( .A(n4229), .B(n4373), .Z(n4233) );
  XNOR U1310 ( .A(n7422), .B(n7562), .Z(n7426) );
  XNOR U1311 ( .A(n7774), .B(n7914), .Z(n7778) );
  XNOR U1312 ( .A(n8302), .B(n8442), .Z(n8306) );
  XNOR U1313 ( .A(n9534), .B(n9674), .Z(n9538) );
  XNOR U1314 ( .A(n13972), .B(n14112), .Z(n13976) );
  XNOR U1315 ( .A(n14324), .B(n14464), .Z(n14328) );
  XNOR U1316 ( .A(n14676), .B(n14816), .Z(n14680) );
  XNOR U1317 ( .A(n15028), .B(n15168), .Z(n15032) );
  XNOR U1318 ( .A(n2613), .B(n2751), .Z(n2617) );
  XNOR U1319 ( .A(n4594), .B(n4732), .Z(n4598) );
  XNOR U1320 ( .A(n6903), .B(n7033), .Z(n6898) );
  XNOR U1321 ( .A(n9891), .B(n10025), .Z(n9895) );
  XNOR U1322 ( .A(n13625), .B(n13759), .Z(n13629) );
  XNOR U1323 ( .A(n15385), .B(n15519), .Z(n15389) );
  XNOR U1324 ( .A(n18646), .B(n18780), .Z(n18650) );
  XNOR U1325 ( .A(n18358), .B(n18492), .Z(n18362) );
  XNOR U1326 ( .A(n18046), .B(n18180), .Z(n18050) );
  XNOR U1327 ( .A(n17710), .B(n17844), .Z(n17714) );
  XNOR U1328 ( .A(n17345), .B(n17482), .Z(n17349) );
  XNOR U1329 ( .A(n1334), .B(n1491), .Z(n1338) );
  XNOR U1330 ( .A(n4959), .B(n5438), .Z(n4963) );
  XNOR U1331 ( .A(n5494), .B(n5621), .Z(n5498) );
  XNOR U1332 ( .A(n5670), .B(n5798), .Z(n5674) );
  XNOR U1333 ( .A(n6029), .B(n5850), .Z(n5852) );
  XNOR U1334 ( .A(n6205), .B(n6026), .Z(n6028) );
  XNOR U1335 ( .A(n6381), .B(n6202), .Z(n6204) );
  XNOR U1336 ( .A(n6557), .B(n6378), .Z(n6380) );
  XNOR U1337 ( .A(n6733), .B(n6554), .Z(n6556) );
  XNOR U1338 ( .A(n6909), .B(n6730), .Z(n6732) );
  XNOR U1339 ( .A(n7085), .B(n6906), .Z(n6908) );
  XNOR U1340 ( .A(n7256), .B(n7384), .Z(n7264) );
  XNOR U1341 ( .A(n8840), .B(n8968), .Z(n8844) );
  XNOR U1342 ( .A(n9192), .B(n9320), .Z(n9196) );
  XNOR U1343 ( .A(n10248), .B(n10376), .Z(n10252) );
  XNOR U1344 ( .A(n10600), .B(n10730), .Z(n10604) );
  XNOR U1345 ( .A(n11170), .B(n10990), .Z(n10992) );
  XNOR U1346 ( .A(n11347), .B(n11167), .Z(n11169) );
  XNOR U1347 ( .A(n11523), .B(n11344), .Z(n11346) );
  XNOR U1348 ( .A(n11699), .B(n11520), .Z(n11522) );
  XNOR U1349 ( .A(n11875), .B(n11696), .Z(n11698) );
  XNOR U1350 ( .A(n12051), .B(n11872), .Z(n11874) );
  XNOR U1351 ( .A(n12227), .B(n12048), .Z(n12050) );
  XNOR U1352 ( .A(n12403), .B(n12224), .Z(n12226) );
  XNOR U1353 ( .A(n12579), .B(n12400), .Z(n12402) );
  XNOR U1354 ( .A(n12578), .B(n12702), .Z(n12573) );
  XNOR U1355 ( .A(n12926), .B(n13054), .Z(n12930) );
  XNOR U1356 ( .A(n13278), .B(n13406), .Z(n13282) );
  XNOR U1357 ( .A(n15742), .B(n15870), .Z(n15746) );
  XNOR U1358 ( .A(n16093), .B(n16220), .Z(n16097) );
  XNOR U1359 ( .A(n16468), .B(n16596), .Z(n16472) );
  XNOR U1360 ( .A(n16645), .B(n16773), .Z(n16649) );
  XNOR U1361 ( .A(n16822), .B(n16950), .Z(n16826) );
  XNOR U1362 ( .A(n16998), .B(n17126), .Z(n17002) );
  XNOR U1363 ( .A(n2081), .B(n2208), .Z(n2085) );
  XNOR U1364 ( .A(n2442), .B(n2569), .Z(n2446) );
  XNOR U1365 ( .A(n3164), .B(n3290), .Z(n3168) );
  XNOR U1366 ( .A(n3524), .B(n3650), .Z(n3528) );
  XNOR U1367 ( .A(n3884), .B(n4010), .Z(n3888) );
  XNOR U1368 ( .A(n4244), .B(n4370), .Z(n4248) );
  XNOR U1369 ( .A(n7613), .B(n7735), .Z(n7617) );
  XNOR U1370 ( .A(n8141), .B(n8263), .Z(n8145) );
  XNOR U1371 ( .A(n8669), .B(n8791), .Z(n8673) );
  XNOR U1372 ( .A(n9549), .B(n9671), .Z(n9553) );
  XNOR U1373 ( .A(n14339), .B(n14461), .Z(n14343) );
  XNOR U1374 ( .A(n14691), .B(n14813), .Z(n14695) );
  XNOR U1375 ( .A(n15043), .B(n15165), .Z(n15047) );
  XNOR U1376 ( .A(n1906), .B(n2026), .Z(n1910) );
  XNOR U1377 ( .A(n2989), .B(n3109), .Z(n2993) );
  XNOR U1378 ( .A(n4609), .B(n4729), .Z(n4613) );
  XNOR U1379 ( .A(n8498), .B(n8614), .Z(n8502) );
  XNOR U1380 ( .A(n9906), .B(n10022), .Z(n9910) );
  XNOR U1381 ( .A(n13992), .B(n14108), .Z(n13996) );
  XNOR U1382 ( .A(n15400), .B(n15516), .Z(n15404) );
  XNOR U1383 ( .A(n18925), .B(n19041), .Z(n18929) );
  XNOR U1384 ( .A(n18661), .B(n18777), .Z(n18665) );
  XNOR U1385 ( .A(n18373), .B(n18489), .Z(n18377) );
  XNOR U1386 ( .A(n18061), .B(n18177), .Z(n18065) );
  XNOR U1387 ( .A(n17725), .B(n17841), .Z(n17729) );
  XNOR U1388 ( .A(n17360), .B(n17479), .Z(n17364) );
  XNOR U1389 ( .A(n1540), .B(n1666), .Z(n1544) );
  XNOR U1390 ( .A(n1159), .B(n1309), .Z(n1163) );
  XNOR U1391 ( .A(n4974), .B(n5432), .Z(n4978) );
  XNOR U1392 ( .A(n5509), .B(n5618), .Z(n5513) );
  XNOR U1393 ( .A(n5685), .B(n5795), .Z(n5689) );
  XNOR U1394 ( .A(n6044), .B(n5865), .Z(n5867) );
  XNOR U1395 ( .A(n6220), .B(n6041), .Z(n6043) );
  XNOR U1396 ( .A(n6396), .B(n6217), .Z(n6219) );
  XNOR U1397 ( .A(n6572), .B(n6393), .Z(n6395) );
  XNOR U1398 ( .A(n6748), .B(n6569), .Z(n6571) );
  XNOR U1399 ( .A(n6924), .B(n6745), .Z(n6747) );
  XNOR U1400 ( .A(n7100), .B(n6921), .Z(n6923) );
  XNOR U1401 ( .A(n7276), .B(n7097), .Z(n7099) );
  XNOR U1402 ( .A(n7452), .B(n7273), .Z(n7275) );
  XNOR U1403 ( .A(n7628), .B(n7449), .Z(n7451) );
  XNOR U1404 ( .A(n9207), .B(n9317), .Z(n9211) );
  XNOR U1405 ( .A(n10263), .B(n10373), .Z(n10267) );
  XNOR U1406 ( .A(n10615), .B(n10727), .Z(n10619) );
  XNOR U1407 ( .A(n11185), .B(n11005), .Z(n11007) );
  XNOR U1408 ( .A(n11362), .B(n11182), .Z(n11184) );
  XNOR U1409 ( .A(n11538), .B(n11359), .Z(n11361) );
  XNOR U1410 ( .A(n11714), .B(n11535), .Z(n11537) );
  XNOR U1411 ( .A(n11890), .B(n11711), .Z(n11713) );
  XNOR U1412 ( .A(n12066), .B(n11887), .Z(n11889) );
  XNOR U1413 ( .A(n12242), .B(n12063), .Z(n12065) );
  XNOR U1414 ( .A(n12418), .B(n12239), .Z(n12241) );
  XNOR U1415 ( .A(n12594), .B(n12415), .Z(n12417) );
  XNOR U1416 ( .A(n12770), .B(n12591), .Z(n12593) );
  XNOR U1417 ( .A(n12946), .B(n12767), .Z(n12769) );
  XNOR U1418 ( .A(n12935), .B(n13050), .Z(n12944) );
  XNOR U1419 ( .A(n13293), .B(n13403), .Z(n13301) );
  XNOR U1420 ( .A(n13645), .B(n13755), .Z(n13649) );
  XNOR U1421 ( .A(n15757), .B(n15867), .Z(n15761) );
  XNOR U1422 ( .A(n16108), .B(n16217), .Z(n16112) );
  XNOR U1423 ( .A(n16483), .B(n16593), .Z(n16487) );
  XNOR U1424 ( .A(n16660), .B(n16770), .Z(n16664) );
  XNOR U1425 ( .A(n16837), .B(n16947), .Z(n16841) );
  XNOR U1426 ( .A(n17013), .B(n17123), .Z(n17017) );
  XNOR U1427 ( .A(n2457), .B(n2566), .Z(n2461) );
  XNOR U1428 ( .A(n2818), .B(n2927), .Z(n2822) );
  XNOR U1429 ( .A(n3539), .B(n3647), .Z(n3543) );
  XNOR U1430 ( .A(n3899), .B(n4007), .Z(n3903) );
  XNOR U1431 ( .A(n4259), .B(n4367), .Z(n4263) );
  XNOR U1432 ( .A(n7808), .B(n7908), .Z(n7803) );
  XNOR U1433 ( .A(n9036), .B(n9140), .Z(n9040) );
  XNOR U1434 ( .A(n9564), .B(n9668), .Z(n9568) );
  XNOR U1435 ( .A(n14706), .B(n14810), .Z(n14710) );
  XNOR U1436 ( .A(n15058), .B(n15162), .Z(n15062) );
  XNOR U1437 ( .A(n1921), .B(n2023), .Z(n1925) );
  XNOR U1438 ( .A(n2282), .B(n2384), .Z(n2286) );
  XNOR U1439 ( .A(n3364), .B(n3466), .Z(n3368) );
  XNOR U1440 ( .A(n4624), .B(n4726), .Z(n4628) );
  XNOR U1441 ( .A(n8161), .B(n8259), .Z(n8169) );
  XNOR U1442 ( .A(n8513), .B(n8611), .Z(n8517) );
  XNOR U1443 ( .A(n8865), .B(n8963), .Z(n8869) );
  XNOR U1444 ( .A(n9921), .B(n10019), .Z(n9925) );
  XNOR U1445 ( .A(n14359), .B(n14457), .Z(n14363) );
  XNOR U1446 ( .A(n15415), .B(n15513), .Z(n15419) );
  XNOR U1447 ( .A(n19396), .B(n19494), .Z(n19400) );
  XNOR U1448 ( .A(n19180), .B(n19278), .Z(n19184) );
  XNOR U1449 ( .A(n18940), .B(n19038), .Z(n18944) );
  XNOR U1450 ( .A(n18676), .B(n18774), .Z(n18680) );
  XNOR U1451 ( .A(n18388), .B(n18486), .Z(n18392) );
  XNOR U1452 ( .A(n18076), .B(n18174), .Z(n18080) );
  XNOR U1453 ( .A(n17740), .B(n17838), .Z(n17744) );
  XNOR U1454 ( .A(n17375), .B(n17476), .Z(n17379) );
  XNOR U1455 ( .A(n1174), .B(n1306), .Z(n1178) );
  XNOR U1456 ( .A(n793), .B(n949), .Z(n797) );
  XNOR U1457 ( .A(n4989), .B(n5426), .Z(n4993) );
  XNOR U1458 ( .A(n5524), .B(n5615), .Z(n5528) );
  XNOR U1459 ( .A(n5700), .B(n5792), .Z(n5704) );
  XNOR U1460 ( .A(n6059), .B(n5880), .Z(n5882) );
  XNOR U1461 ( .A(n6235), .B(n6056), .Z(n6058) );
  XNOR U1462 ( .A(n6411), .B(n6232), .Z(n6234) );
  XNOR U1463 ( .A(n6587), .B(n6408), .Z(n6410) );
  XNOR U1464 ( .A(n6763), .B(n6584), .Z(n6586) );
  XNOR U1465 ( .A(n6939), .B(n6760), .Z(n6762) );
  XNOR U1466 ( .A(n7115), .B(n6936), .Z(n6938) );
  XNOR U1467 ( .A(n7291), .B(n7112), .Z(n7114) );
  XNOR U1468 ( .A(n7467), .B(n7288), .Z(n7290) );
  XNOR U1469 ( .A(n7643), .B(n7464), .Z(n7466) );
  XNOR U1470 ( .A(n7819), .B(n7640), .Z(n7642) );
  XNOR U1471 ( .A(n7995), .B(n7816), .Z(n7818) );
  XNOR U1472 ( .A(n8171), .B(n7992), .Z(n7994) );
  XNOR U1473 ( .A(n10278), .B(n10370), .Z(n10282) );
  XNOR U1474 ( .A(n10630), .B(n10724), .Z(n10634) );
  XNOR U1475 ( .A(n11017), .B(n11109), .Z(n11021) );
  XNOR U1476 ( .A(n11377), .B(n11197), .Z(n11199) );
  XNOR U1477 ( .A(n11553), .B(n11374), .Z(n11376) );
  XNOR U1478 ( .A(n11729), .B(n11550), .Z(n11552) );
  XNOR U1479 ( .A(n11905), .B(n11726), .Z(n11728) );
  XNOR U1480 ( .A(n12081), .B(n11902), .Z(n11904) );
  XNOR U1481 ( .A(n12257), .B(n12078), .Z(n12080) );
  XNOR U1482 ( .A(n12433), .B(n12254), .Z(n12256) );
  XNOR U1483 ( .A(n12609), .B(n12430), .Z(n12432) );
  XNOR U1484 ( .A(n12785), .B(n12606), .Z(n12608) );
  XNOR U1485 ( .A(n12961), .B(n12782), .Z(n12784) );
  XNOR U1486 ( .A(n13137), .B(n12958), .Z(n12960) );
  XNOR U1487 ( .A(n13313), .B(n13134), .Z(n13136) );
  XNOR U1488 ( .A(n13489), .B(n13310), .Z(n13312) );
  XNOR U1489 ( .A(n13665), .B(n13486), .Z(n13488) );
  XNOR U1490 ( .A(n13664), .B(n13752), .Z(n13659) );
  XNOR U1491 ( .A(n14012), .B(n14104), .Z(n14016) );
  XNOR U1492 ( .A(n15772), .B(n15864), .Z(n15776) );
  XNOR U1493 ( .A(n16123), .B(n16214), .Z(n16127) );
  XNOR U1494 ( .A(n16498), .B(n16590), .Z(n16502) );
  XNOR U1495 ( .A(n16675), .B(n16767), .Z(n16679) );
  XNOR U1496 ( .A(n16852), .B(n16944), .Z(n16856) );
  XNOR U1497 ( .A(n17028), .B(n17120), .Z(n17032) );
  XNOR U1498 ( .A(n1204), .B(n1300), .Z(n1208) );
  XNOR U1499 ( .A(n2833), .B(n2924), .Z(n2837) );
  XNOR U1500 ( .A(n3194), .B(n3284), .Z(n3198) );
  XNOR U1501 ( .A(n3914), .B(n4004), .Z(n3918) );
  XNOR U1502 ( .A(n4274), .B(n4364), .Z(n4278) );
  XNOR U1503 ( .A(n9579), .B(n9665), .Z(n9583) );
  XNOR U1504 ( .A(n15073), .B(n15159), .Z(n15077) );
  XNOR U1505 ( .A(n828), .B(n942), .Z(n832) );
  XNOR U1506 ( .A(n1374), .B(n1483), .Z(n1378) );
  XNOR U1507 ( .A(n1936), .B(n2020), .Z(n1940) );
  XNOR U1508 ( .A(n2297), .B(n2381), .Z(n2301) );
  XNOR U1509 ( .A(n2658), .B(n2742), .Z(n2662) );
  XNOR U1510 ( .A(n3739), .B(n3823), .Z(n3743) );
  XNOR U1511 ( .A(n4639), .B(n4723), .Z(n4643) );
  XNOR U1512 ( .A(n8704), .B(n8784), .Z(n8712) );
  XNOR U1513 ( .A(n9056), .B(n9136), .Z(n9060) );
  XNOR U1514 ( .A(n9408), .B(n9488), .Z(n9412) );
  XNOR U1515 ( .A(n9936), .B(n10016), .Z(n9940) );
  XNOR U1516 ( .A(n14726), .B(n14806), .Z(n14730) );
  XNOR U1517 ( .A(n15430), .B(n15510), .Z(n15434) );
  XNOR U1518 ( .A(n19603), .B(n19683), .Z(n19607) );
  XNOR U1519 ( .A(n19411), .B(n19491), .Z(n19415) );
  XNOR U1520 ( .A(n19195), .B(n19275), .Z(n19199) );
  XNOR U1521 ( .A(n18955), .B(n19035), .Z(n18959) );
  XNOR U1522 ( .A(n18691), .B(n18771), .Z(n18695) );
  XNOR U1523 ( .A(n18403), .B(n18483), .Z(n18407) );
  XNOR U1524 ( .A(n18091), .B(n18171), .Z(n18095) );
  XNOR U1525 ( .A(n17755), .B(n17835), .Z(n17759) );
  XNOR U1526 ( .A(n17390), .B(n17473), .Z(n17394) );
  XNOR U1527 ( .A(n998), .B(n1125), .Z(n1002) );
  XNOR U1528 ( .A(n617), .B(n768), .Z(n621) );
  XNOR U1529 ( .A(n853), .B(n937), .Z(n857) );
  XNOR U1530 ( .A(n1580), .B(n1658), .Z(n1584) );
  XNOR U1531 ( .A(n5004), .B(n5420), .Z(n5008) );
  XNOR U1532 ( .A(n5539), .B(n5612), .Z(n5543) );
  XNOR U1533 ( .A(n5715), .B(n5789), .Z(n5719) );
  XNOR U1534 ( .A(n6074), .B(n5895), .Z(n5897) );
  XNOR U1535 ( .A(n6250), .B(n6071), .Z(n6073) );
  XNOR U1536 ( .A(n6426), .B(n6247), .Z(n6249) );
  XNOR U1537 ( .A(n6602), .B(n6423), .Z(n6425) );
  XNOR U1538 ( .A(n6778), .B(n6599), .Z(n6601) );
  XNOR U1539 ( .A(n6954), .B(n6775), .Z(n6777) );
  XNOR U1540 ( .A(n7130), .B(n6951), .Z(n6953) );
  XNOR U1541 ( .A(n7306), .B(n7127), .Z(n7129) );
  XNOR U1542 ( .A(n7482), .B(n7303), .Z(n7305) );
  XNOR U1543 ( .A(n7658), .B(n7479), .Z(n7481) );
  XNOR U1544 ( .A(n7834), .B(n7655), .Z(n7657) );
  XNOR U1545 ( .A(n8010), .B(n7831), .Z(n7833) );
  XNOR U1546 ( .A(n8186), .B(n8007), .Z(n8009) );
  XNOR U1547 ( .A(n8362), .B(n8183), .Z(n8185) );
  XNOR U1548 ( .A(n8538), .B(n8359), .Z(n8361) );
  XNOR U1549 ( .A(n8714), .B(n8535), .Z(n8537) );
  XNOR U1550 ( .A(n10293), .B(n10367), .Z(n10297) );
  XNOR U1551 ( .A(n10645), .B(n10721), .Z(n10649) );
  XNOR U1552 ( .A(n11032), .B(n11106), .Z(n11036) );
  XNOR U1553 ( .A(n11392), .B(n11212), .Z(n11214) );
  XNOR U1554 ( .A(n11568), .B(n11389), .Z(n11391) );
  XNOR U1555 ( .A(n11744), .B(n11565), .Z(n11567) );
  XNOR U1556 ( .A(n11920), .B(n11741), .Z(n11743) );
  XNOR U1557 ( .A(n12096), .B(n11917), .Z(n11919) );
  XNOR U1558 ( .A(n12272), .B(n12093), .Z(n12095) );
  XNOR U1559 ( .A(n12448), .B(n12269), .Z(n12271) );
  XNOR U1560 ( .A(n12624), .B(n12445), .Z(n12447) );
  XNOR U1561 ( .A(n12800), .B(n12621), .Z(n12623) );
  XNOR U1562 ( .A(n12976), .B(n12797), .Z(n12799) );
  XNOR U1563 ( .A(n13152), .B(n12973), .Z(n12975) );
  XNOR U1564 ( .A(n13328), .B(n13149), .Z(n13151) );
  XNOR U1565 ( .A(n13504), .B(n13325), .Z(n13327) );
  XNOR U1566 ( .A(n13680), .B(n13501), .Z(n13503) );
  XNOR U1567 ( .A(n13856), .B(n13677), .Z(n13679) );
  XNOR U1568 ( .A(n14032), .B(n13853), .Z(n13855) );
  XNOR U1569 ( .A(n14021), .B(n14100), .Z(n14030) );
  XNOR U1570 ( .A(n14379), .B(n14453), .Z(n14387) );
  XNOR U1571 ( .A(n15787), .B(n15861), .Z(n15791) );
  XNOR U1572 ( .A(n16138), .B(n16211), .Z(n16142) );
  XNOR U1573 ( .A(n16513), .B(n16587), .Z(n16517) );
  XNOR U1574 ( .A(n16690), .B(n16764), .Z(n16694) );
  XNOR U1575 ( .A(n16867), .B(n16941), .Z(n16871) );
  XNOR U1576 ( .A(n17043), .B(n17117), .Z(n17047) );
  XNOR U1577 ( .A(n1028), .B(n1119), .Z(n1032) );
  XNOR U1578 ( .A(n477), .B(n579), .Z(n481) );
  XNOR U1579 ( .A(n3209), .B(n3281), .Z(n3213) );
  XNOR U1580 ( .A(n3569), .B(n3641), .Z(n3573) );
  XNOR U1581 ( .A(n4289), .B(n4361), .Z(n4293) );
  XNOR U1582 ( .A(n15264), .B(n15332), .Z(n15268) );
  XNOR U1583 ( .A(n652), .B(n761), .Z(n656) );
  XNOR U1584 ( .A(n507), .B(n573), .Z(n511) );
  XNOR U1585 ( .A(n2131), .B(n2198), .Z(n2135) );
  XNOR U1586 ( .A(n2492), .B(n2559), .Z(n2496) );
  XNOR U1587 ( .A(n2853), .B(n2920), .Z(n2857) );
  XNOR U1588 ( .A(n3934), .B(n4000), .Z(n3938) );
  XNOR U1589 ( .A(n4654), .B(n4720), .Z(n4658) );
  XNOR U1590 ( .A(n9075), .B(n9133), .Z(n9070) );
  XNOR U1591 ( .A(n9423), .B(n9485), .Z(n9427) );
  XNOR U1592 ( .A(n9951), .B(n10013), .Z(n9955) );
  XNOR U1593 ( .A(n15093), .B(n15155), .Z(n15097) );
  XNOR U1594 ( .A(n19930), .B(n19992), .Z(n19934) );
  XNOR U1595 ( .A(n19786), .B(n19848), .Z(n19790) );
  XNOR U1596 ( .A(n19618), .B(n19680), .Z(n19622) );
  XNOR U1597 ( .A(n19426), .B(n19488), .Z(n19430) );
  XNOR U1598 ( .A(n19210), .B(n19272), .Z(n19214) );
  XNOR U1599 ( .A(n18970), .B(n19032), .Z(n18974) );
  XNOR U1600 ( .A(n18706), .B(n18768), .Z(n18710) );
  XNOR U1601 ( .A(n18418), .B(n18480), .Z(n18422) );
  XNOR U1602 ( .A(n18106), .B(n18168), .Z(n18110) );
  XNOR U1603 ( .A(n17770), .B(n17832), .Z(n17774) );
  XNOR U1604 ( .A(n17405), .B(n17470), .Z(n17409) );
  XNOR U1605 ( .A(n632), .B(n765), .Z(n636) );
  XNOR U1606 ( .A(n1234), .B(n1294), .Z(n1238) );
  XNOR U1607 ( .A(n1595), .B(n1655), .Z(n1599) );
  XNOR U1608 ( .A(n1956), .B(n2016), .Z(n1960) );
  XNOR U1609 ( .A(n5019), .B(n5414), .Z(n5023) );
  XNOR U1610 ( .A(n5554), .B(n5609), .Z(n5558) );
  XNOR U1611 ( .A(n5730), .B(n5786), .Z(n5734) );
  XNOR U1612 ( .A(n6089), .B(n5910), .Z(n5912) );
  XNOR U1613 ( .A(n6265), .B(n6086), .Z(n6088) );
  XNOR U1614 ( .A(n6441), .B(n6262), .Z(n6264) );
  XNOR U1615 ( .A(n6617), .B(n6438), .Z(n6440) );
  XNOR U1616 ( .A(n6793), .B(n6614), .Z(n6616) );
  XNOR U1617 ( .A(n6969), .B(n6790), .Z(n6792) );
  XNOR U1618 ( .A(n7145), .B(n6966), .Z(n6968) );
  XNOR U1619 ( .A(n7321), .B(n7142), .Z(n7144) );
  XNOR U1620 ( .A(n7497), .B(n7318), .Z(n7320) );
  XNOR U1621 ( .A(n7673), .B(n7494), .Z(n7496) );
  XNOR U1622 ( .A(n7849), .B(n7670), .Z(n7672) );
  XNOR U1623 ( .A(n8025), .B(n7846), .Z(n7848) );
  XNOR U1624 ( .A(n8201), .B(n8022), .Z(n8024) );
  XNOR U1625 ( .A(n8377), .B(n8198), .Z(n8200) );
  XNOR U1626 ( .A(n8553), .B(n8374), .Z(n8376) );
  XNOR U1627 ( .A(n8729), .B(n8550), .Z(n8552) );
  XNOR U1628 ( .A(n8905), .B(n8726), .Z(n8728) );
  XNOR U1629 ( .A(n9081), .B(n8902), .Z(n8904) );
  XNOR U1630 ( .A(n9257), .B(n9078), .Z(n9080) );
  XNOR U1631 ( .A(n9780), .B(n9836), .Z(n9784) );
  XNOR U1632 ( .A(n10308), .B(n10364), .Z(n10312) );
  XNOR U1633 ( .A(n10660), .B(n10718), .Z(n10664) );
  XNOR U1634 ( .A(n11230), .B(n11050), .Z(n11052) );
  XNOR U1635 ( .A(n11407), .B(n11227), .Z(n11229) );
  XNOR U1636 ( .A(n11583), .B(n11404), .Z(n11406) );
  XNOR U1637 ( .A(n11759), .B(n11580), .Z(n11582) );
  XNOR U1638 ( .A(n11935), .B(n11756), .Z(n11758) );
  XNOR U1639 ( .A(n12111), .B(n11932), .Z(n11934) );
  XNOR U1640 ( .A(n12287), .B(n12108), .Z(n12110) );
  XNOR U1641 ( .A(n12463), .B(n12284), .Z(n12286) );
  XNOR U1642 ( .A(n12639), .B(n12460), .Z(n12462) );
  XNOR U1643 ( .A(n12815), .B(n12636), .Z(n12638) );
  XNOR U1644 ( .A(n12991), .B(n12812), .Z(n12814) );
  XNOR U1645 ( .A(n13167), .B(n12988), .Z(n12990) );
  XNOR U1646 ( .A(n13343), .B(n13164), .Z(n13166) );
  XNOR U1647 ( .A(n13519), .B(n13340), .Z(n13342) );
  XNOR U1648 ( .A(n13695), .B(n13516), .Z(n13518) );
  XNOR U1649 ( .A(n13871), .B(n13692), .Z(n13694) );
  XNOR U1650 ( .A(n14047), .B(n13868), .Z(n13870) );
  XNOR U1651 ( .A(n14223), .B(n14044), .Z(n14046) );
  XNOR U1652 ( .A(n14399), .B(n14220), .Z(n14222) );
  XNOR U1653 ( .A(n14575), .B(n14396), .Z(n14398) );
  XNOR U1654 ( .A(n14751), .B(n14572), .Z(n14574) );
  XNOR U1655 ( .A(n14750), .B(n14802), .Z(n14745) );
  XNOR U1656 ( .A(n15802), .B(n15858), .Z(n15806) );
  XNOR U1657 ( .A(n16153), .B(n16208), .Z(n16157) );
  XNOR U1658 ( .A(n16528), .B(n16584), .Z(n16532) );
  XNOR U1659 ( .A(n16705), .B(n16761), .Z(n16709) );
  XNOR U1660 ( .A(n16882), .B(n16938), .Z(n16886) );
  XNOR U1661 ( .A(n17058), .B(n17114), .Z(n17062) );
  XNOR U1662 ( .A(n682), .B(n755), .Z(n686) );
  XNOR U1663 ( .A(n3584), .B(n3638), .Z(n3588) );
  XNOR U1664 ( .A(n15631), .B(n15681), .Z(n15635) );
  XNOR U1665 ( .A(n2688), .B(n2736), .Z(n2692) );
  XNOR U1666 ( .A(n3049), .B(n3097), .Z(n3053) );
  XNOR U1667 ( .A(n3409), .B(n3457), .Z(n3413) );
  XNOR U1668 ( .A(n3949), .B(n3997), .Z(n3953) );
  XNOR U1669 ( .A(n4309), .B(n4357), .Z(n4313) );
  XNOR U1670 ( .A(n4669), .B(n4717), .Z(n4673) );
  XNOR U1671 ( .A(n9618), .B(n9658), .Z(n9613) );
  XNOR U1672 ( .A(n15460), .B(n15504), .Z(n15464) );
  XNOR U1673 ( .A(n20065), .B(n20109), .Z(n20069) );
  XNOR U1674 ( .A(n19945), .B(n19989), .Z(n19949) );
  XNOR U1675 ( .A(n19801), .B(n19845), .Z(n19805) );
  XNOR U1676 ( .A(n19633), .B(n19677), .Z(n19637) );
  XNOR U1677 ( .A(n19441), .B(n19485), .Z(n19445) );
  XNOR U1678 ( .A(n19225), .B(n19269), .Z(n19229) );
  XNOR U1679 ( .A(n18985), .B(n19029), .Z(n18989) );
  XNOR U1680 ( .A(n18721), .B(n18765), .Z(n18725) );
  XNOR U1681 ( .A(n18433), .B(n18477), .Z(n18437) );
  XNOR U1682 ( .A(n18121), .B(n18165), .Z(n18125) );
  XNOR U1683 ( .A(n17785), .B(n17829), .Z(n17789) );
  XNOR U1684 ( .A(n17420), .B(n17467), .Z(n17424) );
  XNOR U1685 ( .A(n527), .B(n569), .Z(n531) );
  XNOR U1686 ( .A(n888), .B(n930), .Z(n892) );
  XNOR U1687 ( .A(n1249), .B(n1291), .Z(n1253) );
  XNOR U1688 ( .A(n1610), .B(n1652), .Z(n1614) );
  XNOR U1689 ( .A(n1971), .B(n2013), .Z(n1975) );
  XNOR U1690 ( .A(n2332), .B(n2374), .Z(n2336) );
  XNOR U1691 ( .A(n5034), .B(n5408), .Z(n5038) );
  XNOR U1692 ( .A(n5569), .B(n5606), .Z(n5573) );
  XNOR U1693 ( .A(n5745), .B(n5783), .Z(n5749) );
  XNOR U1694 ( .A(n6104), .B(n5925), .Z(n5927) );
  XNOR U1695 ( .A(n6280), .B(n6101), .Z(n6103) );
  XNOR U1696 ( .A(n6456), .B(n6277), .Z(n6279) );
  XNOR U1697 ( .A(n6632), .B(n6453), .Z(n6455) );
  XNOR U1698 ( .A(n6808), .B(n6629), .Z(n6631) );
  XNOR U1699 ( .A(n6984), .B(n6805), .Z(n6807) );
  XNOR U1700 ( .A(n7160), .B(n6981), .Z(n6983) );
  XNOR U1701 ( .A(n7336), .B(n7157), .Z(n7159) );
  XNOR U1702 ( .A(n7512), .B(n7333), .Z(n7335) );
  XNOR U1703 ( .A(n7688), .B(n7509), .Z(n7511) );
  XNOR U1704 ( .A(n7864), .B(n7685), .Z(n7687) );
  XNOR U1705 ( .A(n8040), .B(n7861), .Z(n7863) );
  XNOR U1706 ( .A(n8216), .B(n8037), .Z(n8039) );
  XNOR U1707 ( .A(n8392), .B(n8213), .Z(n8215) );
  XNOR U1708 ( .A(n8568), .B(n8389), .Z(n8391) );
  XNOR U1709 ( .A(n8744), .B(n8565), .Z(n8567) );
  XNOR U1710 ( .A(n8920), .B(n8741), .Z(n8743) );
  XNOR U1711 ( .A(n9096), .B(n8917), .Z(n8919) );
  XNOR U1712 ( .A(n9272), .B(n9093), .Z(n9095) );
  XNOR U1713 ( .A(n9448), .B(n9269), .Z(n9271) );
  XNOR U1714 ( .A(n9624), .B(n9445), .Z(n9447) );
  XNOR U1715 ( .A(n9800), .B(n9621), .Z(n9623) );
  XNOR U1716 ( .A(n9971), .B(n10009), .Z(n9979) );
  XNOR U1717 ( .A(n10323), .B(n10361), .Z(n10327) );
  XNOR U1718 ( .A(n10675), .B(n10715), .Z(n10679) );
  XNOR U1719 ( .A(n11062), .B(n11100), .Z(n11066) );
  XNOR U1720 ( .A(n11239), .B(n11277), .Z(n11243) );
  XNOR U1721 ( .A(n11598), .B(n11419), .Z(n11421) );
  XNOR U1722 ( .A(n11774), .B(n11595), .Z(n11597) );
  XNOR U1723 ( .A(n11950), .B(n11771), .Z(n11773) );
  XNOR U1724 ( .A(n12126), .B(n11947), .Z(n11949) );
  XNOR U1725 ( .A(n12302), .B(n12123), .Z(n12125) );
  XNOR U1726 ( .A(n12478), .B(n12299), .Z(n12301) );
  XNOR U1727 ( .A(n12654), .B(n12475), .Z(n12477) );
  XNOR U1728 ( .A(n12830), .B(n12651), .Z(n12653) );
  XNOR U1729 ( .A(n13006), .B(n12827), .Z(n12829) );
  XNOR U1730 ( .A(n13182), .B(n13003), .Z(n13005) );
  XNOR U1731 ( .A(n13358), .B(n13179), .Z(n13181) );
  XNOR U1732 ( .A(n13534), .B(n13355), .Z(n13357) );
  XNOR U1733 ( .A(n13710), .B(n13531), .Z(n13533) );
  XNOR U1734 ( .A(n13886), .B(n13707), .Z(n13709) );
  XNOR U1735 ( .A(n14062), .B(n13883), .Z(n13885) );
  XNOR U1736 ( .A(n14238), .B(n14059), .Z(n14061) );
  XNOR U1737 ( .A(n14414), .B(n14235), .Z(n14237) );
  XNOR U1738 ( .A(n14590), .B(n14411), .Z(n14413) );
  XNOR U1739 ( .A(n14766), .B(n14587), .Z(n14589) );
  XNOR U1740 ( .A(n14942), .B(n14763), .Z(n14765) );
  XNOR U1741 ( .A(n15118), .B(n14939), .Z(n14941) );
  XNOR U1742 ( .A(n15107), .B(n15150), .Z(n15116) );
  XNOR U1743 ( .A(n16168), .B(n16205), .Z(n16172) );
  XNOR U1744 ( .A(n16543), .B(n16581), .Z(n16547) );
  XNOR U1745 ( .A(n16720), .B(n16758), .Z(n16724) );
  XNOR U1746 ( .A(n16897), .B(n16935), .Z(n16901) );
  XNOR U1747 ( .A(n17073), .B(n17111), .Z(n17077) );
  XNOR U1748 ( .A(n3064), .B(n3094), .Z(n3068) );
  XNOR U1749 ( .A(n3424), .B(n3454), .Z(n3428) );
  XNOR U1750 ( .A(n3784), .B(n3814), .Z(n3788) );
  XNOR U1751 ( .A(n4144), .B(n4174), .Z(n4148) );
  XNOR U1752 ( .A(n5761), .B(n5582), .Z(n5584) );
  XNOR U1753 ( .A(n15827), .B(n15853), .Z(n15835) );
  XNOR U1754 ( .A(n20248), .B(n20274), .Z(n20252) );
  XNOR U1755 ( .A(n20176), .B(n20202), .Z(n20180) );
  XNOR U1756 ( .A(n20080), .B(n20106), .Z(n20084) );
  XNOR U1757 ( .A(n19960), .B(n19986), .Z(n19964) );
  XNOR U1758 ( .A(n19816), .B(n19842), .Z(n19820) );
  XNOR U1759 ( .A(n19648), .B(n19674), .Z(n19652) );
  XNOR U1760 ( .A(n19456), .B(n19482), .Z(n19460) );
  XNOR U1761 ( .A(n19240), .B(n19266), .Z(n19244) );
  XNOR U1762 ( .A(n19000), .B(n19026), .Z(n19004) );
  XNOR U1763 ( .A(n18736), .B(n18762), .Z(n18740) );
  XNOR U1764 ( .A(n18448), .B(n18474), .Z(n18452) );
  XNOR U1765 ( .A(n18136), .B(n18162), .Z(n18140) );
  XNOR U1766 ( .A(n17800), .B(n17826), .Z(n17804) );
  XNOR U1767 ( .A(n17435), .B(n17464), .Z(n17439) );
  XNOR U1768 ( .A(n542), .B(n566), .Z(n546) );
  XNOR U1769 ( .A(n903), .B(n927), .Z(n907) );
  XNOR U1770 ( .A(n1264), .B(n1288), .Z(n1268) );
  XNOR U1771 ( .A(n1625), .B(n1649), .Z(n1629) );
  XNOR U1772 ( .A(n1986), .B(n2010), .Z(n1990) );
  XNOR U1773 ( .A(n2347), .B(n2371), .Z(n2351) );
  XNOR U1774 ( .A(n2708), .B(n2732), .Z(n2712) );
  XNOR U1775 ( .A(n4509), .B(n4533), .Z(n4513) );
  XNOR U1776 ( .A(n4869), .B(n4893), .Z(n4873) );
  XNOR U1777 ( .A(n6119), .B(n5940), .Z(n5942) );
  XNOR U1778 ( .A(n6295), .B(n6116), .Z(n6118) );
  XNOR U1779 ( .A(n6471), .B(n6292), .Z(n6294) );
  XNOR U1780 ( .A(n6647), .B(n6468), .Z(n6470) );
  XNOR U1781 ( .A(n6823), .B(n6644), .Z(n6646) );
  XNOR U1782 ( .A(n6999), .B(n6820), .Z(n6822) );
  XNOR U1783 ( .A(n7175), .B(n6996), .Z(n6998) );
  XNOR U1784 ( .A(n7351), .B(n7172), .Z(n7174) );
  XNOR U1785 ( .A(n7527), .B(n7348), .Z(n7350) );
  XNOR U1786 ( .A(n7703), .B(n7524), .Z(n7526) );
  XNOR U1787 ( .A(n7879), .B(n7700), .Z(n7702) );
  XNOR U1788 ( .A(n8055), .B(n7876), .Z(n7878) );
  XNOR U1789 ( .A(n8231), .B(n8052), .Z(n8054) );
  XNOR U1790 ( .A(n8407), .B(n8228), .Z(n8230) );
  XNOR U1791 ( .A(n8583), .B(n8404), .Z(n8406) );
  XNOR U1792 ( .A(n8759), .B(n8580), .Z(n8582) );
  XNOR U1793 ( .A(n8935), .B(n8756), .Z(n8758) );
  XNOR U1794 ( .A(n9111), .B(n8932), .Z(n8934) );
  XNOR U1795 ( .A(n9287), .B(n9108), .Z(n9110) );
  XNOR U1796 ( .A(n9463), .B(n9284), .Z(n9286) );
  XNOR U1797 ( .A(n9639), .B(n9460), .Z(n9462) );
  XNOR U1798 ( .A(n9815), .B(n9636), .Z(n9638) );
  XNOR U1799 ( .A(n9991), .B(n9812), .Z(n9814) );
  XNOR U1800 ( .A(n10167), .B(n9988), .Z(n9990) );
  XNOR U1801 ( .A(n10690), .B(n10712), .Z(n10694) );
  XNOR U1802 ( .A(n11077), .B(n11097), .Z(n11081) );
  XNOR U1803 ( .A(n11254), .B(n11274), .Z(n11258) );
  XNOR U1804 ( .A(n11431), .B(n11451), .Z(n11435) );
  XNOR U1805 ( .A(n11607), .B(n11627), .Z(n11611) );
  XNOR U1806 ( .A(n11783), .B(n11803), .Z(n11787) );
  XNOR U1807 ( .A(n12141), .B(n11962), .Z(n11964) );
  XNOR U1808 ( .A(n12317), .B(n12138), .Z(n12140) );
  XNOR U1809 ( .A(n12493), .B(n12314), .Z(n12316) );
  XNOR U1810 ( .A(n12669), .B(n12490), .Z(n12492) );
  XNOR U1811 ( .A(n12845), .B(n12666), .Z(n12668) );
  XNOR U1812 ( .A(n13021), .B(n12842), .Z(n12844) );
  XNOR U1813 ( .A(n13197), .B(n13018), .Z(n13020) );
  XNOR U1814 ( .A(n13373), .B(n13194), .Z(n13196) );
  XNOR U1815 ( .A(n13549), .B(n13370), .Z(n13372) );
  XNOR U1816 ( .A(n13725), .B(n13546), .Z(n13548) );
  XNOR U1817 ( .A(n13901), .B(n13722), .Z(n13724) );
  XNOR U1818 ( .A(n14077), .B(n13898), .Z(n13900) );
  XNOR U1819 ( .A(n14253), .B(n14074), .Z(n14076) );
  XNOR U1820 ( .A(n14429), .B(n14250), .Z(n14252) );
  XNOR U1821 ( .A(n14605), .B(n14426), .Z(n14428) );
  XNOR U1822 ( .A(n14781), .B(n14602), .Z(n14604) );
  XNOR U1823 ( .A(n14957), .B(n14778), .Z(n14780) );
  XNOR U1824 ( .A(n15133), .B(n14954), .Z(n14956) );
  XNOR U1825 ( .A(n15309), .B(n15130), .Z(n15132) );
  XNOR U1826 ( .A(n15485), .B(n15306), .Z(n15308) );
  XNOR U1827 ( .A(n15661), .B(n15482), .Z(n15484) );
  XNOR U1828 ( .A(n15650), .B(n15675), .Z(n15659) );
  XNOR U1829 ( .A(n16183), .B(n16202), .Z(n16188) );
  XNOR U1830 ( .A(n16558), .B(n16578), .Z(n16562) );
  XNOR U1831 ( .A(n16735), .B(n16755), .Z(n16739) );
  XNOR U1832 ( .A(n16912), .B(n16932), .Z(n16916) );
  XNOR U1833 ( .A(n17088), .B(n17108), .Z(n17092) );
  XNOR U1834 ( .A(n10524), .B(n10345), .Z(n10347) );
  XNOR U1835 ( .A(n10523), .B(n10533), .Z(n10517) );
  XOR U1836 ( .A(n5770), .B(n5777), .Z(n5774) );
  AND U1837 ( .A(n738), .B(n739), .Z(n557) );
  AND U1838 ( .A(n1460), .B(n1461), .Z(n1279) );
  AND U1839 ( .A(n2182), .B(n2183), .Z(n2001) );
  ANDN U1840 ( .B(n3264), .A(n3265), .Z(n3084) );
  ANDN U1841 ( .B(n3984), .A(n3985), .Z(n3804) );
  XNOR U1842 ( .A(n4524), .B(n4526), .Z(n4525) );
  NANDN U1843 ( .A(n4), .B(n3), .Z(n1) );
  XNOR U1844 ( .A(n17499), .B(n17670), .Z(n17504) );
  XNOR U1845 ( .A(n4388), .B(n4557), .Z(n4393) );
  XNOR U1846 ( .A(n6345), .B(n6510), .Z(n6350) );
  XNOR U1847 ( .A(n6873), .B(n7038), .Z(n6878) );
  XNOR U1848 ( .A(n7225), .B(n7390), .Z(n7230) );
  XNOR U1849 ( .A(n9337), .B(n9502), .Z(n9342) );
  XNOR U1850 ( .A(n9689), .B(n9854), .Z(n9694) );
  XNOR U1851 ( .A(n10041), .B(n10206), .Z(n10046) );
  XNOR U1852 ( .A(n10393), .B(n10558), .Z(n10398) );
  XNOR U1853 ( .A(n10747), .B(n10943), .Z(n10752) );
  XNOR U1854 ( .A(n11140), .B(n10960), .Z(n10962) );
  XNOR U1855 ( .A(n11317), .B(n11137), .Z(n11139) );
  XNOR U1856 ( .A(n11493), .B(n11314), .Z(n11315) );
  XNOR U1857 ( .A(n11663), .B(n11828), .Z(n11672) );
  XNOR U1858 ( .A(n12015), .B(n12180), .Z(n12020) );
  XNOR U1859 ( .A(n12367), .B(n12532), .Z(n12372) );
  XNOR U1860 ( .A(n12719), .B(n12884), .Z(n12724) );
  XNOR U1861 ( .A(n16237), .B(n16424), .Z(n16242) );
  XNOR U1862 ( .A(n16621), .B(n16441), .Z(n16443) );
  XNOR U1863 ( .A(n16798), .B(n16618), .Z(n16620) );
  XNOR U1864 ( .A(n16974), .B(n16795), .Z(n16796) );
  XNOR U1865 ( .A(n17144), .B(n17304), .Z(n17153) );
  XNOR U1866 ( .A(n1871), .B(n2033), .Z(n1875) );
  XNOR U1867 ( .A(n2232), .B(n2394), .Z(n2236) );
  XNOR U1868 ( .A(n2593), .B(n2755), .Z(n2597) );
  XNOR U1869 ( .A(n2954), .B(n3116), .Z(n2958) );
  XNOR U1870 ( .A(n3314), .B(n3476), .Z(n3318) );
  XNOR U1871 ( .A(n3674), .B(n3836), .Z(n3678) );
  XNOR U1872 ( .A(n4754), .B(n4916), .Z(n4758) );
  XNOR U1873 ( .A(n5651), .B(n5472), .Z(n5474) );
  XNOR U1874 ( .A(n5828), .B(n5648), .Z(n5650) );
  XNOR U1875 ( .A(n5821), .B(n5980), .Z(n5826) );
  XNOR U1876 ( .A(n6179), .B(n6333), .Z(n6174) );
  XNOR U1877 ( .A(n7583), .B(n7741), .Z(n7587) );
  XNOR U1878 ( .A(n7935), .B(n8093), .Z(n7939) );
  XNOR U1879 ( .A(n4039), .B(n4195), .Z(n4043) );
  XNOR U1880 ( .A(n8292), .B(n8444), .Z(n8296) );
  XNOR U1881 ( .A(n8644), .B(n8796), .Z(n8648) );
  XNOR U1882 ( .A(n8996), .B(n9148), .Z(n9000) );
  XNOR U1883 ( .A(n13434), .B(n13586), .Z(n13438) );
  XNOR U1884 ( .A(n13786), .B(n13938), .Z(n13790) );
  XNOR U1885 ( .A(n14138), .B(n14290), .Z(n14142) );
  XNOR U1886 ( .A(n14490), .B(n14642), .Z(n14494) );
  XNOR U1887 ( .A(n14842), .B(n14994), .Z(n14846) );
  XNOR U1888 ( .A(n15194), .B(n15346), .Z(n15198) );
  XNOR U1889 ( .A(n15546), .B(n15698), .Z(n15550) );
  XNOR U1890 ( .A(n15898), .B(n16049), .Z(n15902) );
  XNOR U1891 ( .A(n18190), .B(n18342), .Z(n18194) );
  XNOR U1892 ( .A(n17866), .B(n18018), .Z(n17870) );
  XNOR U1893 ( .A(n17515), .B(n17667), .Z(n17519) );
  XNOR U1894 ( .A(n1510), .B(n1672), .Z(n1514) );
  XNOR U1895 ( .A(n4404), .B(n4554), .Z(n4408) );
  XNOR U1896 ( .A(n6713), .B(n6859), .Z(n6721) );
  XNOR U1897 ( .A(n7241), .B(n7387), .Z(n7245) );
  XNOR U1898 ( .A(n9353), .B(n9499), .Z(n9357) );
  XNOR U1899 ( .A(n9705), .B(n9851), .Z(n9709) );
  XNOR U1900 ( .A(n10057), .B(n10203), .Z(n10061) );
  XNOR U1901 ( .A(n10409), .B(n10555), .Z(n10413) );
  XNOR U1902 ( .A(n10763), .B(n10937), .Z(n10767) );
  XNOR U1903 ( .A(n11155), .B(n10975), .Z(n10977) );
  XNOR U1904 ( .A(n11149), .B(n11295), .Z(n11153) );
  XNOR U1905 ( .A(n11326), .B(n11472), .Z(n11330) );
  XNOR U1906 ( .A(n11502), .B(n11648), .Z(n11506) );
  XNOR U1907 ( .A(n11678), .B(n11824), .Z(n11682) );
  XNOR U1908 ( .A(n12036), .B(n11857), .Z(n11859) );
  XNOR U1909 ( .A(n12035), .B(n12177), .Z(n12030) );
  XNOR U1910 ( .A(n12383), .B(n12529), .Z(n12387) );
  XNOR U1911 ( .A(n12735), .B(n12881), .Z(n12739) );
  XNOR U1912 ( .A(n13087), .B(n13233), .Z(n13091) );
  XNOR U1913 ( .A(n16253), .B(n16418), .Z(n16257) );
  XNOR U1914 ( .A(n16636), .B(n16456), .Z(n16458) );
  XNOR U1915 ( .A(n16813), .B(n16633), .Z(n16635) );
  XNOR U1916 ( .A(n16989), .B(n16810), .Z(n16812) );
  XNOR U1917 ( .A(n17165), .B(n16986), .Z(n16988) );
  XNOR U1918 ( .A(n17159), .B(n17300), .Z(n17163) );
  XNOR U1919 ( .A(n2247), .B(n2391), .Z(n2251) );
  XNOR U1920 ( .A(n2608), .B(n2752), .Z(n2612) );
  XNOR U1921 ( .A(n2969), .B(n3113), .Z(n2973) );
  XNOR U1922 ( .A(n3329), .B(n3473), .Z(n3333) );
  XNOR U1923 ( .A(n3689), .B(n3833), .Z(n3693) );
  XNOR U1924 ( .A(n4769), .B(n4913), .Z(n4773) );
  XNOR U1925 ( .A(n5666), .B(n5487), .Z(n5489) );
  XNOR U1926 ( .A(n5843), .B(n5663), .Z(n5665) );
  XNOR U1927 ( .A(n5837), .B(n5977), .Z(n5841) );
  XNOR U1928 ( .A(n6013), .B(n6153), .Z(n6017) );
  XNOR U1929 ( .A(n6189), .B(n6329), .Z(n6193) );
  XNOR U1930 ( .A(n6365), .B(n6505), .Z(n6369) );
  XNOR U1931 ( .A(n6536), .B(n6681), .Z(n6545) );
  XNOR U1932 ( .A(n7070), .B(n7210), .Z(n7074) );
  XNOR U1933 ( .A(n7598), .B(n7738), .Z(n7602) );
  XNOR U1934 ( .A(n7950), .B(n8090), .Z(n7954) );
  XNOR U1935 ( .A(n2071), .B(n2210), .Z(n2075) );
  XNOR U1936 ( .A(n4054), .B(n4192), .Z(n4058) );
  XNOR U1937 ( .A(n8307), .B(n8441), .Z(n8311) );
  XNOR U1938 ( .A(n8659), .B(n8793), .Z(n8663) );
  XNOR U1939 ( .A(n9011), .B(n9145), .Z(n9015) );
  XNOR U1940 ( .A(n13801), .B(n13935), .Z(n13805) );
  XNOR U1941 ( .A(n14153), .B(n14287), .Z(n14157) );
  XNOR U1942 ( .A(n14505), .B(n14639), .Z(n14509) );
  XNOR U1943 ( .A(n14857), .B(n14991), .Z(n14861) );
  XNOR U1944 ( .A(n15209), .B(n15343), .Z(n15213) );
  XNOR U1945 ( .A(n15561), .B(n15695), .Z(n15565) );
  XNOR U1946 ( .A(n15913), .B(n16046), .Z(n15917) );
  XNOR U1947 ( .A(n18505), .B(n18639), .Z(n18509) );
  XNOR U1948 ( .A(n18205), .B(n18339), .Z(n18209) );
  XNOR U1949 ( .A(n17881), .B(n18015), .Z(n17885) );
  XNOR U1950 ( .A(n17530), .B(n17664), .Z(n17534) );
  XNOR U1951 ( .A(n1525), .B(n1669), .Z(n1529) );
  XNOR U1952 ( .A(n1143), .B(n1312), .Z(n1148) );
  XNOR U1953 ( .A(n4419), .B(n4551), .Z(n4423) );
  XNOR U1954 ( .A(n9368), .B(n9496), .Z(n9372) );
  XNOR U1955 ( .A(n9720), .B(n9848), .Z(n9724) );
  XNOR U1956 ( .A(n10072), .B(n10200), .Z(n10076) );
  XNOR U1957 ( .A(n10424), .B(n10552), .Z(n10428) );
  XNOR U1958 ( .A(n10778), .B(n10931), .Z(n10782) );
  XNOR U1959 ( .A(n10987), .B(n11115), .Z(n10991) );
  XNOR U1960 ( .A(n11164), .B(n11292), .Z(n11168) );
  XNOR U1961 ( .A(n11341), .B(n11469), .Z(n11345) );
  XNOR U1962 ( .A(n11517), .B(n11645), .Z(n11521) );
  XNOR U1963 ( .A(n11693), .B(n11821), .Z(n11697) );
  XNOR U1964 ( .A(n11869), .B(n11997), .Z(n11873) );
  XNOR U1965 ( .A(n12045), .B(n12173), .Z(n12049) );
  XNOR U1966 ( .A(n12221), .B(n12349), .Z(n12225) );
  XNOR U1967 ( .A(n12392), .B(n12525), .Z(n12401) );
  XNOR U1968 ( .A(n12750), .B(n12878), .Z(n12758) );
  XNOR U1969 ( .A(n13102), .B(n13230), .Z(n13106) );
  XNOR U1970 ( .A(n13454), .B(n13582), .Z(n13458) );
  XNOR U1971 ( .A(n16268), .B(n16412), .Z(n16272) );
  XNOR U1972 ( .A(n16651), .B(n16471), .Z(n16473) );
  XNOR U1973 ( .A(n16828), .B(n16648), .Z(n16650) );
  XNOR U1974 ( .A(n17004), .B(n16825), .Z(n16827) );
  XNOR U1975 ( .A(n17180), .B(n17001), .Z(n17003) );
  XNOR U1976 ( .A(n17174), .B(n17297), .Z(n17178) );
  XNOR U1977 ( .A(n2623), .B(n2749), .Z(n2627) );
  XNOR U1978 ( .A(n2984), .B(n3110), .Z(n2988) );
  XNOR U1979 ( .A(n3344), .B(n3470), .Z(n3348) );
  XNOR U1980 ( .A(n3704), .B(n3830), .Z(n3708) );
  XNOR U1981 ( .A(n4784), .B(n4910), .Z(n4788) );
  XNOR U1982 ( .A(n5681), .B(n5502), .Z(n5504) );
  XNOR U1983 ( .A(n5858), .B(n5678), .Z(n5680) );
  XNOR U1984 ( .A(n5852), .B(n5974), .Z(n5856) );
  XNOR U1985 ( .A(n6028), .B(n6150), .Z(n6032) );
  XNOR U1986 ( .A(n6204), .B(n6326), .Z(n6208) );
  XNOR U1987 ( .A(n6380), .B(n6502), .Z(n6384) );
  XNOR U1988 ( .A(n6556), .B(n6678), .Z(n6560) );
  XNOR U1989 ( .A(n6732), .B(n6854), .Z(n6736) );
  XNOR U1990 ( .A(n6908), .B(n7030), .Z(n6912) );
  XNOR U1991 ( .A(n7079), .B(n7206), .Z(n7088) );
  XNOR U1992 ( .A(n7437), .B(n7559), .Z(n7445) );
  XNOR U1993 ( .A(n7789), .B(n7911), .Z(n7793) );
  XNOR U1994 ( .A(n2086), .B(n2207), .Z(n2090) );
  XNOR U1995 ( .A(n2447), .B(n2568), .Z(n2451) );
  XNOR U1996 ( .A(n4069), .B(n4189), .Z(n4073) );
  XNOR U1997 ( .A(n8146), .B(n8262), .Z(n8150) );
  XNOR U1998 ( .A(n8674), .B(n8790), .Z(n8678) );
  XNOR U1999 ( .A(n9026), .B(n9142), .Z(n9030) );
  XNOR U2000 ( .A(n14168), .B(n14284), .Z(n14172) );
  XNOR U2001 ( .A(n14520), .B(n14636), .Z(n14524) );
  XNOR U2002 ( .A(n14872), .B(n14988), .Z(n14876) );
  XNOR U2003 ( .A(n15224), .B(n15340), .Z(n15228) );
  XNOR U2004 ( .A(n15576), .B(n15692), .Z(n15580) );
  XNOR U2005 ( .A(n15928), .B(n16043), .Z(n15932) );
  XNOR U2006 ( .A(n19048), .B(n19164), .Z(n19052) );
  XNOR U2007 ( .A(n18796), .B(n18912), .Z(n18800) );
  XNOR U2008 ( .A(n18520), .B(n18636), .Z(n18524) );
  XNOR U2009 ( .A(n18220), .B(n18336), .Z(n18224) );
  XNOR U2010 ( .A(n17896), .B(n18012), .Z(n17900) );
  XNOR U2011 ( .A(n17545), .B(n17661), .Z(n17549) );
  XNOR U2012 ( .A(n1349), .B(n1488), .Z(n1353) );
  XNOR U2013 ( .A(n968), .B(n1131), .Z(n972) );
  XNOR U2014 ( .A(n4434), .B(n4548), .Z(n4438) );
  XNOR U2015 ( .A(n8503), .B(n8613), .Z(n8507) );
  XNOR U2016 ( .A(n9383), .B(n9493), .Z(n9387) );
  XNOR U2017 ( .A(n9735), .B(n9845), .Z(n9739) );
  XNOR U2018 ( .A(n10087), .B(n10197), .Z(n10091) );
  XNOR U2019 ( .A(n10439), .B(n10549), .Z(n10443) );
  XNOR U2020 ( .A(n10793), .B(n10925), .Z(n10797) );
  XNOR U2021 ( .A(n11002), .B(n11112), .Z(n11006) );
  XNOR U2022 ( .A(n11179), .B(n11289), .Z(n11183) );
  XNOR U2023 ( .A(n11356), .B(n11466), .Z(n11360) );
  XNOR U2024 ( .A(n11532), .B(n11642), .Z(n11536) );
  XNOR U2025 ( .A(n11708), .B(n11818), .Z(n11712) );
  XNOR U2026 ( .A(n11884), .B(n11994), .Z(n11888) );
  XNOR U2027 ( .A(n12060), .B(n12170), .Z(n12064) );
  XNOR U2028 ( .A(n12236), .B(n12346), .Z(n12240) );
  XNOR U2029 ( .A(n12412), .B(n12522), .Z(n12416) );
  XNOR U2030 ( .A(n12588), .B(n12698), .Z(n12592) );
  XNOR U2031 ( .A(n12764), .B(n12874), .Z(n12768) );
  XNOR U2032 ( .A(n13122), .B(n12943), .Z(n12945) );
  XNOR U2033 ( .A(n13121), .B(n13227), .Z(n13116) );
  XNOR U2034 ( .A(n13469), .B(n13579), .Z(n13473) );
  XNOR U2035 ( .A(n13821), .B(n13931), .Z(n13825) );
  XNOR U2036 ( .A(n16283), .B(n16406), .Z(n16287) );
  XNOR U2037 ( .A(n16666), .B(n16486), .Z(n16488) );
  XNOR U2038 ( .A(n16843), .B(n16663), .Z(n16665) );
  XNOR U2039 ( .A(n17019), .B(n16840), .Z(n16842) );
  XNOR U2040 ( .A(n17195), .B(n17016), .Z(n17018) );
  XNOR U2041 ( .A(n17189), .B(n17294), .Z(n17193) );
  XNOR U2042 ( .A(n1735), .B(n1844), .Z(n1739) );
  XNOR U2043 ( .A(n2999), .B(n3107), .Z(n3003) );
  XNOR U2044 ( .A(n3359), .B(n3467), .Z(n3363) );
  XNOR U2045 ( .A(n3719), .B(n3827), .Z(n3723) );
  XNOR U2046 ( .A(n4799), .B(n4907), .Z(n4803) );
  XNOR U2047 ( .A(n5696), .B(n5517), .Z(n5519) );
  XNOR U2048 ( .A(n5873), .B(n5693), .Z(n5695) );
  XNOR U2049 ( .A(n5867), .B(n5971), .Z(n5871) );
  XNOR U2050 ( .A(n6043), .B(n6147), .Z(n6047) );
  XNOR U2051 ( .A(n6219), .B(n6323), .Z(n6223) );
  XNOR U2052 ( .A(n6395), .B(n6499), .Z(n6399) );
  XNOR U2053 ( .A(n6571), .B(n6675), .Z(n6575) );
  XNOR U2054 ( .A(n6747), .B(n6851), .Z(n6751) );
  XNOR U2055 ( .A(n6923), .B(n7027), .Z(n6927) );
  XNOR U2056 ( .A(n7099), .B(n7203), .Z(n7103) );
  XNOR U2057 ( .A(n7275), .B(n7379), .Z(n7279) );
  XNOR U2058 ( .A(n7451), .B(n7555), .Z(n7455) );
  XNOR U2059 ( .A(n7622), .B(n7731), .Z(n7631) );
  XNOR U2060 ( .A(n7980), .B(n8084), .Z(n7988) );
  XNOR U2061 ( .A(n2101), .B(n2204), .Z(n2105) );
  XNOR U2062 ( .A(n2462), .B(n2565), .Z(n2466) );
  XNOR U2063 ( .A(n2823), .B(n2926), .Z(n2827) );
  XNOR U2064 ( .A(n4084), .B(n4186), .Z(n4088) );
  XNOR U2065 ( .A(n9041), .B(n9139), .Z(n9045) );
  XNOR U2066 ( .A(n14535), .B(n14633), .Z(n14539) );
  XNOR U2067 ( .A(n14887), .B(n14985), .Z(n14891) );
  XNOR U2068 ( .A(n15239), .B(n15337), .Z(n15243) );
  XNOR U2069 ( .A(n15591), .B(n15689), .Z(n15595) );
  XNOR U2070 ( .A(n15943), .B(n16040), .Z(n15947) );
  XNOR U2071 ( .A(n19291), .B(n19389), .Z(n19295) );
  XNOR U2072 ( .A(n19063), .B(n19161), .Z(n19067) );
  XNOR U2073 ( .A(n18811), .B(n18909), .Z(n18815) );
  XNOR U2074 ( .A(n18535), .B(n18633), .Z(n18539) );
  XNOR U2075 ( .A(n18235), .B(n18333), .Z(n18239) );
  XNOR U2076 ( .A(n17911), .B(n18009), .Z(n17915) );
  XNOR U2077 ( .A(n17560), .B(n17658), .Z(n17564) );
  XNOR U2078 ( .A(n983), .B(n1128), .Z(n987) );
  XNOR U2079 ( .A(n601), .B(n771), .Z(n606) );
  XNOR U2080 ( .A(n1384), .B(n1481), .Z(n1388) );
  XNOR U2081 ( .A(n4449), .B(n4545), .Z(n4453) );
  XNOR U2082 ( .A(n8518), .B(n8610), .Z(n8522) );
  XNOR U2083 ( .A(n8870), .B(n8962), .Z(n8874) );
  XNOR U2084 ( .A(n9398), .B(n9490), .Z(n9402) );
  XNOR U2085 ( .A(n9750), .B(n9842), .Z(n9754) );
  XNOR U2086 ( .A(n10102), .B(n10194), .Z(n10106) );
  XNOR U2087 ( .A(n10454), .B(n10546), .Z(n10458) );
  XNOR U2088 ( .A(n10808), .B(n10919), .Z(n10812) );
  XNOR U2089 ( .A(n11200), .B(n11020), .Z(n11022) );
  XNOR U2090 ( .A(n11194), .B(n11286), .Z(n11198) );
  XNOR U2091 ( .A(n11371), .B(n11463), .Z(n11375) );
  XNOR U2092 ( .A(n11547), .B(n11639), .Z(n11551) );
  XNOR U2093 ( .A(n11723), .B(n11815), .Z(n11727) );
  XNOR U2094 ( .A(n11899), .B(n11991), .Z(n11903) );
  XNOR U2095 ( .A(n12075), .B(n12167), .Z(n12079) );
  XNOR U2096 ( .A(n12251), .B(n12343), .Z(n12255) );
  XNOR U2097 ( .A(n12427), .B(n12519), .Z(n12431) );
  XNOR U2098 ( .A(n12603), .B(n12695), .Z(n12607) );
  XNOR U2099 ( .A(n12779), .B(n12871), .Z(n12783) );
  XNOR U2100 ( .A(n12955), .B(n13047), .Z(n12959) );
  XNOR U2101 ( .A(n13131), .B(n13223), .Z(n13135) );
  XNOR U2102 ( .A(n13307), .B(n13399), .Z(n13311) );
  XNOR U2103 ( .A(n13478), .B(n13575), .Z(n13487) );
  XNOR U2104 ( .A(n13836), .B(n13928), .Z(n13844) );
  XNOR U2105 ( .A(n14188), .B(n14280), .Z(n14192) );
  XNOR U2106 ( .A(n16298), .B(n16400), .Z(n16302) );
  XNOR U2107 ( .A(n16681), .B(n16501), .Z(n16503) );
  XNOR U2108 ( .A(n16858), .B(n16678), .Z(n16680) );
  XNOR U2109 ( .A(n17034), .B(n16855), .Z(n16857) );
  XNOR U2110 ( .A(n17210), .B(n17031), .Z(n17033) );
  XNOR U2111 ( .A(n17204), .B(n17291), .Z(n17208) );
  XNOR U2112 ( .A(n1369), .B(n1484), .Z(n1373) );
  XNOR U2113 ( .A(n3374), .B(n3464), .Z(n3378) );
  XNOR U2114 ( .A(n3734), .B(n3824), .Z(n3738) );
  XNOR U2115 ( .A(n4814), .B(n4904), .Z(n4818) );
  XNOR U2116 ( .A(n5711), .B(n5532), .Z(n5534) );
  XNOR U2117 ( .A(n5888), .B(n5708), .Z(n5710) );
  XNOR U2118 ( .A(n5882), .B(n5968), .Z(n5886) );
  XNOR U2119 ( .A(n6058), .B(n6144), .Z(n6062) );
  XNOR U2120 ( .A(n6234), .B(n6320), .Z(n6238) );
  XNOR U2121 ( .A(n6410), .B(n6496), .Z(n6414) );
  XNOR U2122 ( .A(n6586), .B(n6672), .Z(n6590) );
  XNOR U2123 ( .A(n6762), .B(n6848), .Z(n6766) );
  XNOR U2124 ( .A(n6938), .B(n7024), .Z(n6942) );
  XNOR U2125 ( .A(n7114), .B(n7200), .Z(n7118) );
  XNOR U2126 ( .A(n7290), .B(n7376), .Z(n7294) );
  XNOR U2127 ( .A(n7466), .B(n7552), .Z(n7470) );
  XNOR U2128 ( .A(n7642), .B(n7728), .Z(n7646) );
  XNOR U2129 ( .A(n7818), .B(n7904), .Z(n7822) );
  XNOR U2130 ( .A(n7994), .B(n8080), .Z(n7998) );
  XNOR U2131 ( .A(n8351), .B(n8433), .Z(n8346) );
  XNOR U2132 ( .A(n637), .B(n764), .Z(n641) );
  XNOR U2133 ( .A(n2116), .B(n2201), .Z(n2120) );
  XNOR U2134 ( .A(n2477), .B(n2562), .Z(n2481) );
  XNOR U2135 ( .A(n2838), .B(n2923), .Z(n2842) );
  XNOR U2136 ( .A(n3199), .B(n3283), .Z(n3203) );
  XNOR U2137 ( .A(n4099), .B(n4183), .Z(n4103) );
  XNOR U2138 ( .A(n14902), .B(n14982), .Z(n14906) );
  XNOR U2139 ( .A(n15254), .B(n15334), .Z(n15258) );
  XNOR U2140 ( .A(n15606), .B(n15686), .Z(n15610) );
  XNOR U2141 ( .A(n15958), .B(n16037), .Z(n15962) );
  XNOR U2142 ( .A(n19690), .B(n19770), .Z(n19694) );
  XNOR U2143 ( .A(n19510), .B(n19590), .Z(n19514) );
  XNOR U2144 ( .A(n19306), .B(n19386), .Z(n19310) );
  XNOR U2145 ( .A(n19078), .B(n19158), .Z(n19082) );
  XNOR U2146 ( .A(n18826), .B(n18906), .Z(n18830) );
  XNOR U2147 ( .A(n18550), .B(n18630), .Z(n18554) );
  XNOR U2148 ( .A(n18250), .B(n18330), .Z(n18254) );
  XNOR U2149 ( .A(n17926), .B(n18006), .Z(n17930) );
  XNOR U2150 ( .A(n17575), .B(n17655), .Z(n17579) );
  XNOR U2151 ( .A(n1023), .B(n1120), .Z(n1027) );
  XNOR U2152 ( .A(n808), .B(n946), .Z(n812) );
  XNOR U2153 ( .A(n427), .B(n589), .Z(n431) );
  XNOR U2154 ( .A(n1399), .B(n1478), .Z(n1403) );
  XNOR U2155 ( .A(n1760), .B(n1839), .Z(n1764) );
  XNOR U2156 ( .A(n4464), .B(n4542), .Z(n4468) );
  XNOR U2157 ( .A(n8885), .B(n8959), .Z(n8893) );
  XNOR U2158 ( .A(n9237), .B(n9311), .Z(n9241) );
  XNOR U2159 ( .A(n9765), .B(n9839), .Z(n9769) );
  XNOR U2160 ( .A(n10117), .B(n10191), .Z(n10121) );
  XNOR U2161 ( .A(n10469), .B(n10543), .Z(n10473) );
  XNOR U2162 ( .A(n10823), .B(n10913), .Z(n10827) );
  XNOR U2163 ( .A(n11215), .B(n11035), .Z(n11037) );
  XNOR U2164 ( .A(n11209), .B(n11283), .Z(n11213) );
  XNOR U2165 ( .A(n11386), .B(n11460), .Z(n11390) );
  XNOR U2166 ( .A(n11562), .B(n11636), .Z(n11566) );
  XNOR U2167 ( .A(n11738), .B(n11812), .Z(n11742) );
  XNOR U2168 ( .A(n11914), .B(n11988), .Z(n11918) );
  XNOR U2169 ( .A(n12090), .B(n12164), .Z(n12094) );
  XNOR U2170 ( .A(n12266), .B(n12340), .Z(n12270) );
  XNOR U2171 ( .A(n12442), .B(n12516), .Z(n12446) );
  XNOR U2172 ( .A(n12618), .B(n12692), .Z(n12622) );
  XNOR U2173 ( .A(n12794), .B(n12868), .Z(n12798) );
  XNOR U2174 ( .A(n12970), .B(n13044), .Z(n12974) );
  XNOR U2175 ( .A(n13146), .B(n13220), .Z(n13150) );
  XNOR U2176 ( .A(n13322), .B(n13396), .Z(n13326) );
  XNOR U2177 ( .A(n13498), .B(n13572), .Z(n13502) );
  XNOR U2178 ( .A(n13674), .B(n13748), .Z(n13678) );
  XNOR U2179 ( .A(n13850), .B(n13924), .Z(n13854) );
  XNOR U2180 ( .A(n14208), .B(n14029), .Z(n14031) );
  XNOR U2181 ( .A(n14207), .B(n14277), .Z(n14202) );
  XNOR U2182 ( .A(n14555), .B(n14629), .Z(n14559) );
  XNOR U2183 ( .A(n16313), .B(n16394), .Z(n16317) );
  XNOR U2184 ( .A(n16696), .B(n16516), .Z(n16518) );
  XNOR U2185 ( .A(n16873), .B(n16693), .Z(n16695) );
  XNOR U2186 ( .A(n17049), .B(n16870), .Z(n16872) );
  XNOR U2187 ( .A(n17225), .B(n17046), .Z(n17048) );
  XNOR U2188 ( .A(n17219), .B(n17288), .Z(n17223) );
  XNOR U2189 ( .A(n1003), .B(n1124), .Z(n1007) );
  XNOR U2190 ( .A(n858), .B(n936), .Z(n862) );
  XNOR U2191 ( .A(n3749), .B(n3821), .Z(n3753) );
  XNOR U2192 ( .A(n4829), .B(n4901), .Z(n4833) );
  XNOR U2193 ( .A(n5726), .B(n5547), .Z(n5549) );
  XNOR U2194 ( .A(n5903), .B(n5723), .Z(n5725) );
  XNOR U2195 ( .A(n5897), .B(n5965), .Z(n5901) );
  XNOR U2196 ( .A(n6073), .B(n6141), .Z(n6077) );
  XNOR U2197 ( .A(n6249), .B(n6317), .Z(n6253) );
  XNOR U2198 ( .A(n6425), .B(n6493), .Z(n6429) );
  XNOR U2199 ( .A(n6601), .B(n6669), .Z(n6605) );
  XNOR U2200 ( .A(n6777), .B(n6845), .Z(n6781) );
  XNOR U2201 ( .A(n6953), .B(n7021), .Z(n6957) );
  XNOR U2202 ( .A(n7129), .B(n7197), .Z(n7133) );
  XNOR U2203 ( .A(n7305), .B(n7373), .Z(n7309) );
  XNOR U2204 ( .A(n7481), .B(n7549), .Z(n7485) );
  XNOR U2205 ( .A(n7657), .B(n7725), .Z(n7661) );
  XNOR U2206 ( .A(n7833), .B(n7901), .Z(n7837) );
  XNOR U2207 ( .A(n8009), .B(n8077), .Z(n8013) );
  XNOR U2208 ( .A(n8185), .B(n8253), .Z(n8189) );
  XNOR U2209 ( .A(n8361), .B(n8429), .Z(n8365) );
  XNOR U2210 ( .A(n8537), .B(n8605), .Z(n8541) );
  XNOR U2211 ( .A(n8708), .B(n8781), .Z(n8717) );
  XNOR U2212 ( .A(n9594), .B(n9662), .Z(n9598) );
  XNOR U2213 ( .A(n462), .B(n582), .Z(n466) );
  XNOR U2214 ( .A(n2312), .B(n2378), .Z(n2316) );
  XNOR U2215 ( .A(n2673), .B(n2739), .Z(n2677) );
  XNOR U2216 ( .A(n3034), .B(n3100), .Z(n3038) );
  XNOR U2217 ( .A(n3394), .B(n3460), .Z(n3398) );
  XNOR U2218 ( .A(n4114), .B(n4180), .Z(n4118) );
  XNOR U2219 ( .A(n15269), .B(n15331), .Z(n15273) );
  XNOR U2220 ( .A(n15621), .B(n15683), .Z(n15625) );
  XNOR U2221 ( .A(n15973), .B(n16034), .Z(n15977) );
  XNOR U2222 ( .A(n19861), .B(n19923), .Z(n19865) );
  XNOR U2223 ( .A(n19705), .B(n19767), .Z(n19709) );
  XNOR U2224 ( .A(n19525), .B(n19587), .Z(n19529) );
  XNOR U2225 ( .A(n19321), .B(n19383), .Z(n19325) );
  XNOR U2226 ( .A(n19093), .B(n19155), .Z(n19097) );
  XNOR U2227 ( .A(n18841), .B(n18903), .Z(n18845) );
  XNOR U2228 ( .A(n18565), .B(n18627), .Z(n18569) );
  XNOR U2229 ( .A(n18265), .B(n18327), .Z(n18269) );
  XNOR U2230 ( .A(n17941), .B(n18003), .Z(n17945) );
  XNOR U2231 ( .A(n17590), .B(n17652), .Z(n17594) );
  XNOR U2232 ( .A(n657), .B(n760), .Z(n661) );
  XNOR U2233 ( .A(n442), .B(n586), .Z(n446) );
  XNOR U2234 ( .A(n512), .B(n572), .Z(n516) );
  XNOR U2235 ( .A(n1053), .B(n1114), .Z(n1057) );
  XNOR U2236 ( .A(n1414), .B(n1475), .Z(n1418) );
  XNOR U2237 ( .A(n1775), .B(n1836), .Z(n1779) );
  XNOR U2238 ( .A(n2136), .B(n2197), .Z(n2140) );
  XNOR U2239 ( .A(n4479), .B(n4539), .Z(n4483) );
  XNOR U2240 ( .A(n9428), .B(n9484), .Z(n9436) );
  XNOR U2241 ( .A(n10132), .B(n10188), .Z(n10136) );
  XNOR U2242 ( .A(n10484), .B(n10540), .Z(n10488) );
  XNOR U2243 ( .A(n10838), .B(n10907), .Z(n10842) );
  XNOR U2244 ( .A(n11047), .B(n11103), .Z(n11051) );
  XNOR U2245 ( .A(n11224), .B(n11280), .Z(n11228) );
  XNOR U2246 ( .A(n11401), .B(n11457), .Z(n11405) );
  XNOR U2247 ( .A(n11577), .B(n11633), .Z(n11581) );
  XNOR U2248 ( .A(n11753), .B(n11809), .Z(n11757) );
  XNOR U2249 ( .A(n11929), .B(n11985), .Z(n11933) );
  XNOR U2250 ( .A(n12105), .B(n12161), .Z(n12109) );
  XNOR U2251 ( .A(n12281), .B(n12337), .Z(n12285) );
  XNOR U2252 ( .A(n12457), .B(n12513), .Z(n12461) );
  XNOR U2253 ( .A(n12633), .B(n12689), .Z(n12637) );
  XNOR U2254 ( .A(n12809), .B(n12865), .Z(n12813) );
  XNOR U2255 ( .A(n12985), .B(n13041), .Z(n12989) );
  XNOR U2256 ( .A(n13161), .B(n13217), .Z(n13165) );
  XNOR U2257 ( .A(n13337), .B(n13393), .Z(n13341) );
  XNOR U2258 ( .A(n13513), .B(n13569), .Z(n13517) );
  XNOR U2259 ( .A(n13689), .B(n13745), .Z(n13693) );
  XNOR U2260 ( .A(n13865), .B(n13921), .Z(n13869) );
  XNOR U2261 ( .A(n14041), .B(n14097), .Z(n14045) );
  XNOR U2262 ( .A(n14217), .B(n14273), .Z(n14221) );
  XNOR U2263 ( .A(n14393), .B(n14449), .Z(n14397) );
  XNOR U2264 ( .A(n14564), .B(n14625), .Z(n14573) );
  XNOR U2265 ( .A(n14922), .B(n14978), .Z(n14930) );
  XNOR U2266 ( .A(n16328), .B(n16388), .Z(n16332) );
  XNOR U2267 ( .A(n16711), .B(n16531), .Z(n16533) );
  XNOR U2268 ( .A(n16888), .B(n16708), .Z(n16710) );
  XNOR U2269 ( .A(n17064), .B(n16885), .Z(n16887) );
  XNOR U2270 ( .A(n17240), .B(n17061), .Z(n17063) );
  XNOR U2271 ( .A(n17234), .B(n17285), .Z(n17238) );
  XNOR U2272 ( .A(n492), .B(n576), .Z(n496) );
  XNOR U2273 ( .A(n3944), .B(n3998), .Z(n3948) );
  XNOR U2274 ( .A(n4844), .B(n4898), .Z(n4848) );
  XNOR U2275 ( .A(n5741), .B(n5562), .Z(n5564) );
  XNOR U2276 ( .A(n5918), .B(n5738), .Z(n5740) );
  XNOR U2277 ( .A(n5912), .B(n5962), .Z(n5916) );
  XNOR U2278 ( .A(n6088), .B(n6138), .Z(n6092) );
  XNOR U2279 ( .A(n6264), .B(n6314), .Z(n6268) );
  XNOR U2280 ( .A(n6440), .B(n6490), .Z(n6444) );
  XNOR U2281 ( .A(n6616), .B(n6666), .Z(n6620) );
  XNOR U2282 ( .A(n6792), .B(n6842), .Z(n6796) );
  XNOR U2283 ( .A(n6968), .B(n7018), .Z(n6972) );
  XNOR U2284 ( .A(n7144), .B(n7194), .Z(n7148) );
  XNOR U2285 ( .A(n7320), .B(n7370), .Z(n7324) );
  XNOR U2286 ( .A(n7496), .B(n7546), .Z(n7500) );
  XNOR U2287 ( .A(n7672), .B(n7722), .Z(n7676) );
  XNOR U2288 ( .A(n7848), .B(n7898), .Z(n7852) );
  XNOR U2289 ( .A(n8024), .B(n8074), .Z(n8028) );
  XNOR U2290 ( .A(n8200), .B(n8250), .Z(n8204) );
  XNOR U2291 ( .A(n8376), .B(n8426), .Z(n8380) );
  XNOR U2292 ( .A(n8552), .B(n8602), .Z(n8556) );
  XNOR U2293 ( .A(n8728), .B(n8778), .Z(n8732) );
  XNOR U2294 ( .A(n8904), .B(n8954), .Z(n8908) );
  XNOR U2295 ( .A(n9080), .B(n9130), .Z(n9084) );
  XNOR U2296 ( .A(n9251), .B(n9306), .Z(n9260) );
  XNOR U2297 ( .A(n9785), .B(n9835), .Z(n9789) );
  XNOR U2298 ( .A(n687), .B(n754), .Z(n691) );
  XNOR U2299 ( .A(n2868), .B(n2917), .Z(n2872) );
  XNOR U2300 ( .A(n3229), .B(n3277), .Z(n3233) );
  XNOR U2301 ( .A(n3589), .B(n3637), .Z(n3593) );
  XNOR U2302 ( .A(n15636), .B(n15680), .Z(n15640) );
  XNOR U2303 ( .A(n15988), .B(n16031), .Z(n15992) );
  XNOR U2304 ( .A(n20116), .B(n20160), .Z(n20120) );
  XNOR U2305 ( .A(n20008), .B(n20052), .Z(n20012) );
  XNOR U2306 ( .A(n19876), .B(n19920), .Z(n19880) );
  XNOR U2307 ( .A(n19720), .B(n19764), .Z(n19724) );
  XNOR U2308 ( .A(n19540), .B(n19584), .Z(n19544) );
  XNOR U2309 ( .A(n19336), .B(n19380), .Z(n19340) );
  XNOR U2310 ( .A(n19108), .B(n19152), .Z(n19112) );
  XNOR U2311 ( .A(n18856), .B(n18900), .Z(n18860) );
  XNOR U2312 ( .A(n18580), .B(n18624), .Z(n18584) );
  XNOR U2313 ( .A(n18280), .B(n18324), .Z(n18284) );
  XNOR U2314 ( .A(n17956), .B(n18000), .Z(n17960) );
  XNOR U2315 ( .A(n17605), .B(n17649), .Z(n17609) );
  XNOR U2316 ( .A(n707), .B(n750), .Z(n711) );
  XNOR U2317 ( .A(n1068), .B(n1111), .Z(n1072) );
  XNOR U2318 ( .A(n1429), .B(n1472), .Z(n1433) );
  XNOR U2319 ( .A(n1790), .B(n1833), .Z(n1794) );
  XNOR U2320 ( .A(n2151), .B(n2194), .Z(n2155) );
  XNOR U2321 ( .A(n2512), .B(n2555), .Z(n2516) );
  XNOR U2322 ( .A(n4494), .B(n4536), .Z(n4498) );
  XNOR U2323 ( .A(n10499), .B(n10537), .Z(n10503) );
  XNOR U2324 ( .A(n10853), .B(n10901), .Z(n10857) );
  XNOR U2325 ( .A(n11245), .B(n11065), .Z(n11067) );
  XNOR U2326 ( .A(n11422), .B(n11242), .Z(n11244) );
  XNOR U2327 ( .A(n11416), .B(n11454), .Z(n11420) );
  XNOR U2328 ( .A(n11592), .B(n11630), .Z(n11596) );
  XNOR U2329 ( .A(n11768), .B(n11806), .Z(n11772) );
  XNOR U2330 ( .A(n11944), .B(n11982), .Z(n11948) );
  XNOR U2331 ( .A(n12120), .B(n12158), .Z(n12124) );
  XNOR U2332 ( .A(n12296), .B(n12334), .Z(n12300) );
  XNOR U2333 ( .A(n12472), .B(n12510), .Z(n12476) );
  XNOR U2334 ( .A(n12648), .B(n12686), .Z(n12652) );
  XNOR U2335 ( .A(n12824), .B(n12862), .Z(n12828) );
  XNOR U2336 ( .A(n13000), .B(n13038), .Z(n13004) );
  XNOR U2337 ( .A(n13176), .B(n13214), .Z(n13180) );
  XNOR U2338 ( .A(n13352), .B(n13390), .Z(n13356) );
  XNOR U2339 ( .A(n13528), .B(n13566), .Z(n13532) );
  XNOR U2340 ( .A(n13704), .B(n13742), .Z(n13708) );
  XNOR U2341 ( .A(n13880), .B(n13918), .Z(n13884) );
  XNOR U2342 ( .A(n14056), .B(n14094), .Z(n14060) );
  XNOR U2343 ( .A(n14232), .B(n14270), .Z(n14236) );
  XNOR U2344 ( .A(n14408), .B(n14446), .Z(n14412) );
  XNOR U2345 ( .A(n14584), .B(n14622), .Z(n14588) );
  XNOR U2346 ( .A(n14760), .B(n14798), .Z(n14764) );
  XNOR U2347 ( .A(n14936), .B(n14974), .Z(n14940) );
  XNOR U2348 ( .A(n15294), .B(n15115), .Z(n15117) );
  XNOR U2349 ( .A(n15293), .B(n15327), .Z(n15288) );
  XNOR U2350 ( .A(n16343), .B(n16382), .Z(n16347) );
  XNOR U2351 ( .A(n16726), .B(n16546), .Z(n16548) );
  XNOR U2352 ( .A(n16903), .B(n16723), .Z(n16725) );
  XNOR U2353 ( .A(n17079), .B(n16900), .Z(n16902) );
  XNOR U2354 ( .A(n17255), .B(n17076), .Z(n17078) );
  XNOR U2355 ( .A(n17249), .B(n17282), .Z(n17253) );
  XNOR U2356 ( .A(n4139), .B(n4175), .Z(n4143) );
  XNOR U2357 ( .A(n4859), .B(n4895), .Z(n4863) );
  XNOR U2358 ( .A(n5756), .B(n5577), .Z(n5579) );
  XNOR U2359 ( .A(n5933), .B(n5753), .Z(n5755) );
  XNOR U2360 ( .A(n5927), .B(n5959), .Z(n5931) );
  XNOR U2361 ( .A(n6103), .B(n6135), .Z(n6107) );
  XNOR U2362 ( .A(n6279), .B(n6311), .Z(n6283) );
  XNOR U2363 ( .A(n6455), .B(n6487), .Z(n6459) );
  XNOR U2364 ( .A(n6631), .B(n6663), .Z(n6635) );
  XNOR U2365 ( .A(n6807), .B(n6839), .Z(n6811) );
  XNOR U2366 ( .A(n6983), .B(n7015), .Z(n6987) );
  XNOR U2367 ( .A(n7159), .B(n7191), .Z(n7163) );
  XNOR U2368 ( .A(n7335), .B(n7367), .Z(n7339) );
  XNOR U2369 ( .A(n7511), .B(n7543), .Z(n7515) );
  XNOR U2370 ( .A(n7687), .B(n7719), .Z(n7691) );
  XNOR U2371 ( .A(n7863), .B(n7895), .Z(n7867) );
  XNOR U2372 ( .A(n8039), .B(n8071), .Z(n8043) );
  XNOR U2373 ( .A(n8215), .B(n8247), .Z(n8219) );
  XNOR U2374 ( .A(n8391), .B(n8423), .Z(n8395) );
  XNOR U2375 ( .A(n8567), .B(n8599), .Z(n8571) );
  XNOR U2376 ( .A(n8743), .B(n8775), .Z(n8747) );
  XNOR U2377 ( .A(n8919), .B(n8951), .Z(n8923) );
  XNOR U2378 ( .A(n9095), .B(n9127), .Z(n9099) );
  XNOR U2379 ( .A(n9271), .B(n9303), .Z(n9275) );
  XNOR U2380 ( .A(n9447), .B(n9479), .Z(n9451) );
  XNOR U2381 ( .A(n9623), .B(n9655), .Z(n9627) );
  XNOR U2382 ( .A(n9794), .B(n9831), .Z(n9803) );
  XNOR U2383 ( .A(n10152), .B(n10184), .Z(n10160) );
  XNOR U2384 ( .A(n16003), .B(n16028), .Z(n16007) );
  XNOR U2385 ( .A(n20215), .B(n20241), .Z(n20219) );
  XNOR U2386 ( .A(n20131), .B(n20157), .Z(n20135) );
  XNOR U2387 ( .A(n20023), .B(n20049), .Z(n20027) );
  XNOR U2388 ( .A(n19891), .B(n19917), .Z(n19895) );
  XNOR U2389 ( .A(n19735), .B(n19761), .Z(n19739) );
  XNOR U2390 ( .A(n19555), .B(n19581), .Z(n19559) );
  XNOR U2391 ( .A(n19351), .B(n19377), .Z(n19355) );
  XNOR U2392 ( .A(n19123), .B(n19149), .Z(n19127) );
  XNOR U2393 ( .A(n18871), .B(n18897), .Z(n18875) );
  XNOR U2394 ( .A(n18595), .B(n18621), .Z(n18599) );
  XNOR U2395 ( .A(n18295), .B(n18321), .Z(n18299) );
  XNOR U2396 ( .A(n17971), .B(n17997), .Z(n17975) );
  XNOR U2397 ( .A(n17620), .B(n17646), .Z(n17624) );
  XNOR U2398 ( .A(n722), .B(n747), .Z(n726) );
  XNOR U2399 ( .A(n1083), .B(n1108), .Z(n1087) );
  XNOR U2400 ( .A(n1444), .B(n1469), .Z(n1448) );
  XNOR U2401 ( .A(n1805), .B(n1830), .Z(n1809) );
  XNOR U2402 ( .A(n2166), .B(n2191), .Z(n2170) );
  XNOR U2403 ( .A(n2527), .B(n2552), .Z(n2531) );
  XNOR U2404 ( .A(n2888), .B(n2913), .Z(n2892) );
  XNOR U2405 ( .A(n3429), .B(n3453), .Z(n3433) );
  XNOR U2406 ( .A(n3969), .B(n3993), .Z(n3973) );
  XNOR U2407 ( .A(n4689), .B(n4713), .Z(n4693) );
  XNOR U2408 ( .A(n10868), .B(n10895), .Z(n10872) );
  XNOR U2409 ( .A(n11260), .B(n11080), .Z(n11082) );
  XNOR U2410 ( .A(n11437), .B(n11257), .Z(n11259) );
  XNOR U2411 ( .A(n11613), .B(n11434), .Z(n11436) );
  XNOR U2412 ( .A(n11789), .B(n11610), .Z(n11612) );
  XNOR U2413 ( .A(n11965), .B(n11786), .Z(n11788) );
  XNOR U2414 ( .A(n11959), .B(n11979), .Z(n11963) );
  XNOR U2415 ( .A(n12135), .B(n12155), .Z(n12139) );
  XNOR U2416 ( .A(n12311), .B(n12331), .Z(n12315) );
  XNOR U2417 ( .A(n12487), .B(n12507), .Z(n12491) );
  XNOR U2418 ( .A(n12663), .B(n12683), .Z(n12667) );
  XNOR U2419 ( .A(n12839), .B(n12859), .Z(n12843) );
  XNOR U2420 ( .A(n13015), .B(n13035), .Z(n13019) );
  XNOR U2421 ( .A(n13191), .B(n13211), .Z(n13195) );
  XNOR U2422 ( .A(n13367), .B(n13387), .Z(n13371) );
  XNOR U2423 ( .A(n13543), .B(n13563), .Z(n13547) );
  XNOR U2424 ( .A(n13719), .B(n13739), .Z(n13723) );
  XNOR U2425 ( .A(n13895), .B(n13915), .Z(n13899) );
  XNOR U2426 ( .A(n14071), .B(n14091), .Z(n14075) );
  XNOR U2427 ( .A(n14247), .B(n14267), .Z(n14251) );
  XNOR U2428 ( .A(n14423), .B(n14443), .Z(n14427) );
  XNOR U2429 ( .A(n14599), .B(n14619), .Z(n14603) );
  XNOR U2430 ( .A(n14775), .B(n14795), .Z(n14779) );
  XNOR U2431 ( .A(n14951), .B(n14971), .Z(n14955) );
  XNOR U2432 ( .A(n15127), .B(n15147), .Z(n15131) );
  XNOR U2433 ( .A(n15303), .B(n15323), .Z(n15307) );
  XNOR U2434 ( .A(n15479), .B(n15499), .Z(n15483) );
  XNOR U2435 ( .A(n15837), .B(n15658), .Z(n15660) );
  XNOR U2436 ( .A(n15836), .B(n15852), .Z(n15831) );
  XNOR U2437 ( .A(n16358), .B(n16376), .Z(n16364) );
  XNOR U2438 ( .A(n16741), .B(n16561), .Z(n16563) );
  XNOR U2439 ( .A(n16918), .B(n16738), .Z(n16740) );
  XNOR U2440 ( .A(n17094), .B(n16915), .Z(n16917) );
  XNOR U2441 ( .A(n17270), .B(n17091), .Z(n17093) );
  XNOR U2442 ( .A(n17264), .B(n17279), .Z(n17268) );
  XNOR U2443 ( .A(n3254), .B(n3272), .Z(n3263) );
  XNOR U2444 ( .A(n3794), .B(n3812), .Z(n3803) );
  XNOR U2445 ( .A(n4334), .B(n4352), .Z(n4343) );
  XNOR U2446 ( .A(n5054), .B(n5400), .Z(n5062) );
  XNOR U2447 ( .A(n5589), .B(n5602), .Z(n5593) );
  XNOR U2448 ( .A(n5948), .B(n5768), .Z(n5770) );
  XNOR U2449 ( .A(n5942), .B(n5956), .Z(n5946) );
  XNOR U2450 ( .A(n6300), .B(n6121), .Z(n6123) );
  XNOR U2451 ( .A(n6476), .B(n6297), .Z(n6299) );
  XNOR U2452 ( .A(n6470), .B(n6484), .Z(n6474) );
  XNOR U2453 ( .A(n6828), .B(n6649), .Z(n6651) );
  XNOR U2454 ( .A(n7004), .B(n6825), .Z(n6827) );
  XNOR U2455 ( .A(n6998), .B(n7012), .Z(n7002) );
  XNOR U2456 ( .A(n7356), .B(n7177), .Z(n7179) );
  XNOR U2457 ( .A(n7532), .B(n7353), .Z(n7355) );
  XNOR U2458 ( .A(n7526), .B(n7540), .Z(n7530) );
  XNOR U2459 ( .A(n7884), .B(n7705), .Z(n7707) );
  XNOR U2460 ( .A(n8060), .B(n7881), .Z(n7883) );
  XNOR U2461 ( .A(n8054), .B(n8068), .Z(n8058) );
  XNOR U2462 ( .A(n8412), .B(n8233), .Z(n8235) );
  XNOR U2463 ( .A(n8588), .B(n8409), .Z(n8411) );
  XNOR U2464 ( .A(n8582), .B(n8596), .Z(n8586) );
  XNOR U2465 ( .A(n8940), .B(n8761), .Z(n8763) );
  XNOR U2466 ( .A(n9116), .B(n8937), .Z(n8939) );
  XNOR U2467 ( .A(n9110), .B(n9124), .Z(n9114) );
  XNOR U2468 ( .A(n9468), .B(n9289), .Z(n9291) );
  XNOR U2469 ( .A(n9644), .B(n9465), .Z(n9467) );
  XNOR U2470 ( .A(n9638), .B(n9652), .Z(n9642) );
  XNOR U2471 ( .A(n9996), .B(n9817), .Z(n9819) );
  XNOR U2472 ( .A(n10172), .B(n9993), .Z(n9995) );
  XNOR U2473 ( .A(n10166), .B(n10180), .Z(n10170) );
  XNOR U2474 ( .A(n10337), .B(n10356), .Z(n10346) );
  XNOR U2475 ( .A(n10695), .B(n10711), .Z(n10703) );
  NAND U2476 ( .A(n919), .B(n918), .Z(n737) );
  NAND U2477 ( .A(n1641), .B(n1640), .Z(n1459) );
  NAND U2478 ( .A(n2363), .B(n2362), .Z(n2181) );
  ANDN U2479 ( .B(n2904), .A(n2905), .Z(n2723) );
  XNOR U2480 ( .A(n3444), .B(n3446), .Z(n3445) );
  XNOR U2481 ( .A(n3984), .B(n3986), .Z(n3985) );
  XNOR U2482 ( .A(n4704), .B(n4706), .Z(n4705) );
  AND U2483 ( .A(n5), .B(n6), .Z(n3) );
  XNOR U2484 ( .A(n1865), .B(n2034), .Z(n1870) );
  XNOR U2485 ( .A(n4568), .B(n4737), .Z(n4573) );
  XNOR U2486 ( .A(n5997), .B(n6158), .Z(n5993) );
  XNOR U2487 ( .A(n7753), .B(n7918), .Z(n7758) );
  XNOR U2488 ( .A(n8105), .B(n8270), .Z(n8110) );
  XNOR U2489 ( .A(n9865), .B(n10030), .Z(n9870) );
  XNOR U2490 ( .A(n12895), .B(n13060), .Z(n12900) );
  XNOR U2491 ( .A(n13247), .B(n13412), .Z(n13252) );
  XNOR U2492 ( .A(n13599), .B(n13764), .Z(n13604) );
  XNOR U2493 ( .A(n13951), .B(n14116), .Z(n13956) );
  XNOR U2494 ( .A(n14303), .B(n14468), .Z(n14308) );
  XNOR U2495 ( .A(n14655), .B(n14820), .Z(n14660) );
  XNOR U2496 ( .A(n15007), .B(n15172), .Z(n15012) );
  XNOR U2497 ( .A(n15359), .B(n15524), .Z(n15364) );
  XNOR U2498 ( .A(n17685), .B(n17849), .Z(n17689) );
  XNOR U2499 ( .A(n17321), .B(n17487), .Z(n17329) );
  XNOR U2500 ( .A(n4934), .B(n5448), .Z(n4938) );
  XNOR U2501 ( .A(n5469), .B(n5626), .Z(n5473) );
  XNOR U2502 ( .A(n5645), .B(n5803), .Z(n5649) );
  XNOR U2503 ( .A(n6004), .B(n5825), .Z(n5827) );
  XNOR U2504 ( .A(n6180), .B(n6001), .Z(n6003) );
  XNOR U2505 ( .A(n6351), .B(n6509), .Z(n6359) );
  XNOR U2506 ( .A(n6703), .B(n6861), .Z(n6707) );
  XNOR U2507 ( .A(n8463), .B(n8621), .Z(n8467) );
  XNOR U2508 ( .A(n8815), .B(n8973), .Z(n8819) );
  XNOR U2509 ( .A(n9167), .B(n9325), .Z(n9171) );
  XNOR U2510 ( .A(n10223), .B(n10381), .Z(n10227) );
  XNOR U2511 ( .A(n10575), .B(n10735), .Z(n10579) );
  XNOR U2512 ( .A(n11145), .B(n10965), .Z(n10967) );
  XNOR U2513 ( .A(n11322), .B(n11142), .Z(n11144) );
  XNOR U2514 ( .A(n11498), .B(n11319), .Z(n11321) );
  XNOR U2515 ( .A(n11674), .B(n11495), .Z(n11497) );
  XNOR U2516 ( .A(n11673), .B(n11827), .Z(n11668) );
  XNOR U2517 ( .A(n12021), .B(n12179), .Z(n12025) );
  XNOR U2518 ( .A(n12373), .B(n12531), .Z(n12377) );
  XNOR U2519 ( .A(n12725), .B(n12883), .Z(n12729) );
  XNOR U2520 ( .A(n15717), .B(n15875), .Z(n15721) );
  XNOR U2521 ( .A(n16068), .B(n16225), .Z(n16072) );
  XNOR U2522 ( .A(n16443), .B(n16601), .Z(n16447) );
  XNOR U2523 ( .A(n16620), .B(n16778), .Z(n16624) );
  XNOR U2524 ( .A(n16796), .B(n16955), .Z(n16801) );
  XNOR U2525 ( .A(n16968), .B(n17131), .Z(n16977) );
  XNOR U2526 ( .A(n2417), .B(n2574), .Z(n2421) );
  XNOR U2527 ( .A(n2778), .B(n2935), .Z(n2782) );
  XNOR U2528 ( .A(n3139), .B(n3295), .Z(n3143) );
  XNOR U2529 ( .A(n3499), .B(n3655), .Z(n3503) );
  XNOR U2530 ( .A(n3859), .B(n4015), .Z(n3863) );
  XNOR U2531 ( .A(n4219), .B(n4375), .Z(n4223) );
  XNOR U2532 ( .A(n7060), .B(n7212), .Z(n7064) );
  XNOR U2533 ( .A(n7412), .B(n7564), .Z(n7416) );
  XNOR U2534 ( .A(n9524), .B(n9676), .Z(n9528) );
  XNOR U2535 ( .A(n1881), .B(n2031), .Z(n1885) );
  XNOR U2536 ( .A(n2242), .B(n2392), .Z(n2246) );
  XNOR U2537 ( .A(n4584), .B(n4734), .Z(n4588) );
  XNOR U2538 ( .A(n7769), .B(n7915), .Z(n7773) );
  XNOR U2539 ( .A(n8121), .B(n8267), .Z(n8125) );
  XNOR U2540 ( .A(n9881), .B(n10027), .Z(n9885) );
  XNOR U2541 ( .A(n13263), .B(n13409), .Z(n13267) );
  XNOR U2542 ( .A(n13615), .B(n13761), .Z(n13619) );
  XNOR U2543 ( .A(n13967), .B(n14113), .Z(n13971) );
  XNOR U2544 ( .A(n14319), .B(n14465), .Z(n14323) );
  XNOR U2545 ( .A(n14671), .B(n14817), .Z(n14675) );
  XNOR U2546 ( .A(n15023), .B(n15169), .Z(n15027) );
  XNOR U2547 ( .A(n15375), .B(n15521), .Z(n15379) );
  XNOR U2548 ( .A(n18348), .B(n18494), .Z(n18352) );
  XNOR U2549 ( .A(n18036), .B(n18182), .Z(n18040) );
  XNOR U2550 ( .A(n17700), .B(n17846), .Z(n17704) );
  XNOR U2551 ( .A(n17335), .B(n17484), .Z(n17339) );
  XNOR U2552 ( .A(n1323), .B(n1493), .Z(n1328) );
  XNOR U2553 ( .A(n4949), .B(n5442), .Z(n4953) );
  XNOR U2554 ( .A(n5484), .B(n5623), .Z(n5488) );
  XNOR U2555 ( .A(n5660), .B(n5800), .Z(n5664) );
  XNOR U2556 ( .A(n6019), .B(n5840), .Z(n5842) );
  XNOR U2557 ( .A(n6195), .B(n6016), .Z(n6018) );
  XNOR U2558 ( .A(n6371), .B(n6192), .Z(n6194) );
  XNOR U2559 ( .A(n6547), .B(n6368), .Z(n6370) );
  XNOR U2560 ( .A(n6723), .B(n6544), .Z(n6546) );
  XNOR U2561 ( .A(n6722), .B(n6858), .Z(n6717) );
  XNOR U2562 ( .A(n8478), .B(n8618), .Z(n8482) );
  XNOR U2563 ( .A(n8830), .B(n8970), .Z(n8834) );
  XNOR U2564 ( .A(n9182), .B(n9322), .Z(n9186) );
  XNOR U2565 ( .A(n10238), .B(n10378), .Z(n10242) );
  XNOR U2566 ( .A(n10590), .B(n10732), .Z(n10594) );
  XNOR U2567 ( .A(n10977), .B(n11117), .Z(n10981) );
  XNOR U2568 ( .A(n11154), .B(n11294), .Z(n11158) );
  XNOR U2569 ( .A(n11513), .B(n11334), .Z(n11336) );
  XNOR U2570 ( .A(n11689), .B(n11510), .Z(n11512) );
  XNOR U2571 ( .A(n11865), .B(n11686), .Z(n11688) );
  XNOR U2572 ( .A(n12041), .B(n11862), .Z(n11864) );
  XNOR U2573 ( .A(n12030), .B(n12175), .Z(n12039) );
  XNOR U2574 ( .A(n12388), .B(n12528), .Z(n12396) );
  XNOR U2575 ( .A(n12740), .B(n12880), .Z(n12744) );
  XNOR U2576 ( .A(n13092), .B(n13232), .Z(n13096) );
  XNOR U2577 ( .A(n15732), .B(n15872), .Z(n15736) );
  XNOR U2578 ( .A(n16083), .B(n16222), .Z(n16087) );
  XNOR U2579 ( .A(n16458), .B(n16598), .Z(n16462) );
  XNOR U2580 ( .A(n16635), .B(n16775), .Z(n16639) );
  XNOR U2581 ( .A(n16812), .B(n16952), .Z(n16816) );
  XNOR U2582 ( .A(n16988), .B(n17128), .Z(n16992) );
  XNOR U2583 ( .A(n2793), .B(n2932), .Z(n2797) );
  XNOR U2584 ( .A(n3154), .B(n3292), .Z(n3158) );
  XNOR U2585 ( .A(n3514), .B(n3652), .Z(n3518) );
  XNOR U2586 ( .A(n3874), .B(n4012), .Z(n3878) );
  XNOR U2587 ( .A(n4234), .B(n4372), .Z(n4238) );
  XNOR U2588 ( .A(n7075), .B(n7209), .Z(n7083) );
  XNOR U2589 ( .A(n7427), .B(n7561), .Z(n7431) );
  XNOR U2590 ( .A(n9539), .B(n9673), .Z(n9543) );
  XNOR U2591 ( .A(n1896), .B(n2028), .Z(n1900) );
  XNOR U2592 ( .A(n2257), .B(n2389), .Z(n2261) );
  XNOR U2593 ( .A(n2618), .B(n2750), .Z(n2622) );
  XNOR U2594 ( .A(n4599), .B(n4731), .Z(n4603) );
  XNOR U2595 ( .A(n7784), .B(n7912), .Z(n7788) );
  XNOR U2596 ( .A(n8136), .B(n8264), .Z(n8140) );
  XNOR U2597 ( .A(n9896), .B(n10024), .Z(n9900) );
  XNOR U2598 ( .A(n13630), .B(n13758), .Z(n13634) );
  XNOR U2599 ( .A(n13982), .B(n14110), .Z(n13986) );
  XNOR U2600 ( .A(n14334), .B(n14462), .Z(n14338) );
  XNOR U2601 ( .A(n14686), .B(n14814), .Z(n14690) );
  XNOR U2602 ( .A(n15038), .B(n15166), .Z(n15042) );
  XNOR U2603 ( .A(n15390), .B(n15518), .Z(n15394) );
  XNOR U2604 ( .A(n18651), .B(n18779), .Z(n18655) );
  XNOR U2605 ( .A(n18363), .B(n18491), .Z(n18367) );
  XNOR U2606 ( .A(n18051), .B(n18179), .Z(n18055) );
  XNOR U2607 ( .A(n17715), .B(n17843), .Z(n17719) );
  XNOR U2608 ( .A(n17350), .B(n17481), .Z(n17354) );
  XNOR U2609 ( .A(n1530), .B(n1668), .Z(n1534) );
  XNOR U2610 ( .A(n1149), .B(n1311), .Z(n1153) );
  XNOR U2611 ( .A(n4964), .B(n5436), .Z(n4968) );
  XNOR U2612 ( .A(n5499), .B(n5620), .Z(n5503) );
  XNOR U2613 ( .A(n5675), .B(n5797), .Z(n5679) );
  XNOR U2614 ( .A(n6034), .B(n5855), .Z(n5857) );
  XNOR U2615 ( .A(n6210), .B(n6031), .Z(n6033) );
  XNOR U2616 ( .A(n6386), .B(n6207), .Z(n6209) );
  XNOR U2617 ( .A(n6562), .B(n6383), .Z(n6385) );
  XNOR U2618 ( .A(n6738), .B(n6559), .Z(n6561) );
  XNOR U2619 ( .A(n6914), .B(n6735), .Z(n6737) );
  XNOR U2620 ( .A(n7090), .B(n6911), .Z(n6913) );
  XNOR U2621 ( .A(n7266), .B(n7087), .Z(n7089) );
  XNOR U2622 ( .A(n8493), .B(n8615), .Z(n8497) );
  XNOR U2623 ( .A(n8845), .B(n8967), .Z(n8849) );
  XNOR U2624 ( .A(n9197), .B(n9319), .Z(n9201) );
  XNOR U2625 ( .A(n10253), .B(n10375), .Z(n10257) );
  XNOR U2626 ( .A(n10605), .B(n10729), .Z(n10609) );
  XNOR U2627 ( .A(n11175), .B(n10995), .Z(n10997) );
  XNOR U2628 ( .A(n11352), .B(n11172), .Z(n11174) );
  XNOR U2629 ( .A(n11528), .B(n11349), .Z(n11351) );
  XNOR U2630 ( .A(n11704), .B(n11525), .Z(n11527) );
  XNOR U2631 ( .A(n11880), .B(n11701), .Z(n11703) );
  XNOR U2632 ( .A(n12056), .B(n11877), .Z(n11879) );
  XNOR U2633 ( .A(n12232), .B(n12053), .Z(n12055) );
  XNOR U2634 ( .A(n12408), .B(n12229), .Z(n12231) );
  XNOR U2635 ( .A(n12584), .B(n12405), .Z(n12407) );
  XNOR U2636 ( .A(n12760), .B(n12581), .Z(n12583) );
  XNOR U2637 ( .A(n12759), .B(n12877), .Z(n12754) );
  XNOR U2638 ( .A(n13107), .B(n13229), .Z(n13111) );
  XNOR U2639 ( .A(n13459), .B(n13581), .Z(n13463) );
  XNOR U2640 ( .A(n15747), .B(n15869), .Z(n15751) );
  XNOR U2641 ( .A(n16098), .B(n16219), .Z(n16102) );
  XNOR U2642 ( .A(n16473), .B(n16595), .Z(n16477) );
  XNOR U2643 ( .A(n16650), .B(n16772), .Z(n16654) );
  XNOR U2644 ( .A(n16827), .B(n16949), .Z(n16831) );
  XNOR U2645 ( .A(n17003), .B(n17125), .Z(n17007) );
  XNOR U2646 ( .A(n3169), .B(n3289), .Z(n3173) );
  XNOR U2647 ( .A(n3529), .B(n3649), .Z(n3533) );
  XNOR U2648 ( .A(n3889), .B(n4009), .Z(n3893) );
  XNOR U2649 ( .A(n4249), .B(n4369), .Z(n4253) );
  XNOR U2650 ( .A(n7446), .B(n7558), .Z(n7441) );
  XNOR U2651 ( .A(n9554), .B(n9670), .Z(n9558) );
  XNOR U2652 ( .A(n1911), .B(n2025), .Z(n1915) );
  XNOR U2653 ( .A(n2272), .B(n2386), .Z(n2276) );
  XNOR U2654 ( .A(n2633), .B(n2747), .Z(n2637) );
  XNOR U2655 ( .A(n2994), .B(n3108), .Z(n2998) );
  XNOR U2656 ( .A(n4614), .B(n4728), .Z(n4618) );
  XNOR U2657 ( .A(n7799), .B(n7909), .Z(n7807) );
  XNOR U2658 ( .A(n8151), .B(n8261), .Z(n8155) );
  XNOR U2659 ( .A(n9911), .B(n10021), .Z(n9915) );
  XNOR U2660 ( .A(n13997), .B(n14107), .Z(n14001) );
  XNOR U2661 ( .A(n14349), .B(n14459), .Z(n14353) );
  XNOR U2662 ( .A(n14701), .B(n14811), .Z(n14705) );
  XNOR U2663 ( .A(n15053), .B(n15163), .Z(n15057) );
  XNOR U2664 ( .A(n15405), .B(n15515), .Z(n15409) );
  XNOR U2665 ( .A(n19170), .B(n19280), .Z(n19174) );
  XNOR U2666 ( .A(n18930), .B(n19040), .Z(n18934) );
  XNOR U2667 ( .A(n18666), .B(n18776), .Z(n18670) );
  XNOR U2668 ( .A(n18378), .B(n18488), .Z(n18382) );
  XNOR U2669 ( .A(n18066), .B(n18176), .Z(n18070) );
  XNOR U2670 ( .A(n17730), .B(n17840), .Z(n17734) );
  XNOR U2671 ( .A(n17365), .B(n17478), .Z(n17369) );
  XNOR U2672 ( .A(n1164), .B(n1308), .Z(n1168) );
  XNOR U2673 ( .A(n782), .B(n951), .Z(n787) );
  XNOR U2674 ( .A(n4979), .B(n5430), .Z(n4983) );
  XNOR U2675 ( .A(n5514), .B(n5617), .Z(n5518) );
  XNOR U2676 ( .A(n5690), .B(n5794), .Z(n5694) );
  XNOR U2677 ( .A(n6049), .B(n5870), .Z(n5872) );
  XNOR U2678 ( .A(n6225), .B(n6046), .Z(n6048) );
  XNOR U2679 ( .A(n6401), .B(n6222), .Z(n6224) );
  XNOR U2680 ( .A(n6577), .B(n6398), .Z(n6400) );
  XNOR U2681 ( .A(n6753), .B(n6574), .Z(n6576) );
  XNOR U2682 ( .A(n6929), .B(n6750), .Z(n6752) );
  XNOR U2683 ( .A(n7105), .B(n6926), .Z(n6928) );
  XNOR U2684 ( .A(n7281), .B(n7102), .Z(n7104) );
  XNOR U2685 ( .A(n7457), .B(n7278), .Z(n7280) );
  XNOR U2686 ( .A(n7633), .B(n7454), .Z(n7456) );
  XNOR U2687 ( .A(n7809), .B(n7630), .Z(n7632) );
  XNOR U2688 ( .A(n8508), .B(n8612), .Z(n8512) );
  XNOR U2689 ( .A(n8860), .B(n8964), .Z(n8864) );
  XNOR U2690 ( .A(n9212), .B(n9316), .Z(n9216) );
  XNOR U2691 ( .A(n10268), .B(n10372), .Z(n10272) );
  XNOR U2692 ( .A(n10620), .B(n10726), .Z(n10624) );
  XNOR U2693 ( .A(n11190), .B(n11010), .Z(n11012) );
  XNOR U2694 ( .A(n11367), .B(n11187), .Z(n11189) );
  XNOR U2695 ( .A(n11543), .B(n11364), .Z(n11366) );
  XNOR U2696 ( .A(n11719), .B(n11540), .Z(n11542) );
  XNOR U2697 ( .A(n11895), .B(n11716), .Z(n11718) );
  XNOR U2698 ( .A(n12071), .B(n11892), .Z(n11894) );
  XNOR U2699 ( .A(n12247), .B(n12068), .Z(n12070) );
  XNOR U2700 ( .A(n12423), .B(n12244), .Z(n12246) );
  XNOR U2701 ( .A(n12599), .B(n12420), .Z(n12422) );
  XNOR U2702 ( .A(n12775), .B(n12596), .Z(n12598) );
  XNOR U2703 ( .A(n12951), .B(n12772), .Z(n12774) );
  XNOR U2704 ( .A(n13127), .B(n12948), .Z(n12950) );
  XNOR U2705 ( .A(n13116), .B(n13225), .Z(n13125) );
  XNOR U2706 ( .A(n13474), .B(n13578), .Z(n13482) );
  XNOR U2707 ( .A(n13826), .B(n13930), .Z(n13830) );
  XNOR U2708 ( .A(n15762), .B(n15866), .Z(n15766) );
  XNOR U2709 ( .A(n16113), .B(n16216), .Z(n16117) );
  XNOR U2710 ( .A(n16488), .B(n16592), .Z(n16492) );
  XNOR U2711 ( .A(n16665), .B(n16769), .Z(n16669) );
  XNOR U2712 ( .A(n16842), .B(n16946), .Z(n16846) );
  XNOR U2713 ( .A(n17018), .B(n17122), .Z(n17022) );
  XNOR U2714 ( .A(n3544), .B(n3646), .Z(n3548) );
  XNOR U2715 ( .A(n3904), .B(n4006), .Z(n3908) );
  XNOR U2716 ( .A(n4264), .B(n4366), .Z(n4268) );
  XNOR U2717 ( .A(n9569), .B(n9667), .Z(n9573) );
  XNOR U2718 ( .A(n1364), .B(n1485), .Z(n1368) );
  XNOR U2719 ( .A(n1565), .B(n1661), .Z(n1569) );
  XNOR U2720 ( .A(n1926), .B(n2022), .Z(n1930) );
  XNOR U2721 ( .A(n2287), .B(n2383), .Z(n2291) );
  XNOR U2722 ( .A(n2648), .B(n2744), .Z(n2652) );
  XNOR U2723 ( .A(n3009), .B(n3105), .Z(n3013) );
  XNOR U2724 ( .A(n3369), .B(n3465), .Z(n3373) );
  XNOR U2725 ( .A(n4629), .B(n4725), .Z(n4633) );
  XNOR U2726 ( .A(n8170), .B(n8258), .Z(n8165) );
  XNOR U2727 ( .A(n9926), .B(n10018), .Z(n9930) );
  XNOR U2728 ( .A(n14364), .B(n14456), .Z(n14368) );
  XNOR U2729 ( .A(n14716), .B(n14808), .Z(n14720) );
  XNOR U2730 ( .A(n15068), .B(n15160), .Z(n15072) );
  XNOR U2731 ( .A(n15420), .B(n15512), .Z(n15424) );
  XNOR U2732 ( .A(n19401), .B(n19493), .Z(n19405) );
  XNOR U2733 ( .A(n19185), .B(n19277), .Z(n19189) );
  XNOR U2734 ( .A(n18945), .B(n19037), .Z(n18949) );
  XNOR U2735 ( .A(n18681), .B(n18773), .Z(n18685) );
  XNOR U2736 ( .A(n18393), .B(n18485), .Z(n18397) );
  XNOR U2737 ( .A(n18081), .B(n18173), .Z(n18085) );
  XNOR U2738 ( .A(n17745), .B(n17837), .Z(n17749) );
  XNOR U2739 ( .A(n17380), .B(n17475), .Z(n17384) );
  XNOR U2740 ( .A(n988), .B(n1127), .Z(n992) );
  XNOR U2741 ( .A(n607), .B(n770), .Z(n611) );
  XNOR U2742 ( .A(n4994), .B(n5424), .Z(n4998) );
  XNOR U2743 ( .A(n5529), .B(n5614), .Z(n5533) );
  XNOR U2744 ( .A(n5705), .B(n5791), .Z(n5709) );
  XNOR U2745 ( .A(n6064), .B(n5885), .Z(n5887) );
  XNOR U2746 ( .A(n6240), .B(n6061), .Z(n6063) );
  XNOR U2747 ( .A(n6416), .B(n6237), .Z(n6239) );
  XNOR U2748 ( .A(n6592), .B(n6413), .Z(n6415) );
  XNOR U2749 ( .A(n6768), .B(n6589), .Z(n6591) );
  XNOR U2750 ( .A(n6944), .B(n6765), .Z(n6767) );
  XNOR U2751 ( .A(n7120), .B(n6941), .Z(n6943) );
  XNOR U2752 ( .A(n7296), .B(n7117), .Z(n7119) );
  XNOR U2753 ( .A(n7472), .B(n7293), .Z(n7295) );
  XNOR U2754 ( .A(n7648), .B(n7469), .Z(n7471) );
  XNOR U2755 ( .A(n7824), .B(n7645), .Z(n7647) );
  XNOR U2756 ( .A(n8000), .B(n7821), .Z(n7823) );
  XNOR U2757 ( .A(n8176), .B(n7997), .Z(n7999) );
  XNOR U2758 ( .A(n8352), .B(n8173), .Z(n8175) );
  XNOR U2759 ( .A(n8523), .B(n8609), .Z(n8531) );
  XNOR U2760 ( .A(n8875), .B(n8961), .Z(n8879) );
  XNOR U2761 ( .A(n9227), .B(n9313), .Z(n9231) );
  XNOR U2762 ( .A(n10283), .B(n10369), .Z(n10287) );
  XNOR U2763 ( .A(n10635), .B(n10723), .Z(n10639) );
  XNOR U2764 ( .A(n11205), .B(n11025), .Z(n11027) );
  XNOR U2765 ( .A(n11382), .B(n11202), .Z(n11204) );
  XNOR U2766 ( .A(n11558), .B(n11379), .Z(n11381) );
  XNOR U2767 ( .A(n11734), .B(n11555), .Z(n11557) );
  XNOR U2768 ( .A(n11910), .B(n11731), .Z(n11733) );
  XNOR U2769 ( .A(n12086), .B(n11907), .Z(n11909) );
  XNOR U2770 ( .A(n12262), .B(n12083), .Z(n12085) );
  XNOR U2771 ( .A(n12438), .B(n12259), .Z(n12261) );
  XNOR U2772 ( .A(n12614), .B(n12435), .Z(n12437) );
  XNOR U2773 ( .A(n12790), .B(n12611), .Z(n12613) );
  XNOR U2774 ( .A(n12966), .B(n12787), .Z(n12789) );
  XNOR U2775 ( .A(n13142), .B(n12963), .Z(n12965) );
  XNOR U2776 ( .A(n13318), .B(n13139), .Z(n13141) );
  XNOR U2777 ( .A(n13494), .B(n13315), .Z(n13317) );
  XNOR U2778 ( .A(n13670), .B(n13491), .Z(n13493) );
  XNOR U2779 ( .A(n13846), .B(n13667), .Z(n13669) );
  XNOR U2780 ( .A(n13845), .B(n13927), .Z(n13840) );
  XNOR U2781 ( .A(n14193), .B(n14279), .Z(n14197) );
  XNOR U2782 ( .A(n15777), .B(n15863), .Z(n15781) );
  XNOR U2783 ( .A(n16128), .B(n16213), .Z(n16132) );
  XNOR U2784 ( .A(n16503), .B(n16589), .Z(n16507) );
  XNOR U2785 ( .A(n16680), .B(n16766), .Z(n16684) );
  XNOR U2786 ( .A(n16857), .B(n16943), .Z(n16861) );
  XNOR U2787 ( .A(n17033), .B(n17119), .Z(n17037) );
  XNOR U2788 ( .A(n1018), .B(n1121), .Z(n1022) );
  XNOR U2789 ( .A(n3919), .B(n4003), .Z(n3923) );
  XNOR U2790 ( .A(n4279), .B(n4363), .Z(n4283) );
  XNOR U2791 ( .A(n9584), .B(n9664), .Z(n9588) );
  XNOR U2792 ( .A(n642), .B(n763), .Z(n646) );
  XNOR U2793 ( .A(n1189), .B(n1303), .Z(n1193) );
  XNOR U2794 ( .A(n1941), .B(n2019), .Z(n1945) );
  XNOR U2795 ( .A(n2302), .B(n2380), .Z(n2306) );
  XNOR U2796 ( .A(n2663), .B(n2741), .Z(n2667) );
  XNOR U2797 ( .A(n3024), .B(n3102), .Z(n3028) );
  XNOR U2798 ( .A(n3384), .B(n3462), .Z(n3388) );
  XNOR U2799 ( .A(n3744), .B(n3822), .Z(n3748) );
  XNOR U2800 ( .A(n4644), .B(n4722), .Z(n4648) );
  XNOR U2801 ( .A(n9941), .B(n10015), .Z(n9945) );
  XNOR U2802 ( .A(n14731), .B(n14805), .Z(n14735) );
  XNOR U2803 ( .A(n15083), .B(n15157), .Z(n15087) );
  XNOR U2804 ( .A(n15435), .B(n15509), .Z(n15439) );
  XNOR U2805 ( .A(n19776), .B(n19850), .Z(n19780) );
  XNOR U2806 ( .A(n19608), .B(n19682), .Z(n19612) );
  XNOR U2807 ( .A(n19416), .B(n19490), .Z(n19420) );
  XNOR U2808 ( .A(n19200), .B(n19274), .Z(n19204) );
  XNOR U2809 ( .A(n18960), .B(n19034), .Z(n18964) );
  XNOR U2810 ( .A(n18696), .B(n18770), .Z(n18700) );
  XNOR U2811 ( .A(n18408), .B(n18482), .Z(n18412) );
  XNOR U2812 ( .A(n18096), .B(n18170), .Z(n18100) );
  XNOR U2813 ( .A(n17760), .B(n17834), .Z(n17764) );
  XNOR U2814 ( .A(n17395), .B(n17472), .Z(n17399) );
  XNOR U2815 ( .A(n813), .B(n945), .Z(n817) );
  XNOR U2816 ( .A(n432), .B(n588), .Z(n436) );
  XNOR U2817 ( .A(n1043), .B(n1116), .Z(n1047) );
  XNOR U2818 ( .A(n1404), .B(n1477), .Z(n1408) );
  XNOR U2819 ( .A(n1765), .B(n1838), .Z(n1769) );
  XNOR U2820 ( .A(n5009), .B(n5418), .Z(n5013) );
  XNOR U2821 ( .A(n5544), .B(n5611), .Z(n5548) );
  XNOR U2822 ( .A(n5720), .B(n5788), .Z(n5724) );
  XNOR U2823 ( .A(n6079), .B(n5900), .Z(n5902) );
  XNOR U2824 ( .A(n6255), .B(n6076), .Z(n6078) );
  XNOR U2825 ( .A(n6431), .B(n6252), .Z(n6254) );
  XNOR U2826 ( .A(n6607), .B(n6428), .Z(n6430) );
  XNOR U2827 ( .A(n6783), .B(n6604), .Z(n6606) );
  XNOR U2828 ( .A(n6959), .B(n6780), .Z(n6782) );
  XNOR U2829 ( .A(n7135), .B(n6956), .Z(n6958) );
  XNOR U2830 ( .A(n7311), .B(n7132), .Z(n7134) );
  XNOR U2831 ( .A(n7487), .B(n7308), .Z(n7310) );
  XNOR U2832 ( .A(n7663), .B(n7484), .Z(n7486) );
  XNOR U2833 ( .A(n7839), .B(n7660), .Z(n7662) );
  XNOR U2834 ( .A(n8015), .B(n7836), .Z(n7838) );
  XNOR U2835 ( .A(n8191), .B(n8012), .Z(n8014) );
  XNOR U2836 ( .A(n8367), .B(n8188), .Z(n8190) );
  XNOR U2837 ( .A(n8543), .B(n8364), .Z(n8366) );
  XNOR U2838 ( .A(n8719), .B(n8540), .Z(n8542) );
  XNOR U2839 ( .A(n8895), .B(n8716), .Z(n8718) );
  XNOR U2840 ( .A(n8894), .B(n8958), .Z(n8889) );
  XNOR U2841 ( .A(n9242), .B(n9310), .Z(n9246) );
  XNOR U2842 ( .A(n10298), .B(n10366), .Z(n10302) );
  XNOR U2843 ( .A(n10650), .B(n10720), .Z(n10654) );
  XNOR U2844 ( .A(n11037), .B(n11105), .Z(n11041) );
  XNOR U2845 ( .A(n11214), .B(n11282), .Z(n11218) );
  XNOR U2846 ( .A(n11573), .B(n11394), .Z(n11396) );
  XNOR U2847 ( .A(n11749), .B(n11570), .Z(n11572) );
  XNOR U2848 ( .A(n11925), .B(n11746), .Z(n11748) );
  XNOR U2849 ( .A(n12101), .B(n11922), .Z(n11924) );
  XNOR U2850 ( .A(n12277), .B(n12098), .Z(n12100) );
  XNOR U2851 ( .A(n12453), .B(n12274), .Z(n12276) );
  XNOR U2852 ( .A(n12629), .B(n12450), .Z(n12452) );
  XNOR U2853 ( .A(n12805), .B(n12626), .Z(n12628) );
  XNOR U2854 ( .A(n12981), .B(n12802), .Z(n12804) );
  XNOR U2855 ( .A(n13157), .B(n12978), .Z(n12980) );
  XNOR U2856 ( .A(n13333), .B(n13154), .Z(n13156) );
  XNOR U2857 ( .A(n13509), .B(n13330), .Z(n13332) );
  XNOR U2858 ( .A(n13685), .B(n13506), .Z(n13508) );
  XNOR U2859 ( .A(n13861), .B(n13682), .Z(n13684) );
  XNOR U2860 ( .A(n14037), .B(n13858), .Z(n13860) );
  XNOR U2861 ( .A(n14213), .B(n14034), .Z(n14036) );
  XNOR U2862 ( .A(n14202), .B(n14275), .Z(n14211) );
  XNOR U2863 ( .A(n14560), .B(n14628), .Z(n14568) );
  XNOR U2864 ( .A(n15792), .B(n15860), .Z(n15796) );
  XNOR U2865 ( .A(n16143), .B(n16210), .Z(n16147) );
  XNOR U2866 ( .A(n16518), .B(n16586), .Z(n16522) );
  XNOR U2867 ( .A(n16695), .B(n16763), .Z(n16699) );
  XNOR U2868 ( .A(n16872), .B(n16940), .Z(n16876) );
  XNOR U2869 ( .A(n17048), .B(n17116), .Z(n17052) );
  XNOR U2870 ( .A(n843), .B(n939), .Z(n847) );
  XNOR U2871 ( .A(n482), .B(n578), .Z(n486) );
  XNOR U2872 ( .A(n4294), .B(n4360), .Z(n4298) );
  XNOR U2873 ( .A(n9599), .B(n9661), .Z(n9603) );
  XNOR U2874 ( .A(n467), .B(n581), .Z(n471) );
  XNOR U2875 ( .A(n2317), .B(n2377), .Z(n2321) );
  XNOR U2876 ( .A(n2678), .B(n2738), .Z(n2682) );
  XNOR U2877 ( .A(n3039), .B(n3099), .Z(n3043) );
  XNOR U2878 ( .A(n3399), .B(n3459), .Z(n3403) );
  XNOR U2879 ( .A(n3759), .B(n3819), .Z(n3763) );
  XNOR U2880 ( .A(n4119), .B(n4179), .Z(n4123) );
  XNOR U2881 ( .A(n4659), .B(n4719), .Z(n4663) );
  XNOR U2882 ( .A(n9956), .B(n10012), .Z(n9960) );
  XNOR U2883 ( .A(n15098), .B(n15154), .Z(n15102) );
  XNOR U2884 ( .A(n15450), .B(n15506), .Z(n15454) );
  XNOR U2885 ( .A(n19935), .B(n19991), .Z(n19939) );
  XNOR U2886 ( .A(n19791), .B(n19847), .Z(n19795) );
  XNOR U2887 ( .A(n19623), .B(n19679), .Z(n19627) );
  XNOR U2888 ( .A(n19431), .B(n19487), .Z(n19435) );
  XNOR U2889 ( .A(n19215), .B(n19271), .Z(n19219) );
  XNOR U2890 ( .A(n18975), .B(n19031), .Z(n18979) );
  XNOR U2891 ( .A(n18711), .B(n18767), .Z(n18715) );
  XNOR U2892 ( .A(n18423), .B(n18479), .Z(n18427) );
  XNOR U2893 ( .A(n18111), .B(n18167), .Z(n18115) );
  XNOR U2894 ( .A(n17775), .B(n17831), .Z(n17779) );
  XNOR U2895 ( .A(n17410), .B(n17469), .Z(n17414) );
  XNOR U2896 ( .A(n447), .B(n585), .Z(n451) );
  XNOR U2897 ( .A(n697), .B(n752), .Z(n701) );
  XNOR U2898 ( .A(n1058), .B(n1113), .Z(n1062) );
  XNOR U2899 ( .A(n1419), .B(n1474), .Z(n1423) );
  XNOR U2900 ( .A(n1780), .B(n1835), .Z(n1784) );
  XNOR U2901 ( .A(n2141), .B(n2196), .Z(n2145) );
  XNOR U2902 ( .A(n5024), .B(n5412), .Z(n5028) );
  XNOR U2903 ( .A(n5559), .B(n5608), .Z(n5563) );
  XNOR U2904 ( .A(n5735), .B(n5785), .Z(n5739) );
  XNOR U2905 ( .A(n6094), .B(n5915), .Z(n5917) );
  XNOR U2906 ( .A(n6270), .B(n6091), .Z(n6093) );
  XNOR U2907 ( .A(n6446), .B(n6267), .Z(n6269) );
  XNOR U2908 ( .A(n6622), .B(n6443), .Z(n6445) );
  XNOR U2909 ( .A(n6798), .B(n6619), .Z(n6621) );
  XNOR U2910 ( .A(n6974), .B(n6795), .Z(n6797) );
  XNOR U2911 ( .A(n7150), .B(n6971), .Z(n6973) );
  XNOR U2912 ( .A(n7326), .B(n7147), .Z(n7149) );
  XNOR U2913 ( .A(n7502), .B(n7323), .Z(n7325) );
  XNOR U2914 ( .A(n7678), .B(n7499), .Z(n7501) );
  XNOR U2915 ( .A(n7854), .B(n7675), .Z(n7677) );
  XNOR U2916 ( .A(n8030), .B(n7851), .Z(n7853) );
  XNOR U2917 ( .A(n8206), .B(n8027), .Z(n8029) );
  XNOR U2918 ( .A(n8382), .B(n8203), .Z(n8205) );
  XNOR U2919 ( .A(n8558), .B(n8379), .Z(n8381) );
  XNOR U2920 ( .A(n8734), .B(n8555), .Z(n8557) );
  XNOR U2921 ( .A(n8910), .B(n8731), .Z(n8733) );
  XNOR U2922 ( .A(n9086), .B(n8907), .Z(n8909) );
  XNOR U2923 ( .A(n9262), .B(n9083), .Z(n9085) );
  XNOR U2924 ( .A(n9438), .B(n9259), .Z(n9261) );
  XNOR U2925 ( .A(n9437), .B(n9483), .Z(n9432) );
  XNOR U2926 ( .A(n10313), .B(n10363), .Z(n10317) );
  XNOR U2927 ( .A(n10665), .B(n10717), .Z(n10669) );
  XNOR U2928 ( .A(n11235), .B(n11055), .Z(n11057) );
  XNOR U2929 ( .A(n11412), .B(n11232), .Z(n11234) );
  XNOR U2930 ( .A(n11588), .B(n11409), .Z(n11411) );
  XNOR U2931 ( .A(n11764), .B(n11585), .Z(n11587) );
  XNOR U2932 ( .A(n11940), .B(n11761), .Z(n11763) );
  XNOR U2933 ( .A(n12116), .B(n11937), .Z(n11939) );
  XNOR U2934 ( .A(n12292), .B(n12113), .Z(n12115) );
  XNOR U2935 ( .A(n12468), .B(n12289), .Z(n12291) );
  XNOR U2936 ( .A(n12644), .B(n12465), .Z(n12467) );
  XNOR U2937 ( .A(n12820), .B(n12641), .Z(n12643) );
  XNOR U2938 ( .A(n12996), .B(n12817), .Z(n12819) );
  XNOR U2939 ( .A(n13172), .B(n12993), .Z(n12995) );
  XNOR U2940 ( .A(n13348), .B(n13169), .Z(n13171) );
  XNOR U2941 ( .A(n13524), .B(n13345), .Z(n13347) );
  XNOR U2942 ( .A(n13700), .B(n13521), .Z(n13523) );
  XNOR U2943 ( .A(n13876), .B(n13697), .Z(n13699) );
  XNOR U2944 ( .A(n14052), .B(n13873), .Z(n13875) );
  XNOR U2945 ( .A(n14228), .B(n14049), .Z(n14051) );
  XNOR U2946 ( .A(n14404), .B(n14225), .Z(n14227) );
  XNOR U2947 ( .A(n14580), .B(n14401), .Z(n14403) );
  XNOR U2948 ( .A(n14756), .B(n14577), .Z(n14579) );
  XNOR U2949 ( .A(n14932), .B(n14753), .Z(n14755) );
  XNOR U2950 ( .A(n14931), .B(n14977), .Z(n14926) );
  XNOR U2951 ( .A(n15807), .B(n15857), .Z(n15811) );
  XNOR U2952 ( .A(n16158), .B(n16207), .Z(n16162) );
  XNOR U2953 ( .A(n16533), .B(n16583), .Z(n16537) );
  XNOR U2954 ( .A(n16710), .B(n16760), .Z(n16714) );
  XNOR U2955 ( .A(n16887), .B(n16937), .Z(n16891) );
  XNOR U2956 ( .A(n17063), .B(n17113), .Z(n17067) );
  XNOR U2957 ( .A(n497), .B(n575), .Z(n501) );
  XNOR U2958 ( .A(n9790), .B(n9834), .Z(n9798) );
  XNOR U2959 ( .A(n2693), .B(n2735), .Z(n2697) );
  XNOR U2960 ( .A(n3054), .B(n3096), .Z(n3058) );
  XNOR U2961 ( .A(n3414), .B(n3456), .Z(n3418) );
  XNOR U2962 ( .A(n3774), .B(n3816), .Z(n3778) );
  XNOR U2963 ( .A(n4134), .B(n4176), .Z(n4138) );
  XNOR U2964 ( .A(n4674), .B(n4716), .Z(n4678) );
  XNOR U2965 ( .A(n15465), .B(n15503), .Z(n15473) );
  XNOR U2966 ( .A(n20166), .B(n20204), .Z(n20170) );
  XNOR U2967 ( .A(n20070), .B(n20108), .Z(n20074) );
  XNOR U2968 ( .A(n19950), .B(n19988), .Z(n19954) );
  XNOR U2969 ( .A(n19806), .B(n19844), .Z(n19810) );
  XNOR U2970 ( .A(n19638), .B(n19676), .Z(n19642) );
  XNOR U2971 ( .A(n19446), .B(n19484), .Z(n19450) );
  XNOR U2972 ( .A(n19230), .B(n19268), .Z(n19234) );
  XNOR U2973 ( .A(n18990), .B(n19028), .Z(n18994) );
  XNOR U2974 ( .A(n18726), .B(n18764), .Z(n18730) );
  XNOR U2975 ( .A(n18438), .B(n18476), .Z(n18442) );
  XNOR U2976 ( .A(n18126), .B(n18164), .Z(n18130) );
  XNOR U2977 ( .A(n17790), .B(n17828), .Z(n17794) );
  XNOR U2978 ( .A(n17425), .B(n17466), .Z(n17429) );
  XNOR U2979 ( .A(n712), .B(n749), .Z(n716) );
  XNOR U2980 ( .A(n1073), .B(n1110), .Z(n1077) );
  XNOR U2981 ( .A(n1434), .B(n1471), .Z(n1438) );
  XNOR U2982 ( .A(n1795), .B(n1832), .Z(n1799) );
  XNOR U2983 ( .A(n2156), .B(n2193), .Z(n2160) );
  XNOR U2984 ( .A(n2517), .B(n2554), .Z(n2521) );
  XNOR U2985 ( .A(n4499), .B(n4535), .Z(n4503) );
  XNOR U2986 ( .A(n5039), .B(n5406), .Z(n5043) );
  XNOR U2987 ( .A(n5574), .B(n5605), .Z(n5578) );
  XNOR U2988 ( .A(n5750), .B(n5782), .Z(n5754) );
  XNOR U2989 ( .A(n6109), .B(n5930), .Z(n5932) );
  XNOR U2990 ( .A(n6285), .B(n6106), .Z(n6108) );
  XNOR U2991 ( .A(n6461), .B(n6282), .Z(n6284) );
  XNOR U2992 ( .A(n6637), .B(n6458), .Z(n6460) );
  XNOR U2993 ( .A(n6813), .B(n6634), .Z(n6636) );
  XNOR U2994 ( .A(n6989), .B(n6810), .Z(n6812) );
  XNOR U2995 ( .A(n7165), .B(n6986), .Z(n6988) );
  XNOR U2996 ( .A(n7341), .B(n7162), .Z(n7164) );
  XNOR U2997 ( .A(n7517), .B(n7338), .Z(n7340) );
  XNOR U2998 ( .A(n7693), .B(n7514), .Z(n7516) );
  XNOR U2999 ( .A(n7869), .B(n7690), .Z(n7692) );
  XNOR U3000 ( .A(n8045), .B(n7866), .Z(n7868) );
  XNOR U3001 ( .A(n8221), .B(n8042), .Z(n8044) );
  XNOR U3002 ( .A(n8397), .B(n8218), .Z(n8220) );
  XNOR U3003 ( .A(n8573), .B(n8394), .Z(n8396) );
  XNOR U3004 ( .A(n8749), .B(n8570), .Z(n8572) );
  XNOR U3005 ( .A(n8925), .B(n8746), .Z(n8748) );
  XNOR U3006 ( .A(n9101), .B(n8922), .Z(n8924) );
  XNOR U3007 ( .A(n9277), .B(n9098), .Z(n9100) );
  XNOR U3008 ( .A(n9453), .B(n9274), .Z(n9276) );
  XNOR U3009 ( .A(n9629), .B(n9450), .Z(n9452) );
  XNOR U3010 ( .A(n9805), .B(n9626), .Z(n9628) );
  XNOR U3011 ( .A(n9981), .B(n9802), .Z(n9804) );
  XNOR U3012 ( .A(n10328), .B(n10360), .Z(n10332) );
  XNOR U3013 ( .A(n10680), .B(n10714), .Z(n10684) );
  XNOR U3014 ( .A(n11067), .B(n11099), .Z(n11071) );
  XNOR U3015 ( .A(n11244), .B(n11276), .Z(n11248) );
  XNOR U3016 ( .A(n11421), .B(n11453), .Z(n11425) );
  XNOR U3017 ( .A(n11779), .B(n11600), .Z(n11602) );
  XNOR U3018 ( .A(n11955), .B(n11776), .Z(n11778) );
  XNOR U3019 ( .A(n12131), .B(n11952), .Z(n11954) );
  XNOR U3020 ( .A(n12307), .B(n12128), .Z(n12130) );
  XNOR U3021 ( .A(n12483), .B(n12304), .Z(n12306) );
  XNOR U3022 ( .A(n12659), .B(n12480), .Z(n12482) );
  XNOR U3023 ( .A(n12835), .B(n12656), .Z(n12658) );
  XNOR U3024 ( .A(n13011), .B(n12832), .Z(n12834) );
  XNOR U3025 ( .A(n13187), .B(n13008), .Z(n13010) );
  XNOR U3026 ( .A(n13363), .B(n13184), .Z(n13186) );
  XNOR U3027 ( .A(n13539), .B(n13360), .Z(n13362) );
  XNOR U3028 ( .A(n13715), .B(n13536), .Z(n13538) );
  XNOR U3029 ( .A(n13891), .B(n13712), .Z(n13714) );
  XNOR U3030 ( .A(n14067), .B(n13888), .Z(n13890) );
  XNOR U3031 ( .A(n14243), .B(n14064), .Z(n14066) );
  XNOR U3032 ( .A(n14419), .B(n14240), .Z(n14242) );
  XNOR U3033 ( .A(n14595), .B(n14416), .Z(n14418) );
  XNOR U3034 ( .A(n14771), .B(n14592), .Z(n14594) );
  XNOR U3035 ( .A(n14947), .B(n14768), .Z(n14770) );
  XNOR U3036 ( .A(n15123), .B(n14944), .Z(n14946) );
  XNOR U3037 ( .A(n15299), .B(n15120), .Z(n15122) );
  XNOR U3038 ( .A(n15288), .B(n15325), .Z(n15297) );
  XNOR U3039 ( .A(n15822), .B(n15854), .Z(n15826) );
  XNOR U3040 ( .A(n16173), .B(n16204), .Z(n16177) );
  XNOR U3041 ( .A(n16548), .B(n16580), .Z(n16552) );
  XNOR U3042 ( .A(n16725), .B(n16757), .Z(n16729) );
  XNOR U3043 ( .A(n16902), .B(n16934), .Z(n16906) );
  XNOR U3044 ( .A(n17078), .B(n17110), .Z(n17082) );
  XNOR U3045 ( .A(n10161), .B(n10183), .Z(n10156) );
  XNOR U3046 ( .A(n3069), .B(n3093), .Z(n3073) );
  XNOR U3047 ( .A(n3609), .B(n3633), .Z(n3613) );
  XNOR U3048 ( .A(n4149), .B(n4173), .Z(n4153) );
  XNOR U3049 ( .A(n20280), .B(n20311), .Z(n20289) );
  XNOR U3050 ( .A(n20220), .B(n20240), .Z(n20229) );
  XNOR U3051 ( .A(n20136), .B(n20156), .Z(n20145) );
  XNOR U3052 ( .A(n20028), .B(n20048), .Z(n20037) );
  XNOR U3053 ( .A(n19896), .B(n19916), .Z(n19905) );
  XNOR U3054 ( .A(n19740), .B(n19760), .Z(n19749) );
  XNOR U3055 ( .A(n19560), .B(n19580), .Z(n19569) );
  XNOR U3056 ( .A(n19356), .B(n19376), .Z(n19365) );
  XNOR U3057 ( .A(n19128), .B(n19148), .Z(n19137) );
  XNOR U3058 ( .A(n18876), .B(n18896), .Z(n18885) );
  XNOR U3059 ( .A(n18600), .B(n18620), .Z(n18609) );
  XNOR U3060 ( .A(n18300), .B(n18320), .Z(n18309) );
  XNOR U3061 ( .A(n17976), .B(n17996), .Z(n17985) );
  XNOR U3062 ( .A(n17625), .B(n17645), .Z(n17634) );
  XNOR U3063 ( .A(n727), .B(n746), .Z(n736) );
  XNOR U3064 ( .A(n1088), .B(n1107), .Z(n1097) );
  XNOR U3065 ( .A(n1449), .B(n1468), .Z(n1458) );
  XNOR U3066 ( .A(n1810), .B(n1829), .Z(n1819) );
  XNOR U3067 ( .A(n2171), .B(n2190), .Z(n2180) );
  XNOR U3068 ( .A(n2532), .B(n2551), .Z(n2541) );
  XNOR U3069 ( .A(n2893), .B(n2912), .Z(n2902) );
  XNOR U3070 ( .A(n3434), .B(n3452), .Z(n3443) );
  XNOR U3071 ( .A(n3974), .B(n3992), .Z(n3983) );
  XNOR U3072 ( .A(n4514), .B(n4532), .Z(n4523) );
  XNOR U3073 ( .A(n4874), .B(n4892), .Z(n4883) );
  XNOR U3074 ( .A(n5765), .B(n5779), .Z(n5769) );
  XNOR U3075 ( .A(n6124), .B(n5945), .Z(n5947) );
  XNOR U3076 ( .A(n6118), .B(n6132), .Z(n6122) );
  XNOR U3077 ( .A(n6294), .B(n6308), .Z(n6298) );
  XNOR U3078 ( .A(n6652), .B(n6473), .Z(n6475) );
  XNOR U3079 ( .A(n6646), .B(n6660), .Z(n6650) );
  XNOR U3080 ( .A(n6822), .B(n6836), .Z(n6826) );
  XNOR U3081 ( .A(n7180), .B(n7001), .Z(n7003) );
  XNOR U3082 ( .A(n7174), .B(n7188), .Z(n7178) );
  XNOR U3083 ( .A(n7350), .B(n7364), .Z(n7354) );
  XNOR U3084 ( .A(n7708), .B(n7529), .Z(n7531) );
  XNOR U3085 ( .A(n7702), .B(n7716), .Z(n7706) );
  XNOR U3086 ( .A(n7878), .B(n7892), .Z(n7882) );
  XNOR U3087 ( .A(n8236), .B(n8057), .Z(n8059) );
  XNOR U3088 ( .A(n8230), .B(n8244), .Z(n8234) );
  XNOR U3089 ( .A(n8406), .B(n8420), .Z(n8410) );
  XNOR U3090 ( .A(n8764), .B(n8585), .Z(n8587) );
  XNOR U3091 ( .A(n8758), .B(n8772), .Z(n8762) );
  XNOR U3092 ( .A(n8934), .B(n8948), .Z(n8938) );
  XNOR U3093 ( .A(n9292), .B(n9113), .Z(n9115) );
  XNOR U3094 ( .A(n9286), .B(n9300), .Z(n9290) );
  XNOR U3095 ( .A(n9462), .B(n9476), .Z(n9466) );
  XNOR U3096 ( .A(n9820), .B(n9641), .Z(n9643) );
  XNOR U3097 ( .A(n9814), .B(n9828), .Z(n9818) );
  XNOR U3098 ( .A(n9990), .B(n10004), .Z(n9994) );
  XNOR U3099 ( .A(n10348), .B(n10169), .Z(n10171) );
  XNOR U3100 ( .A(n10873), .B(n10886), .Z(n10879) );
  XNOR U3101 ( .A(n11086), .B(n11085), .Z(n10889) );
  XNOR U3102 ( .A(n11259), .B(n11264), .Z(n11094) );
  XNOR U3103 ( .A(n11440), .B(n11439), .Z(n11269) );
  XNOR U3104 ( .A(n11612), .B(n11617), .Z(n11448) );
  XNOR U3105 ( .A(n11792), .B(n11791), .Z(n11622) );
  XNOR U3106 ( .A(n11964), .B(n11969), .Z(n11800) );
  XNOR U3107 ( .A(n12144), .B(n12143), .Z(n11974) );
  XNOR U3108 ( .A(n12316), .B(n12321), .Z(n12152) );
  XNOR U3109 ( .A(n12496), .B(n12495), .Z(n12326) );
  XNOR U3110 ( .A(n12668), .B(n12673), .Z(n12504) );
  XNOR U3111 ( .A(n12848), .B(n12847), .Z(n12678) );
  XNOR U3112 ( .A(n13020), .B(n13025), .Z(n12856) );
  XNOR U3113 ( .A(n13200), .B(n13199), .Z(n13030) );
  XNOR U3114 ( .A(n13372), .B(n13377), .Z(n13208) );
  XNOR U3115 ( .A(n13552), .B(n13551), .Z(n13382) );
  XNOR U3116 ( .A(n13724), .B(n13729), .Z(n13560) );
  XNOR U3117 ( .A(n13904), .B(n13903), .Z(n13734) );
  XNOR U3118 ( .A(n14076), .B(n14081), .Z(n13912) );
  XNOR U3119 ( .A(n14256), .B(n14255), .Z(n14086) );
  XNOR U3120 ( .A(n14428), .B(n14433), .Z(n14264) );
  XNOR U3121 ( .A(n14608), .B(n14607), .Z(n14438) );
  XNOR U3122 ( .A(n14780), .B(n14785), .Z(n14616) );
  XNOR U3123 ( .A(n14960), .B(n14959), .Z(n14790) );
  XNOR U3124 ( .A(n15132), .B(n15137), .Z(n14968) );
  XNOR U3125 ( .A(n15312), .B(n15311), .Z(n15142) );
  XNOR U3126 ( .A(n15484), .B(n15489), .Z(n15320) );
  XNOR U3127 ( .A(n15664), .B(n15663), .Z(n15494) );
  XNOR U3128 ( .A(n15831), .B(n15841), .Z(n15672) );
  XNOR U3129 ( .A(n16361), .B(n16360), .Z(n16193) );
  XNOR U3130 ( .A(n16563), .B(n16568), .Z(n16369) );
  XNOR U3131 ( .A(n16744), .B(n16743), .Z(n16573) );
  XNOR U3132 ( .A(n16917), .B(n16922), .Z(n16752) );
  XNOR U3133 ( .A(n17097), .B(n17096), .Z(n16927) );
  XNOR U3134 ( .A(n17269), .B(n17274), .Z(n17105) );
  XOR U3135 ( .A(n5594), .B(n5601), .Z(n5598) );
  XOR U3136 ( .A(n10517), .B(n10530), .Z(n10528) );
  AND U3137 ( .A(n1099), .B(n1100), .Z(n918) );
  AND U3138 ( .A(n1821), .B(n1822), .Z(n1640) );
  AND U3139 ( .A(n2543), .B(n2544), .Z(n2362) );
  XNOR U3140 ( .A(n3084), .B(n3086), .Z(n3085) );
  XNOR U3141 ( .A(n3624), .B(n3626), .Z(n3625) );
  XNOR U3142 ( .A(n4164), .B(n4166), .Z(n4165) );
  NOR U3143 ( .A(n2), .B(n1), .Z(n4884) );
  AND U3144 ( .A(n7), .B(n8), .Z(n5) );
  XNOR U3145 ( .A(n2045), .B(n2215), .Z(n2050) );
  XNOR U3146 ( .A(n2406), .B(n2576), .Z(n2411) );
  XNOR U3147 ( .A(n2767), .B(n2937), .Z(n2772) );
  XNOR U3148 ( .A(n3128), .B(n3297), .Z(n3133) );
  XNOR U3149 ( .A(n3488), .B(n3657), .Z(n3493) );
  XNOR U3150 ( .A(n3848), .B(n4017), .Z(n3853) );
  XNOR U3151 ( .A(n4208), .B(n4377), .Z(n4213) );
  XNOR U3152 ( .A(n6169), .B(n6334), .Z(n6178) );
  XNOR U3153 ( .A(n6521), .B(n6686), .Z(n6526) );
  XNOR U3154 ( .A(n8281), .B(n8446), .Z(n8286) );
  XNOR U3155 ( .A(n8633), .B(n8798), .Z(n8638) );
  XNOR U3156 ( .A(n8985), .B(n9150), .Z(n8990) );
  XNOR U3157 ( .A(n13071), .B(n13236), .Z(n13076) );
  XNOR U3158 ( .A(n17856), .B(n18020), .Z(n17860) );
  XNOR U3159 ( .A(n17505), .B(n17669), .Z(n17509) );
  XNOR U3160 ( .A(n4574), .B(n4736), .Z(n4578) );
  XNOR U3161 ( .A(n6879), .B(n7037), .Z(n6883) );
  XNOR U3162 ( .A(n7231), .B(n7389), .Z(n7235) );
  XNOR U3163 ( .A(n9343), .B(n9501), .Z(n9347) );
  XNOR U3164 ( .A(n9695), .B(n9853), .Z(n9699) );
  XNOR U3165 ( .A(n10047), .B(n10205), .Z(n10051) );
  XNOR U3166 ( .A(n10399), .B(n10557), .Z(n10403) );
  XNOR U3167 ( .A(n10753), .B(n10941), .Z(n10757) );
  XNOR U3168 ( .A(n10962), .B(n11120), .Z(n10966) );
  XNOR U3169 ( .A(n11139), .B(n11297), .Z(n11143) );
  XNOR U3170 ( .A(n11315), .B(n11474), .Z(n11320) );
  XNOR U3171 ( .A(n11487), .B(n11650), .Z(n11496) );
  XNOR U3172 ( .A(n11845), .B(n12003), .Z(n11853) );
  XNOR U3173 ( .A(n12197), .B(n12355), .Z(n12201) );
  XNOR U3174 ( .A(n12549), .B(n12707), .Z(n12553) );
  XNOR U3175 ( .A(n12901), .B(n13059), .Z(n12905) );
  XNOR U3176 ( .A(n13781), .B(n13939), .Z(n13785) );
  XNOR U3177 ( .A(n14133), .B(n14291), .Z(n14137) );
  XNOR U3178 ( .A(n14485), .B(n14643), .Z(n14489) );
  XNOR U3179 ( .A(n14837), .B(n14995), .Z(n14841) );
  XNOR U3180 ( .A(n15189), .B(n15347), .Z(n15193) );
  XNOR U3181 ( .A(n15541), .B(n15699), .Z(n15545) );
  XNOR U3182 ( .A(n15893), .B(n16050), .Z(n15897) );
  XNOR U3183 ( .A(n16243), .B(n16422), .Z(n16247) );
  XNOR U3184 ( .A(n16626), .B(n16446), .Z(n16448) );
  XNOR U3185 ( .A(n16803), .B(n16623), .Z(n16625) );
  XNOR U3186 ( .A(n16979), .B(n16800), .Z(n16802) );
  XNOR U3187 ( .A(n17155), .B(n16976), .Z(n16978) );
  XNOR U3188 ( .A(n17154), .B(n17303), .Z(n17149) );
  XNOR U3189 ( .A(n1695), .B(n1852), .Z(n1699) );
  XNOR U3190 ( .A(n4939), .B(n5446), .Z(n4943) );
  XNOR U3191 ( .A(n5474), .B(n5625), .Z(n5478) );
  XNOR U3192 ( .A(n5650), .B(n5802), .Z(n5654) );
  XNOR U3193 ( .A(n6009), .B(n5830), .Z(n5832) );
  XNOR U3194 ( .A(n6185), .B(n6006), .Z(n6008) );
  XNOR U3195 ( .A(n6361), .B(n6182), .Z(n6184) );
  XNOR U3196 ( .A(n7588), .B(n7740), .Z(n7592) );
  XNOR U3197 ( .A(n7940), .B(n8092), .Z(n7944) );
  XNOR U3198 ( .A(n13610), .B(n13762), .Z(n13614) );
  XNOR U3199 ( .A(n2061), .B(n2212), .Z(n2065) );
  XNOR U3200 ( .A(n2422), .B(n2573), .Z(n2426) );
  XNOR U3201 ( .A(n2783), .B(n2934), .Z(n2787) );
  XNOR U3202 ( .A(n3144), .B(n3294), .Z(n3148) );
  XNOR U3203 ( .A(n3504), .B(n3654), .Z(n3508) );
  XNOR U3204 ( .A(n3864), .B(n4014), .Z(n3868) );
  XNOR U3205 ( .A(n4224), .B(n4374), .Z(n4228) );
  XNOR U3206 ( .A(n6541), .B(n6683), .Z(n6536) );
  XNOR U3207 ( .A(n8297), .B(n8443), .Z(n8301) );
  XNOR U3208 ( .A(n8649), .B(n8795), .Z(n8653) );
  XNOR U3209 ( .A(n9001), .B(n9147), .Z(n9005) );
  XNOR U3210 ( .A(n13439), .B(n13585), .Z(n13443) );
  XNOR U3211 ( .A(n18195), .B(n18341), .Z(n18199) );
  XNOR U3212 ( .A(n17871), .B(n18017), .Z(n17875) );
  XNOR U3213 ( .A(n17520), .B(n17666), .Z(n17524) );
  XNOR U3214 ( .A(n4589), .B(n4733), .Z(n4593) );
  XNOR U3215 ( .A(n6894), .B(n7034), .Z(n6902) );
  XNOR U3216 ( .A(n7246), .B(n7386), .Z(n7250) );
  XNOR U3217 ( .A(n9358), .B(n9498), .Z(n9362) );
  XNOR U3218 ( .A(n9710), .B(n9850), .Z(n9714) );
  XNOR U3219 ( .A(n10062), .B(n10202), .Z(n10066) );
  XNOR U3220 ( .A(n10414), .B(n10554), .Z(n10418) );
  XNOR U3221 ( .A(n10768), .B(n10935), .Z(n10772) );
  XNOR U3222 ( .A(n11160), .B(n10980), .Z(n10982) );
  XNOR U3223 ( .A(n11337), .B(n11157), .Z(n11159) );
  XNOR U3224 ( .A(n11331), .B(n11471), .Z(n11335) );
  XNOR U3225 ( .A(n11507), .B(n11647), .Z(n11511) );
  XNOR U3226 ( .A(n11683), .B(n11823), .Z(n11687) );
  XNOR U3227 ( .A(n11859), .B(n11999), .Z(n11863) );
  XNOR U3228 ( .A(n12217), .B(n12038), .Z(n12040) );
  XNOR U3229 ( .A(n12216), .B(n12352), .Z(n12211) );
  XNOR U3230 ( .A(n12564), .B(n12704), .Z(n12568) );
  XNOR U3231 ( .A(n12916), .B(n13056), .Z(n12920) );
  XNOR U3232 ( .A(n13268), .B(n13408), .Z(n13272) );
  XNOR U3233 ( .A(n14148), .B(n14288), .Z(n14152) );
  XNOR U3234 ( .A(n14500), .B(n14640), .Z(n14504) );
  XNOR U3235 ( .A(n14852), .B(n14992), .Z(n14856) );
  XNOR U3236 ( .A(n15204), .B(n15344), .Z(n15208) );
  XNOR U3237 ( .A(n15556), .B(n15696), .Z(n15560) );
  XNOR U3238 ( .A(n15908), .B(n16047), .Z(n15912) );
  XNOR U3239 ( .A(n16258), .B(n16416), .Z(n16262) );
  XNOR U3240 ( .A(n16641), .B(n16461), .Z(n16463) );
  XNOR U3241 ( .A(n16818), .B(n16638), .Z(n16640) );
  XNOR U3242 ( .A(n16994), .B(n16815), .Z(n16817) );
  XNOR U3243 ( .A(n17170), .B(n16991), .Z(n16993) );
  XNOR U3244 ( .A(n17164), .B(n17299), .Z(n17168) );
  XNOR U3245 ( .A(n1329), .B(n1492), .Z(n1333) );
  XNOR U3246 ( .A(n1710), .B(n1849), .Z(n1714) );
  XNOR U3247 ( .A(n4954), .B(n5440), .Z(n4958) );
  XNOR U3248 ( .A(n5489), .B(n5622), .Z(n5493) );
  XNOR U3249 ( .A(n5665), .B(n5799), .Z(n5669) );
  XNOR U3250 ( .A(n6024), .B(n5845), .Z(n5847) );
  XNOR U3251 ( .A(n6200), .B(n6021), .Z(n6023) );
  XNOR U3252 ( .A(n6376), .B(n6197), .Z(n6199) );
  XNOR U3253 ( .A(n6552), .B(n6373), .Z(n6375) );
  XNOR U3254 ( .A(n6728), .B(n6549), .Z(n6551) );
  XNOR U3255 ( .A(n6904), .B(n6725), .Z(n6727) );
  XNOR U3256 ( .A(n7603), .B(n7737), .Z(n7607) );
  XNOR U3257 ( .A(n7955), .B(n8089), .Z(n7959) );
  XNOR U3258 ( .A(n13977), .B(n14111), .Z(n13981) );
  XNOR U3259 ( .A(n2076), .B(n2209), .Z(n2080) );
  XNOR U3260 ( .A(n2437), .B(n2570), .Z(n2441) );
  XNOR U3261 ( .A(n2798), .B(n2931), .Z(n2802) );
  XNOR U3262 ( .A(n3159), .B(n3291), .Z(n3163) );
  XNOR U3263 ( .A(n3519), .B(n3651), .Z(n3523) );
  XNOR U3264 ( .A(n3879), .B(n4011), .Z(n3883) );
  XNOR U3265 ( .A(n4239), .B(n4371), .Z(n4243) );
  XNOR U3266 ( .A(n8312), .B(n8440), .Z(n8316) );
  XNOR U3267 ( .A(n8664), .B(n8792), .Z(n8668) );
  XNOR U3268 ( .A(n9016), .B(n9144), .Z(n9020) );
  XNOR U3269 ( .A(n13806), .B(n13934), .Z(n13810) );
  XNOR U3270 ( .A(n18786), .B(n18914), .Z(n18790) );
  XNOR U3271 ( .A(n18510), .B(n18638), .Z(n18514) );
  XNOR U3272 ( .A(n18210), .B(n18338), .Z(n18214) );
  XNOR U3273 ( .A(n17886), .B(n18014), .Z(n17890) );
  XNOR U3274 ( .A(n17535), .B(n17663), .Z(n17539) );
  XNOR U3275 ( .A(n4604), .B(n4730), .Z(n4608) );
  XNOR U3276 ( .A(n7265), .B(n7383), .Z(n7260) );
  XNOR U3277 ( .A(n9373), .B(n9495), .Z(n9377) );
  XNOR U3278 ( .A(n9725), .B(n9847), .Z(n9729) );
  XNOR U3279 ( .A(n10077), .B(n10199), .Z(n10081) );
  XNOR U3280 ( .A(n10429), .B(n10551), .Z(n10433) );
  XNOR U3281 ( .A(n10783), .B(n10929), .Z(n10787) );
  XNOR U3282 ( .A(n10992), .B(n11114), .Z(n10996) );
  XNOR U3283 ( .A(n11169), .B(n11291), .Z(n11173) );
  XNOR U3284 ( .A(n11346), .B(n11468), .Z(n11350) );
  XNOR U3285 ( .A(n11522), .B(n11644), .Z(n11526) );
  XNOR U3286 ( .A(n11698), .B(n11820), .Z(n11702) );
  XNOR U3287 ( .A(n11874), .B(n11996), .Z(n11878) );
  XNOR U3288 ( .A(n12050), .B(n12172), .Z(n12054) );
  XNOR U3289 ( .A(n12226), .B(n12348), .Z(n12230) );
  XNOR U3290 ( .A(n12402), .B(n12524), .Z(n12406) );
  XNOR U3291 ( .A(n12573), .B(n12700), .Z(n12582) );
  XNOR U3292 ( .A(n12931), .B(n13053), .Z(n12939) );
  XNOR U3293 ( .A(n13283), .B(n13405), .Z(n13287) );
  XNOR U3294 ( .A(n13635), .B(n13757), .Z(n13639) );
  XNOR U3295 ( .A(n14515), .B(n14637), .Z(n14519) );
  XNOR U3296 ( .A(n14867), .B(n14989), .Z(n14871) );
  XNOR U3297 ( .A(n15219), .B(n15341), .Z(n15223) );
  XNOR U3298 ( .A(n15571), .B(n15693), .Z(n15575) );
  XNOR U3299 ( .A(n15923), .B(n16044), .Z(n15927) );
  XNOR U3300 ( .A(n16273), .B(n16410), .Z(n16277) );
  XNOR U3301 ( .A(n16656), .B(n16476), .Z(n16478) );
  XNOR U3302 ( .A(n16833), .B(n16653), .Z(n16655) );
  XNOR U3303 ( .A(n17009), .B(n16830), .Z(n16832) );
  XNOR U3304 ( .A(n17185), .B(n17006), .Z(n17008) );
  XNOR U3305 ( .A(n17179), .B(n17296), .Z(n17183) );
  XNOR U3306 ( .A(n1344), .B(n1489), .Z(n1348) );
  XNOR U3307 ( .A(n962), .B(n1132), .Z(n967) );
  XNOR U3308 ( .A(n1725), .B(n1846), .Z(n1729) );
  XNOR U3309 ( .A(n4969), .B(n5434), .Z(n4973) );
  XNOR U3310 ( .A(n5504), .B(n5619), .Z(n5508) );
  XNOR U3311 ( .A(n5680), .B(n5796), .Z(n5684) );
  XNOR U3312 ( .A(n6039), .B(n5860), .Z(n5862) );
  XNOR U3313 ( .A(n6215), .B(n6036), .Z(n6038) );
  XNOR U3314 ( .A(n6391), .B(n6212), .Z(n6214) );
  XNOR U3315 ( .A(n6567), .B(n6388), .Z(n6390) );
  XNOR U3316 ( .A(n6743), .B(n6564), .Z(n6566) );
  XNOR U3317 ( .A(n6919), .B(n6740), .Z(n6742) );
  XNOR U3318 ( .A(n7095), .B(n6916), .Z(n6918) );
  XNOR U3319 ( .A(n7271), .B(n7092), .Z(n7094) );
  XNOR U3320 ( .A(n7447), .B(n7268), .Z(n7270) );
  XNOR U3321 ( .A(n7618), .B(n7734), .Z(n7626) );
  XNOR U3322 ( .A(n7970), .B(n8086), .Z(n7974) );
  XNOR U3323 ( .A(n14344), .B(n14460), .Z(n14348) );
  XNOR U3324 ( .A(n2091), .B(n2206), .Z(n2095) );
  XNOR U3325 ( .A(n2452), .B(n2567), .Z(n2456) );
  XNOR U3326 ( .A(n2813), .B(n2928), .Z(n2817) );
  XNOR U3327 ( .A(n3174), .B(n3288), .Z(n3178) );
  XNOR U3328 ( .A(n3534), .B(n3648), .Z(n3538) );
  XNOR U3329 ( .A(n3894), .B(n4008), .Z(n3898) );
  XNOR U3330 ( .A(n4254), .B(n4368), .Z(n4258) );
  XNOR U3331 ( .A(n8327), .B(n8437), .Z(n8331) );
  XNOR U3332 ( .A(n8679), .B(n8789), .Z(n8683) );
  XNOR U3333 ( .A(n9031), .B(n9141), .Z(n9035) );
  XNOR U3334 ( .A(n14173), .B(n14283), .Z(n14177) );
  XNOR U3335 ( .A(n19053), .B(n19163), .Z(n19057) );
  XNOR U3336 ( .A(n18801), .B(n18911), .Z(n18805) );
  XNOR U3337 ( .A(n18525), .B(n18635), .Z(n18529) );
  XNOR U3338 ( .A(n18225), .B(n18335), .Z(n18229) );
  XNOR U3339 ( .A(n17901), .B(n18011), .Z(n17905) );
  XNOR U3340 ( .A(n17550), .B(n17660), .Z(n17554) );
  XNOR U3341 ( .A(n4619), .B(n4727), .Z(n4623) );
  XNOR U3342 ( .A(n9388), .B(n9492), .Z(n9392) );
  XNOR U3343 ( .A(n9740), .B(n9844), .Z(n9744) );
  XNOR U3344 ( .A(n10092), .B(n10196), .Z(n10096) );
  XNOR U3345 ( .A(n10444), .B(n10548), .Z(n10448) );
  XNOR U3346 ( .A(n10798), .B(n10923), .Z(n10802) );
  XNOR U3347 ( .A(n11007), .B(n11111), .Z(n11011) );
  XNOR U3348 ( .A(n11184), .B(n11288), .Z(n11188) );
  XNOR U3349 ( .A(n11361), .B(n11465), .Z(n11365) );
  XNOR U3350 ( .A(n11537), .B(n11641), .Z(n11541) );
  XNOR U3351 ( .A(n11713), .B(n11817), .Z(n11717) );
  XNOR U3352 ( .A(n11889), .B(n11993), .Z(n11893) );
  XNOR U3353 ( .A(n12065), .B(n12169), .Z(n12069) );
  XNOR U3354 ( .A(n12241), .B(n12345), .Z(n12245) );
  XNOR U3355 ( .A(n12417), .B(n12521), .Z(n12421) );
  XNOR U3356 ( .A(n12593), .B(n12697), .Z(n12597) );
  XNOR U3357 ( .A(n12769), .B(n12873), .Z(n12773) );
  XNOR U3358 ( .A(n12945), .B(n13049), .Z(n12949) );
  XNOR U3359 ( .A(n13303), .B(n13124), .Z(n13126) );
  XNOR U3360 ( .A(n13302), .B(n13402), .Z(n13297) );
  XNOR U3361 ( .A(n13650), .B(n13754), .Z(n13654) );
  XNOR U3362 ( .A(n14002), .B(n14106), .Z(n14006) );
  XNOR U3363 ( .A(n14882), .B(n14986), .Z(n14886) );
  XNOR U3364 ( .A(n15234), .B(n15338), .Z(n15238) );
  XNOR U3365 ( .A(n15586), .B(n15690), .Z(n15590) );
  XNOR U3366 ( .A(n15938), .B(n16041), .Z(n15942) );
  XNOR U3367 ( .A(n16288), .B(n16404), .Z(n16292) );
  XNOR U3368 ( .A(n16671), .B(n16491), .Z(n16493) );
  XNOR U3369 ( .A(n16848), .B(n16668), .Z(n16670) );
  XNOR U3370 ( .A(n17024), .B(n16845), .Z(n16847) );
  XNOR U3371 ( .A(n17200), .B(n17021), .Z(n17023) );
  XNOR U3372 ( .A(n17194), .B(n17293), .Z(n17198) );
  XNOR U3373 ( .A(n1550), .B(n1664), .Z(n1554) );
  XNOR U3374 ( .A(n1169), .B(n1307), .Z(n1173) );
  XNOR U3375 ( .A(n788), .B(n950), .Z(n792) );
  XNOR U3376 ( .A(n4984), .B(n5428), .Z(n4988) );
  XNOR U3377 ( .A(n5519), .B(n5616), .Z(n5523) );
  XNOR U3378 ( .A(n5695), .B(n5793), .Z(n5699) );
  XNOR U3379 ( .A(n6054), .B(n5875), .Z(n5877) );
  XNOR U3380 ( .A(n6230), .B(n6051), .Z(n6053) );
  XNOR U3381 ( .A(n6406), .B(n6227), .Z(n6229) );
  XNOR U3382 ( .A(n6582), .B(n6403), .Z(n6405) );
  XNOR U3383 ( .A(n6758), .B(n6579), .Z(n6581) );
  XNOR U3384 ( .A(n6934), .B(n6755), .Z(n6757) );
  XNOR U3385 ( .A(n7110), .B(n6931), .Z(n6933) );
  XNOR U3386 ( .A(n7286), .B(n7107), .Z(n7109) );
  XNOR U3387 ( .A(n7462), .B(n7283), .Z(n7285) );
  XNOR U3388 ( .A(n7638), .B(n7459), .Z(n7461) );
  XNOR U3389 ( .A(n7814), .B(n7635), .Z(n7637) );
  XNOR U3390 ( .A(n7990), .B(n7811), .Z(n7813) );
  XNOR U3391 ( .A(n7989), .B(n8083), .Z(n7984) );
  XNOR U3392 ( .A(n14711), .B(n14809), .Z(n14715) );
  XNOR U3393 ( .A(n1745), .B(n1842), .Z(n1749) );
  XNOR U3394 ( .A(n2106), .B(n2203), .Z(n2110) );
  XNOR U3395 ( .A(n2467), .B(n2564), .Z(n2471) );
  XNOR U3396 ( .A(n2828), .B(n2925), .Z(n2832) );
  XNOR U3397 ( .A(n3189), .B(n3285), .Z(n3193) );
  XNOR U3398 ( .A(n3549), .B(n3645), .Z(n3553) );
  XNOR U3399 ( .A(n3909), .B(n4005), .Z(n3913) );
  XNOR U3400 ( .A(n4269), .B(n4365), .Z(n4273) );
  XNOR U3401 ( .A(n8342), .B(n8434), .Z(n8350) );
  XNOR U3402 ( .A(n8694), .B(n8786), .Z(n8698) );
  XNOR U3403 ( .A(n9046), .B(n9138), .Z(n9050) );
  XNOR U3404 ( .A(n14540), .B(n14632), .Z(n14544) );
  XNOR U3405 ( .A(n19500), .B(n19592), .Z(n19504) );
  XNOR U3406 ( .A(n19296), .B(n19388), .Z(n19300) );
  XNOR U3407 ( .A(n19068), .B(n19160), .Z(n19072) );
  XNOR U3408 ( .A(n18816), .B(n18908), .Z(n18820) );
  XNOR U3409 ( .A(n18540), .B(n18632), .Z(n18544) );
  XNOR U3410 ( .A(n18240), .B(n18332), .Z(n18244) );
  XNOR U3411 ( .A(n17916), .B(n18008), .Z(n17920) );
  XNOR U3412 ( .A(n17565), .B(n17657), .Z(n17569) );
  XNOR U3413 ( .A(n1013), .B(n1122), .Z(n1017) );
  XNOR U3414 ( .A(n1570), .B(n1660), .Z(n1574) );
  XNOR U3415 ( .A(n4634), .B(n4724), .Z(n4638) );
  XNOR U3416 ( .A(n9403), .B(n9489), .Z(n9407) );
  XNOR U3417 ( .A(n9755), .B(n9841), .Z(n9759) );
  XNOR U3418 ( .A(n10107), .B(n10193), .Z(n10111) );
  XNOR U3419 ( .A(n10459), .B(n10545), .Z(n10463) );
  XNOR U3420 ( .A(n10813), .B(n10917), .Z(n10817) );
  XNOR U3421 ( .A(n11022), .B(n11108), .Z(n11026) );
  XNOR U3422 ( .A(n11199), .B(n11285), .Z(n11203) );
  XNOR U3423 ( .A(n11376), .B(n11462), .Z(n11380) );
  XNOR U3424 ( .A(n11552), .B(n11638), .Z(n11556) );
  XNOR U3425 ( .A(n11728), .B(n11814), .Z(n11732) );
  XNOR U3426 ( .A(n11904), .B(n11990), .Z(n11908) );
  XNOR U3427 ( .A(n12080), .B(n12166), .Z(n12084) );
  XNOR U3428 ( .A(n12256), .B(n12342), .Z(n12260) );
  XNOR U3429 ( .A(n12432), .B(n12518), .Z(n12436) );
  XNOR U3430 ( .A(n12608), .B(n12694), .Z(n12612) );
  XNOR U3431 ( .A(n12784), .B(n12870), .Z(n12788) );
  XNOR U3432 ( .A(n12960), .B(n13046), .Z(n12964) );
  XNOR U3433 ( .A(n13136), .B(n13222), .Z(n13140) );
  XNOR U3434 ( .A(n13312), .B(n13398), .Z(n13316) );
  XNOR U3435 ( .A(n13488), .B(n13574), .Z(n13492) );
  XNOR U3436 ( .A(n13659), .B(n13750), .Z(n13668) );
  XNOR U3437 ( .A(n14017), .B(n14103), .Z(n14025) );
  XNOR U3438 ( .A(n14369), .B(n14455), .Z(n14373) );
  XNOR U3439 ( .A(n15249), .B(n15335), .Z(n15253) );
  XNOR U3440 ( .A(n15601), .B(n15687), .Z(n15605) );
  XNOR U3441 ( .A(n15953), .B(n16038), .Z(n15957) );
  XNOR U3442 ( .A(n16303), .B(n16398), .Z(n16307) );
  XNOR U3443 ( .A(n16686), .B(n16506), .Z(n16508) );
  XNOR U3444 ( .A(n16863), .B(n16683), .Z(n16685) );
  XNOR U3445 ( .A(n17039), .B(n16860), .Z(n16862) );
  XNOR U3446 ( .A(n17215), .B(n17036), .Z(n17038) );
  XNOR U3447 ( .A(n17209), .B(n17290), .Z(n17213) );
  XNOR U3448 ( .A(n1184), .B(n1304), .Z(n1188) );
  XNOR U3449 ( .A(n803), .B(n947), .Z(n807) );
  XNOR U3450 ( .A(n421), .B(n590), .Z(n426) );
  XNOR U3451 ( .A(n4999), .B(n5422), .Z(n5003) );
  XNOR U3452 ( .A(n5534), .B(n5613), .Z(n5538) );
  XNOR U3453 ( .A(n5710), .B(n5790), .Z(n5714) );
  XNOR U3454 ( .A(n6069), .B(n5890), .Z(n5892) );
  XNOR U3455 ( .A(n6245), .B(n6066), .Z(n6068) );
  XNOR U3456 ( .A(n6421), .B(n6242), .Z(n6244) );
  XNOR U3457 ( .A(n6597), .B(n6418), .Z(n6420) );
  XNOR U3458 ( .A(n6773), .B(n6594), .Z(n6596) );
  XNOR U3459 ( .A(n6949), .B(n6770), .Z(n6772) );
  XNOR U3460 ( .A(n7125), .B(n6946), .Z(n6948) );
  XNOR U3461 ( .A(n7301), .B(n7122), .Z(n7124) );
  XNOR U3462 ( .A(n7477), .B(n7298), .Z(n7300) );
  XNOR U3463 ( .A(n7653), .B(n7474), .Z(n7476) );
  XNOR U3464 ( .A(n7829), .B(n7650), .Z(n7652) );
  XNOR U3465 ( .A(n8005), .B(n7826), .Z(n7828) );
  XNOR U3466 ( .A(n8181), .B(n8002), .Z(n8004) );
  XNOR U3467 ( .A(n8357), .B(n8178), .Z(n8180) );
  XNOR U3468 ( .A(n8533), .B(n8354), .Z(n8356) );
  XNOR U3469 ( .A(n15078), .B(n15158), .Z(n15082) );
  XNOR U3470 ( .A(n2121), .B(n2200), .Z(n2125) );
  XNOR U3471 ( .A(n2482), .B(n2561), .Z(n2486) );
  XNOR U3472 ( .A(n2843), .B(n2922), .Z(n2847) );
  XNOR U3473 ( .A(n3204), .B(n3282), .Z(n3208) );
  XNOR U3474 ( .A(n3564), .B(n3642), .Z(n3568) );
  XNOR U3475 ( .A(n3924), .B(n4002), .Z(n3928) );
  XNOR U3476 ( .A(n4284), .B(n4362), .Z(n4288) );
  XNOR U3477 ( .A(n8713), .B(n8783), .Z(n8708) );
  XNOR U3478 ( .A(n9061), .B(n9135), .Z(n9065) );
  XNOR U3479 ( .A(n14907), .B(n14981), .Z(n14911) );
  XNOR U3480 ( .A(n19695), .B(n19769), .Z(n19699) );
  XNOR U3481 ( .A(n19515), .B(n19589), .Z(n19519) );
  XNOR U3482 ( .A(n19311), .B(n19385), .Z(n19315) );
  XNOR U3483 ( .A(n19083), .B(n19157), .Z(n19087) );
  XNOR U3484 ( .A(n18831), .B(n18905), .Z(n18835) );
  XNOR U3485 ( .A(n18555), .B(n18629), .Z(n18559) );
  XNOR U3486 ( .A(n18255), .B(n18329), .Z(n18259) );
  XNOR U3487 ( .A(n17931), .B(n18005), .Z(n17935) );
  XNOR U3488 ( .A(n17580), .B(n17654), .Z(n17584) );
  XNOR U3489 ( .A(n838), .B(n940), .Z(n842) );
  XNOR U3490 ( .A(n457), .B(n583), .Z(n461) );
  XNOR U3491 ( .A(n1224), .B(n1296), .Z(n1228) );
  XNOR U3492 ( .A(n1585), .B(n1657), .Z(n1589) );
  XNOR U3493 ( .A(n1946), .B(n2018), .Z(n1950) );
  XNOR U3494 ( .A(n4649), .B(n4721), .Z(n4653) );
  XNOR U3495 ( .A(n9418), .B(n9486), .Z(n9422) );
  XNOR U3496 ( .A(n9770), .B(n9838), .Z(n9774) );
  XNOR U3497 ( .A(n10122), .B(n10190), .Z(n10126) );
  XNOR U3498 ( .A(n10474), .B(n10542), .Z(n10478) );
  XNOR U3499 ( .A(n10828), .B(n10911), .Z(n10832) );
  XNOR U3500 ( .A(n11220), .B(n11040), .Z(n11042) );
  XNOR U3501 ( .A(n11397), .B(n11217), .Z(n11219) );
  XNOR U3502 ( .A(n11391), .B(n11459), .Z(n11395) );
  XNOR U3503 ( .A(n11567), .B(n11635), .Z(n11571) );
  XNOR U3504 ( .A(n11743), .B(n11811), .Z(n11747) );
  XNOR U3505 ( .A(n11919), .B(n11987), .Z(n11923) );
  XNOR U3506 ( .A(n12095), .B(n12163), .Z(n12099) );
  XNOR U3507 ( .A(n12271), .B(n12339), .Z(n12275) );
  XNOR U3508 ( .A(n12447), .B(n12515), .Z(n12451) );
  XNOR U3509 ( .A(n12623), .B(n12691), .Z(n12627) );
  XNOR U3510 ( .A(n12799), .B(n12867), .Z(n12803) );
  XNOR U3511 ( .A(n12975), .B(n13043), .Z(n12979) );
  XNOR U3512 ( .A(n13151), .B(n13219), .Z(n13155) );
  XNOR U3513 ( .A(n13327), .B(n13395), .Z(n13331) );
  XNOR U3514 ( .A(n13503), .B(n13571), .Z(n13507) );
  XNOR U3515 ( .A(n13679), .B(n13747), .Z(n13683) );
  XNOR U3516 ( .A(n13855), .B(n13923), .Z(n13859) );
  XNOR U3517 ( .A(n14031), .B(n14099), .Z(n14035) );
  XNOR U3518 ( .A(n14389), .B(n14210), .Z(n14212) );
  XNOR U3519 ( .A(n14388), .B(n14452), .Z(n14383) );
  XNOR U3520 ( .A(n14736), .B(n14804), .Z(n14740) );
  XNOR U3521 ( .A(n15616), .B(n15684), .Z(n15620) );
  XNOR U3522 ( .A(n15968), .B(n16035), .Z(n15972) );
  XNOR U3523 ( .A(n16318), .B(n16392), .Z(n16322) );
  XNOR U3524 ( .A(n16701), .B(n16521), .Z(n16523) );
  XNOR U3525 ( .A(n16878), .B(n16698), .Z(n16700) );
  XNOR U3526 ( .A(n17054), .B(n16875), .Z(n16877) );
  XNOR U3527 ( .A(n17230), .B(n17051), .Z(n17053) );
  XNOR U3528 ( .A(n17224), .B(n17287), .Z(n17228) );
  XNOR U3529 ( .A(n818), .B(n944), .Z(n822) );
  XNOR U3530 ( .A(n437), .B(n587), .Z(n441) );
  XNOR U3531 ( .A(n863), .B(n935), .Z(n867) );
  XNOR U3532 ( .A(n5014), .B(n5416), .Z(n5018) );
  XNOR U3533 ( .A(n5549), .B(n5610), .Z(n5553) );
  XNOR U3534 ( .A(n5725), .B(n5787), .Z(n5729) );
  XNOR U3535 ( .A(n6084), .B(n5905), .Z(n5907) );
  XNOR U3536 ( .A(n6260), .B(n6081), .Z(n6083) );
  XNOR U3537 ( .A(n6436), .B(n6257), .Z(n6259) );
  XNOR U3538 ( .A(n6612), .B(n6433), .Z(n6435) );
  XNOR U3539 ( .A(n6788), .B(n6609), .Z(n6611) );
  XNOR U3540 ( .A(n6964), .B(n6785), .Z(n6787) );
  XNOR U3541 ( .A(n7140), .B(n6961), .Z(n6963) );
  XNOR U3542 ( .A(n7316), .B(n7137), .Z(n7139) );
  XNOR U3543 ( .A(n7492), .B(n7313), .Z(n7315) );
  XNOR U3544 ( .A(n7668), .B(n7489), .Z(n7491) );
  XNOR U3545 ( .A(n7844), .B(n7665), .Z(n7667) );
  XNOR U3546 ( .A(n8020), .B(n7841), .Z(n7843) );
  XNOR U3547 ( .A(n8196), .B(n8017), .Z(n8019) );
  XNOR U3548 ( .A(n8372), .B(n8193), .Z(n8195) );
  XNOR U3549 ( .A(n8548), .B(n8369), .Z(n8371) );
  XNOR U3550 ( .A(n8724), .B(n8545), .Z(n8547) );
  XNOR U3551 ( .A(n8900), .B(n8721), .Z(n8723) );
  XNOR U3552 ( .A(n9076), .B(n8897), .Z(n8899) );
  XNOR U3553 ( .A(n15445), .B(n15507), .Z(n15449) );
  XNOR U3554 ( .A(n487), .B(n577), .Z(n491) );
  XNOR U3555 ( .A(n2497), .B(n2558), .Z(n2501) );
  XNOR U3556 ( .A(n2858), .B(n2919), .Z(n2862) );
  XNOR U3557 ( .A(n3219), .B(n3279), .Z(n3223) );
  XNOR U3558 ( .A(n3579), .B(n3639), .Z(n3583) );
  XNOR U3559 ( .A(n3939), .B(n3999), .Z(n3943) );
  XNOR U3560 ( .A(n4299), .B(n4359), .Z(n4303) );
  XNOR U3561 ( .A(n9256), .B(n9308), .Z(n9251) );
  XNOR U3562 ( .A(n15274), .B(n15330), .Z(n15278) );
  XNOR U3563 ( .A(n19998), .B(n20054), .Z(n20002) );
  XNOR U3564 ( .A(n19866), .B(n19922), .Z(n19870) );
  XNOR U3565 ( .A(n19710), .B(n19766), .Z(n19714) );
  XNOR U3566 ( .A(n19530), .B(n19586), .Z(n19534) );
  XNOR U3567 ( .A(n19326), .B(n19382), .Z(n19330) );
  XNOR U3568 ( .A(n19098), .B(n19154), .Z(n19102) );
  XNOR U3569 ( .A(n18846), .B(n18902), .Z(n18850) );
  XNOR U3570 ( .A(n18570), .B(n18626), .Z(n18574) );
  XNOR U3571 ( .A(n18270), .B(n18326), .Z(n18274) );
  XNOR U3572 ( .A(n17946), .B(n18002), .Z(n17950) );
  XNOR U3573 ( .A(n17595), .B(n17651), .Z(n17599) );
  XNOR U3574 ( .A(n472), .B(n580), .Z(n476) );
  XNOR U3575 ( .A(n517), .B(n571), .Z(n521) );
  XNOR U3576 ( .A(n878), .B(n932), .Z(n882) );
  XNOR U3577 ( .A(n1239), .B(n1293), .Z(n1243) );
  XNOR U3578 ( .A(n1600), .B(n1654), .Z(n1604) );
  XNOR U3579 ( .A(n1961), .B(n2015), .Z(n1965) );
  XNOR U3580 ( .A(n2322), .B(n2376), .Z(n2326) );
  XNOR U3581 ( .A(n4664), .B(n4718), .Z(n4668) );
  XNOR U3582 ( .A(n9609), .B(n9659), .Z(n9617) );
  XNOR U3583 ( .A(n9961), .B(n10011), .Z(n9965) );
  XNOR U3584 ( .A(n10489), .B(n10539), .Z(n10493) );
  XNOR U3585 ( .A(n10843), .B(n10905), .Z(n10847) );
  XNOR U3586 ( .A(n11052), .B(n11102), .Z(n11056) );
  XNOR U3587 ( .A(n11229), .B(n11279), .Z(n11233) );
  XNOR U3588 ( .A(n11406), .B(n11456), .Z(n11410) );
  XNOR U3589 ( .A(n11582), .B(n11632), .Z(n11586) );
  XNOR U3590 ( .A(n11758), .B(n11808), .Z(n11762) );
  XNOR U3591 ( .A(n11934), .B(n11984), .Z(n11938) );
  XNOR U3592 ( .A(n12110), .B(n12160), .Z(n12114) );
  XNOR U3593 ( .A(n12286), .B(n12336), .Z(n12290) );
  XNOR U3594 ( .A(n12462), .B(n12512), .Z(n12466) );
  XNOR U3595 ( .A(n12638), .B(n12688), .Z(n12642) );
  XNOR U3596 ( .A(n12814), .B(n12864), .Z(n12818) );
  XNOR U3597 ( .A(n12990), .B(n13040), .Z(n12994) );
  XNOR U3598 ( .A(n13166), .B(n13216), .Z(n13170) );
  XNOR U3599 ( .A(n13342), .B(n13392), .Z(n13346) );
  XNOR U3600 ( .A(n13518), .B(n13568), .Z(n13522) );
  XNOR U3601 ( .A(n13694), .B(n13744), .Z(n13698) );
  XNOR U3602 ( .A(n13870), .B(n13920), .Z(n13874) );
  XNOR U3603 ( .A(n14046), .B(n14096), .Z(n14050) );
  XNOR U3604 ( .A(n14222), .B(n14272), .Z(n14226) );
  XNOR U3605 ( .A(n14398), .B(n14448), .Z(n14402) );
  XNOR U3606 ( .A(n14574), .B(n14624), .Z(n14578) );
  XNOR U3607 ( .A(n14745), .B(n14800), .Z(n14754) );
  XNOR U3608 ( .A(n15103), .B(n15153), .Z(n15111) );
  XNOR U3609 ( .A(n15983), .B(n16032), .Z(n15987) );
  XNOR U3610 ( .A(n16333), .B(n16386), .Z(n16337) );
  XNOR U3611 ( .A(n16716), .B(n16536), .Z(n16538) );
  XNOR U3612 ( .A(n16893), .B(n16713), .Z(n16715) );
  XNOR U3613 ( .A(n17069), .B(n16890), .Z(n16892) );
  XNOR U3614 ( .A(n17245), .B(n17066), .Z(n17068) );
  XNOR U3615 ( .A(n17239), .B(n17284), .Z(n17243) );
  XNOR U3616 ( .A(n250), .B(n394), .Z(n262) );
  XNOR U3617 ( .A(n5029), .B(n5410), .Z(n5033) );
  XNOR U3618 ( .A(n5564), .B(n5607), .Z(n5568) );
  XNOR U3619 ( .A(n5740), .B(n5784), .Z(n5744) );
  XNOR U3620 ( .A(n6099), .B(n5920), .Z(n5922) );
  XNOR U3621 ( .A(n6275), .B(n6096), .Z(n6098) );
  XNOR U3622 ( .A(n6451), .B(n6272), .Z(n6274) );
  XNOR U3623 ( .A(n6627), .B(n6448), .Z(n6450) );
  XNOR U3624 ( .A(n6803), .B(n6624), .Z(n6626) );
  XNOR U3625 ( .A(n6979), .B(n6800), .Z(n6802) );
  XNOR U3626 ( .A(n7155), .B(n6976), .Z(n6978) );
  XNOR U3627 ( .A(n7331), .B(n7152), .Z(n7154) );
  XNOR U3628 ( .A(n7507), .B(n7328), .Z(n7330) );
  XNOR U3629 ( .A(n7683), .B(n7504), .Z(n7506) );
  XNOR U3630 ( .A(n7859), .B(n7680), .Z(n7682) );
  XNOR U3631 ( .A(n8035), .B(n7856), .Z(n7858) );
  XNOR U3632 ( .A(n8211), .B(n8032), .Z(n8034) );
  XNOR U3633 ( .A(n8387), .B(n8208), .Z(n8210) );
  XNOR U3634 ( .A(n8563), .B(n8384), .Z(n8386) );
  XNOR U3635 ( .A(n8739), .B(n8560), .Z(n8562) );
  XNOR U3636 ( .A(n8915), .B(n8736), .Z(n8738) );
  XNOR U3637 ( .A(n9091), .B(n8912), .Z(n8914) );
  XNOR U3638 ( .A(n9267), .B(n9088), .Z(n9090) );
  XNOR U3639 ( .A(n9443), .B(n9264), .Z(n9266) );
  XNOR U3640 ( .A(n9619), .B(n9440), .Z(n9442) );
  XNOR U3641 ( .A(n10318), .B(n10362), .Z(n10322) );
  XNOR U3642 ( .A(n15812), .B(n15856), .Z(n15816) );
  XNOR U3643 ( .A(n502), .B(n574), .Z(n506) );
  XNOR U3644 ( .A(n2873), .B(n2916), .Z(n2877) );
  XNOR U3645 ( .A(n3234), .B(n3276), .Z(n3238) );
  XNOR U3646 ( .A(n3594), .B(n3636), .Z(n3598) );
  XNOR U3647 ( .A(n3954), .B(n3996), .Z(n3958) );
  XNOR U3648 ( .A(n4314), .B(n4356), .Z(n4318) );
  XNOR U3649 ( .A(n15641), .B(n15679), .Z(n15645) );
  XNOR U3650 ( .A(n20121), .B(n20159), .Z(n20125) );
  XNOR U3651 ( .A(n20013), .B(n20051), .Z(n20017) );
  XNOR U3652 ( .A(n19881), .B(n19919), .Z(n19885) );
  XNOR U3653 ( .A(n19725), .B(n19763), .Z(n19729) );
  XNOR U3654 ( .A(n19545), .B(n19583), .Z(n19549) );
  XNOR U3655 ( .A(n19341), .B(n19379), .Z(n19345) );
  XNOR U3656 ( .A(n19113), .B(n19151), .Z(n19117) );
  XNOR U3657 ( .A(n18861), .B(n18899), .Z(n18865) );
  XNOR U3658 ( .A(n18585), .B(n18623), .Z(n18589) );
  XNOR U3659 ( .A(n18285), .B(n18323), .Z(n18289) );
  XNOR U3660 ( .A(n17961), .B(n17999), .Z(n17965) );
  XNOR U3661 ( .A(n17610), .B(n17648), .Z(n17614) );
  XNOR U3662 ( .A(n532), .B(n568), .Z(n536) );
  XNOR U3663 ( .A(n893), .B(n929), .Z(n897) );
  XNOR U3664 ( .A(n1254), .B(n1290), .Z(n1258) );
  XNOR U3665 ( .A(n1615), .B(n1651), .Z(n1619) );
  XNOR U3666 ( .A(n1976), .B(n2012), .Z(n1980) );
  XNOR U3667 ( .A(n2337), .B(n2373), .Z(n2341) );
  XNOR U3668 ( .A(n2698), .B(n2734), .Z(n2702) );
  XNOR U3669 ( .A(n4679), .B(n4715), .Z(n4683) );
  XNOR U3670 ( .A(n9980), .B(n10008), .Z(n9975) );
  XNOR U3671 ( .A(n10858), .B(n10899), .Z(n10862) );
  XNOR U3672 ( .A(n11250), .B(n11070), .Z(n11072) );
  XNOR U3673 ( .A(n11427), .B(n11247), .Z(n11249) );
  XNOR U3674 ( .A(n11603), .B(n11424), .Z(n11426) );
  XNOR U3675 ( .A(n11597), .B(n11629), .Z(n11601) );
  XNOR U3676 ( .A(n11773), .B(n11805), .Z(n11777) );
  XNOR U3677 ( .A(n11949), .B(n11981), .Z(n11953) );
  XNOR U3678 ( .A(n12125), .B(n12157), .Z(n12129) );
  XNOR U3679 ( .A(n12301), .B(n12333), .Z(n12305) );
  XNOR U3680 ( .A(n12477), .B(n12509), .Z(n12481) );
  XNOR U3681 ( .A(n12653), .B(n12685), .Z(n12657) );
  XNOR U3682 ( .A(n12829), .B(n12861), .Z(n12833) );
  XNOR U3683 ( .A(n13005), .B(n13037), .Z(n13009) );
  XNOR U3684 ( .A(n13181), .B(n13213), .Z(n13185) );
  XNOR U3685 ( .A(n13357), .B(n13389), .Z(n13361) );
  XNOR U3686 ( .A(n13533), .B(n13565), .Z(n13537) );
  XNOR U3687 ( .A(n13709), .B(n13741), .Z(n13713) );
  XNOR U3688 ( .A(n13885), .B(n13917), .Z(n13889) );
  XNOR U3689 ( .A(n14061), .B(n14093), .Z(n14065) );
  XNOR U3690 ( .A(n14237), .B(n14269), .Z(n14241) );
  XNOR U3691 ( .A(n14413), .B(n14445), .Z(n14417) );
  XNOR U3692 ( .A(n14589), .B(n14621), .Z(n14593) );
  XNOR U3693 ( .A(n14765), .B(n14797), .Z(n14769) );
  XNOR U3694 ( .A(n14941), .B(n14973), .Z(n14945) );
  XNOR U3695 ( .A(n15117), .B(n15149), .Z(n15121) );
  XNOR U3696 ( .A(n15475), .B(n15296), .Z(n15298) );
  XNOR U3697 ( .A(n15474), .B(n15502), .Z(n15469) );
  XNOR U3698 ( .A(n16348), .B(n16380), .Z(n16352) );
  XNOR U3699 ( .A(n16731), .B(n16551), .Z(n16553) );
  XNOR U3700 ( .A(n16908), .B(n16728), .Z(n16730) );
  XNOR U3701 ( .A(n17084), .B(n16905), .Z(n16907) );
  XNOR U3702 ( .A(n17260), .B(n17081), .Z(n17083) );
  XNOR U3703 ( .A(n17254), .B(n17281), .Z(n17258) );
  XNOR U3704 ( .A(n5044), .B(n5404), .Z(n5048) );
  XNOR U3705 ( .A(n5579), .B(n5604), .Z(n5583) );
  XNOR U3706 ( .A(n5755), .B(n5781), .Z(n5759) );
  XNOR U3707 ( .A(n6114), .B(n5935), .Z(n5937) );
  XNOR U3708 ( .A(n6290), .B(n6111), .Z(n6113) );
  XNOR U3709 ( .A(n6466), .B(n6287), .Z(n6289) );
  XNOR U3710 ( .A(n6642), .B(n6463), .Z(n6465) );
  XNOR U3711 ( .A(n6818), .B(n6639), .Z(n6641) );
  XNOR U3712 ( .A(n6994), .B(n6815), .Z(n6817) );
  XNOR U3713 ( .A(n7170), .B(n6991), .Z(n6993) );
  XNOR U3714 ( .A(n7346), .B(n7167), .Z(n7169) );
  XNOR U3715 ( .A(n7522), .B(n7343), .Z(n7345) );
  XNOR U3716 ( .A(n7698), .B(n7519), .Z(n7521) );
  XNOR U3717 ( .A(n7874), .B(n7695), .Z(n7697) );
  XNOR U3718 ( .A(n8050), .B(n7871), .Z(n7873) );
  XNOR U3719 ( .A(n8226), .B(n8047), .Z(n8049) );
  XNOR U3720 ( .A(n8402), .B(n8223), .Z(n8225) );
  XNOR U3721 ( .A(n8578), .B(n8399), .Z(n8401) );
  XNOR U3722 ( .A(n8754), .B(n8575), .Z(n8577) );
  XNOR U3723 ( .A(n8930), .B(n8751), .Z(n8753) );
  XNOR U3724 ( .A(n9106), .B(n8927), .Z(n8929) );
  XNOR U3725 ( .A(n9282), .B(n9103), .Z(n9105) );
  XNOR U3726 ( .A(n9458), .B(n9279), .Z(n9281) );
  XNOR U3727 ( .A(n9634), .B(n9455), .Z(n9457) );
  XNOR U3728 ( .A(n9810), .B(n9631), .Z(n9633) );
  XNOR U3729 ( .A(n9986), .B(n9807), .Z(n9809) );
  XNOR U3730 ( .A(n10162), .B(n9983), .Z(n9985) );
  XNOR U3731 ( .A(n10333), .B(n10359), .Z(n10341) );
  XNOR U3732 ( .A(n10685), .B(n10713), .Z(n10689) );
  XNOR U3733 ( .A(n16178), .B(n16203), .Z(n16182) );
  XNOR U3734 ( .A(n3249), .B(n3273), .Z(n3253) );
  XNOR U3735 ( .A(n3789), .B(n3813), .Z(n3793) );
  XNOR U3736 ( .A(n4329), .B(n4353), .Z(n4333) );
  XNOR U3737 ( .A(n16008), .B(n16027), .Z(n16013) );
  XNOR U3738 ( .A(n20253), .B(n20273), .Z(n20262) );
  XNOR U3739 ( .A(n20181), .B(n20201), .Z(n20190) );
  XNOR U3740 ( .A(n20085), .B(n20105), .Z(n20094) );
  XNOR U3741 ( .A(n19965), .B(n19985), .Z(n19974) );
  XNOR U3742 ( .A(n19821), .B(n19841), .Z(n19830) );
  XNOR U3743 ( .A(n19653), .B(n19673), .Z(n19662) );
  XNOR U3744 ( .A(n19461), .B(n19481), .Z(n19470) );
  XNOR U3745 ( .A(n19245), .B(n19265), .Z(n19254) );
  XNOR U3746 ( .A(n19005), .B(n19025), .Z(n19014) );
  XNOR U3747 ( .A(n18741), .B(n18761), .Z(n18750) );
  XNOR U3748 ( .A(n18453), .B(n18473), .Z(n18462) );
  XNOR U3749 ( .A(n18141), .B(n18161), .Z(n18150) );
  XNOR U3750 ( .A(n17805), .B(n17825), .Z(n17814) );
  XNOR U3751 ( .A(n17440), .B(n17463), .Z(n17445) );
  XNOR U3752 ( .A(n547), .B(n565), .Z(n556) );
  XNOR U3753 ( .A(n908), .B(n926), .Z(n917) );
  XNOR U3754 ( .A(n1269), .B(n1287), .Z(n1278) );
  XNOR U3755 ( .A(n1630), .B(n1648), .Z(n1639) );
  XNOR U3756 ( .A(n1991), .B(n2009), .Z(n2000) );
  XNOR U3757 ( .A(n2352), .B(n2370), .Z(n2361) );
  XNOR U3758 ( .A(n2713), .B(n2731), .Z(n2722) );
  XNOR U3759 ( .A(n3074), .B(n3092), .Z(n3083) );
  XNOR U3760 ( .A(n3614), .B(n3632), .Z(n3623) );
  XNOR U3761 ( .A(n4154), .B(n4172), .Z(n4163) );
  XNOR U3762 ( .A(n4694), .B(n4712), .Z(n4703) );
  XNOR U3763 ( .A(n5771), .B(n5592), .Z(n5594) );
  XNOR U3764 ( .A(n11082), .B(n11087), .Z(n10891) );
  XNOR U3765 ( .A(n11263), .B(n11262), .Z(n11092) );
  XNOR U3766 ( .A(n11436), .B(n11441), .Z(n11271) );
  XNOR U3767 ( .A(n11616), .B(n11615), .Z(n11446) );
  XNOR U3768 ( .A(n11788), .B(n11793), .Z(n11624) );
  XNOR U3769 ( .A(n11968), .B(n11967), .Z(n11798) );
  XNOR U3770 ( .A(n12140), .B(n12145), .Z(n11976) );
  XNOR U3771 ( .A(n12320), .B(n12319), .Z(n12150) );
  XNOR U3772 ( .A(n12492), .B(n12497), .Z(n12328) );
  XNOR U3773 ( .A(n12672), .B(n12671), .Z(n12502) );
  XNOR U3774 ( .A(n12844), .B(n12849), .Z(n12680) );
  XNOR U3775 ( .A(n13024), .B(n13023), .Z(n12854) );
  XNOR U3776 ( .A(n13196), .B(n13201), .Z(n13032) );
  XNOR U3777 ( .A(n13376), .B(n13375), .Z(n13206) );
  XNOR U3778 ( .A(n13548), .B(n13553), .Z(n13384) );
  XNOR U3779 ( .A(n13728), .B(n13727), .Z(n13558) );
  XNOR U3780 ( .A(n13900), .B(n13905), .Z(n13736) );
  XNOR U3781 ( .A(n14080), .B(n14079), .Z(n13910) );
  XNOR U3782 ( .A(n14252), .B(n14257), .Z(n14088) );
  XNOR U3783 ( .A(n14432), .B(n14431), .Z(n14262) );
  XNOR U3784 ( .A(n14604), .B(n14609), .Z(n14440) );
  XNOR U3785 ( .A(n14784), .B(n14783), .Z(n14614) );
  XNOR U3786 ( .A(n14956), .B(n14961), .Z(n14792) );
  XNOR U3787 ( .A(n15136), .B(n15135), .Z(n14966) );
  XNOR U3788 ( .A(n15308), .B(n15313), .Z(n15144) );
  XNOR U3789 ( .A(n15488), .B(n15487), .Z(n15318) );
  XNOR U3790 ( .A(n15660), .B(n15665), .Z(n15496) );
  XNOR U3791 ( .A(n15840), .B(n15839), .Z(n15670) );
  XNOR U3792 ( .A(n16567), .B(n16566), .Z(n16367) );
  XNOR U3793 ( .A(n16740), .B(n16745), .Z(n16575) );
  XNOR U3794 ( .A(n16921), .B(n16920), .Z(n16750) );
  XNOR U3795 ( .A(n17093), .B(n17098), .Z(n16929) );
  XNOR U3796 ( .A(n17273), .B(n17272), .Z(n17103) );
  XOR U3797 ( .A(n5063), .B(n5399), .Z(n5057) );
  XOR U3798 ( .A(n5947), .B(n5954), .Z(n5952) );
  XOR U3799 ( .A(n6123), .B(n6130), .Z(n6128) );
  XOR U3800 ( .A(n6299), .B(n6306), .Z(n6304) );
  XOR U3801 ( .A(n6475), .B(n6482), .Z(n6480) );
  XOR U3802 ( .A(n6651), .B(n6658), .Z(n6656) );
  XOR U3803 ( .A(n6827), .B(n6834), .Z(n6832) );
  XOR U3804 ( .A(n7003), .B(n7010), .Z(n7008) );
  XOR U3805 ( .A(n7179), .B(n7186), .Z(n7184) );
  XOR U3806 ( .A(n7355), .B(n7362), .Z(n7360) );
  XOR U3807 ( .A(n7531), .B(n7538), .Z(n7536) );
  XOR U3808 ( .A(n7707), .B(n7714), .Z(n7712) );
  XOR U3809 ( .A(n7883), .B(n7890), .Z(n7888) );
  XOR U3810 ( .A(n8059), .B(n8066), .Z(n8064) );
  XOR U3811 ( .A(n8235), .B(n8242), .Z(n8240) );
  XOR U3812 ( .A(n8411), .B(n8418), .Z(n8416) );
  XOR U3813 ( .A(n8587), .B(n8594), .Z(n8592) );
  XOR U3814 ( .A(n8763), .B(n8770), .Z(n8768) );
  XOR U3815 ( .A(n8939), .B(n8946), .Z(n8944) );
  XOR U3816 ( .A(n9115), .B(n9122), .Z(n9120) );
  XOR U3817 ( .A(n9291), .B(n9298), .Z(n9296) );
  XOR U3818 ( .A(n9467), .B(n9474), .Z(n9472) );
  XOR U3819 ( .A(n9643), .B(n9650), .Z(n9648) );
  XOR U3820 ( .A(n9819), .B(n9826), .Z(n9824) );
  XOR U3821 ( .A(n9995), .B(n10002), .Z(n10000) );
  XOR U3822 ( .A(n10171), .B(n10178), .Z(n10176) );
  XOR U3823 ( .A(n10347), .B(n10354), .Z(n10352) );
  XOR U3824 ( .A(n10703), .B(n10707), .Z(n10699) );
  XOR U3825 ( .A(n10887), .B(n10892), .Z(n10880) );
  XOR U3826 ( .A(n16365), .B(n16370), .Z(n16196) );
  XNOR U3827 ( .A(n20300), .B(n20297), .Z(n20299) );
  NAND U3828 ( .A(n1280), .B(n1279), .Z(n1098) );
  NAND U3829 ( .A(n2002), .B(n2001), .Z(n1820) );
  NAND U3830 ( .A(n2724), .B(n2723), .Z(n2542) );
  XNOR U3831 ( .A(n3264), .B(n3266), .Z(n3265) );
  XNOR U3832 ( .A(n3804), .B(n3806), .Z(n3805) );
  XNOR U3833 ( .A(n4344), .B(n4346), .Z(n4345) );
  XNOR U3834 ( .A(n4884), .B(n4886), .Z(n4885) );
  XOR U3835 ( .A(n5071), .B(n5), .Z(n5070) );
  NAND U3836 ( .A(n558), .B(n557), .Z(n311) );
  XNOR U3837 ( .A(n1), .B(n2), .Z(swire[99]) );
  XOR U3838 ( .A(n3), .B(n4), .Z(swire[98]) );
  XNOR U3839 ( .A(n5), .B(n6), .Z(swire[97]) );
  XNOR U3840 ( .A(n7), .B(n8), .Z(swire[96]) );
  XOR U3841 ( .A(n9), .B(n10), .Z(swire[95]) );
  XOR U3842 ( .A(n11), .B(n12), .Z(swire[94]) );
  XOR U3843 ( .A(n13), .B(n14), .Z(swire[93]) );
  XOR U3844 ( .A(n15), .B(n16), .Z(swire[92]) );
  XOR U3845 ( .A(n17), .B(n18), .Z(swire[91]) );
  XOR U3846 ( .A(n19), .B(n20), .Z(swire[90]) );
  XOR U3847 ( .A(n21), .B(n22), .Z(swire[89]) );
  XOR U3848 ( .A(n23), .B(n24), .Z(swire[88]) );
  XOR U3849 ( .A(n25), .B(n26), .Z(swire[87]) );
  XOR U3850 ( .A(n27), .B(n28), .Z(swire[86]) );
  XOR U3851 ( .A(n29), .B(n30), .Z(swire[85]) );
  XOR U3852 ( .A(n31), .B(n32), .Z(swire[84]) );
  XOR U3853 ( .A(n33), .B(n34), .Z(swire[83]) );
  XOR U3854 ( .A(n35), .B(n36), .Z(swire[82]) );
  XOR U3855 ( .A(n37), .B(n38), .Z(swire[81]) );
  XOR U3856 ( .A(n39), .B(n40), .Z(swire[80]) );
  XOR U3857 ( .A(n41), .B(n42), .Z(swire[79]) );
  XOR U3858 ( .A(n43), .B(n44), .Z(swire[78]) );
  XOR U3859 ( .A(n45), .B(n46), .Z(swire[77]) );
  XOR U3860 ( .A(n47), .B(n48), .Z(swire[76]) );
  XOR U3861 ( .A(n49), .B(n50), .Z(swire[75]) );
  XOR U3862 ( .A(n51), .B(n52), .Z(swire[74]) );
  XOR U3863 ( .A(n53), .B(n54), .Z(swire[73]) );
  XOR U3864 ( .A(n55), .B(n56), .Z(swire[72]) );
  XOR U3865 ( .A(n57), .B(n58), .Z(swire[71]) );
  XOR U3866 ( .A(n59), .B(n60), .Z(swire[70]) );
  XOR U3867 ( .A(n61), .B(n62), .Z(swire[69]) );
  XOR U3868 ( .A(n63), .B(n64), .Z(swire[68]) );
  XOR U3869 ( .A(n65), .B(n66), .Z(swire[67]) );
  XOR U3870 ( .A(n67), .B(n68), .Z(swire[66]) );
  XOR U3871 ( .A(n69), .B(n70), .Z(swire[65]) );
  XOR U3872 ( .A(n71), .B(n72), .Z(swire[64]) );
  XOR U3873 ( .A(n73), .B(n74), .Z(swire[63]) );
  XOR U3874 ( .A(n75), .B(n76), .Z(swire[62]) );
  XOR U3875 ( .A(n77), .B(n78), .Z(swire[61]) );
  XOR U3876 ( .A(n79), .B(n80), .Z(swire[60]) );
  XOR U3877 ( .A(n81), .B(n82), .Z(swire[59]) );
  XOR U3878 ( .A(n83), .B(n84), .Z(swire[58]) );
  XOR U3879 ( .A(n85), .B(n86), .Z(swire[57]) );
  XOR U3880 ( .A(n87), .B(n88), .Z(swire[56]) );
  XOR U3881 ( .A(n89), .B(n90), .Z(swire[55]) );
  XOR U3882 ( .A(n91), .B(n92), .Z(swire[54]) );
  XOR U3883 ( .A(n93), .B(n94), .Z(swire[53]) );
  XOR U3884 ( .A(n95), .B(n96), .Z(swire[52]) );
  XOR U3885 ( .A(n97), .B(n98), .Z(swire[51]) );
  XOR U3886 ( .A(n99), .B(n100), .Z(swire[50]) );
  XOR U3887 ( .A(n101), .B(n102), .Z(swire[49]) );
  XOR U3888 ( .A(n103), .B(n104), .Z(swire[48]) );
  XOR U3889 ( .A(n105), .B(n106), .Z(swire[47]) );
  XOR U3890 ( .A(n107), .B(n108), .Z(swire[46]) );
  XOR U3891 ( .A(n109), .B(n110), .Z(swire[45]) );
  XOR U3892 ( .A(n111), .B(n112), .Z(swire[44]) );
  XOR U3893 ( .A(n113), .B(n114), .Z(swire[43]) );
  XOR U3894 ( .A(n115), .B(n116), .Z(swire[42]) );
  XOR U3895 ( .A(n117), .B(n118), .Z(swire[41]) );
  XOR U3896 ( .A(n119), .B(n120), .Z(swire[40]) );
  XOR U3897 ( .A(n121), .B(n122), .Z(swire[39]) );
  XOR U3898 ( .A(n123), .B(n124), .Z(swire[38]) );
  XOR U3899 ( .A(n125), .B(n126), .Z(swire[37]) );
  XOR U3900 ( .A(n127), .B(n128), .Z(swire[36]) );
  XOR U3901 ( .A(n129), .B(n130), .Z(swire[35]) );
  XOR U3902 ( .A(n131), .B(n132), .Z(swire[34]) );
  XOR U3903 ( .A(n133), .B(n134), .Z(swire[33]) );
  XOR U3904 ( .A(n135), .B(n136), .Z(swire[32]) );
  XOR U3905 ( .A(n137), .B(n138), .Z(swire[127]) );
  XOR U3906 ( .A(n139), .B(n140), .Z(n138) );
  XOR U3907 ( .A(n141), .B(n142), .Z(n140) );
  XOR U3908 ( .A(n143), .B(n144), .Z(n142) );
  XOR U3909 ( .A(n145), .B(n146), .Z(n144) );
  XNOR U3910 ( .A(n147), .B(n148), .Z(n146) );
  AND U3911 ( .A(b[1]), .B(a[126]), .Z(n148) );
  XOR U3912 ( .A(n149), .B(n150), .Z(n145) );
  XOR U3913 ( .A(n151), .B(n152), .Z(n150) );
  XOR U3914 ( .A(n153), .B(n154), .Z(n152) );
  AND U3915 ( .A(b[7]), .B(a[120]), .Z(n154) );
  AND U3916 ( .A(b[8]), .B(a[119]), .Z(n153) );
  XOR U3917 ( .A(n155), .B(n156), .Z(n151) );
  XOR U3918 ( .A(n157), .B(n158), .Z(n156) );
  XOR U3919 ( .A(n159), .B(n160), .Z(n158) );
  XOR U3920 ( .A(n161), .B(n162), .Z(n160) );
  XOR U3921 ( .A(n163), .B(n164), .Z(n162) );
  XOR U3922 ( .A(n165), .B(n166), .Z(n164) );
  AND U3923 ( .A(b[20]), .B(a[107]), .Z(n166) );
  AND U3924 ( .A(b[25]), .B(a[102]), .Z(n165) );
  XOR U3925 ( .A(n167), .B(n168), .Z(n163) );
  AND U3926 ( .A(b[26]), .B(a[101]), .Z(n168) );
  AND U3927 ( .A(b[27]), .B(a[100]), .Z(n167) );
  XOR U3928 ( .A(n169), .B(n170), .Z(n161) );
  XOR U3929 ( .A(n171), .B(n172), .Z(n170) );
  AND U3930 ( .A(b[28]), .B(a[99]), .Z(n172) );
  AND U3931 ( .A(b[29]), .B(a[98]), .Z(n171) );
  XOR U3932 ( .A(n173), .B(n174), .Z(n169) );
  AND U3933 ( .A(b[30]), .B(a[97]), .Z(n174) );
  AND U3934 ( .A(b[31]), .B(a[96]), .Z(n173) );
  AND U3935 ( .A(b[13]), .B(a[114]), .Z(n159) );
  XOR U3936 ( .A(n175), .B(n176), .Z(n157) );
  AND U3937 ( .A(b[14]), .B(a[113]), .Z(n176) );
  AND U3938 ( .A(b[19]), .B(a[108]), .Z(n175) );
  XOR U3939 ( .A(n177), .B(n178), .Z(n155) );
  XOR U3940 ( .A(n179), .B(n180), .Z(n178) );
  AND U3941 ( .A(b[21]), .B(a[106]), .Z(n180) );
  AND U3942 ( .A(b[22]), .B(a[105]), .Z(n179) );
  XOR U3943 ( .A(n181), .B(n182), .Z(n177) );
  AND U3944 ( .A(b[23]), .B(a[104]), .Z(n182) );
  AND U3945 ( .A(b[24]), .B(a[103]), .Z(n181) );
  XOR U3946 ( .A(n183), .B(n184), .Z(n149) );
  XOR U3947 ( .A(n185), .B(n186), .Z(n184) );
  AND U3948 ( .A(b[15]), .B(a[112]), .Z(n186) );
  AND U3949 ( .A(b[16]), .B(a[111]), .Z(n185) );
  XOR U3950 ( .A(n187), .B(n188), .Z(n183) );
  AND U3951 ( .A(b[17]), .B(a[110]), .Z(n188) );
  AND U3952 ( .A(b[18]), .B(a[109]), .Z(n187) );
  XOR U3953 ( .A(n189), .B(n190), .Z(n143) );
  XOR U3954 ( .A(n191), .B(n192), .Z(n190) );
  AND U3955 ( .A(b[9]), .B(a[118]), .Z(n192) );
  AND U3956 ( .A(b[10]), .B(a[117]), .Z(n191) );
  XOR U3957 ( .A(n193), .B(n194), .Z(n189) );
  AND U3958 ( .A(b[11]), .B(a[116]), .Z(n194) );
  AND U3959 ( .A(b[12]), .B(a[115]), .Z(n193) );
  AND U3960 ( .A(a[127]), .B(b[0]), .Z(n141) );
  XNOR U3961 ( .A(n195), .B(n147), .Z(n139) );
  OR U3962 ( .A(n196), .B(n197), .Z(n147) );
  AND U3963 ( .A(b[2]), .B(a[125]), .Z(n195) );
  XOR U3964 ( .A(n198), .B(n199), .Z(n137) );
  XOR U3965 ( .A(n200), .B(n201), .Z(n199) );
  AND U3966 ( .A(b[3]), .B(a[124]), .Z(n201) );
  AND U3967 ( .A(b[4]), .B(a[123]), .Z(n200) );
  XOR U3968 ( .A(n202), .B(n203), .Z(n198) );
  AND U3969 ( .A(b[5]), .B(a[122]), .Z(n203) );
  AND U3970 ( .A(b[6]), .B(a[121]), .Z(n202) );
  XOR U3971 ( .A(n196), .B(n197), .Z(swire[126]) );
  XOR U3972 ( .A(n204), .B(n205), .Z(n197) );
  XNOR U3973 ( .A(n206), .B(n207), .Z(n205) );
  XOR U3974 ( .A(n208), .B(n209), .Z(n207) );
  XOR U3975 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U3976 ( .A(n212), .B(n206), .Z(n211) );
  XOR U3977 ( .A(n213), .B(n214), .Z(n210) );
  XOR U3978 ( .A(n215), .B(n216), .Z(n214) );
  XOR U3979 ( .A(n217), .B(n218), .Z(n216) );
  XOR U3980 ( .A(n219), .B(n220), .Z(n218) );
  AND U3981 ( .A(b[7]), .B(a[119]), .Z(n219) );
  XOR U3982 ( .A(n221), .B(n222), .Z(n217) );
  XOR U3983 ( .A(n223), .B(n224), .Z(n222) );
  XOR U3984 ( .A(n225), .B(n226), .Z(n224) );
  XOR U3985 ( .A(n227), .B(n228), .Z(n226) );
  AND U3986 ( .A(b[13]), .B(a[113]), .Z(n227) );
  XOR U3987 ( .A(n229), .B(n230), .Z(n225) );
  XOR U3988 ( .A(n231), .B(n232), .Z(n230) );
  XOR U3989 ( .A(n233), .B(n234), .Z(n232) );
  XOR U3990 ( .A(n235), .B(n236), .Z(n234) );
  AND U3991 ( .A(b[19]), .B(a[107]), .Z(n235) );
  XOR U3992 ( .A(n237), .B(n238), .Z(n233) );
  AND U3993 ( .A(b[24]), .B(a[102]), .Z(n237) );
  XOR U3994 ( .A(n236), .B(n239), .Z(n231) );
  XOR U3995 ( .A(n238), .B(n240), .Z(n239) );
  XOR U3996 ( .A(n241), .B(n242), .Z(n240) );
  XOR U3997 ( .A(n243), .B(n244), .Z(n242) );
  XOR U3998 ( .A(n245), .B(n246), .Z(n244) );
  XOR U3999 ( .A(n247), .B(n245), .Z(n246) );
  AND U4000 ( .A(b[25]), .B(a[101]), .Z(n247) );
  XOR U4001 ( .A(n248), .B(n249), .Z(n245) );
  ANDN U4002 ( .B(n250), .A(n251), .Z(n248) );
  XOR U4003 ( .A(n252), .B(n253), .Z(n243) );
  AND U4004 ( .A(b[26]), .B(a[100]), .Z(n253) );
  AND U4005 ( .A(b[27]), .B(a[99]), .Z(n252) );
  XOR U4006 ( .A(n254), .B(n255), .Z(n241) );
  XOR U4007 ( .A(n256), .B(n257), .Z(n255) );
  AND U4008 ( .A(b[28]), .B(a[98]), .Z(n257) );
  AND U4009 ( .A(b[29]), .B(a[97]), .Z(n256) );
  XOR U4010 ( .A(n258), .B(n259), .Z(n254) );
  AND U4011 ( .A(b[30]), .B(a[96]), .Z(n259) );
  AND U4012 ( .A(b[31]), .B(a[95]), .Z(n258) );
  XOR U4013 ( .A(n260), .B(n261), .Z(n238) );
  AND U4014 ( .A(n262), .B(n263), .Z(n260) );
  XOR U4015 ( .A(n264), .B(n265), .Z(n236) );
  ANDN U4016 ( .B(n266), .A(n267), .Z(n264) );
  XOR U4017 ( .A(n268), .B(n269), .Z(n229) );
  XOR U4018 ( .A(n270), .B(n271), .Z(n269) );
  AND U4019 ( .A(b[20]), .B(a[106]), .Z(n271) );
  AND U4020 ( .A(b[21]), .B(a[105]), .Z(n270) );
  XOR U4021 ( .A(n272), .B(n273), .Z(n268) );
  AND U4022 ( .A(b[22]), .B(a[104]), .Z(n273) );
  AND U4023 ( .A(b[23]), .B(a[103]), .Z(n272) );
  XOR U4024 ( .A(n274), .B(n228), .Z(n223) );
  XOR U4025 ( .A(n275), .B(n276), .Z(n228) );
  ANDN U4026 ( .B(n277), .A(n278), .Z(n275) );
  AND U4027 ( .A(b[14]), .B(a[112]), .Z(n274) );
  XOR U4028 ( .A(n279), .B(n280), .Z(n221) );
  XOR U4029 ( .A(n281), .B(n282), .Z(n280) );
  AND U4030 ( .A(b[15]), .B(a[111]), .Z(n282) );
  AND U4031 ( .A(b[16]), .B(a[110]), .Z(n281) );
  XOR U4032 ( .A(n283), .B(n284), .Z(n279) );
  AND U4033 ( .A(b[17]), .B(a[109]), .Z(n284) );
  AND U4034 ( .A(b[18]), .B(a[108]), .Z(n283) );
  XOR U4035 ( .A(n285), .B(n220), .Z(n215) );
  XOR U4036 ( .A(n286), .B(n287), .Z(n220) );
  ANDN U4037 ( .B(n288), .A(n289), .Z(n286) );
  AND U4038 ( .A(b[8]), .B(a[118]), .Z(n285) );
  XOR U4039 ( .A(n290), .B(n291), .Z(n213) );
  XOR U4040 ( .A(n292), .B(n293), .Z(n291) );
  AND U4041 ( .A(b[9]), .B(a[117]), .Z(n293) );
  AND U4042 ( .A(b[10]), .B(a[116]), .Z(n292) );
  XOR U4043 ( .A(n294), .B(n295), .Z(n290) );
  AND U4044 ( .A(b[11]), .B(a[115]), .Z(n295) );
  AND U4045 ( .A(b[12]), .B(a[114]), .Z(n294) );
  XOR U4046 ( .A(n296), .B(n297), .Z(n208) );
  XOR U4047 ( .A(n298), .B(n299), .Z(n297) );
  AND U4048 ( .A(b[3]), .B(a[123]), .Z(n299) );
  AND U4049 ( .A(b[4]), .B(a[122]), .Z(n298) );
  XOR U4050 ( .A(n300), .B(n301), .Z(n296) );
  AND U4051 ( .A(b[5]), .B(a[121]), .Z(n301) );
  AND U4052 ( .A(b[6]), .B(a[120]), .Z(n300) );
  XOR U4053 ( .A(n302), .B(n303), .Z(n206) );
  OR U4054 ( .A(n304), .B(n305), .Z(n303) );
  XOR U4055 ( .A(n306), .B(n307), .Z(n204) );
  XNOR U4056 ( .A(n308), .B(n212), .Z(n307) );
  NANDN U4057 ( .A(n309), .B(n310), .Z(n212) );
  AND U4058 ( .A(b[2]), .B(a[124]), .Z(n308) );
  AND U4059 ( .A(b[1]), .B(a[125]), .Z(n306) );
  NAND U4060 ( .A(a[126]), .B(b[0]), .Z(n196) );
  XNOR U4061 ( .A(n311), .B(n312), .Z(swire[125]) );
  XOR U4062 ( .A(n310), .B(n313), .Z(n312) );
  XOR U4063 ( .A(n309), .B(n311), .Z(n313) );
  NAND U4064 ( .A(a[125]), .B(b[0]), .Z(n309) );
  XOR U4065 ( .A(n304), .B(n305), .Z(n310) );
  XOR U4066 ( .A(n302), .B(n314), .Z(n305) );
  NAND U4067 ( .A(b[1]), .B(a[124]), .Z(n314) );
  XOR U4068 ( .A(n315), .B(n316), .Z(n304) );
  XOR U4069 ( .A(n302), .B(n317), .Z(n316) );
  XOR U4070 ( .A(n318), .B(n319), .Z(n317) );
  AND U4071 ( .A(b[2]), .B(a[123]), .Z(n318) );
  ANDN U4072 ( .B(n320), .A(n321), .Z(n302) );
  XOR U4073 ( .A(n322), .B(n323), .Z(n315) );
  XNOR U4074 ( .A(n319), .B(n324), .Z(n323) );
  XOR U4075 ( .A(n325), .B(n326), .Z(n324) );
  XOR U4076 ( .A(n327), .B(n328), .Z(n326) );
  XOR U4077 ( .A(n329), .B(n330), .Z(n328) );
  XOR U4078 ( .A(n331), .B(n332), .Z(n330) );
  XOR U4079 ( .A(n288), .B(n333), .Z(n332) );
  XNOR U4080 ( .A(n334), .B(n289), .Z(n333) );
  XOR U4081 ( .A(n335), .B(n336), .Z(n289) );
  XOR U4082 ( .A(n287), .B(n337), .Z(n336) );
  XOR U4083 ( .A(n338), .B(n339), .Z(n337) );
  XOR U4084 ( .A(n340), .B(n341), .Z(n339) );
  XOR U4085 ( .A(n342), .B(n343), .Z(n341) );
  XOR U4086 ( .A(n344), .B(n345), .Z(n343) );
  XOR U4087 ( .A(n346), .B(n347), .Z(n345) );
  XOR U4088 ( .A(n348), .B(n349), .Z(n347) );
  XOR U4089 ( .A(n350), .B(n351), .Z(n349) );
  XOR U4090 ( .A(n352), .B(n353), .Z(n351) );
  XOR U4091 ( .A(n277), .B(n354), .Z(n353) );
  XOR U4092 ( .A(n355), .B(n278), .Z(n354) );
  XOR U4093 ( .A(n356), .B(n357), .Z(n278) );
  XOR U4094 ( .A(n276), .B(n358), .Z(n357) );
  XOR U4095 ( .A(n359), .B(n360), .Z(n358) );
  XOR U4096 ( .A(n361), .B(n362), .Z(n360) );
  XOR U4097 ( .A(n363), .B(n364), .Z(n362) );
  XOR U4098 ( .A(n365), .B(n366), .Z(n364) );
  XOR U4099 ( .A(n367), .B(n368), .Z(n366) );
  XOR U4100 ( .A(n369), .B(n370), .Z(n368) );
  XOR U4101 ( .A(n371), .B(n372), .Z(n370) );
  XOR U4102 ( .A(n373), .B(n374), .Z(n372) );
  XOR U4103 ( .A(n266), .B(n375), .Z(n374) );
  XOR U4104 ( .A(n376), .B(n267), .Z(n375) );
  XOR U4105 ( .A(n377), .B(n378), .Z(n267) );
  XOR U4106 ( .A(n265), .B(n379), .Z(n378) );
  XOR U4107 ( .A(n380), .B(n381), .Z(n379) );
  XOR U4108 ( .A(n382), .B(n383), .Z(n381) );
  XOR U4109 ( .A(n384), .B(n385), .Z(n383) );
  XOR U4110 ( .A(n386), .B(n387), .Z(n385) );
  XOR U4111 ( .A(n388), .B(n389), .Z(n387) );
  XOR U4112 ( .A(n390), .B(n391), .Z(n389) );
  XOR U4113 ( .A(n263), .B(n392), .Z(n391) );
  XNOR U4114 ( .A(n393), .B(n262), .Z(n392) );
  XOR U4115 ( .A(n261), .B(n251), .Z(n394) );
  XOR U4116 ( .A(n395), .B(n396), .Z(n251) );
  XOR U4117 ( .A(n249), .B(n397), .Z(n396) );
  XOR U4118 ( .A(n398), .B(n399), .Z(n397) );
  XOR U4119 ( .A(n400), .B(n401), .Z(n399) );
  XOR U4120 ( .A(n402), .B(n403), .Z(n401) );
  XOR U4121 ( .A(n404), .B(n405), .Z(n403) );
  XOR U4122 ( .A(n406), .B(n407), .Z(n405) );
  XOR U4123 ( .A(n408), .B(n409), .Z(n407) );
  XOR U4124 ( .A(n410), .B(n411), .Z(n409) );
  XOR U4125 ( .A(n412), .B(n413), .Z(n411) );
  XOR U4126 ( .A(n414), .B(n415), .Z(n413) );
  XOR U4127 ( .A(n416), .B(n417), .Z(n415) );
  NAND U4128 ( .A(b[30]), .B(a[95]), .Z(n417) );
  AND U4129 ( .A(a[94]), .B(b[31]), .Z(n416) );
  XOR U4130 ( .A(n418), .B(n414), .Z(n410) );
  XOR U4131 ( .A(n419), .B(n420), .Z(n414) );
  ANDN U4132 ( .B(n421), .A(n422), .Z(n419) );
  AND U4133 ( .A(b[29]), .B(a[96]), .Z(n418) );
  XOR U4134 ( .A(n423), .B(n412), .Z(n406) );
  XOR U4135 ( .A(n424), .B(n425), .Z(n412) );
  AND U4136 ( .A(n426), .B(n427), .Z(n424) );
  AND U4137 ( .A(b[28]), .B(a[97]), .Z(n423) );
  XOR U4138 ( .A(n428), .B(n408), .Z(n402) );
  XOR U4139 ( .A(n429), .B(n430), .Z(n408) );
  AND U4140 ( .A(n431), .B(n432), .Z(n429) );
  AND U4141 ( .A(b[27]), .B(a[98]), .Z(n428) );
  XOR U4142 ( .A(n433), .B(n404), .Z(n398) );
  XOR U4143 ( .A(n434), .B(n435), .Z(n404) );
  AND U4144 ( .A(n436), .B(n437), .Z(n434) );
  AND U4145 ( .A(b[26]), .B(a[99]), .Z(n433) );
  XOR U4146 ( .A(n438), .B(n400), .Z(n395) );
  XOR U4147 ( .A(n439), .B(n440), .Z(n400) );
  AND U4148 ( .A(n441), .B(n442), .Z(n439) );
  AND U4149 ( .A(b[25]), .B(a[100]), .Z(n438) );
  XOR U4150 ( .A(n443), .B(n249), .Z(n250) );
  XOR U4151 ( .A(n444), .B(n445), .Z(n249) );
  AND U4152 ( .A(n446), .B(n447), .Z(n444) );
  AND U4153 ( .A(b[24]), .B(a[101]), .Z(n443) );
  XOR U4154 ( .A(n448), .B(n261), .Z(n263) );
  XOR U4155 ( .A(n449), .B(n450), .Z(n261) );
  AND U4156 ( .A(n451), .B(n452), .Z(n449) );
  AND U4157 ( .A(b[23]), .B(a[102]), .Z(n448) );
  XOR U4158 ( .A(n453), .B(n393), .Z(n388) );
  XOR U4159 ( .A(n454), .B(n455), .Z(n393) );
  AND U4160 ( .A(n456), .B(n457), .Z(n454) );
  AND U4161 ( .A(b[22]), .B(a[103]), .Z(n453) );
  XOR U4162 ( .A(n458), .B(n390), .Z(n384) );
  XOR U4163 ( .A(n459), .B(n460), .Z(n390) );
  AND U4164 ( .A(n461), .B(n462), .Z(n459) );
  AND U4165 ( .A(b[21]), .B(a[104]), .Z(n458) );
  XOR U4166 ( .A(n463), .B(n386), .Z(n380) );
  XOR U4167 ( .A(n464), .B(n465), .Z(n386) );
  AND U4168 ( .A(n466), .B(n467), .Z(n464) );
  AND U4169 ( .A(b[20]), .B(a[105]), .Z(n463) );
  XOR U4170 ( .A(n468), .B(n382), .Z(n377) );
  XOR U4171 ( .A(n469), .B(n470), .Z(n382) );
  AND U4172 ( .A(n471), .B(n472), .Z(n469) );
  AND U4173 ( .A(b[19]), .B(a[106]), .Z(n468) );
  XOR U4174 ( .A(n473), .B(n265), .Z(n266) );
  XOR U4175 ( .A(n474), .B(n475), .Z(n265) );
  AND U4176 ( .A(n476), .B(n477), .Z(n474) );
  AND U4177 ( .A(b[18]), .B(a[107]), .Z(n473) );
  XOR U4178 ( .A(n478), .B(n376), .Z(n371) );
  XOR U4179 ( .A(n479), .B(n480), .Z(n376) );
  AND U4180 ( .A(n481), .B(n482), .Z(n479) );
  AND U4181 ( .A(b[17]), .B(a[108]), .Z(n478) );
  XOR U4182 ( .A(n483), .B(n373), .Z(n367) );
  XOR U4183 ( .A(n484), .B(n485), .Z(n373) );
  AND U4184 ( .A(n486), .B(n487), .Z(n484) );
  AND U4185 ( .A(b[16]), .B(a[109]), .Z(n483) );
  XOR U4186 ( .A(n488), .B(n369), .Z(n363) );
  XOR U4187 ( .A(n489), .B(n490), .Z(n369) );
  AND U4188 ( .A(n491), .B(n492), .Z(n489) );
  AND U4189 ( .A(b[15]), .B(a[110]), .Z(n488) );
  XOR U4190 ( .A(n493), .B(n365), .Z(n359) );
  XOR U4191 ( .A(n494), .B(n495), .Z(n365) );
  AND U4192 ( .A(n496), .B(n497), .Z(n494) );
  AND U4193 ( .A(b[14]), .B(a[111]), .Z(n493) );
  XOR U4194 ( .A(n498), .B(n361), .Z(n356) );
  XOR U4195 ( .A(n499), .B(n500), .Z(n361) );
  AND U4196 ( .A(n501), .B(n502), .Z(n499) );
  AND U4197 ( .A(b[13]), .B(a[112]), .Z(n498) );
  XOR U4198 ( .A(n503), .B(n276), .Z(n277) );
  XOR U4199 ( .A(n504), .B(n505), .Z(n276) );
  AND U4200 ( .A(n506), .B(n507), .Z(n504) );
  AND U4201 ( .A(b[12]), .B(a[113]), .Z(n503) );
  XOR U4202 ( .A(n508), .B(n355), .Z(n350) );
  XOR U4203 ( .A(n509), .B(n510), .Z(n355) );
  AND U4204 ( .A(n511), .B(n512), .Z(n509) );
  AND U4205 ( .A(b[11]), .B(a[114]), .Z(n508) );
  XOR U4206 ( .A(n513), .B(n352), .Z(n346) );
  XOR U4207 ( .A(n514), .B(n515), .Z(n352) );
  AND U4208 ( .A(n516), .B(n517), .Z(n514) );
  AND U4209 ( .A(b[10]), .B(a[115]), .Z(n513) );
  XOR U4210 ( .A(n518), .B(n348), .Z(n342) );
  XOR U4211 ( .A(n519), .B(n520), .Z(n348) );
  AND U4212 ( .A(n521), .B(n522), .Z(n519) );
  AND U4213 ( .A(b[9]), .B(a[116]), .Z(n518) );
  XOR U4214 ( .A(n523), .B(n344), .Z(n338) );
  XOR U4215 ( .A(n524), .B(n525), .Z(n344) );
  AND U4216 ( .A(n526), .B(n527), .Z(n524) );
  AND U4217 ( .A(b[8]), .B(a[117]), .Z(n523) );
  XOR U4218 ( .A(n528), .B(n340), .Z(n335) );
  XOR U4219 ( .A(n529), .B(n530), .Z(n340) );
  AND U4220 ( .A(n531), .B(n532), .Z(n529) );
  AND U4221 ( .A(b[7]), .B(a[118]), .Z(n528) );
  XOR U4222 ( .A(n533), .B(n287), .Z(n288) );
  XOR U4223 ( .A(n534), .B(n535), .Z(n287) );
  AND U4224 ( .A(n536), .B(n537), .Z(n534) );
  AND U4225 ( .A(b[6]), .B(a[119]), .Z(n533) );
  XOR U4226 ( .A(n538), .B(n334), .Z(n329) );
  XOR U4227 ( .A(n539), .B(n540), .Z(n334) );
  AND U4228 ( .A(n541), .B(n542), .Z(n539) );
  AND U4229 ( .A(b[5]), .B(a[120]), .Z(n538) );
  XOR U4230 ( .A(n543), .B(n331), .Z(n325) );
  XOR U4231 ( .A(n544), .B(n545), .Z(n331) );
  AND U4232 ( .A(n546), .B(n547), .Z(n544) );
  AND U4233 ( .A(b[4]), .B(a[121]), .Z(n543) );
  XNOR U4234 ( .A(n548), .B(n549), .Z(n319) );
  NANDN U4235 ( .A(n550), .B(n551), .Z(n549) );
  XOR U4236 ( .A(n552), .B(n327), .Z(n322) );
  XNOR U4237 ( .A(n553), .B(n554), .Z(n327) );
  AND U4238 ( .A(n555), .B(n556), .Z(n553) );
  AND U4239 ( .A(b[3]), .B(a[122]), .Z(n552) );
  XNOR U4240 ( .A(n557), .B(n558), .Z(swire[124]) );
  XOR U4241 ( .A(n320), .B(n559), .Z(n558) );
  XOR U4242 ( .A(n321), .B(n557), .Z(n559) );
  NAND U4243 ( .A(a[124]), .B(b[0]), .Z(n321) );
  XNOR U4244 ( .A(n550), .B(n551), .Z(n320) );
  XOR U4245 ( .A(n548), .B(n560), .Z(n551) );
  NAND U4246 ( .A(b[1]), .B(a[123]), .Z(n560) );
  XOR U4247 ( .A(n556), .B(n561), .Z(n550) );
  XOR U4248 ( .A(n548), .B(n555), .Z(n561) );
  XNOR U4249 ( .A(n562), .B(n554), .Z(n555) );
  AND U4250 ( .A(b[2]), .B(a[122]), .Z(n562) );
  NANDN U4251 ( .A(n563), .B(n564), .Z(n548) );
  XOR U4252 ( .A(n554), .B(n546), .Z(n565) );
  XNOR U4253 ( .A(n545), .B(n541), .Z(n566) );
  XNOR U4254 ( .A(n540), .B(n536), .Z(n567) );
  XNOR U4255 ( .A(n535), .B(n531), .Z(n568) );
  XNOR U4256 ( .A(n530), .B(n526), .Z(n569) );
  XNOR U4257 ( .A(n525), .B(n521), .Z(n570) );
  XNOR U4258 ( .A(n520), .B(n516), .Z(n571) );
  XNOR U4259 ( .A(n515), .B(n511), .Z(n572) );
  XNOR U4260 ( .A(n510), .B(n506), .Z(n573) );
  XNOR U4261 ( .A(n505), .B(n501), .Z(n574) );
  XNOR U4262 ( .A(n500), .B(n496), .Z(n575) );
  XNOR U4263 ( .A(n495), .B(n491), .Z(n576) );
  XNOR U4264 ( .A(n490), .B(n486), .Z(n577) );
  XNOR U4265 ( .A(n485), .B(n481), .Z(n578) );
  XNOR U4266 ( .A(n480), .B(n476), .Z(n579) );
  XNOR U4267 ( .A(n475), .B(n471), .Z(n580) );
  XNOR U4268 ( .A(n470), .B(n466), .Z(n581) );
  XNOR U4269 ( .A(n465), .B(n461), .Z(n582) );
  XNOR U4270 ( .A(n460), .B(n456), .Z(n583) );
  XNOR U4271 ( .A(n455), .B(n451), .Z(n584) );
  XNOR U4272 ( .A(n450), .B(n446), .Z(n585) );
  XNOR U4273 ( .A(n445), .B(n441), .Z(n586) );
  XNOR U4274 ( .A(n440), .B(n436), .Z(n587) );
  XNOR U4275 ( .A(n435), .B(n431), .Z(n588) );
  XNOR U4276 ( .A(n430), .B(n426), .Z(n589) );
  XOR U4277 ( .A(n425), .B(n422), .Z(n590) );
  XOR U4278 ( .A(n591), .B(n592), .Z(n422) );
  XOR U4279 ( .A(n420), .B(n593), .Z(n592) );
  XOR U4280 ( .A(n594), .B(n595), .Z(n593) );
  XOR U4281 ( .A(n596), .B(n597), .Z(n595) );
  NAND U4282 ( .A(a[94]), .B(b[30]), .Z(n597) );
  AND U4283 ( .A(a[93]), .B(b[31]), .Z(n596) );
  XOR U4284 ( .A(n598), .B(n594), .Z(n591) );
  XOR U4285 ( .A(n599), .B(n600), .Z(n594) );
  ANDN U4286 ( .B(n601), .A(n602), .Z(n599) );
  AND U4287 ( .A(b[29]), .B(a[95]), .Z(n598) );
  XOR U4288 ( .A(n603), .B(n420), .Z(n421) );
  XOR U4289 ( .A(n604), .B(n605), .Z(n420) );
  AND U4290 ( .A(n606), .B(n607), .Z(n604) );
  AND U4291 ( .A(b[28]), .B(a[96]), .Z(n603) );
  XOR U4292 ( .A(n608), .B(n425), .Z(n427) );
  XOR U4293 ( .A(n609), .B(n610), .Z(n425) );
  AND U4294 ( .A(n611), .B(n612), .Z(n609) );
  AND U4295 ( .A(b[27]), .B(a[97]), .Z(n608) );
  XOR U4296 ( .A(n613), .B(n430), .Z(n432) );
  XOR U4297 ( .A(n614), .B(n615), .Z(n430) );
  AND U4298 ( .A(n616), .B(n617), .Z(n614) );
  AND U4299 ( .A(b[26]), .B(a[98]), .Z(n613) );
  XOR U4300 ( .A(n618), .B(n435), .Z(n437) );
  XOR U4301 ( .A(n619), .B(n620), .Z(n435) );
  AND U4302 ( .A(n621), .B(n622), .Z(n619) );
  AND U4303 ( .A(b[25]), .B(a[99]), .Z(n618) );
  XOR U4304 ( .A(n623), .B(n440), .Z(n442) );
  XOR U4305 ( .A(n624), .B(n625), .Z(n440) );
  AND U4306 ( .A(n626), .B(n627), .Z(n624) );
  AND U4307 ( .A(b[24]), .B(a[100]), .Z(n623) );
  XOR U4308 ( .A(n628), .B(n445), .Z(n447) );
  XOR U4309 ( .A(n629), .B(n630), .Z(n445) );
  AND U4310 ( .A(n631), .B(n632), .Z(n629) );
  AND U4311 ( .A(b[23]), .B(a[101]), .Z(n628) );
  XOR U4312 ( .A(n633), .B(n450), .Z(n452) );
  XOR U4313 ( .A(n634), .B(n635), .Z(n450) );
  AND U4314 ( .A(n636), .B(n637), .Z(n634) );
  AND U4315 ( .A(b[22]), .B(a[102]), .Z(n633) );
  XOR U4316 ( .A(n638), .B(n455), .Z(n457) );
  XOR U4317 ( .A(n639), .B(n640), .Z(n455) );
  AND U4318 ( .A(n641), .B(n642), .Z(n639) );
  AND U4319 ( .A(b[21]), .B(a[103]), .Z(n638) );
  XOR U4320 ( .A(n643), .B(n460), .Z(n462) );
  XOR U4321 ( .A(n644), .B(n645), .Z(n460) );
  AND U4322 ( .A(n646), .B(n647), .Z(n644) );
  AND U4323 ( .A(b[20]), .B(a[104]), .Z(n643) );
  XOR U4324 ( .A(n648), .B(n465), .Z(n467) );
  XOR U4325 ( .A(n649), .B(n650), .Z(n465) );
  AND U4326 ( .A(n651), .B(n652), .Z(n649) );
  AND U4327 ( .A(b[19]), .B(a[105]), .Z(n648) );
  XOR U4328 ( .A(n653), .B(n470), .Z(n472) );
  XOR U4329 ( .A(n654), .B(n655), .Z(n470) );
  AND U4330 ( .A(n656), .B(n657), .Z(n654) );
  AND U4331 ( .A(b[18]), .B(a[106]), .Z(n653) );
  XOR U4332 ( .A(n658), .B(n475), .Z(n477) );
  XOR U4333 ( .A(n659), .B(n660), .Z(n475) );
  AND U4334 ( .A(n661), .B(n662), .Z(n659) );
  AND U4335 ( .A(b[17]), .B(a[107]), .Z(n658) );
  XOR U4336 ( .A(n663), .B(n480), .Z(n482) );
  XOR U4337 ( .A(n664), .B(n665), .Z(n480) );
  AND U4338 ( .A(n666), .B(n667), .Z(n664) );
  AND U4339 ( .A(b[16]), .B(a[108]), .Z(n663) );
  XOR U4340 ( .A(n668), .B(n485), .Z(n487) );
  XOR U4341 ( .A(n669), .B(n670), .Z(n485) );
  AND U4342 ( .A(n671), .B(n672), .Z(n669) );
  AND U4343 ( .A(b[15]), .B(a[109]), .Z(n668) );
  XOR U4344 ( .A(n673), .B(n490), .Z(n492) );
  XOR U4345 ( .A(n674), .B(n675), .Z(n490) );
  AND U4346 ( .A(n676), .B(n677), .Z(n674) );
  AND U4347 ( .A(b[14]), .B(a[110]), .Z(n673) );
  XOR U4348 ( .A(n678), .B(n495), .Z(n497) );
  XOR U4349 ( .A(n679), .B(n680), .Z(n495) );
  AND U4350 ( .A(n681), .B(n682), .Z(n679) );
  AND U4351 ( .A(b[13]), .B(a[111]), .Z(n678) );
  XOR U4352 ( .A(n683), .B(n500), .Z(n502) );
  XOR U4353 ( .A(n684), .B(n685), .Z(n500) );
  AND U4354 ( .A(n686), .B(n687), .Z(n684) );
  AND U4355 ( .A(b[12]), .B(a[112]), .Z(n683) );
  XOR U4356 ( .A(n688), .B(n505), .Z(n507) );
  XOR U4357 ( .A(n689), .B(n690), .Z(n505) );
  AND U4358 ( .A(n691), .B(n692), .Z(n689) );
  AND U4359 ( .A(b[11]), .B(a[113]), .Z(n688) );
  XOR U4360 ( .A(n693), .B(n510), .Z(n512) );
  XOR U4361 ( .A(n694), .B(n695), .Z(n510) );
  AND U4362 ( .A(n696), .B(n697), .Z(n694) );
  AND U4363 ( .A(b[10]), .B(a[114]), .Z(n693) );
  XOR U4364 ( .A(n698), .B(n515), .Z(n517) );
  XOR U4365 ( .A(n699), .B(n700), .Z(n515) );
  AND U4366 ( .A(n701), .B(n702), .Z(n699) );
  AND U4367 ( .A(b[9]), .B(a[115]), .Z(n698) );
  XOR U4368 ( .A(n703), .B(n520), .Z(n522) );
  XOR U4369 ( .A(n704), .B(n705), .Z(n520) );
  AND U4370 ( .A(n706), .B(n707), .Z(n704) );
  AND U4371 ( .A(b[8]), .B(a[116]), .Z(n703) );
  XOR U4372 ( .A(n708), .B(n525), .Z(n527) );
  XOR U4373 ( .A(n709), .B(n710), .Z(n525) );
  AND U4374 ( .A(n711), .B(n712), .Z(n709) );
  AND U4375 ( .A(b[7]), .B(a[117]), .Z(n708) );
  XOR U4376 ( .A(n713), .B(n530), .Z(n532) );
  XOR U4377 ( .A(n714), .B(n715), .Z(n530) );
  AND U4378 ( .A(n716), .B(n717), .Z(n714) );
  AND U4379 ( .A(b[6]), .B(a[118]), .Z(n713) );
  XOR U4380 ( .A(n718), .B(n535), .Z(n537) );
  XOR U4381 ( .A(n719), .B(n720), .Z(n535) );
  AND U4382 ( .A(n721), .B(n722), .Z(n719) );
  AND U4383 ( .A(b[5]), .B(a[119]), .Z(n718) );
  XOR U4384 ( .A(n723), .B(n540), .Z(n542) );
  XOR U4385 ( .A(n724), .B(n725), .Z(n540) );
  AND U4386 ( .A(n726), .B(n727), .Z(n724) );
  AND U4387 ( .A(b[4]), .B(a[120]), .Z(n723) );
  XNOR U4388 ( .A(n728), .B(n729), .Z(n554) );
  NANDN U4389 ( .A(n730), .B(n731), .Z(n729) );
  XOR U4390 ( .A(n732), .B(n545), .Z(n547) );
  XNOR U4391 ( .A(n733), .B(n734), .Z(n545) );
  AND U4392 ( .A(n735), .B(n736), .Z(n733) );
  AND U4393 ( .A(b[3]), .B(a[121]), .Z(n732) );
  XOR U4394 ( .A(n737), .B(n738), .Z(swire[123]) );
  XOR U4395 ( .A(n564), .B(n740), .Z(n738) );
  XOR U4396 ( .A(n563), .B(n739), .Z(n740) );
  IV U4397 ( .A(n737), .Z(n739) );
  NAND U4398 ( .A(a[123]), .B(b[0]), .Z(n563) );
  XNOR U4399 ( .A(n730), .B(n731), .Z(n564) );
  XOR U4400 ( .A(n728), .B(n741), .Z(n731) );
  NAND U4401 ( .A(b[1]), .B(a[122]), .Z(n741) );
  XOR U4402 ( .A(n736), .B(n742), .Z(n730) );
  XOR U4403 ( .A(n728), .B(n735), .Z(n742) );
  XNOR U4404 ( .A(n743), .B(n734), .Z(n735) );
  AND U4405 ( .A(b[2]), .B(a[121]), .Z(n743) );
  NANDN U4406 ( .A(n744), .B(n745), .Z(n728) );
  XOR U4407 ( .A(n734), .B(n726), .Z(n746) );
  XNOR U4408 ( .A(n725), .B(n721), .Z(n747) );
  XNOR U4409 ( .A(n720), .B(n716), .Z(n748) );
  XNOR U4410 ( .A(n715), .B(n711), .Z(n749) );
  XNOR U4411 ( .A(n710), .B(n706), .Z(n750) );
  XNOR U4412 ( .A(n705), .B(n701), .Z(n751) );
  XNOR U4413 ( .A(n700), .B(n696), .Z(n752) );
  XNOR U4414 ( .A(n695), .B(n691), .Z(n753) );
  XNOR U4415 ( .A(n690), .B(n686), .Z(n754) );
  XNOR U4416 ( .A(n685), .B(n681), .Z(n755) );
  XNOR U4417 ( .A(n680), .B(n676), .Z(n756) );
  XNOR U4418 ( .A(n675), .B(n671), .Z(n757) );
  XNOR U4419 ( .A(n670), .B(n666), .Z(n758) );
  XNOR U4420 ( .A(n665), .B(n661), .Z(n759) );
  XNOR U4421 ( .A(n660), .B(n656), .Z(n760) );
  XNOR U4422 ( .A(n655), .B(n651), .Z(n761) );
  XNOR U4423 ( .A(n650), .B(n646), .Z(n762) );
  XNOR U4424 ( .A(n645), .B(n641), .Z(n763) );
  XNOR U4425 ( .A(n640), .B(n636), .Z(n764) );
  XNOR U4426 ( .A(n635), .B(n631), .Z(n765) );
  XNOR U4427 ( .A(n630), .B(n626), .Z(n766) );
  XNOR U4428 ( .A(n625), .B(n621), .Z(n767) );
  XNOR U4429 ( .A(n620), .B(n616), .Z(n768) );
  XNOR U4430 ( .A(n615), .B(n611), .Z(n769) );
  XNOR U4431 ( .A(n610), .B(n606), .Z(n770) );
  XOR U4432 ( .A(n605), .B(n602), .Z(n771) );
  XOR U4433 ( .A(n772), .B(n773), .Z(n602) );
  XOR U4434 ( .A(n600), .B(n774), .Z(n773) );
  XOR U4435 ( .A(n775), .B(n776), .Z(n774) );
  XOR U4436 ( .A(n777), .B(n778), .Z(n776) );
  NAND U4437 ( .A(a[93]), .B(b[30]), .Z(n778) );
  AND U4438 ( .A(a[92]), .B(b[31]), .Z(n777) );
  XOR U4439 ( .A(n779), .B(n775), .Z(n772) );
  XOR U4440 ( .A(n780), .B(n781), .Z(n775) );
  ANDN U4441 ( .B(n782), .A(n783), .Z(n780) );
  AND U4442 ( .A(a[94]), .B(b[29]), .Z(n779) );
  XOR U4443 ( .A(n784), .B(n600), .Z(n601) );
  XOR U4444 ( .A(n785), .B(n786), .Z(n600) );
  AND U4445 ( .A(n787), .B(n788), .Z(n785) );
  AND U4446 ( .A(b[28]), .B(a[95]), .Z(n784) );
  XOR U4447 ( .A(n789), .B(n605), .Z(n607) );
  XOR U4448 ( .A(n790), .B(n791), .Z(n605) );
  AND U4449 ( .A(n792), .B(n793), .Z(n790) );
  AND U4450 ( .A(b[27]), .B(a[96]), .Z(n789) );
  XOR U4451 ( .A(n794), .B(n610), .Z(n612) );
  XOR U4452 ( .A(n795), .B(n796), .Z(n610) );
  AND U4453 ( .A(n797), .B(n798), .Z(n795) );
  AND U4454 ( .A(b[26]), .B(a[97]), .Z(n794) );
  XOR U4455 ( .A(n799), .B(n615), .Z(n617) );
  XOR U4456 ( .A(n800), .B(n801), .Z(n615) );
  AND U4457 ( .A(n802), .B(n803), .Z(n800) );
  AND U4458 ( .A(b[25]), .B(a[98]), .Z(n799) );
  XOR U4459 ( .A(n804), .B(n620), .Z(n622) );
  XOR U4460 ( .A(n805), .B(n806), .Z(n620) );
  AND U4461 ( .A(n807), .B(n808), .Z(n805) );
  AND U4462 ( .A(b[24]), .B(a[99]), .Z(n804) );
  XOR U4463 ( .A(n809), .B(n625), .Z(n627) );
  XOR U4464 ( .A(n810), .B(n811), .Z(n625) );
  AND U4465 ( .A(n812), .B(n813), .Z(n810) );
  AND U4466 ( .A(b[23]), .B(a[100]), .Z(n809) );
  XOR U4467 ( .A(n814), .B(n630), .Z(n632) );
  XOR U4468 ( .A(n815), .B(n816), .Z(n630) );
  AND U4469 ( .A(n817), .B(n818), .Z(n815) );
  AND U4470 ( .A(b[22]), .B(a[101]), .Z(n814) );
  XOR U4471 ( .A(n819), .B(n635), .Z(n637) );
  XOR U4472 ( .A(n820), .B(n821), .Z(n635) );
  AND U4473 ( .A(n822), .B(n823), .Z(n820) );
  AND U4474 ( .A(b[21]), .B(a[102]), .Z(n819) );
  XOR U4475 ( .A(n824), .B(n640), .Z(n642) );
  XOR U4476 ( .A(n825), .B(n826), .Z(n640) );
  AND U4477 ( .A(n827), .B(n828), .Z(n825) );
  AND U4478 ( .A(b[20]), .B(a[103]), .Z(n824) );
  XOR U4479 ( .A(n829), .B(n645), .Z(n647) );
  XOR U4480 ( .A(n830), .B(n831), .Z(n645) );
  AND U4481 ( .A(n832), .B(n833), .Z(n830) );
  AND U4482 ( .A(b[19]), .B(a[104]), .Z(n829) );
  XOR U4483 ( .A(n834), .B(n650), .Z(n652) );
  XOR U4484 ( .A(n835), .B(n836), .Z(n650) );
  AND U4485 ( .A(n837), .B(n838), .Z(n835) );
  AND U4486 ( .A(b[18]), .B(a[105]), .Z(n834) );
  XOR U4487 ( .A(n839), .B(n655), .Z(n657) );
  XOR U4488 ( .A(n840), .B(n841), .Z(n655) );
  AND U4489 ( .A(n842), .B(n843), .Z(n840) );
  AND U4490 ( .A(b[17]), .B(a[106]), .Z(n839) );
  XOR U4491 ( .A(n844), .B(n660), .Z(n662) );
  XOR U4492 ( .A(n845), .B(n846), .Z(n660) );
  AND U4493 ( .A(n847), .B(n848), .Z(n845) );
  AND U4494 ( .A(b[16]), .B(a[107]), .Z(n844) );
  XOR U4495 ( .A(n849), .B(n665), .Z(n667) );
  XOR U4496 ( .A(n850), .B(n851), .Z(n665) );
  AND U4497 ( .A(n852), .B(n853), .Z(n850) );
  AND U4498 ( .A(b[15]), .B(a[108]), .Z(n849) );
  XOR U4499 ( .A(n854), .B(n670), .Z(n672) );
  XOR U4500 ( .A(n855), .B(n856), .Z(n670) );
  AND U4501 ( .A(n857), .B(n858), .Z(n855) );
  AND U4502 ( .A(b[14]), .B(a[109]), .Z(n854) );
  XOR U4503 ( .A(n859), .B(n675), .Z(n677) );
  XOR U4504 ( .A(n860), .B(n861), .Z(n675) );
  AND U4505 ( .A(n862), .B(n863), .Z(n860) );
  AND U4506 ( .A(b[13]), .B(a[110]), .Z(n859) );
  XOR U4507 ( .A(n864), .B(n680), .Z(n682) );
  XOR U4508 ( .A(n865), .B(n866), .Z(n680) );
  AND U4509 ( .A(n867), .B(n868), .Z(n865) );
  AND U4510 ( .A(b[12]), .B(a[111]), .Z(n864) );
  XOR U4511 ( .A(n869), .B(n685), .Z(n687) );
  XOR U4512 ( .A(n870), .B(n871), .Z(n685) );
  AND U4513 ( .A(n872), .B(n873), .Z(n870) );
  AND U4514 ( .A(b[11]), .B(a[112]), .Z(n869) );
  XOR U4515 ( .A(n874), .B(n690), .Z(n692) );
  XOR U4516 ( .A(n875), .B(n876), .Z(n690) );
  AND U4517 ( .A(n877), .B(n878), .Z(n875) );
  AND U4518 ( .A(b[10]), .B(a[113]), .Z(n874) );
  XOR U4519 ( .A(n879), .B(n695), .Z(n697) );
  XOR U4520 ( .A(n880), .B(n881), .Z(n695) );
  AND U4521 ( .A(n882), .B(n883), .Z(n880) );
  AND U4522 ( .A(b[9]), .B(a[114]), .Z(n879) );
  XOR U4523 ( .A(n884), .B(n700), .Z(n702) );
  XOR U4524 ( .A(n885), .B(n886), .Z(n700) );
  AND U4525 ( .A(n887), .B(n888), .Z(n885) );
  AND U4526 ( .A(b[8]), .B(a[115]), .Z(n884) );
  XOR U4527 ( .A(n889), .B(n705), .Z(n707) );
  XOR U4528 ( .A(n890), .B(n891), .Z(n705) );
  AND U4529 ( .A(n892), .B(n893), .Z(n890) );
  AND U4530 ( .A(b[7]), .B(a[116]), .Z(n889) );
  XOR U4531 ( .A(n894), .B(n710), .Z(n712) );
  XOR U4532 ( .A(n895), .B(n896), .Z(n710) );
  AND U4533 ( .A(n897), .B(n898), .Z(n895) );
  AND U4534 ( .A(b[6]), .B(a[117]), .Z(n894) );
  XOR U4535 ( .A(n899), .B(n715), .Z(n717) );
  XOR U4536 ( .A(n900), .B(n901), .Z(n715) );
  AND U4537 ( .A(n902), .B(n903), .Z(n900) );
  AND U4538 ( .A(b[5]), .B(a[118]), .Z(n899) );
  XOR U4539 ( .A(n904), .B(n720), .Z(n722) );
  XOR U4540 ( .A(n905), .B(n906), .Z(n720) );
  AND U4541 ( .A(n907), .B(n908), .Z(n905) );
  AND U4542 ( .A(b[4]), .B(a[119]), .Z(n904) );
  XNOR U4543 ( .A(n909), .B(n910), .Z(n734) );
  NANDN U4544 ( .A(n911), .B(n912), .Z(n910) );
  XOR U4545 ( .A(n913), .B(n725), .Z(n727) );
  XNOR U4546 ( .A(n914), .B(n915), .Z(n725) );
  AND U4547 ( .A(n916), .B(n917), .Z(n914) );
  AND U4548 ( .A(b[3]), .B(a[120]), .Z(n913) );
  XNOR U4549 ( .A(n918), .B(n919), .Z(swire[122]) );
  XOR U4550 ( .A(n745), .B(n920), .Z(n919) );
  XOR U4551 ( .A(n744), .B(n918), .Z(n920) );
  NAND U4552 ( .A(a[122]), .B(b[0]), .Z(n744) );
  XNOR U4553 ( .A(n911), .B(n912), .Z(n745) );
  XOR U4554 ( .A(n909), .B(n921), .Z(n912) );
  NAND U4555 ( .A(b[1]), .B(a[121]), .Z(n921) );
  XOR U4556 ( .A(n917), .B(n922), .Z(n911) );
  XOR U4557 ( .A(n909), .B(n916), .Z(n922) );
  XNOR U4558 ( .A(n923), .B(n915), .Z(n916) );
  AND U4559 ( .A(b[2]), .B(a[120]), .Z(n923) );
  NANDN U4560 ( .A(n924), .B(n925), .Z(n909) );
  XOR U4561 ( .A(n915), .B(n907), .Z(n926) );
  XNOR U4562 ( .A(n906), .B(n902), .Z(n927) );
  XNOR U4563 ( .A(n901), .B(n897), .Z(n928) );
  XNOR U4564 ( .A(n896), .B(n892), .Z(n929) );
  XNOR U4565 ( .A(n891), .B(n887), .Z(n930) );
  XNOR U4566 ( .A(n886), .B(n882), .Z(n931) );
  XNOR U4567 ( .A(n881), .B(n877), .Z(n932) );
  XNOR U4568 ( .A(n876), .B(n872), .Z(n933) );
  XNOR U4569 ( .A(n871), .B(n867), .Z(n934) );
  XNOR U4570 ( .A(n866), .B(n862), .Z(n935) );
  XNOR U4571 ( .A(n861), .B(n857), .Z(n936) );
  XNOR U4572 ( .A(n856), .B(n852), .Z(n937) );
  XNOR U4573 ( .A(n851), .B(n847), .Z(n938) );
  XNOR U4574 ( .A(n846), .B(n842), .Z(n939) );
  XNOR U4575 ( .A(n841), .B(n837), .Z(n940) );
  XNOR U4576 ( .A(n836), .B(n832), .Z(n941) );
  XNOR U4577 ( .A(n831), .B(n827), .Z(n942) );
  XNOR U4578 ( .A(n826), .B(n822), .Z(n943) );
  XNOR U4579 ( .A(n821), .B(n817), .Z(n944) );
  XNOR U4580 ( .A(n816), .B(n812), .Z(n945) );
  XNOR U4581 ( .A(n811), .B(n807), .Z(n946) );
  XNOR U4582 ( .A(n806), .B(n802), .Z(n947) );
  XNOR U4583 ( .A(n801), .B(n797), .Z(n948) );
  XNOR U4584 ( .A(n796), .B(n792), .Z(n949) );
  XNOR U4585 ( .A(n791), .B(n787), .Z(n950) );
  XOR U4586 ( .A(n786), .B(n783), .Z(n951) );
  XOR U4587 ( .A(n952), .B(n953), .Z(n783) );
  XOR U4588 ( .A(n781), .B(n954), .Z(n953) );
  XOR U4589 ( .A(n955), .B(n956), .Z(n954) );
  XOR U4590 ( .A(n957), .B(n958), .Z(n956) );
  NAND U4591 ( .A(a[92]), .B(b[30]), .Z(n958) );
  AND U4592 ( .A(a[91]), .B(b[31]), .Z(n957) );
  XOR U4593 ( .A(n959), .B(n955), .Z(n952) );
  XOR U4594 ( .A(n960), .B(n961), .Z(n955) );
  ANDN U4595 ( .B(n962), .A(n963), .Z(n960) );
  AND U4596 ( .A(a[93]), .B(b[29]), .Z(n959) );
  XOR U4597 ( .A(n964), .B(n781), .Z(n782) );
  XOR U4598 ( .A(n965), .B(n966), .Z(n781) );
  AND U4599 ( .A(n967), .B(n968), .Z(n965) );
  AND U4600 ( .A(a[94]), .B(b[28]), .Z(n964) );
  XOR U4601 ( .A(n969), .B(n786), .Z(n788) );
  XOR U4602 ( .A(n970), .B(n971), .Z(n786) );
  AND U4603 ( .A(n972), .B(n973), .Z(n970) );
  AND U4604 ( .A(b[27]), .B(a[95]), .Z(n969) );
  XOR U4605 ( .A(n974), .B(n791), .Z(n793) );
  XOR U4606 ( .A(n975), .B(n976), .Z(n791) );
  AND U4607 ( .A(n977), .B(n978), .Z(n975) );
  AND U4608 ( .A(b[26]), .B(a[96]), .Z(n974) );
  XOR U4609 ( .A(n979), .B(n796), .Z(n798) );
  XOR U4610 ( .A(n980), .B(n981), .Z(n796) );
  AND U4611 ( .A(n982), .B(n983), .Z(n980) );
  AND U4612 ( .A(b[25]), .B(a[97]), .Z(n979) );
  XOR U4613 ( .A(n984), .B(n801), .Z(n803) );
  XOR U4614 ( .A(n985), .B(n986), .Z(n801) );
  AND U4615 ( .A(n987), .B(n988), .Z(n985) );
  AND U4616 ( .A(b[24]), .B(a[98]), .Z(n984) );
  XOR U4617 ( .A(n989), .B(n806), .Z(n808) );
  XOR U4618 ( .A(n990), .B(n991), .Z(n806) );
  AND U4619 ( .A(n992), .B(n993), .Z(n990) );
  AND U4620 ( .A(b[23]), .B(a[99]), .Z(n989) );
  XOR U4621 ( .A(n994), .B(n811), .Z(n813) );
  XOR U4622 ( .A(n995), .B(n996), .Z(n811) );
  AND U4623 ( .A(n997), .B(n998), .Z(n995) );
  AND U4624 ( .A(b[22]), .B(a[100]), .Z(n994) );
  XOR U4625 ( .A(n999), .B(n816), .Z(n818) );
  XOR U4626 ( .A(n1000), .B(n1001), .Z(n816) );
  AND U4627 ( .A(n1002), .B(n1003), .Z(n1000) );
  AND U4628 ( .A(b[21]), .B(a[101]), .Z(n999) );
  XOR U4629 ( .A(n1004), .B(n821), .Z(n823) );
  XOR U4630 ( .A(n1005), .B(n1006), .Z(n821) );
  AND U4631 ( .A(n1007), .B(n1008), .Z(n1005) );
  AND U4632 ( .A(b[20]), .B(a[102]), .Z(n1004) );
  XOR U4633 ( .A(n1009), .B(n826), .Z(n828) );
  XOR U4634 ( .A(n1010), .B(n1011), .Z(n826) );
  AND U4635 ( .A(n1012), .B(n1013), .Z(n1010) );
  AND U4636 ( .A(b[19]), .B(a[103]), .Z(n1009) );
  XOR U4637 ( .A(n1014), .B(n831), .Z(n833) );
  XOR U4638 ( .A(n1015), .B(n1016), .Z(n831) );
  AND U4639 ( .A(n1017), .B(n1018), .Z(n1015) );
  AND U4640 ( .A(b[18]), .B(a[104]), .Z(n1014) );
  XOR U4641 ( .A(n1019), .B(n836), .Z(n838) );
  XOR U4642 ( .A(n1020), .B(n1021), .Z(n836) );
  AND U4643 ( .A(n1022), .B(n1023), .Z(n1020) );
  AND U4644 ( .A(b[17]), .B(a[105]), .Z(n1019) );
  XOR U4645 ( .A(n1024), .B(n841), .Z(n843) );
  XOR U4646 ( .A(n1025), .B(n1026), .Z(n841) );
  AND U4647 ( .A(n1027), .B(n1028), .Z(n1025) );
  AND U4648 ( .A(b[16]), .B(a[106]), .Z(n1024) );
  XOR U4649 ( .A(n1029), .B(n846), .Z(n848) );
  XOR U4650 ( .A(n1030), .B(n1031), .Z(n846) );
  AND U4651 ( .A(n1032), .B(n1033), .Z(n1030) );
  AND U4652 ( .A(b[15]), .B(a[107]), .Z(n1029) );
  XOR U4653 ( .A(n1034), .B(n851), .Z(n853) );
  XOR U4654 ( .A(n1035), .B(n1036), .Z(n851) );
  AND U4655 ( .A(n1037), .B(n1038), .Z(n1035) );
  AND U4656 ( .A(b[14]), .B(a[108]), .Z(n1034) );
  XOR U4657 ( .A(n1039), .B(n856), .Z(n858) );
  XOR U4658 ( .A(n1040), .B(n1041), .Z(n856) );
  AND U4659 ( .A(n1042), .B(n1043), .Z(n1040) );
  AND U4660 ( .A(b[13]), .B(a[109]), .Z(n1039) );
  XOR U4661 ( .A(n1044), .B(n861), .Z(n863) );
  XOR U4662 ( .A(n1045), .B(n1046), .Z(n861) );
  AND U4663 ( .A(n1047), .B(n1048), .Z(n1045) );
  AND U4664 ( .A(b[12]), .B(a[110]), .Z(n1044) );
  XOR U4665 ( .A(n1049), .B(n866), .Z(n868) );
  XOR U4666 ( .A(n1050), .B(n1051), .Z(n866) );
  AND U4667 ( .A(n1052), .B(n1053), .Z(n1050) );
  AND U4668 ( .A(b[11]), .B(a[111]), .Z(n1049) );
  XOR U4669 ( .A(n1054), .B(n871), .Z(n873) );
  XOR U4670 ( .A(n1055), .B(n1056), .Z(n871) );
  AND U4671 ( .A(n1057), .B(n1058), .Z(n1055) );
  AND U4672 ( .A(b[10]), .B(a[112]), .Z(n1054) );
  XOR U4673 ( .A(n1059), .B(n876), .Z(n878) );
  XOR U4674 ( .A(n1060), .B(n1061), .Z(n876) );
  AND U4675 ( .A(n1062), .B(n1063), .Z(n1060) );
  AND U4676 ( .A(b[9]), .B(a[113]), .Z(n1059) );
  XOR U4677 ( .A(n1064), .B(n881), .Z(n883) );
  XOR U4678 ( .A(n1065), .B(n1066), .Z(n881) );
  AND U4679 ( .A(n1067), .B(n1068), .Z(n1065) );
  AND U4680 ( .A(b[8]), .B(a[114]), .Z(n1064) );
  XOR U4681 ( .A(n1069), .B(n886), .Z(n888) );
  XOR U4682 ( .A(n1070), .B(n1071), .Z(n886) );
  AND U4683 ( .A(n1072), .B(n1073), .Z(n1070) );
  AND U4684 ( .A(b[7]), .B(a[115]), .Z(n1069) );
  XOR U4685 ( .A(n1074), .B(n891), .Z(n893) );
  XOR U4686 ( .A(n1075), .B(n1076), .Z(n891) );
  AND U4687 ( .A(n1077), .B(n1078), .Z(n1075) );
  AND U4688 ( .A(b[6]), .B(a[116]), .Z(n1074) );
  XOR U4689 ( .A(n1079), .B(n896), .Z(n898) );
  XOR U4690 ( .A(n1080), .B(n1081), .Z(n896) );
  AND U4691 ( .A(n1082), .B(n1083), .Z(n1080) );
  AND U4692 ( .A(b[5]), .B(a[117]), .Z(n1079) );
  XOR U4693 ( .A(n1084), .B(n901), .Z(n903) );
  XOR U4694 ( .A(n1085), .B(n1086), .Z(n901) );
  AND U4695 ( .A(n1087), .B(n1088), .Z(n1085) );
  AND U4696 ( .A(b[4]), .B(a[118]), .Z(n1084) );
  XNOR U4697 ( .A(n1089), .B(n1090), .Z(n915) );
  NANDN U4698 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U4699 ( .A(n1093), .B(n906), .Z(n908) );
  XNOR U4700 ( .A(n1094), .B(n1095), .Z(n906) );
  AND U4701 ( .A(n1096), .B(n1097), .Z(n1094) );
  AND U4702 ( .A(b[3]), .B(a[119]), .Z(n1093) );
  XOR U4703 ( .A(n1098), .B(n1099), .Z(swire[121]) );
  XOR U4704 ( .A(n925), .B(n1101), .Z(n1099) );
  XOR U4705 ( .A(n924), .B(n1100), .Z(n1101) );
  IV U4706 ( .A(n1098), .Z(n1100) );
  NAND U4707 ( .A(a[121]), .B(b[0]), .Z(n924) );
  XNOR U4708 ( .A(n1091), .B(n1092), .Z(n925) );
  XOR U4709 ( .A(n1089), .B(n1102), .Z(n1092) );
  NAND U4710 ( .A(b[1]), .B(a[120]), .Z(n1102) );
  XOR U4711 ( .A(n1097), .B(n1103), .Z(n1091) );
  XOR U4712 ( .A(n1089), .B(n1096), .Z(n1103) );
  XNOR U4713 ( .A(n1104), .B(n1095), .Z(n1096) );
  AND U4714 ( .A(b[2]), .B(a[119]), .Z(n1104) );
  NANDN U4715 ( .A(n1105), .B(n1106), .Z(n1089) );
  XOR U4716 ( .A(n1095), .B(n1087), .Z(n1107) );
  XNOR U4717 ( .A(n1086), .B(n1082), .Z(n1108) );
  XNOR U4718 ( .A(n1081), .B(n1077), .Z(n1109) );
  XNOR U4719 ( .A(n1076), .B(n1072), .Z(n1110) );
  XNOR U4720 ( .A(n1071), .B(n1067), .Z(n1111) );
  XNOR U4721 ( .A(n1066), .B(n1062), .Z(n1112) );
  XNOR U4722 ( .A(n1061), .B(n1057), .Z(n1113) );
  XNOR U4723 ( .A(n1056), .B(n1052), .Z(n1114) );
  XNOR U4724 ( .A(n1051), .B(n1047), .Z(n1115) );
  XNOR U4725 ( .A(n1046), .B(n1042), .Z(n1116) );
  XNOR U4726 ( .A(n1041), .B(n1037), .Z(n1117) );
  XNOR U4727 ( .A(n1036), .B(n1032), .Z(n1118) );
  XNOR U4728 ( .A(n1031), .B(n1027), .Z(n1119) );
  XNOR U4729 ( .A(n1026), .B(n1022), .Z(n1120) );
  XNOR U4730 ( .A(n1021), .B(n1017), .Z(n1121) );
  XNOR U4731 ( .A(n1016), .B(n1012), .Z(n1122) );
  XNOR U4732 ( .A(n1011), .B(n1007), .Z(n1123) );
  XNOR U4733 ( .A(n1006), .B(n1002), .Z(n1124) );
  XNOR U4734 ( .A(n1001), .B(n997), .Z(n1125) );
  XNOR U4735 ( .A(n996), .B(n992), .Z(n1126) );
  XNOR U4736 ( .A(n991), .B(n987), .Z(n1127) );
  XNOR U4737 ( .A(n986), .B(n982), .Z(n1128) );
  XNOR U4738 ( .A(n981), .B(n977), .Z(n1129) );
  XNOR U4739 ( .A(n976), .B(n972), .Z(n1130) );
  XNOR U4740 ( .A(n971), .B(n967), .Z(n1131) );
  XOR U4741 ( .A(n966), .B(n963), .Z(n1132) );
  XOR U4742 ( .A(n1133), .B(n1134), .Z(n963) );
  XOR U4743 ( .A(n961), .B(n1135), .Z(n1134) );
  XOR U4744 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U4745 ( .A(n1138), .B(n1139), .Z(n1137) );
  NAND U4746 ( .A(a[91]), .B(b[30]), .Z(n1139) );
  AND U4747 ( .A(a[90]), .B(b[31]), .Z(n1138) );
  XOR U4748 ( .A(n1140), .B(n1136), .Z(n1133) );
  XOR U4749 ( .A(n1141), .B(n1142), .Z(n1136) );
  ANDN U4750 ( .B(n1143), .A(n1144), .Z(n1141) );
  AND U4751 ( .A(a[92]), .B(b[29]), .Z(n1140) );
  XOR U4752 ( .A(n1145), .B(n961), .Z(n962) );
  XOR U4753 ( .A(n1146), .B(n1147), .Z(n961) );
  AND U4754 ( .A(n1148), .B(n1149), .Z(n1146) );
  AND U4755 ( .A(a[93]), .B(b[28]), .Z(n1145) );
  XOR U4756 ( .A(n1150), .B(n966), .Z(n968) );
  XOR U4757 ( .A(n1151), .B(n1152), .Z(n966) );
  AND U4758 ( .A(n1153), .B(n1154), .Z(n1151) );
  AND U4759 ( .A(a[94]), .B(b[27]), .Z(n1150) );
  XOR U4760 ( .A(n1155), .B(n971), .Z(n973) );
  XOR U4761 ( .A(n1156), .B(n1157), .Z(n971) );
  AND U4762 ( .A(n1158), .B(n1159), .Z(n1156) );
  AND U4763 ( .A(b[26]), .B(a[95]), .Z(n1155) );
  XOR U4764 ( .A(n1160), .B(n976), .Z(n978) );
  XOR U4765 ( .A(n1161), .B(n1162), .Z(n976) );
  AND U4766 ( .A(n1163), .B(n1164), .Z(n1161) );
  AND U4767 ( .A(b[25]), .B(a[96]), .Z(n1160) );
  XOR U4768 ( .A(n1165), .B(n981), .Z(n983) );
  XOR U4769 ( .A(n1166), .B(n1167), .Z(n981) );
  AND U4770 ( .A(n1168), .B(n1169), .Z(n1166) );
  AND U4771 ( .A(b[24]), .B(a[97]), .Z(n1165) );
  XOR U4772 ( .A(n1170), .B(n986), .Z(n988) );
  XOR U4773 ( .A(n1171), .B(n1172), .Z(n986) );
  AND U4774 ( .A(n1173), .B(n1174), .Z(n1171) );
  AND U4775 ( .A(b[23]), .B(a[98]), .Z(n1170) );
  XOR U4776 ( .A(n1175), .B(n991), .Z(n993) );
  XOR U4777 ( .A(n1176), .B(n1177), .Z(n991) );
  AND U4778 ( .A(n1178), .B(n1179), .Z(n1176) );
  AND U4779 ( .A(b[22]), .B(a[99]), .Z(n1175) );
  XOR U4780 ( .A(n1180), .B(n996), .Z(n998) );
  XOR U4781 ( .A(n1181), .B(n1182), .Z(n996) );
  AND U4782 ( .A(n1183), .B(n1184), .Z(n1181) );
  AND U4783 ( .A(b[21]), .B(a[100]), .Z(n1180) );
  XOR U4784 ( .A(n1185), .B(n1001), .Z(n1003) );
  XOR U4785 ( .A(n1186), .B(n1187), .Z(n1001) );
  AND U4786 ( .A(n1188), .B(n1189), .Z(n1186) );
  AND U4787 ( .A(b[20]), .B(a[101]), .Z(n1185) );
  XOR U4788 ( .A(n1190), .B(n1006), .Z(n1008) );
  XOR U4789 ( .A(n1191), .B(n1192), .Z(n1006) );
  AND U4790 ( .A(n1193), .B(n1194), .Z(n1191) );
  AND U4791 ( .A(b[19]), .B(a[102]), .Z(n1190) );
  XOR U4792 ( .A(n1195), .B(n1011), .Z(n1013) );
  XOR U4793 ( .A(n1196), .B(n1197), .Z(n1011) );
  AND U4794 ( .A(n1198), .B(n1199), .Z(n1196) );
  AND U4795 ( .A(b[18]), .B(a[103]), .Z(n1195) );
  XOR U4796 ( .A(n1200), .B(n1016), .Z(n1018) );
  XOR U4797 ( .A(n1201), .B(n1202), .Z(n1016) );
  AND U4798 ( .A(n1203), .B(n1204), .Z(n1201) );
  AND U4799 ( .A(b[17]), .B(a[104]), .Z(n1200) );
  XOR U4800 ( .A(n1205), .B(n1021), .Z(n1023) );
  XOR U4801 ( .A(n1206), .B(n1207), .Z(n1021) );
  AND U4802 ( .A(n1208), .B(n1209), .Z(n1206) );
  AND U4803 ( .A(b[16]), .B(a[105]), .Z(n1205) );
  XOR U4804 ( .A(n1210), .B(n1026), .Z(n1028) );
  XOR U4805 ( .A(n1211), .B(n1212), .Z(n1026) );
  AND U4806 ( .A(n1213), .B(n1214), .Z(n1211) );
  AND U4807 ( .A(b[15]), .B(a[106]), .Z(n1210) );
  XOR U4808 ( .A(n1215), .B(n1031), .Z(n1033) );
  XOR U4809 ( .A(n1216), .B(n1217), .Z(n1031) );
  AND U4810 ( .A(n1218), .B(n1219), .Z(n1216) );
  AND U4811 ( .A(b[14]), .B(a[107]), .Z(n1215) );
  XOR U4812 ( .A(n1220), .B(n1036), .Z(n1038) );
  XOR U4813 ( .A(n1221), .B(n1222), .Z(n1036) );
  AND U4814 ( .A(n1223), .B(n1224), .Z(n1221) );
  AND U4815 ( .A(b[13]), .B(a[108]), .Z(n1220) );
  XOR U4816 ( .A(n1225), .B(n1041), .Z(n1043) );
  XOR U4817 ( .A(n1226), .B(n1227), .Z(n1041) );
  AND U4818 ( .A(n1228), .B(n1229), .Z(n1226) );
  AND U4819 ( .A(b[12]), .B(a[109]), .Z(n1225) );
  XOR U4820 ( .A(n1230), .B(n1046), .Z(n1048) );
  XOR U4821 ( .A(n1231), .B(n1232), .Z(n1046) );
  AND U4822 ( .A(n1233), .B(n1234), .Z(n1231) );
  AND U4823 ( .A(b[11]), .B(a[110]), .Z(n1230) );
  XOR U4824 ( .A(n1235), .B(n1051), .Z(n1053) );
  XOR U4825 ( .A(n1236), .B(n1237), .Z(n1051) );
  AND U4826 ( .A(n1238), .B(n1239), .Z(n1236) );
  AND U4827 ( .A(b[10]), .B(a[111]), .Z(n1235) );
  XOR U4828 ( .A(n1240), .B(n1056), .Z(n1058) );
  XOR U4829 ( .A(n1241), .B(n1242), .Z(n1056) );
  AND U4830 ( .A(n1243), .B(n1244), .Z(n1241) );
  AND U4831 ( .A(b[9]), .B(a[112]), .Z(n1240) );
  XOR U4832 ( .A(n1245), .B(n1061), .Z(n1063) );
  XOR U4833 ( .A(n1246), .B(n1247), .Z(n1061) );
  AND U4834 ( .A(n1248), .B(n1249), .Z(n1246) );
  AND U4835 ( .A(b[8]), .B(a[113]), .Z(n1245) );
  XOR U4836 ( .A(n1250), .B(n1066), .Z(n1068) );
  XOR U4837 ( .A(n1251), .B(n1252), .Z(n1066) );
  AND U4838 ( .A(n1253), .B(n1254), .Z(n1251) );
  AND U4839 ( .A(b[7]), .B(a[114]), .Z(n1250) );
  XOR U4840 ( .A(n1255), .B(n1071), .Z(n1073) );
  XOR U4841 ( .A(n1256), .B(n1257), .Z(n1071) );
  AND U4842 ( .A(n1258), .B(n1259), .Z(n1256) );
  AND U4843 ( .A(b[6]), .B(a[115]), .Z(n1255) );
  XOR U4844 ( .A(n1260), .B(n1076), .Z(n1078) );
  XOR U4845 ( .A(n1261), .B(n1262), .Z(n1076) );
  AND U4846 ( .A(n1263), .B(n1264), .Z(n1261) );
  AND U4847 ( .A(b[5]), .B(a[116]), .Z(n1260) );
  XOR U4848 ( .A(n1265), .B(n1081), .Z(n1083) );
  XOR U4849 ( .A(n1266), .B(n1267), .Z(n1081) );
  AND U4850 ( .A(n1268), .B(n1269), .Z(n1266) );
  AND U4851 ( .A(b[4]), .B(a[117]), .Z(n1265) );
  XNOR U4852 ( .A(n1270), .B(n1271), .Z(n1095) );
  NANDN U4853 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U4854 ( .A(n1274), .B(n1086), .Z(n1088) );
  XNOR U4855 ( .A(n1275), .B(n1276), .Z(n1086) );
  AND U4856 ( .A(n1277), .B(n1278), .Z(n1275) );
  AND U4857 ( .A(b[3]), .B(a[118]), .Z(n1274) );
  XNOR U4858 ( .A(n1279), .B(n1280), .Z(swire[120]) );
  XOR U4859 ( .A(n1106), .B(n1281), .Z(n1280) );
  XOR U4860 ( .A(n1105), .B(n1279), .Z(n1281) );
  NAND U4861 ( .A(a[120]), .B(b[0]), .Z(n1105) );
  XNOR U4862 ( .A(n1272), .B(n1273), .Z(n1106) );
  XOR U4863 ( .A(n1270), .B(n1282), .Z(n1273) );
  NAND U4864 ( .A(b[1]), .B(a[119]), .Z(n1282) );
  XOR U4865 ( .A(n1278), .B(n1283), .Z(n1272) );
  XOR U4866 ( .A(n1270), .B(n1277), .Z(n1283) );
  XNOR U4867 ( .A(n1284), .B(n1276), .Z(n1277) );
  AND U4868 ( .A(b[2]), .B(a[118]), .Z(n1284) );
  NANDN U4869 ( .A(n1285), .B(n1286), .Z(n1270) );
  XOR U4870 ( .A(n1276), .B(n1268), .Z(n1287) );
  XNOR U4871 ( .A(n1267), .B(n1263), .Z(n1288) );
  XNOR U4872 ( .A(n1262), .B(n1258), .Z(n1289) );
  XNOR U4873 ( .A(n1257), .B(n1253), .Z(n1290) );
  XNOR U4874 ( .A(n1252), .B(n1248), .Z(n1291) );
  XNOR U4875 ( .A(n1247), .B(n1243), .Z(n1292) );
  XNOR U4876 ( .A(n1242), .B(n1238), .Z(n1293) );
  XNOR U4877 ( .A(n1237), .B(n1233), .Z(n1294) );
  XNOR U4878 ( .A(n1232), .B(n1228), .Z(n1295) );
  XNOR U4879 ( .A(n1227), .B(n1223), .Z(n1296) );
  XNOR U4880 ( .A(n1222), .B(n1218), .Z(n1297) );
  XNOR U4881 ( .A(n1217), .B(n1213), .Z(n1298) );
  XNOR U4882 ( .A(n1212), .B(n1208), .Z(n1299) );
  XNOR U4883 ( .A(n1207), .B(n1203), .Z(n1300) );
  XNOR U4884 ( .A(n1202), .B(n1198), .Z(n1301) );
  XNOR U4885 ( .A(n1197), .B(n1193), .Z(n1302) );
  XNOR U4886 ( .A(n1192), .B(n1188), .Z(n1303) );
  XNOR U4887 ( .A(n1187), .B(n1183), .Z(n1304) );
  XNOR U4888 ( .A(n1182), .B(n1178), .Z(n1305) );
  XNOR U4889 ( .A(n1177), .B(n1173), .Z(n1306) );
  XNOR U4890 ( .A(n1172), .B(n1168), .Z(n1307) );
  XNOR U4891 ( .A(n1167), .B(n1163), .Z(n1308) );
  XNOR U4892 ( .A(n1162), .B(n1158), .Z(n1309) );
  XNOR U4893 ( .A(n1157), .B(n1153), .Z(n1310) );
  XNOR U4894 ( .A(n1152), .B(n1148), .Z(n1311) );
  XOR U4895 ( .A(n1147), .B(n1144), .Z(n1312) );
  XOR U4896 ( .A(n1313), .B(n1314), .Z(n1144) );
  XOR U4897 ( .A(n1142), .B(n1315), .Z(n1314) );
  XOR U4898 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U4899 ( .A(n1318), .B(n1319), .Z(n1317) );
  NAND U4900 ( .A(a[90]), .B(b[30]), .Z(n1319) );
  AND U4901 ( .A(a[89]), .B(b[31]), .Z(n1318) );
  XOR U4902 ( .A(n1320), .B(n1316), .Z(n1313) );
  XOR U4903 ( .A(n1321), .B(n1322), .Z(n1316) );
  ANDN U4904 ( .B(n1323), .A(n1324), .Z(n1321) );
  AND U4905 ( .A(a[91]), .B(b[29]), .Z(n1320) );
  XOR U4906 ( .A(n1325), .B(n1142), .Z(n1143) );
  XOR U4907 ( .A(n1326), .B(n1327), .Z(n1142) );
  AND U4908 ( .A(n1328), .B(n1329), .Z(n1326) );
  AND U4909 ( .A(a[92]), .B(b[28]), .Z(n1325) );
  XOR U4910 ( .A(n1330), .B(n1147), .Z(n1149) );
  XOR U4911 ( .A(n1331), .B(n1332), .Z(n1147) );
  AND U4912 ( .A(n1333), .B(n1334), .Z(n1331) );
  AND U4913 ( .A(a[93]), .B(b[27]), .Z(n1330) );
  XOR U4914 ( .A(n1335), .B(n1152), .Z(n1154) );
  XOR U4915 ( .A(n1336), .B(n1337), .Z(n1152) );
  AND U4916 ( .A(n1338), .B(n1339), .Z(n1336) );
  AND U4917 ( .A(a[94]), .B(b[26]), .Z(n1335) );
  XOR U4918 ( .A(n1340), .B(n1157), .Z(n1159) );
  XOR U4919 ( .A(n1341), .B(n1342), .Z(n1157) );
  AND U4920 ( .A(n1343), .B(n1344), .Z(n1341) );
  AND U4921 ( .A(b[25]), .B(a[95]), .Z(n1340) );
  XOR U4922 ( .A(n1345), .B(n1162), .Z(n1164) );
  XOR U4923 ( .A(n1346), .B(n1347), .Z(n1162) );
  AND U4924 ( .A(n1348), .B(n1349), .Z(n1346) );
  AND U4925 ( .A(b[24]), .B(a[96]), .Z(n1345) );
  XOR U4926 ( .A(n1350), .B(n1167), .Z(n1169) );
  XOR U4927 ( .A(n1351), .B(n1352), .Z(n1167) );
  AND U4928 ( .A(n1353), .B(n1354), .Z(n1351) );
  AND U4929 ( .A(b[23]), .B(a[97]), .Z(n1350) );
  XOR U4930 ( .A(n1355), .B(n1172), .Z(n1174) );
  XOR U4931 ( .A(n1356), .B(n1357), .Z(n1172) );
  AND U4932 ( .A(n1358), .B(n1359), .Z(n1356) );
  AND U4933 ( .A(b[22]), .B(a[98]), .Z(n1355) );
  XOR U4934 ( .A(n1360), .B(n1177), .Z(n1179) );
  XOR U4935 ( .A(n1361), .B(n1362), .Z(n1177) );
  AND U4936 ( .A(n1363), .B(n1364), .Z(n1361) );
  AND U4937 ( .A(b[21]), .B(a[99]), .Z(n1360) );
  XOR U4938 ( .A(n1365), .B(n1182), .Z(n1184) );
  XOR U4939 ( .A(n1366), .B(n1367), .Z(n1182) );
  AND U4940 ( .A(n1368), .B(n1369), .Z(n1366) );
  AND U4941 ( .A(b[20]), .B(a[100]), .Z(n1365) );
  XOR U4942 ( .A(n1370), .B(n1187), .Z(n1189) );
  XOR U4943 ( .A(n1371), .B(n1372), .Z(n1187) );
  AND U4944 ( .A(n1373), .B(n1374), .Z(n1371) );
  AND U4945 ( .A(b[19]), .B(a[101]), .Z(n1370) );
  XOR U4946 ( .A(n1375), .B(n1192), .Z(n1194) );
  XOR U4947 ( .A(n1376), .B(n1377), .Z(n1192) );
  AND U4948 ( .A(n1378), .B(n1379), .Z(n1376) );
  AND U4949 ( .A(b[18]), .B(a[102]), .Z(n1375) );
  XOR U4950 ( .A(n1380), .B(n1197), .Z(n1199) );
  XOR U4951 ( .A(n1381), .B(n1382), .Z(n1197) );
  AND U4952 ( .A(n1383), .B(n1384), .Z(n1381) );
  AND U4953 ( .A(b[17]), .B(a[103]), .Z(n1380) );
  XOR U4954 ( .A(n1385), .B(n1202), .Z(n1204) );
  XOR U4955 ( .A(n1386), .B(n1387), .Z(n1202) );
  AND U4956 ( .A(n1388), .B(n1389), .Z(n1386) );
  AND U4957 ( .A(b[16]), .B(a[104]), .Z(n1385) );
  XOR U4958 ( .A(n1390), .B(n1207), .Z(n1209) );
  XOR U4959 ( .A(n1391), .B(n1392), .Z(n1207) );
  AND U4960 ( .A(n1393), .B(n1394), .Z(n1391) );
  AND U4961 ( .A(b[15]), .B(a[105]), .Z(n1390) );
  XOR U4962 ( .A(n1395), .B(n1212), .Z(n1214) );
  XOR U4963 ( .A(n1396), .B(n1397), .Z(n1212) );
  AND U4964 ( .A(n1398), .B(n1399), .Z(n1396) );
  AND U4965 ( .A(b[14]), .B(a[106]), .Z(n1395) );
  XOR U4966 ( .A(n1400), .B(n1217), .Z(n1219) );
  XOR U4967 ( .A(n1401), .B(n1402), .Z(n1217) );
  AND U4968 ( .A(n1403), .B(n1404), .Z(n1401) );
  AND U4969 ( .A(b[13]), .B(a[107]), .Z(n1400) );
  XOR U4970 ( .A(n1405), .B(n1222), .Z(n1224) );
  XOR U4971 ( .A(n1406), .B(n1407), .Z(n1222) );
  AND U4972 ( .A(n1408), .B(n1409), .Z(n1406) );
  AND U4973 ( .A(b[12]), .B(a[108]), .Z(n1405) );
  XOR U4974 ( .A(n1410), .B(n1227), .Z(n1229) );
  XOR U4975 ( .A(n1411), .B(n1412), .Z(n1227) );
  AND U4976 ( .A(n1413), .B(n1414), .Z(n1411) );
  AND U4977 ( .A(b[11]), .B(a[109]), .Z(n1410) );
  XOR U4978 ( .A(n1415), .B(n1232), .Z(n1234) );
  XOR U4979 ( .A(n1416), .B(n1417), .Z(n1232) );
  AND U4980 ( .A(n1418), .B(n1419), .Z(n1416) );
  AND U4981 ( .A(b[10]), .B(a[110]), .Z(n1415) );
  XOR U4982 ( .A(n1420), .B(n1237), .Z(n1239) );
  XOR U4983 ( .A(n1421), .B(n1422), .Z(n1237) );
  AND U4984 ( .A(n1423), .B(n1424), .Z(n1421) );
  AND U4985 ( .A(b[9]), .B(a[111]), .Z(n1420) );
  XOR U4986 ( .A(n1425), .B(n1242), .Z(n1244) );
  XOR U4987 ( .A(n1426), .B(n1427), .Z(n1242) );
  AND U4988 ( .A(n1428), .B(n1429), .Z(n1426) );
  AND U4989 ( .A(b[8]), .B(a[112]), .Z(n1425) );
  XOR U4990 ( .A(n1430), .B(n1247), .Z(n1249) );
  XOR U4991 ( .A(n1431), .B(n1432), .Z(n1247) );
  AND U4992 ( .A(n1433), .B(n1434), .Z(n1431) );
  AND U4993 ( .A(b[7]), .B(a[113]), .Z(n1430) );
  XOR U4994 ( .A(n1435), .B(n1252), .Z(n1254) );
  XOR U4995 ( .A(n1436), .B(n1437), .Z(n1252) );
  AND U4996 ( .A(n1438), .B(n1439), .Z(n1436) );
  AND U4997 ( .A(b[6]), .B(a[114]), .Z(n1435) );
  XOR U4998 ( .A(n1440), .B(n1257), .Z(n1259) );
  XOR U4999 ( .A(n1441), .B(n1442), .Z(n1257) );
  AND U5000 ( .A(n1443), .B(n1444), .Z(n1441) );
  AND U5001 ( .A(b[5]), .B(a[115]), .Z(n1440) );
  XOR U5002 ( .A(n1445), .B(n1262), .Z(n1264) );
  XOR U5003 ( .A(n1446), .B(n1447), .Z(n1262) );
  AND U5004 ( .A(n1448), .B(n1449), .Z(n1446) );
  AND U5005 ( .A(b[4]), .B(a[116]), .Z(n1445) );
  XNOR U5006 ( .A(n1450), .B(n1451), .Z(n1276) );
  NANDN U5007 ( .A(n1452), .B(n1453), .Z(n1451) );
  XOR U5008 ( .A(n1454), .B(n1267), .Z(n1269) );
  XNOR U5009 ( .A(n1455), .B(n1456), .Z(n1267) );
  AND U5010 ( .A(n1457), .B(n1458), .Z(n1455) );
  AND U5011 ( .A(b[3]), .B(a[117]), .Z(n1454) );
  XOR U5012 ( .A(n1459), .B(n1460), .Z(swire[119]) );
  XOR U5013 ( .A(n1286), .B(n1462), .Z(n1460) );
  XOR U5014 ( .A(n1285), .B(n1461), .Z(n1462) );
  IV U5015 ( .A(n1459), .Z(n1461) );
  NAND U5016 ( .A(a[119]), .B(b[0]), .Z(n1285) );
  XNOR U5017 ( .A(n1452), .B(n1453), .Z(n1286) );
  XOR U5018 ( .A(n1450), .B(n1463), .Z(n1453) );
  NAND U5019 ( .A(b[1]), .B(a[118]), .Z(n1463) );
  XOR U5020 ( .A(n1458), .B(n1464), .Z(n1452) );
  XOR U5021 ( .A(n1450), .B(n1457), .Z(n1464) );
  XNOR U5022 ( .A(n1465), .B(n1456), .Z(n1457) );
  AND U5023 ( .A(b[2]), .B(a[117]), .Z(n1465) );
  NANDN U5024 ( .A(n1466), .B(n1467), .Z(n1450) );
  XOR U5025 ( .A(n1456), .B(n1448), .Z(n1468) );
  XNOR U5026 ( .A(n1447), .B(n1443), .Z(n1469) );
  XNOR U5027 ( .A(n1442), .B(n1438), .Z(n1470) );
  XNOR U5028 ( .A(n1437), .B(n1433), .Z(n1471) );
  XNOR U5029 ( .A(n1432), .B(n1428), .Z(n1472) );
  XNOR U5030 ( .A(n1427), .B(n1423), .Z(n1473) );
  XNOR U5031 ( .A(n1422), .B(n1418), .Z(n1474) );
  XNOR U5032 ( .A(n1417), .B(n1413), .Z(n1475) );
  XNOR U5033 ( .A(n1412), .B(n1408), .Z(n1476) );
  XNOR U5034 ( .A(n1407), .B(n1403), .Z(n1477) );
  XNOR U5035 ( .A(n1402), .B(n1398), .Z(n1478) );
  XNOR U5036 ( .A(n1397), .B(n1393), .Z(n1479) );
  XNOR U5037 ( .A(n1392), .B(n1388), .Z(n1480) );
  XNOR U5038 ( .A(n1387), .B(n1383), .Z(n1481) );
  XNOR U5039 ( .A(n1382), .B(n1378), .Z(n1482) );
  XNOR U5040 ( .A(n1377), .B(n1373), .Z(n1483) );
  XNOR U5041 ( .A(n1372), .B(n1368), .Z(n1484) );
  XNOR U5042 ( .A(n1367), .B(n1363), .Z(n1485) );
  XNOR U5043 ( .A(n1362), .B(n1358), .Z(n1486) );
  XNOR U5044 ( .A(n1357), .B(n1353), .Z(n1487) );
  XNOR U5045 ( .A(n1352), .B(n1348), .Z(n1488) );
  XNOR U5046 ( .A(n1347), .B(n1343), .Z(n1489) );
  XNOR U5047 ( .A(n1342), .B(n1338), .Z(n1490) );
  XNOR U5048 ( .A(n1337), .B(n1333), .Z(n1491) );
  XNOR U5049 ( .A(n1332), .B(n1328), .Z(n1492) );
  XOR U5050 ( .A(n1327), .B(n1324), .Z(n1493) );
  XOR U5051 ( .A(n1494), .B(n1495), .Z(n1324) );
  XOR U5052 ( .A(n1322), .B(n1496), .Z(n1495) );
  XOR U5053 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U5054 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U5055 ( .A(a[89]), .B(b[30]), .Z(n1500) );
  AND U5056 ( .A(a[88]), .B(b[31]), .Z(n1499) );
  XOR U5057 ( .A(n1501), .B(n1497), .Z(n1494) );
  XOR U5058 ( .A(n1502), .B(n1503), .Z(n1497) );
  ANDN U5059 ( .B(n1504), .A(n1505), .Z(n1502) );
  AND U5060 ( .A(a[90]), .B(b[29]), .Z(n1501) );
  XOR U5061 ( .A(n1506), .B(n1322), .Z(n1323) );
  XOR U5062 ( .A(n1507), .B(n1508), .Z(n1322) );
  AND U5063 ( .A(n1509), .B(n1510), .Z(n1507) );
  AND U5064 ( .A(a[91]), .B(b[28]), .Z(n1506) );
  XOR U5065 ( .A(n1511), .B(n1327), .Z(n1329) );
  XOR U5066 ( .A(n1512), .B(n1513), .Z(n1327) );
  AND U5067 ( .A(n1514), .B(n1515), .Z(n1512) );
  AND U5068 ( .A(a[92]), .B(b[27]), .Z(n1511) );
  XOR U5069 ( .A(n1516), .B(n1332), .Z(n1334) );
  XOR U5070 ( .A(n1517), .B(n1518), .Z(n1332) );
  AND U5071 ( .A(n1519), .B(n1520), .Z(n1517) );
  AND U5072 ( .A(a[93]), .B(b[26]), .Z(n1516) );
  XOR U5073 ( .A(n1521), .B(n1337), .Z(n1339) );
  XOR U5074 ( .A(n1522), .B(n1523), .Z(n1337) );
  AND U5075 ( .A(n1524), .B(n1525), .Z(n1522) );
  AND U5076 ( .A(a[94]), .B(b[25]), .Z(n1521) );
  XOR U5077 ( .A(n1526), .B(n1342), .Z(n1344) );
  XOR U5078 ( .A(n1527), .B(n1528), .Z(n1342) );
  AND U5079 ( .A(n1529), .B(n1530), .Z(n1527) );
  AND U5080 ( .A(b[24]), .B(a[95]), .Z(n1526) );
  XOR U5081 ( .A(n1531), .B(n1347), .Z(n1349) );
  XOR U5082 ( .A(n1532), .B(n1533), .Z(n1347) );
  AND U5083 ( .A(n1534), .B(n1535), .Z(n1532) );
  AND U5084 ( .A(b[23]), .B(a[96]), .Z(n1531) );
  XOR U5085 ( .A(n1536), .B(n1352), .Z(n1354) );
  XOR U5086 ( .A(n1537), .B(n1538), .Z(n1352) );
  AND U5087 ( .A(n1539), .B(n1540), .Z(n1537) );
  AND U5088 ( .A(b[22]), .B(a[97]), .Z(n1536) );
  XOR U5089 ( .A(n1541), .B(n1357), .Z(n1359) );
  XOR U5090 ( .A(n1542), .B(n1543), .Z(n1357) );
  AND U5091 ( .A(n1544), .B(n1545), .Z(n1542) );
  AND U5092 ( .A(b[21]), .B(a[98]), .Z(n1541) );
  XOR U5093 ( .A(n1546), .B(n1362), .Z(n1364) );
  XOR U5094 ( .A(n1547), .B(n1548), .Z(n1362) );
  AND U5095 ( .A(n1549), .B(n1550), .Z(n1547) );
  AND U5096 ( .A(b[20]), .B(a[99]), .Z(n1546) );
  XOR U5097 ( .A(n1551), .B(n1367), .Z(n1369) );
  XOR U5098 ( .A(n1552), .B(n1553), .Z(n1367) );
  AND U5099 ( .A(n1554), .B(n1555), .Z(n1552) );
  AND U5100 ( .A(b[19]), .B(a[100]), .Z(n1551) );
  XOR U5101 ( .A(n1556), .B(n1372), .Z(n1374) );
  XOR U5102 ( .A(n1557), .B(n1558), .Z(n1372) );
  AND U5103 ( .A(n1559), .B(n1560), .Z(n1557) );
  AND U5104 ( .A(b[18]), .B(a[101]), .Z(n1556) );
  XOR U5105 ( .A(n1561), .B(n1377), .Z(n1379) );
  XOR U5106 ( .A(n1562), .B(n1563), .Z(n1377) );
  AND U5107 ( .A(n1564), .B(n1565), .Z(n1562) );
  AND U5108 ( .A(b[17]), .B(a[102]), .Z(n1561) );
  XOR U5109 ( .A(n1566), .B(n1382), .Z(n1384) );
  XOR U5110 ( .A(n1567), .B(n1568), .Z(n1382) );
  AND U5111 ( .A(n1569), .B(n1570), .Z(n1567) );
  AND U5112 ( .A(b[16]), .B(a[103]), .Z(n1566) );
  XOR U5113 ( .A(n1571), .B(n1387), .Z(n1389) );
  XOR U5114 ( .A(n1572), .B(n1573), .Z(n1387) );
  AND U5115 ( .A(n1574), .B(n1575), .Z(n1572) );
  AND U5116 ( .A(b[15]), .B(a[104]), .Z(n1571) );
  XOR U5117 ( .A(n1576), .B(n1392), .Z(n1394) );
  XOR U5118 ( .A(n1577), .B(n1578), .Z(n1392) );
  AND U5119 ( .A(n1579), .B(n1580), .Z(n1577) );
  AND U5120 ( .A(b[14]), .B(a[105]), .Z(n1576) );
  XOR U5121 ( .A(n1581), .B(n1397), .Z(n1399) );
  XOR U5122 ( .A(n1582), .B(n1583), .Z(n1397) );
  AND U5123 ( .A(n1584), .B(n1585), .Z(n1582) );
  AND U5124 ( .A(b[13]), .B(a[106]), .Z(n1581) );
  XOR U5125 ( .A(n1586), .B(n1402), .Z(n1404) );
  XOR U5126 ( .A(n1587), .B(n1588), .Z(n1402) );
  AND U5127 ( .A(n1589), .B(n1590), .Z(n1587) );
  AND U5128 ( .A(b[12]), .B(a[107]), .Z(n1586) );
  XOR U5129 ( .A(n1591), .B(n1407), .Z(n1409) );
  XOR U5130 ( .A(n1592), .B(n1593), .Z(n1407) );
  AND U5131 ( .A(n1594), .B(n1595), .Z(n1592) );
  AND U5132 ( .A(b[11]), .B(a[108]), .Z(n1591) );
  XOR U5133 ( .A(n1596), .B(n1412), .Z(n1414) );
  XOR U5134 ( .A(n1597), .B(n1598), .Z(n1412) );
  AND U5135 ( .A(n1599), .B(n1600), .Z(n1597) );
  AND U5136 ( .A(b[10]), .B(a[109]), .Z(n1596) );
  XOR U5137 ( .A(n1601), .B(n1417), .Z(n1419) );
  XOR U5138 ( .A(n1602), .B(n1603), .Z(n1417) );
  AND U5139 ( .A(n1604), .B(n1605), .Z(n1602) );
  AND U5140 ( .A(b[9]), .B(a[110]), .Z(n1601) );
  XOR U5141 ( .A(n1606), .B(n1422), .Z(n1424) );
  XOR U5142 ( .A(n1607), .B(n1608), .Z(n1422) );
  AND U5143 ( .A(n1609), .B(n1610), .Z(n1607) );
  AND U5144 ( .A(b[8]), .B(a[111]), .Z(n1606) );
  XOR U5145 ( .A(n1611), .B(n1427), .Z(n1429) );
  XOR U5146 ( .A(n1612), .B(n1613), .Z(n1427) );
  AND U5147 ( .A(n1614), .B(n1615), .Z(n1612) );
  AND U5148 ( .A(b[7]), .B(a[112]), .Z(n1611) );
  XOR U5149 ( .A(n1616), .B(n1432), .Z(n1434) );
  XOR U5150 ( .A(n1617), .B(n1618), .Z(n1432) );
  AND U5151 ( .A(n1619), .B(n1620), .Z(n1617) );
  AND U5152 ( .A(b[6]), .B(a[113]), .Z(n1616) );
  XOR U5153 ( .A(n1621), .B(n1437), .Z(n1439) );
  XOR U5154 ( .A(n1622), .B(n1623), .Z(n1437) );
  AND U5155 ( .A(n1624), .B(n1625), .Z(n1622) );
  AND U5156 ( .A(b[5]), .B(a[114]), .Z(n1621) );
  XOR U5157 ( .A(n1626), .B(n1442), .Z(n1444) );
  XOR U5158 ( .A(n1627), .B(n1628), .Z(n1442) );
  AND U5159 ( .A(n1629), .B(n1630), .Z(n1627) );
  AND U5160 ( .A(b[4]), .B(a[115]), .Z(n1626) );
  XNOR U5161 ( .A(n1631), .B(n1632), .Z(n1456) );
  NANDN U5162 ( .A(n1633), .B(n1634), .Z(n1632) );
  XOR U5163 ( .A(n1635), .B(n1447), .Z(n1449) );
  XNOR U5164 ( .A(n1636), .B(n1637), .Z(n1447) );
  AND U5165 ( .A(n1638), .B(n1639), .Z(n1636) );
  AND U5166 ( .A(b[3]), .B(a[116]), .Z(n1635) );
  XNOR U5167 ( .A(n1640), .B(n1641), .Z(swire[118]) );
  XOR U5168 ( .A(n1467), .B(n1642), .Z(n1641) );
  XOR U5169 ( .A(n1466), .B(n1640), .Z(n1642) );
  NAND U5170 ( .A(a[118]), .B(b[0]), .Z(n1466) );
  XNOR U5171 ( .A(n1633), .B(n1634), .Z(n1467) );
  XOR U5172 ( .A(n1631), .B(n1643), .Z(n1634) );
  NAND U5173 ( .A(b[1]), .B(a[117]), .Z(n1643) );
  XOR U5174 ( .A(n1639), .B(n1644), .Z(n1633) );
  XOR U5175 ( .A(n1631), .B(n1638), .Z(n1644) );
  XNOR U5176 ( .A(n1645), .B(n1637), .Z(n1638) );
  AND U5177 ( .A(b[2]), .B(a[116]), .Z(n1645) );
  NANDN U5178 ( .A(n1646), .B(n1647), .Z(n1631) );
  XOR U5179 ( .A(n1637), .B(n1629), .Z(n1648) );
  XNOR U5180 ( .A(n1628), .B(n1624), .Z(n1649) );
  XNOR U5181 ( .A(n1623), .B(n1619), .Z(n1650) );
  XNOR U5182 ( .A(n1618), .B(n1614), .Z(n1651) );
  XNOR U5183 ( .A(n1613), .B(n1609), .Z(n1652) );
  XNOR U5184 ( .A(n1608), .B(n1604), .Z(n1653) );
  XNOR U5185 ( .A(n1603), .B(n1599), .Z(n1654) );
  XNOR U5186 ( .A(n1598), .B(n1594), .Z(n1655) );
  XNOR U5187 ( .A(n1593), .B(n1589), .Z(n1656) );
  XNOR U5188 ( .A(n1588), .B(n1584), .Z(n1657) );
  XNOR U5189 ( .A(n1583), .B(n1579), .Z(n1658) );
  XNOR U5190 ( .A(n1578), .B(n1574), .Z(n1659) );
  XNOR U5191 ( .A(n1573), .B(n1569), .Z(n1660) );
  XNOR U5192 ( .A(n1568), .B(n1564), .Z(n1661) );
  XNOR U5193 ( .A(n1563), .B(n1559), .Z(n1662) );
  XNOR U5194 ( .A(n1558), .B(n1554), .Z(n1663) );
  XNOR U5195 ( .A(n1553), .B(n1549), .Z(n1664) );
  XNOR U5196 ( .A(n1548), .B(n1544), .Z(n1665) );
  XNOR U5197 ( .A(n1543), .B(n1539), .Z(n1666) );
  XNOR U5198 ( .A(n1538), .B(n1534), .Z(n1667) );
  XNOR U5199 ( .A(n1533), .B(n1529), .Z(n1668) );
  XNOR U5200 ( .A(n1528), .B(n1524), .Z(n1669) );
  XNOR U5201 ( .A(n1523), .B(n1519), .Z(n1670) );
  XNOR U5202 ( .A(n1518), .B(n1514), .Z(n1671) );
  XNOR U5203 ( .A(n1513), .B(n1509), .Z(n1672) );
  XOR U5204 ( .A(n1508), .B(n1505), .Z(n1673) );
  XOR U5205 ( .A(n1674), .B(n1675), .Z(n1505) );
  XOR U5206 ( .A(n1503), .B(n1676), .Z(n1675) );
  XOR U5207 ( .A(n1677), .B(n1678), .Z(n1676) );
  XOR U5208 ( .A(n1679), .B(n1680), .Z(n1678) );
  NAND U5209 ( .A(a[88]), .B(b[30]), .Z(n1680) );
  AND U5210 ( .A(a[87]), .B(b[31]), .Z(n1679) );
  XOR U5211 ( .A(n1681), .B(n1677), .Z(n1674) );
  XOR U5212 ( .A(n1682), .B(n1683), .Z(n1677) );
  ANDN U5213 ( .B(n1684), .A(n1685), .Z(n1682) );
  AND U5214 ( .A(a[89]), .B(b[29]), .Z(n1681) );
  XOR U5215 ( .A(n1686), .B(n1503), .Z(n1504) );
  XOR U5216 ( .A(n1687), .B(n1688), .Z(n1503) );
  AND U5217 ( .A(n1689), .B(n1690), .Z(n1687) );
  AND U5218 ( .A(a[90]), .B(b[28]), .Z(n1686) );
  XOR U5219 ( .A(n1691), .B(n1508), .Z(n1510) );
  XOR U5220 ( .A(n1692), .B(n1693), .Z(n1508) );
  AND U5221 ( .A(n1694), .B(n1695), .Z(n1692) );
  AND U5222 ( .A(a[91]), .B(b[27]), .Z(n1691) );
  XOR U5223 ( .A(n1696), .B(n1513), .Z(n1515) );
  XOR U5224 ( .A(n1697), .B(n1698), .Z(n1513) );
  AND U5225 ( .A(n1699), .B(n1700), .Z(n1697) );
  AND U5226 ( .A(a[92]), .B(b[26]), .Z(n1696) );
  XOR U5227 ( .A(n1701), .B(n1518), .Z(n1520) );
  XOR U5228 ( .A(n1702), .B(n1703), .Z(n1518) );
  AND U5229 ( .A(n1704), .B(n1705), .Z(n1702) );
  AND U5230 ( .A(a[93]), .B(b[25]), .Z(n1701) );
  XOR U5231 ( .A(n1706), .B(n1523), .Z(n1525) );
  XOR U5232 ( .A(n1707), .B(n1708), .Z(n1523) );
  AND U5233 ( .A(n1709), .B(n1710), .Z(n1707) );
  AND U5234 ( .A(a[94]), .B(b[24]), .Z(n1706) );
  XOR U5235 ( .A(n1711), .B(n1528), .Z(n1530) );
  XOR U5236 ( .A(n1712), .B(n1713), .Z(n1528) );
  AND U5237 ( .A(n1714), .B(n1715), .Z(n1712) );
  AND U5238 ( .A(b[23]), .B(a[95]), .Z(n1711) );
  XOR U5239 ( .A(n1716), .B(n1533), .Z(n1535) );
  XOR U5240 ( .A(n1717), .B(n1718), .Z(n1533) );
  AND U5241 ( .A(n1719), .B(n1720), .Z(n1717) );
  AND U5242 ( .A(b[22]), .B(a[96]), .Z(n1716) );
  XOR U5243 ( .A(n1721), .B(n1538), .Z(n1540) );
  XOR U5244 ( .A(n1722), .B(n1723), .Z(n1538) );
  AND U5245 ( .A(n1724), .B(n1725), .Z(n1722) );
  AND U5246 ( .A(b[21]), .B(a[97]), .Z(n1721) );
  XOR U5247 ( .A(n1726), .B(n1543), .Z(n1545) );
  XOR U5248 ( .A(n1727), .B(n1728), .Z(n1543) );
  AND U5249 ( .A(n1729), .B(n1730), .Z(n1727) );
  AND U5250 ( .A(b[20]), .B(a[98]), .Z(n1726) );
  XOR U5251 ( .A(n1731), .B(n1548), .Z(n1550) );
  XOR U5252 ( .A(n1732), .B(n1733), .Z(n1548) );
  AND U5253 ( .A(n1734), .B(n1735), .Z(n1732) );
  AND U5254 ( .A(b[19]), .B(a[99]), .Z(n1731) );
  XOR U5255 ( .A(n1736), .B(n1553), .Z(n1555) );
  XOR U5256 ( .A(n1737), .B(n1738), .Z(n1553) );
  AND U5257 ( .A(n1739), .B(n1740), .Z(n1737) );
  AND U5258 ( .A(b[18]), .B(a[100]), .Z(n1736) );
  XOR U5259 ( .A(n1741), .B(n1558), .Z(n1560) );
  XOR U5260 ( .A(n1742), .B(n1743), .Z(n1558) );
  AND U5261 ( .A(n1744), .B(n1745), .Z(n1742) );
  AND U5262 ( .A(b[17]), .B(a[101]), .Z(n1741) );
  XOR U5263 ( .A(n1746), .B(n1563), .Z(n1565) );
  XOR U5264 ( .A(n1747), .B(n1748), .Z(n1563) );
  AND U5265 ( .A(n1749), .B(n1750), .Z(n1747) );
  AND U5266 ( .A(b[16]), .B(a[102]), .Z(n1746) );
  XOR U5267 ( .A(n1751), .B(n1568), .Z(n1570) );
  XOR U5268 ( .A(n1752), .B(n1753), .Z(n1568) );
  AND U5269 ( .A(n1754), .B(n1755), .Z(n1752) );
  AND U5270 ( .A(b[15]), .B(a[103]), .Z(n1751) );
  XOR U5271 ( .A(n1756), .B(n1573), .Z(n1575) );
  XOR U5272 ( .A(n1757), .B(n1758), .Z(n1573) );
  AND U5273 ( .A(n1759), .B(n1760), .Z(n1757) );
  AND U5274 ( .A(b[14]), .B(a[104]), .Z(n1756) );
  XOR U5275 ( .A(n1761), .B(n1578), .Z(n1580) );
  XOR U5276 ( .A(n1762), .B(n1763), .Z(n1578) );
  AND U5277 ( .A(n1764), .B(n1765), .Z(n1762) );
  AND U5278 ( .A(b[13]), .B(a[105]), .Z(n1761) );
  XOR U5279 ( .A(n1766), .B(n1583), .Z(n1585) );
  XOR U5280 ( .A(n1767), .B(n1768), .Z(n1583) );
  AND U5281 ( .A(n1769), .B(n1770), .Z(n1767) );
  AND U5282 ( .A(b[12]), .B(a[106]), .Z(n1766) );
  XOR U5283 ( .A(n1771), .B(n1588), .Z(n1590) );
  XOR U5284 ( .A(n1772), .B(n1773), .Z(n1588) );
  AND U5285 ( .A(n1774), .B(n1775), .Z(n1772) );
  AND U5286 ( .A(b[11]), .B(a[107]), .Z(n1771) );
  XOR U5287 ( .A(n1776), .B(n1593), .Z(n1595) );
  XOR U5288 ( .A(n1777), .B(n1778), .Z(n1593) );
  AND U5289 ( .A(n1779), .B(n1780), .Z(n1777) );
  AND U5290 ( .A(b[10]), .B(a[108]), .Z(n1776) );
  XOR U5291 ( .A(n1781), .B(n1598), .Z(n1600) );
  XOR U5292 ( .A(n1782), .B(n1783), .Z(n1598) );
  AND U5293 ( .A(n1784), .B(n1785), .Z(n1782) );
  AND U5294 ( .A(b[9]), .B(a[109]), .Z(n1781) );
  XOR U5295 ( .A(n1786), .B(n1603), .Z(n1605) );
  XOR U5296 ( .A(n1787), .B(n1788), .Z(n1603) );
  AND U5297 ( .A(n1789), .B(n1790), .Z(n1787) );
  AND U5298 ( .A(b[8]), .B(a[110]), .Z(n1786) );
  XOR U5299 ( .A(n1791), .B(n1608), .Z(n1610) );
  XOR U5300 ( .A(n1792), .B(n1793), .Z(n1608) );
  AND U5301 ( .A(n1794), .B(n1795), .Z(n1792) );
  AND U5302 ( .A(b[7]), .B(a[111]), .Z(n1791) );
  XOR U5303 ( .A(n1796), .B(n1613), .Z(n1615) );
  XOR U5304 ( .A(n1797), .B(n1798), .Z(n1613) );
  AND U5305 ( .A(n1799), .B(n1800), .Z(n1797) );
  AND U5306 ( .A(b[6]), .B(a[112]), .Z(n1796) );
  XOR U5307 ( .A(n1801), .B(n1618), .Z(n1620) );
  XOR U5308 ( .A(n1802), .B(n1803), .Z(n1618) );
  AND U5309 ( .A(n1804), .B(n1805), .Z(n1802) );
  AND U5310 ( .A(b[5]), .B(a[113]), .Z(n1801) );
  XOR U5311 ( .A(n1806), .B(n1623), .Z(n1625) );
  XOR U5312 ( .A(n1807), .B(n1808), .Z(n1623) );
  AND U5313 ( .A(n1809), .B(n1810), .Z(n1807) );
  AND U5314 ( .A(b[4]), .B(a[114]), .Z(n1806) );
  XNOR U5315 ( .A(n1811), .B(n1812), .Z(n1637) );
  NANDN U5316 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U5317 ( .A(n1815), .B(n1628), .Z(n1630) );
  XNOR U5318 ( .A(n1816), .B(n1817), .Z(n1628) );
  AND U5319 ( .A(n1818), .B(n1819), .Z(n1816) );
  AND U5320 ( .A(b[3]), .B(a[115]), .Z(n1815) );
  XOR U5321 ( .A(n1820), .B(n1821), .Z(swire[117]) );
  XOR U5322 ( .A(n1647), .B(n1823), .Z(n1821) );
  XOR U5323 ( .A(n1646), .B(n1822), .Z(n1823) );
  IV U5324 ( .A(n1820), .Z(n1822) );
  NAND U5325 ( .A(a[117]), .B(b[0]), .Z(n1646) );
  XNOR U5326 ( .A(n1813), .B(n1814), .Z(n1647) );
  XOR U5327 ( .A(n1811), .B(n1824), .Z(n1814) );
  NAND U5328 ( .A(b[1]), .B(a[116]), .Z(n1824) );
  XOR U5329 ( .A(n1819), .B(n1825), .Z(n1813) );
  XOR U5330 ( .A(n1811), .B(n1818), .Z(n1825) );
  XNOR U5331 ( .A(n1826), .B(n1817), .Z(n1818) );
  AND U5332 ( .A(b[2]), .B(a[115]), .Z(n1826) );
  NANDN U5333 ( .A(n1827), .B(n1828), .Z(n1811) );
  XOR U5334 ( .A(n1817), .B(n1809), .Z(n1829) );
  XNOR U5335 ( .A(n1808), .B(n1804), .Z(n1830) );
  XNOR U5336 ( .A(n1803), .B(n1799), .Z(n1831) );
  XNOR U5337 ( .A(n1798), .B(n1794), .Z(n1832) );
  XNOR U5338 ( .A(n1793), .B(n1789), .Z(n1833) );
  XNOR U5339 ( .A(n1788), .B(n1784), .Z(n1834) );
  XNOR U5340 ( .A(n1783), .B(n1779), .Z(n1835) );
  XNOR U5341 ( .A(n1778), .B(n1774), .Z(n1836) );
  XNOR U5342 ( .A(n1773), .B(n1769), .Z(n1837) );
  XNOR U5343 ( .A(n1768), .B(n1764), .Z(n1838) );
  XNOR U5344 ( .A(n1763), .B(n1759), .Z(n1839) );
  XNOR U5345 ( .A(n1758), .B(n1754), .Z(n1840) );
  XNOR U5346 ( .A(n1753), .B(n1749), .Z(n1841) );
  XNOR U5347 ( .A(n1748), .B(n1744), .Z(n1842) );
  XNOR U5348 ( .A(n1743), .B(n1739), .Z(n1843) );
  XNOR U5349 ( .A(n1738), .B(n1734), .Z(n1844) );
  XNOR U5350 ( .A(n1733), .B(n1729), .Z(n1845) );
  XNOR U5351 ( .A(n1728), .B(n1724), .Z(n1846) );
  XNOR U5352 ( .A(n1723), .B(n1719), .Z(n1847) );
  XNOR U5353 ( .A(n1718), .B(n1714), .Z(n1848) );
  XNOR U5354 ( .A(n1713), .B(n1709), .Z(n1849) );
  XNOR U5355 ( .A(n1708), .B(n1704), .Z(n1850) );
  XNOR U5356 ( .A(n1703), .B(n1699), .Z(n1851) );
  XNOR U5357 ( .A(n1698), .B(n1694), .Z(n1852) );
  XNOR U5358 ( .A(n1693), .B(n1689), .Z(n1853) );
  XOR U5359 ( .A(n1688), .B(n1685), .Z(n1854) );
  XOR U5360 ( .A(n1855), .B(n1856), .Z(n1685) );
  XOR U5361 ( .A(n1683), .B(n1857), .Z(n1856) );
  XOR U5362 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U5363 ( .A(n1860), .B(n1861), .Z(n1859) );
  NAND U5364 ( .A(a[87]), .B(b[30]), .Z(n1861) );
  AND U5365 ( .A(a[86]), .B(b[31]), .Z(n1860) );
  XOR U5366 ( .A(n1862), .B(n1858), .Z(n1855) );
  XOR U5367 ( .A(n1863), .B(n1864), .Z(n1858) );
  ANDN U5368 ( .B(n1865), .A(n1866), .Z(n1863) );
  AND U5369 ( .A(a[88]), .B(b[29]), .Z(n1862) );
  XOR U5370 ( .A(n1867), .B(n1683), .Z(n1684) );
  XOR U5371 ( .A(n1868), .B(n1869), .Z(n1683) );
  AND U5372 ( .A(n1870), .B(n1871), .Z(n1868) );
  AND U5373 ( .A(a[89]), .B(b[28]), .Z(n1867) );
  XOR U5374 ( .A(n1872), .B(n1688), .Z(n1690) );
  XOR U5375 ( .A(n1873), .B(n1874), .Z(n1688) );
  AND U5376 ( .A(n1875), .B(n1876), .Z(n1873) );
  AND U5377 ( .A(a[90]), .B(b[27]), .Z(n1872) );
  XOR U5378 ( .A(n1877), .B(n1693), .Z(n1695) );
  XOR U5379 ( .A(n1878), .B(n1879), .Z(n1693) );
  AND U5380 ( .A(n1880), .B(n1881), .Z(n1878) );
  AND U5381 ( .A(a[91]), .B(b[26]), .Z(n1877) );
  XOR U5382 ( .A(n1882), .B(n1698), .Z(n1700) );
  XOR U5383 ( .A(n1883), .B(n1884), .Z(n1698) );
  AND U5384 ( .A(n1885), .B(n1886), .Z(n1883) );
  AND U5385 ( .A(a[92]), .B(b[25]), .Z(n1882) );
  XOR U5386 ( .A(n1887), .B(n1703), .Z(n1705) );
  XOR U5387 ( .A(n1888), .B(n1889), .Z(n1703) );
  AND U5388 ( .A(n1890), .B(n1891), .Z(n1888) );
  AND U5389 ( .A(a[93]), .B(b[24]), .Z(n1887) );
  XOR U5390 ( .A(n1892), .B(n1708), .Z(n1710) );
  XOR U5391 ( .A(n1893), .B(n1894), .Z(n1708) );
  AND U5392 ( .A(n1895), .B(n1896), .Z(n1893) );
  AND U5393 ( .A(a[94]), .B(b[23]), .Z(n1892) );
  XOR U5394 ( .A(n1897), .B(n1713), .Z(n1715) );
  XOR U5395 ( .A(n1898), .B(n1899), .Z(n1713) );
  AND U5396 ( .A(n1900), .B(n1901), .Z(n1898) );
  AND U5397 ( .A(b[22]), .B(a[95]), .Z(n1897) );
  XOR U5398 ( .A(n1902), .B(n1718), .Z(n1720) );
  XOR U5399 ( .A(n1903), .B(n1904), .Z(n1718) );
  AND U5400 ( .A(n1905), .B(n1906), .Z(n1903) );
  AND U5401 ( .A(b[21]), .B(a[96]), .Z(n1902) );
  XOR U5402 ( .A(n1907), .B(n1723), .Z(n1725) );
  XOR U5403 ( .A(n1908), .B(n1909), .Z(n1723) );
  AND U5404 ( .A(n1910), .B(n1911), .Z(n1908) );
  AND U5405 ( .A(b[20]), .B(a[97]), .Z(n1907) );
  XOR U5406 ( .A(n1912), .B(n1728), .Z(n1730) );
  XOR U5407 ( .A(n1913), .B(n1914), .Z(n1728) );
  AND U5408 ( .A(n1915), .B(n1916), .Z(n1913) );
  AND U5409 ( .A(b[19]), .B(a[98]), .Z(n1912) );
  XOR U5410 ( .A(n1917), .B(n1733), .Z(n1735) );
  XOR U5411 ( .A(n1918), .B(n1919), .Z(n1733) );
  AND U5412 ( .A(n1920), .B(n1921), .Z(n1918) );
  AND U5413 ( .A(b[18]), .B(a[99]), .Z(n1917) );
  XOR U5414 ( .A(n1922), .B(n1738), .Z(n1740) );
  XOR U5415 ( .A(n1923), .B(n1924), .Z(n1738) );
  AND U5416 ( .A(n1925), .B(n1926), .Z(n1923) );
  AND U5417 ( .A(b[17]), .B(a[100]), .Z(n1922) );
  XOR U5418 ( .A(n1927), .B(n1743), .Z(n1745) );
  XOR U5419 ( .A(n1928), .B(n1929), .Z(n1743) );
  AND U5420 ( .A(n1930), .B(n1931), .Z(n1928) );
  AND U5421 ( .A(b[16]), .B(a[101]), .Z(n1927) );
  XOR U5422 ( .A(n1932), .B(n1748), .Z(n1750) );
  XOR U5423 ( .A(n1933), .B(n1934), .Z(n1748) );
  AND U5424 ( .A(n1935), .B(n1936), .Z(n1933) );
  AND U5425 ( .A(b[15]), .B(a[102]), .Z(n1932) );
  XOR U5426 ( .A(n1937), .B(n1753), .Z(n1755) );
  XOR U5427 ( .A(n1938), .B(n1939), .Z(n1753) );
  AND U5428 ( .A(n1940), .B(n1941), .Z(n1938) );
  AND U5429 ( .A(b[14]), .B(a[103]), .Z(n1937) );
  XOR U5430 ( .A(n1942), .B(n1758), .Z(n1760) );
  XOR U5431 ( .A(n1943), .B(n1944), .Z(n1758) );
  AND U5432 ( .A(n1945), .B(n1946), .Z(n1943) );
  AND U5433 ( .A(b[13]), .B(a[104]), .Z(n1942) );
  XOR U5434 ( .A(n1947), .B(n1763), .Z(n1765) );
  XOR U5435 ( .A(n1948), .B(n1949), .Z(n1763) );
  AND U5436 ( .A(n1950), .B(n1951), .Z(n1948) );
  AND U5437 ( .A(b[12]), .B(a[105]), .Z(n1947) );
  XOR U5438 ( .A(n1952), .B(n1768), .Z(n1770) );
  XOR U5439 ( .A(n1953), .B(n1954), .Z(n1768) );
  AND U5440 ( .A(n1955), .B(n1956), .Z(n1953) );
  AND U5441 ( .A(b[11]), .B(a[106]), .Z(n1952) );
  XOR U5442 ( .A(n1957), .B(n1773), .Z(n1775) );
  XOR U5443 ( .A(n1958), .B(n1959), .Z(n1773) );
  AND U5444 ( .A(n1960), .B(n1961), .Z(n1958) );
  AND U5445 ( .A(b[10]), .B(a[107]), .Z(n1957) );
  XOR U5446 ( .A(n1962), .B(n1778), .Z(n1780) );
  XOR U5447 ( .A(n1963), .B(n1964), .Z(n1778) );
  AND U5448 ( .A(n1965), .B(n1966), .Z(n1963) );
  AND U5449 ( .A(b[9]), .B(a[108]), .Z(n1962) );
  XOR U5450 ( .A(n1967), .B(n1783), .Z(n1785) );
  XOR U5451 ( .A(n1968), .B(n1969), .Z(n1783) );
  AND U5452 ( .A(n1970), .B(n1971), .Z(n1968) );
  AND U5453 ( .A(b[8]), .B(a[109]), .Z(n1967) );
  XOR U5454 ( .A(n1972), .B(n1788), .Z(n1790) );
  XOR U5455 ( .A(n1973), .B(n1974), .Z(n1788) );
  AND U5456 ( .A(n1975), .B(n1976), .Z(n1973) );
  AND U5457 ( .A(b[7]), .B(a[110]), .Z(n1972) );
  XOR U5458 ( .A(n1977), .B(n1793), .Z(n1795) );
  XOR U5459 ( .A(n1978), .B(n1979), .Z(n1793) );
  AND U5460 ( .A(n1980), .B(n1981), .Z(n1978) );
  AND U5461 ( .A(b[6]), .B(a[111]), .Z(n1977) );
  XOR U5462 ( .A(n1982), .B(n1798), .Z(n1800) );
  XOR U5463 ( .A(n1983), .B(n1984), .Z(n1798) );
  AND U5464 ( .A(n1985), .B(n1986), .Z(n1983) );
  AND U5465 ( .A(b[5]), .B(a[112]), .Z(n1982) );
  XOR U5466 ( .A(n1987), .B(n1803), .Z(n1805) );
  XOR U5467 ( .A(n1988), .B(n1989), .Z(n1803) );
  AND U5468 ( .A(n1990), .B(n1991), .Z(n1988) );
  AND U5469 ( .A(b[4]), .B(a[113]), .Z(n1987) );
  XNOR U5470 ( .A(n1992), .B(n1993), .Z(n1817) );
  NANDN U5471 ( .A(n1994), .B(n1995), .Z(n1993) );
  XOR U5472 ( .A(n1996), .B(n1808), .Z(n1810) );
  XNOR U5473 ( .A(n1997), .B(n1998), .Z(n1808) );
  AND U5474 ( .A(n1999), .B(n2000), .Z(n1997) );
  AND U5475 ( .A(b[3]), .B(a[114]), .Z(n1996) );
  XNOR U5476 ( .A(n2001), .B(n2002), .Z(swire[116]) );
  XOR U5477 ( .A(n1828), .B(n2003), .Z(n2002) );
  XOR U5478 ( .A(n1827), .B(n2001), .Z(n2003) );
  NAND U5479 ( .A(a[116]), .B(b[0]), .Z(n1827) );
  XNOR U5480 ( .A(n1994), .B(n1995), .Z(n1828) );
  XOR U5481 ( .A(n1992), .B(n2004), .Z(n1995) );
  NAND U5482 ( .A(b[1]), .B(a[115]), .Z(n2004) );
  XOR U5483 ( .A(n2000), .B(n2005), .Z(n1994) );
  XOR U5484 ( .A(n1992), .B(n1999), .Z(n2005) );
  XNOR U5485 ( .A(n2006), .B(n1998), .Z(n1999) );
  AND U5486 ( .A(b[2]), .B(a[114]), .Z(n2006) );
  NANDN U5487 ( .A(n2007), .B(n2008), .Z(n1992) );
  XOR U5488 ( .A(n1998), .B(n1990), .Z(n2009) );
  XNOR U5489 ( .A(n1989), .B(n1985), .Z(n2010) );
  XNOR U5490 ( .A(n1984), .B(n1980), .Z(n2011) );
  XNOR U5491 ( .A(n1979), .B(n1975), .Z(n2012) );
  XNOR U5492 ( .A(n1974), .B(n1970), .Z(n2013) );
  XNOR U5493 ( .A(n1969), .B(n1965), .Z(n2014) );
  XNOR U5494 ( .A(n1964), .B(n1960), .Z(n2015) );
  XNOR U5495 ( .A(n1959), .B(n1955), .Z(n2016) );
  XNOR U5496 ( .A(n1954), .B(n1950), .Z(n2017) );
  XNOR U5497 ( .A(n1949), .B(n1945), .Z(n2018) );
  XNOR U5498 ( .A(n1944), .B(n1940), .Z(n2019) );
  XNOR U5499 ( .A(n1939), .B(n1935), .Z(n2020) );
  XNOR U5500 ( .A(n1934), .B(n1930), .Z(n2021) );
  XNOR U5501 ( .A(n1929), .B(n1925), .Z(n2022) );
  XNOR U5502 ( .A(n1924), .B(n1920), .Z(n2023) );
  XNOR U5503 ( .A(n1919), .B(n1915), .Z(n2024) );
  XNOR U5504 ( .A(n1914), .B(n1910), .Z(n2025) );
  XNOR U5505 ( .A(n1909), .B(n1905), .Z(n2026) );
  XNOR U5506 ( .A(n1904), .B(n1900), .Z(n2027) );
  XNOR U5507 ( .A(n1899), .B(n1895), .Z(n2028) );
  XNOR U5508 ( .A(n1894), .B(n1890), .Z(n2029) );
  XNOR U5509 ( .A(n1889), .B(n1885), .Z(n2030) );
  XNOR U5510 ( .A(n1884), .B(n1880), .Z(n2031) );
  XNOR U5511 ( .A(n1879), .B(n1875), .Z(n2032) );
  XNOR U5512 ( .A(n1874), .B(n1870), .Z(n2033) );
  XOR U5513 ( .A(n1869), .B(n1866), .Z(n2034) );
  XOR U5514 ( .A(n2035), .B(n2036), .Z(n1866) );
  XOR U5515 ( .A(n1864), .B(n2037), .Z(n2036) );
  XOR U5516 ( .A(n2038), .B(n2039), .Z(n2037) );
  XOR U5517 ( .A(n2040), .B(n2041), .Z(n2039) );
  NAND U5518 ( .A(a[86]), .B(b[30]), .Z(n2041) );
  AND U5519 ( .A(a[85]), .B(b[31]), .Z(n2040) );
  XOR U5520 ( .A(n2042), .B(n2038), .Z(n2035) );
  XOR U5521 ( .A(n2043), .B(n2044), .Z(n2038) );
  ANDN U5522 ( .B(n2045), .A(n2046), .Z(n2043) );
  AND U5523 ( .A(a[87]), .B(b[29]), .Z(n2042) );
  XOR U5524 ( .A(n2047), .B(n1864), .Z(n1865) );
  XOR U5525 ( .A(n2048), .B(n2049), .Z(n1864) );
  AND U5526 ( .A(n2050), .B(n2051), .Z(n2048) );
  AND U5527 ( .A(a[88]), .B(b[28]), .Z(n2047) );
  XOR U5528 ( .A(n2052), .B(n1869), .Z(n1871) );
  XOR U5529 ( .A(n2053), .B(n2054), .Z(n1869) );
  AND U5530 ( .A(n2055), .B(n2056), .Z(n2053) );
  AND U5531 ( .A(a[89]), .B(b[27]), .Z(n2052) );
  XOR U5532 ( .A(n2057), .B(n1874), .Z(n1876) );
  XOR U5533 ( .A(n2058), .B(n2059), .Z(n1874) );
  AND U5534 ( .A(n2060), .B(n2061), .Z(n2058) );
  AND U5535 ( .A(a[90]), .B(b[26]), .Z(n2057) );
  XOR U5536 ( .A(n2062), .B(n1879), .Z(n1881) );
  XOR U5537 ( .A(n2063), .B(n2064), .Z(n1879) );
  AND U5538 ( .A(n2065), .B(n2066), .Z(n2063) );
  AND U5539 ( .A(a[91]), .B(b[25]), .Z(n2062) );
  XOR U5540 ( .A(n2067), .B(n1884), .Z(n1886) );
  XOR U5541 ( .A(n2068), .B(n2069), .Z(n1884) );
  AND U5542 ( .A(n2070), .B(n2071), .Z(n2068) );
  AND U5543 ( .A(a[92]), .B(b[24]), .Z(n2067) );
  XOR U5544 ( .A(n2072), .B(n1889), .Z(n1891) );
  XOR U5545 ( .A(n2073), .B(n2074), .Z(n1889) );
  AND U5546 ( .A(n2075), .B(n2076), .Z(n2073) );
  AND U5547 ( .A(a[93]), .B(b[23]), .Z(n2072) );
  XOR U5548 ( .A(n2077), .B(n1894), .Z(n1896) );
  XOR U5549 ( .A(n2078), .B(n2079), .Z(n1894) );
  AND U5550 ( .A(n2080), .B(n2081), .Z(n2078) );
  AND U5551 ( .A(a[94]), .B(b[22]), .Z(n2077) );
  XOR U5552 ( .A(n2082), .B(n1899), .Z(n1901) );
  XOR U5553 ( .A(n2083), .B(n2084), .Z(n1899) );
  AND U5554 ( .A(n2085), .B(n2086), .Z(n2083) );
  AND U5555 ( .A(b[21]), .B(a[95]), .Z(n2082) );
  XOR U5556 ( .A(n2087), .B(n1904), .Z(n1906) );
  XOR U5557 ( .A(n2088), .B(n2089), .Z(n1904) );
  AND U5558 ( .A(n2090), .B(n2091), .Z(n2088) );
  AND U5559 ( .A(b[20]), .B(a[96]), .Z(n2087) );
  XOR U5560 ( .A(n2092), .B(n1909), .Z(n1911) );
  XOR U5561 ( .A(n2093), .B(n2094), .Z(n1909) );
  AND U5562 ( .A(n2095), .B(n2096), .Z(n2093) );
  AND U5563 ( .A(b[19]), .B(a[97]), .Z(n2092) );
  XOR U5564 ( .A(n2097), .B(n1914), .Z(n1916) );
  XOR U5565 ( .A(n2098), .B(n2099), .Z(n1914) );
  AND U5566 ( .A(n2100), .B(n2101), .Z(n2098) );
  AND U5567 ( .A(b[18]), .B(a[98]), .Z(n2097) );
  XOR U5568 ( .A(n2102), .B(n1919), .Z(n1921) );
  XOR U5569 ( .A(n2103), .B(n2104), .Z(n1919) );
  AND U5570 ( .A(n2105), .B(n2106), .Z(n2103) );
  AND U5571 ( .A(b[17]), .B(a[99]), .Z(n2102) );
  XOR U5572 ( .A(n2107), .B(n1924), .Z(n1926) );
  XOR U5573 ( .A(n2108), .B(n2109), .Z(n1924) );
  AND U5574 ( .A(n2110), .B(n2111), .Z(n2108) );
  AND U5575 ( .A(b[16]), .B(a[100]), .Z(n2107) );
  XOR U5576 ( .A(n2112), .B(n1929), .Z(n1931) );
  XOR U5577 ( .A(n2113), .B(n2114), .Z(n1929) );
  AND U5578 ( .A(n2115), .B(n2116), .Z(n2113) );
  AND U5579 ( .A(b[15]), .B(a[101]), .Z(n2112) );
  XOR U5580 ( .A(n2117), .B(n1934), .Z(n1936) );
  XOR U5581 ( .A(n2118), .B(n2119), .Z(n1934) );
  AND U5582 ( .A(n2120), .B(n2121), .Z(n2118) );
  AND U5583 ( .A(b[14]), .B(a[102]), .Z(n2117) );
  XOR U5584 ( .A(n2122), .B(n1939), .Z(n1941) );
  XOR U5585 ( .A(n2123), .B(n2124), .Z(n1939) );
  AND U5586 ( .A(n2125), .B(n2126), .Z(n2123) );
  AND U5587 ( .A(b[13]), .B(a[103]), .Z(n2122) );
  XOR U5588 ( .A(n2127), .B(n1944), .Z(n1946) );
  XOR U5589 ( .A(n2128), .B(n2129), .Z(n1944) );
  AND U5590 ( .A(n2130), .B(n2131), .Z(n2128) );
  AND U5591 ( .A(b[12]), .B(a[104]), .Z(n2127) );
  XOR U5592 ( .A(n2132), .B(n1949), .Z(n1951) );
  XOR U5593 ( .A(n2133), .B(n2134), .Z(n1949) );
  AND U5594 ( .A(n2135), .B(n2136), .Z(n2133) );
  AND U5595 ( .A(b[11]), .B(a[105]), .Z(n2132) );
  XOR U5596 ( .A(n2137), .B(n1954), .Z(n1956) );
  XOR U5597 ( .A(n2138), .B(n2139), .Z(n1954) );
  AND U5598 ( .A(n2140), .B(n2141), .Z(n2138) );
  AND U5599 ( .A(b[10]), .B(a[106]), .Z(n2137) );
  XOR U5600 ( .A(n2142), .B(n1959), .Z(n1961) );
  XOR U5601 ( .A(n2143), .B(n2144), .Z(n1959) );
  AND U5602 ( .A(n2145), .B(n2146), .Z(n2143) );
  AND U5603 ( .A(b[9]), .B(a[107]), .Z(n2142) );
  XOR U5604 ( .A(n2147), .B(n1964), .Z(n1966) );
  XOR U5605 ( .A(n2148), .B(n2149), .Z(n1964) );
  AND U5606 ( .A(n2150), .B(n2151), .Z(n2148) );
  AND U5607 ( .A(b[8]), .B(a[108]), .Z(n2147) );
  XOR U5608 ( .A(n2152), .B(n1969), .Z(n1971) );
  XOR U5609 ( .A(n2153), .B(n2154), .Z(n1969) );
  AND U5610 ( .A(n2155), .B(n2156), .Z(n2153) );
  AND U5611 ( .A(b[7]), .B(a[109]), .Z(n2152) );
  XOR U5612 ( .A(n2157), .B(n1974), .Z(n1976) );
  XOR U5613 ( .A(n2158), .B(n2159), .Z(n1974) );
  AND U5614 ( .A(n2160), .B(n2161), .Z(n2158) );
  AND U5615 ( .A(b[6]), .B(a[110]), .Z(n2157) );
  XOR U5616 ( .A(n2162), .B(n1979), .Z(n1981) );
  XOR U5617 ( .A(n2163), .B(n2164), .Z(n1979) );
  AND U5618 ( .A(n2165), .B(n2166), .Z(n2163) );
  AND U5619 ( .A(b[5]), .B(a[111]), .Z(n2162) );
  XOR U5620 ( .A(n2167), .B(n1984), .Z(n1986) );
  XOR U5621 ( .A(n2168), .B(n2169), .Z(n1984) );
  AND U5622 ( .A(n2170), .B(n2171), .Z(n2168) );
  AND U5623 ( .A(b[4]), .B(a[112]), .Z(n2167) );
  XNOR U5624 ( .A(n2172), .B(n2173), .Z(n1998) );
  NANDN U5625 ( .A(n2174), .B(n2175), .Z(n2173) );
  XOR U5626 ( .A(n2176), .B(n1989), .Z(n1991) );
  XNOR U5627 ( .A(n2177), .B(n2178), .Z(n1989) );
  AND U5628 ( .A(n2179), .B(n2180), .Z(n2177) );
  AND U5629 ( .A(b[3]), .B(a[113]), .Z(n2176) );
  XOR U5630 ( .A(n2181), .B(n2182), .Z(swire[115]) );
  XOR U5631 ( .A(n2008), .B(n2184), .Z(n2182) );
  XOR U5632 ( .A(n2007), .B(n2183), .Z(n2184) );
  IV U5633 ( .A(n2181), .Z(n2183) );
  NAND U5634 ( .A(a[115]), .B(b[0]), .Z(n2007) );
  XNOR U5635 ( .A(n2174), .B(n2175), .Z(n2008) );
  XOR U5636 ( .A(n2172), .B(n2185), .Z(n2175) );
  NAND U5637 ( .A(b[1]), .B(a[114]), .Z(n2185) );
  XOR U5638 ( .A(n2180), .B(n2186), .Z(n2174) );
  XOR U5639 ( .A(n2172), .B(n2179), .Z(n2186) );
  XNOR U5640 ( .A(n2187), .B(n2178), .Z(n2179) );
  AND U5641 ( .A(b[2]), .B(a[113]), .Z(n2187) );
  NANDN U5642 ( .A(n2188), .B(n2189), .Z(n2172) );
  XOR U5643 ( .A(n2178), .B(n2170), .Z(n2190) );
  XNOR U5644 ( .A(n2169), .B(n2165), .Z(n2191) );
  XNOR U5645 ( .A(n2164), .B(n2160), .Z(n2192) );
  XNOR U5646 ( .A(n2159), .B(n2155), .Z(n2193) );
  XNOR U5647 ( .A(n2154), .B(n2150), .Z(n2194) );
  XNOR U5648 ( .A(n2149), .B(n2145), .Z(n2195) );
  XNOR U5649 ( .A(n2144), .B(n2140), .Z(n2196) );
  XNOR U5650 ( .A(n2139), .B(n2135), .Z(n2197) );
  XNOR U5651 ( .A(n2134), .B(n2130), .Z(n2198) );
  XNOR U5652 ( .A(n2129), .B(n2125), .Z(n2199) );
  XNOR U5653 ( .A(n2124), .B(n2120), .Z(n2200) );
  XNOR U5654 ( .A(n2119), .B(n2115), .Z(n2201) );
  XNOR U5655 ( .A(n2114), .B(n2110), .Z(n2202) );
  XNOR U5656 ( .A(n2109), .B(n2105), .Z(n2203) );
  XNOR U5657 ( .A(n2104), .B(n2100), .Z(n2204) );
  XNOR U5658 ( .A(n2099), .B(n2095), .Z(n2205) );
  XNOR U5659 ( .A(n2094), .B(n2090), .Z(n2206) );
  XNOR U5660 ( .A(n2089), .B(n2085), .Z(n2207) );
  XNOR U5661 ( .A(n2084), .B(n2080), .Z(n2208) );
  XNOR U5662 ( .A(n2079), .B(n2075), .Z(n2209) );
  XNOR U5663 ( .A(n2074), .B(n2070), .Z(n2210) );
  XNOR U5664 ( .A(n2069), .B(n2065), .Z(n2211) );
  XNOR U5665 ( .A(n2064), .B(n2060), .Z(n2212) );
  XNOR U5666 ( .A(n2059), .B(n2055), .Z(n2213) );
  XNOR U5667 ( .A(n2054), .B(n2050), .Z(n2214) );
  XOR U5668 ( .A(n2049), .B(n2046), .Z(n2215) );
  XOR U5669 ( .A(n2216), .B(n2217), .Z(n2046) );
  XOR U5670 ( .A(n2044), .B(n2218), .Z(n2217) );
  XOR U5671 ( .A(n2219), .B(n2220), .Z(n2218) );
  XOR U5672 ( .A(n2221), .B(n2222), .Z(n2220) );
  NAND U5673 ( .A(a[85]), .B(b[30]), .Z(n2222) );
  AND U5674 ( .A(a[84]), .B(b[31]), .Z(n2221) );
  XOR U5675 ( .A(n2223), .B(n2219), .Z(n2216) );
  XOR U5676 ( .A(n2224), .B(n2225), .Z(n2219) );
  ANDN U5677 ( .B(n2226), .A(n2227), .Z(n2224) );
  AND U5678 ( .A(a[86]), .B(b[29]), .Z(n2223) );
  XOR U5679 ( .A(n2228), .B(n2044), .Z(n2045) );
  XOR U5680 ( .A(n2229), .B(n2230), .Z(n2044) );
  AND U5681 ( .A(n2231), .B(n2232), .Z(n2229) );
  AND U5682 ( .A(a[87]), .B(b[28]), .Z(n2228) );
  XOR U5683 ( .A(n2233), .B(n2049), .Z(n2051) );
  XOR U5684 ( .A(n2234), .B(n2235), .Z(n2049) );
  AND U5685 ( .A(n2236), .B(n2237), .Z(n2234) );
  AND U5686 ( .A(a[88]), .B(b[27]), .Z(n2233) );
  XOR U5687 ( .A(n2238), .B(n2054), .Z(n2056) );
  XOR U5688 ( .A(n2239), .B(n2240), .Z(n2054) );
  AND U5689 ( .A(n2241), .B(n2242), .Z(n2239) );
  AND U5690 ( .A(a[89]), .B(b[26]), .Z(n2238) );
  XOR U5691 ( .A(n2243), .B(n2059), .Z(n2061) );
  XOR U5692 ( .A(n2244), .B(n2245), .Z(n2059) );
  AND U5693 ( .A(n2246), .B(n2247), .Z(n2244) );
  AND U5694 ( .A(a[90]), .B(b[25]), .Z(n2243) );
  XOR U5695 ( .A(n2248), .B(n2064), .Z(n2066) );
  XOR U5696 ( .A(n2249), .B(n2250), .Z(n2064) );
  AND U5697 ( .A(n2251), .B(n2252), .Z(n2249) );
  AND U5698 ( .A(a[91]), .B(b[24]), .Z(n2248) );
  XOR U5699 ( .A(n2253), .B(n2069), .Z(n2071) );
  XOR U5700 ( .A(n2254), .B(n2255), .Z(n2069) );
  AND U5701 ( .A(n2256), .B(n2257), .Z(n2254) );
  AND U5702 ( .A(a[92]), .B(b[23]), .Z(n2253) );
  XOR U5703 ( .A(n2258), .B(n2074), .Z(n2076) );
  XOR U5704 ( .A(n2259), .B(n2260), .Z(n2074) );
  AND U5705 ( .A(n2261), .B(n2262), .Z(n2259) );
  AND U5706 ( .A(a[93]), .B(b[22]), .Z(n2258) );
  XOR U5707 ( .A(n2263), .B(n2079), .Z(n2081) );
  XOR U5708 ( .A(n2264), .B(n2265), .Z(n2079) );
  AND U5709 ( .A(n2266), .B(n2267), .Z(n2264) );
  AND U5710 ( .A(a[94]), .B(b[21]), .Z(n2263) );
  XOR U5711 ( .A(n2268), .B(n2084), .Z(n2086) );
  XOR U5712 ( .A(n2269), .B(n2270), .Z(n2084) );
  AND U5713 ( .A(n2271), .B(n2272), .Z(n2269) );
  AND U5714 ( .A(b[20]), .B(a[95]), .Z(n2268) );
  XOR U5715 ( .A(n2273), .B(n2089), .Z(n2091) );
  XOR U5716 ( .A(n2274), .B(n2275), .Z(n2089) );
  AND U5717 ( .A(n2276), .B(n2277), .Z(n2274) );
  AND U5718 ( .A(b[19]), .B(a[96]), .Z(n2273) );
  XOR U5719 ( .A(n2278), .B(n2094), .Z(n2096) );
  XOR U5720 ( .A(n2279), .B(n2280), .Z(n2094) );
  AND U5721 ( .A(n2281), .B(n2282), .Z(n2279) );
  AND U5722 ( .A(b[18]), .B(a[97]), .Z(n2278) );
  XOR U5723 ( .A(n2283), .B(n2099), .Z(n2101) );
  XOR U5724 ( .A(n2284), .B(n2285), .Z(n2099) );
  AND U5725 ( .A(n2286), .B(n2287), .Z(n2284) );
  AND U5726 ( .A(b[17]), .B(a[98]), .Z(n2283) );
  XOR U5727 ( .A(n2288), .B(n2104), .Z(n2106) );
  XOR U5728 ( .A(n2289), .B(n2290), .Z(n2104) );
  AND U5729 ( .A(n2291), .B(n2292), .Z(n2289) );
  AND U5730 ( .A(b[16]), .B(a[99]), .Z(n2288) );
  XOR U5731 ( .A(n2293), .B(n2109), .Z(n2111) );
  XOR U5732 ( .A(n2294), .B(n2295), .Z(n2109) );
  AND U5733 ( .A(n2296), .B(n2297), .Z(n2294) );
  AND U5734 ( .A(b[15]), .B(a[100]), .Z(n2293) );
  XOR U5735 ( .A(n2298), .B(n2114), .Z(n2116) );
  XOR U5736 ( .A(n2299), .B(n2300), .Z(n2114) );
  AND U5737 ( .A(n2301), .B(n2302), .Z(n2299) );
  AND U5738 ( .A(b[14]), .B(a[101]), .Z(n2298) );
  XOR U5739 ( .A(n2303), .B(n2119), .Z(n2121) );
  XOR U5740 ( .A(n2304), .B(n2305), .Z(n2119) );
  AND U5741 ( .A(n2306), .B(n2307), .Z(n2304) );
  AND U5742 ( .A(b[13]), .B(a[102]), .Z(n2303) );
  XOR U5743 ( .A(n2308), .B(n2124), .Z(n2126) );
  XOR U5744 ( .A(n2309), .B(n2310), .Z(n2124) );
  AND U5745 ( .A(n2311), .B(n2312), .Z(n2309) );
  AND U5746 ( .A(b[12]), .B(a[103]), .Z(n2308) );
  XOR U5747 ( .A(n2313), .B(n2129), .Z(n2131) );
  XOR U5748 ( .A(n2314), .B(n2315), .Z(n2129) );
  AND U5749 ( .A(n2316), .B(n2317), .Z(n2314) );
  AND U5750 ( .A(b[11]), .B(a[104]), .Z(n2313) );
  XOR U5751 ( .A(n2318), .B(n2134), .Z(n2136) );
  XOR U5752 ( .A(n2319), .B(n2320), .Z(n2134) );
  AND U5753 ( .A(n2321), .B(n2322), .Z(n2319) );
  AND U5754 ( .A(b[10]), .B(a[105]), .Z(n2318) );
  XOR U5755 ( .A(n2323), .B(n2139), .Z(n2141) );
  XOR U5756 ( .A(n2324), .B(n2325), .Z(n2139) );
  AND U5757 ( .A(n2326), .B(n2327), .Z(n2324) );
  AND U5758 ( .A(b[9]), .B(a[106]), .Z(n2323) );
  XOR U5759 ( .A(n2328), .B(n2144), .Z(n2146) );
  XOR U5760 ( .A(n2329), .B(n2330), .Z(n2144) );
  AND U5761 ( .A(n2331), .B(n2332), .Z(n2329) );
  AND U5762 ( .A(b[8]), .B(a[107]), .Z(n2328) );
  XOR U5763 ( .A(n2333), .B(n2149), .Z(n2151) );
  XOR U5764 ( .A(n2334), .B(n2335), .Z(n2149) );
  AND U5765 ( .A(n2336), .B(n2337), .Z(n2334) );
  AND U5766 ( .A(b[7]), .B(a[108]), .Z(n2333) );
  XOR U5767 ( .A(n2338), .B(n2154), .Z(n2156) );
  XOR U5768 ( .A(n2339), .B(n2340), .Z(n2154) );
  AND U5769 ( .A(n2341), .B(n2342), .Z(n2339) );
  AND U5770 ( .A(b[6]), .B(a[109]), .Z(n2338) );
  XOR U5771 ( .A(n2343), .B(n2159), .Z(n2161) );
  XOR U5772 ( .A(n2344), .B(n2345), .Z(n2159) );
  AND U5773 ( .A(n2346), .B(n2347), .Z(n2344) );
  AND U5774 ( .A(b[5]), .B(a[110]), .Z(n2343) );
  XOR U5775 ( .A(n2348), .B(n2164), .Z(n2166) );
  XOR U5776 ( .A(n2349), .B(n2350), .Z(n2164) );
  AND U5777 ( .A(n2351), .B(n2352), .Z(n2349) );
  AND U5778 ( .A(b[4]), .B(a[111]), .Z(n2348) );
  XNOR U5779 ( .A(n2353), .B(n2354), .Z(n2178) );
  NANDN U5780 ( .A(n2355), .B(n2356), .Z(n2354) );
  XOR U5781 ( .A(n2357), .B(n2169), .Z(n2171) );
  XNOR U5782 ( .A(n2358), .B(n2359), .Z(n2169) );
  AND U5783 ( .A(n2360), .B(n2361), .Z(n2358) );
  AND U5784 ( .A(b[3]), .B(a[112]), .Z(n2357) );
  XNOR U5785 ( .A(n2362), .B(n2363), .Z(swire[114]) );
  XOR U5786 ( .A(n2189), .B(n2364), .Z(n2363) );
  XOR U5787 ( .A(n2188), .B(n2362), .Z(n2364) );
  NAND U5788 ( .A(a[114]), .B(b[0]), .Z(n2188) );
  XNOR U5789 ( .A(n2355), .B(n2356), .Z(n2189) );
  XOR U5790 ( .A(n2353), .B(n2365), .Z(n2356) );
  NAND U5791 ( .A(b[1]), .B(a[113]), .Z(n2365) );
  XOR U5792 ( .A(n2361), .B(n2366), .Z(n2355) );
  XOR U5793 ( .A(n2353), .B(n2360), .Z(n2366) );
  XNOR U5794 ( .A(n2367), .B(n2359), .Z(n2360) );
  AND U5795 ( .A(b[2]), .B(a[112]), .Z(n2367) );
  NANDN U5796 ( .A(n2368), .B(n2369), .Z(n2353) );
  XOR U5797 ( .A(n2359), .B(n2351), .Z(n2370) );
  XNOR U5798 ( .A(n2350), .B(n2346), .Z(n2371) );
  XNOR U5799 ( .A(n2345), .B(n2341), .Z(n2372) );
  XNOR U5800 ( .A(n2340), .B(n2336), .Z(n2373) );
  XNOR U5801 ( .A(n2335), .B(n2331), .Z(n2374) );
  XNOR U5802 ( .A(n2330), .B(n2326), .Z(n2375) );
  XNOR U5803 ( .A(n2325), .B(n2321), .Z(n2376) );
  XNOR U5804 ( .A(n2320), .B(n2316), .Z(n2377) );
  XNOR U5805 ( .A(n2315), .B(n2311), .Z(n2378) );
  XNOR U5806 ( .A(n2310), .B(n2306), .Z(n2379) );
  XNOR U5807 ( .A(n2305), .B(n2301), .Z(n2380) );
  XNOR U5808 ( .A(n2300), .B(n2296), .Z(n2381) );
  XNOR U5809 ( .A(n2295), .B(n2291), .Z(n2382) );
  XNOR U5810 ( .A(n2290), .B(n2286), .Z(n2383) );
  XNOR U5811 ( .A(n2285), .B(n2281), .Z(n2384) );
  XNOR U5812 ( .A(n2280), .B(n2276), .Z(n2385) );
  XNOR U5813 ( .A(n2275), .B(n2271), .Z(n2386) );
  XNOR U5814 ( .A(n2270), .B(n2266), .Z(n2387) );
  XNOR U5815 ( .A(n2265), .B(n2261), .Z(n2388) );
  XNOR U5816 ( .A(n2260), .B(n2256), .Z(n2389) );
  XNOR U5817 ( .A(n2255), .B(n2251), .Z(n2390) );
  XNOR U5818 ( .A(n2250), .B(n2246), .Z(n2391) );
  XNOR U5819 ( .A(n2245), .B(n2241), .Z(n2392) );
  XNOR U5820 ( .A(n2240), .B(n2236), .Z(n2393) );
  XNOR U5821 ( .A(n2235), .B(n2231), .Z(n2394) );
  XOR U5822 ( .A(n2230), .B(n2227), .Z(n2395) );
  XOR U5823 ( .A(n2396), .B(n2397), .Z(n2227) );
  XOR U5824 ( .A(n2225), .B(n2398), .Z(n2397) );
  XOR U5825 ( .A(n2399), .B(n2400), .Z(n2398) );
  XOR U5826 ( .A(n2401), .B(n2402), .Z(n2400) );
  NAND U5827 ( .A(a[84]), .B(b[30]), .Z(n2402) );
  AND U5828 ( .A(a[83]), .B(b[31]), .Z(n2401) );
  XOR U5829 ( .A(n2403), .B(n2399), .Z(n2396) );
  XOR U5830 ( .A(n2404), .B(n2405), .Z(n2399) );
  ANDN U5831 ( .B(n2406), .A(n2407), .Z(n2404) );
  AND U5832 ( .A(a[85]), .B(b[29]), .Z(n2403) );
  XOR U5833 ( .A(n2408), .B(n2225), .Z(n2226) );
  XOR U5834 ( .A(n2409), .B(n2410), .Z(n2225) );
  AND U5835 ( .A(n2411), .B(n2412), .Z(n2409) );
  AND U5836 ( .A(a[86]), .B(b[28]), .Z(n2408) );
  XOR U5837 ( .A(n2413), .B(n2230), .Z(n2232) );
  XOR U5838 ( .A(n2414), .B(n2415), .Z(n2230) );
  AND U5839 ( .A(n2416), .B(n2417), .Z(n2414) );
  AND U5840 ( .A(a[87]), .B(b[27]), .Z(n2413) );
  XOR U5841 ( .A(n2418), .B(n2235), .Z(n2237) );
  XOR U5842 ( .A(n2419), .B(n2420), .Z(n2235) );
  AND U5843 ( .A(n2421), .B(n2422), .Z(n2419) );
  AND U5844 ( .A(a[88]), .B(b[26]), .Z(n2418) );
  XOR U5845 ( .A(n2423), .B(n2240), .Z(n2242) );
  XOR U5846 ( .A(n2424), .B(n2425), .Z(n2240) );
  AND U5847 ( .A(n2426), .B(n2427), .Z(n2424) );
  AND U5848 ( .A(a[89]), .B(b[25]), .Z(n2423) );
  XOR U5849 ( .A(n2428), .B(n2245), .Z(n2247) );
  XOR U5850 ( .A(n2429), .B(n2430), .Z(n2245) );
  AND U5851 ( .A(n2431), .B(n2432), .Z(n2429) );
  AND U5852 ( .A(a[90]), .B(b[24]), .Z(n2428) );
  XOR U5853 ( .A(n2433), .B(n2250), .Z(n2252) );
  XOR U5854 ( .A(n2434), .B(n2435), .Z(n2250) );
  AND U5855 ( .A(n2436), .B(n2437), .Z(n2434) );
  AND U5856 ( .A(a[91]), .B(b[23]), .Z(n2433) );
  XOR U5857 ( .A(n2438), .B(n2255), .Z(n2257) );
  XOR U5858 ( .A(n2439), .B(n2440), .Z(n2255) );
  AND U5859 ( .A(n2441), .B(n2442), .Z(n2439) );
  AND U5860 ( .A(a[92]), .B(b[22]), .Z(n2438) );
  XOR U5861 ( .A(n2443), .B(n2260), .Z(n2262) );
  XOR U5862 ( .A(n2444), .B(n2445), .Z(n2260) );
  AND U5863 ( .A(n2446), .B(n2447), .Z(n2444) );
  AND U5864 ( .A(a[93]), .B(b[21]), .Z(n2443) );
  XOR U5865 ( .A(n2448), .B(n2265), .Z(n2267) );
  XOR U5866 ( .A(n2449), .B(n2450), .Z(n2265) );
  AND U5867 ( .A(n2451), .B(n2452), .Z(n2449) );
  AND U5868 ( .A(a[94]), .B(b[20]), .Z(n2448) );
  XOR U5869 ( .A(n2453), .B(n2270), .Z(n2272) );
  XOR U5870 ( .A(n2454), .B(n2455), .Z(n2270) );
  AND U5871 ( .A(n2456), .B(n2457), .Z(n2454) );
  AND U5872 ( .A(b[19]), .B(a[95]), .Z(n2453) );
  XOR U5873 ( .A(n2458), .B(n2275), .Z(n2277) );
  XOR U5874 ( .A(n2459), .B(n2460), .Z(n2275) );
  AND U5875 ( .A(n2461), .B(n2462), .Z(n2459) );
  AND U5876 ( .A(b[18]), .B(a[96]), .Z(n2458) );
  XOR U5877 ( .A(n2463), .B(n2280), .Z(n2282) );
  XOR U5878 ( .A(n2464), .B(n2465), .Z(n2280) );
  AND U5879 ( .A(n2466), .B(n2467), .Z(n2464) );
  AND U5880 ( .A(b[17]), .B(a[97]), .Z(n2463) );
  XOR U5881 ( .A(n2468), .B(n2285), .Z(n2287) );
  XOR U5882 ( .A(n2469), .B(n2470), .Z(n2285) );
  AND U5883 ( .A(n2471), .B(n2472), .Z(n2469) );
  AND U5884 ( .A(b[16]), .B(a[98]), .Z(n2468) );
  XOR U5885 ( .A(n2473), .B(n2290), .Z(n2292) );
  XOR U5886 ( .A(n2474), .B(n2475), .Z(n2290) );
  AND U5887 ( .A(n2476), .B(n2477), .Z(n2474) );
  AND U5888 ( .A(b[15]), .B(a[99]), .Z(n2473) );
  XOR U5889 ( .A(n2478), .B(n2295), .Z(n2297) );
  XOR U5890 ( .A(n2479), .B(n2480), .Z(n2295) );
  AND U5891 ( .A(n2481), .B(n2482), .Z(n2479) );
  AND U5892 ( .A(b[14]), .B(a[100]), .Z(n2478) );
  XOR U5893 ( .A(n2483), .B(n2300), .Z(n2302) );
  XOR U5894 ( .A(n2484), .B(n2485), .Z(n2300) );
  AND U5895 ( .A(n2486), .B(n2487), .Z(n2484) );
  AND U5896 ( .A(b[13]), .B(a[101]), .Z(n2483) );
  XOR U5897 ( .A(n2488), .B(n2305), .Z(n2307) );
  XOR U5898 ( .A(n2489), .B(n2490), .Z(n2305) );
  AND U5899 ( .A(n2491), .B(n2492), .Z(n2489) );
  AND U5900 ( .A(b[12]), .B(a[102]), .Z(n2488) );
  XOR U5901 ( .A(n2493), .B(n2310), .Z(n2312) );
  XOR U5902 ( .A(n2494), .B(n2495), .Z(n2310) );
  AND U5903 ( .A(n2496), .B(n2497), .Z(n2494) );
  AND U5904 ( .A(b[11]), .B(a[103]), .Z(n2493) );
  XOR U5905 ( .A(n2498), .B(n2315), .Z(n2317) );
  XOR U5906 ( .A(n2499), .B(n2500), .Z(n2315) );
  AND U5907 ( .A(n2501), .B(n2502), .Z(n2499) );
  AND U5908 ( .A(b[10]), .B(a[104]), .Z(n2498) );
  XOR U5909 ( .A(n2503), .B(n2320), .Z(n2322) );
  XOR U5910 ( .A(n2504), .B(n2505), .Z(n2320) );
  AND U5911 ( .A(n2506), .B(n2507), .Z(n2504) );
  AND U5912 ( .A(b[9]), .B(a[105]), .Z(n2503) );
  XOR U5913 ( .A(n2508), .B(n2325), .Z(n2327) );
  XOR U5914 ( .A(n2509), .B(n2510), .Z(n2325) );
  AND U5915 ( .A(n2511), .B(n2512), .Z(n2509) );
  AND U5916 ( .A(b[8]), .B(a[106]), .Z(n2508) );
  XOR U5917 ( .A(n2513), .B(n2330), .Z(n2332) );
  XOR U5918 ( .A(n2514), .B(n2515), .Z(n2330) );
  AND U5919 ( .A(n2516), .B(n2517), .Z(n2514) );
  AND U5920 ( .A(b[7]), .B(a[107]), .Z(n2513) );
  XOR U5921 ( .A(n2518), .B(n2335), .Z(n2337) );
  XOR U5922 ( .A(n2519), .B(n2520), .Z(n2335) );
  AND U5923 ( .A(n2521), .B(n2522), .Z(n2519) );
  AND U5924 ( .A(b[6]), .B(a[108]), .Z(n2518) );
  XOR U5925 ( .A(n2523), .B(n2340), .Z(n2342) );
  XOR U5926 ( .A(n2524), .B(n2525), .Z(n2340) );
  AND U5927 ( .A(n2526), .B(n2527), .Z(n2524) );
  AND U5928 ( .A(b[5]), .B(a[109]), .Z(n2523) );
  XOR U5929 ( .A(n2528), .B(n2345), .Z(n2347) );
  XOR U5930 ( .A(n2529), .B(n2530), .Z(n2345) );
  AND U5931 ( .A(n2531), .B(n2532), .Z(n2529) );
  AND U5932 ( .A(b[4]), .B(a[110]), .Z(n2528) );
  XNOR U5933 ( .A(n2533), .B(n2534), .Z(n2359) );
  NANDN U5934 ( .A(n2535), .B(n2536), .Z(n2534) );
  XOR U5935 ( .A(n2537), .B(n2350), .Z(n2352) );
  XNOR U5936 ( .A(n2538), .B(n2539), .Z(n2350) );
  AND U5937 ( .A(n2540), .B(n2541), .Z(n2538) );
  AND U5938 ( .A(b[3]), .B(a[111]), .Z(n2537) );
  XOR U5939 ( .A(n2542), .B(n2543), .Z(swire[113]) );
  XOR U5940 ( .A(n2369), .B(n2545), .Z(n2543) );
  XOR U5941 ( .A(n2368), .B(n2544), .Z(n2545) );
  IV U5942 ( .A(n2542), .Z(n2544) );
  NAND U5943 ( .A(a[113]), .B(b[0]), .Z(n2368) );
  XNOR U5944 ( .A(n2535), .B(n2536), .Z(n2369) );
  XOR U5945 ( .A(n2533), .B(n2546), .Z(n2536) );
  NAND U5946 ( .A(b[1]), .B(a[112]), .Z(n2546) );
  XOR U5947 ( .A(n2541), .B(n2547), .Z(n2535) );
  XOR U5948 ( .A(n2533), .B(n2540), .Z(n2547) );
  XNOR U5949 ( .A(n2548), .B(n2539), .Z(n2540) );
  AND U5950 ( .A(b[2]), .B(a[111]), .Z(n2548) );
  NANDN U5951 ( .A(n2549), .B(n2550), .Z(n2533) );
  XOR U5952 ( .A(n2539), .B(n2531), .Z(n2551) );
  XNOR U5953 ( .A(n2530), .B(n2526), .Z(n2552) );
  XNOR U5954 ( .A(n2525), .B(n2521), .Z(n2553) );
  XNOR U5955 ( .A(n2520), .B(n2516), .Z(n2554) );
  XNOR U5956 ( .A(n2515), .B(n2511), .Z(n2555) );
  XNOR U5957 ( .A(n2510), .B(n2506), .Z(n2556) );
  XNOR U5958 ( .A(n2505), .B(n2501), .Z(n2557) );
  XNOR U5959 ( .A(n2500), .B(n2496), .Z(n2558) );
  XNOR U5960 ( .A(n2495), .B(n2491), .Z(n2559) );
  XNOR U5961 ( .A(n2490), .B(n2486), .Z(n2560) );
  XNOR U5962 ( .A(n2485), .B(n2481), .Z(n2561) );
  XNOR U5963 ( .A(n2480), .B(n2476), .Z(n2562) );
  XNOR U5964 ( .A(n2475), .B(n2471), .Z(n2563) );
  XNOR U5965 ( .A(n2470), .B(n2466), .Z(n2564) );
  XNOR U5966 ( .A(n2465), .B(n2461), .Z(n2565) );
  XNOR U5967 ( .A(n2460), .B(n2456), .Z(n2566) );
  XNOR U5968 ( .A(n2455), .B(n2451), .Z(n2567) );
  XNOR U5969 ( .A(n2450), .B(n2446), .Z(n2568) );
  XNOR U5970 ( .A(n2445), .B(n2441), .Z(n2569) );
  XNOR U5971 ( .A(n2440), .B(n2436), .Z(n2570) );
  XNOR U5972 ( .A(n2435), .B(n2431), .Z(n2571) );
  XNOR U5973 ( .A(n2430), .B(n2426), .Z(n2572) );
  XNOR U5974 ( .A(n2425), .B(n2421), .Z(n2573) );
  XNOR U5975 ( .A(n2420), .B(n2416), .Z(n2574) );
  XNOR U5976 ( .A(n2415), .B(n2411), .Z(n2575) );
  XOR U5977 ( .A(n2410), .B(n2407), .Z(n2576) );
  XOR U5978 ( .A(n2577), .B(n2578), .Z(n2407) );
  XOR U5979 ( .A(n2405), .B(n2579), .Z(n2578) );
  XOR U5980 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U5981 ( .A(n2582), .B(n2583), .Z(n2581) );
  NAND U5982 ( .A(a[83]), .B(b[30]), .Z(n2583) );
  AND U5983 ( .A(a[82]), .B(b[31]), .Z(n2582) );
  XOR U5984 ( .A(n2584), .B(n2580), .Z(n2577) );
  XOR U5985 ( .A(n2585), .B(n2586), .Z(n2580) );
  ANDN U5986 ( .B(n2587), .A(n2588), .Z(n2585) );
  AND U5987 ( .A(a[84]), .B(b[29]), .Z(n2584) );
  XOR U5988 ( .A(n2589), .B(n2405), .Z(n2406) );
  XOR U5989 ( .A(n2590), .B(n2591), .Z(n2405) );
  AND U5990 ( .A(n2592), .B(n2593), .Z(n2590) );
  AND U5991 ( .A(a[85]), .B(b[28]), .Z(n2589) );
  XOR U5992 ( .A(n2594), .B(n2410), .Z(n2412) );
  XOR U5993 ( .A(n2595), .B(n2596), .Z(n2410) );
  AND U5994 ( .A(n2597), .B(n2598), .Z(n2595) );
  AND U5995 ( .A(a[86]), .B(b[27]), .Z(n2594) );
  XOR U5996 ( .A(n2599), .B(n2415), .Z(n2417) );
  XOR U5997 ( .A(n2600), .B(n2601), .Z(n2415) );
  AND U5998 ( .A(n2602), .B(n2603), .Z(n2600) );
  AND U5999 ( .A(a[87]), .B(b[26]), .Z(n2599) );
  XOR U6000 ( .A(n2604), .B(n2420), .Z(n2422) );
  XOR U6001 ( .A(n2605), .B(n2606), .Z(n2420) );
  AND U6002 ( .A(n2607), .B(n2608), .Z(n2605) );
  AND U6003 ( .A(a[88]), .B(b[25]), .Z(n2604) );
  XOR U6004 ( .A(n2609), .B(n2425), .Z(n2427) );
  XOR U6005 ( .A(n2610), .B(n2611), .Z(n2425) );
  AND U6006 ( .A(n2612), .B(n2613), .Z(n2610) );
  AND U6007 ( .A(a[89]), .B(b[24]), .Z(n2609) );
  XOR U6008 ( .A(n2614), .B(n2430), .Z(n2432) );
  XOR U6009 ( .A(n2615), .B(n2616), .Z(n2430) );
  AND U6010 ( .A(n2617), .B(n2618), .Z(n2615) );
  AND U6011 ( .A(a[90]), .B(b[23]), .Z(n2614) );
  XOR U6012 ( .A(n2619), .B(n2435), .Z(n2437) );
  XOR U6013 ( .A(n2620), .B(n2621), .Z(n2435) );
  AND U6014 ( .A(n2622), .B(n2623), .Z(n2620) );
  AND U6015 ( .A(a[91]), .B(b[22]), .Z(n2619) );
  XOR U6016 ( .A(n2624), .B(n2440), .Z(n2442) );
  XOR U6017 ( .A(n2625), .B(n2626), .Z(n2440) );
  AND U6018 ( .A(n2627), .B(n2628), .Z(n2625) );
  AND U6019 ( .A(a[92]), .B(b[21]), .Z(n2624) );
  XOR U6020 ( .A(n2629), .B(n2445), .Z(n2447) );
  XOR U6021 ( .A(n2630), .B(n2631), .Z(n2445) );
  AND U6022 ( .A(n2632), .B(n2633), .Z(n2630) );
  AND U6023 ( .A(a[93]), .B(b[20]), .Z(n2629) );
  XOR U6024 ( .A(n2634), .B(n2450), .Z(n2452) );
  XOR U6025 ( .A(n2635), .B(n2636), .Z(n2450) );
  AND U6026 ( .A(n2637), .B(n2638), .Z(n2635) );
  AND U6027 ( .A(a[94]), .B(b[19]), .Z(n2634) );
  XOR U6028 ( .A(n2639), .B(n2455), .Z(n2457) );
  XOR U6029 ( .A(n2640), .B(n2641), .Z(n2455) );
  AND U6030 ( .A(n2642), .B(n2643), .Z(n2640) );
  AND U6031 ( .A(b[18]), .B(a[95]), .Z(n2639) );
  XOR U6032 ( .A(n2644), .B(n2460), .Z(n2462) );
  XOR U6033 ( .A(n2645), .B(n2646), .Z(n2460) );
  AND U6034 ( .A(n2647), .B(n2648), .Z(n2645) );
  AND U6035 ( .A(b[17]), .B(a[96]), .Z(n2644) );
  XOR U6036 ( .A(n2649), .B(n2465), .Z(n2467) );
  XOR U6037 ( .A(n2650), .B(n2651), .Z(n2465) );
  AND U6038 ( .A(n2652), .B(n2653), .Z(n2650) );
  AND U6039 ( .A(b[16]), .B(a[97]), .Z(n2649) );
  XOR U6040 ( .A(n2654), .B(n2470), .Z(n2472) );
  XOR U6041 ( .A(n2655), .B(n2656), .Z(n2470) );
  AND U6042 ( .A(n2657), .B(n2658), .Z(n2655) );
  AND U6043 ( .A(b[15]), .B(a[98]), .Z(n2654) );
  XOR U6044 ( .A(n2659), .B(n2475), .Z(n2477) );
  XOR U6045 ( .A(n2660), .B(n2661), .Z(n2475) );
  AND U6046 ( .A(n2662), .B(n2663), .Z(n2660) );
  AND U6047 ( .A(b[14]), .B(a[99]), .Z(n2659) );
  XOR U6048 ( .A(n2664), .B(n2480), .Z(n2482) );
  XOR U6049 ( .A(n2665), .B(n2666), .Z(n2480) );
  AND U6050 ( .A(n2667), .B(n2668), .Z(n2665) );
  AND U6051 ( .A(b[13]), .B(a[100]), .Z(n2664) );
  XOR U6052 ( .A(n2669), .B(n2485), .Z(n2487) );
  XOR U6053 ( .A(n2670), .B(n2671), .Z(n2485) );
  AND U6054 ( .A(n2672), .B(n2673), .Z(n2670) );
  AND U6055 ( .A(b[12]), .B(a[101]), .Z(n2669) );
  XOR U6056 ( .A(n2674), .B(n2490), .Z(n2492) );
  XOR U6057 ( .A(n2675), .B(n2676), .Z(n2490) );
  AND U6058 ( .A(n2677), .B(n2678), .Z(n2675) );
  AND U6059 ( .A(b[11]), .B(a[102]), .Z(n2674) );
  XOR U6060 ( .A(n2679), .B(n2495), .Z(n2497) );
  XOR U6061 ( .A(n2680), .B(n2681), .Z(n2495) );
  AND U6062 ( .A(n2682), .B(n2683), .Z(n2680) );
  AND U6063 ( .A(b[10]), .B(a[103]), .Z(n2679) );
  XOR U6064 ( .A(n2684), .B(n2500), .Z(n2502) );
  XOR U6065 ( .A(n2685), .B(n2686), .Z(n2500) );
  AND U6066 ( .A(n2687), .B(n2688), .Z(n2685) );
  AND U6067 ( .A(b[9]), .B(a[104]), .Z(n2684) );
  XOR U6068 ( .A(n2689), .B(n2505), .Z(n2507) );
  XOR U6069 ( .A(n2690), .B(n2691), .Z(n2505) );
  AND U6070 ( .A(n2692), .B(n2693), .Z(n2690) );
  AND U6071 ( .A(b[8]), .B(a[105]), .Z(n2689) );
  XOR U6072 ( .A(n2694), .B(n2510), .Z(n2512) );
  XOR U6073 ( .A(n2695), .B(n2696), .Z(n2510) );
  AND U6074 ( .A(n2697), .B(n2698), .Z(n2695) );
  AND U6075 ( .A(b[7]), .B(a[106]), .Z(n2694) );
  XOR U6076 ( .A(n2699), .B(n2515), .Z(n2517) );
  XOR U6077 ( .A(n2700), .B(n2701), .Z(n2515) );
  AND U6078 ( .A(n2702), .B(n2703), .Z(n2700) );
  AND U6079 ( .A(b[6]), .B(a[107]), .Z(n2699) );
  XOR U6080 ( .A(n2704), .B(n2520), .Z(n2522) );
  XOR U6081 ( .A(n2705), .B(n2706), .Z(n2520) );
  AND U6082 ( .A(n2707), .B(n2708), .Z(n2705) );
  AND U6083 ( .A(b[5]), .B(a[108]), .Z(n2704) );
  XOR U6084 ( .A(n2709), .B(n2525), .Z(n2527) );
  XOR U6085 ( .A(n2710), .B(n2711), .Z(n2525) );
  AND U6086 ( .A(n2712), .B(n2713), .Z(n2710) );
  AND U6087 ( .A(b[4]), .B(a[109]), .Z(n2709) );
  XNOR U6088 ( .A(n2714), .B(n2715), .Z(n2539) );
  NANDN U6089 ( .A(n2716), .B(n2717), .Z(n2715) );
  XOR U6090 ( .A(n2718), .B(n2530), .Z(n2532) );
  XNOR U6091 ( .A(n2719), .B(n2720), .Z(n2530) );
  AND U6092 ( .A(n2721), .B(n2722), .Z(n2719) );
  AND U6093 ( .A(b[3]), .B(a[110]), .Z(n2718) );
  XNOR U6094 ( .A(n2723), .B(n2724), .Z(swire[112]) );
  XOR U6095 ( .A(n2550), .B(n2725), .Z(n2724) );
  XOR U6096 ( .A(n2549), .B(n2723), .Z(n2725) );
  NAND U6097 ( .A(a[112]), .B(b[0]), .Z(n2549) );
  XNOR U6098 ( .A(n2716), .B(n2717), .Z(n2550) );
  XOR U6099 ( .A(n2714), .B(n2726), .Z(n2717) );
  NAND U6100 ( .A(b[1]), .B(a[111]), .Z(n2726) );
  XOR U6101 ( .A(n2722), .B(n2727), .Z(n2716) );
  XOR U6102 ( .A(n2714), .B(n2721), .Z(n2727) );
  XNOR U6103 ( .A(n2728), .B(n2720), .Z(n2721) );
  AND U6104 ( .A(b[2]), .B(a[110]), .Z(n2728) );
  NANDN U6105 ( .A(n2729), .B(n2730), .Z(n2714) );
  XOR U6106 ( .A(n2720), .B(n2712), .Z(n2731) );
  XNOR U6107 ( .A(n2711), .B(n2707), .Z(n2732) );
  XNOR U6108 ( .A(n2706), .B(n2702), .Z(n2733) );
  XNOR U6109 ( .A(n2701), .B(n2697), .Z(n2734) );
  XNOR U6110 ( .A(n2696), .B(n2692), .Z(n2735) );
  XNOR U6111 ( .A(n2691), .B(n2687), .Z(n2736) );
  XNOR U6112 ( .A(n2686), .B(n2682), .Z(n2737) );
  XNOR U6113 ( .A(n2681), .B(n2677), .Z(n2738) );
  XNOR U6114 ( .A(n2676), .B(n2672), .Z(n2739) );
  XNOR U6115 ( .A(n2671), .B(n2667), .Z(n2740) );
  XNOR U6116 ( .A(n2666), .B(n2662), .Z(n2741) );
  XNOR U6117 ( .A(n2661), .B(n2657), .Z(n2742) );
  XNOR U6118 ( .A(n2656), .B(n2652), .Z(n2743) );
  XNOR U6119 ( .A(n2651), .B(n2647), .Z(n2744) );
  XNOR U6120 ( .A(n2646), .B(n2642), .Z(n2745) );
  XNOR U6121 ( .A(n2641), .B(n2637), .Z(n2746) );
  XNOR U6122 ( .A(n2636), .B(n2632), .Z(n2747) );
  XNOR U6123 ( .A(n2631), .B(n2627), .Z(n2748) );
  XNOR U6124 ( .A(n2626), .B(n2622), .Z(n2749) );
  XNOR U6125 ( .A(n2621), .B(n2617), .Z(n2750) );
  XNOR U6126 ( .A(n2616), .B(n2612), .Z(n2751) );
  XNOR U6127 ( .A(n2611), .B(n2607), .Z(n2752) );
  XNOR U6128 ( .A(n2606), .B(n2602), .Z(n2753) );
  XNOR U6129 ( .A(n2601), .B(n2597), .Z(n2754) );
  XNOR U6130 ( .A(n2596), .B(n2592), .Z(n2755) );
  XOR U6131 ( .A(n2591), .B(n2588), .Z(n2756) );
  XOR U6132 ( .A(n2757), .B(n2758), .Z(n2588) );
  XOR U6133 ( .A(n2586), .B(n2759), .Z(n2758) );
  XOR U6134 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U6135 ( .A(n2762), .B(n2763), .Z(n2761) );
  NAND U6136 ( .A(a[82]), .B(b[30]), .Z(n2763) );
  AND U6137 ( .A(a[81]), .B(b[31]), .Z(n2762) );
  XOR U6138 ( .A(n2764), .B(n2760), .Z(n2757) );
  XOR U6139 ( .A(n2765), .B(n2766), .Z(n2760) );
  ANDN U6140 ( .B(n2767), .A(n2768), .Z(n2765) );
  AND U6141 ( .A(a[83]), .B(b[29]), .Z(n2764) );
  XOR U6142 ( .A(n2769), .B(n2586), .Z(n2587) );
  XOR U6143 ( .A(n2770), .B(n2771), .Z(n2586) );
  AND U6144 ( .A(n2772), .B(n2773), .Z(n2770) );
  AND U6145 ( .A(a[84]), .B(b[28]), .Z(n2769) );
  XOR U6146 ( .A(n2774), .B(n2591), .Z(n2593) );
  XOR U6147 ( .A(n2775), .B(n2776), .Z(n2591) );
  AND U6148 ( .A(n2777), .B(n2778), .Z(n2775) );
  AND U6149 ( .A(a[85]), .B(b[27]), .Z(n2774) );
  XOR U6150 ( .A(n2779), .B(n2596), .Z(n2598) );
  XOR U6151 ( .A(n2780), .B(n2781), .Z(n2596) );
  AND U6152 ( .A(n2782), .B(n2783), .Z(n2780) );
  AND U6153 ( .A(a[86]), .B(b[26]), .Z(n2779) );
  XOR U6154 ( .A(n2784), .B(n2601), .Z(n2603) );
  XOR U6155 ( .A(n2785), .B(n2786), .Z(n2601) );
  AND U6156 ( .A(n2787), .B(n2788), .Z(n2785) );
  AND U6157 ( .A(a[87]), .B(b[25]), .Z(n2784) );
  XOR U6158 ( .A(n2789), .B(n2606), .Z(n2608) );
  XOR U6159 ( .A(n2790), .B(n2791), .Z(n2606) );
  AND U6160 ( .A(n2792), .B(n2793), .Z(n2790) );
  AND U6161 ( .A(a[88]), .B(b[24]), .Z(n2789) );
  XOR U6162 ( .A(n2794), .B(n2611), .Z(n2613) );
  XOR U6163 ( .A(n2795), .B(n2796), .Z(n2611) );
  AND U6164 ( .A(n2797), .B(n2798), .Z(n2795) );
  AND U6165 ( .A(a[89]), .B(b[23]), .Z(n2794) );
  XOR U6166 ( .A(n2799), .B(n2616), .Z(n2618) );
  XOR U6167 ( .A(n2800), .B(n2801), .Z(n2616) );
  AND U6168 ( .A(n2802), .B(n2803), .Z(n2800) );
  AND U6169 ( .A(a[90]), .B(b[22]), .Z(n2799) );
  XOR U6170 ( .A(n2804), .B(n2621), .Z(n2623) );
  XOR U6171 ( .A(n2805), .B(n2806), .Z(n2621) );
  AND U6172 ( .A(n2807), .B(n2808), .Z(n2805) );
  AND U6173 ( .A(a[91]), .B(b[21]), .Z(n2804) );
  XOR U6174 ( .A(n2809), .B(n2626), .Z(n2628) );
  XOR U6175 ( .A(n2810), .B(n2811), .Z(n2626) );
  AND U6176 ( .A(n2812), .B(n2813), .Z(n2810) );
  AND U6177 ( .A(a[92]), .B(b[20]), .Z(n2809) );
  XOR U6178 ( .A(n2814), .B(n2631), .Z(n2633) );
  XOR U6179 ( .A(n2815), .B(n2816), .Z(n2631) );
  AND U6180 ( .A(n2817), .B(n2818), .Z(n2815) );
  AND U6181 ( .A(a[93]), .B(b[19]), .Z(n2814) );
  XOR U6182 ( .A(n2819), .B(n2636), .Z(n2638) );
  XOR U6183 ( .A(n2820), .B(n2821), .Z(n2636) );
  AND U6184 ( .A(n2822), .B(n2823), .Z(n2820) );
  AND U6185 ( .A(a[94]), .B(b[18]), .Z(n2819) );
  XOR U6186 ( .A(n2824), .B(n2641), .Z(n2643) );
  XOR U6187 ( .A(n2825), .B(n2826), .Z(n2641) );
  AND U6188 ( .A(n2827), .B(n2828), .Z(n2825) );
  AND U6189 ( .A(b[17]), .B(a[95]), .Z(n2824) );
  XOR U6190 ( .A(n2829), .B(n2646), .Z(n2648) );
  XOR U6191 ( .A(n2830), .B(n2831), .Z(n2646) );
  AND U6192 ( .A(n2832), .B(n2833), .Z(n2830) );
  AND U6193 ( .A(b[16]), .B(a[96]), .Z(n2829) );
  XOR U6194 ( .A(n2834), .B(n2651), .Z(n2653) );
  XOR U6195 ( .A(n2835), .B(n2836), .Z(n2651) );
  AND U6196 ( .A(n2837), .B(n2838), .Z(n2835) );
  AND U6197 ( .A(b[15]), .B(a[97]), .Z(n2834) );
  XOR U6198 ( .A(n2839), .B(n2656), .Z(n2658) );
  XOR U6199 ( .A(n2840), .B(n2841), .Z(n2656) );
  AND U6200 ( .A(n2842), .B(n2843), .Z(n2840) );
  AND U6201 ( .A(b[14]), .B(a[98]), .Z(n2839) );
  XOR U6202 ( .A(n2844), .B(n2661), .Z(n2663) );
  XOR U6203 ( .A(n2845), .B(n2846), .Z(n2661) );
  AND U6204 ( .A(n2847), .B(n2848), .Z(n2845) );
  AND U6205 ( .A(b[13]), .B(a[99]), .Z(n2844) );
  XOR U6206 ( .A(n2849), .B(n2666), .Z(n2668) );
  XOR U6207 ( .A(n2850), .B(n2851), .Z(n2666) );
  AND U6208 ( .A(n2852), .B(n2853), .Z(n2850) );
  AND U6209 ( .A(b[12]), .B(a[100]), .Z(n2849) );
  XOR U6210 ( .A(n2854), .B(n2671), .Z(n2673) );
  XOR U6211 ( .A(n2855), .B(n2856), .Z(n2671) );
  AND U6212 ( .A(n2857), .B(n2858), .Z(n2855) );
  AND U6213 ( .A(b[11]), .B(a[101]), .Z(n2854) );
  XOR U6214 ( .A(n2859), .B(n2676), .Z(n2678) );
  XOR U6215 ( .A(n2860), .B(n2861), .Z(n2676) );
  AND U6216 ( .A(n2862), .B(n2863), .Z(n2860) );
  AND U6217 ( .A(b[10]), .B(a[102]), .Z(n2859) );
  XOR U6218 ( .A(n2864), .B(n2681), .Z(n2683) );
  XOR U6219 ( .A(n2865), .B(n2866), .Z(n2681) );
  AND U6220 ( .A(n2867), .B(n2868), .Z(n2865) );
  AND U6221 ( .A(b[9]), .B(a[103]), .Z(n2864) );
  XOR U6222 ( .A(n2869), .B(n2686), .Z(n2688) );
  XOR U6223 ( .A(n2870), .B(n2871), .Z(n2686) );
  AND U6224 ( .A(n2872), .B(n2873), .Z(n2870) );
  AND U6225 ( .A(b[8]), .B(a[104]), .Z(n2869) );
  XOR U6226 ( .A(n2874), .B(n2691), .Z(n2693) );
  XOR U6227 ( .A(n2875), .B(n2876), .Z(n2691) );
  AND U6228 ( .A(n2877), .B(n2878), .Z(n2875) );
  AND U6229 ( .A(b[7]), .B(a[105]), .Z(n2874) );
  XOR U6230 ( .A(n2879), .B(n2696), .Z(n2698) );
  XOR U6231 ( .A(n2880), .B(n2881), .Z(n2696) );
  AND U6232 ( .A(n2882), .B(n2883), .Z(n2880) );
  AND U6233 ( .A(b[6]), .B(a[106]), .Z(n2879) );
  XOR U6234 ( .A(n2884), .B(n2701), .Z(n2703) );
  XOR U6235 ( .A(n2885), .B(n2886), .Z(n2701) );
  AND U6236 ( .A(n2887), .B(n2888), .Z(n2885) );
  AND U6237 ( .A(b[5]), .B(a[107]), .Z(n2884) );
  XOR U6238 ( .A(n2889), .B(n2706), .Z(n2708) );
  XOR U6239 ( .A(n2890), .B(n2891), .Z(n2706) );
  AND U6240 ( .A(n2892), .B(n2893), .Z(n2890) );
  AND U6241 ( .A(b[4]), .B(a[108]), .Z(n2889) );
  XNOR U6242 ( .A(n2894), .B(n2895), .Z(n2720) );
  NANDN U6243 ( .A(n2896), .B(n2897), .Z(n2895) );
  XOR U6244 ( .A(n2898), .B(n2711), .Z(n2713) );
  XNOR U6245 ( .A(n2899), .B(n2900), .Z(n2711) );
  AND U6246 ( .A(n2901), .B(n2902), .Z(n2899) );
  AND U6247 ( .A(b[3]), .B(a[109]), .Z(n2898) );
  XNOR U6248 ( .A(n2903), .B(n2905), .Z(swire[111]) );
  XOR U6249 ( .A(n2903), .B(n2906), .Z(n2905) );
  XOR U6250 ( .A(n2729), .B(n2730), .Z(n2906) );
  XNOR U6251 ( .A(n2896), .B(n2897), .Z(n2730) );
  XOR U6252 ( .A(n2894), .B(n2907), .Z(n2897) );
  NAND U6253 ( .A(b[1]), .B(a[110]), .Z(n2907) );
  XOR U6254 ( .A(n2902), .B(n2908), .Z(n2896) );
  XOR U6255 ( .A(n2894), .B(n2901), .Z(n2908) );
  XNOR U6256 ( .A(n2909), .B(n2900), .Z(n2901) );
  AND U6257 ( .A(b[2]), .B(a[109]), .Z(n2909) );
  NANDN U6258 ( .A(n2910), .B(n2911), .Z(n2894) );
  XOR U6259 ( .A(n2900), .B(n2892), .Z(n2912) );
  XNOR U6260 ( .A(n2891), .B(n2887), .Z(n2913) );
  XNOR U6261 ( .A(n2886), .B(n2882), .Z(n2914) );
  XNOR U6262 ( .A(n2881), .B(n2877), .Z(n2915) );
  XNOR U6263 ( .A(n2876), .B(n2872), .Z(n2916) );
  XNOR U6264 ( .A(n2871), .B(n2867), .Z(n2917) );
  XNOR U6265 ( .A(n2866), .B(n2862), .Z(n2918) );
  XNOR U6266 ( .A(n2861), .B(n2857), .Z(n2919) );
  XNOR U6267 ( .A(n2856), .B(n2852), .Z(n2920) );
  XNOR U6268 ( .A(n2851), .B(n2847), .Z(n2921) );
  XNOR U6269 ( .A(n2846), .B(n2842), .Z(n2922) );
  XNOR U6270 ( .A(n2841), .B(n2837), .Z(n2923) );
  XNOR U6271 ( .A(n2836), .B(n2832), .Z(n2924) );
  XNOR U6272 ( .A(n2831), .B(n2827), .Z(n2925) );
  XNOR U6273 ( .A(n2826), .B(n2822), .Z(n2926) );
  XNOR U6274 ( .A(n2821), .B(n2817), .Z(n2927) );
  XNOR U6275 ( .A(n2816), .B(n2812), .Z(n2928) );
  XNOR U6276 ( .A(n2811), .B(n2807), .Z(n2929) );
  XNOR U6277 ( .A(n2806), .B(n2802), .Z(n2930) );
  XNOR U6278 ( .A(n2801), .B(n2797), .Z(n2931) );
  XNOR U6279 ( .A(n2796), .B(n2792), .Z(n2932) );
  XNOR U6280 ( .A(n2791), .B(n2787), .Z(n2933) );
  XNOR U6281 ( .A(n2786), .B(n2782), .Z(n2934) );
  XNOR U6282 ( .A(n2781), .B(n2777), .Z(n2935) );
  XNOR U6283 ( .A(n2776), .B(n2772), .Z(n2936) );
  XOR U6284 ( .A(n2771), .B(n2768), .Z(n2937) );
  XOR U6285 ( .A(n2938), .B(n2939), .Z(n2768) );
  XOR U6286 ( .A(n2766), .B(n2940), .Z(n2939) );
  XOR U6287 ( .A(n2941), .B(n2942), .Z(n2940) );
  XOR U6288 ( .A(n2943), .B(n2944), .Z(n2942) );
  NAND U6289 ( .A(a[81]), .B(b[30]), .Z(n2944) );
  AND U6290 ( .A(a[80]), .B(b[31]), .Z(n2943) );
  XOR U6291 ( .A(n2945), .B(n2941), .Z(n2938) );
  XOR U6292 ( .A(n2946), .B(n2947), .Z(n2941) );
  ANDN U6293 ( .B(n2948), .A(n2949), .Z(n2946) );
  AND U6294 ( .A(a[82]), .B(b[29]), .Z(n2945) );
  XOR U6295 ( .A(n2950), .B(n2766), .Z(n2767) );
  XOR U6296 ( .A(n2951), .B(n2952), .Z(n2766) );
  AND U6297 ( .A(n2953), .B(n2954), .Z(n2951) );
  AND U6298 ( .A(a[83]), .B(b[28]), .Z(n2950) );
  XOR U6299 ( .A(n2955), .B(n2771), .Z(n2773) );
  XOR U6300 ( .A(n2956), .B(n2957), .Z(n2771) );
  AND U6301 ( .A(n2958), .B(n2959), .Z(n2956) );
  AND U6302 ( .A(a[84]), .B(b[27]), .Z(n2955) );
  XOR U6303 ( .A(n2960), .B(n2776), .Z(n2778) );
  XOR U6304 ( .A(n2961), .B(n2962), .Z(n2776) );
  AND U6305 ( .A(n2963), .B(n2964), .Z(n2961) );
  AND U6306 ( .A(a[85]), .B(b[26]), .Z(n2960) );
  XOR U6307 ( .A(n2965), .B(n2781), .Z(n2783) );
  XOR U6308 ( .A(n2966), .B(n2967), .Z(n2781) );
  AND U6309 ( .A(n2968), .B(n2969), .Z(n2966) );
  AND U6310 ( .A(a[86]), .B(b[25]), .Z(n2965) );
  XOR U6311 ( .A(n2970), .B(n2786), .Z(n2788) );
  XOR U6312 ( .A(n2971), .B(n2972), .Z(n2786) );
  AND U6313 ( .A(n2973), .B(n2974), .Z(n2971) );
  AND U6314 ( .A(a[87]), .B(b[24]), .Z(n2970) );
  XOR U6315 ( .A(n2975), .B(n2791), .Z(n2793) );
  XOR U6316 ( .A(n2976), .B(n2977), .Z(n2791) );
  AND U6317 ( .A(n2978), .B(n2979), .Z(n2976) );
  AND U6318 ( .A(a[88]), .B(b[23]), .Z(n2975) );
  XOR U6319 ( .A(n2980), .B(n2796), .Z(n2798) );
  XOR U6320 ( .A(n2981), .B(n2982), .Z(n2796) );
  AND U6321 ( .A(n2983), .B(n2984), .Z(n2981) );
  AND U6322 ( .A(a[89]), .B(b[22]), .Z(n2980) );
  XOR U6323 ( .A(n2985), .B(n2801), .Z(n2803) );
  XOR U6324 ( .A(n2986), .B(n2987), .Z(n2801) );
  AND U6325 ( .A(n2988), .B(n2989), .Z(n2986) );
  AND U6326 ( .A(a[90]), .B(b[21]), .Z(n2985) );
  XOR U6327 ( .A(n2990), .B(n2806), .Z(n2808) );
  XOR U6328 ( .A(n2991), .B(n2992), .Z(n2806) );
  AND U6329 ( .A(n2993), .B(n2994), .Z(n2991) );
  AND U6330 ( .A(a[91]), .B(b[20]), .Z(n2990) );
  XOR U6331 ( .A(n2995), .B(n2811), .Z(n2813) );
  XOR U6332 ( .A(n2996), .B(n2997), .Z(n2811) );
  AND U6333 ( .A(n2998), .B(n2999), .Z(n2996) );
  AND U6334 ( .A(a[92]), .B(b[19]), .Z(n2995) );
  XOR U6335 ( .A(n3000), .B(n2816), .Z(n2818) );
  XOR U6336 ( .A(n3001), .B(n3002), .Z(n2816) );
  AND U6337 ( .A(n3003), .B(n3004), .Z(n3001) );
  AND U6338 ( .A(a[93]), .B(b[18]), .Z(n3000) );
  XOR U6339 ( .A(n3005), .B(n2821), .Z(n2823) );
  XOR U6340 ( .A(n3006), .B(n3007), .Z(n2821) );
  AND U6341 ( .A(n3008), .B(n3009), .Z(n3006) );
  AND U6342 ( .A(a[94]), .B(b[17]), .Z(n3005) );
  XOR U6343 ( .A(n3010), .B(n2826), .Z(n2828) );
  XOR U6344 ( .A(n3011), .B(n3012), .Z(n2826) );
  AND U6345 ( .A(n3013), .B(n3014), .Z(n3011) );
  AND U6346 ( .A(b[16]), .B(a[95]), .Z(n3010) );
  XOR U6347 ( .A(n3015), .B(n2831), .Z(n2833) );
  XOR U6348 ( .A(n3016), .B(n3017), .Z(n2831) );
  AND U6349 ( .A(n3018), .B(n3019), .Z(n3016) );
  AND U6350 ( .A(b[15]), .B(a[96]), .Z(n3015) );
  XOR U6351 ( .A(n3020), .B(n2836), .Z(n2838) );
  XOR U6352 ( .A(n3021), .B(n3022), .Z(n2836) );
  AND U6353 ( .A(n3023), .B(n3024), .Z(n3021) );
  AND U6354 ( .A(b[14]), .B(a[97]), .Z(n3020) );
  XOR U6355 ( .A(n3025), .B(n2841), .Z(n2843) );
  XOR U6356 ( .A(n3026), .B(n3027), .Z(n2841) );
  AND U6357 ( .A(n3028), .B(n3029), .Z(n3026) );
  AND U6358 ( .A(b[13]), .B(a[98]), .Z(n3025) );
  XOR U6359 ( .A(n3030), .B(n2846), .Z(n2848) );
  XOR U6360 ( .A(n3031), .B(n3032), .Z(n2846) );
  AND U6361 ( .A(n3033), .B(n3034), .Z(n3031) );
  AND U6362 ( .A(b[12]), .B(a[99]), .Z(n3030) );
  XOR U6363 ( .A(n3035), .B(n2851), .Z(n2853) );
  XOR U6364 ( .A(n3036), .B(n3037), .Z(n2851) );
  AND U6365 ( .A(n3038), .B(n3039), .Z(n3036) );
  AND U6366 ( .A(b[11]), .B(a[100]), .Z(n3035) );
  XOR U6367 ( .A(n3040), .B(n2856), .Z(n2858) );
  XOR U6368 ( .A(n3041), .B(n3042), .Z(n2856) );
  AND U6369 ( .A(n3043), .B(n3044), .Z(n3041) );
  AND U6370 ( .A(b[10]), .B(a[101]), .Z(n3040) );
  XOR U6371 ( .A(n3045), .B(n2861), .Z(n2863) );
  XOR U6372 ( .A(n3046), .B(n3047), .Z(n2861) );
  AND U6373 ( .A(n3048), .B(n3049), .Z(n3046) );
  AND U6374 ( .A(b[9]), .B(a[102]), .Z(n3045) );
  XOR U6375 ( .A(n3050), .B(n2866), .Z(n2868) );
  XOR U6376 ( .A(n3051), .B(n3052), .Z(n2866) );
  AND U6377 ( .A(n3053), .B(n3054), .Z(n3051) );
  AND U6378 ( .A(b[8]), .B(a[103]), .Z(n3050) );
  XOR U6379 ( .A(n3055), .B(n2871), .Z(n2873) );
  XOR U6380 ( .A(n3056), .B(n3057), .Z(n2871) );
  AND U6381 ( .A(n3058), .B(n3059), .Z(n3056) );
  AND U6382 ( .A(b[7]), .B(a[104]), .Z(n3055) );
  XOR U6383 ( .A(n3060), .B(n2876), .Z(n2878) );
  XOR U6384 ( .A(n3061), .B(n3062), .Z(n2876) );
  AND U6385 ( .A(n3063), .B(n3064), .Z(n3061) );
  AND U6386 ( .A(b[6]), .B(a[105]), .Z(n3060) );
  XOR U6387 ( .A(n3065), .B(n2881), .Z(n2883) );
  XOR U6388 ( .A(n3066), .B(n3067), .Z(n2881) );
  AND U6389 ( .A(n3068), .B(n3069), .Z(n3066) );
  AND U6390 ( .A(b[5]), .B(a[106]), .Z(n3065) );
  XOR U6391 ( .A(n3070), .B(n2886), .Z(n2888) );
  XOR U6392 ( .A(n3071), .B(n3072), .Z(n2886) );
  AND U6393 ( .A(n3073), .B(n3074), .Z(n3071) );
  AND U6394 ( .A(b[4]), .B(a[107]), .Z(n3070) );
  XNOR U6395 ( .A(n3075), .B(n3076), .Z(n2900) );
  NANDN U6396 ( .A(n3077), .B(n3078), .Z(n3076) );
  XOR U6397 ( .A(n3079), .B(n2891), .Z(n2893) );
  XNOR U6398 ( .A(n3080), .B(n3081), .Z(n2891) );
  AND U6399 ( .A(n3082), .B(n3083), .Z(n3080) );
  AND U6400 ( .A(b[3]), .B(a[108]), .Z(n3079) );
  NAND U6401 ( .A(a[111]), .B(b[0]), .Z(n2729) );
  IV U6402 ( .A(n2904), .Z(n2903) );
  XOR U6403 ( .A(n3084), .B(n3085), .Z(swire[110]) );
  XOR U6404 ( .A(n2910), .B(n2911), .Z(n3086) );
  XNOR U6405 ( .A(n3077), .B(n3078), .Z(n2911) );
  XOR U6406 ( .A(n3075), .B(n3087), .Z(n3078) );
  NAND U6407 ( .A(b[1]), .B(a[109]), .Z(n3087) );
  XOR U6408 ( .A(n3083), .B(n3088), .Z(n3077) );
  XOR U6409 ( .A(n3075), .B(n3082), .Z(n3088) );
  XNOR U6410 ( .A(n3089), .B(n3081), .Z(n3082) );
  AND U6411 ( .A(b[2]), .B(a[108]), .Z(n3089) );
  NANDN U6412 ( .A(n3090), .B(n3091), .Z(n3075) );
  XOR U6413 ( .A(n3081), .B(n3073), .Z(n3092) );
  XNOR U6414 ( .A(n3072), .B(n3068), .Z(n3093) );
  XNOR U6415 ( .A(n3067), .B(n3063), .Z(n3094) );
  XNOR U6416 ( .A(n3062), .B(n3058), .Z(n3095) );
  XNOR U6417 ( .A(n3057), .B(n3053), .Z(n3096) );
  XNOR U6418 ( .A(n3052), .B(n3048), .Z(n3097) );
  XNOR U6419 ( .A(n3047), .B(n3043), .Z(n3098) );
  XNOR U6420 ( .A(n3042), .B(n3038), .Z(n3099) );
  XNOR U6421 ( .A(n3037), .B(n3033), .Z(n3100) );
  XNOR U6422 ( .A(n3032), .B(n3028), .Z(n3101) );
  XNOR U6423 ( .A(n3027), .B(n3023), .Z(n3102) );
  XNOR U6424 ( .A(n3022), .B(n3018), .Z(n3103) );
  XNOR U6425 ( .A(n3017), .B(n3013), .Z(n3104) );
  XNOR U6426 ( .A(n3012), .B(n3008), .Z(n3105) );
  XNOR U6427 ( .A(n3007), .B(n3003), .Z(n3106) );
  XNOR U6428 ( .A(n3002), .B(n2998), .Z(n3107) );
  XNOR U6429 ( .A(n2997), .B(n2993), .Z(n3108) );
  XNOR U6430 ( .A(n2992), .B(n2988), .Z(n3109) );
  XNOR U6431 ( .A(n2987), .B(n2983), .Z(n3110) );
  XNOR U6432 ( .A(n2982), .B(n2978), .Z(n3111) );
  XNOR U6433 ( .A(n2977), .B(n2973), .Z(n3112) );
  XNOR U6434 ( .A(n2972), .B(n2968), .Z(n3113) );
  XNOR U6435 ( .A(n2967), .B(n2963), .Z(n3114) );
  XNOR U6436 ( .A(n2962), .B(n2958), .Z(n3115) );
  XNOR U6437 ( .A(n2957), .B(n2953), .Z(n3116) );
  XOR U6438 ( .A(n2952), .B(n2949), .Z(n3117) );
  XOR U6439 ( .A(n3118), .B(n3119), .Z(n2949) );
  XOR U6440 ( .A(n2947), .B(n3120), .Z(n3119) );
  XOR U6441 ( .A(n3121), .B(n3122), .Z(n3120) );
  XOR U6442 ( .A(n3123), .B(n3124), .Z(n3122) );
  NAND U6443 ( .A(a[80]), .B(b[30]), .Z(n3124) );
  AND U6444 ( .A(a[79]), .B(b[31]), .Z(n3123) );
  XOR U6445 ( .A(n3125), .B(n3121), .Z(n3118) );
  XOR U6446 ( .A(n3126), .B(n3127), .Z(n3121) );
  ANDN U6447 ( .B(n3128), .A(n3129), .Z(n3126) );
  AND U6448 ( .A(a[81]), .B(b[29]), .Z(n3125) );
  XOR U6449 ( .A(n3130), .B(n2947), .Z(n2948) );
  XOR U6450 ( .A(n3131), .B(n3132), .Z(n2947) );
  AND U6451 ( .A(n3133), .B(n3134), .Z(n3131) );
  AND U6452 ( .A(a[82]), .B(b[28]), .Z(n3130) );
  XOR U6453 ( .A(n3135), .B(n2952), .Z(n2954) );
  XOR U6454 ( .A(n3136), .B(n3137), .Z(n2952) );
  AND U6455 ( .A(n3138), .B(n3139), .Z(n3136) );
  AND U6456 ( .A(a[83]), .B(b[27]), .Z(n3135) );
  XOR U6457 ( .A(n3140), .B(n2957), .Z(n2959) );
  XOR U6458 ( .A(n3141), .B(n3142), .Z(n2957) );
  AND U6459 ( .A(n3143), .B(n3144), .Z(n3141) );
  AND U6460 ( .A(a[84]), .B(b[26]), .Z(n3140) );
  XOR U6461 ( .A(n3145), .B(n2962), .Z(n2964) );
  XOR U6462 ( .A(n3146), .B(n3147), .Z(n2962) );
  AND U6463 ( .A(n3148), .B(n3149), .Z(n3146) );
  AND U6464 ( .A(a[85]), .B(b[25]), .Z(n3145) );
  XOR U6465 ( .A(n3150), .B(n2967), .Z(n2969) );
  XOR U6466 ( .A(n3151), .B(n3152), .Z(n2967) );
  AND U6467 ( .A(n3153), .B(n3154), .Z(n3151) );
  AND U6468 ( .A(a[86]), .B(b[24]), .Z(n3150) );
  XOR U6469 ( .A(n3155), .B(n2972), .Z(n2974) );
  XOR U6470 ( .A(n3156), .B(n3157), .Z(n2972) );
  AND U6471 ( .A(n3158), .B(n3159), .Z(n3156) );
  AND U6472 ( .A(a[87]), .B(b[23]), .Z(n3155) );
  XOR U6473 ( .A(n3160), .B(n2977), .Z(n2979) );
  XOR U6474 ( .A(n3161), .B(n3162), .Z(n2977) );
  AND U6475 ( .A(n3163), .B(n3164), .Z(n3161) );
  AND U6476 ( .A(a[88]), .B(b[22]), .Z(n3160) );
  XOR U6477 ( .A(n3165), .B(n2982), .Z(n2984) );
  XOR U6478 ( .A(n3166), .B(n3167), .Z(n2982) );
  AND U6479 ( .A(n3168), .B(n3169), .Z(n3166) );
  AND U6480 ( .A(a[89]), .B(b[21]), .Z(n3165) );
  XOR U6481 ( .A(n3170), .B(n2987), .Z(n2989) );
  XOR U6482 ( .A(n3171), .B(n3172), .Z(n2987) );
  AND U6483 ( .A(n3173), .B(n3174), .Z(n3171) );
  AND U6484 ( .A(a[90]), .B(b[20]), .Z(n3170) );
  XOR U6485 ( .A(n3175), .B(n2992), .Z(n2994) );
  XOR U6486 ( .A(n3176), .B(n3177), .Z(n2992) );
  AND U6487 ( .A(n3178), .B(n3179), .Z(n3176) );
  AND U6488 ( .A(a[91]), .B(b[19]), .Z(n3175) );
  XOR U6489 ( .A(n3180), .B(n2997), .Z(n2999) );
  XOR U6490 ( .A(n3181), .B(n3182), .Z(n2997) );
  AND U6491 ( .A(n3183), .B(n3184), .Z(n3181) );
  AND U6492 ( .A(a[92]), .B(b[18]), .Z(n3180) );
  XOR U6493 ( .A(n3185), .B(n3002), .Z(n3004) );
  XOR U6494 ( .A(n3186), .B(n3187), .Z(n3002) );
  AND U6495 ( .A(n3188), .B(n3189), .Z(n3186) );
  AND U6496 ( .A(a[93]), .B(b[17]), .Z(n3185) );
  XOR U6497 ( .A(n3190), .B(n3007), .Z(n3009) );
  XOR U6498 ( .A(n3191), .B(n3192), .Z(n3007) );
  AND U6499 ( .A(n3193), .B(n3194), .Z(n3191) );
  AND U6500 ( .A(a[94]), .B(b[16]), .Z(n3190) );
  XOR U6501 ( .A(n3195), .B(n3012), .Z(n3014) );
  XOR U6502 ( .A(n3196), .B(n3197), .Z(n3012) );
  AND U6503 ( .A(n3198), .B(n3199), .Z(n3196) );
  AND U6504 ( .A(b[15]), .B(a[95]), .Z(n3195) );
  XOR U6505 ( .A(n3200), .B(n3017), .Z(n3019) );
  XOR U6506 ( .A(n3201), .B(n3202), .Z(n3017) );
  AND U6507 ( .A(n3203), .B(n3204), .Z(n3201) );
  AND U6508 ( .A(b[14]), .B(a[96]), .Z(n3200) );
  XOR U6509 ( .A(n3205), .B(n3022), .Z(n3024) );
  XOR U6510 ( .A(n3206), .B(n3207), .Z(n3022) );
  AND U6511 ( .A(n3208), .B(n3209), .Z(n3206) );
  AND U6512 ( .A(b[13]), .B(a[97]), .Z(n3205) );
  XOR U6513 ( .A(n3210), .B(n3027), .Z(n3029) );
  XOR U6514 ( .A(n3211), .B(n3212), .Z(n3027) );
  AND U6515 ( .A(n3213), .B(n3214), .Z(n3211) );
  AND U6516 ( .A(b[12]), .B(a[98]), .Z(n3210) );
  XOR U6517 ( .A(n3215), .B(n3032), .Z(n3034) );
  XOR U6518 ( .A(n3216), .B(n3217), .Z(n3032) );
  AND U6519 ( .A(n3218), .B(n3219), .Z(n3216) );
  AND U6520 ( .A(b[11]), .B(a[99]), .Z(n3215) );
  XOR U6521 ( .A(n3220), .B(n3037), .Z(n3039) );
  XOR U6522 ( .A(n3221), .B(n3222), .Z(n3037) );
  AND U6523 ( .A(n3223), .B(n3224), .Z(n3221) );
  AND U6524 ( .A(b[10]), .B(a[100]), .Z(n3220) );
  XOR U6525 ( .A(n3225), .B(n3042), .Z(n3044) );
  XOR U6526 ( .A(n3226), .B(n3227), .Z(n3042) );
  AND U6527 ( .A(n3228), .B(n3229), .Z(n3226) );
  AND U6528 ( .A(b[9]), .B(a[101]), .Z(n3225) );
  XOR U6529 ( .A(n3230), .B(n3047), .Z(n3049) );
  XOR U6530 ( .A(n3231), .B(n3232), .Z(n3047) );
  AND U6531 ( .A(n3233), .B(n3234), .Z(n3231) );
  AND U6532 ( .A(b[8]), .B(a[102]), .Z(n3230) );
  XOR U6533 ( .A(n3235), .B(n3052), .Z(n3054) );
  XOR U6534 ( .A(n3236), .B(n3237), .Z(n3052) );
  AND U6535 ( .A(n3238), .B(n3239), .Z(n3236) );
  AND U6536 ( .A(b[7]), .B(a[103]), .Z(n3235) );
  XOR U6537 ( .A(n3240), .B(n3057), .Z(n3059) );
  XOR U6538 ( .A(n3241), .B(n3242), .Z(n3057) );
  AND U6539 ( .A(n3243), .B(n3244), .Z(n3241) );
  AND U6540 ( .A(b[6]), .B(a[104]), .Z(n3240) );
  XOR U6541 ( .A(n3245), .B(n3062), .Z(n3064) );
  XOR U6542 ( .A(n3246), .B(n3247), .Z(n3062) );
  AND U6543 ( .A(n3248), .B(n3249), .Z(n3246) );
  AND U6544 ( .A(b[5]), .B(a[105]), .Z(n3245) );
  XOR U6545 ( .A(n3250), .B(n3067), .Z(n3069) );
  XOR U6546 ( .A(n3251), .B(n3252), .Z(n3067) );
  AND U6547 ( .A(n3253), .B(n3254), .Z(n3251) );
  AND U6548 ( .A(b[4]), .B(a[106]), .Z(n3250) );
  XNOR U6549 ( .A(n3255), .B(n3256), .Z(n3081) );
  NANDN U6550 ( .A(n3257), .B(n3258), .Z(n3256) );
  XOR U6551 ( .A(n3259), .B(n3072), .Z(n3074) );
  XNOR U6552 ( .A(n3260), .B(n3261), .Z(n3072) );
  AND U6553 ( .A(n3262), .B(n3263), .Z(n3260) );
  AND U6554 ( .A(b[3]), .B(a[107]), .Z(n3259) );
  NAND U6555 ( .A(a[110]), .B(b[0]), .Z(n2910) );
  XOR U6556 ( .A(n3264), .B(n3265), .Z(swire[109]) );
  XOR U6557 ( .A(n3090), .B(n3091), .Z(n3266) );
  XNOR U6558 ( .A(n3257), .B(n3258), .Z(n3091) );
  XOR U6559 ( .A(n3255), .B(n3267), .Z(n3258) );
  NAND U6560 ( .A(b[1]), .B(a[108]), .Z(n3267) );
  XOR U6561 ( .A(n3263), .B(n3268), .Z(n3257) );
  XOR U6562 ( .A(n3255), .B(n3262), .Z(n3268) );
  XNOR U6563 ( .A(n3269), .B(n3261), .Z(n3262) );
  AND U6564 ( .A(b[2]), .B(a[107]), .Z(n3269) );
  NANDN U6565 ( .A(n3270), .B(n3271), .Z(n3255) );
  XOR U6566 ( .A(n3261), .B(n3253), .Z(n3272) );
  XNOR U6567 ( .A(n3252), .B(n3248), .Z(n3273) );
  XNOR U6568 ( .A(n3247), .B(n3243), .Z(n3274) );
  XNOR U6569 ( .A(n3242), .B(n3238), .Z(n3275) );
  XNOR U6570 ( .A(n3237), .B(n3233), .Z(n3276) );
  XNOR U6571 ( .A(n3232), .B(n3228), .Z(n3277) );
  XNOR U6572 ( .A(n3227), .B(n3223), .Z(n3278) );
  XNOR U6573 ( .A(n3222), .B(n3218), .Z(n3279) );
  XNOR U6574 ( .A(n3217), .B(n3213), .Z(n3280) );
  XNOR U6575 ( .A(n3212), .B(n3208), .Z(n3281) );
  XNOR U6576 ( .A(n3207), .B(n3203), .Z(n3282) );
  XNOR U6577 ( .A(n3202), .B(n3198), .Z(n3283) );
  XNOR U6578 ( .A(n3197), .B(n3193), .Z(n3284) );
  XNOR U6579 ( .A(n3192), .B(n3188), .Z(n3285) );
  XNOR U6580 ( .A(n3187), .B(n3183), .Z(n3286) );
  XNOR U6581 ( .A(n3182), .B(n3178), .Z(n3287) );
  XNOR U6582 ( .A(n3177), .B(n3173), .Z(n3288) );
  XNOR U6583 ( .A(n3172), .B(n3168), .Z(n3289) );
  XNOR U6584 ( .A(n3167), .B(n3163), .Z(n3290) );
  XNOR U6585 ( .A(n3162), .B(n3158), .Z(n3291) );
  XNOR U6586 ( .A(n3157), .B(n3153), .Z(n3292) );
  XNOR U6587 ( .A(n3152), .B(n3148), .Z(n3293) );
  XNOR U6588 ( .A(n3147), .B(n3143), .Z(n3294) );
  XNOR U6589 ( .A(n3142), .B(n3138), .Z(n3295) );
  XNOR U6590 ( .A(n3137), .B(n3133), .Z(n3296) );
  XOR U6591 ( .A(n3132), .B(n3129), .Z(n3297) );
  XOR U6592 ( .A(n3298), .B(n3299), .Z(n3129) );
  XOR U6593 ( .A(n3127), .B(n3300), .Z(n3299) );
  XOR U6594 ( .A(n3301), .B(n3302), .Z(n3300) );
  XOR U6595 ( .A(n3303), .B(n3304), .Z(n3302) );
  NAND U6596 ( .A(a[79]), .B(b[30]), .Z(n3304) );
  AND U6597 ( .A(a[78]), .B(b[31]), .Z(n3303) );
  XOR U6598 ( .A(n3305), .B(n3301), .Z(n3298) );
  XOR U6599 ( .A(n3306), .B(n3307), .Z(n3301) );
  ANDN U6600 ( .B(n3308), .A(n3309), .Z(n3306) );
  AND U6601 ( .A(a[80]), .B(b[29]), .Z(n3305) );
  XOR U6602 ( .A(n3310), .B(n3127), .Z(n3128) );
  XOR U6603 ( .A(n3311), .B(n3312), .Z(n3127) );
  AND U6604 ( .A(n3313), .B(n3314), .Z(n3311) );
  AND U6605 ( .A(a[81]), .B(b[28]), .Z(n3310) );
  XOR U6606 ( .A(n3315), .B(n3132), .Z(n3134) );
  XOR U6607 ( .A(n3316), .B(n3317), .Z(n3132) );
  AND U6608 ( .A(n3318), .B(n3319), .Z(n3316) );
  AND U6609 ( .A(a[82]), .B(b[27]), .Z(n3315) );
  XOR U6610 ( .A(n3320), .B(n3137), .Z(n3139) );
  XOR U6611 ( .A(n3321), .B(n3322), .Z(n3137) );
  AND U6612 ( .A(n3323), .B(n3324), .Z(n3321) );
  AND U6613 ( .A(a[83]), .B(b[26]), .Z(n3320) );
  XOR U6614 ( .A(n3325), .B(n3142), .Z(n3144) );
  XOR U6615 ( .A(n3326), .B(n3327), .Z(n3142) );
  AND U6616 ( .A(n3328), .B(n3329), .Z(n3326) );
  AND U6617 ( .A(a[84]), .B(b[25]), .Z(n3325) );
  XOR U6618 ( .A(n3330), .B(n3147), .Z(n3149) );
  XOR U6619 ( .A(n3331), .B(n3332), .Z(n3147) );
  AND U6620 ( .A(n3333), .B(n3334), .Z(n3331) );
  AND U6621 ( .A(a[85]), .B(b[24]), .Z(n3330) );
  XOR U6622 ( .A(n3335), .B(n3152), .Z(n3154) );
  XOR U6623 ( .A(n3336), .B(n3337), .Z(n3152) );
  AND U6624 ( .A(n3338), .B(n3339), .Z(n3336) );
  AND U6625 ( .A(a[86]), .B(b[23]), .Z(n3335) );
  XOR U6626 ( .A(n3340), .B(n3157), .Z(n3159) );
  XOR U6627 ( .A(n3341), .B(n3342), .Z(n3157) );
  AND U6628 ( .A(n3343), .B(n3344), .Z(n3341) );
  AND U6629 ( .A(a[87]), .B(b[22]), .Z(n3340) );
  XOR U6630 ( .A(n3345), .B(n3162), .Z(n3164) );
  XOR U6631 ( .A(n3346), .B(n3347), .Z(n3162) );
  AND U6632 ( .A(n3348), .B(n3349), .Z(n3346) );
  AND U6633 ( .A(a[88]), .B(b[21]), .Z(n3345) );
  XOR U6634 ( .A(n3350), .B(n3167), .Z(n3169) );
  XOR U6635 ( .A(n3351), .B(n3352), .Z(n3167) );
  AND U6636 ( .A(n3353), .B(n3354), .Z(n3351) );
  AND U6637 ( .A(a[89]), .B(b[20]), .Z(n3350) );
  XOR U6638 ( .A(n3355), .B(n3172), .Z(n3174) );
  XOR U6639 ( .A(n3356), .B(n3357), .Z(n3172) );
  AND U6640 ( .A(n3358), .B(n3359), .Z(n3356) );
  AND U6641 ( .A(a[90]), .B(b[19]), .Z(n3355) );
  XOR U6642 ( .A(n3360), .B(n3177), .Z(n3179) );
  XOR U6643 ( .A(n3361), .B(n3362), .Z(n3177) );
  AND U6644 ( .A(n3363), .B(n3364), .Z(n3361) );
  AND U6645 ( .A(a[91]), .B(b[18]), .Z(n3360) );
  XOR U6646 ( .A(n3365), .B(n3182), .Z(n3184) );
  XOR U6647 ( .A(n3366), .B(n3367), .Z(n3182) );
  AND U6648 ( .A(n3368), .B(n3369), .Z(n3366) );
  AND U6649 ( .A(a[92]), .B(b[17]), .Z(n3365) );
  XOR U6650 ( .A(n3370), .B(n3187), .Z(n3189) );
  XOR U6651 ( .A(n3371), .B(n3372), .Z(n3187) );
  AND U6652 ( .A(n3373), .B(n3374), .Z(n3371) );
  AND U6653 ( .A(a[93]), .B(b[16]), .Z(n3370) );
  XOR U6654 ( .A(n3375), .B(n3192), .Z(n3194) );
  XOR U6655 ( .A(n3376), .B(n3377), .Z(n3192) );
  AND U6656 ( .A(n3378), .B(n3379), .Z(n3376) );
  AND U6657 ( .A(a[94]), .B(b[15]), .Z(n3375) );
  XOR U6658 ( .A(n3380), .B(n3197), .Z(n3199) );
  XOR U6659 ( .A(n3381), .B(n3382), .Z(n3197) );
  AND U6660 ( .A(n3383), .B(n3384), .Z(n3381) );
  AND U6661 ( .A(b[14]), .B(a[95]), .Z(n3380) );
  XOR U6662 ( .A(n3385), .B(n3202), .Z(n3204) );
  XOR U6663 ( .A(n3386), .B(n3387), .Z(n3202) );
  AND U6664 ( .A(n3388), .B(n3389), .Z(n3386) );
  AND U6665 ( .A(b[13]), .B(a[96]), .Z(n3385) );
  XOR U6666 ( .A(n3390), .B(n3207), .Z(n3209) );
  XOR U6667 ( .A(n3391), .B(n3392), .Z(n3207) );
  AND U6668 ( .A(n3393), .B(n3394), .Z(n3391) );
  AND U6669 ( .A(b[12]), .B(a[97]), .Z(n3390) );
  XOR U6670 ( .A(n3395), .B(n3212), .Z(n3214) );
  XOR U6671 ( .A(n3396), .B(n3397), .Z(n3212) );
  AND U6672 ( .A(n3398), .B(n3399), .Z(n3396) );
  AND U6673 ( .A(b[11]), .B(a[98]), .Z(n3395) );
  XOR U6674 ( .A(n3400), .B(n3217), .Z(n3219) );
  XOR U6675 ( .A(n3401), .B(n3402), .Z(n3217) );
  AND U6676 ( .A(n3403), .B(n3404), .Z(n3401) );
  AND U6677 ( .A(b[10]), .B(a[99]), .Z(n3400) );
  XOR U6678 ( .A(n3405), .B(n3222), .Z(n3224) );
  XOR U6679 ( .A(n3406), .B(n3407), .Z(n3222) );
  AND U6680 ( .A(n3408), .B(n3409), .Z(n3406) );
  AND U6681 ( .A(b[9]), .B(a[100]), .Z(n3405) );
  XOR U6682 ( .A(n3410), .B(n3227), .Z(n3229) );
  XOR U6683 ( .A(n3411), .B(n3412), .Z(n3227) );
  AND U6684 ( .A(n3413), .B(n3414), .Z(n3411) );
  AND U6685 ( .A(b[8]), .B(a[101]), .Z(n3410) );
  XOR U6686 ( .A(n3415), .B(n3232), .Z(n3234) );
  XOR U6687 ( .A(n3416), .B(n3417), .Z(n3232) );
  AND U6688 ( .A(n3418), .B(n3419), .Z(n3416) );
  AND U6689 ( .A(b[7]), .B(a[102]), .Z(n3415) );
  XOR U6690 ( .A(n3420), .B(n3237), .Z(n3239) );
  XOR U6691 ( .A(n3421), .B(n3422), .Z(n3237) );
  AND U6692 ( .A(n3423), .B(n3424), .Z(n3421) );
  AND U6693 ( .A(b[6]), .B(a[103]), .Z(n3420) );
  XOR U6694 ( .A(n3425), .B(n3242), .Z(n3244) );
  XOR U6695 ( .A(n3426), .B(n3427), .Z(n3242) );
  AND U6696 ( .A(n3428), .B(n3429), .Z(n3426) );
  AND U6697 ( .A(b[5]), .B(a[104]), .Z(n3425) );
  XOR U6698 ( .A(n3430), .B(n3247), .Z(n3249) );
  XOR U6699 ( .A(n3431), .B(n3432), .Z(n3247) );
  AND U6700 ( .A(n3433), .B(n3434), .Z(n3431) );
  AND U6701 ( .A(b[4]), .B(a[105]), .Z(n3430) );
  XNOR U6702 ( .A(n3435), .B(n3436), .Z(n3261) );
  NANDN U6703 ( .A(n3437), .B(n3438), .Z(n3436) );
  XOR U6704 ( .A(n3439), .B(n3252), .Z(n3254) );
  XNOR U6705 ( .A(n3440), .B(n3441), .Z(n3252) );
  AND U6706 ( .A(n3442), .B(n3443), .Z(n3440) );
  AND U6707 ( .A(b[3]), .B(a[106]), .Z(n3439) );
  NAND U6708 ( .A(a[109]), .B(b[0]), .Z(n3090) );
  XOR U6709 ( .A(n3444), .B(n3445), .Z(swire[108]) );
  XOR U6710 ( .A(n3270), .B(n3271), .Z(n3446) );
  XNOR U6711 ( .A(n3437), .B(n3438), .Z(n3271) );
  XOR U6712 ( .A(n3435), .B(n3447), .Z(n3438) );
  NAND U6713 ( .A(b[1]), .B(a[107]), .Z(n3447) );
  XOR U6714 ( .A(n3443), .B(n3448), .Z(n3437) );
  XOR U6715 ( .A(n3435), .B(n3442), .Z(n3448) );
  XNOR U6716 ( .A(n3449), .B(n3441), .Z(n3442) );
  AND U6717 ( .A(b[2]), .B(a[106]), .Z(n3449) );
  NANDN U6718 ( .A(n3450), .B(n3451), .Z(n3435) );
  XOR U6719 ( .A(n3441), .B(n3433), .Z(n3452) );
  XNOR U6720 ( .A(n3432), .B(n3428), .Z(n3453) );
  XNOR U6721 ( .A(n3427), .B(n3423), .Z(n3454) );
  XNOR U6722 ( .A(n3422), .B(n3418), .Z(n3455) );
  XNOR U6723 ( .A(n3417), .B(n3413), .Z(n3456) );
  XNOR U6724 ( .A(n3412), .B(n3408), .Z(n3457) );
  XNOR U6725 ( .A(n3407), .B(n3403), .Z(n3458) );
  XNOR U6726 ( .A(n3402), .B(n3398), .Z(n3459) );
  XNOR U6727 ( .A(n3397), .B(n3393), .Z(n3460) );
  XNOR U6728 ( .A(n3392), .B(n3388), .Z(n3461) );
  XNOR U6729 ( .A(n3387), .B(n3383), .Z(n3462) );
  XNOR U6730 ( .A(n3382), .B(n3378), .Z(n3463) );
  XNOR U6731 ( .A(n3377), .B(n3373), .Z(n3464) );
  XNOR U6732 ( .A(n3372), .B(n3368), .Z(n3465) );
  XNOR U6733 ( .A(n3367), .B(n3363), .Z(n3466) );
  XNOR U6734 ( .A(n3362), .B(n3358), .Z(n3467) );
  XNOR U6735 ( .A(n3357), .B(n3353), .Z(n3468) );
  XNOR U6736 ( .A(n3352), .B(n3348), .Z(n3469) );
  XNOR U6737 ( .A(n3347), .B(n3343), .Z(n3470) );
  XNOR U6738 ( .A(n3342), .B(n3338), .Z(n3471) );
  XNOR U6739 ( .A(n3337), .B(n3333), .Z(n3472) );
  XNOR U6740 ( .A(n3332), .B(n3328), .Z(n3473) );
  XNOR U6741 ( .A(n3327), .B(n3323), .Z(n3474) );
  XNOR U6742 ( .A(n3322), .B(n3318), .Z(n3475) );
  XNOR U6743 ( .A(n3317), .B(n3313), .Z(n3476) );
  XOR U6744 ( .A(n3312), .B(n3309), .Z(n3477) );
  XOR U6745 ( .A(n3478), .B(n3479), .Z(n3309) );
  XOR U6746 ( .A(n3307), .B(n3480), .Z(n3479) );
  XOR U6747 ( .A(n3481), .B(n3482), .Z(n3480) );
  XOR U6748 ( .A(n3483), .B(n3484), .Z(n3482) );
  NAND U6749 ( .A(a[78]), .B(b[30]), .Z(n3484) );
  AND U6750 ( .A(a[77]), .B(b[31]), .Z(n3483) );
  XOR U6751 ( .A(n3485), .B(n3481), .Z(n3478) );
  XOR U6752 ( .A(n3486), .B(n3487), .Z(n3481) );
  ANDN U6753 ( .B(n3488), .A(n3489), .Z(n3486) );
  AND U6754 ( .A(a[79]), .B(b[29]), .Z(n3485) );
  XOR U6755 ( .A(n3490), .B(n3307), .Z(n3308) );
  XOR U6756 ( .A(n3491), .B(n3492), .Z(n3307) );
  AND U6757 ( .A(n3493), .B(n3494), .Z(n3491) );
  AND U6758 ( .A(a[80]), .B(b[28]), .Z(n3490) );
  XOR U6759 ( .A(n3495), .B(n3312), .Z(n3314) );
  XOR U6760 ( .A(n3496), .B(n3497), .Z(n3312) );
  AND U6761 ( .A(n3498), .B(n3499), .Z(n3496) );
  AND U6762 ( .A(a[81]), .B(b[27]), .Z(n3495) );
  XOR U6763 ( .A(n3500), .B(n3317), .Z(n3319) );
  XOR U6764 ( .A(n3501), .B(n3502), .Z(n3317) );
  AND U6765 ( .A(n3503), .B(n3504), .Z(n3501) );
  AND U6766 ( .A(a[82]), .B(b[26]), .Z(n3500) );
  XOR U6767 ( .A(n3505), .B(n3322), .Z(n3324) );
  XOR U6768 ( .A(n3506), .B(n3507), .Z(n3322) );
  AND U6769 ( .A(n3508), .B(n3509), .Z(n3506) );
  AND U6770 ( .A(a[83]), .B(b[25]), .Z(n3505) );
  XOR U6771 ( .A(n3510), .B(n3327), .Z(n3329) );
  XOR U6772 ( .A(n3511), .B(n3512), .Z(n3327) );
  AND U6773 ( .A(n3513), .B(n3514), .Z(n3511) );
  AND U6774 ( .A(a[84]), .B(b[24]), .Z(n3510) );
  XOR U6775 ( .A(n3515), .B(n3332), .Z(n3334) );
  XOR U6776 ( .A(n3516), .B(n3517), .Z(n3332) );
  AND U6777 ( .A(n3518), .B(n3519), .Z(n3516) );
  AND U6778 ( .A(a[85]), .B(b[23]), .Z(n3515) );
  XOR U6779 ( .A(n3520), .B(n3337), .Z(n3339) );
  XOR U6780 ( .A(n3521), .B(n3522), .Z(n3337) );
  AND U6781 ( .A(n3523), .B(n3524), .Z(n3521) );
  AND U6782 ( .A(a[86]), .B(b[22]), .Z(n3520) );
  XOR U6783 ( .A(n3525), .B(n3342), .Z(n3344) );
  XOR U6784 ( .A(n3526), .B(n3527), .Z(n3342) );
  AND U6785 ( .A(n3528), .B(n3529), .Z(n3526) );
  AND U6786 ( .A(a[87]), .B(b[21]), .Z(n3525) );
  XOR U6787 ( .A(n3530), .B(n3347), .Z(n3349) );
  XOR U6788 ( .A(n3531), .B(n3532), .Z(n3347) );
  AND U6789 ( .A(n3533), .B(n3534), .Z(n3531) );
  AND U6790 ( .A(a[88]), .B(b[20]), .Z(n3530) );
  XOR U6791 ( .A(n3535), .B(n3352), .Z(n3354) );
  XOR U6792 ( .A(n3536), .B(n3537), .Z(n3352) );
  AND U6793 ( .A(n3538), .B(n3539), .Z(n3536) );
  AND U6794 ( .A(a[89]), .B(b[19]), .Z(n3535) );
  XOR U6795 ( .A(n3540), .B(n3357), .Z(n3359) );
  XOR U6796 ( .A(n3541), .B(n3542), .Z(n3357) );
  AND U6797 ( .A(n3543), .B(n3544), .Z(n3541) );
  AND U6798 ( .A(a[90]), .B(b[18]), .Z(n3540) );
  XOR U6799 ( .A(n3545), .B(n3362), .Z(n3364) );
  XOR U6800 ( .A(n3546), .B(n3547), .Z(n3362) );
  AND U6801 ( .A(n3548), .B(n3549), .Z(n3546) );
  AND U6802 ( .A(a[91]), .B(b[17]), .Z(n3545) );
  XOR U6803 ( .A(n3550), .B(n3367), .Z(n3369) );
  XOR U6804 ( .A(n3551), .B(n3552), .Z(n3367) );
  AND U6805 ( .A(n3553), .B(n3554), .Z(n3551) );
  AND U6806 ( .A(a[92]), .B(b[16]), .Z(n3550) );
  XOR U6807 ( .A(n3555), .B(n3372), .Z(n3374) );
  XOR U6808 ( .A(n3556), .B(n3557), .Z(n3372) );
  AND U6809 ( .A(n3558), .B(n3559), .Z(n3556) );
  AND U6810 ( .A(a[93]), .B(b[15]), .Z(n3555) );
  XOR U6811 ( .A(n3560), .B(n3377), .Z(n3379) );
  XOR U6812 ( .A(n3561), .B(n3562), .Z(n3377) );
  AND U6813 ( .A(n3563), .B(n3564), .Z(n3561) );
  AND U6814 ( .A(a[94]), .B(b[14]), .Z(n3560) );
  XOR U6815 ( .A(n3565), .B(n3382), .Z(n3384) );
  XOR U6816 ( .A(n3566), .B(n3567), .Z(n3382) );
  AND U6817 ( .A(n3568), .B(n3569), .Z(n3566) );
  AND U6818 ( .A(b[13]), .B(a[95]), .Z(n3565) );
  XOR U6819 ( .A(n3570), .B(n3387), .Z(n3389) );
  XOR U6820 ( .A(n3571), .B(n3572), .Z(n3387) );
  AND U6821 ( .A(n3573), .B(n3574), .Z(n3571) );
  AND U6822 ( .A(b[12]), .B(a[96]), .Z(n3570) );
  XOR U6823 ( .A(n3575), .B(n3392), .Z(n3394) );
  XOR U6824 ( .A(n3576), .B(n3577), .Z(n3392) );
  AND U6825 ( .A(n3578), .B(n3579), .Z(n3576) );
  AND U6826 ( .A(b[11]), .B(a[97]), .Z(n3575) );
  XOR U6827 ( .A(n3580), .B(n3397), .Z(n3399) );
  XOR U6828 ( .A(n3581), .B(n3582), .Z(n3397) );
  AND U6829 ( .A(n3583), .B(n3584), .Z(n3581) );
  AND U6830 ( .A(b[10]), .B(a[98]), .Z(n3580) );
  XOR U6831 ( .A(n3585), .B(n3402), .Z(n3404) );
  XOR U6832 ( .A(n3586), .B(n3587), .Z(n3402) );
  AND U6833 ( .A(n3588), .B(n3589), .Z(n3586) );
  AND U6834 ( .A(b[9]), .B(a[99]), .Z(n3585) );
  XOR U6835 ( .A(n3590), .B(n3407), .Z(n3409) );
  XOR U6836 ( .A(n3591), .B(n3592), .Z(n3407) );
  AND U6837 ( .A(n3593), .B(n3594), .Z(n3591) );
  AND U6838 ( .A(b[8]), .B(a[100]), .Z(n3590) );
  XOR U6839 ( .A(n3595), .B(n3412), .Z(n3414) );
  XOR U6840 ( .A(n3596), .B(n3597), .Z(n3412) );
  AND U6841 ( .A(n3598), .B(n3599), .Z(n3596) );
  AND U6842 ( .A(b[7]), .B(a[101]), .Z(n3595) );
  XOR U6843 ( .A(n3600), .B(n3417), .Z(n3419) );
  XOR U6844 ( .A(n3601), .B(n3602), .Z(n3417) );
  AND U6845 ( .A(n3603), .B(n3604), .Z(n3601) );
  AND U6846 ( .A(b[6]), .B(a[102]), .Z(n3600) );
  XOR U6847 ( .A(n3605), .B(n3422), .Z(n3424) );
  XOR U6848 ( .A(n3606), .B(n3607), .Z(n3422) );
  AND U6849 ( .A(n3608), .B(n3609), .Z(n3606) );
  AND U6850 ( .A(b[5]), .B(a[103]), .Z(n3605) );
  XOR U6851 ( .A(n3610), .B(n3427), .Z(n3429) );
  XOR U6852 ( .A(n3611), .B(n3612), .Z(n3427) );
  AND U6853 ( .A(n3613), .B(n3614), .Z(n3611) );
  AND U6854 ( .A(b[4]), .B(a[104]), .Z(n3610) );
  XNOR U6855 ( .A(n3615), .B(n3616), .Z(n3441) );
  NANDN U6856 ( .A(n3617), .B(n3618), .Z(n3616) );
  XOR U6857 ( .A(n3619), .B(n3432), .Z(n3434) );
  XNOR U6858 ( .A(n3620), .B(n3621), .Z(n3432) );
  AND U6859 ( .A(n3622), .B(n3623), .Z(n3620) );
  AND U6860 ( .A(b[3]), .B(a[105]), .Z(n3619) );
  NAND U6861 ( .A(a[108]), .B(b[0]), .Z(n3270) );
  XOR U6862 ( .A(n3624), .B(n3625), .Z(swire[107]) );
  XOR U6863 ( .A(n3450), .B(n3451), .Z(n3626) );
  XNOR U6864 ( .A(n3617), .B(n3618), .Z(n3451) );
  XOR U6865 ( .A(n3615), .B(n3627), .Z(n3618) );
  NAND U6866 ( .A(b[1]), .B(a[106]), .Z(n3627) );
  XOR U6867 ( .A(n3623), .B(n3628), .Z(n3617) );
  XOR U6868 ( .A(n3615), .B(n3622), .Z(n3628) );
  XNOR U6869 ( .A(n3629), .B(n3621), .Z(n3622) );
  AND U6870 ( .A(b[2]), .B(a[105]), .Z(n3629) );
  NANDN U6871 ( .A(n3630), .B(n3631), .Z(n3615) );
  XOR U6872 ( .A(n3621), .B(n3613), .Z(n3632) );
  XNOR U6873 ( .A(n3612), .B(n3608), .Z(n3633) );
  XNOR U6874 ( .A(n3607), .B(n3603), .Z(n3634) );
  XNOR U6875 ( .A(n3602), .B(n3598), .Z(n3635) );
  XNOR U6876 ( .A(n3597), .B(n3593), .Z(n3636) );
  XNOR U6877 ( .A(n3592), .B(n3588), .Z(n3637) );
  XNOR U6878 ( .A(n3587), .B(n3583), .Z(n3638) );
  XNOR U6879 ( .A(n3582), .B(n3578), .Z(n3639) );
  XNOR U6880 ( .A(n3577), .B(n3573), .Z(n3640) );
  XNOR U6881 ( .A(n3572), .B(n3568), .Z(n3641) );
  XNOR U6882 ( .A(n3567), .B(n3563), .Z(n3642) );
  XNOR U6883 ( .A(n3562), .B(n3558), .Z(n3643) );
  XNOR U6884 ( .A(n3557), .B(n3553), .Z(n3644) );
  XNOR U6885 ( .A(n3552), .B(n3548), .Z(n3645) );
  XNOR U6886 ( .A(n3547), .B(n3543), .Z(n3646) );
  XNOR U6887 ( .A(n3542), .B(n3538), .Z(n3647) );
  XNOR U6888 ( .A(n3537), .B(n3533), .Z(n3648) );
  XNOR U6889 ( .A(n3532), .B(n3528), .Z(n3649) );
  XNOR U6890 ( .A(n3527), .B(n3523), .Z(n3650) );
  XNOR U6891 ( .A(n3522), .B(n3518), .Z(n3651) );
  XNOR U6892 ( .A(n3517), .B(n3513), .Z(n3652) );
  XNOR U6893 ( .A(n3512), .B(n3508), .Z(n3653) );
  XNOR U6894 ( .A(n3507), .B(n3503), .Z(n3654) );
  XNOR U6895 ( .A(n3502), .B(n3498), .Z(n3655) );
  XNOR U6896 ( .A(n3497), .B(n3493), .Z(n3656) );
  XOR U6897 ( .A(n3492), .B(n3489), .Z(n3657) );
  XOR U6898 ( .A(n3658), .B(n3659), .Z(n3489) );
  XOR U6899 ( .A(n3487), .B(n3660), .Z(n3659) );
  XOR U6900 ( .A(n3661), .B(n3662), .Z(n3660) );
  XOR U6901 ( .A(n3663), .B(n3664), .Z(n3662) );
  NAND U6902 ( .A(a[77]), .B(b[30]), .Z(n3664) );
  AND U6903 ( .A(a[76]), .B(b[31]), .Z(n3663) );
  XOR U6904 ( .A(n3665), .B(n3661), .Z(n3658) );
  XOR U6905 ( .A(n3666), .B(n3667), .Z(n3661) );
  ANDN U6906 ( .B(n3668), .A(n3669), .Z(n3666) );
  AND U6907 ( .A(a[78]), .B(b[29]), .Z(n3665) );
  XOR U6908 ( .A(n3670), .B(n3487), .Z(n3488) );
  XOR U6909 ( .A(n3671), .B(n3672), .Z(n3487) );
  AND U6910 ( .A(n3673), .B(n3674), .Z(n3671) );
  AND U6911 ( .A(a[79]), .B(b[28]), .Z(n3670) );
  XOR U6912 ( .A(n3675), .B(n3492), .Z(n3494) );
  XOR U6913 ( .A(n3676), .B(n3677), .Z(n3492) );
  AND U6914 ( .A(n3678), .B(n3679), .Z(n3676) );
  AND U6915 ( .A(a[80]), .B(b[27]), .Z(n3675) );
  XOR U6916 ( .A(n3680), .B(n3497), .Z(n3499) );
  XOR U6917 ( .A(n3681), .B(n3682), .Z(n3497) );
  AND U6918 ( .A(n3683), .B(n3684), .Z(n3681) );
  AND U6919 ( .A(a[81]), .B(b[26]), .Z(n3680) );
  XOR U6920 ( .A(n3685), .B(n3502), .Z(n3504) );
  XOR U6921 ( .A(n3686), .B(n3687), .Z(n3502) );
  AND U6922 ( .A(n3688), .B(n3689), .Z(n3686) );
  AND U6923 ( .A(a[82]), .B(b[25]), .Z(n3685) );
  XOR U6924 ( .A(n3690), .B(n3507), .Z(n3509) );
  XOR U6925 ( .A(n3691), .B(n3692), .Z(n3507) );
  AND U6926 ( .A(n3693), .B(n3694), .Z(n3691) );
  AND U6927 ( .A(a[83]), .B(b[24]), .Z(n3690) );
  XOR U6928 ( .A(n3695), .B(n3512), .Z(n3514) );
  XOR U6929 ( .A(n3696), .B(n3697), .Z(n3512) );
  AND U6930 ( .A(n3698), .B(n3699), .Z(n3696) );
  AND U6931 ( .A(a[84]), .B(b[23]), .Z(n3695) );
  XOR U6932 ( .A(n3700), .B(n3517), .Z(n3519) );
  XOR U6933 ( .A(n3701), .B(n3702), .Z(n3517) );
  AND U6934 ( .A(n3703), .B(n3704), .Z(n3701) );
  AND U6935 ( .A(a[85]), .B(b[22]), .Z(n3700) );
  XOR U6936 ( .A(n3705), .B(n3522), .Z(n3524) );
  XOR U6937 ( .A(n3706), .B(n3707), .Z(n3522) );
  AND U6938 ( .A(n3708), .B(n3709), .Z(n3706) );
  AND U6939 ( .A(a[86]), .B(b[21]), .Z(n3705) );
  XOR U6940 ( .A(n3710), .B(n3527), .Z(n3529) );
  XOR U6941 ( .A(n3711), .B(n3712), .Z(n3527) );
  AND U6942 ( .A(n3713), .B(n3714), .Z(n3711) );
  AND U6943 ( .A(a[87]), .B(b[20]), .Z(n3710) );
  XOR U6944 ( .A(n3715), .B(n3532), .Z(n3534) );
  XOR U6945 ( .A(n3716), .B(n3717), .Z(n3532) );
  AND U6946 ( .A(n3718), .B(n3719), .Z(n3716) );
  AND U6947 ( .A(a[88]), .B(b[19]), .Z(n3715) );
  XOR U6948 ( .A(n3720), .B(n3537), .Z(n3539) );
  XOR U6949 ( .A(n3721), .B(n3722), .Z(n3537) );
  AND U6950 ( .A(n3723), .B(n3724), .Z(n3721) );
  AND U6951 ( .A(a[89]), .B(b[18]), .Z(n3720) );
  XOR U6952 ( .A(n3725), .B(n3542), .Z(n3544) );
  XOR U6953 ( .A(n3726), .B(n3727), .Z(n3542) );
  AND U6954 ( .A(n3728), .B(n3729), .Z(n3726) );
  AND U6955 ( .A(a[90]), .B(b[17]), .Z(n3725) );
  XOR U6956 ( .A(n3730), .B(n3547), .Z(n3549) );
  XOR U6957 ( .A(n3731), .B(n3732), .Z(n3547) );
  AND U6958 ( .A(n3733), .B(n3734), .Z(n3731) );
  AND U6959 ( .A(a[91]), .B(b[16]), .Z(n3730) );
  XOR U6960 ( .A(n3735), .B(n3552), .Z(n3554) );
  XOR U6961 ( .A(n3736), .B(n3737), .Z(n3552) );
  AND U6962 ( .A(n3738), .B(n3739), .Z(n3736) );
  AND U6963 ( .A(a[92]), .B(b[15]), .Z(n3735) );
  XOR U6964 ( .A(n3740), .B(n3557), .Z(n3559) );
  XOR U6965 ( .A(n3741), .B(n3742), .Z(n3557) );
  AND U6966 ( .A(n3743), .B(n3744), .Z(n3741) );
  AND U6967 ( .A(a[93]), .B(b[14]), .Z(n3740) );
  XOR U6968 ( .A(n3745), .B(n3562), .Z(n3564) );
  XOR U6969 ( .A(n3746), .B(n3747), .Z(n3562) );
  AND U6970 ( .A(n3748), .B(n3749), .Z(n3746) );
  AND U6971 ( .A(a[94]), .B(b[13]), .Z(n3745) );
  XOR U6972 ( .A(n3750), .B(n3567), .Z(n3569) );
  XOR U6973 ( .A(n3751), .B(n3752), .Z(n3567) );
  AND U6974 ( .A(n3753), .B(n3754), .Z(n3751) );
  AND U6975 ( .A(b[12]), .B(a[95]), .Z(n3750) );
  XOR U6976 ( .A(n3755), .B(n3572), .Z(n3574) );
  XOR U6977 ( .A(n3756), .B(n3757), .Z(n3572) );
  AND U6978 ( .A(n3758), .B(n3759), .Z(n3756) );
  AND U6979 ( .A(b[11]), .B(a[96]), .Z(n3755) );
  XOR U6980 ( .A(n3760), .B(n3577), .Z(n3579) );
  XOR U6981 ( .A(n3761), .B(n3762), .Z(n3577) );
  AND U6982 ( .A(n3763), .B(n3764), .Z(n3761) );
  AND U6983 ( .A(b[10]), .B(a[97]), .Z(n3760) );
  XOR U6984 ( .A(n3765), .B(n3582), .Z(n3584) );
  XOR U6985 ( .A(n3766), .B(n3767), .Z(n3582) );
  AND U6986 ( .A(n3768), .B(n3769), .Z(n3766) );
  AND U6987 ( .A(b[9]), .B(a[98]), .Z(n3765) );
  XOR U6988 ( .A(n3770), .B(n3587), .Z(n3589) );
  XOR U6989 ( .A(n3771), .B(n3772), .Z(n3587) );
  AND U6990 ( .A(n3773), .B(n3774), .Z(n3771) );
  AND U6991 ( .A(b[8]), .B(a[99]), .Z(n3770) );
  XOR U6992 ( .A(n3775), .B(n3592), .Z(n3594) );
  XOR U6993 ( .A(n3776), .B(n3777), .Z(n3592) );
  AND U6994 ( .A(n3778), .B(n3779), .Z(n3776) );
  AND U6995 ( .A(b[7]), .B(a[100]), .Z(n3775) );
  XOR U6996 ( .A(n3780), .B(n3597), .Z(n3599) );
  XOR U6997 ( .A(n3781), .B(n3782), .Z(n3597) );
  AND U6998 ( .A(n3783), .B(n3784), .Z(n3781) );
  AND U6999 ( .A(b[6]), .B(a[101]), .Z(n3780) );
  XOR U7000 ( .A(n3785), .B(n3602), .Z(n3604) );
  XOR U7001 ( .A(n3786), .B(n3787), .Z(n3602) );
  AND U7002 ( .A(n3788), .B(n3789), .Z(n3786) );
  AND U7003 ( .A(b[5]), .B(a[102]), .Z(n3785) );
  XOR U7004 ( .A(n3790), .B(n3607), .Z(n3609) );
  XOR U7005 ( .A(n3791), .B(n3792), .Z(n3607) );
  AND U7006 ( .A(n3793), .B(n3794), .Z(n3791) );
  AND U7007 ( .A(b[4]), .B(a[103]), .Z(n3790) );
  XNOR U7008 ( .A(n3795), .B(n3796), .Z(n3621) );
  NANDN U7009 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U7010 ( .A(n3799), .B(n3612), .Z(n3614) );
  XNOR U7011 ( .A(n3800), .B(n3801), .Z(n3612) );
  AND U7012 ( .A(n3802), .B(n3803), .Z(n3800) );
  AND U7013 ( .A(b[3]), .B(a[104]), .Z(n3799) );
  NAND U7014 ( .A(a[107]), .B(b[0]), .Z(n3450) );
  XOR U7015 ( .A(n3804), .B(n3805), .Z(swire[106]) );
  XOR U7016 ( .A(n3630), .B(n3631), .Z(n3806) );
  XNOR U7017 ( .A(n3797), .B(n3798), .Z(n3631) );
  XOR U7018 ( .A(n3795), .B(n3807), .Z(n3798) );
  NAND U7019 ( .A(b[1]), .B(a[105]), .Z(n3807) );
  XOR U7020 ( .A(n3803), .B(n3808), .Z(n3797) );
  XOR U7021 ( .A(n3795), .B(n3802), .Z(n3808) );
  XNOR U7022 ( .A(n3809), .B(n3801), .Z(n3802) );
  AND U7023 ( .A(b[2]), .B(a[104]), .Z(n3809) );
  NANDN U7024 ( .A(n3810), .B(n3811), .Z(n3795) );
  XOR U7025 ( .A(n3801), .B(n3793), .Z(n3812) );
  XNOR U7026 ( .A(n3792), .B(n3788), .Z(n3813) );
  XNOR U7027 ( .A(n3787), .B(n3783), .Z(n3814) );
  XNOR U7028 ( .A(n3782), .B(n3778), .Z(n3815) );
  XNOR U7029 ( .A(n3777), .B(n3773), .Z(n3816) );
  XNOR U7030 ( .A(n3772), .B(n3768), .Z(n3817) );
  XNOR U7031 ( .A(n3767), .B(n3763), .Z(n3818) );
  XNOR U7032 ( .A(n3762), .B(n3758), .Z(n3819) );
  XNOR U7033 ( .A(n3757), .B(n3753), .Z(n3820) );
  XNOR U7034 ( .A(n3752), .B(n3748), .Z(n3821) );
  XNOR U7035 ( .A(n3747), .B(n3743), .Z(n3822) );
  XNOR U7036 ( .A(n3742), .B(n3738), .Z(n3823) );
  XNOR U7037 ( .A(n3737), .B(n3733), .Z(n3824) );
  XNOR U7038 ( .A(n3732), .B(n3728), .Z(n3825) );
  XNOR U7039 ( .A(n3727), .B(n3723), .Z(n3826) );
  XNOR U7040 ( .A(n3722), .B(n3718), .Z(n3827) );
  XNOR U7041 ( .A(n3717), .B(n3713), .Z(n3828) );
  XNOR U7042 ( .A(n3712), .B(n3708), .Z(n3829) );
  XNOR U7043 ( .A(n3707), .B(n3703), .Z(n3830) );
  XNOR U7044 ( .A(n3702), .B(n3698), .Z(n3831) );
  XNOR U7045 ( .A(n3697), .B(n3693), .Z(n3832) );
  XNOR U7046 ( .A(n3692), .B(n3688), .Z(n3833) );
  XNOR U7047 ( .A(n3687), .B(n3683), .Z(n3834) );
  XNOR U7048 ( .A(n3682), .B(n3678), .Z(n3835) );
  XNOR U7049 ( .A(n3677), .B(n3673), .Z(n3836) );
  XOR U7050 ( .A(n3672), .B(n3669), .Z(n3837) );
  XOR U7051 ( .A(n3838), .B(n3839), .Z(n3669) );
  XOR U7052 ( .A(n3667), .B(n3840), .Z(n3839) );
  XOR U7053 ( .A(n3841), .B(n3842), .Z(n3840) );
  XOR U7054 ( .A(n3843), .B(n3844), .Z(n3842) );
  NAND U7055 ( .A(a[76]), .B(b[30]), .Z(n3844) );
  AND U7056 ( .A(a[75]), .B(b[31]), .Z(n3843) );
  XOR U7057 ( .A(n3845), .B(n3841), .Z(n3838) );
  XOR U7058 ( .A(n3846), .B(n3847), .Z(n3841) );
  ANDN U7059 ( .B(n3848), .A(n3849), .Z(n3846) );
  AND U7060 ( .A(a[77]), .B(b[29]), .Z(n3845) );
  XOR U7061 ( .A(n3850), .B(n3667), .Z(n3668) );
  XOR U7062 ( .A(n3851), .B(n3852), .Z(n3667) );
  AND U7063 ( .A(n3853), .B(n3854), .Z(n3851) );
  AND U7064 ( .A(a[78]), .B(b[28]), .Z(n3850) );
  XOR U7065 ( .A(n3855), .B(n3672), .Z(n3674) );
  XOR U7066 ( .A(n3856), .B(n3857), .Z(n3672) );
  AND U7067 ( .A(n3858), .B(n3859), .Z(n3856) );
  AND U7068 ( .A(a[79]), .B(b[27]), .Z(n3855) );
  XOR U7069 ( .A(n3860), .B(n3677), .Z(n3679) );
  XOR U7070 ( .A(n3861), .B(n3862), .Z(n3677) );
  AND U7071 ( .A(n3863), .B(n3864), .Z(n3861) );
  AND U7072 ( .A(a[80]), .B(b[26]), .Z(n3860) );
  XOR U7073 ( .A(n3865), .B(n3682), .Z(n3684) );
  XOR U7074 ( .A(n3866), .B(n3867), .Z(n3682) );
  AND U7075 ( .A(n3868), .B(n3869), .Z(n3866) );
  AND U7076 ( .A(a[81]), .B(b[25]), .Z(n3865) );
  XOR U7077 ( .A(n3870), .B(n3687), .Z(n3689) );
  XOR U7078 ( .A(n3871), .B(n3872), .Z(n3687) );
  AND U7079 ( .A(n3873), .B(n3874), .Z(n3871) );
  AND U7080 ( .A(a[82]), .B(b[24]), .Z(n3870) );
  XOR U7081 ( .A(n3875), .B(n3692), .Z(n3694) );
  XOR U7082 ( .A(n3876), .B(n3877), .Z(n3692) );
  AND U7083 ( .A(n3878), .B(n3879), .Z(n3876) );
  AND U7084 ( .A(a[83]), .B(b[23]), .Z(n3875) );
  XOR U7085 ( .A(n3880), .B(n3697), .Z(n3699) );
  XOR U7086 ( .A(n3881), .B(n3882), .Z(n3697) );
  AND U7087 ( .A(n3883), .B(n3884), .Z(n3881) );
  AND U7088 ( .A(a[84]), .B(b[22]), .Z(n3880) );
  XOR U7089 ( .A(n3885), .B(n3702), .Z(n3704) );
  XOR U7090 ( .A(n3886), .B(n3887), .Z(n3702) );
  AND U7091 ( .A(n3888), .B(n3889), .Z(n3886) );
  AND U7092 ( .A(a[85]), .B(b[21]), .Z(n3885) );
  XOR U7093 ( .A(n3890), .B(n3707), .Z(n3709) );
  XOR U7094 ( .A(n3891), .B(n3892), .Z(n3707) );
  AND U7095 ( .A(n3893), .B(n3894), .Z(n3891) );
  AND U7096 ( .A(a[86]), .B(b[20]), .Z(n3890) );
  XOR U7097 ( .A(n3895), .B(n3712), .Z(n3714) );
  XOR U7098 ( .A(n3896), .B(n3897), .Z(n3712) );
  AND U7099 ( .A(n3898), .B(n3899), .Z(n3896) );
  AND U7100 ( .A(a[87]), .B(b[19]), .Z(n3895) );
  XOR U7101 ( .A(n3900), .B(n3717), .Z(n3719) );
  XOR U7102 ( .A(n3901), .B(n3902), .Z(n3717) );
  AND U7103 ( .A(n3903), .B(n3904), .Z(n3901) );
  AND U7104 ( .A(a[88]), .B(b[18]), .Z(n3900) );
  XOR U7105 ( .A(n3905), .B(n3722), .Z(n3724) );
  XOR U7106 ( .A(n3906), .B(n3907), .Z(n3722) );
  AND U7107 ( .A(n3908), .B(n3909), .Z(n3906) );
  AND U7108 ( .A(a[89]), .B(b[17]), .Z(n3905) );
  XOR U7109 ( .A(n3910), .B(n3727), .Z(n3729) );
  XOR U7110 ( .A(n3911), .B(n3912), .Z(n3727) );
  AND U7111 ( .A(n3913), .B(n3914), .Z(n3911) );
  AND U7112 ( .A(a[90]), .B(b[16]), .Z(n3910) );
  XOR U7113 ( .A(n3915), .B(n3732), .Z(n3734) );
  XOR U7114 ( .A(n3916), .B(n3917), .Z(n3732) );
  AND U7115 ( .A(n3918), .B(n3919), .Z(n3916) );
  AND U7116 ( .A(a[91]), .B(b[15]), .Z(n3915) );
  XOR U7117 ( .A(n3920), .B(n3737), .Z(n3739) );
  XOR U7118 ( .A(n3921), .B(n3922), .Z(n3737) );
  AND U7119 ( .A(n3923), .B(n3924), .Z(n3921) );
  AND U7120 ( .A(a[92]), .B(b[14]), .Z(n3920) );
  XOR U7121 ( .A(n3925), .B(n3742), .Z(n3744) );
  XOR U7122 ( .A(n3926), .B(n3927), .Z(n3742) );
  AND U7123 ( .A(n3928), .B(n3929), .Z(n3926) );
  AND U7124 ( .A(a[93]), .B(b[13]), .Z(n3925) );
  XOR U7125 ( .A(n3930), .B(n3747), .Z(n3749) );
  XOR U7126 ( .A(n3931), .B(n3932), .Z(n3747) );
  AND U7127 ( .A(n3933), .B(n3934), .Z(n3931) );
  AND U7128 ( .A(a[94]), .B(b[12]), .Z(n3930) );
  XOR U7129 ( .A(n3935), .B(n3752), .Z(n3754) );
  XOR U7130 ( .A(n3936), .B(n3937), .Z(n3752) );
  AND U7131 ( .A(n3938), .B(n3939), .Z(n3936) );
  AND U7132 ( .A(b[11]), .B(a[95]), .Z(n3935) );
  XOR U7133 ( .A(n3940), .B(n3757), .Z(n3759) );
  XOR U7134 ( .A(n3941), .B(n3942), .Z(n3757) );
  AND U7135 ( .A(n3943), .B(n3944), .Z(n3941) );
  AND U7136 ( .A(b[10]), .B(a[96]), .Z(n3940) );
  XOR U7137 ( .A(n3945), .B(n3762), .Z(n3764) );
  XOR U7138 ( .A(n3946), .B(n3947), .Z(n3762) );
  AND U7139 ( .A(n3948), .B(n3949), .Z(n3946) );
  AND U7140 ( .A(b[9]), .B(a[97]), .Z(n3945) );
  XOR U7141 ( .A(n3950), .B(n3767), .Z(n3769) );
  XOR U7142 ( .A(n3951), .B(n3952), .Z(n3767) );
  AND U7143 ( .A(n3953), .B(n3954), .Z(n3951) );
  AND U7144 ( .A(b[8]), .B(a[98]), .Z(n3950) );
  XOR U7145 ( .A(n3955), .B(n3772), .Z(n3774) );
  XOR U7146 ( .A(n3956), .B(n3957), .Z(n3772) );
  AND U7147 ( .A(n3958), .B(n3959), .Z(n3956) );
  AND U7148 ( .A(b[7]), .B(a[99]), .Z(n3955) );
  XOR U7149 ( .A(n3960), .B(n3777), .Z(n3779) );
  XOR U7150 ( .A(n3961), .B(n3962), .Z(n3777) );
  AND U7151 ( .A(n3963), .B(n3964), .Z(n3961) );
  AND U7152 ( .A(b[6]), .B(a[100]), .Z(n3960) );
  XOR U7153 ( .A(n3965), .B(n3782), .Z(n3784) );
  XOR U7154 ( .A(n3966), .B(n3967), .Z(n3782) );
  AND U7155 ( .A(n3968), .B(n3969), .Z(n3966) );
  AND U7156 ( .A(b[5]), .B(a[101]), .Z(n3965) );
  XOR U7157 ( .A(n3970), .B(n3787), .Z(n3789) );
  XOR U7158 ( .A(n3971), .B(n3972), .Z(n3787) );
  AND U7159 ( .A(n3973), .B(n3974), .Z(n3971) );
  AND U7160 ( .A(b[4]), .B(a[102]), .Z(n3970) );
  XNOR U7161 ( .A(n3975), .B(n3976), .Z(n3801) );
  NANDN U7162 ( .A(n3977), .B(n3978), .Z(n3976) );
  XOR U7163 ( .A(n3979), .B(n3792), .Z(n3794) );
  XNOR U7164 ( .A(n3980), .B(n3981), .Z(n3792) );
  AND U7165 ( .A(n3982), .B(n3983), .Z(n3980) );
  AND U7166 ( .A(b[3]), .B(a[103]), .Z(n3979) );
  NAND U7167 ( .A(a[106]), .B(b[0]), .Z(n3630) );
  XOR U7168 ( .A(n3984), .B(n3985), .Z(swire[105]) );
  XOR U7169 ( .A(n3810), .B(n3811), .Z(n3986) );
  XNOR U7170 ( .A(n3977), .B(n3978), .Z(n3811) );
  XOR U7171 ( .A(n3975), .B(n3987), .Z(n3978) );
  NAND U7172 ( .A(b[1]), .B(a[104]), .Z(n3987) );
  XOR U7173 ( .A(n3983), .B(n3988), .Z(n3977) );
  XOR U7174 ( .A(n3975), .B(n3982), .Z(n3988) );
  XNOR U7175 ( .A(n3989), .B(n3981), .Z(n3982) );
  AND U7176 ( .A(b[2]), .B(a[103]), .Z(n3989) );
  NANDN U7177 ( .A(n3990), .B(n3991), .Z(n3975) );
  XOR U7178 ( .A(n3981), .B(n3973), .Z(n3992) );
  XNOR U7179 ( .A(n3972), .B(n3968), .Z(n3993) );
  XNOR U7180 ( .A(n3967), .B(n3963), .Z(n3994) );
  XNOR U7181 ( .A(n3962), .B(n3958), .Z(n3995) );
  XNOR U7182 ( .A(n3957), .B(n3953), .Z(n3996) );
  XNOR U7183 ( .A(n3952), .B(n3948), .Z(n3997) );
  XNOR U7184 ( .A(n3947), .B(n3943), .Z(n3998) );
  XNOR U7185 ( .A(n3942), .B(n3938), .Z(n3999) );
  XNOR U7186 ( .A(n3937), .B(n3933), .Z(n4000) );
  XNOR U7187 ( .A(n3932), .B(n3928), .Z(n4001) );
  XNOR U7188 ( .A(n3927), .B(n3923), .Z(n4002) );
  XNOR U7189 ( .A(n3922), .B(n3918), .Z(n4003) );
  XNOR U7190 ( .A(n3917), .B(n3913), .Z(n4004) );
  XNOR U7191 ( .A(n3912), .B(n3908), .Z(n4005) );
  XNOR U7192 ( .A(n3907), .B(n3903), .Z(n4006) );
  XNOR U7193 ( .A(n3902), .B(n3898), .Z(n4007) );
  XNOR U7194 ( .A(n3897), .B(n3893), .Z(n4008) );
  XNOR U7195 ( .A(n3892), .B(n3888), .Z(n4009) );
  XNOR U7196 ( .A(n3887), .B(n3883), .Z(n4010) );
  XNOR U7197 ( .A(n3882), .B(n3878), .Z(n4011) );
  XNOR U7198 ( .A(n3877), .B(n3873), .Z(n4012) );
  XNOR U7199 ( .A(n3872), .B(n3868), .Z(n4013) );
  XNOR U7200 ( .A(n3867), .B(n3863), .Z(n4014) );
  XNOR U7201 ( .A(n3862), .B(n3858), .Z(n4015) );
  XNOR U7202 ( .A(n3857), .B(n3853), .Z(n4016) );
  XOR U7203 ( .A(n3852), .B(n3849), .Z(n4017) );
  XOR U7204 ( .A(n4018), .B(n4019), .Z(n3849) );
  XOR U7205 ( .A(n3847), .B(n4020), .Z(n4019) );
  XOR U7206 ( .A(n4021), .B(n4022), .Z(n4020) );
  XOR U7207 ( .A(n4023), .B(n4024), .Z(n4022) );
  NAND U7208 ( .A(a[75]), .B(b[30]), .Z(n4024) );
  AND U7209 ( .A(a[74]), .B(b[31]), .Z(n4023) );
  XOR U7210 ( .A(n4025), .B(n4021), .Z(n4018) );
  XOR U7211 ( .A(n4026), .B(n4027), .Z(n4021) );
  ANDN U7212 ( .B(n4028), .A(n4029), .Z(n4026) );
  AND U7213 ( .A(a[76]), .B(b[29]), .Z(n4025) );
  XOR U7214 ( .A(n4030), .B(n3847), .Z(n3848) );
  XOR U7215 ( .A(n4031), .B(n4032), .Z(n3847) );
  AND U7216 ( .A(n4033), .B(n4034), .Z(n4031) );
  AND U7217 ( .A(a[77]), .B(b[28]), .Z(n4030) );
  XOR U7218 ( .A(n4035), .B(n3852), .Z(n3854) );
  XOR U7219 ( .A(n4036), .B(n4037), .Z(n3852) );
  AND U7220 ( .A(n4038), .B(n4039), .Z(n4036) );
  AND U7221 ( .A(a[78]), .B(b[27]), .Z(n4035) );
  XOR U7222 ( .A(n4040), .B(n3857), .Z(n3859) );
  XOR U7223 ( .A(n4041), .B(n4042), .Z(n3857) );
  AND U7224 ( .A(n4043), .B(n4044), .Z(n4041) );
  AND U7225 ( .A(a[79]), .B(b[26]), .Z(n4040) );
  XOR U7226 ( .A(n4045), .B(n3862), .Z(n3864) );
  XOR U7227 ( .A(n4046), .B(n4047), .Z(n3862) );
  AND U7228 ( .A(n4048), .B(n4049), .Z(n4046) );
  AND U7229 ( .A(a[80]), .B(b[25]), .Z(n4045) );
  XOR U7230 ( .A(n4050), .B(n3867), .Z(n3869) );
  XOR U7231 ( .A(n4051), .B(n4052), .Z(n3867) );
  AND U7232 ( .A(n4053), .B(n4054), .Z(n4051) );
  AND U7233 ( .A(a[81]), .B(b[24]), .Z(n4050) );
  XOR U7234 ( .A(n4055), .B(n3872), .Z(n3874) );
  XOR U7235 ( .A(n4056), .B(n4057), .Z(n3872) );
  AND U7236 ( .A(n4058), .B(n4059), .Z(n4056) );
  AND U7237 ( .A(a[82]), .B(b[23]), .Z(n4055) );
  XOR U7238 ( .A(n4060), .B(n3877), .Z(n3879) );
  XOR U7239 ( .A(n4061), .B(n4062), .Z(n3877) );
  AND U7240 ( .A(n4063), .B(n4064), .Z(n4061) );
  AND U7241 ( .A(a[83]), .B(b[22]), .Z(n4060) );
  XOR U7242 ( .A(n4065), .B(n3882), .Z(n3884) );
  XOR U7243 ( .A(n4066), .B(n4067), .Z(n3882) );
  AND U7244 ( .A(n4068), .B(n4069), .Z(n4066) );
  AND U7245 ( .A(a[84]), .B(b[21]), .Z(n4065) );
  XOR U7246 ( .A(n4070), .B(n3887), .Z(n3889) );
  XOR U7247 ( .A(n4071), .B(n4072), .Z(n3887) );
  AND U7248 ( .A(n4073), .B(n4074), .Z(n4071) );
  AND U7249 ( .A(a[85]), .B(b[20]), .Z(n4070) );
  XOR U7250 ( .A(n4075), .B(n3892), .Z(n3894) );
  XOR U7251 ( .A(n4076), .B(n4077), .Z(n3892) );
  AND U7252 ( .A(n4078), .B(n4079), .Z(n4076) );
  AND U7253 ( .A(a[86]), .B(b[19]), .Z(n4075) );
  XOR U7254 ( .A(n4080), .B(n3897), .Z(n3899) );
  XOR U7255 ( .A(n4081), .B(n4082), .Z(n3897) );
  AND U7256 ( .A(n4083), .B(n4084), .Z(n4081) );
  AND U7257 ( .A(a[87]), .B(b[18]), .Z(n4080) );
  XOR U7258 ( .A(n4085), .B(n3902), .Z(n3904) );
  XOR U7259 ( .A(n4086), .B(n4087), .Z(n3902) );
  AND U7260 ( .A(n4088), .B(n4089), .Z(n4086) );
  AND U7261 ( .A(a[88]), .B(b[17]), .Z(n4085) );
  XOR U7262 ( .A(n4090), .B(n3907), .Z(n3909) );
  XOR U7263 ( .A(n4091), .B(n4092), .Z(n3907) );
  AND U7264 ( .A(n4093), .B(n4094), .Z(n4091) );
  AND U7265 ( .A(a[89]), .B(b[16]), .Z(n4090) );
  XOR U7266 ( .A(n4095), .B(n3912), .Z(n3914) );
  XOR U7267 ( .A(n4096), .B(n4097), .Z(n3912) );
  AND U7268 ( .A(n4098), .B(n4099), .Z(n4096) );
  AND U7269 ( .A(a[90]), .B(b[15]), .Z(n4095) );
  XOR U7270 ( .A(n4100), .B(n3917), .Z(n3919) );
  XOR U7271 ( .A(n4101), .B(n4102), .Z(n3917) );
  AND U7272 ( .A(n4103), .B(n4104), .Z(n4101) );
  AND U7273 ( .A(a[91]), .B(b[14]), .Z(n4100) );
  XOR U7274 ( .A(n4105), .B(n3922), .Z(n3924) );
  XOR U7275 ( .A(n4106), .B(n4107), .Z(n3922) );
  AND U7276 ( .A(n4108), .B(n4109), .Z(n4106) );
  AND U7277 ( .A(a[92]), .B(b[13]), .Z(n4105) );
  XOR U7278 ( .A(n4110), .B(n3927), .Z(n3929) );
  XOR U7279 ( .A(n4111), .B(n4112), .Z(n3927) );
  AND U7280 ( .A(n4113), .B(n4114), .Z(n4111) );
  AND U7281 ( .A(a[93]), .B(b[12]), .Z(n4110) );
  XOR U7282 ( .A(n4115), .B(n3932), .Z(n3934) );
  XOR U7283 ( .A(n4116), .B(n4117), .Z(n3932) );
  AND U7284 ( .A(n4118), .B(n4119), .Z(n4116) );
  AND U7285 ( .A(a[94]), .B(b[11]), .Z(n4115) );
  XOR U7286 ( .A(n4120), .B(n3937), .Z(n3939) );
  XOR U7287 ( .A(n4121), .B(n4122), .Z(n3937) );
  AND U7288 ( .A(n4123), .B(n4124), .Z(n4121) );
  AND U7289 ( .A(b[10]), .B(a[95]), .Z(n4120) );
  XOR U7290 ( .A(n4125), .B(n3942), .Z(n3944) );
  XOR U7291 ( .A(n4126), .B(n4127), .Z(n3942) );
  AND U7292 ( .A(n4128), .B(n4129), .Z(n4126) );
  AND U7293 ( .A(b[9]), .B(a[96]), .Z(n4125) );
  XOR U7294 ( .A(n4130), .B(n3947), .Z(n3949) );
  XOR U7295 ( .A(n4131), .B(n4132), .Z(n3947) );
  AND U7296 ( .A(n4133), .B(n4134), .Z(n4131) );
  AND U7297 ( .A(b[8]), .B(a[97]), .Z(n4130) );
  XOR U7298 ( .A(n4135), .B(n3952), .Z(n3954) );
  XOR U7299 ( .A(n4136), .B(n4137), .Z(n3952) );
  AND U7300 ( .A(n4138), .B(n4139), .Z(n4136) );
  AND U7301 ( .A(b[7]), .B(a[98]), .Z(n4135) );
  XOR U7302 ( .A(n4140), .B(n3957), .Z(n3959) );
  XOR U7303 ( .A(n4141), .B(n4142), .Z(n3957) );
  AND U7304 ( .A(n4143), .B(n4144), .Z(n4141) );
  AND U7305 ( .A(b[6]), .B(a[99]), .Z(n4140) );
  XOR U7306 ( .A(n4145), .B(n3962), .Z(n3964) );
  XOR U7307 ( .A(n4146), .B(n4147), .Z(n3962) );
  AND U7308 ( .A(n4148), .B(n4149), .Z(n4146) );
  AND U7309 ( .A(b[5]), .B(a[100]), .Z(n4145) );
  XOR U7310 ( .A(n4150), .B(n3967), .Z(n3969) );
  XOR U7311 ( .A(n4151), .B(n4152), .Z(n3967) );
  AND U7312 ( .A(n4153), .B(n4154), .Z(n4151) );
  AND U7313 ( .A(b[4]), .B(a[101]), .Z(n4150) );
  XNOR U7314 ( .A(n4155), .B(n4156), .Z(n3981) );
  NANDN U7315 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U7316 ( .A(n4159), .B(n3972), .Z(n3974) );
  XNOR U7317 ( .A(n4160), .B(n4161), .Z(n3972) );
  AND U7318 ( .A(n4162), .B(n4163), .Z(n4160) );
  AND U7319 ( .A(b[3]), .B(a[102]), .Z(n4159) );
  NAND U7320 ( .A(a[105]), .B(b[0]), .Z(n3810) );
  XOR U7321 ( .A(n4164), .B(n4165), .Z(swire[104]) );
  XOR U7322 ( .A(n3990), .B(n3991), .Z(n4166) );
  XNOR U7323 ( .A(n4157), .B(n4158), .Z(n3991) );
  XOR U7324 ( .A(n4155), .B(n4167), .Z(n4158) );
  NAND U7325 ( .A(b[1]), .B(a[103]), .Z(n4167) );
  XOR U7326 ( .A(n4163), .B(n4168), .Z(n4157) );
  XOR U7327 ( .A(n4155), .B(n4162), .Z(n4168) );
  XNOR U7328 ( .A(n4169), .B(n4161), .Z(n4162) );
  AND U7329 ( .A(b[2]), .B(a[102]), .Z(n4169) );
  NANDN U7330 ( .A(n4170), .B(n4171), .Z(n4155) );
  XOR U7331 ( .A(n4161), .B(n4153), .Z(n4172) );
  XNOR U7332 ( .A(n4152), .B(n4148), .Z(n4173) );
  XNOR U7333 ( .A(n4147), .B(n4143), .Z(n4174) );
  XNOR U7334 ( .A(n4142), .B(n4138), .Z(n4175) );
  XNOR U7335 ( .A(n4137), .B(n4133), .Z(n4176) );
  XNOR U7336 ( .A(n4132), .B(n4128), .Z(n4177) );
  XNOR U7337 ( .A(n4127), .B(n4123), .Z(n4178) );
  XNOR U7338 ( .A(n4122), .B(n4118), .Z(n4179) );
  XNOR U7339 ( .A(n4117), .B(n4113), .Z(n4180) );
  XNOR U7340 ( .A(n4112), .B(n4108), .Z(n4181) );
  XNOR U7341 ( .A(n4107), .B(n4103), .Z(n4182) );
  XNOR U7342 ( .A(n4102), .B(n4098), .Z(n4183) );
  XNOR U7343 ( .A(n4097), .B(n4093), .Z(n4184) );
  XNOR U7344 ( .A(n4092), .B(n4088), .Z(n4185) );
  XNOR U7345 ( .A(n4087), .B(n4083), .Z(n4186) );
  XNOR U7346 ( .A(n4082), .B(n4078), .Z(n4187) );
  XNOR U7347 ( .A(n4077), .B(n4073), .Z(n4188) );
  XNOR U7348 ( .A(n4072), .B(n4068), .Z(n4189) );
  XNOR U7349 ( .A(n4067), .B(n4063), .Z(n4190) );
  XNOR U7350 ( .A(n4062), .B(n4058), .Z(n4191) );
  XNOR U7351 ( .A(n4057), .B(n4053), .Z(n4192) );
  XNOR U7352 ( .A(n4052), .B(n4048), .Z(n4193) );
  XNOR U7353 ( .A(n4047), .B(n4043), .Z(n4194) );
  XNOR U7354 ( .A(n4042), .B(n4038), .Z(n4195) );
  XNOR U7355 ( .A(n4037), .B(n4033), .Z(n4196) );
  XOR U7356 ( .A(n4032), .B(n4029), .Z(n4197) );
  XOR U7357 ( .A(n4198), .B(n4199), .Z(n4029) );
  XOR U7358 ( .A(n4027), .B(n4200), .Z(n4199) );
  XOR U7359 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U7360 ( .A(n4203), .B(n4204), .Z(n4202) );
  NAND U7361 ( .A(a[74]), .B(b[30]), .Z(n4204) );
  AND U7362 ( .A(a[73]), .B(b[31]), .Z(n4203) );
  XOR U7363 ( .A(n4205), .B(n4201), .Z(n4198) );
  XOR U7364 ( .A(n4206), .B(n4207), .Z(n4201) );
  ANDN U7365 ( .B(n4208), .A(n4209), .Z(n4206) );
  AND U7366 ( .A(a[75]), .B(b[29]), .Z(n4205) );
  XOR U7367 ( .A(n4210), .B(n4027), .Z(n4028) );
  XOR U7368 ( .A(n4211), .B(n4212), .Z(n4027) );
  AND U7369 ( .A(n4213), .B(n4214), .Z(n4211) );
  AND U7370 ( .A(a[76]), .B(b[28]), .Z(n4210) );
  XOR U7371 ( .A(n4215), .B(n4032), .Z(n4034) );
  XOR U7372 ( .A(n4216), .B(n4217), .Z(n4032) );
  AND U7373 ( .A(n4218), .B(n4219), .Z(n4216) );
  AND U7374 ( .A(a[77]), .B(b[27]), .Z(n4215) );
  XOR U7375 ( .A(n4220), .B(n4037), .Z(n4039) );
  XOR U7376 ( .A(n4221), .B(n4222), .Z(n4037) );
  AND U7377 ( .A(n4223), .B(n4224), .Z(n4221) );
  AND U7378 ( .A(a[78]), .B(b[26]), .Z(n4220) );
  XOR U7379 ( .A(n4225), .B(n4042), .Z(n4044) );
  XOR U7380 ( .A(n4226), .B(n4227), .Z(n4042) );
  AND U7381 ( .A(n4228), .B(n4229), .Z(n4226) );
  AND U7382 ( .A(a[79]), .B(b[25]), .Z(n4225) );
  XOR U7383 ( .A(n4230), .B(n4047), .Z(n4049) );
  XOR U7384 ( .A(n4231), .B(n4232), .Z(n4047) );
  AND U7385 ( .A(n4233), .B(n4234), .Z(n4231) );
  AND U7386 ( .A(a[80]), .B(b[24]), .Z(n4230) );
  XOR U7387 ( .A(n4235), .B(n4052), .Z(n4054) );
  XOR U7388 ( .A(n4236), .B(n4237), .Z(n4052) );
  AND U7389 ( .A(n4238), .B(n4239), .Z(n4236) );
  AND U7390 ( .A(a[81]), .B(b[23]), .Z(n4235) );
  XOR U7391 ( .A(n4240), .B(n4057), .Z(n4059) );
  XOR U7392 ( .A(n4241), .B(n4242), .Z(n4057) );
  AND U7393 ( .A(n4243), .B(n4244), .Z(n4241) );
  AND U7394 ( .A(a[82]), .B(b[22]), .Z(n4240) );
  XOR U7395 ( .A(n4245), .B(n4062), .Z(n4064) );
  XOR U7396 ( .A(n4246), .B(n4247), .Z(n4062) );
  AND U7397 ( .A(n4248), .B(n4249), .Z(n4246) );
  AND U7398 ( .A(a[83]), .B(b[21]), .Z(n4245) );
  XOR U7399 ( .A(n4250), .B(n4067), .Z(n4069) );
  XOR U7400 ( .A(n4251), .B(n4252), .Z(n4067) );
  AND U7401 ( .A(n4253), .B(n4254), .Z(n4251) );
  AND U7402 ( .A(a[84]), .B(b[20]), .Z(n4250) );
  XOR U7403 ( .A(n4255), .B(n4072), .Z(n4074) );
  XOR U7404 ( .A(n4256), .B(n4257), .Z(n4072) );
  AND U7405 ( .A(n4258), .B(n4259), .Z(n4256) );
  AND U7406 ( .A(a[85]), .B(b[19]), .Z(n4255) );
  XOR U7407 ( .A(n4260), .B(n4077), .Z(n4079) );
  XOR U7408 ( .A(n4261), .B(n4262), .Z(n4077) );
  AND U7409 ( .A(n4263), .B(n4264), .Z(n4261) );
  AND U7410 ( .A(a[86]), .B(b[18]), .Z(n4260) );
  XOR U7411 ( .A(n4265), .B(n4082), .Z(n4084) );
  XOR U7412 ( .A(n4266), .B(n4267), .Z(n4082) );
  AND U7413 ( .A(n4268), .B(n4269), .Z(n4266) );
  AND U7414 ( .A(a[87]), .B(b[17]), .Z(n4265) );
  XOR U7415 ( .A(n4270), .B(n4087), .Z(n4089) );
  XOR U7416 ( .A(n4271), .B(n4272), .Z(n4087) );
  AND U7417 ( .A(n4273), .B(n4274), .Z(n4271) );
  AND U7418 ( .A(a[88]), .B(b[16]), .Z(n4270) );
  XOR U7419 ( .A(n4275), .B(n4092), .Z(n4094) );
  XOR U7420 ( .A(n4276), .B(n4277), .Z(n4092) );
  AND U7421 ( .A(n4278), .B(n4279), .Z(n4276) );
  AND U7422 ( .A(a[89]), .B(b[15]), .Z(n4275) );
  XOR U7423 ( .A(n4280), .B(n4097), .Z(n4099) );
  XOR U7424 ( .A(n4281), .B(n4282), .Z(n4097) );
  AND U7425 ( .A(n4283), .B(n4284), .Z(n4281) );
  AND U7426 ( .A(a[90]), .B(b[14]), .Z(n4280) );
  XOR U7427 ( .A(n4285), .B(n4102), .Z(n4104) );
  XOR U7428 ( .A(n4286), .B(n4287), .Z(n4102) );
  AND U7429 ( .A(n4288), .B(n4289), .Z(n4286) );
  AND U7430 ( .A(a[91]), .B(b[13]), .Z(n4285) );
  XOR U7431 ( .A(n4290), .B(n4107), .Z(n4109) );
  XOR U7432 ( .A(n4291), .B(n4292), .Z(n4107) );
  AND U7433 ( .A(n4293), .B(n4294), .Z(n4291) );
  AND U7434 ( .A(a[92]), .B(b[12]), .Z(n4290) );
  XOR U7435 ( .A(n4295), .B(n4112), .Z(n4114) );
  XOR U7436 ( .A(n4296), .B(n4297), .Z(n4112) );
  AND U7437 ( .A(n4298), .B(n4299), .Z(n4296) );
  AND U7438 ( .A(a[93]), .B(b[11]), .Z(n4295) );
  XOR U7439 ( .A(n4300), .B(n4117), .Z(n4119) );
  XOR U7440 ( .A(n4301), .B(n4302), .Z(n4117) );
  AND U7441 ( .A(n4303), .B(n4304), .Z(n4301) );
  AND U7442 ( .A(a[94]), .B(b[10]), .Z(n4300) );
  XOR U7443 ( .A(n4305), .B(n4122), .Z(n4124) );
  XOR U7444 ( .A(n4306), .B(n4307), .Z(n4122) );
  AND U7445 ( .A(n4308), .B(n4309), .Z(n4306) );
  AND U7446 ( .A(b[9]), .B(a[95]), .Z(n4305) );
  XOR U7447 ( .A(n4310), .B(n4127), .Z(n4129) );
  XOR U7448 ( .A(n4311), .B(n4312), .Z(n4127) );
  AND U7449 ( .A(n4313), .B(n4314), .Z(n4311) );
  AND U7450 ( .A(b[8]), .B(a[96]), .Z(n4310) );
  XOR U7451 ( .A(n4315), .B(n4132), .Z(n4134) );
  XOR U7452 ( .A(n4316), .B(n4317), .Z(n4132) );
  AND U7453 ( .A(n4318), .B(n4319), .Z(n4316) );
  AND U7454 ( .A(b[7]), .B(a[97]), .Z(n4315) );
  XOR U7455 ( .A(n4320), .B(n4137), .Z(n4139) );
  XOR U7456 ( .A(n4321), .B(n4322), .Z(n4137) );
  AND U7457 ( .A(n4323), .B(n4324), .Z(n4321) );
  AND U7458 ( .A(b[6]), .B(a[98]), .Z(n4320) );
  XOR U7459 ( .A(n4325), .B(n4142), .Z(n4144) );
  XOR U7460 ( .A(n4326), .B(n4327), .Z(n4142) );
  AND U7461 ( .A(n4328), .B(n4329), .Z(n4326) );
  AND U7462 ( .A(b[5]), .B(a[99]), .Z(n4325) );
  XOR U7463 ( .A(n4330), .B(n4147), .Z(n4149) );
  XOR U7464 ( .A(n4331), .B(n4332), .Z(n4147) );
  AND U7465 ( .A(n4333), .B(n4334), .Z(n4331) );
  AND U7466 ( .A(b[4]), .B(a[100]), .Z(n4330) );
  XNOR U7467 ( .A(n4335), .B(n4336), .Z(n4161) );
  NANDN U7468 ( .A(n4337), .B(n4338), .Z(n4336) );
  XOR U7469 ( .A(n4339), .B(n4152), .Z(n4154) );
  XNOR U7470 ( .A(n4340), .B(n4341), .Z(n4152) );
  AND U7471 ( .A(n4342), .B(n4343), .Z(n4340) );
  AND U7472 ( .A(b[3]), .B(a[101]), .Z(n4339) );
  NAND U7473 ( .A(a[104]), .B(b[0]), .Z(n3990) );
  XOR U7474 ( .A(n4344), .B(n4345), .Z(swire[103]) );
  XOR U7475 ( .A(n4170), .B(n4171), .Z(n4346) );
  XNOR U7476 ( .A(n4337), .B(n4338), .Z(n4171) );
  XOR U7477 ( .A(n4335), .B(n4347), .Z(n4338) );
  NAND U7478 ( .A(b[1]), .B(a[102]), .Z(n4347) );
  XOR U7479 ( .A(n4343), .B(n4348), .Z(n4337) );
  XOR U7480 ( .A(n4335), .B(n4342), .Z(n4348) );
  XNOR U7481 ( .A(n4349), .B(n4341), .Z(n4342) );
  AND U7482 ( .A(b[2]), .B(a[101]), .Z(n4349) );
  NANDN U7483 ( .A(n4350), .B(n4351), .Z(n4335) );
  XOR U7484 ( .A(n4341), .B(n4333), .Z(n4352) );
  XNOR U7485 ( .A(n4332), .B(n4328), .Z(n4353) );
  XNOR U7486 ( .A(n4327), .B(n4323), .Z(n4354) );
  XNOR U7487 ( .A(n4322), .B(n4318), .Z(n4355) );
  XNOR U7488 ( .A(n4317), .B(n4313), .Z(n4356) );
  XNOR U7489 ( .A(n4312), .B(n4308), .Z(n4357) );
  XNOR U7490 ( .A(n4307), .B(n4303), .Z(n4358) );
  XNOR U7491 ( .A(n4302), .B(n4298), .Z(n4359) );
  XNOR U7492 ( .A(n4297), .B(n4293), .Z(n4360) );
  XNOR U7493 ( .A(n4292), .B(n4288), .Z(n4361) );
  XNOR U7494 ( .A(n4287), .B(n4283), .Z(n4362) );
  XNOR U7495 ( .A(n4282), .B(n4278), .Z(n4363) );
  XNOR U7496 ( .A(n4277), .B(n4273), .Z(n4364) );
  XNOR U7497 ( .A(n4272), .B(n4268), .Z(n4365) );
  XNOR U7498 ( .A(n4267), .B(n4263), .Z(n4366) );
  XNOR U7499 ( .A(n4262), .B(n4258), .Z(n4367) );
  XNOR U7500 ( .A(n4257), .B(n4253), .Z(n4368) );
  XNOR U7501 ( .A(n4252), .B(n4248), .Z(n4369) );
  XNOR U7502 ( .A(n4247), .B(n4243), .Z(n4370) );
  XNOR U7503 ( .A(n4242), .B(n4238), .Z(n4371) );
  XNOR U7504 ( .A(n4237), .B(n4233), .Z(n4372) );
  XNOR U7505 ( .A(n4232), .B(n4228), .Z(n4373) );
  XNOR U7506 ( .A(n4227), .B(n4223), .Z(n4374) );
  XNOR U7507 ( .A(n4222), .B(n4218), .Z(n4375) );
  XNOR U7508 ( .A(n4217), .B(n4213), .Z(n4376) );
  XOR U7509 ( .A(n4212), .B(n4209), .Z(n4377) );
  XOR U7510 ( .A(n4378), .B(n4379), .Z(n4209) );
  XOR U7511 ( .A(n4207), .B(n4380), .Z(n4379) );
  XOR U7512 ( .A(n4381), .B(n4382), .Z(n4380) );
  XOR U7513 ( .A(n4383), .B(n4384), .Z(n4382) );
  NAND U7514 ( .A(a[73]), .B(b[30]), .Z(n4384) );
  AND U7515 ( .A(a[72]), .B(b[31]), .Z(n4383) );
  XOR U7516 ( .A(n4385), .B(n4381), .Z(n4378) );
  XOR U7517 ( .A(n4386), .B(n4387), .Z(n4381) );
  ANDN U7518 ( .B(n4388), .A(n4389), .Z(n4386) );
  AND U7519 ( .A(a[74]), .B(b[29]), .Z(n4385) );
  XOR U7520 ( .A(n4390), .B(n4207), .Z(n4208) );
  XOR U7521 ( .A(n4391), .B(n4392), .Z(n4207) );
  AND U7522 ( .A(n4393), .B(n4394), .Z(n4391) );
  AND U7523 ( .A(a[75]), .B(b[28]), .Z(n4390) );
  XOR U7524 ( .A(n4395), .B(n4212), .Z(n4214) );
  XOR U7525 ( .A(n4396), .B(n4397), .Z(n4212) );
  AND U7526 ( .A(n4398), .B(n4399), .Z(n4396) );
  AND U7527 ( .A(a[76]), .B(b[27]), .Z(n4395) );
  XOR U7528 ( .A(n4400), .B(n4217), .Z(n4219) );
  XOR U7529 ( .A(n4401), .B(n4402), .Z(n4217) );
  AND U7530 ( .A(n4403), .B(n4404), .Z(n4401) );
  AND U7531 ( .A(a[77]), .B(b[26]), .Z(n4400) );
  XOR U7532 ( .A(n4405), .B(n4222), .Z(n4224) );
  XOR U7533 ( .A(n4406), .B(n4407), .Z(n4222) );
  AND U7534 ( .A(n4408), .B(n4409), .Z(n4406) );
  AND U7535 ( .A(a[78]), .B(b[25]), .Z(n4405) );
  XOR U7536 ( .A(n4410), .B(n4227), .Z(n4229) );
  XOR U7537 ( .A(n4411), .B(n4412), .Z(n4227) );
  AND U7538 ( .A(n4413), .B(n4414), .Z(n4411) );
  AND U7539 ( .A(a[79]), .B(b[24]), .Z(n4410) );
  XOR U7540 ( .A(n4415), .B(n4232), .Z(n4234) );
  XOR U7541 ( .A(n4416), .B(n4417), .Z(n4232) );
  AND U7542 ( .A(n4418), .B(n4419), .Z(n4416) );
  AND U7543 ( .A(a[80]), .B(b[23]), .Z(n4415) );
  XOR U7544 ( .A(n4420), .B(n4237), .Z(n4239) );
  XOR U7545 ( .A(n4421), .B(n4422), .Z(n4237) );
  AND U7546 ( .A(n4423), .B(n4424), .Z(n4421) );
  AND U7547 ( .A(a[81]), .B(b[22]), .Z(n4420) );
  XOR U7548 ( .A(n4425), .B(n4242), .Z(n4244) );
  XOR U7549 ( .A(n4426), .B(n4427), .Z(n4242) );
  AND U7550 ( .A(n4428), .B(n4429), .Z(n4426) );
  AND U7551 ( .A(a[82]), .B(b[21]), .Z(n4425) );
  XOR U7552 ( .A(n4430), .B(n4247), .Z(n4249) );
  XOR U7553 ( .A(n4431), .B(n4432), .Z(n4247) );
  AND U7554 ( .A(n4433), .B(n4434), .Z(n4431) );
  AND U7555 ( .A(a[83]), .B(b[20]), .Z(n4430) );
  XOR U7556 ( .A(n4435), .B(n4252), .Z(n4254) );
  XOR U7557 ( .A(n4436), .B(n4437), .Z(n4252) );
  AND U7558 ( .A(n4438), .B(n4439), .Z(n4436) );
  AND U7559 ( .A(a[84]), .B(b[19]), .Z(n4435) );
  XOR U7560 ( .A(n4440), .B(n4257), .Z(n4259) );
  XOR U7561 ( .A(n4441), .B(n4442), .Z(n4257) );
  AND U7562 ( .A(n4443), .B(n4444), .Z(n4441) );
  AND U7563 ( .A(a[85]), .B(b[18]), .Z(n4440) );
  XOR U7564 ( .A(n4445), .B(n4262), .Z(n4264) );
  XOR U7565 ( .A(n4446), .B(n4447), .Z(n4262) );
  AND U7566 ( .A(n4448), .B(n4449), .Z(n4446) );
  AND U7567 ( .A(a[86]), .B(b[17]), .Z(n4445) );
  XOR U7568 ( .A(n4450), .B(n4267), .Z(n4269) );
  XOR U7569 ( .A(n4451), .B(n4452), .Z(n4267) );
  AND U7570 ( .A(n4453), .B(n4454), .Z(n4451) );
  AND U7571 ( .A(a[87]), .B(b[16]), .Z(n4450) );
  XOR U7572 ( .A(n4455), .B(n4272), .Z(n4274) );
  XOR U7573 ( .A(n4456), .B(n4457), .Z(n4272) );
  AND U7574 ( .A(n4458), .B(n4459), .Z(n4456) );
  AND U7575 ( .A(a[88]), .B(b[15]), .Z(n4455) );
  XOR U7576 ( .A(n4460), .B(n4277), .Z(n4279) );
  XOR U7577 ( .A(n4461), .B(n4462), .Z(n4277) );
  AND U7578 ( .A(n4463), .B(n4464), .Z(n4461) );
  AND U7579 ( .A(a[89]), .B(b[14]), .Z(n4460) );
  XOR U7580 ( .A(n4465), .B(n4282), .Z(n4284) );
  XOR U7581 ( .A(n4466), .B(n4467), .Z(n4282) );
  AND U7582 ( .A(n4468), .B(n4469), .Z(n4466) );
  AND U7583 ( .A(a[90]), .B(b[13]), .Z(n4465) );
  XOR U7584 ( .A(n4470), .B(n4287), .Z(n4289) );
  XOR U7585 ( .A(n4471), .B(n4472), .Z(n4287) );
  AND U7586 ( .A(n4473), .B(n4474), .Z(n4471) );
  AND U7587 ( .A(a[91]), .B(b[12]), .Z(n4470) );
  XOR U7588 ( .A(n4475), .B(n4292), .Z(n4294) );
  XOR U7589 ( .A(n4476), .B(n4477), .Z(n4292) );
  AND U7590 ( .A(n4478), .B(n4479), .Z(n4476) );
  AND U7591 ( .A(a[92]), .B(b[11]), .Z(n4475) );
  XOR U7592 ( .A(n4480), .B(n4297), .Z(n4299) );
  XOR U7593 ( .A(n4481), .B(n4482), .Z(n4297) );
  AND U7594 ( .A(n4483), .B(n4484), .Z(n4481) );
  AND U7595 ( .A(a[93]), .B(b[10]), .Z(n4480) );
  XOR U7596 ( .A(n4485), .B(n4302), .Z(n4304) );
  XOR U7597 ( .A(n4486), .B(n4487), .Z(n4302) );
  AND U7598 ( .A(n4488), .B(n4489), .Z(n4486) );
  AND U7599 ( .A(a[94]), .B(b[9]), .Z(n4485) );
  XOR U7600 ( .A(n4490), .B(n4307), .Z(n4309) );
  XOR U7601 ( .A(n4491), .B(n4492), .Z(n4307) );
  AND U7602 ( .A(n4493), .B(n4494), .Z(n4491) );
  AND U7603 ( .A(b[8]), .B(a[95]), .Z(n4490) );
  XOR U7604 ( .A(n4495), .B(n4312), .Z(n4314) );
  XOR U7605 ( .A(n4496), .B(n4497), .Z(n4312) );
  AND U7606 ( .A(n4498), .B(n4499), .Z(n4496) );
  AND U7607 ( .A(b[7]), .B(a[96]), .Z(n4495) );
  XOR U7608 ( .A(n4500), .B(n4317), .Z(n4319) );
  XOR U7609 ( .A(n4501), .B(n4502), .Z(n4317) );
  AND U7610 ( .A(n4503), .B(n4504), .Z(n4501) );
  AND U7611 ( .A(b[6]), .B(a[97]), .Z(n4500) );
  XOR U7612 ( .A(n4505), .B(n4322), .Z(n4324) );
  XOR U7613 ( .A(n4506), .B(n4507), .Z(n4322) );
  AND U7614 ( .A(n4508), .B(n4509), .Z(n4506) );
  AND U7615 ( .A(b[5]), .B(a[98]), .Z(n4505) );
  XOR U7616 ( .A(n4510), .B(n4327), .Z(n4329) );
  XOR U7617 ( .A(n4511), .B(n4512), .Z(n4327) );
  AND U7618 ( .A(n4513), .B(n4514), .Z(n4511) );
  AND U7619 ( .A(b[4]), .B(a[99]), .Z(n4510) );
  XNOR U7620 ( .A(n4515), .B(n4516), .Z(n4341) );
  NANDN U7621 ( .A(n4517), .B(n4518), .Z(n4516) );
  XOR U7622 ( .A(n4519), .B(n4332), .Z(n4334) );
  XNOR U7623 ( .A(n4520), .B(n4521), .Z(n4332) );
  AND U7624 ( .A(n4522), .B(n4523), .Z(n4520) );
  AND U7625 ( .A(b[3]), .B(a[100]), .Z(n4519) );
  NAND U7626 ( .A(a[103]), .B(b[0]), .Z(n4170) );
  XOR U7627 ( .A(n4524), .B(n4525), .Z(swire[102]) );
  XOR U7628 ( .A(n4350), .B(n4351), .Z(n4526) );
  XNOR U7629 ( .A(n4517), .B(n4518), .Z(n4351) );
  XOR U7630 ( .A(n4515), .B(n4527), .Z(n4518) );
  NAND U7631 ( .A(b[1]), .B(a[101]), .Z(n4527) );
  XOR U7632 ( .A(n4523), .B(n4528), .Z(n4517) );
  XOR U7633 ( .A(n4515), .B(n4522), .Z(n4528) );
  XNOR U7634 ( .A(n4529), .B(n4521), .Z(n4522) );
  AND U7635 ( .A(b[2]), .B(a[100]), .Z(n4529) );
  NANDN U7636 ( .A(n4530), .B(n4531), .Z(n4515) );
  XOR U7637 ( .A(n4521), .B(n4513), .Z(n4532) );
  XNOR U7638 ( .A(n4512), .B(n4508), .Z(n4533) );
  XNOR U7639 ( .A(n4507), .B(n4503), .Z(n4534) );
  XNOR U7640 ( .A(n4502), .B(n4498), .Z(n4535) );
  XNOR U7641 ( .A(n4497), .B(n4493), .Z(n4536) );
  XNOR U7642 ( .A(n4492), .B(n4488), .Z(n4537) );
  XNOR U7643 ( .A(n4487), .B(n4483), .Z(n4538) );
  XNOR U7644 ( .A(n4482), .B(n4478), .Z(n4539) );
  XNOR U7645 ( .A(n4477), .B(n4473), .Z(n4540) );
  XNOR U7646 ( .A(n4472), .B(n4468), .Z(n4541) );
  XNOR U7647 ( .A(n4467), .B(n4463), .Z(n4542) );
  XNOR U7648 ( .A(n4462), .B(n4458), .Z(n4543) );
  XNOR U7649 ( .A(n4457), .B(n4453), .Z(n4544) );
  XNOR U7650 ( .A(n4452), .B(n4448), .Z(n4545) );
  XNOR U7651 ( .A(n4447), .B(n4443), .Z(n4546) );
  XNOR U7652 ( .A(n4442), .B(n4438), .Z(n4547) );
  XNOR U7653 ( .A(n4437), .B(n4433), .Z(n4548) );
  XNOR U7654 ( .A(n4432), .B(n4428), .Z(n4549) );
  XNOR U7655 ( .A(n4427), .B(n4423), .Z(n4550) );
  XNOR U7656 ( .A(n4422), .B(n4418), .Z(n4551) );
  XNOR U7657 ( .A(n4417), .B(n4413), .Z(n4552) );
  XNOR U7658 ( .A(n4412), .B(n4408), .Z(n4553) );
  XNOR U7659 ( .A(n4407), .B(n4403), .Z(n4554) );
  XNOR U7660 ( .A(n4402), .B(n4398), .Z(n4555) );
  XNOR U7661 ( .A(n4397), .B(n4393), .Z(n4556) );
  XOR U7662 ( .A(n4392), .B(n4389), .Z(n4557) );
  XOR U7663 ( .A(n4558), .B(n4559), .Z(n4389) );
  XOR U7664 ( .A(n4387), .B(n4560), .Z(n4559) );
  XOR U7665 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U7666 ( .A(n4563), .B(n4564), .Z(n4562) );
  NAND U7667 ( .A(a[72]), .B(b[30]), .Z(n4564) );
  AND U7668 ( .A(a[71]), .B(b[31]), .Z(n4563) );
  XOR U7669 ( .A(n4565), .B(n4561), .Z(n4558) );
  XOR U7670 ( .A(n4566), .B(n4567), .Z(n4561) );
  ANDN U7671 ( .B(n4568), .A(n4569), .Z(n4566) );
  AND U7672 ( .A(a[73]), .B(b[29]), .Z(n4565) );
  XOR U7673 ( .A(n4570), .B(n4387), .Z(n4388) );
  XOR U7674 ( .A(n4571), .B(n4572), .Z(n4387) );
  AND U7675 ( .A(n4573), .B(n4574), .Z(n4571) );
  AND U7676 ( .A(a[74]), .B(b[28]), .Z(n4570) );
  XOR U7677 ( .A(n4575), .B(n4392), .Z(n4394) );
  XOR U7678 ( .A(n4576), .B(n4577), .Z(n4392) );
  AND U7679 ( .A(n4578), .B(n4579), .Z(n4576) );
  AND U7680 ( .A(a[75]), .B(b[27]), .Z(n4575) );
  XOR U7681 ( .A(n4580), .B(n4397), .Z(n4399) );
  XOR U7682 ( .A(n4581), .B(n4582), .Z(n4397) );
  AND U7683 ( .A(n4583), .B(n4584), .Z(n4581) );
  AND U7684 ( .A(a[76]), .B(b[26]), .Z(n4580) );
  XOR U7685 ( .A(n4585), .B(n4402), .Z(n4404) );
  XOR U7686 ( .A(n4586), .B(n4587), .Z(n4402) );
  AND U7687 ( .A(n4588), .B(n4589), .Z(n4586) );
  AND U7688 ( .A(a[77]), .B(b[25]), .Z(n4585) );
  XOR U7689 ( .A(n4590), .B(n4407), .Z(n4409) );
  XOR U7690 ( .A(n4591), .B(n4592), .Z(n4407) );
  AND U7691 ( .A(n4593), .B(n4594), .Z(n4591) );
  AND U7692 ( .A(a[78]), .B(b[24]), .Z(n4590) );
  XOR U7693 ( .A(n4595), .B(n4412), .Z(n4414) );
  XOR U7694 ( .A(n4596), .B(n4597), .Z(n4412) );
  AND U7695 ( .A(n4598), .B(n4599), .Z(n4596) );
  AND U7696 ( .A(a[79]), .B(b[23]), .Z(n4595) );
  XOR U7697 ( .A(n4600), .B(n4417), .Z(n4419) );
  XOR U7698 ( .A(n4601), .B(n4602), .Z(n4417) );
  AND U7699 ( .A(n4603), .B(n4604), .Z(n4601) );
  AND U7700 ( .A(a[80]), .B(b[22]), .Z(n4600) );
  XOR U7701 ( .A(n4605), .B(n4422), .Z(n4424) );
  XOR U7702 ( .A(n4606), .B(n4607), .Z(n4422) );
  AND U7703 ( .A(n4608), .B(n4609), .Z(n4606) );
  AND U7704 ( .A(a[81]), .B(b[21]), .Z(n4605) );
  XOR U7705 ( .A(n4610), .B(n4427), .Z(n4429) );
  XOR U7706 ( .A(n4611), .B(n4612), .Z(n4427) );
  AND U7707 ( .A(n4613), .B(n4614), .Z(n4611) );
  AND U7708 ( .A(a[82]), .B(b[20]), .Z(n4610) );
  XOR U7709 ( .A(n4615), .B(n4432), .Z(n4434) );
  XOR U7710 ( .A(n4616), .B(n4617), .Z(n4432) );
  AND U7711 ( .A(n4618), .B(n4619), .Z(n4616) );
  AND U7712 ( .A(a[83]), .B(b[19]), .Z(n4615) );
  XOR U7713 ( .A(n4620), .B(n4437), .Z(n4439) );
  XOR U7714 ( .A(n4621), .B(n4622), .Z(n4437) );
  AND U7715 ( .A(n4623), .B(n4624), .Z(n4621) );
  AND U7716 ( .A(a[84]), .B(b[18]), .Z(n4620) );
  XOR U7717 ( .A(n4625), .B(n4442), .Z(n4444) );
  XOR U7718 ( .A(n4626), .B(n4627), .Z(n4442) );
  AND U7719 ( .A(n4628), .B(n4629), .Z(n4626) );
  AND U7720 ( .A(a[85]), .B(b[17]), .Z(n4625) );
  XOR U7721 ( .A(n4630), .B(n4447), .Z(n4449) );
  XOR U7722 ( .A(n4631), .B(n4632), .Z(n4447) );
  AND U7723 ( .A(n4633), .B(n4634), .Z(n4631) );
  AND U7724 ( .A(a[86]), .B(b[16]), .Z(n4630) );
  XOR U7725 ( .A(n4635), .B(n4452), .Z(n4454) );
  XOR U7726 ( .A(n4636), .B(n4637), .Z(n4452) );
  AND U7727 ( .A(n4638), .B(n4639), .Z(n4636) );
  AND U7728 ( .A(a[87]), .B(b[15]), .Z(n4635) );
  XOR U7729 ( .A(n4640), .B(n4457), .Z(n4459) );
  XOR U7730 ( .A(n4641), .B(n4642), .Z(n4457) );
  AND U7731 ( .A(n4643), .B(n4644), .Z(n4641) );
  AND U7732 ( .A(a[88]), .B(b[14]), .Z(n4640) );
  XOR U7733 ( .A(n4645), .B(n4462), .Z(n4464) );
  XOR U7734 ( .A(n4646), .B(n4647), .Z(n4462) );
  AND U7735 ( .A(n4648), .B(n4649), .Z(n4646) );
  AND U7736 ( .A(a[89]), .B(b[13]), .Z(n4645) );
  XOR U7737 ( .A(n4650), .B(n4467), .Z(n4469) );
  XOR U7738 ( .A(n4651), .B(n4652), .Z(n4467) );
  AND U7739 ( .A(n4653), .B(n4654), .Z(n4651) );
  AND U7740 ( .A(a[90]), .B(b[12]), .Z(n4650) );
  XOR U7741 ( .A(n4655), .B(n4472), .Z(n4474) );
  XOR U7742 ( .A(n4656), .B(n4657), .Z(n4472) );
  AND U7743 ( .A(n4658), .B(n4659), .Z(n4656) );
  AND U7744 ( .A(a[91]), .B(b[11]), .Z(n4655) );
  XOR U7745 ( .A(n4660), .B(n4477), .Z(n4479) );
  XOR U7746 ( .A(n4661), .B(n4662), .Z(n4477) );
  AND U7747 ( .A(n4663), .B(n4664), .Z(n4661) );
  AND U7748 ( .A(a[92]), .B(b[10]), .Z(n4660) );
  XOR U7749 ( .A(n4665), .B(n4482), .Z(n4484) );
  XOR U7750 ( .A(n4666), .B(n4667), .Z(n4482) );
  AND U7751 ( .A(n4668), .B(n4669), .Z(n4666) );
  AND U7752 ( .A(a[93]), .B(b[9]), .Z(n4665) );
  XOR U7753 ( .A(n4670), .B(n4487), .Z(n4489) );
  XOR U7754 ( .A(n4671), .B(n4672), .Z(n4487) );
  AND U7755 ( .A(n4673), .B(n4674), .Z(n4671) );
  AND U7756 ( .A(a[94]), .B(b[8]), .Z(n4670) );
  XOR U7757 ( .A(n4675), .B(n4492), .Z(n4494) );
  XOR U7758 ( .A(n4676), .B(n4677), .Z(n4492) );
  AND U7759 ( .A(n4678), .B(n4679), .Z(n4676) );
  AND U7760 ( .A(b[7]), .B(a[95]), .Z(n4675) );
  XOR U7761 ( .A(n4680), .B(n4497), .Z(n4499) );
  XOR U7762 ( .A(n4681), .B(n4682), .Z(n4497) );
  AND U7763 ( .A(n4683), .B(n4684), .Z(n4681) );
  AND U7764 ( .A(b[6]), .B(a[96]), .Z(n4680) );
  XOR U7765 ( .A(n4685), .B(n4502), .Z(n4504) );
  XOR U7766 ( .A(n4686), .B(n4687), .Z(n4502) );
  AND U7767 ( .A(n4688), .B(n4689), .Z(n4686) );
  AND U7768 ( .A(b[5]), .B(a[97]), .Z(n4685) );
  XOR U7769 ( .A(n4690), .B(n4507), .Z(n4509) );
  XOR U7770 ( .A(n4691), .B(n4692), .Z(n4507) );
  AND U7771 ( .A(n4693), .B(n4694), .Z(n4691) );
  AND U7772 ( .A(b[4]), .B(a[98]), .Z(n4690) );
  XNOR U7773 ( .A(n4695), .B(n4696), .Z(n4521) );
  NANDN U7774 ( .A(n4697), .B(n4698), .Z(n4696) );
  XOR U7775 ( .A(n4699), .B(n4512), .Z(n4514) );
  XNOR U7776 ( .A(n4700), .B(n4701), .Z(n4512) );
  AND U7777 ( .A(n4702), .B(n4703), .Z(n4700) );
  AND U7778 ( .A(b[3]), .B(a[99]), .Z(n4699) );
  NAND U7779 ( .A(a[102]), .B(b[0]), .Z(n4350) );
  XOR U7780 ( .A(n4704), .B(n4705), .Z(swire[101]) );
  XOR U7781 ( .A(n4530), .B(n4531), .Z(n4706) );
  XNOR U7782 ( .A(n4697), .B(n4698), .Z(n4531) );
  XOR U7783 ( .A(n4695), .B(n4707), .Z(n4698) );
  NAND U7784 ( .A(b[1]), .B(a[100]), .Z(n4707) );
  XOR U7785 ( .A(n4703), .B(n4708), .Z(n4697) );
  XOR U7786 ( .A(n4695), .B(n4702), .Z(n4708) );
  XNOR U7787 ( .A(n4709), .B(n4701), .Z(n4702) );
  AND U7788 ( .A(b[2]), .B(a[99]), .Z(n4709) );
  NANDN U7789 ( .A(n4710), .B(n4711), .Z(n4695) );
  XOR U7790 ( .A(n4701), .B(n4693), .Z(n4712) );
  XNOR U7791 ( .A(n4692), .B(n4688), .Z(n4713) );
  XNOR U7792 ( .A(n4687), .B(n4683), .Z(n4714) );
  XNOR U7793 ( .A(n4682), .B(n4678), .Z(n4715) );
  XNOR U7794 ( .A(n4677), .B(n4673), .Z(n4716) );
  XNOR U7795 ( .A(n4672), .B(n4668), .Z(n4717) );
  XNOR U7796 ( .A(n4667), .B(n4663), .Z(n4718) );
  XNOR U7797 ( .A(n4662), .B(n4658), .Z(n4719) );
  XNOR U7798 ( .A(n4657), .B(n4653), .Z(n4720) );
  XNOR U7799 ( .A(n4652), .B(n4648), .Z(n4721) );
  XNOR U7800 ( .A(n4647), .B(n4643), .Z(n4722) );
  XNOR U7801 ( .A(n4642), .B(n4638), .Z(n4723) );
  XNOR U7802 ( .A(n4637), .B(n4633), .Z(n4724) );
  XNOR U7803 ( .A(n4632), .B(n4628), .Z(n4725) );
  XNOR U7804 ( .A(n4627), .B(n4623), .Z(n4726) );
  XNOR U7805 ( .A(n4622), .B(n4618), .Z(n4727) );
  XNOR U7806 ( .A(n4617), .B(n4613), .Z(n4728) );
  XNOR U7807 ( .A(n4612), .B(n4608), .Z(n4729) );
  XNOR U7808 ( .A(n4607), .B(n4603), .Z(n4730) );
  XNOR U7809 ( .A(n4602), .B(n4598), .Z(n4731) );
  XNOR U7810 ( .A(n4597), .B(n4593), .Z(n4732) );
  XNOR U7811 ( .A(n4592), .B(n4588), .Z(n4733) );
  XNOR U7812 ( .A(n4587), .B(n4583), .Z(n4734) );
  XNOR U7813 ( .A(n4582), .B(n4578), .Z(n4735) );
  XNOR U7814 ( .A(n4577), .B(n4573), .Z(n4736) );
  XOR U7815 ( .A(n4572), .B(n4569), .Z(n4737) );
  XOR U7816 ( .A(n4738), .B(n4739), .Z(n4569) );
  XOR U7817 ( .A(n4567), .B(n4740), .Z(n4739) );
  XOR U7818 ( .A(n4741), .B(n4742), .Z(n4740) );
  XOR U7819 ( .A(n4743), .B(n4744), .Z(n4742) );
  NAND U7820 ( .A(a[71]), .B(b[30]), .Z(n4744) );
  AND U7821 ( .A(a[70]), .B(b[31]), .Z(n4743) );
  XOR U7822 ( .A(n4745), .B(n4741), .Z(n4738) );
  XOR U7823 ( .A(n4746), .B(n4747), .Z(n4741) );
  ANDN U7824 ( .B(n4748), .A(n4749), .Z(n4746) );
  AND U7825 ( .A(a[72]), .B(b[29]), .Z(n4745) );
  XOR U7826 ( .A(n4750), .B(n4567), .Z(n4568) );
  XOR U7827 ( .A(n4751), .B(n4752), .Z(n4567) );
  AND U7828 ( .A(n4753), .B(n4754), .Z(n4751) );
  AND U7829 ( .A(a[73]), .B(b[28]), .Z(n4750) );
  XOR U7830 ( .A(n4755), .B(n4572), .Z(n4574) );
  XOR U7831 ( .A(n4756), .B(n4757), .Z(n4572) );
  AND U7832 ( .A(n4758), .B(n4759), .Z(n4756) );
  AND U7833 ( .A(a[74]), .B(b[27]), .Z(n4755) );
  XOR U7834 ( .A(n4760), .B(n4577), .Z(n4579) );
  XOR U7835 ( .A(n4761), .B(n4762), .Z(n4577) );
  AND U7836 ( .A(n4763), .B(n4764), .Z(n4761) );
  AND U7837 ( .A(a[75]), .B(b[26]), .Z(n4760) );
  XOR U7838 ( .A(n4765), .B(n4582), .Z(n4584) );
  XOR U7839 ( .A(n4766), .B(n4767), .Z(n4582) );
  AND U7840 ( .A(n4768), .B(n4769), .Z(n4766) );
  AND U7841 ( .A(a[76]), .B(b[25]), .Z(n4765) );
  XOR U7842 ( .A(n4770), .B(n4587), .Z(n4589) );
  XOR U7843 ( .A(n4771), .B(n4772), .Z(n4587) );
  AND U7844 ( .A(n4773), .B(n4774), .Z(n4771) );
  AND U7845 ( .A(a[77]), .B(b[24]), .Z(n4770) );
  XOR U7846 ( .A(n4775), .B(n4592), .Z(n4594) );
  XOR U7847 ( .A(n4776), .B(n4777), .Z(n4592) );
  AND U7848 ( .A(n4778), .B(n4779), .Z(n4776) );
  AND U7849 ( .A(a[78]), .B(b[23]), .Z(n4775) );
  XOR U7850 ( .A(n4780), .B(n4597), .Z(n4599) );
  XOR U7851 ( .A(n4781), .B(n4782), .Z(n4597) );
  AND U7852 ( .A(n4783), .B(n4784), .Z(n4781) );
  AND U7853 ( .A(a[79]), .B(b[22]), .Z(n4780) );
  XOR U7854 ( .A(n4785), .B(n4602), .Z(n4604) );
  XOR U7855 ( .A(n4786), .B(n4787), .Z(n4602) );
  AND U7856 ( .A(n4788), .B(n4789), .Z(n4786) );
  AND U7857 ( .A(a[80]), .B(b[21]), .Z(n4785) );
  XOR U7858 ( .A(n4790), .B(n4607), .Z(n4609) );
  XOR U7859 ( .A(n4791), .B(n4792), .Z(n4607) );
  AND U7860 ( .A(n4793), .B(n4794), .Z(n4791) );
  AND U7861 ( .A(a[81]), .B(b[20]), .Z(n4790) );
  XOR U7862 ( .A(n4795), .B(n4612), .Z(n4614) );
  XOR U7863 ( .A(n4796), .B(n4797), .Z(n4612) );
  AND U7864 ( .A(n4798), .B(n4799), .Z(n4796) );
  AND U7865 ( .A(a[82]), .B(b[19]), .Z(n4795) );
  XOR U7866 ( .A(n4800), .B(n4617), .Z(n4619) );
  XOR U7867 ( .A(n4801), .B(n4802), .Z(n4617) );
  AND U7868 ( .A(n4803), .B(n4804), .Z(n4801) );
  AND U7869 ( .A(a[83]), .B(b[18]), .Z(n4800) );
  XOR U7870 ( .A(n4805), .B(n4622), .Z(n4624) );
  XOR U7871 ( .A(n4806), .B(n4807), .Z(n4622) );
  AND U7872 ( .A(n4808), .B(n4809), .Z(n4806) );
  AND U7873 ( .A(a[84]), .B(b[17]), .Z(n4805) );
  XOR U7874 ( .A(n4810), .B(n4627), .Z(n4629) );
  XOR U7875 ( .A(n4811), .B(n4812), .Z(n4627) );
  AND U7876 ( .A(n4813), .B(n4814), .Z(n4811) );
  AND U7877 ( .A(a[85]), .B(b[16]), .Z(n4810) );
  XOR U7878 ( .A(n4815), .B(n4632), .Z(n4634) );
  XOR U7879 ( .A(n4816), .B(n4817), .Z(n4632) );
  AND U7880 ( .A(n4818), .B(n4819), .Z(n4816) );
  AND U7881 ( .A(a[86]), .B(b[15]), .Z(n4815) );
  XOR U7882 ( .A(n4820), .B(n4637), .Z(n4639) );
  XOR U7883 ( .A(n4821), .B(n4822), .Z(n4637) );
  AND U7884 ( .A(n4823), .B(n4824), .Z(n4821) );
  AND U7885 ( .A(a[87]), .B(b[14]), .Z(n4820) );
  XOR U7886 ( .A(n4825), .B(n4642), .Z(n4644) );
  XOR U7887 ( .A(n4826), .B(n4827), .Z(n4642) );
  AND U7888 ( .A(n4828), .B(n4829), .Z(n4826) );
  AND U7889 ( .A(a[88]), .B(b[13]), .Z(n4825) );
  XOR U7890 ( .A(n4830), .B(n4647), .Z(n4649) );
  XOR U7891 ( .A(n4831), .B(n4832), .Z(n4647) );
  AND U7892 ( .A(n4833), .B(n4834), .Z(n4831) );
  AND U7893 ( .A(a[89]), .B(b[12]), .Z(n4830) );
  XOR U7894 ( .A(n4835), .B(n4652), .Z(n4654) );
  XOR U7895 ( .A(n4836), .B(n4837), .Z(n4652) );
  AND U7896 ( .A(n4838), .B(n4839), .Z(n4836) );
  AND U7897 ( .A(a[90]), .B(b[11]), .Z(n4835) );
  XOR U7898 ( .A(n4840), .B(n4657), .Z(n4659) );
  XOR U7899 ( .A(n4841), .B(n4842), .Z(n4657) );
  AND U7900 ( .A(n4843), .B(n4844), .Z(n4841) );
  AND U7901 ( .A(a[91]), .B(b[10]), .Z(n4840) );
  XOR U7902 ( .A(n4845), .B(n4662), .Z(n4664) );
  XOR U7903 ( .A(n4846), .B(n4847), .Z(n4662) );
  AND U7904 ( .A(n4848), .B(n4849), .Z(n4846) );
  AND U7905 ( .A(a[92]), .B(b[9]), .Z(n4845) );
  XOR U7906 ( .A(n4850), .B(n4667), .Z(n4669) );
  XOR U7907 ( .A(n4851), .B(n4852), .Z(n4667) );
  AND U7908 ( .A(n4853), .B(n4854), .Z(n4851) );
  AND U7909 ( .A(a[93]), .B(b[8]), .Z(n4850) );
  XOR U7910 ( .A(n4855), .B(n4672), .Z(n4674) );
  XOR U7911 ( .A(n4856), .B(n4857), .Z(n4672) );
  AND U7912 ( .A(n4858), .B(n4859), .Z(n4856) );
  AND U7913 ( .A(a[94]), .B(b[7]), .Z(n4855) );
  XOR U7914 ( .A(n4860), .B(n4677), .Z(n4679) );
  XOR U7915 ( .A(n4861), .B(n4862), .Z(n4677) );
  AND U7916 ( .A(n4863), .B(n4864), .Z(n4861) );
  AND U7917 ( .A(b[6]), .B(a[95]), .Z(n4860) );
  XOR U7918 ( .A(n4865), .B(n4682), .Z(n4684) );
  XOR U7919 ( .A(n4866), .B(n4867), .Z(n4682) );
  AND U7920 ( .A(n4868), .B(n4869), .Z(n4866) );
  AND U7921 ( .A(b[5]), .B(a[96]), .Z(n4865) );
  XOR U7922 ( .A(n4870), .B(n4687), .Z(n4689) );
  XOR U7923 ( .A(n4871), .B(n4872), .Z(n4687) );
  AND U7924 ( .A(n4873), .B(n4874), .Z(n4871) );
  AND U7925 ( .A(b[4]), .B(a[97]), .Z(n4870) );
  XNOR U7926 ( .A(n4875), .B(n4876), .Z(n4701) );
  NANDN U7927 ( .A(n4877), .B(n4878), .Z(n4876) );
  XOR U7928 ( .A(n4879), .B(n4692), .Z(n4694) );
  XNOR U7929 ( .A(n4880), .B(n4881), .Z(n4692) );
  AND U7930 ( .A(n4882), .B(n4883), .Z(n4880) );
  AND U7931 ( .A(b[3]), .B(a[98]), .Z(n4879) );
  NAND U7932 ( .A(a[101]), .B(b[0]), .Z(n4530) );
  XOR U7933 ( .A(n4884), .B(n4885), .Z(swire[100]) );
  XOR U7934 ( .A(n4710), .B(n4711), .Z(n4886) );
  XNOR U7935 ( .A(n4877), .B(n4878), .Z(n4711) );
  XOR U7936 ( .A(n4875), .B(n4887), .Z(n4878) );
  NAND U7937 ( .A(b[1]), .B(a[99]), .Z(n4887) );
  XOR U7938 ( .A(n4883), .B(n4888), .Z(n4877) );
  XOR U7939 ( .A(n4875), .B(n4882), .Z(n4888) );
  XNOR U7940 ( .A(n4889), .B(n4881), .Z(n4882) );
  AND U7941 ( .A(b[2]), .B(a[98]), .Z(n4889) );
  OR U7942 ( .A(n4890), .B(n4891), .Z(n4875) );
  XOR U7943 ( .A(n4881), .B(n4873), .Z(n4892) );
  XNOR U7944 ( .A(n4872), .B(n4868), .Z(n4893) );
  XNOR U7945 ( .A(n4867), .B(n4863), .Z(n4894) );
  XNOR U7946 ( .A(n4862), .B(n4858), .Z(n4895) );
  XNOR U7947 ( .A(n4857), .B(n4853), .Z(n4896) );
  XNOR U7948 ( .A(n4852), .B(n4848), .Z(n4897) );
  XNOR U7949 ( .A(n4847), .B(n4843), .Z(n4898) );
  XNOR U7950 ( .A(n4842), .B(n4838), .Z(n4899) );
  XNOR U7951 ( .A(n4837), .B(n4833), .Z(n4900) );
  XNOR U7952 ( .A(n4832), .B(n4828), .Z(n4901) );
  XNOR U7953 ( .A(n4827), .B(n4823), .Z(n4902) );
  XNOR U7954 ( .A(n4822), .B(n4818), .Z(n4903) );
  XNOR U7955 ( .A(n4817), .B(n4813), .Z(n4904) );
  XNOR U7956 ( .A(n4812), .B(n4808), .Z(n4905) );
  XNOR U7957 ( .A(n4807), .B(n4803), .Z(n4906) );
  XNOR U7958 ( .A(n4802), .B(n4798), .Z(n4907) );
  XNOR U7959 ( .A(n4797), .B(n4793), .Z(n4908) );
  XNOR U7960 ( .A(n4792), .B(n4788), .Z(n4909) );
  XNOR U7961 ( .A(n4787), .B(n4783), .Z(n4910) );
  XNOR U7962 ( .A(n4782), .B(n4778), .Z(n4911) );
  XNOR U7963 ( .A(n4777), .B(n4773), .Z(n4912) );
  XNOR U7964 ( .A(n4772), .B(n4768), .Z(n4913) );
  XNOR U7965 ( .A(n4767), .B(n4763), .Z(n4914) );
  XNOR U7966 ( .A(n4762), .B(n4758), .Z(n4915) );
  XNOR U7967 ( .A(n4757), .B(n4753), .Z(n4916) );
  XOR U7968 ( .A(n4752), .B(n4749), .Z(n4917) );
  XOR U7969 ( .A(n4918), .B(n4919), .Z(n4749) );
  XOR U7970 ( .A(n4747), .B(n4920), .Z(n4919) );
  XNOR U7971 ( .A(n4921), .B(n4922), .Z(n4920) );
  XOR U7972 ( .A(n4923), .B(n4924), .Z(n4922) );
  NAND U7973 ( .A(a[70]), .B(b[30]), .Z(n4924) );
  AND U7974 ( .A(a[69]), .B(b[31]), .Z(n4923) );
  XNOR U7975 ( .A(n4925), .B(n4921), .Z(n4918) );
  XNOR U7976 ( .A(n4926), .B(n4927), .Z(n4921) );
  ANDN U7977 ( .B(n4928), .A(n4929), .Z(n4926) );
  AND U7978 ( .A(a[71]), .B(b[29]), .Z(n4925) );
  XOR U7979 ( .A(n4930), .B(n4747), .Z(n4748) );
  XOR U7980 ( .A(n4931), .B(n4932), .Z(n4747) );
  AND U7981 ( .A(n4933), .B(n4934), .Z(n4931) );
  AND U7982 ( .A(a[72]), .B(b[28]), .Z(n4930) );
  XOR U7983 ( .A(n4935), .B(n4752), .Z(n4754) );
  XOR U7984 ( .A(n4936), .B(n4937), .Z(n4752) );
  AND U7985 ( .A(n4938), .B(n4939), .Z(n4936) );
  AND U7986 ( .A(a[73]), .B(b[27]), .Z(n4935) );
  XOR U7987 ( .A(n4940), .B(n4757), .Z(n4759) );
  XOR U7988 ( .A(n4941), .B(n4942), .Z(n4757) );
  AND U7989 ( .A(n4943), .B(n4944), .Z(n4941) );
  AND U7990 ( .A(a[74]), .B(b[26]), .Z(n4940) );
  XOR U7991 ( .A(n4945), .B(n4762), .Z(n4764) );
  XOR U7992 ( .A(n4946), .B(n4947), .Z(n4762) );
  AND U7993 ( .A(n4948), .B(n4949), .Z(n4946) );
  AND U7994 ( .A(a[75]), .B(b[25]), .Z(n4945) );
  XOR U7995 ( .A(n4950), .B(n4767), .Z(n4769) );
  XOR U7996 ( .A(n4951), .B(n4952), .Z(n4767) );
  AND U7997 ( .A(n4953), .B(n4954), .Z(n4951) );
  AND U7998 ( .A(a[76]), .B(b[24]), .Z(n4950) );
  XOR U7999 ( .A(n4955), .B(n4772), .Z(n4774) );
  XOR U8000 ( .A(n4956), .B(n4957), .Z(n4772) );
  AND U8001 ( .A(n4958), .B(n4959), .Z(n4956) );
  AND U8002 ( .A(a[77]), .B(b[23]), .Z(n4955) );
  XOR U8003 ( .A(n4960), .B(n4777), .Z(n4779) );
  XOR U8004 ( .A(n4961), .B(n4962), .Z(n4777) );
  AND U8005 ( .A(n4963), .B(n4964), .Z(n4961) );
  AND U8006 ( .A(a[78]), .B(b[22]), .Z(n4960) );
  XOR U8007 ( .A(n4965), .B(n4782), .Z(n4784) );
  XOR U8008 ( .A(n4966), .B(n4967), .Z(n4782) );
  AND U8009 ( .A(n4968), .B(n4969), .Z(n4966) );
  AND U8010 ( .A(a[79]), .B(b[21]), .Z(n4965) );
  XOR U8011 ( .A(n4970), .B(n4787), .Z(n4789) );
  XOR U8012 ( .A(n4971), .B(n4972), .Z(n4787) );
  AND U8013 ( .A(n4973), .B(n4974), .Z(n4971) );
  AND U8014 ( .A(a[80]), .B(b[20]), .Z(n4970) );
  XOR U8015 ( .A(n4975), .B(n4792), .Z(n4794) );
  XOR U8016 ( .A(n4976), .B(n4977), .Z(n4792) );
  AND U8017 ( .A(n4978), .B(n4979), .Z(n4976) );
  AND U8018 ( .A(a[81]), .B(b[19]), .Z(n4975) );
  XOR U8019 ( .A(n4980), .B(n4797), .Z(n4799) );
  XOR U8020 ( .A(n4981), .B(n4982), .Z(n4797) );
  AND U8021 ( .A(n4983), .B(n4984), .Z(n4981) );
  AND U8022 ( .A(a[82]), .B(b[18]), .Z(n4980) );
  XOR U8023 ( .A(n4985), .B(n4802), .Z(n4804) );
  XOR U8024 ( .A(n4986), .B(n4987), .Z(n4802) );
  AND U8025 ( .A(n4988), .B(n4989), .Z(n4986) );
  AND U8026 ( .A(a[83]), .B(b[17]), .Z(n4985) );
  XOR U8027 ( .A(n4990), .B(n4807), .Z(n4809) );
  XOR U8028 ( .A(n4991), .B(n4992), .Z(n4807) );
  AND U8029 ( .A(n4993), .B(n4994), .Z(n4991) );
  AND U8030 ( .A(a[84]), .B(b[16]), .Z(n4990) );
  XOR U8031 ( .A(n4995), .B(n4812), .Z(n4814) );
  XOR U8032 ( .A(n4996), .B(n4997), .Z(n4812) );
  AND U8033 ( .A(n4998), .B(n4999), .Z(n4996) );
  AND U8034 ( .A(a[85]), .B(b[15]), .Z(n4995) );
  XOR U8035 ( .A(n5000), .B(n4817), .Z(n4819) );
  XOR U8036 ( .A(n5001), .B(n5002), .Z(n4817) );
  AND U8037 ( .A(n5003), .B(n5004), .Z(n5001) );
  AND U8038 ( .A(a[86]), .B(b[14]), .Z(n5000) );
  XOR U8039 ( .A(n5005), .B(n4822), .Z(n4824) );
  XOR U8040 ( .A(n5006), .B(n5007), .Z(n4822) );
  AND U8041 ( .A(n5008), .B(n5009), .Z(n5006) );
  AND U8042 ( .A(a[87]), .B(b[13]), .Z(n5005) );
  XOR U8043 ( .A(n5010), .B(n4827), .Z(n4829) );
  XOR U8044 ( .A(n5011), .B(n5012), .Z(n4827) );
  AND U8045 ( .A(n5013), .B(n5014), .Z(n5011) );
  AND U8046 ( .A(a[88]), .B(b[12]), .Z(n5010) );
  XOR U8047 ( .A(n5015), .B(n4832), .Z(n4834) );
  XOR U8048 ( .A(n5016), .B(n5017), .Z(n4832) );
  AND U8049 ( .A(n5018), .B(n5019), .Z(n5016) );
  AND U8050 ( .A(a[89]), .B(b[11]), .Z(n5015) );
  XOR U8051 ( .A(n5020), .B(n4837), .Z(n4839) );
  XOR U8052 ( .A(n5021), .B(n5022), .Z(n4837) );
  AND U8053 ( .A(n5023), .B(n5024), .Z(n5021) );
  AND U8054 ( .A(a[90]), .B(b[10]), .Z(n5020) );
  XOR U8055 ( .A(n5025), .B(n4842), .Z(n4844) );
  XOR U8056 ( .A(n5026), .B(n5027), .Z(n4842) );
  AND U8057 ( .A(n5028), .B(n5029), .Z(n5026) );
  AND U8058 ( .A(a[91]), .B(b[9]), .Z(n5025) );
  XOR U8059 ( .A(n5030), .B(n4847), .Z(n4849) );
  XOR U8060 ( .A(n5031), .B(n5032), .Z(n4847) );
  AND U8061 ( .A(n5033), .B(n5034), .Z(n5031) );
  AND U8062 ( .A(a[92]), .B(b[8]), .Z(n5030) );
  XOR U8063 ( .A(n5035), .B(n4852), .Z(n4854) );
  XOR U8064 ( .A(n5036), .B(n5037), .Z(n4852) );
  AND U8065 ( .A(n5038), .B(n5039), .Z(n5036) );
  AND U8066 ( .A(a[93]), .B(b[7]), .Z(n5035) );
  XOR U8067 ( .A(n5040), .B(n4857), .Z(n4859) );
  XOR U8068 ( .A(n5041), .B(n5042), .Z(n4857) );
  AND U8069 ( .A(n5043), .B(n5044), .Z(n5041) );
  AND U8070 ( .A(a[94]), .B(b[6]), .Z(n5040) );
  XOR U8071 ( .A(n5045), .B(n4862), .Z(n4864) );
  XOR U8072 ( .A(n5046), .B(n5047), .Z(n4862) );
  AND U8073 ( .A(n5048), .B(n5049), .Z(n5046) );
  AND U8074 ( .A(b[5]), .B(a[95]), .Z(n5045) );
  XOR U8075 ( .A(n5050), .B(n4867), .Z(n4869) );
  XOR U8076 ( .A(n5051), .B(n5052), .Z(n4867) );
  AND U8077 ( .A(n5053), .B(n5054), .Z(n5051) );
  AND U8078 ( .A(b[4]), .B(a[96]), .Z(n5050) );
  XNOR U8079 ( .A(n5055), .B(n5056), .Z(n4881) );
  NANDN U8080 ( .A(n5057), .B(n5058), .Z(n5056) );
  XOR U8081 ( .A(n5059), .B(n4872), .Z(n4874) );
  XOR U8082 ( .A(n5060), .B(n5061), .Z(n4872) );
  AND U8083 ( .A(n5062), .B(n5063), .Z(n5060) );
  AND U8084 ( .A(b[3]), .B(a[97]), .Z(n5059) );
  NAND U8085 ( .A(a[100]), .B(b[0]), .Z(n4710) );
  XOR U8086 ( .A(n4891), .B(n5064), .Z(n2) );
  XNOR U8087 ( .A(n4890), .B(n1), .Z(n5064) );
  XOR U8088 ( .A(n5066), .B(n5067), .Z(n4) );
  XNOR U8089 ( .A(n5068), .B(n5065), .Z(n5067) );
  IV U8090 ( .A(n3), .Z(n5065) );
  XNOR U8091 ( .A(n5069), .B(n5070), .Z(n6) );
  XOR U8092 ( .A(n5072), .B(n5073), .Z(n8) );
  XOR U8093 ( .A(n5074), .B(n7), .Z(n5073) );
  XNOR U8094 ( .A(n5075), .B(n5076), .Z(n7) );
  NOR U8095 ( .A(n10), .B(n9), .Z(n5075) );
  XOR U8096 ( .A(n5077), .B(n5078), .Z(n9) );
  XNOR U8097 ( .A(n5079), .B(n5076), .Z(n5078) );
  XOR U8098 ( .A(sreg[223]), .B(n5076), .Z(n10) );
  XOR U8099 ( .A(n5080), .B(n5081), .Z(n5076) );
  NOR U8100 ( .A(n12), .B(n11), .Z(n5080) );
  XOR U8101 ( .A(n5082), .B(n5083), .Z(n11) );
  XNOR U8102 ( .A(n5084), .B(n5081), .Z(n5083) );
  XOR U8103 ( .A(sreg[222]), .B(n5081), .Z(n12) );
  XOR U8104 ( .A(n5085), .B(n5086), .Z(n5081) );
  NOR U8105 ( .A(n14), .B(n13), .Z(n5085) );
  XOR U8106 ( .A(n5087), .B(n5088), .Z(n13) );
  XNOR U8107 ( .A(n5089), .B(n5086), .Z(n5088) );
  XOR U8108 ( .A(sreg[221]), .B(n5086), .Z(n14) );
  XOR U8109 ( .A(n5090), .B(n5091), .Z(n5086) );
  NOR U8110 ( .A(n16), .B(n15), .Z(n5090) );
  XOR U8111 ( .A(n5092), .B(n5093), .Z(n15) );
  XNOR U8112 ( .A(n5094), .B(n5091), .Z(n5093) );
  XOR U8113 ( .A(sreg[220]), .B(n5091), .Z(n16) );
  XOR U8114 ( .A(n5095), .B(n5096), .Z(n5091) );
  NOR U8115 ( .A(n18), .B(n17), .Z(n5095) );
  XOR U8116 ( .A(n5097), .B(n5098), .Z(n17) );
  XNOR U8117 ( .A(n5099), .B(n5096), .Z(n5098) );
  XOR U8118 ( .A(sreg[219]), .B(n5096), .Z(n18) );
  XOR U8119 ( .A(n5100), .B(n5101), .Z(n5096) );
  NOR U8120 ( .A(n20), .B(n19), .Z(n5100) );
  XOR U8121 ( .A(n5102), .B(n5103), .Z(n19) );
  XNOR U8122 ( .A(n5104), .B(n5101), .Z(n5103) );
  XOR U8123 ( .A(sreg[218]), .B(n5101), .Z(n20) );
  XOR U8124 ( .A(n5105), .B(n5106), .Z(n5101) );
  NOR U8125 ( .A(n22), .B(n21), .Z(n5105) );
  XOR U8126 ( .A(n5107), .B(n5108), .Z(n21) );
  XNOR U8127 ( .A(n5109), .B(n5106), .Z(n5108) );
  XOR U8128 ( .A(sreg[217]), .B(n5106), .Z(n22) );
  XOR U8129 ( .A(n5110), .B(n5111), .Z(n5106) );
  NOR U8130 ( .A(n24), .B(n23), .Z(n5110) );
  XOR U8131 ( .A(n5112), .B(n5113), .Z(n23) );
  XNOR U8132 ( .A(n5114), .B(n5111), .Z(n5113) );
  XOR U8133 ( .A(sreg[216]), .B(n5111), .Z(n24) );
  XOR U8134 ( .A(n5115), .B(n5116), .Z(n5111) );
  NOR U8135 ( .A(n26), .B(n25), .Z(n5115) );
  XOR U8136 ( .A(n5117), .B(n5118), .Z(n25) );
  XNOR U8137 ( .A(n5119), .B(n5116), .Z(n5118) );
  XOR U8138 ( .A(sreg[215]), .B(n5116), .Z(n26) );
  XOR U8139 ( .A(n5120), .B(n5121), .Z(n5116) );
  NOR U8140 ( .A(n28), .B(n27), .Z(n5120) );
  XOR U8141 ( .A(n5122), .B(n5123), .Z(n27) );
  XNOR U8142 ( .A(n5124), .B(n5121), .Z(n5123) );
  XOR U8143 ( .A(sreg[214]), .B(n5121), .Z(n28) );
  XOR U8144 ( .A(n5125), .B(n5126), .Z(n5121) );
  NOR U8145 ( .A(n30), .B(n29), .Z(n5125) );
  XOR U8146 ( .A(n5127), .B(n5128), .Z(n29) );
  XNOR U8147 ( .A(n5129), .B(n5126), .Z(n5128) );
  XOR U8148 ( .A(sreg[213]), .B(n5126), .Z(n30) );
  XOR U8149 ( .A(n5130), .B(n5131), .Z(n5126) );
  NOR U8150 ( .A(n32), .B(n31), .Z(n5130) );
  XOR U8151 ( .A(n5132), .B(n5133), .Z(n31) );
  XNOR U8152 ( .A(n5134), .B(n5131), .Z(n5133) );
  XOR U8153 ( .A(sreg[212]), .B(n5131), .Z(n32) );
  XOR U8154 ( .A(n5135), .B(n5136), .Z(n5131) );
  NOR U8155 ( .A(n34), .B(n33), .Z(n5135) );
  XOR U8156 ( .A(n5137), .B(n5138), .Z(n33) );
  XNOR U8157 ( .A(n5139), .B(n5136), .Z(n5138) );
  XOR U8158 ( .A(sreg[211]), .B(n5136), .Z(n34) );
  XOR U8159 ( .A(n5140), .B(n5141), .Z(n5136) );
  NOR U8160 ( .A(n36), .B(n35), .Z(n5140) );
  XOR U8161 ( .A(n5142), .B(n5143), .Z(n35) );
  XNOR U8162 ( .A(n5144), .B(n5141), .Z(n5143) );
  XOR U8163 ( .A(sreg[210]), .B(n5141), .Z(n36) );
  XOR U8164 ( .A(n5145), .B(n5146), .Z(n5141) );
  NOR U8165 ( .A(n38), .B(n37), .Z(n5145) );
  XOR U8166 ( .A(n5147), .B(n5148), .Z(n37) );
  XNOR U8167 ( .A(n5149), .B(n5146), .Z(n5148) );
  XOR U8168 ( .A(sreg[209]), .B(n5146), .Z(n38) );
  XOR U8169 ( .A(n5150), .B(n5151), .Z(n5146) );
  NOR U8170 ( .A(n40), .B(n39), .Z(n5150) );
  XOR U8171 ( .A(n5152), .B(n5153), .Z(n39) );
  XNOR U8172 ( .A(n5154), .B(n5151), .Z(n5153) );
  XOR U8173 ( .A(sreg[208]), .B(n5151), .Z(n40) );
  XOR U8174 ( .A(n5155), .B(n5156), .Z(n5151) );
  NOR U8175 ( .A(n42), .B(n41), .Z(n5155) );
  XOR U8176 ( .A(n5157), .B(n5158), .Z(n41) );
  XNOR U8177 ( .A(n5159), .B(n5156), .Z(n5158) );
  XOR U8178 ( .A(sreg[207]), .B(n5156), .Z(n42) );
  XOR U8179 ( .A(n5160), .B(n5161), .Z(n5156) );
  NOR U8180 ( .A(n44), .B(n43), .Z(n5160) );
  XOR U8181 ( .A(n5162), .B(n5163), .Z(n43) );
  XNOR U8182 ( .A(n5164), .B(n5161), .Z(n5163) );
  XOR U8183 ( .A(sreg[206]), .B(n5161), .Z(n44) );
  XOR U8184 ( .A(n5165), .B(n5166), .Z(n5161) );
  NOR U8185 ( .A(n46), .B(n45), .Z(n5165) );
  XOR U8186 ( .A(n5167), .B(n5168), .Z(n45) );
  XNOR U8187 ( .A(n5169), .B(n5166), .Z(n5168) );
  XOR U8188 ( .A(sreg[205]), .B(n5166), .Z(n46) );
  XOR U8189 ( .A(n5170), .B(n5171), .Z(n5166) );
  NOR U8190 ( .A(n48), .B(n47), .Z(n5170) );
  XOR U8191 ( .A(n5172), .B(n5173), .Z(n47) );
  XNOR U8192 ( .A(n5174), .B(n5171), .Z(n5173) );
  XOR U8193 ( .A(sreg[204]), .B(n5171), .Z(n48) );
  XOR U8194 ( .A(n5175), .B(n5176), .Z(n5171) );
  NOR U8195 ( .A(n50), .B(n49), .Z(n5175) );
  XOR U8196 ( .A(n5177), .B(n5178), .Z(n49) );
  XNOR U8197 ( .A(n5179), .B(n5176), .Z(n5178) );
  XOR U8198 ( .A(sreg[203]), .B(n5176), .Z(n50) );
  XOR U8199 ( .A(n5180), .B(n5181), .Z(n5176) );
  NOR U8200 ( .A(n52), .B(n51), .Z(n5180) );
  XOR U8201 ( .A(n5182), .B(n5183), .Z(n51) );
  XNOR U8202 ( .A(n5184), .B(n5181), .Z(n5183) );
  XOR U8203 ( .A(sreg[202]), .B(n5181), .Z(n52) );
  XOR U8204 ( .A(n5185), .B(n5186), .Z(n5181) );
  NOR U8205 ( .A(n54), .B(n53), .Z(n5185) );
  XOR U8206 ( .A(n5187), .B(n5188), .Z(n53) );
  XNOR U8207 ( .A(n5189), .B(n5186), .Z(n5188) );
  XOR U8208 ( .A(sreg[201]), .B(n5186), .Z(n54) );
  XOR U8209 ( .A(n5190), .B(n5191), .Z(n5186) );
  NOR U8210 ( .A(n56), .B(n55), .Z(n5190) );
  XOR U8211 ( .A(n5192), .B(n5193), .Z(n55) );
  XNOR U8212 ( .A(n5194), .B(n5191), .Z(n5193) );
  XOR U8213 ( .A(sreg[200]), .B(n5191), .Z(n56) );
  XOR U8214 ( .A(n5195), .B(n5196), .Z(n5191) );
  NOR U8215 ( .A(n58), .B(n57), .Z(n5195) );
  XOR U8216 ( .A(n5197), .B(n5198), .Z(n57) );
  XNOR U8217 ( .A(n5199), .B(n5196), .Z(n5198) );
  XOR U8218 ( .A(sreg[199]), .B(n5196), .Z(n58) );
  XOR U8219 ( .A(n5200), .B(n5201), .Z(n5196) );
  NOR U8220 ( .A(n60), .B(n59), .Z(n5200) );
  XOR U8221 ( .A(n5202), .B(n5203), .Z(n59) );
  XNOR U8222 ( .A(n5204), .B(n5201), .Z(n5203) );
  XOR U8223 ( .A(sreg[198]), .B(n5201), .Z(n60) );
  XOR U8224 ( .A(n5205), .B(n5206), .Z(n5201) );
  NOR U8225 ( .A(n62), .B(n61), .Z(n5205) );
  XOR U8226 ( .A(n5207), .B(n5208), .Z(n61) );
  XNOR U8227 ( .A(n5209), .B(n5206), .Z(n5208) );
  XOR U8228 ( .A(sreg[197]), .B(n5206), .Z(n62) );
  XOR U8229 ( .A(n5210), .B(n5211), .Z(n5206) );
  NOR U8230 ( .A(n64), .B(n63), .Z(n5210) );
  XOR U8231 ( .A(n5212), .B(n5213), .Z(n63) );
  XNOR U8232 ( .A(n5214), .B(n5211), .Z(n5213) );
  XOR U8233 ( .A(sreg[196]), .B(n5211), .Z(n64) );
  XOR U8234 ( .A(n5215), .B(n5216), .Z(n5211) );
  NOR U8235 ( .A(n66), .B(n65), .Z(n5215) );
  XOR U8236 ( .A(n5217), .B(n5218), .Z(n65) );
  XNOR U8237 ( .A(n5219), .B(n5216), .Z(n5218) );
  XOR U8238 ( .A(sreg[195]), .B(n5216), .Z(n66) );
  XOR U8239 ( .A(n5220), .B(n5221), .Z(n5216) );
  NOR U8240 ( .A(n68), .B(n67), .Z(n5220) );
  XOR U8241 ( .A(n5222), .B(n5223), .Z(n67) );
  XNOR U8242 ( .A(n5224), .B(n5221), .Z(n5223) );
  XOR U8243 ( .A(sreg[194]), .B(n5221), .Z(n68) );
  XOR U8244 ( .A(n5225), .B(n5226), .Z(n5221) );
  NOR U8245 ( .A(n70), .B(n69), .Z(n5225) );
  XOR U8246 ( .A(n5227), .B(n5228), .Z(n69) );
  XNOR U8247 ( .A(n5229), .B(n5226), .Z(n5228) );
  XOR U8248 ( .A(sreg[193]), .B(n5226), .Z(n70) );
  XOR U8249 ( .A(n5230), .B(n5231), .Z(n5226) );
  NOR U8250 ( .A(n72), .B(n71), .Z(n5230) );
  XOR U8251 ( .A(n5232), .B(n5233), .Z(n71) );
  XNOR U8252 ( .A(n5234), .B(n5231), .Z(n5233) );
  XOR U8253 ( .A(sreg[192]), .B(n5231), .Z(n72) );
  XOR U8254 ( .A(n5235), .B(n5236), .Z(n5231) );
  NOR U8255 ( .A(n74), .B(n73), .Z(n5235) );
  XOR U8256 ( .A(n5237), .B(n5238), .Z(n73) );
  XNOR U8257 ( .A(n5239), .B(n5236), .Z(n5238) );
  XOR U8258 ( .A(sreg[191]), .B(n5236), .Z(n74) );
  XOR U8259 ( .A(n5240), .B(n5241), .Z(n5236) );
  NOR U8260 ( .A(n76), .B(n75), .Z(n5240) );
  XOR U8261 ( .A(n5242), .B(n5243), .Z(n75) );
  XNOR U8262 ( .A(n5244), .B(n5241), .Z(n5243) );
  XOR U8263 ( .A(sreg[190]), .B(n5241), .Z(n76) );
  XOR U8264 ( .A(n5245), .B(n5246), .Z(n5241) );
  NOR U8265 ( .A(n78), .B(n77), .Z(n5245) );
  XOR U8266 ( .A(n5247), .B(n5248), .Z(n77) );
  XNOR U8267 ( .A(n5249), .B(n5246), .Z(n5248) );
  XOR U8268 ( .A(sreg[189]), .B(n5246), .Z(n78) );
  XOR U8269 ( .A(n5250), .B(n5251), .Z(n5246) );
  NOR U8270 ( .A(n80), .B(n79), .Z(n5250) );
  XOR U8271 ( .A(n5252), .B(n5253), .Z(n79) );
  XNOR U8272 ( .A(n5254), .B(n5251), .Z(n5253) );
  XOR U8273 ( .A(sreg[188]), .B(n5251), .Z(n80) );
  XOR U8274 ( .A(n5255), .B(n5256), .Z(n5251) );
  NOR U8275 ( .A(n82), .B(n81), .Z(n5255) );
  XOR U8276 ( .A(n5257), .B(n5258), .Z(n81) );
  XNOR U8277 ( .A(n5259), .B(n5256), .Z(n5258) );
  XOR U8278 ( .A(sreg[187]), .B(n5256), .Z(n82) );
  XOR U8279 ( .A(n5260), .B(n5261), .Z(n5256) );
  NOR U8280 ( .A(n84), .B(n83), .Z(n5260) );
  XOR U8281 ( .A(n5262), .B(n5263), .Z(n83) );
  XNOR U8282 ( .A(n5264), .B(n5261), .Z(n5263) );
  XOR U8283 ( .A(sreg[186]), .B(n5261), .Z(n84) );
  XOR U8284 ( .A(n5265), .B(n5266), .Z(n5261) );
  NOR U8285 ( .A(n86), .B(n85), .Z(n5265) );
  XOR U8286 ( .A(n5267), .B(n5268), .Z(n85) );
  XNOR U8287 ( .A(n5269), .B(n5266), .Z(n5268) );
  XOR U8288 ( .A(sreg[185]), .B(n5266), .Z(n86) );
  XOR U8289 ( .A(n5270), .B(n5271), .Z(n5266) );
  NOR U8290 ( .A(n88), .B(n87), .Z(n5270) );
  XOR U8291 ( .A(n5272), .B(n5273), .Z(n87) );
  XNOR U8292 ( .A(n5274), .B(n5271), .Z(n5273) );
  XOR U8293 ( .A(sreg[184]), .B(n5271), .Z(n88) );
  XOR U8294 ( .A(n5275), .B(n5276), .Z(n5271) );
  NOR U8295 ( .A(n90), .B(n89), .Z(n5275) );
  XOR U8296 ( .A(n5277), .B(n5278), .Z(n89) );
  XNOR U8297 ( .A(n5279), .B(n5276), .Z(n5278) );
  XOR U8298 ( .A(sreg[183]), .B(n5276), .Z(n90) );
  XOR U8299 ( .A(n5280), .B(n5281), .Z(n5276) );
  NOR U8300 ( .A(n92), .B(n91), .Z(n5280) );
  XOR U8301 ( .A(n5282), .B(n5283), .Z(n91) );
  XNOR U8302 ( .A(n5284), .B(n5281), .Z(n5283) );
  XOR U8303 ( .A(sreg[182]), .B(n5281), .Z(n92) );
  XOR U8304 ( .A(n5285), .B(n5286), .Z(n5281) );
  NOR U8305 ( .A(n94), .B(n93), .Z(n5285) );
  XOR U8306 ( .A(n5287), .B(n5288), .Z(n93) );
  XNOR U8307 ( .A(n5289), .B(n5286), .Z(n5288) );
  XOR U8308 ( .A(sreg[181]), .B(n5286), .Z(n94) );
  XOR U8309 ( .A(n5290), .B(n5291), .Z(n5286) );
  NOR U8310 ( .A(n96), .B(n95), .Z(n5290) );
  XOR U8311 ( .A(n5292), .B(n5293), .Z(n95) );
  XNOR U8312 ( .A(n5294), .B(n5291), .Z(n5293) );
  XOR U8313 ( .A(sreg[180]), .B(n5291), .Z(n96) );
  XOR U8314 ( .A(n5295), .B(n5296), .Z(n5291) );
  NOR U8315 ( .A(n98), .B(n97), .Z(n5295) );
  XOR U8316 ( .A(n5297), .B(n5298), .Z(n97) );
  XNOR U8317 ( .A(n5299), .B(n5296), .Z(n5298) );
  XOR U8318 ( .A(sreg[179]), .B(n5296), .Z(n98) );
  XOR U8319 ( .A(n5300), .B(n5301), .Z(n5296) );
  NOR U8320 ( .A(n100), .B(n99), .Z(n5300) );
  XOR U8321 ( .A(n5302), .B(n5303), .Z(n99) );
  XNOR U8322 ( .A(n5304), .B(n5301), .Z(n5303) );
  XOR U8323 ( .A(sreg[178]), .B(n5301), .Z(n100) );
  XOR U8324 ( .A(n5305), .B(n5306), .Z(n5301) );
  NOR U8325 ( .A(n102), .B(n101), .Z(n5305) );
  XOR U8326 ( .A(n5307), .B(n5308), .Z(n101) );
  XNOR U8327 ( .A(n5309), .B(n5306), .Z(n5308) );
  XOR U8328 ( .A(sreg[177]), .B(n5306), .Z(n102) );
  XOR U8329 ( .A(n5310), .B(n5311), .Z(n5306) );
  NOR U8330 ( .A(n104), .B(n103), .Z(n5310) );
  XOR U8331 ( .A(n5312), .B(n5313), .Z(n103) );
  XNOR U8332 ( .A(n5314), .B(n5311), .Z(n5313) );
  XOR U8333 ( .A(sreg[176]), .B(n5311), .Z(n104) );
  XOR U8334 ( .A(n5315), .B(n5316), .Z(n5311) );
  NOR U8335 ( .A(n106), .B(n105), .Z(n5315) );
  XOR U8336 ( .A(n5317), .B(n5318), .Z(n105) );
  XNOR U8337 ( .A(n5319), .B(n5316), .Z(n5318) );
  XOR U8338 ( .A(sreg[175]), .B(n5316), .Z(n106) );
  XOR U8339 ( .A(n5320), .B(n5321), .Z(n5316) );
  NOR U8340 ( .A(n108), .B(n107), .Z(n5320) );
  XOR U8341 ( .A(n5322), .B(n5323), .Z(n107) );
  XNOR U8342 ( .A(n5324), .B(n5321), .Z(n5323) );
  XOR U8343 ( .A(sreg[174]), .B(n5321), .Z(n108) );
  XOR U8344 ( .A(n5325), .B(n5326), .Z(n5321) );
  NOR U8345 ( .A(n110), .B(n109), .Z(n5325) );
  XOR U8346 ( .A(n5327), .B(n5328), .Z(n109) );
  XNOR U8347 ( .A(n5329), .B(n5326), .Z(n5328) );
  XOR U8348 ( .A(sreg[173]), .B(n5326), .Z(n110) );
  XOR U8349 ( .A(n5330), .B(n5331), .Z(n5326) );
  NOR U8350 ( .A(n112), .B(n111), .Z(n5330) );
  XOR U8351 ( .A(n5332), .B(n5333), .Z(n111) );
  XNOR U8352 ( .A(n5334), .B(n5331), .Z(n5333) );
  XOR U8353 ( .A(sreg[172]), .B(n5331), .Z(n112) );
  XOR U8354 ( .A(n5335), .B(n5336), .Z(n5331) );
  NOR U8355 ( .A(n114), .B(n113), .Z(n5335) );
  XOR U8356 ( .A(n5337), .B(n5338), .Z(n113) );
  XNOR U8357 ( .A(n5339), .B(n5336), .Z(n5338) );
  XOR U8358 ( .A(sreg[171]), .B(n5336), .Z(n114) );
  XOR U8359 ( .A(n5340), .B(n5341), .Z(n5336) );
  NOR U8360 ( .A(n116), .B(n115), .Z(n5340) );
  XOR U8361 ( .A(n5342), .B(n5343), .Z(n115) );
  XNOR U8362 ( .A(n5344), .B(n5341), .Z(n5343) );
  XOR U8363 ( .A(sreg[170]), .B(n5341), .Z(n116) );
  XOR U8364 ( .A(n5345), .B(n5346), .Z(n5341) );
  NOR U8365 ( .A(n118), .B(n117), .Z(n5345) );
  XOR U8366 ( .A(n5347), .B(n5348), .Z(n117) );
  XNOR U8367 ( .A(n5349), .B(n5346), .Z(n5348) );
  XOR U8368 ( .A(sreg[169]), .B(n5346), .Z(n118) );
  XOR U8369 ( .A(n5350), .B(n5351), .Z(n5346) );
  NOR U8370 ( .A(n120), .B(n119), .Z(n5350) );
  XOR U8371 ( .A(n5352), .B(n5353), .Z(n119) );
  XNOR U8372 ( .A(n5354), .B(n5351), .Z(n5353) );
  XOR U8373 ( .A(sreg[168]), .B(n5351), .Z(n120) );
  XOR U8374 ( .A(n5355), .B(n5356), .Z(n5351) );
  NOR U8375 ( .A(n122), .B(n121), .Z(n5355) );
  XOR U8376 ( .A(n5357), .B(n5358), .Z(n121) );
  XNOR U8377 ( .A(n5359), .B(n5356), .Z(n5358) );
  XOR U8378 ( .A(sreg[167]), .B(n5356), .Z(n122) );
  XOR U8379 ( .A(n5360), .B(n5361), .Z(n5356) );
  NOR U8380 ( .A(n124), .B(n123), .Z(n5360) );
  XOR U8381 ( .A(n5362), .B(n5363), .Z(n123) );
  XNOR U8382 ( .A(n5364), .B(n5361), .Z(n5363) );
  XOR U8383 ( .A(sreg[166]), .B(n5361), .Z(n124) );
  XOR U8384 ( .A(n5365), .B(n5366), .Z(n5361) );
  NOR U8385 ( .A(n126), .B(n125), .Z(n5365) );
  XOR U8386 ( .A(n5367), .B(n5368), .Z(n125) );
  XNOR U8387 ( .A(n5369), .B(n5366), .Z(n5368) );
  XOR U8388 ( .A(sreg[165]), .B(n5366), .Z(n126) );
  XOR U8389 ( .A(n5370), .B(n5371), .Z(n5366) );
  NOR U8390 ( .A(n128), .B(n127), .Z(n5370) );
  XOR U8391 ( .A(n5372), .B(n5373), .Z(n127) );
  XNOR U8392 ( .A(n5374), .B(n5371), .Z(n5373) );
  XOR U8393 ( .A(sreg[164]), .B(n5371), .Z(n128) );
  XOR U8394 ( .A(n5375), .B(n5376), .Z(n5371) );
  NOR U8395 ( .A(n130), .B(n129), .Z(n5375) );
  XOR U8396 ( .A(n5377), .B(n5378), .Z(n129) );
  XNOR U8397 ( .A(n5379), .B(n5376), .Z(n5378) );
  XOR U8398 ( .A(sreg[163]), .B(n5376), .Z(n130) );
  XOR U8399 ( .A(n5380), .B(n5381), .Z(n5376) );
  NOR U8400 ( .A(n132), .B(n131), .Z(n5380) );
  XOR U8401 ( .A(n5382), .B(n5383), .Z(n131) );
  XNOR U8402 ( .A(n5384), .B(n5381), .Z(n5383) );
  XOR U8403 ( .A(sreg[162]), .B(n5381), .Z(n132) );
  XOR U8404 ( .A(n5385), .B(n5386), .Z(n5381) );
  NOR U8405 ( .A(n134), .B(n133), .Z(n5385) );
  XOR U8406 ( .A(n5387), .B(n5388), .Z(n133) );
  XNOR U8407 ( .A(n5389), .B(n5386), .Z(n5388) );
  XOR U8408 ( .A(sreg[161]), .B(n5386), .Z(n134) );
  XOR U8409 ( .A(n5390), .B(n5391), .Z(n5386) );
  NOR U8410 ( .A(n136), .B(n135), .Z(n5390) );
  XOR U8411 ( .A(n5392), .B(n5393), .Z(n135) );
  XNOR U8412 ( .A(n5394), .B(n5391), .Z(n5393) );
  XOR U8413 ( .A(sreg[160]), .B(n5391), .Z(n136) );
  XOR U8414 ( .A(n5395), .B(n5396), .Z(n5391) );
  NOR U8415 ( .A(n5397), .B(n5398), .Z(n5395) );
  NAND U8416 ( .A(a[99]), .B(b[0]), .Z(n4890) );
  XOR U8417 ( .A(n5058), .B(n5057), .Z(n4891) );
  XOR U8418 ( .A(n5055), .B(n5062), .Z(n5399) );
  XOR U8419 ( .A(n5053), .B(n5401), .Z(n5400) );
  XOR U8420 ( .A(n5048), .B(n5403), .Z(n5402) );
  XOR U8421 ( .A(n5043), .B(n5405), .Z(n5404) );
  XOR U8422 ( .A(n5038), .B(n5407), .Z(n5406) );
  XOR U8423 ( .A(n5033), .B(n5409), .Z(n5408) );
  XOR U8424 ( .A(n5028), .B(n5411), .Z(n5410) );
  XOR U8425 ( .A(n5023), .B(n5413), .Z(n5412) );
  XOR U8426 ( .A(n5018), .B(n5415), .Z(n5414) );
  XOR U8427 ( .A(n5013), .B(n5417), .Z(n5416) );
  XOR U8428 ( .A(n5008), .B(n5419), .Z(n5418) );
  XOR U8429 ( .A(n5003), .B(n5421), .Z(n5420) );
  XOR U8430 ( .A(n4998), .B(n5423), .Z(n5422) );
  XOR U8431 ( .A(n4993), .B(n5425), .Z(n5424) );
  XOR U8432 ( .A(n4988), .B(n5427), .Z(n5426) );
  XOR U8433 ( .A(n4983), .B(n5429), .Z(n5428) );
  XOR U8434 ( .A(n4978), .B(n5431), .Z(n5430) );
  XOR U8435 ( .A(n4973), .B(n5433), .Z(n5432) );
  XOR U8436 ( .A(n4968), .B(n5435), .Z(n5434) );
  XOR U8437 ( .A(n4963), .B(n5437), .Z(n5436) );
  XOR U8438 ( .A(n4958), .B(n5439), .Z(n5438) );
  XOR U8439 ( .A(n4953), .B(n5441), .Z(n5440) );
  XOR U8440 ( .A(n4948), .B(n5443), .Z(n5442) );
  XOR U8441 ( .A(n4943), .B(n5445), .Z(n5444) );
  XOR U8442 ( .A(n4938), .B(n5447), .Z(n5446) );
  XOR U8443 ( .A(n4933), .B(n5449), .Z(n5448) );
  XNOR U8444 ( .A(n4929), .B(n5451), .Z(n5450) );
  XOR U8445 ( .A(n5452), .B(n5453), .Z(n4929) );
  XOR U8446 ( .A(n5454), .B(n5455), .Z(n5453) );
  XNOR U8447 ( .A(n5456), .B(n5457), .Z(n5454) );
  XOR U8448 ( .A(n5458), .B(n5459), .Z(n5457) );
  AND U8449 ( .A(b[31]), .B(a[68]), .Z(n5459) );
  AND U8450 ( .A(a[69]), .B(b[30]), .Z(n5458) );
  XNOR U8451 ( .A(n5460), .B(n5456), .Z(n5452) );
  XNOR U8452 ( .A(n5461), .B(n5462), .Z(n5456) );
  ANDN U8453 ( .B(n5463), .A(n5464), .Z(n5461) );
  AND U8454 ( .A(a[70]), .B(b[29]), .Z(n5460) );
  XOR U8455 ( .A(n5465), .B(n4927), .Z(n4928) );
  IV U8456 ( .A(n5455), .Z(n4927) );
  XOR U8457 ( .A(n5466), .B(n5467), .Z(n5455) );
  AND U8458 ( .A(n5468), .B(n5469), .Z(n5466) );
  AND U8459 ( .A(a[71]), .B(b[28]), .Z(n5465) );
  XOR U8460 ( .A(n5470), .B(n4932), .Z(n4934) );
  IV U8461 ( .A(n5451), .Z(n4932) );
  XOR U8462 ( .A(n5471), .B(n5472), .Z(n5451) );
  AND U8463 ( .A(n5473), .B(n5474), .Z(n5471) );
  AND U8464 ( .A(a[72]), .B(b[27]), .Z(n5470) );
  XOR U8465 ( .A(n5475), .B(n4937), .Z(n4939) );
  IV U8466 ( .A(n5449), .Z(n4937) );
  XOR U8467 ( .A(n5476), .B(n5477), .Z(n5449) );
  AND U8468 ( .A(n5478), .B(n5479), .Z(n5476) );
  AND U8469 ( .A(a[73]), .B(b[26]), .Z(n5475) );
  XOR U8470 ( .A(n5480), .B(n4942), .Z(n4944) );
  IV U8471 ( .A(n5447), .Z(n4942) );
  XOR U8472 ( .A(n5481), .B(n5482), .Z(n5447) );
  AND U8473 ( .A(n5483), .B(n5484), .Z(n5481) );
  AND U8474 ( .A(a[74]), .B(b[25]), .Z(n5480) );
  XOR U8475 ( .A(n5485), .B(n4947), .Z(n4949) );
  IV U8476 ( .A(n5445), .Z(n4947) );
  XOR U8477 ( .A(n5486), .B(n5487), .Z(n5445) );
  AND U8478 ( .A(n5488), .B(n5489), .Z(n5486) );
  AND U8479 ( .A(a[75]), .B(b[24]), .Z(n5485) );
  XOR U8480 ( .A(n5490), .B(n4952), .Z(n4954) );
  IV U8481 ( .A(n5443), .Z(n4952) );
  XOR U8482 ( .A(n5491), .B(n5492), .Z(n5443) );
  AND U8483 ( .A(n5493), .B(n5494), .Z(n5491) );
  AND U8484 ( .A(a[76]), .B(b[23]), .Z(n5490) );
  XOR U8485 ( .A(n5495), .B(n4957), .Z(n4959) );
  IV U8486 ( .A(n5441), .Z(n4957) );
  XOR U8487 ( .A(n5496), .B(n5497), .Z(n5441) );
  AND U8488 ( .A(n5498), .B(n5499), .Z(n5496) );
  AND U8489 ( .A(a[77]), .B(b[22]), .Z(n5495) );
  XOR U8490 ( .A(n5500), .B(n4962), .Z(n4964) );
  IV U8491 ( .A(n5439), .Z(n4962) );
  XOR U8492 ( .A(n5501), .B(n5502), .Z(n5439) );
  AND U8493 ( .A(n5503), .B(n5504), .Z(n5501) );
  AND U8494 ( .A(a[78]), .B(b[21]), .Z(n5500) );
  XOR U8495 ( .A(n5505), .B(n4967), .Z(n4969) );
  IV U8496 ( .A(n5437), .Z(n4967) );
  XOR U8497 ( .A(n5506), .B(n5507), .Z(n5437) );
  AND U8498 ( .A(n5508), .B(n5509), .Z(n5506) );
  AND U8499 ( .A(a[79]), .B(b[20]), .Z(n5505) );
  XOR U8500 ( .A(n5510), .B(n4972), .Z(n4974) );
  IV U8501 ( .A(n5435), .Z(n4972) );
  XOR U8502 ( .A(n5511), .B(n5512), .Z(n5435) );
  AND U8503 ( .A(n5513), .B(n5514), .Z(n5511) );
  AND U8504 ( .A(a[80]), .B(b[19]), .Z(n5510) );
  XOR U8505 ( .A(n5515), .B(n4977), .Z(n4979) );
  IV U8506 ( .A(n5433), .Z(n4977) );
  XOR U8507 ( .A(n5516), .B(n5517), .Z(n5433) );
  AND U8508 ( .A(n5518), .B(n5519), .Z(n5516) );
  AND U8509 ( .A(a[81]), .B(b[18]), .Z(n5515) );
  XOR U8510 ( .A(n5520), .B(n4982), .Z(n4984) );
  IV U8511 ( .A(n5431), .Z(n4982) );
  XOR U8512 ( .A(n5521), .B(n5522), .Z(n5431) );
  AND U8513 ( .A(n5523), .B(n5524), .Z(n5521) );
  AND U8514 ( .A(a[82]), .B(b[17]), .Z(n5520) );
  XOR U8515 ( .A(n5525), .B(n4987), .Z(n4989) );
  IV U8516 ( .A(n5429), .Z(n4987) );
  XOR U8517 ( .A(n5526), .B(n5527), .Z(n5429) );
  AND U8518 ( .A(n5528), .B(n5529), .Z(n5526) );
  AND U8519 ( .A(a[83]), .B(b[16]), .Z(n5525) );
  XOR U8520 ( .A(n5530), .B(n4992), .Z(n4994) );
  IV U8521 ( .A(n5427), .Z(n4992) );
  XOR U8522 ( .A(n5531), .B(n5532), .Z(n5427) );
  AND U8523 ( .A(n5533), .B(n5534), .Z(n5531) );
  AND U8524 ( .A(a[84]), .B(b[15]), .Z(n5530) );
  XOR U8525 ( .A(n5535), .B(n4997), .Z(n4999) );
  IV U8526 ( .A(n5425), .Z(n4997) );
  XOR U8527 ( .A(n5536), .B(n5537), .Z(n5425) );
  AND U8528 ( .A(n5538), .B(n5539), .Z(n5536) );
  AND U8529 ( .A(a[85]), .B(b[14]), .Z(n5535) );
  XOR U8530 ( .A(n5540), .B(n5002), .Z(n5004) );
  IV U8531 ( .A(n5423), .Z(n5002) );
  XOR U8532 ( .A(n5541), .B(n5542), .Z(n5423) );
  AND U8533 ( .A(n5543), .B(n5544), .Z(n5541) );
  AND U8534 ( .A(a[86]), .B(b[13]), .Z(n5540) );
  XOR U8535 ( .A(n5545), .B(n5007), .Z(n5009) );
  IV U8536 ( .A(n5421), .Z(n5007) );
  XOR U8537 ( .A(n5546), .B(n5547), .Z(n5421) );
  AND U8538 ( .A(n5548), .B(n5549), .Z(n5546) );
  AND U8539 ( .A(a[87]), .B(b[12]), .Z(n5545) );
  XOR U8540 ( .A(n5550), .B(n5012), .Z(n5014) );
  IV U8541 ( .A(n5419), .Z(n5012) );
  XOR U8542 ( .A(n5551), .B(n5552), .Z(n5419) );
  AND U8543 ( .A(n5553), .B(n5554), .Z(n5551) );
  AND U8544 ( .A(a[88]), .B(b[11]), .Z(n5550) );
  XOR U8545 ( .A(n5555), .B(n5017), .Z(n5019) );
  IV U8546 ( .A(n5417), .Z(n5017) );
  XOR U8547 ( .A(n5556), .B(n5557), .Z(n5417) );
  AND U8548 ( .A(n5558), .B(n5559), .Z(n5556) );
  AND U8549 ( .A(a[89]), .B(b[10]), .Z(n5555) );
  XOR U8550 ( .A(n5560), .B(n5022), .Z(n5024) );
  IV U8551 ( .A(n5415), .Z(n5022) );
  XOR U8552 ( .A(n5561), .B(n5562), .Z(n5415) );
  AND U8553 ( .A(n5563), .B(n5564), .Z(n5561) );
  AND U8554 ( .A(a[90]), .B(b[9]), .Z(n5560) );
  XOR U8555 ( .A(n5565), .B(n5027), .Z(n5029) );
  IV U8556 ( .A(n5413), .Z(n5027) );
  XOR U8557 ( .A(n5566), .B(n5567), .Z(n5413) );
  AND U8558 ( .A(n5568), .B(n5569), .Z(n5566) );
  AND U8559 ( .A(a[91]), .B(b[8]), .Z(n5565) );
  XOR U8560 ( .A(n5570), .B(n5032), .Z(n5034) );
  IV U8561 ( .A(n5411), .Z(n5032) );
  XOR U8562 ( .A(n5571), .B(n5572), .Z(n5411) );
  AND U8563 ( .A(n5573), .B(n5574), .Z(n5571) );
  AND U8564 ( .A(a[92]), .B(b[7]), .Z(n5570) );
  XOR U8565 ( .A(n5575), .B(n5037), .Z(n5039) );
  IV U8566 ( .A(n5409), .Z(n5037) );
  XOR U8567 ( .A(n5576), .B(n5577), .Z(n5409) );
  AND U8568 ( .A(n5578), .B(n5579), .Z(n5576) );
  AND U8569 ( .A(a[93]), .B(b[6]), .Z(n5575) );
  XOR U8570 ( .A(n5580), .B(n5042), .Z(n5044) );
  IV U8571 ( .A(n5407), .Z(n5042) );
  XOR U8572 ( .A(n5581), .B(n5582), .Z(n5407) );
  AND U8573 ( .A(n5583), .B(n5584), .Z(n5581) );
  AND U8574 ( .A(a[94]), .B(b[5]), .Z(n5580) );
  XOR U8575 ( .A(n5585), .B(n5047), .Z(n5049) );
  IV U8576 ( .A(n5405), .Z(n5047) );
  XOR U8577 ( .A(n5586), .B(n5587), .Z(n5405) );
  AND U8578 ( .A(n5588), .B(n5589), .Z(n5586) );
  AND U8579 ( .A(b[4]), .B(a[95]), .Z(n5585) );
  XOR U8580 ( .A(n5590), .B(n5052), .Z(n5054) );
  IV U8581 ( .A(n5403), .Z(n5052) );
  XOR U8582 ( .A(n5591), .B(n5592), .Z(n5403) );
  AND U8583 ( .A(n5593), .B(n5594), .Z(n5591) );
  AND U8584 ( .A(b[3]), .B(a[96]), .Z(n5590) );
  XOR U8585 ( .A(n5595), .B(n5061), .Z(n5063) );
  IV U8586 ( .A(n5401), .Z(n5061) );
  XNOR U8587 ( .A(n5596), .B(n5597), .Z(n5401) );
  NANDN U8588 ( .A(n5598), .B(n5599), .Z(n5597) );
  AND U8589 ( .A(b[2]), .B(a[97]), .Z(n5595) );
  XOR U8590 ( .A(n5055), .B(n5600), .Z(n5058) );
  NAND U8591 ( .A(b[1]), .B(a[98]), .Z(n5600) );
  OR U8592 ( .A(n5068), .B(n5066), .Z(n5055) );
  XOR U8593 ( .A(n5599), .B(n5598), .Z(n5066) );
  XOR U8594 ( .A(n5596), .B(n5593), .Z(n5601) );
  XOR U8595 ( .A(n5588), .B(n5592), .Z(n5602) );
  XOR U8596 ( .A(n5583), .B(n5587), .Z(n5603) );
  XOR U8597 ( .A(n5578), .B(n5582), .Z(n5604) );
  XOR U8598 ( .A(n5573), .B(n5577), .Z(n5605) );
  XOR U8599 ( .A(n5568), .B(n5572), .Z(n5606) );
  XOR U8600 ( .A(n5563), .B(n5567), .Z(n5607) );
  XOR U8601 ( .A(n5558), .B(n5562), .Z(n5608) );
  XOR U8602 ( .A(n5553), .B(n5557), .Z(n5609) );
  XOR U8603 ( .A(n5548), .B(n5552), .Z(n5610) );
  XOR U8604 ( .A(n5543), .B(n5547), .Z(n5611) );
  XOR U8605 ( .A(n5538), .B(n5542), .Z(n5612) );
  XOR U8606 ( .A(n5533), .B(n5537), .Z(n5613) );
  XOR U8607 ( .A(n5528), .B(n5532), .Z(n5614) );
  XOR U8608 ( .A(n5523), .B(n5527), .Z(n5615) );
  XOR U8609 ( .A(n5518), .B(n5522), .Z(n5616) );
  XOR U8610 ( .A(n5513), .B(n5517), .Z(n5617) );
  XOR U8611 ( .A(n5508), .B(n5512), .Z(n5618) );
  XOR U8612 ( .A(n5503), .B(n5507), .Z(n5619) );
  XOR U8613 ( .A(n5498), .B(n5502), .Z(n5620) );
  XOR U8614 ( .A(n5493), .B(n5497), .Z(n5621) );
  XOR U8615 ( .A(n5488), .B(n5492), .Z(n5622) );
  XOR U8616 ( .A(n5483), .B(n5487), .Z(n5623) );
  XOR U8617 ( .A(n5478), .B(n5482), .Z(n5624) );
  XOR U8618 ( .A(n5473), .B(n5477), .Z(n5625) );
  XOR U8619 ( .A(n5468), .B(n5472), .Z(n5626) );
  XNOR U8620 ( .A(n5464), .B(n5467), .Z(n5627) );
  XOR U8621 ( .A(n5628), .B(n5629), .Z(n5464) );
  XOR U8622 ( .A(n5630), .B(n5631), .Z(n5629) );
  XNOR U8623 ( .A(n5632), .B(n5633), .Z(n5630) );
  XOR U8624 ( .A(n5634), .B(n5635), .Z(n5633) );
  AND U8625 ( .A(b[30]), .B(a[68]), .Z(n5635) );
  AND U8626 ( .A(a[67]), .B(b[31]), .Z(n5634) );
  XNOR U8627 ( .A(n5636), .B(n5632), .Z(n5628) );
  XNOR U8628 ( .A(n5637), .B(n5638), .Z(n5632) );
  ANDN U8629 ( .B(n5639), .A(n5640), .Z(n5637) );
  AND U8630 ( .A(a[69]), .B(b[29]), .Z(n5636) );
  XOR U8631 ( .A(n5641), .B(n5462), .Z(n5463) );
  IV U8632 ( .A(n5631), .Z(n5462) );
  XOR U8633 ( .A(n5642), .B(n5643), .Z(n5631) );
  AND U8634 ( .A(n5644), .B(n5645), .Z(n5642) );
  AND U8635 ( .A(a[70]), .B(b[28]), .Z(n5641) );
  XOR U8636 ( .A(n5647), .B(n5648), .Z(n5467) );
  AND U8637 ( .A(n5649), .B(n5650), .Z(n5647) );
  AND U8638 ( .A(a[71]), .B(b[27]), .Z(n5646) );
  XOR U8639 ( .A(n5652), .B(n5653), .Z(n5472) );
  AND U8640 ( .A(n5654), .B(n5655), .Z(n5652) );
  AND U8641 ( .A(a[72]), .B(b[26]), .Z(n5651) );
  XOR U8642 ( .A(n5657), .B(n5658), .Z(n5477) );
  AND U8643 ( .A(n5659), .B(n5660), .Z(n5657) );
  AND U8644 ( .A(a[73]), .B(b[25]), .Z(n5656) );
  XOR U8645 ( .A(n5662), .B(n5663), .Z(n5482) );
  AND U8646 ( .A(n5664), .B(n5665), .Z(n5662) );
  AND U8647 ( .A(a[74]), .B(b[24]), .Z(n5661) );
  XOR U8648 ( .A(n5667), .B(n5668), .Z(n5487) );
  AND U8649 ( .A(n5669), .B(n5670), .Z(n5667) );
  AND U8650 ( .A(a[75]), .B(b[23]), .Z(n5666) );
  XOR U8651 ( .A(n5672), .B(n5673), .Z(n5492) );
  AND U8652 ( .A(n5674), .B(n5675), .Z(n5672) );
  AND U8653 ( .A(a[76]), .B(b[22]), .Z(n5671) );
  XOR U8654 ( .A(n5677), .B(n5678), .Z(n5497) );
  AND U8655 ( .A(n5679), .B(n5680), .Z(n5677) );
  AND U8656 ( .A(a[77]), .B(b[21]), .Z(n5676) );
  XOR U8657 ( .A(n5682), .B(n5683), .Z(n5502) );
  AND U8658 ( .A(n5684), .B(n5685), .Z(n5682) );
  AND U8659 ( .A(a[78]), .B(b[20]), .Z(n5681) );
  XOR U8660 ( .A(n5687), .B(n5688), .Z(n5507) );
  AND U8661 ( .A(n5689), .B(n5690), .Z(n5687) );
  AND U8662 ( .A(a[79]), .B(b[19]), .Z(n5686) );
  XOR U8663 ( .A(n5692), .B(n5693), .Z(n5512) );
  AND U8664 ( .A(n5694), .B(n5695), .Z(n5692) );
  AND U8665 ( .A(a[80]), .B(b[18]), .Z(n5691) );
  XOR U8666 ( .A(n5697), .B(n5698), .Z(n5517) );
  AND U8667 ( .A(n5699), .B(n5700), .Z(n5697) );
  AND U8668 ( .A(a[81]), .B(b[17]), .Z(n5696) );
  XOR U8669 ( .A(n5702), .B(n5703), .Z(n5522) );
  AND U8670 ( .A(n5704), .B(n5705), .Z(n5702) );
  AND U8671 ( .A(a[82]), .B(b[16]), .Z(n5701) );
  XOR U8672 ( .A(n5707), .B(n5708), .Z(n5527) );
  AND U8673 ( .A(n5709), .B(n5710), .Z(n5707) );
  AND U8674 ( .A(a[83]), .B(b[15]), .Z(n5706) );
  XOR U8675 ( .A(n5712), .B(n5713), .Z(n5532) );
  AND U8676 ( .A(n5714), .B(n5715), .Z(n5712) );
  AND U8677 ( .A(a[84]), .B(b[14]), .Z(n5711) );
  XOR U8678 ( .A(n5717), .B(n5718), .Z(n5537) );
  AND U8679 ( .A(n5719), .B(n5720), .Z(n5717) );
  AND U8680 ( .A(a[85]), .B(b[13]), .Z(n5716) );
  XOR U8681 ( .A(n5722), .B(n5723), .Z(n5542) );
  AND U8682 ( .A(n5724), .B(n5725), .Z(n5722) );
  AND U8683 ( .A(a[86]), .B(b[12]), .Z(n5721) );
  XOR U8684 ( .A(n5727), .B(n5728), .Z(n5547) );
  AND U8685 ( .A(n5729), .B(n5730), .Z(n5727) );
  AND U8686 ( .A(a[87]), .B(b[11]), .Z(n5726) );
  XOR U8687 ( .A(n5732), .B(n5733), .Z(n5552) );
  AND U8688 ( .A(n5734), .B(n5735), .Z(n5732) );
  AND U8689 ( .A(a[88]), .B(b[10]), .Z(n5731) );
  XOR U8690 ( .A(n5737), .B(n5738), .Z(n5557) );
  AND U8691 ( .A(n5739), .B(n5740), .Z(n5737) );
  AND U8692 ( .A(a[89]), .B(b[9]), .Z(n5736) );
  XOR U8693 ( .A(n5742), .B(n5743), .Z(n5562) );
  AND U8694 ( .A(n5744), .B(n5745), .Z(n5742) );
  AND U8695 ( .A(a[90]), .B(b[8]), .Z(n5741) );
  XOR U8696 ( .A(n5747), .B(n5748), .Z(n5567) );
  AND U8697 ( .A(n5749), .B(n5750), .Z(n5747) );
  AND U8698 ( .A(a[91]), .B(b[7]), .Z(n5746) );
  XOR U8699 ( .A(n5752), .B(n5753), .Z(n5572) );
  AND U8700 ( .A(n5754), .B(n5755), .Z(n5752) );
  AND U8701 ( .A(a[92]), .B(b[6]), .Z(n5751) );
  XOR U8702 ( .A(n5757), .B(n5758), .Z(n5577) );
  AND U8703 ( .A(n5759), .B(n5760), .Z(n5757) );
  AND U8704 ( .A(a[93]), .B(b[5]), .Z(n5756) );
  XOR U8705 ( .A(n5762), .B(n5763), .Z(n5582) );
  AND U8706 ( .A(n5764), .B(n5765), .Z(n5762) );
  AND U8707 ( .A(a[94]), .B(b[4]), .Z(n5761) );
  XOR U8708 ( .A(n5767), .B(n5768), .Z(n5587) );
  AND U8709 ( .A(n5769), .B(n5770), .Z(n5767) );
  AND U8710 ( .A(b[3]), .B(a[95]), .Z(n5766) );
  XOR U8711 ( .A(n5772), .B(n5773), .Z(n5592) );
  NANDN U8712 ( .A(n5774), .B(n5775), .Z(n5773) );
  AND U8713 ( .A(b[2]), .B(a[96]), .Z(n5771) );
  XOR U8714 ( .A(n5596), .B(n5776), .Z(n5599) );
  NAND U8715 ( .A(b[1]), .B(a[97]), .Z(n5776) );
  OR U8716 ( .A(n5071), .B(n5069), .Z(n5596) );
  XOR U8717 ( .A(n5775), .B(n5774), .Z(n5069) );
  XOR U8718 ( .A(n5778), .B(n5769), .Z(n5777) );
  XOR U8719 ( .A(n5764), .B(n5768), .Z(n5779) );
  XOR U8720 ( .A(n5759), .B(n5763), .Z(n5780) );
  XOR U8721 ( .A(n5754), .B(n5758), .Z(n5781) );
  XOR U8722 ( .A(n5749), .B(n5753), .Z(n5782) );
  XOR U8723 ( .A(n5744), .B(n5748), .Z(n5783) );
  XOR U8724 ( .A(n5739), .B(n5743), .Z(n5784) );
  XOR U8725 ( .A(n5734), .B(n5738), .Z(n5785) );
  XOR U8726 ( .A(n5729), .B(n5733), .Z(n5786) );
  XOR U8727 ( .A(n5724), .B(n5728), .Z(n5787) );
  XOR U8728 ( .A(n5719), .B(n5723), .Z(n5788) );
  XOR U8729 ( .A(n5714), .B(n5718), .Z(n5789) );
  XOR U8730 ( .A(n5709), .B(n5713), .Z(n5790) );
  XOR U8731 ( .A(n5704), .B(n5708), .Z(n5791) );
  XOR U8732 ( .A(n5699), .B(n5703), .Z(n5792) );
  XOR U8733 ( .A(n5694), .B(n5698), .Z(n5793) );
  XOR U8734 ( .A(n5689), .B(n5693), .Z(n5794) );
  XOR U8735 ( .A(n5684), .B(n5688), .Z(n5795) );
  XOR U8736 ( .A(n5679), .B(n5683), .Z(n5796) );
  XOR U8737 ( .A(n5674), .B(n5678), .Z(n5797) );
  XOR U8738 ( .A(n5669), .B(n5673), .Z(n5798) );
  XOR U8739 ( .A(n5664), .B(n5668), .Z(n5799) );
  XOR U8740 ( .A(n5659), .B(n5663), .Z(n5800) );
  XOR U8741 ( .A(n5654), .B(n5658), .Z(n5801) );
  XOR U8742 ( .A(n5649), .B(n5653), .Z(n5802) );
  XOR U8743 ( .A(n5644), .B(n5648), .Z(n5803) );
  XNOR U8744 ( .A(n5640), .B(n5643), .Z(n5804) );
  XOR U8745 ( .A(n5805), .B(n5806), .Z(n5640) );
  XOR U8746 ( .A(n5807), .B(n5808), .Z(n5806) );
  XOR U8747 ( .A(n5809), .B(n5810), .Z(n5807) );
  AND U8748 ( .A(b[29]), .B(a[68]), .Z(n5809) );
  XOR U8749 ( .A(n5810), .B(n5811), .Z(n5805) );
  XOR U8750 ( .A(n5812), .B(n5813), .Z(n5811) );
  AND U8751 ( .A(a[67]), .B(b[30]), .Z(n5813) );
  AND U8752 ( .A(a[66]), .B(b[31]), .Z(n5812) );
  XOR U8753 ( .A(n5814), .B(n5815), .Z(n5810) );
  ANDN U8754 ( .B(n5816), .A(n5817), .Z(n5814) );
  XOR U8755 ( .A(n5818), .B(n5638), .Z(n5639) );
  IV U8756 ( .A(n5808), .Z(n5638) );
  XOR U8757 ( .A(n5819), .B(n5820), .Z(n5808) );
  ANDN U8758 ( .B(n5821), .A(n5822), .Z(n5819) );
  AND U8759 ( .A(a[69]), .B(b[28]), .Z(n5818) );
  XOR U8760 ( .A(n5824), .B(n5825), .Z(n5643) );
  AND U8761 ( .A(n5826), .B(n5827), .Z(n5824) );
  AND U8762 ( .A(a[70]), .B(b[27]), .Z(n5823) );
  XOR U8763 ( .A(n5829), .B(n5830), .Z(n5648) );
  AND U8764 ( .A(n5831), .B(n5832), .Z(n5829) );
  AND U8765 ( .A(a[71]), .B(b[26]), .Z(n5828) );
  XOR U8766 ( .A(n5834), .B(n5835), .Z(n5653) );
  AND U8767 ( .A(n5836), .B(n5837), .Z(n5834) );
  AND U8768 ( .A(a[72]), .B(b[25]), .Z(n5833) );
  XOR U8769 ( .A(n5839), .B(n5840), .Z(n5658) );
  AND U8770 ( .A(n5841), .B(n5842), .Z(n5839) );
  AND U8771 ( .A(a[73]), .B(b[24]), .Z(n5838) );
  XOR U8772 ( .A(n5844), .B(n5845), .Z(n5663) );
  AND U8773 ( .A(n5846), .B(n5847), .Z(n5844) );
  AND U8774 ( .A(a[74]), .B(b[23]), .Z(n5843) );
  XOR U8775 ( .A(n5849), .B(n5850), .Z(n5668) );
  AND U8776 ( .A(n5851), .B(n5852), .Z(n5849) );
  AND U8777 ( .A(a[75]), .B(b[22]), .Z(n5848) );
  XOR U8778 ( .A(n5854), .B(n5855), .Z(n5673) );
  AND U8779 ( .A(n5856), .B(n5857), .Z(n5854) );
  AND U8780 ( .A(a[76]), .B(b[21]), .Z(n5853) );
  XOR U8781 ( .A(n5859), .B(n5860), .Z(n5678) );
  AND U8782 ( .A(n5861), .B(n5862), .Z(n5859) );
  AND U8783 ( .A(a[77]), .B(b[20]), .Z(n5858) );
  XOR U8784 ( .A(n5864), .B(n5865), .Z(n5683) );
  AND U8785 ( .A(n5866), .B(n5867), .Z(n5864) );
  AND U8786 ( .A(a[78]), .B(b[19]), .Z(n5863) );
  XOR U8787 ( .A(n5869), .B(n5870), .Z(n5688) );
  AND U8788 ( .A(n5871), .B(n5872), .Z(n5869) );
  AND U8789 ( .A(a[79]), .B(b[18]), .Z(n5868) );
  XOR U8790 ( .A(n5874), .B(n5875), .Z(n5693) );
  AND U8791 ( .A(n5876), .B(n5877), .Z(n5874) );
  AND U8792 ( .A(a[80]), .B(b[17]), .Z(n5873) );
  XOR U8793 ( .A(n5879), .B(n5880), .Z(n5698) );
  AND U8794 ( .A(n5881), .B(n5882), .Z(n5879) );
  AND U8795 ( .A(a[81]), .B(b[16]), .Z(n5878) );
  XOR U8796 ( .A(n5884), .B(n5885), .Z(n5703) );
  AND U8797 ( .A(n5886), .B(n5887), .Z(n5884) );
  AND U8798 ( .A(a[82]), .B(b[15]), .Z(n5883) );
  XOR U8799 ( .A(n5889), .B(n5890), .Z(n5708) );
  AND U8800 ( .A(n5891), .B(n5892), .Z(n5889) );
  AND U8801 ( .A(a[83]), .B(b[14]), .Z(n5888) );
  XOR U8802 ( .A(n5894), .B(n5895), .Z(n5713) );
  AND U8803 ( .A(n5896), .B(n5897), .Z(n5894) );
  AND U8804 ( .A(a[84]), .B(b[13]), .Z(n5893) );
  XOR U8805 ( .A(n5899), .B(n5900), .Z(n5718) );
  AND U8806 ( .A(n5901), .B(n5902), .Z(n5899) );
  AND U8807 ( .A(a[85]), .B(b[12]), .Z(n5898) );
  XOR U8808 ( .A(n5904), .B(n5905), .Z(n5723) );
  AND U8809 ( .A(n5906), .B(n5907), .Z(n5904) );
  AND U8810 ( .A(a[86]), .B(b[11]), .Z(n5903) );
  XOR U8811 ( .A(n5909), .B(n5910), .Z(n5728) );
  AND U8812 ( .A(n5911), .B(n5912), .Z(n5909) );
  AND U8813 ( .A(a[87]), .B(b[10]), .Z(n5908) );
  XOR U8814 ( .A(n5914), .B(n5915), .Z(n5733) );
  AND U8815 ( .A(n5916), .B(n5917), .Z(n5914) );
  AND U8816 ( .A(a[88]), .B(b[9]), .Z(n5913) );
  XOR U8817 ( .A(n5919), .B(n5920), .Z(n5738) );
  AND U8818 ( .A(n5921), .B(n5922), .Z(n5919) );
  AND U8819 ( .A(a[89]), .B(b[8]), .Z(n5918) );
  XOR U8820 ( .A(n5924), .B(n5925), .Z(n5743) );
  AND U8821 ( .A(n5926), .B(n5927), .Z(n5924) );
  AND U8822 ( .A(a[90]), .B(b[7]), .Z(n5923) );
  XOR U8823 ( .A(n5929), .B(n5930), .Z(n5748) );
  AND U8824 ( .A(n5931), .B(n5932), .Z(n5929) );
  AND U8825 ( .A(a[91]), .B(b[6]), .Z(n5928) );
  XOR U8826 ( .A(n5934), .B(n5935), .Z(n5753) );
  AND U8827 ( .A(n5936), .B(n5937), .Z(n5934) );
  AND U8828 ( .A(a[92]), .B(b[5]), .Z(n5933) );
  XOR U8829 ( .A(n5939), .B(n5940), .Z(n5758) );
  AND U8830 ( .A(n5941), .B(n5942), .Z(n5939) );
  AND U8831 ( .A(a[93]), .B(b[4]), .Z(n5938) );
  XOR U8832 ( .A(n5944), .B(n5945), .Z(n5763) );
  AND U8833 ( .A(n5946), .B(n5947), .Z(n5944) );
  AND U8834 ( .A(a[94]), .B(b[3]), .Z(n5943) );
  IV U8835 ( .A(n5772), .Z(n5778) );
  XOR U8836 ( .A(n5949), .B(n5950), .Z(n5768) );
  OR U8837 ( .A(n5951), .B(n5952), .Z(n5950) );
  AND U8838 ( .A(b[2]), .B(a[95]), .Z(n5948) );
  XNOR U8839 ( .A(n5772), .B(n5953), .Z(n5775) );
  NAND U8840 ( .A(b[1]), .B(a[96]), .Z(n5953) );
  ANDN U8841 ( .B(n5072), .A(n5074), .Z(n5772) );
  NAND U8842 ( .A(a[96]), .B(b[0]), .Z(n5074) );
  XOR U8843 ( .A(n5951), .B(n5952), .Z(n5072) );
  XOR U8844 ( .A(n5955), .B(n5946), .Z(n5954) );
  XOR U8845 ( .A(n5941), .B(n5945), .Z(n5956) );
  XOR U8846 ( .A(n5936), .B(n5940), .Z(n5957) );
  XOR U8847 ( .A(n5931), .B(n5935), .Z(n5958) );
  XOR U8848 ( .A(n5926), .B(n5930), .Z(n5959) );
  XOR U8849 ( .A(n5921), .B(n5925), .Z(n5960) );
  XOR U8850 ( .A(n5916), .B(n5920), .Z(n5961) );
  XOR U8851 ( .A(n5911), .B(n5915), .Z(n5962) );
  XOR U8852 ( .A(n5906), .B(n5910), .Z(n5963) );
  XOR U8853 ( .A(n5901), .B(n5905), .Z(n5964) );
  XOR U8854 ( .A(n5896), .B(n5900), .Z(n5965) );
  XOR U8855 ( .A(n5891), .B(n5895), .Z(n5966) );
  XOR U8856 ( .A(n5886), .B(n5890), .Z(n5967) );
  XOR U8857 ( .A(n5881), .B(n5885), .Z(n5968) );
  XOR U8858 ( .A(n5876), .B(n5880), .Z(n5969) );
  XOR U8859 ( .A(n5871), .B(n5875), .Z(n5970) );
  XOR U8860 ( .A(n5866), .B(n5870), .Z(n5971) );
  XOR U8861 ( .A(n5861), .B(n5865), .Z(n5972) );
  XOR U8862 ( .A(n5856), .B(n5860), .Z(n5973) );
  XOR U8863 ( .A(n5851), .B(n5855), .Z(n5974) );
  XOR U8864 ( .A(n5846), .B(n5850), .Z(n5975) );
  XOR U8865 ( .A(n5841), .B(n5845), .Z(n5976) );
  XOR U8866 ( .A(n5836), .B(n5840), .Z(n5977) );
  XOR U8867 ( .A(n5831), .B(n5835), .Z(n5978) );
  XOR U8868 ( .A(n5826), .B(n5830), .Z(n5979) );
  XNOR U8869 ( .A(n5822), .B(n5825), .Z(n5980) );
  XNOR U8870 ( .A(n5817), .B(n5981), .Z(n5822) );
  XOR U8871 ( .A(n5816), .B(n5820), .Z(n5981) );
  XOR U8872 ( .A(n5982), .B(n5815), .Z(n5816) );
  AND U8873 ( .A(b[28]), .B(a[68]), .Z(n5982) );
  XOR U8874 ( .A(n5983), .B(n5984), .Z(n5817) );
  XOR U8875 ( .A(n5815), .B(n5985), .Z(n5984) );
  XOR U8876 ( .A(n5986), .B(n5987), .Z(n5985) );
  XOR U8877 ( .A(n5988), .B(n5989), .Z(n5987) );
  NAND U8878 ( .A(a[66]), .B(b[30]), .Z(n5989) );
  AND U8879 ( .A(a[65]), .B(b[31]), .Z(n5988) );
  XOR U8880 ( .A(n5990), .B(n5991), .Z(n5815) );
  AND U8881 ( .A(n5992), .B(n5993), .Z(n5990) );
  XOR U8882 ( .A(n5994), .B(n5986), .Z(n5983) );
  XOR U8883 ( .A(n5995), .B(n5996), .Z(n5986) );
  ANDN U8884 ( .B(n5997), .A(n5998), .Z(n5995) );
  AND U8885 ( .A(a[67]), .B(b[29]), .Z(n5994) );
  XOR U8886 ( .A(n6000), .B(n6001), .Z(n5820) );
  AND U8887 ( .A(n6002), .B(n6003), .Z(n6000) );
  AND U8888 ( .A(a[69]), .B(b[27]), .Z(n5999) );
  XOR U8889 ( .A(n6005), .B(n6006), .Z(n5825) );
  AND U8890 ( .A(n6007), .B(n6008), .Z(n6005) );
  AND U8891 ( .A(a[70]), .B(b[26]), .Z(n6004) );
  XOR U8892 ( .A(n6010), .B(n6011), .Z(n5830) );
  AND U8893 ( .A(n6012), .B(n6013), .Z(n6010) );
  AND U8894 ( .A(a[71]), .B(b[25]), .Z(n6009) );
  XOR U8895 ( .A(n6015), .B(n6016), .Z(n5835) );
  AND U8896 ( .A(n6017), .B(n6018), .Z(n6015) );
  AND U8897 ( .A(a[72]), .B(b[24]), .Z(n6014) );
  XOR U8898 ( .A(n6020), .B(n6021), .Z(n5840) );
  AND U8899 ( .A(n6022), .B(n6023), .Z(n6020) );
  AND U8900 ( .A(a[73]), .B(b[23]), .Z(n6019) );
  XOR U8901 ( .A(n6025), .B(n6026), .Z(n5845) );
  AND U8902 ( .A(n6027), .B(n6028), .Z(n6025) );
  AND U8903 ( .A(a[74]), .B(b[22]), .Z(n6024) );
  XOR U8904 ( .A(n6030), .B(n6031), .Z(n5850) );
  AND U8905 ( .A(n6032), .B(n6033), .Z(n6030) );
  AND U8906 ( .A(a[75]), .B(b[21]), .Z(n6029) );
  XOR U8907 ( .A(n6035), .B(n6036), .Z(n5855) );
  AND U8908 ( .A(n6037), .B(n6038), .Z(n6035) );
  AND U8909 ( .A(a[76]), .B(b[20]), .Z(n6034) );
  XOR U8910 ( .A(n6040), .B(n6041), .Z(n5860) );
  AND U8911 ( .A(n6042), .B(n6043), .Z(n6040) );
  AND U8912 ( .A(a[77]), .B(b[19]), .Z(n6039) );
  XOR U8913 ( .A(n6045), .B(n6046), .Z(n5865) );
  AND U8914 ( .A(n6047), .B(n6048), .Z(n6045) );
  AND U8915 ( .A(a[78]), .B(b[18]), .Z(n6044) );
  XOR U8916 ( .A(n6050), .B(n6051), .Z(n5870) );
  AND U8917 ( .A(n6052), .B(n6053), .Z(n6050) );
  AND U8918 ( .A(a[79]), .B(b[17]), .Z(n6049) );
  XOR U8919 ( .A(n6055), .B(n6056), .Z(n5875) );
  AND U8920 ( .A(n6057), .B(n6058), .Z(n6055) );
  AND U8921 ( .A(a[80]), .B(b[16]), .Z(n6054) );
  XOR U8922 ( .A(n6060), .B(n6061), .Z(n5880) );
  AND U8923 ( .A(n6062), .B(n6063), .Z(n6060) );
  AND U8924 ( .A(a[81]), .B(b[15]), .Z(n6059) );
  XOR U8925 ( .A(n6065), .B(n6066), .Z(n5885) );
  AND U8926 ( .A(n6067), .B(n6068), .Z(n6065) );
  AND U8927 ( .A(a[82]), .B(b[14]), .Z(n6064) );
  XOR U8928 ( .A(n6070), .B(n6071), .Z(n5890) );
  AND U8929 ( .A(n6072), .B(n6073), .Z(n6070) );
  AND U8930 ( .A(a[83]), .B(b[13]), .Z(n6069) );
  XOR U8931 ( .A(n6075), .B(n6076), .Z(n5895) );
  AND U8932 ( .A(n6077), .B(n6078), .Z(n6075) );
  AND U8933 ( .A(a[84]), .B(b[12]), .Z(n6074) );
  XOR U8934 ( .A(n6080), .B(n6081), .Z(n5900) );
  AND U8935 ( .A(n6082), .B(n6083), .Z(n6080) );
  AND U8936 ( .A(a[85]), .B(b[11]), .Z(n6079) );
  XOR U8937 ( .A(n6085), .B(n6086), .Z(n5905) );
  AND U8938 ( .A(n6087), .B(n6088), .Z(n6085) );
  AND U8939 ( .A(a[86]), .B(b[10]), .Z(n6084) );
  XOR U8940 ( .A(n6090), .B(n6091), .Z(n5910) );
  AND U8941 ( .A(n6092), .B(n6093), .Z(n6090) );
  AND U8942 ( .A(a[87]), .B(b[9]), .Z(n6089) );
  XOR U8943 ( .A(n6095), .B(n6096), .Z(n5915) );
  AND U8944 ( .A(n6097), .B(n6098), .Z(n6095) );
  AND U8945 ( .A(a[88]), .B(b[8]), .Z(n6094) );
  XOR U8946 ( .A(n6100), .B(n6101), .Z(n5920) );
  AND U8947 ( .A(n6102), .B(n6103), .Z(n6100) );
  AND U8948 ( .A(a[89]), .B(b[7]), .Z(n6099) );
  XOR U8949 ( .A(n6105), .B(n6106), .Z(n5925) );
  AND U8950 ( .A(n6107), .B(n6108), .Z(n6105) );
  AND U8951 ( .A(a[90]), .B(b[6]), .Z(n6104) );
  XOR U8952 ( .A(n6110), .B(n6111), .Z(n5930) );
  AND U8953 ( .A(n6112), .B(n6113), .Z(n6110) );
  AND U8954 ( .A(a[91]), .B(b[5]), .Z(n6109) );
  XOR U8955 ( .A(n6115), .B(n6116), .Z(n5935) );
  AND U8956 ( .A(n6117), .B(n6118), .Z(n6115) );
  AND U8957 ( .A(a[92]), .B(b[4]), .Z(n6114) );
  XOR U8958 ( .A(n6120), .B(n6121), .Z(n5940) );
  AND U8959 ( .A(n6122), .B(n6123), .Z(n6120) );
  AND U8960 ( .A(a[93]), .B(b[3]), .Z(n6119) );
  XOR U8961 ( .A(n6125), .B(n6126), .Z(n5945) );
  OR U8962 ( .A(n6127), .B(n6128), .Z(n6126) );
  AND U8963 ( .A(a[94]), .B(b[2]), .Z(n6124) );
  XNOR U8964 ( .A(n5955), .B(n6129), .Z(n5951) );
  NAND U8965 ( .A(b[1]), .B(a[95]), .Z(n6129) );
  IV U8966 ( .A(n5949), .Z(n5955) );
  ANDN U8967 ( .B(n5077), .A(n5079), .Z(n5949) );
  NAND U8968 ( .A(a[95]), .B(b[0]), .Z(n5079) );
  XOR U8969 ( .A(n6127), .B(n6128), .Z(n5077) );
  XOR U8970 ( .A(n6131), .B(n6122), .Z(n6130) );
  XOR U8971 ( .A(n6117), .B(n6121), .Z(n6132) );
  XOR U8972 ( .A(n6112), .B(n6116), .Z(n6133) );
  XOR U8973 ( .A(n6107), .B(n6111), .Z(n6134) );
  XOR U8974 ( .A(n6102), .B(n6106), .Z(n6135) );
  XOR U8975 ( .A(n6097), .B(n6101), .Z(n6136) );
  XOR U8976 ( .A(n6092), .B(n6096), .Z(n6137) );
  XOR U8977 ( .A(n6087), .B(n6091), .Z(n6138) );
  XOR U8978 ( .A(n6082), .B(n6086), .Z(n6139) );
  XOR U8979 ( .A(n6077), .B(n6081), .Z(n6140) );
  XOR U8980 ( .A(n6072), .B(n6076), .Z(n6141) );
  XOR U8981 ( .A(n6067), .B(n6071), .Z(n6142) );
  XOR U8982 ( .A(n6062), .B(n6066), .Z(n6143) );
  XOR U8983 ( .A(n6057), .B(n6061), .Z(n6144) );
  XOR U8984 ( .A(n6052), .B(n6056), .Z(n6145) );
  XOR U8985 ( .A(n6047), .B(n6051), .Z(n6146) );
  XOR U8986 ( .A(n6042), .B(n6046), .Z(n6147) );
  XOR U8987 ( .A(n6037), .B(n6041), .Z(n6148) );
  XOR U8988 ( .A(n6032), .B(n6036), .Z(n6149) );
  XOR U8989 ( .A(n6027), .B(n6031), .Z(n6150) );
  XOR U8990 ( .A(n6022), .B(n6026), .Z(n6151) );
  XOR U8991 ( .A(n6017), .B(n6021), .Z(n6152) );
  XOR U8992 ( .A(n6012), .B(n6016), .Z(n6153) );
  XOR U8993 ( .A(n6007), .B(n6011), .Z(n6154) );
  XOR U8994 ( .A(n6002), .B(n6006), .Z(n6155) );
  XOR U8995 ( .A(n5992), .B(n6001), .Z(n6156) );
  XOR U8996 ( .A(n6157), .B(n5991), .Z(n5992) );
  AND U8997 ( .A(b[27]), .B(a[68]), .Z(n6157) );
  XOR U8998 ( .A(n5991), .B(n5998), .Z(n6158) );
  XOR U8999 ( .A(n6159), .B(n6160), .Z(n5998) );
  XOR U9000 ( .A(n5996), .B(n6161), .Z(n6160) );
  XOR U9001 ( .A(n6162), .B(n6163), .Z(n6161) );
  XOR U9002 ( .A(n6164), .B(n6165), .Z(n6163) );
  NAND U9003 ( .A(a[65]), .B(b[30]), .Z(n6165) );
  AND U9004 ( .A(a[64]), .B(b[31]), .Z(n6164) );
  XOR U9005 ( .A(n6166), .B(n6162), .Z(n6159) );
  XOR U9006 ( .A(n6167), .B(n6168), .Z(n6162) );
  ANDN U9007 ( .B(n6169), .A(n6170), .Z(n6167) );
  AND U9008 ( .A(a[66]), .B(b[29]), .Z(n6166) );
  XOR U9009 ( .A(n6171), .B(n6172), .Z(n5991) );
  AND U9010 ( .A(n6173), .B(n6174), .Z(n6171) );
  XOR U9011 ( .A(n6175), .B(n5996), .Z(n5997) );
  XOR U9012 ( .A(n6176), .B(n6177), .Z(n5996) );
  AND U9013 ( .A(n6178), .B(n6179), .Z(n6176) );
  AND U9014 ( .A(a[67]), .B(b[28]), .Z(n6175) );
  XOR U9015 ( .A(n6181), .B(n6182), .Z(n6001) );
  AND U9016 ( .A(n6183), .B(n6184), .Z(n6181) );
  AND U9017 ( .A(a[69]), .B(b[26]), .Z(n6180) );
  XOR U9018 ( .A(n6186), .B(n6187), .Z(n6006) );
  AND U9019 ( .A(n6188), .B(n6189), .Z(n6186) );
  AND U9020 ( .A(a[70]), .B(b[25]), .Z(n6185) );
  XOR U9021 ( .A(n6191), .B(n6192), .Z(n6011) );
  AND U9022 ( .A(n6193), .B(n6194), .Z(n6191) );
  AND U9023 ( .A(a[71]), .B(b[24]), .Z(n6190) );
  XOR U9024 ( .A(n6196), .B(n6197), .Z(n6016) );
  AND U9025 ( .A(n6198), .B(n6199), .Z(n6196) );
  AND U9026 ( .A(a[72]), .B(b[23]), .Z(n6195) );
  XOR U9027 ( .A(n6201), .B(n6202), .Z(n6021) );
  AND U9028 ( .A(n6203), .B(n6204), .Z(n6201) );
  AND U9029 ( .A(a[73]), .B(b[22]), .Z(n6200) );
  XOR U9030 ( .A(n6206), .B(n6207), .Z(n6026) );
  AND U9031 ( .A(n6208), .B(n6209), .Z(n6206) );
  AND U9032 ( .A(a[74]), .B(b[21]), .Z(n6205) );
  XOR U9033 ( .A(n6211), .B(n6212), .Z(n6031) );
  AND U9034 ( .A(n6213), .B(n6214), .Z(n6211) );
  AND U9035 ( .A(a[75]), .B(b[20]), .Z(n6210) );
  XOR U9036 ( .A(n6216), .B(n6217), .Z(n6036) );
  AND U9037 ( .A(n6218), .B(n6219), .Z(n6216) );
  AND U9038 ( .A(a[76]), .B(b[19]), .Z(n6215) );
  XOR U9039 ( .A(n6221), .B(n6222), .Z(n6041) );
  AND U9040 ( .A(n6223), .B(n6224), .Z(n6221) );
  AND U9041 ( .A(a[77]), .B(b[18]), .Z(n6220) );
  XOR U9042 ( .A(n6226), .B(n6227), .Z(n6046) );
  AND U9043 ( .A(n6228), .B(n6229), .Z(n6226) );
  AND U9044 ( .A(a[78]), .B(b[17]), .Z(n6225) );
  XOR U9045 ( .A(n6231), .B(n6232), .Z(n6051) );
  AND U9046 ( .A(n6233), .B(n6234), .Z(n6231) );
  AND U9047 ( .A(a[79]), .B(b[16]), .Z(n6230) );
  XOR U9048 ( .A(n6236), .B(n6237), .Z(n6056) );
  AND U9049 ( .A(n6238), .B(n6239), .Z(n6236) );
  AND U9050 ( .A(a[80]), .B(b[15]), .Z(n6235) );
  XOR U9051 ( .A(n6241), .B(n6242), .Z(n6061) );
  AND U9052 ( .A(n6243), .B(n6244), .Z(n6241) );
  AND U9053 ( .A(a[81]), .B(b[14]), .Z(n6240) );
  XOR U9054 ( .A(n6246), .B(n6247), .Z(n6066) );
  AND U9055 ( .A(n6248), .B(n6249), .Z(n6246) );
  AND U9056 ( .A(a[82]), .B(b[13]), .Z(n6245) );
  XOR U9057 ( .A(n6251), .B(n6252), .Z(n6071) );
  AND U9058 ( .A(n6253), .B(n6254), .Z(n6251) );
  AND U9059 ( .A(a[83]), .B(b[12]), .Z(n6250) );
  XOR U9060 ( .A(n6256), .B(n6257), .Z(n6076) );
  AND U9061 ( .A(n6258), .B(n6259), .Z(n6256) );
  AND U9062 ( .A(a[84]), .B(b[11]), .Z(n6255) );
  XOR U9063 ( .A(n6261), .B(n6262), .Z(n6081) );
  AND U9064 ( .A(n6263), .B(n6264), .Z(n6261) );
  AND U9065 ( .A(a[85]), .B(b[10]), .Z(n6260) );
  XOR U9066 ( .A(n6266), .B(n6267), .Z(n6086) );
  AND U9067 ( .A(n6268), .B(n6269), .Z(n6266) );
  AND U9068 ( .A(a[86]), .B(b[9]), .Z(n6265) );
  XOR U9069 ( .A(n6271), .B(n6272), .Z(n6091) );
  AND U9070 ( .A(n6273), .B(n6274), .Z(n6271) );
  AND U9071 ( .A(a[87]), .B(b[8]), .Z(n6270) );
  XOR U9072 ( .A(n6276), .B(n6277), .Z(n6096) );
  AND U9073 ( .A(n6278), .B(n6279), .Z(n6276) );
  AND U9074 ( .A(a[88]), .B(b[7]), .Z(n6275) );
  XOR U9075 ( .A(n6281), .B(n6282), .Z(n6101) );
  AND U9076 ( .A(n6283), .B(n6284), .Z(n6281) );
  AND U9077 ( .A(a[89]), .B(b[6]), .Z(n6280) );
  XOR U9078 ( .A(n6286), .B(n6287), .Z(n6106) );
  AND U9079 ( .A(n6288), .B(n6289), .Z(n6286) );
  AND U9080 ( .A(a[90]), .B(b[5]), .Z(n6285) );
  XOR U9081 ( .A(n6291), .B(n6292), .Z(n6111) );
  AND U9082 ( .A(n6293), .B(n6294), .Z(n6291) );
  AND U9083 ( .A(a[91]), .B(b[4]), .Z(n6290) );
  XOR U9084 ( .A(n6296), .B(n6297), .Z(n6116) );
  AND U9085 ( .A(n6298), .B(n6299), .Z(n6296) );
  AND U9086 ( .A(a[92]), .B(b[3]), .Z(n6295) );
  XOR U9087 ( .A(n6301), .B(n6302), .Z(n6121) );
  OR U9088 ( .A(n6303), .B(n6304), .Z(n6302) );
  AND U9089 ( .A(a[93]), .B(b[2]), .Z(n6300) );
  XNOR U9090 ( .A(n6131), .B(n6305), .Z(n6127) );
  NAND U9091 ( .A(a[94]), .B(b[1]), .Z(n6305) );
  IV U9092 ( .A(n6125), .Z(n6131) );
  ANDN U9093 ( .B(n5082), .A(n5084), .Z(n6125) );
  NAND U9094 ( .A(b[0]), .B(a[94]), .Z(n5084) );
  XOR U9095 ( .A(n6303), .B(n6304), .Z(n5082) );
  XOR U9096 ( .A(n6307), .B(n6298), .Z(n6306) );
  XOR U9097 ( .A(n6293), .B(n6297), .Z(n6308) );
  XOR U9098 ( .A(n6288), .B(n6292), .Z(n6309) );
  XOR U9099 ( .A(n6283), .B(n6287), .Z(n6310) );
  XOR U9100 ( .A(n6278), .B(n6282), .Z(n6311) );
  XOR U9101 ( .A(n6273), .B(n6277), .Z(n6312) );
  XOR U9102 ( .A(n6268), .B(n6272), .Z(n6313) );
  XOR U9103 ( .A(n6263), .B(n6267), .Z(n6314) );
  XOR U9104 ( .A(n6258), .B(n6262), .Z(n6315) );
  XOR U9105 ( .A(n6253), .B(n6257), .Z(n6316) );
  XOR U9106 ( .A(n6248), .B(n6252), .Z(n6317) );
  XOR U9107 ( .A(n6243), .B(n6247), .Z(n6318) );
  XOR U9108 ( .A(n6238), .B(n6242), .Z(n6319) );
  XOR U9109 ( .A(n6233), .B(n6237), .Z(n6320) );
  XOR U9110 ( .A(n6228), .B(n6232), .Z(n6321) );
  XOR U9111 ( .A(n6223), .B(n6227), .Z(n6322) );
  XOR U9112 ( .A(n6218), .B(n6222), .Z(n6323) );
  XOR U9113 ( .A(n6213), .B(n6217), .Z(n6324) );
  XOR U9114 ( .A(n6208), .B(n6212), .Z(n6325) );
  XOR U9115 ( .A(n6203), .B(n6207), .Z(n6326) );
  XOR U9116 ( .A(n6198), .B(n6202), .Z(n6327) );
  XOR U9117 ( .A(n6193), .B(n6197), .Z(n6328) );
  XOR U9118 ( .A(n6188), .B(n6192), .Z(n6329) );
  XOR U9119 ( .A(n6183), .B(n6187), .Z(n6330) );
  XOR U9120 ( .A(n6173), .B(n6182), .Z(n6331) );
  XOR U9121 ( .A(n6332), .B(n6172), .Z(n6173) );
  AND U9122 ( .A(b[26]), .B(a[68]), .Z(n6332) );
  XNOR U9123 ( .A(n6172), .B(n6178), .Z(n6333) );
  XOR U9124 ( .A(n6177), .B(n6170), .Z(n6334) );
  XOR U9125 ( .A(n6335), .B(n6336), .Z(n6170) );
  XOR U9126 ( .A(n6168), .B(n6337), .Z(n6336) );
  XOR U9127 ( .A(n6338), .B(n6339), .Z(n6337) );
  XOR U9128 ( .A(n6340), .B(n6341), .Z(n6339) );
  NAND U9129 ( .A(a[64]), .B(b[30]), .Z(n6341) );
  AND U9130 ( .A(a[63]), .B(b[31]), .Z(n6340) );
  XOR U9131 ( .A(n6342), .B(n6338), .Z(n6335) );
  XOR U9132 ( .A(n6343), .B(n6344), .Z(n6338) );
  ANDN U9133 ( .B(n6345), .A(n6346), .Z(n6343) );
  AND U9134 ( .A(a[65]), .B(b[29]), .Z(n6342) );
  XOR U9135 ( .A(n6347), .B(n6168), .Z(n6169) );
  XOR U9136 ( .A(n6348), .B(n6349), .Z(n6168) );
  AND U9137 ( .A(n6350), .B(n6351), .Z(n6348) );
  AND U9138 ( .A(a[66]), .B(b[28]), .Z(n6347) );
  XOR U9139 ( .A(n6352), .B(n6353), .Z(n6172) );
  AND U9140 ( .A(n6354), .B(n6355), .Z(n6352) );
  XOR U9141 ( .A(n6356), .B(n6177), .Z(n6179) );
  XOR U9142 ( .A(n6357), .B(n6358), .Z(n6177) );
  AND U9143 ( .A(n6359), .B(n6360), .Z(n6357) );
  AND U9144 ( .A(a[67]), .B(b[27]), .Z(n6356) );
  XOR U9145 ( .A(n6362), .B(n6363), .Z(n6182) );
  AND U9146 ( .A(n6364), .B(n6365), .Z(n6362) );
  AND U9147 ( .A(a[69]), .B(b[25]), .Z(n6361) );
  XOR U9148 ( .A(n6367), .B(n6368), .Z(n6187) );
  AND U9149 ( .A(n6369), .B(n6370), .Z(n6367) );
  AND U9150 ( .A(a[70]), .B(b[24]), .Z(n6366) );
  XOR U9151 ( .A(n6372), .B(n6373), .Z(n6192) );
  AND U9152 ( .A(n6374), .B(n6375), .Z(n6372) );
  AND U9153 ( .A(a[71]), .B(b[23]), .Z(n6371) );
  XOR U9154 ( .A(n6377), .B(n6378), .Z(n6197) );
  AND U9155 ( .A(n6379), .B(n6380), .Z(n6377) );
  AND U9156 ( .A(a[72]), .B(b[22]), .Z(n6376) );
  XOR U9157 ( .A(n6382), .B(n6383), .Z(n6202) );
  AND U9158 ( .A(n6384), .B(n6385), .Z(n6382) );
  AND U9159 ( .A(a[73]), .B(b[21]), .Z(n6381) );
  XOR U9160 ( .A(n6387), .B(n6388), .Z(n6207) );
  AND U9161 ( .A(n6389), .B(n6390), .Z(n6387) );
  AND U9162 ( .A(a[74]), .B(b[20]), .Z(n6386) );
  XOR U9163 ( .A(n6392), .B(n6393), .Z(n6212) );
  AND U9164 ( .A(n6394), .B(n6395), .Z(n6392) );
  AND U9165 ( .A(a[75]), .B(b[19]), .Z(n6391) );
  XOR U9166 ( .A(n6397), .B(n6398), .Z(n6217) );
  AND U9167 ( .A(n6399), .B(n6400), .Z(n6397) );
  AND U9168 ( .A(a[76]), .B(b[18]), .Z(n6396) );
  XOR U9169 ( .A(n6402), .B(n6403), .Z(n6222) );
  AND U9170 ( .A(n6404), .B(n6405), .Z(n6402) );
  AND U9171 ( .A(a[77]), .B(b[17]), .Z(n6401) );
  XOR U9172 ( .A(n6407), .B(n6408), .Z(n6227) );
  AND U9173 ( .A(n6409), .B(n6410), .Z(n6407) );
  AND U9174 ( .A(a[78]), .B(b[16]), .Z(n6406) );
  XOR U9175 ( .A(n6412), .B(n6413), .Z(n6232) );
  AND U9176 ( .A(n6414), .B(n6415), .Z(n6412) );
  AND U9177 ( .A(a[79]), .B(b[15]), .Z(n6411) );
  XOR U9178 ( .A(n6417), .B(n6418), .Z(n6237) );
  AND U9179 ( .A(n6419), .B(n6420), .Z(n6417) );
  AND U9180 ( .A(a[80]), .B(b[14]), .Z(n6416) );
  XOR U9181 ( .A(n6422), .B(n6423), .Z(n6242) );
  AND U9182 ( .A(n6424), .B(n6425), .Z(n6422) );
  AND U9183 ( .A(a[81]), .B(b[13]), .Z(n6421) );
  XOR U9184 ( .A(n6427), .B(n6428), .Z(n6247) );
  AND U9185 ( .A(n6429), .B(n6430), .Z(n6427) );
  AND U9186 ( .A(a[82]), .B(b[12]), .Z(n6426) );
  XOR U9187 ( .A(n6432), .B(n6433), .Z(n6252) );
  AND U9188 ( .A(n6434), .B(n6435), .Z(n6432) );
  AND U9189 ( .A(a[83]), .B(b[11]), .Z(n6431) );
  XOR U9190 ( .A(n6437), .B(n6438), .Z(n6257) );
  AND U9191 ( .A(n6439), .B(n6440), .Z(n6437) );
  AND U9192 ( .A(a[84]), .B(b[10]), .Z(n6436) );
  XOR U9193 ( .A(n6442), .B(n6443), .Z(n6262) );
  AND U9194 ( .A(n6444), .B(n6445), .Z(n6442) );
  AND U9195 ( .A(a[85]), .B(b[9]), .Z(n6441) );
  XOR U9196 ( .A(n6447), .B(n6448), .Z(n6267) );
  AND U9197 ( .A(n6449), .B(n6450), .Z(n6447) );
  AND U9198 ( .A(a[86]), .B(b[8]), .Z(n6446) );
  XOR U9199 ( .A(n6452), .B(n6453), .Z(n6272) );
  AND U9200 ( .A(n6454), .B(n6455), .Z(n6452) );
  AND U9201 ( .A(a[87]), .B(b[7]), .Z(n6451) );
  XOR U9202 ( .A(n6457), .B(n6458), .Z(n6277) );
  AND U9203 ( .A(n6459), .B(n6460), .Z(n6457) );
  AND U9204 ( .A(a[88]), .B(b[6]), .Z(n6456) );
  XOR U9205 ( .A(n6462), .B(n6463), .Z(n6282) );
  AND U9206 ( .A(n6464), .B(n6465), .Z(n6462) );
  AND U9207 ( .A(a[89]), .B(b[5]), .Z(n6461) );
  XOR U9208 ( .A(n6467), .B(n6468), .Z(n6287) );
  AND U9209 ( .A(n6469), .B(n6470), .Z(n6467) );
  AND U9210 ( .A(a[90]), .B(b[4]), .Z(n6466) );
  XOR U9211 ( .A(n6472), .B(n6473), .Z(n6292) );
  AND U9212 ( .A(n6474), .B(n6475), .Z(n6472) );
  AND U9213 ( .A(a[91]), .B(b[3]), .Z(n6471) );
  XOR U9214 ( .A(n6477), .B(n6478), .Z(n6297) );
  OR U9215 ( .A(n6479), .B(n6480), .Z(n6478) );
  AND U9216 ( .A(a[92]), .B(b[2]), .Z(n6476) );
  XNOR U9217 ( .A(n6307), .B(n6481), .Z(n6303) );
  NAND U9218 ( .A(a[93]), .B(b[1]), .Z(n6481) );
  IV U9219 ( .A(n6301), .Z(n6307) );
  ANDN U9220 ( .B(n5087), .A(n5089), .Z(n6301) );
  NAND U9221 ( .A(a[93]), .B(b[0]), .Z(n5089) );
  XOR U9222 ( .A(n6479), .B(n6480), .Z(n5087) );
  XOR U9223 ( .A(n6483), .B(n6474), .Z(n6482) );
  XOR U9224 ( .A(n6469), .B(n6473), .Z(n6484) );
  XOR U9225 ( .A(n6464), .B(n6468), .Z(n6485) );
  XOR U9226 ( .A(n6459), .B(n6463), .Z(n6486) );
  XOR U9227 ( .A(n6454), .B(n6458), .Z(n6487) );
  XOR U9228 ( .A(n6449), .B(n6453), .Z(n6488) );
  XOR U9229 ( .A(n6444), .B(n6448), .Z(n6489) );
  XOR U9230 ( .A(n6439), .B(n6443), .Z(n6490) );
  XOR U9231 ( .A(n6434), .B(n6438), .Z(n6491) );
  XOR U9232 ( .A(n6429), .B(n6433), .Z(n6492) );
  XOR U9233 ( .A(n6424), .B(n6428), .Z(n6493) );
  XOR U9234 ( .A(n6419), .B(n6423), .Z(n6494) );
  XOR U9235 ( .A(n6414), .B(n6418), .Z(n6495) );
  XOR U9236 ( .A(n6409), .B(n6413), .Z(n6496) );
  XOR U9237 ( .A(n6404), .B(n6408), .Z(n6497) );
  XOR U9238 ( .A(n6399), .B(n6403), .Z(n6498) );
  XOR U9239 ( .A(n6394), .B(n6398), .Z(n6499) );
  XOR U9240 ( .A(n6389), .B(n6393), .Z(n6500) );
  XOR U9241 ( .A(n6384), .B(n6388), .Z(n6501) );
  XOR U9242 ( .A(n6379), .B(n6383), .Z(n6502) );
  XOR U9243 ( .A(n6374), .B(n6378), .Z(n6503) );
  XOR U9244 ( .A(n6369), .B(n6373), .Z(n6504) );
  XOR U9245 ( .A(n6364), .B(n6368), .Z(n6505) );
  XOR U9246 ( .A(n6354), .B(n6363), .Z(n6506) );
  XOR U9247 ( .A(n6507), .B(n6353), .Z(n6354) );
  AND U9248 ( .A(b[25]), .B(a[68]), .Z(n6507) );
  XNOR U9249 ( .A(n6353), .B(n6359), .Z(n6508) );
  XNOR U9250 ( .A(n6358), .B(n6350), .Z(n6509) );
  XOR U9251 ( .A(n6349), .B(n6346), .Z(n6510) );
  XOR U9252 ( .A(n6511), .B(n6512), .Z(n6346) );
  XOR U9253 ( .A(n6344), .B(n6513), .Z(n6512) );
  XOR U9254 ( .A(n6514), .B(n6515), .Z(n6513) );
  XOR U9255 ( .A(n6516), .B(n6517), .Z(n6515) );
  NAND U9256 ( .A(a[63]), .B(b[30]), .Z(n6517) );
  AND U9257 ( .A(a[62]), .B(b[31]), .Z(n6516) );
  XOR U9258 ( .A(n6518), .B(n6514), .Z(n6511) );
  XOR U9259 ( .A(n6519), .B(n6520), .Z(n6514) );
  ANDN U9260 ( .B(n6521), .A(n6522), .Z(n6519) );
  AND U9261 ( .A(a[64]), .B(b[29]), .Z(n6518) );
  XOR U9262 ( .A(n6523), .B(n6344), .Z(n6345) );
  XOR U9263 ( .A(n6524), .B(n6525), .Z(n6344) );
  AND U9264 ( .A(n6526), .B(n6527), .Z(n6524) );
  AND U9265 ( .A(a[65]), .B(b[28]), .Z(n6523) );
  XOR U9266 ( .A(n6528), .B(n6349), .Z(n6351) );
  XOR U9267 ( .A(n6529), .B(n6530), .Z(n6349) );
  AND U9268 ( .A(n6531), .B(n6532), .Z(n6529) );
  AND U9269 ( .A(a[66]), .B(b[27]), .Z(n6528) );
  XOR U9270 ( .A(n6533), .B(n6534), .Z(n6353) );
  AND U9271 ( .A(n6535), .B(n6536), .Z(n6533) );
  XOR U9272 ( .A(n6537), .B(n6358), .Z(n6360) );
  XOR U9273 ( .A(n6538), .B(n6539), .Z(n6358) );
  AND U9274 ( .A(n6540), .B(n6541), .Z(n6538) );
  AND U9275 ( .A(a[67]), .B(b[26]), .Z(n6537) );
  XOR U9276 ( .A(n6543), .B(n6544), .Z(n6363) );
  AND U9277 ( .A(n6545), .B(n6546), .Z(n6543) );
  AND U9278 ( .A(a[69]), .B(b[24]), .Z(n6542) );
  XOR U9279 ( .A(n6548), .B(n6549), .Z(n6368) );
  AND U9280 ( .A(n6550), .B(n6551), .Z(n6548) );
  AND U9281 ( .A(a[70]), .B(b[23]), .Z(n6547) );
  XOR U9282 ( .A(n6553), .B(n6554), .Z(n6373) );
  AND U9283 ( .A(n6555), .B(n6556), .Z(n6553) );
  AND U9284 ( .A(a[71]), .B(b[22]), .Z(n6552) );
  XOR U9285 ( .A(n6558), .B(n6559), .Z(n6378) );
  AND U9286 ( .A(n6560), .B(n6561), .Z(n6558) );
  AND U9287 ( .A(a[72]), .B(b[21]), .Z(n6557) );
  XOR U9288 ( .A(n6563), .B(n6564), .Z(n6383) );
  AND U9289 ( .A(n6565), .B(n6566), .Z(n6563) );
  AND U9290 ( .A(a[73]), .B(b[20]), .Z(n6562) );
  XOR U9291 ( .A(n6568), .B(n6569), .Z(n6388) );
  AND U9292 ( .A(n6570), .B(n6571), .Z(n6568) );
  AND U9293 ( .A(a[74]), .B(b[19]), .Z(n6567) );
  XOR U9294 ( .A(n6573), .B(n6574), .Z(n6393) );
  AND U9295 ( .A(n6575), .B(n6576), .Z(n6573) );
  AND U9296 ( .A(a[75]), .B(b[18]), .Z(n6572) );
  XOR U9297 ( .A(n6578), .B(n6579), .Z(n6398) );
  AND U9298 ( .A(n6580), .B(n6581), .Z(n6578) );
  AND U9299 ( .A(a[76]), .B(b[17]), .Z(n6577) );
  XOR U9300 ( .A(n6583), .B(n6584), .Z(n6403) );
  AND U9301 ( .A(n6585), .B(n6586), .Z(n6583) );
  AND U9302 ( .A(a[77]), .B(b[16]), .Z(n6582) );
  XOR U9303 ( .A(n6588), .B(n6589), .Z(n6408) );
  AND U9304 ( .A(n6590), .B(n6591), .Z(n6588) );
  AND U9305 ( .A(a[78]), .B(b[15]), .Z(n6587) );
  XOR U9306 ( .A(n6593), .B(n6594), .Z(n6413) );
  AND U9307 ( .A(n6595), .B(n6596), .Z(n6593) );
  AND U9308 ( .A(a[79]), .B(b[14]), .Z(n6592) );
  XOR U9309 ( .A(n6598), .B(n6599), .Z(n6418) );
  AND U9310 ( .A(n6600), .B(n6601), .Z(n6598) );
  AND U9311 ( .A(a[80]), .B(b[13]), .Z(n6597) );
  XOR U9312 ( .A(n6603), .B(n6604), .Z(n6423) );
  AND U9313 ( .A(n6605), .B(n6606), .Z(n6603) );
  AND U9314 ( .A(a[81]), .B(b[12]), .Z(n6602) );
  XOR U9315 ( .A(n6608), .B(n6609), .Z(n6428) );
  AND U9316 ( .A(n6610), .B(n6611), .Z(n6608) );
  AND U9317 ( .A(a[82]), .B(b[11]), .Z(n6607) );
  XOR U9318 ( .A(n6613), .B(n6614), .Z(n6433) );
  AND U9319 ( .A(n6615), .B(n6616), .Z(n6613) );
  AND U9320 ( .A(a[83]), .B(b[10]), .Z(n6612) );
  XOR U9321 ( .A(n6618), .B(n6619), .Z(n6438) );
  AND U9322 ( .A(n6620), .B(n6621), .Z(n6618) );
  AND U9323 ( .A(a[84]), .B(b[9]), .Z(n6617) );
  XOR U9324 ( .A(n6623), .B(n6624), .Z(n6443) );
  AND U9325 ( .A(n6625), .B(n6626), .Z(n6623) );
  AND U9326 ( .A(a[85]), .B(b[8]), .Z(n6622) );
  XOR U9327 ( .A(n6628), .B(n6629), .Z(n6448) );
  AND U9328 ( .A(n6630), .B(n6631), .Z(n6628) );
  AND U9329 ( .A(a[86]), .B(b[7]), .Z(n6627) );
  XOR U9330 ( .A(n6633), .B(n6634), .Z(n6453) );
  AND U9331 ( .A(n6635), .B(n6636), .Z(n6633) );
  AND U9332 ( .A(a[87]), .B(b[6]), .Z(n6632) );
  XOR U9333 ( .A(n6638), .B(n6639), .Z(n6458) );
  AND U9334 ( .A(n6640), .B(n6641), .Z(n6638) );
  AND U9335 ( .A(a[88]), .B(b[5]), .Z(n6637) );
  XOR U9336 ( .A(n6643), .B(n6644), .Z(n6463) );
  AND U9337 ( .A(n6645), .B(n6646), .Z(n6643) );
  AND U9338 ( .A(a[89]), .B(b[4]), .Z(n6642) );
  XOR U9339 ( .A(n6648), .B(n6649), .Z(n6468) );
  AND U9340 ( .A(n6650), .B(n6651), .Z(n6648) );
  AND U9341 ( .A(a[90]), .B(b[3]), .Z(n6647) );
  XOR U9342 ( .A(n6653), .B(n6654), .Z(n6473) );
  OR U9343 ( .A(n6655), .B(n6656), .Z(n6654) );
  AND U9344 ( .A(a[91]), .B(b[2]), .Z(n6652) );
  XNOR U9345 ( .A(n6483), .B(n6657), .Z(n6479) );
  NAND U9346 ( .A(a[92]), .B(b[1]), .Z(n6657) );
  IV U9347 ( .A(n6477), .Z(n6483) );
  ANDN U9348 ( .B(n5092), .A(n5094), .Z(n6477) );
  NAND U9349 ( .A(a[92]), .B(b[0]), .Z(n5094) );
  XOR U9350 ( .A(n6655), .B(n6656), .Z(n5092) );
  XOR U9351 ( .A(n6659), .B(n6650), .Z(n6658) );
  XOR U9352 ( .A(n6645), .B(n6649), .Z(n6660) );
  XOR U9353 ( .A(n6640), .B(n6644), .Z(n6661) );
  XOR U9354 ( .A(n6635), .B(n6639), .Z(n6662) );
  XOR U9355 ( .A(n6630), .B(n6634), .Z(n6663) );
  XOR U9356 ( .A(n6625), .B(n6629), .Z(n6664) );
  XOR U9357 ( .A(n6620), .B(n6624), .Z(n6665) );
  XOR U9358 ( .A(n6615), .B(n6619), .Z(n6666) );
  XOR U9359 ( .A(n6610), .B(n6614), .Z(n6667) );
  XOR U9360 ( .A(n6605), .B(n6609), .Z(n6668) );
  XOR U9361 ( .A(n6600), .B(n6604), .Z(n6669) );
  XOR U9362 ( .A(n6595), .B(n6599), .Z(n6670) );
  XOR U9363 ( .A(n6590), .B(n6594), .Z(n6671) );
  XOR U9364 ( .A(n6585), .B(n6589), .Z(n6672) );
  XOR U9365 ( .A(n6580), .B(n6584), .Z(n6673) );
  XOR U9366 ( .A(n6575), .B(n6579), .Z(n6674) );
  XOR U9367 ( .A(n6570), .B(n6574), .Z(n6675) );
  XOR U9368 ( .A(n6565), .B(n6569), .Z(n6676) );
  XOR U9369 ( .A(n6560), .B(n6564), .Z(n6677) );
  XOR U9370 ( .A(n6555), .B(n6559), .Z(n6678) );
  XOR U9371 ( .A(n6550), .B(n6554), .Z(n6679) );
  XOR U9372 ( .A(n6545), .B(n6549), .Z(n6680) );
  XOR U9373 ( .A(n6535), .B(n6544), .Z(n6681) );
  XOR U9374 ( .A(n6682), .B(n6534), .Z(n6535) );
  AND U9375 ( .A(b[24]), .B(a[68]), .Z(n6682) );
  XNOR U9376 ( .A(n6534), .B(n6540), .Z(n6683) );
  XNOR U9377 ( .A(n6539), .B(n6531), .Z(n6684) );
  XNOR U9378 ( .A(n6530), .B(n6526), .Z(n6685) );
  XOR U9379 ( .A(n6525), .B(n6522), .Z(n6686) );
  XOR U9380 ( .A(n6687), .B(n6688), .Z(n6522) );
  XOR U9381 ( .A(n6520), .B(n6689), .Z(n6688) );
  XOR U9382 ( .A(n6690), .B(n6691), .Z(n6689) );
  XOR U9383 ( .A(n6692), .B(n6693), .Z(n6691) );
  NAND U9384 ( .A(a[62]), .B(b[30]), .Z(n6693) );
  AND U9385 ( .A(a[61]), .B(b[31]), .Z(n6692) );
  XOR U9386 ( .A(n6694), .B(n6690), .Z(n6687) );
  XOR U9387 ( .A(n6695), .B(n6696), .Z(n6690) );
  ANDN U9388 ( .B(n6697), .A(n6698), .Z(n6695) );
  AND U9389 ( .A(a[63]), .B(b[29]), .Z(n6694) );
  XOR U9390 ( .A(n6699), .B(n6520), .Z(n6521) );
  XOR U9391 ( .A(n6700), .B(n6701), .Z(n6520) );
  AND U9392 ( .A(n6702), .B(n6703), .Z(n6700) );
  AND U9393 ( .A(a[64]), .B(b[28]), .Z(n6699) );
  XOR U9394 ( .A(n6704), .B(n6525), .Z(n6527) );
  XOR U9395 ( .A(n6705), .B(n6706), .Z(n6525) );
  AND U9396 ( .A(n6707), .B(n6708), .Z(n6705) );
  AND U9397 ( .A(a[65]), .B(b[27]), .Z(n6704) );
  XOR U9398 ( .A(n6709), .B(n6530), .Z(n6532) );
  XOR U9399 ( .A(n6710), .B(n6711), .Z(n6530) );
  AND U9400 ( .A(n6712), .B(n6713), .Z(n6710) );
  AND U9401 ( .A(a[66]), .B(b[26]), .Z(n6709) );
  XOR U9402 ( .A(n6714), .B(n6715), .Z(n6534) );
  AND U9403 ( .A(n6716), .B(n6717), .Z(n6714) );
  XOR U9404 ( .A(n6718), .B(n6539), .Z(n6541) );
  XOR U9405 ( .A(n6719), .B(n6720), .Z(n6539) );
  AND U9406 ( .A(n6721), .B(n6722), .Z(n6719) );
  AND U9407 ( .A(a[67]), .B(b[25]), .Z(n6718) );
  XOR U9408 ( .A(n6724), .B(n6725), .Z(n6544) );
  AND U9409 ( .A(n6726), .B(n6727), .Z(n6724) );
  AND U9410 ( .A(a[69]), .B(b[23]), .Z(n6723) );
  XOR U9411 ( .A(n6729), .B(n6730), .Z(n6549) );
  AND U9412 ( .A(n6731), .B(n6732), .Z(n6729) );
  AND U9413 ( .A(a[70]), .B(b[22]), .Z(n6728) );
  XOR U9414 ( .A(n6734), .B(n6735), .Z(n6554) );
  AND U9415 ( .A(n6736), .B(n6737), .Z(n6734) );
  AND U9416 ( .A(a[71]), .B(b[21]), .Z(n6733) );
  XOR U9417 ( .A(n6739), .B(n6740), .Z(n6559) );
  AND U9418 ( .A(n6741), .B(n6742), .Z(n6739) );
  AND U9419 ( .A(a[72]), .B(b[20]), .Z(n6738) );
  XOR U9420 ( .A(n6744), .B(n6745), .Z(n6564) );
  AND U9421 ( .A(n6746), .B(n6747), .Z(n6744) );
  AND U9422 ( .A(a[73]), .B(b[19]), .Z(n6743) );
  XOR U9423 ( .A(n6749), .B(n6750), .Z(n6569) );
  AND U9424 ( .A(n6751), .B(n6752), .Z(n6749) );
  AND U9425 ( .A(a[74]), .B(b[18]), .Z(n6748) );
  XOR U9426 ( .A(n6754), .B(n6755), .Z(n6574) );
  AND U9427 ( .A(n6756), .B(n6757), .Z(n6754) );
  AND U9428 ( .A(a[75]), .B(b[17]), .Z(n6753) );
  XOR U9429 ( .A(n6759), .B(n6760), .Z(n6579) );
  AND U9430 ( .A(n6761), .B(n6762), .Z(n6759) );
  AND U9431 ( .A(a[76]), .B(b[16]), .Z(n6758) );
  XOR U9432 ( .A(n6764), .B(n6765), .Z(n6584) );
  AND U9433 ( .A(n6766), .B(n6767), .Z(n6764) );
  AND U9434 ( .A(a[77]), .B(b[15]), .Z(n6763) );
  XOR U9435 ( .A(n6769), .B(n6770), .Z(n6589) );
  AND U9436 ( .A(n6771), .B(n6772), .Z(n6769) );
  AND U9437 ( .A(a[78]), .B(b[14]), .Z(n6768) );
  XOR U9438 ( .A(n6774), .B(n6775), .Z(n6594) );
  AND U9439 ( .A(n6776), .B(n6777), .Z(n6774) );
  AND U9440 ( .A(a[79]), .B(b[13]), .Z(n6773) );
  XOR U9441 ( .A(n6779), .B(n6780), .Z(n6599) );
  AND U9442 ( .A(n6781), .B(n6782), .Z(n6779) );
  AND U9443 ( .A(a[80]), .B(b[12]), .Z(n6778) );
  XOR U9444 ( .A(n6784), .B(n6785), .Z(n6604) );
  AND U9445 ( .A(n6786), .B(n6787), .Z(n6784) );
  AND U9446 ( .A(a[81]), .B(b[11]), .Z(n6783) );
  XOR U9447 ( .A(n6789), .B(n6790), .Z(n6609) );
  AND U9448 ( .A(n6791), .B(n6792), .Z(n6789) );
  AND U9449 ( .A(a[82]), .B(b[10]), .Z(n6788) );
  XOR U9450 ( .A(n6794), .B(n6795), .Z(n6614) );
  AND U9451 ( .A(n6796), .B(n6797), .Z(n6794) );
  AND U9452 ( .A(a[83]), .B(b[9]), .Z(n6793) );
  XOR U9453 ( .A(n6799), .B(n6800), .Z(n6619) );
  AND U9454 ( .A(n6801), .B(n6802), .Z(n6799) );
  AND U9455 ( .A(a[84]), .B(b[8]), .Z(n6798) );
  XOR U9456 ( .A(n6804), .B(n6805), .Z(n6624) );
  AND U9457 ( .A(n6806), .B(n6807), .Z(n6804) );
  AND U9458 ( .A(a[85]), .B(b[7]), .Z(n6803) );
  XOR U9459 ( .A(n6809), .B(n6810), .Z(n6629) );
  AND U9460 ( .A(n6811), .B(n6812), .Z(n6809) );
  AND U9461 ( .A(a[86]), .B(b[6]), .Z(n6808) );
  XOR U9462 ( .A(n6814), .B(n6815), .Z(n6634) );
  AND U9463 ( .A(n6816), .B(n6817), .Z(n6814) );
  AND U9464 ( .A(a[87]), .B(b[5]), .Z(n6813) );
  XOR U9465 ( .A(n6819), .B(n6820), .Z(n6639) );
  AND U9466 ( .A(n6821), .B(n6822), .Z(n6819) );
  AND U9467 ( .A(a[88]), .B(b[4]), .Z(n6818) );
  XOR U9468 ( .A(n6824), .B(n6825), .Z(n6644) );
  AND U9469 ( .A(n6826), .B(n6827), .Z(n6824) );
  AND U9470 ( .A(a[89]), .B(b[3]), .Z(n6823) );
  XOR U9471 ( .A(n6829), .B(n6830), .Z(n6649) );
  OR U9472 ( .A(n6831), .B(n6832), .Z(n6830) );
  AND U9473 ( .A(a[90]), .B(b[2]), .Z(n6828) );
  XNOR U9474 ( .A(n6659), .B(n6833), .Z(n6655) );
  NAND U9475 ( .A(a[91]), .B(b[1]), .Z(n6833) );
  IV U9476 ( .A(n6653), .Z(n6659) );
  ANDN U9477 ( .B(n5097), .A(n5099), .Z(n6653) );
  NAND U9478 ( .A(a[91]), .B(b[0]), .Z(n5099) );
  XOR U9479 ( .A(n6831), .B(n6832), .Z(n5097) );
  XOR U9480 ( .A(n6835), .B(n6826), .Z(n6834) );
  XOR U9481 ( .A(n6821), .B(n6825), .Z(n6836) );
  XOR U9482 ( .A(n6816), .B(n6820), .Z(n6837) );
  XOR U9483 ( .A(n6811), .B(n6815), .Z(n6838) );
  XOR U9484 ( .A(n6806), .B(n6810), .Z(n6839) );
  XOR U9485 ( .A(n6801), .B(n6805), .Z(n6840) );
  XOR U9486 ( .A(n6796), .B(n6800), .Z(n6841) );
  XOR U9487 ( .A(n6791), .B(n6795), .Z(n6842) );
  XOR U9488 ( .A(n6786), .B(n6790), .Z(n6843) );
  XOR U9489 ( .A(n6781), .B(n6785), .Z(n6844) );
  XOR U9490 ( .A(n6776), .B(n6780), .Z(n6845) );
  XOR U9491 ( .A(n6771), .B(n6775), .Z(n6846) );
  XOR U9492 ( .A(n6766), .B(n6770), .Z(n6847) );
  XOR U9493 ( .A(n6761), .B(n6765), .Z(n6848) );
  XOR U9494 ( .A(n6756), .B(n6760), .Z(n6849) );
  XOR U9495 ( .A(n6751), .B(n6755), .Z(n6850) );
  XOR U9496 ( .A(n6746), .B(n6750), .Z(n6851) );
  XOR U9497 ( .A(n6741), .B(n6745), .Z(n6852) );
  XOR U9498 ( .A(n6736), .B(n6740), .Z(n6853) );
  XOR U9499 ( .A(n6731), .B(n6735), .Z(n6854) );
  XOR U9500 ( .A(n6726), .B(n6730), .Z(n6855) );
  XOR U9501 ( .A(n6716), .B(n6725), .Z(n6856) );
  XOR U9502 ( .A(n6857), .B(n6715), .Z(n6716) );
  AND U9503 ( .A(b[23]), .B(a[68]), .Z(n6857) );
  XNOR U9504 ( .A(n6715), .B(n6721), .Z(n6858) );
  XNOR U9505 ( .A(n6720), .B(n6712), .Z(n6859) );
  XNOR U9506 ( .A(n6711), .B(n6707), .Z(n6860) );
  XNOR U9507 ( .A(n6706), .B(n6702), .Z(n6861) );
  XOR U9508 ( .A(n6701), .B(n6698), .Z(n6862) );
  XOR U9509 ( .A(n6863), .B(n6864), .Z(n6698) );
  XOR U9510 ( .A(n6696), .B(n6865), .Z(n6864) );
  XOR U9511 ( .A(n6866), .B(n6867), .Z(n6865) );
  XOR U9512 ( .A(n6868), .B(n6869), .Z(n6867) );
  NAND U9513 ( .A(a[61]), .B(b[30]), .Z(n6869) );
  AND U9514 ( .A(a[60]), .B(b[31]), .Z(n6868) );
  XOR U9515 ( .A(n6870), .B(n6866), .Z(n6863) );
  XOR U9516 ( .A(n6871), .B(n6872), .Z(n6866) );
  ANDN U9517 ( .B(n6873), .A(n6874), .Z(n6871) );
  AND U9518 ( .A(a[62]), .B(b[29]), .Z(n6870) );
  XOR U9519 ( .A(n6875), .B(n6696), .Z(n6697) );
  XOR U9520 ( .A(n6876), .B(n6877), .Z(n6696) );
  AND U9521 ( .A(n6878), .B(n6879), .Z(n6876) );
  AND U9522 ( .A(a[63]), .B(b[28]), .Z(n6875) );
  XOR U9523 ( .A(n6880), .B(n6701), .Z(n6703) );
  XOR U9524 ( .A(n6881), .B(n6882), .Z(n6701) );
  AND U9525 ( .A(n6883), .B(n6884), .Z(n6881) );
  AND U9526 ( .A(a[64]), .B(b[27]), .Z(n6880) );
  XOR U9527 ( .A(n6885), .B(n6706), .Z(n6708) );
  XOR U9528 ( .A(n6886), .B(n6887), .Z(n6706) );
  AND U9529 ( .A(n6888), .B(n6889), .Z(n6886) );
  AND U9530 ( .A(a[65]), .B(b[26]), .Z(n6885) );
  XOR U9531 ( .A(n6890), .B(n6711), .Z(n6713) );
  XOR U9532 ( .A(n6891), .B(n6892), .Z(n6711) );
  AND U9533 ( .A(n6893), .B(n6894), .Z(n6891) );
  AND U9534 ( .A(a[66]), .B(b[25]), .Z(n6890) );
  XOR U9535 ( .A(n6895), .B(n6896), .Z(n6715) );
  AND U9536 ( .A(n6897), .B(n6898), .Z(n6895) );
  XOR U9537 ( .A(n6899), .B(n6720), .Z(n6722) );
  XOR U9538 ( .A(n6900), .B(n6901), .Z(n6720) );
  AND U9539 ( .A(n6902), .B(n6903), .Z(n6900) );
  AND U9540 ( .A(a[67]), .B(b[24]), .Z(n6899) );
  XOR U9541 ( .A(n6905), .B(n6906), .Z(n6725) );
  AND U9542 ( .A(n6907), .B(n6908), .Z(n6905) );
  AND U9543 ( .A(a[69]), .B(b[22]), .Z(n6904) );
  XOR U9544 ( .A(n6910), .B(n6911), .Z(n6730) );
  AND U9545 ( .A(n6912), .B(n6913), .Z(n6910) );
  AND U9546 ( .A(a[70]), .B(b[21]), .Z(n6909) );
  XOR U9547 ( .A(n6915), .B(n6916), .Z(n6735) );
  AND U9548 ( .A(n6917), .B(n6918), .Z(n6915) );
  AND U9549 ( .A(a[71]), .B(b[20]), .Z(n6914) );
  XOR U9550 ( .A(n6920), .B(n6921), .Z(n6740) );
  AND U9551 ( .A(n6922), .B(n6923), .Z(n6920) );
  AND U9552 ( .A(a[72]), .B(b[19]), .Z(n6919) );
  XOR U9553 ( .A(n6925), .B(n6926), .Z(n6745) );
  AND U9554 ( .A(n6927), .B(n6928), .Z(n6925) );
  AND U9555 ( .A(a[73]), .B(b[18]), .Z(n6924) );
  XOR U9556 ( .A(n6930), .B(n6931), .Z(n6750) );
  AND U9557 ( .A(n6932), .B(n6933), .Z(n6930) );
  AND U9558 ( .A(a[74]), .B(b[17]), .Z(n6929) );
  XOR U9559 ( .A(n6935), .B(n6936), .Z(n6755) );
  AND U9560 ( .A(n6937), .B(n6938), .Z(n6935) );
  AND U9561 ( .A(a[75]), .B(b[16]), .Z(n6934) );
  XOR U9562 ( .A(n6940), .B(n6941), .Z(n6760) );
  AND U9563 ( .A(n6942), .B(n6943), .Z(n6940) );
  AND U9564 ( .A(a[76]), .B(b[15]), .Z(n6939) );
  XOR U9565 ( .A(n6945), .B(n6946), .Z(n6765) );
  AND U9566 ( .A(n6947), .B(n6948), .Z(n6945) );
  AND U9567 ( .A(a[77]), .B(b[14]), .Z(n6944) );
  XOR U9568 ( .A(n6950), .B(n6951), .Z(n6770) );
  AND U9569 ( .A(n6952), .B(n6953), .Z(n6950) );
  AND U9570 ( .A(a[78]), .B(b[13]), .Z(n6949) );
  XOR U9571 ( .A(n6955), .B(n6956), .Z(n6775) );
  AND U9572 ( .A(n6957), .B(n6958), .Z(n6955) );
  AND U9573 ( .A(a[79]), .B(b[12]), .Z(n6954) );
  XOR U9574 ( .A(n6960), .B(n6961), .Z(n6780) );
  AND U9575 ( .A(n6962), .B(n6963), .Z(n6960) );
  AND U9576 ( .A(a[80]), .B(b[11]), .Z(n6959) );
  XOR U9577 ( .A(n6965), .B(n6966), .Z(n6785) );
  AND U9578 ( .A(n6967), .B(n6968), .Z(n6965) );
  AND U9579 ( .A(a[81]), .B(b[10]), .Z(n6964) );
  XOR U9580 ( .A(n6970), .B(n6971), .Z(n6790) );
  AND U9581 ( .A(n6972), .B(n6973), .Z(n6970) );
  AND U9582 ( .A(a[82]), .B(b[9]), .Z(n6969) );
  XOR U9583 ( .A(n6975), .B(n6976), .Z(n6795) );
  AND U9584 ( .A(n6977), .B(n6978), .Z(n6975) );
  AND U9585 ( .A(a[83]), .B(b[8]), .Z(n6974) );
  XOR U9586 ( .A(n6980), .B(n6981), .Z(n6800) );
  AND U9587 ( .A(n6982), .B(n6983), .Z(n6980) );
  AND U9588 ( .A(a[84]), .B(b[7]), .Z(n6979) );
  XOR U9589 ( .A(n6985), .B(n6986), .Z(n6805) );
  AND U9590 ( .A(n6987), .B(n6988), .Z(n6985) );
  AND U9591 ( .A(a[85]), .B(b[6]), .Z(n6984) );
  XOR U9592 ( .A(n6990), .B(n6991), .Z(n6810) );
  AND U9593 ( .A(n6992), .B(n6993), .Z(n6990) );
  AND U9594 ( .A(a[86]), .B(b[5]), .Z(n6989) );
  XOR U9595 ( .A(n6995), .B(n6996), .Z(n6815) );
  AND U9596 ( .A(n6997), .B(n6998), .Z(n6995) );
  AND U9597 ( .A(a[87]), .B(b[4]), .Z(n6994) );
  XOR U9598 ( .A(n7000), .B(n7001), .Z(n6820) );
  AND U9599 ( .A(n7002), .B(n7003), .Z(n7000) );
  AND U9600 ( .A(a[88]), .B(b[3]), .Z(n6999) );
  XOR U9601 ( .A(n7005), .B(n7006), .Z(n6825) );
  OR U9602 ( .A(n7007), .B(n7008), .Z(n7006) );
  AND U9603 ( .A(a[89]), .B(b[2]), .Z(n7004) );
  XNOR U9604 ( .A(n6835), .B(n7009), .Z(n6831) );
  NAND U9605 ( .A(a[90]), .B(b[1]), .Z(n7009) );
  IV U9606 ( .A(n6829), .Z(n6835) );
  ANDN U9607 ( .B(n5102), .A(n5104), .Z(n6829) );
  NAND U9608 ( .A(a[90]), .B(b[0]), .Z(n5104) );
  XOR U9609 ( .A(n7007), .B(n7008), .Z(n5102) );
  XOR U9610 ( .A(n7011), .B(n7002), .Z(n7010) );
  XOR U9611 ( .A(n6997), .B(n7001), .Z(n7012) );
  XOR U9612 ( .A(n6992), .B(n6996), .Z(n7013) );
  XOR U9613 ( .A(n6987), .B(n6991), .Z(n7014) );
  XOR U9614 ( .A(n6982), .B(n6986), .Z(n7015) );
  XOR U9615 ( .A(n6977), .B(n6981), .Z(n7016) );
  XOR U9616 ( .A(n6972), .B(n6976), .Z(n7017) );
  XOR U9617 ( .A(n6967), .B(n6971), .Z(n7018) );
  XOR U9618 ( .A(n6962), .B(n6966), .Z(n7019) );
  XOR U9619 ( .A(n6957), .B(n6961), .Z(n7020) );
  XOR U9620 ( .A(n6952), .B(n6956), .Z(n7021) );
  XOR U9621 ( .A(n6947), .B(n6951), .Z(n7022) );
  XOR U9622 ( .A(n6942), .B(n6946), .Z(n7023) );
  XOR U9623 ( .A(n6937), .B(n6941), .Z(n7024) );
  XOR U9624 ( .A(n6932), .B(n6936), .Z(n7025) );
  XOR U9625 ( .A(n6927), .B(n6931), .Z(n7026) );
  XOR U9626 ( .A(n6922), .B(n6926), .Z(n7027) );
  XOR U9627 ( .A(n6917), .B(n6921), .Z(n7028) );
  XOR U9628 ( .A(n6912), .B(n6916), .Z(n7029) );
  XOR U9629 ( .A(n6907), .B(n6911), .Z(n7030) );
  XOR U9630 ( .A(n6897), .B(n6906), .Z(n7031) );
  XOR U9631 ( .A(n7032), .B(n6896), .Z(n6897) );
  AND U9632 ( .A(b[22]), .B(a[68]), .Z(n7032) );
  XNOR U9633 ( .A(n6896), .B(n6902), .Z(n7033) );
  XNOR U9634 ( .A(n6901), .B(n6893), .Z(n7034) );
  XNOR U9635 ( .A(n6892), .B(n6888), .Z(n7035) );
  XNOR U9636 ( .A(n6887), .B(n6883), .Z(n7036) );
  XNOR U9637 ( .A(n6882), .B(n6878), .Z(n7037) );
  XOR U9638 ( .A(n6877), .B(n6874), .Z(n7038) );
  XOR U9639 ( .A(n7039), .B(n7040), .Z(n6874) );
  XOR U9640 ( .A(n6872), .B(n7041), .Z(n7040) );
  XOR U9641 ( .A(n7042), .B(n7043), .Z(n7041) );
  XOR U9642 ( .A(n7044), .B(n7045), .Z(n7043) );
  NAND U9643 ( .A(a[60]), .B(b[30]), .Z(n7045) );
  AND U9644 ( .A(a[59]), .B(b[31]), .Z(n7044) );
  XOR U9645 ( .A(n7046), .B(n7042), .Z(n7039) );
  XOR U9646 ( .A(n7047), .B(n7048), .Z(n7042) );
  ANDN U9647 ( .B(n7049), .A(n7050), .Z(n7047) );
  AND U9648 ( .A(a[61]), .B(b[29]), .Z(n7046) );
  XOR U9649 ( .A(n7051), .B(n6872), .Z(n6873) );
  XOR U9650 ( .A(n7052), .B(n7053), .Z(n6872) );
  AND U9651 ( .A(n7054), .B(n7055), .Z(n7052) );
  AND U9652 ( .A(a[62]), .B(b[28]), .Z(n7051) );
  XOR U9653 ( .A(n7056), .B(n6877), .Z(n6879) );
  XOR U9654 ( .A(n7057), .B(n7058), .Z(n6877) );
  AND U9655 ( .A(n7059), .B(n7060), .Z(n7057) );
  AND U9656 ( .A(a[63]), .B(b[27]), .Z(n7056) );
  XOR U9657 ( .A(n7061), .B(n6882), .Z(n6884) );
  XOR U9658 ( .A(n7062), .B(n7063), .Z(n6882) );
  AND U9659 ( .A(n7064), .B(n7065), .Z(n7062) );
  AND U9660 ( .A(a[64]), .B(b[26]), .Z(n7061) );
  XOR U9661 ( .A(n7066), .B(n6887), .Z(n6889) );
  XOR U9662 ( .A(n7067), .B(n7068), .Z(n6887) );
  AND U9663 ( .A(n7069), .B(n7070), .Z(n7067) );
  AND U9664 ( .A(a[65]), .B(b[25]), .Z(n7066) );
  XOR U9665 ( .A(n7071), .B(n6892), .Z(n6894) );
  XOR U9666 ( .A(n7072), .B(n7073), .Z(n6892) );
  AND U9667 ( .A(n7074), .B(n7075), .Z(n7072) );
  AND U9668 ( .A(a[66]), .B(b[24]), .Z(n7071) );
  XOR U9669 ( .A(n7076), .B(n7077), .Z(n6896) );
  AND U9670 ( .A(n7078), .B(n7079), .Z(n7076) );
  XOR U9671 ( .A(n7080), .B(n6901), .Z(n6903) );
  XOR U9672 ( .A(n7081), .B(n7082), .Z(n6901) );
  AND U9673 ( .A(n7083), .B(n7084), .Z(n7081) );
  AND U9674 ( .A(a[67]), .B(b[23]), .Z(n7080) );
  XOR U9675 ( .A(n7086), .B(n7087), .Z(n6906) );
  AND U9676 ( .A(n7088), .B(n7089), .Z(n7086) );
  AND U9677 ( .A(a[69]), .B(b[21]), .Z(n7085) );
  XOR U9678 ( .A(n7091), .B(n7092), .Z(n6911) );
  AND U9679 ( .A(n7093), .B(n7094), .Z(n7091) );
  AND U9680 ( .A(a[70]), .B(b[20]), .Z(n7090) );
  XOR U9681 ( .A(n7096), .B(n7097), .Z(n6916) );
  AND U9682 ( .A(n7098), .B(n7099), .Z(n7096) );
  AND U9683 ( .A(a[71]), .B(b[19]), .Z(n7095) );
  XOR U9684 ( .A(n7101), .B(n7102), .Z(n6921) );
  AND U9685 ( .A(n7103), .B(n7104), .Z(n7101) );
  AND U9686 ( .A(a[72]), .B(b[18]), .Z(n7100) );
  XOR U9687 ( .A(n7106), .B(n7107), .Z(n6926) );
  AND U9688 ( .A(n7108), .B(n7109), .Z(n7106) );
  AND U9689 ( .A(a[73]), .B(b[17]), .Z(n7105) );
  XOR U9690 ( .A(n7111), .B(n7112), .Z(n6931) );
  AND U9691 ( .A(n7113), .B(n7114), .Z(n7111) );
  AND U9692 ( .A(a[74]), .B(b[16]), .Z(n7110) );
  XOR U9693 ( .A(n7116), .B(n7117), .Z(n6936) );
  AND U9694 ( .A(n7118), .B(n7119), .Z(n7116) );
  AND U9695 ( .A(a[75]), .B(b[15]), .Z(n7115) );
  XOR U9696 ( .A(n7121), .B(n7122), .Z(n6941) );
  AND U9697 ( .A(n7123), .B(n7124), .Z(n7121) );
  AND U9698 ( .A(a[76]), .B(b[14]), .Z(n7120) );
  XOR U9699 ( .A(n7126), .B(n7127), .Z(n6946) );
  AND U9700 ( .A(n7128), .B(n7129), .Z(n7126) );
  AND U9701 ( .A(a[77]), .B(b[13]), .Z(n7125) );
  XOR U9702 ( .A(n7131), .B(n7132), .Z(n6951) );
  AND U9703 ( .A(n7133), .B(n7134), .Z(n7131) );
  AND U9704 ( .A(a[78]), .B(b[12]), .Z(n7130) );
  XOR U9705 ( .A(n7136), .B(n7137), .Z(n6956) );
  AND U9706 ( .A(n7138), .B(n7139), .Z(n7136) );
  AND U9707 ( .A(a[79]), .B(b[11]), .Z(n7135) );
  XOR U9708 ( .A(n7141), .B(n7142), .Z(n6961) );
  AND U9709 ( .A(n7143), .B(n7144), .Z(n7141) );
  AND U9710 ( .A(a[80]), .B(b[10]), .Z(n7140) );
  XOR U9711 ( .A(n7146), .B(n7147), .Z(n6966) );
  AND U9712 ( .A(n7148), .B(n7149), .Z(n7146) );
  AND U9713 ( .A(a[81]), .B(b[9]), .Z(n7145) );
  XOR U9714 ( .A(n7151), .B(n7152), .Z(n6971) );
  AND U9715 ( .A(n7153), .B(n7154), .Z(n7151) );
  AND U9716 ( .A(a[82]), .B(b[8]), .Z(n7150) );
  XOR U9717 ( .A(n7156), .B(n7157), .Z(n6976) );
  AND U9718 ( .A(n7158), .B(n7159), .Z(n7156) );
  AND U9719 ( .A(a[83]), .B(b[7]), .Z(n7155) );
  XOR U9720 ( .A(n7161), .B(n7162), .Z(n6981) );
  AND U9721 ( .A(n7163), .B(n7164), .Z(n7161) );
  AND U9722 ( .A(a[84]), .B(b[6]), .Z(n7160) );
  XOR U9723 ( .A(n7166), .B(n7167), .Z(n6986) );
  AND U9724 ( .A(n7168), .B(n7169), .Z(n7166) );
  AND U9725 ( .A(a[85]), .B(b[5]), .Z(n7165) );
  XOR U9726 ( .A(n7171), .B(n7172), .Z(n6991) );
  AND U9727 ( .A(n7173), .B(n7174), .Z(n7171) );
  AND U9728 ( .A(a[86]), .B(b[4]), .Z(n7170) );
  XOR U9729 ( .A(n7176), .B(n7177), .Z(n6996) );
  AND U9730 ( .A(n7178), .B(n7179), .Z(n7176) );
  AND U9731 ( .A(a[87]), .B(b[3]), .Z(n7175) );
  XOR U9732 ( .A(n7181), .B(n7182), .Z(n7001) );
  OR U9733 ( .A(n7183), .B(n7184), .Z(n7182) );
  AND U9734 ( .A(a[88]), .B(b[2]), .Z(n7180) );
  XNOR U9735 ( .A(n7011), .B(n7185), .Z(n7007) );
  NAND U9736 ( .A(a[89]), .B(b[1]), .Z(n7185) );
  IV U9737 ( .A(n7005), .Z(n7011) );
  ANDN U9738 ( .B(n5107), .A(n5109), .Z(n7005) );
  NAND U9739 ( .A(a[89]), .B(b[0]), .Z(n5109) );
  XOR U9740 ( .A(n7183), .B(n7184), .Z(n5107) );
  XOR U9741 ( .A(n7187), .B(n7178), .Z(n7186) );
  XOR U9742 ( .A(n7173), .B(n7177), .Z(n7188) );
  XOR U9743 ( .A(n7168), .B(n7172), .Z(n7189) );
  XOR U9744 ( .A(n7163), .B(n7167), .Z(n7190) );
  XOR U9745 ( .A(n7158), .B(n7162), .Z(n7191) );
  XOR U9746 ( .A(n7153), .B(n7157), .Z(n7192) );
  XOR U9747 ( .A(n7148), .B(n7152), .Z(n7193) );
  XOR U9748 ( .A(n7143), .B(n7147), .Z(n7194) );
  XOR U9749 ( .A(n7138), .B(n7142), .Z(n7195) );
  XOR U9750 ( .A(n7133), .B(n7137), .Z(n7196) );
  XOR U9751 ( .A(n7128), .B(n7132), .Z(n7197) );
  XOR U9752 ( .A(n7123), .B(n7127), .Z(n7198) );
  XOR U9753 ( .A(n7118), .B(n7122), .Z(n7199) );
  XOR U9754 ( .A(n7113), .B(n7117), .Z(n7200) );
  XOR U9755 ( .A(n7108), .B(n7112), .Z(n7201) );
  XOR U9756 ( .A(n7103), .B(n7107), .Z(n7202) );
  XOR U9757 ( .A(n7098), .B(n7102), .Z(n7203) );
  XOR U9758 ( .A(n7093), .B(n7097), .Z(n7204) );
  XOR U9759 ( .A(n7088), .B(n7092), .Z(n7205) );
  XOR U9760 ( .A(n7078), .B(n7087), .Z(n7206) );
  XOR U9761 ( .A(n7207), .B(n7077), .Z(n7078) );
  AND U9762 ( .A(b[21]), .B(a[68]), .Z(n7207) );
  XNOR U9763 ( .A(n7077), .B(n7083), .Z(n7208) );
  XNOR U9764 ( .A(n7082), .B(n7074), .Z(n7209) );
  XNOR U9765 ( .A(n7073), .B(n7069), .Z(n7210) );
  XNOR U9766 ( .A(n7068), .B(n7064), .Z(n7211) );
  XNOR U9767 ( .A(n7063), .B(n7059), .Z(n7212) );
  XNOR U9768 ( .A(n7058), .B(n7054), .Z(n7213) );
  XOR U9769 ( .A(n7053), .B(n7050), .Z(n7214) );
  XOR U9770 ( .A(n7215), .B(n7216), .Z(n7050) );
  XOR U9771 ( .A(n7048), .B(n7217), .Z(n7216) );
  XOR U9772 ( .A(n7218), .B(n7219), .Z(n7217) );
  XOR U9773 ( .A(n7220), .B(n7221), .Z(n7219) );
  NAND U9774 ( .A(a[59]), .B(b[30]), .Z(n7221) );
  AND U9775 ( .A(a[58]), .B(b[31]), .Z(n7220) );
  XOR U9776 ( .A(n7222), .B(n7218), .Z(n7215) );
  XOR U9777 ( .A(n7223), .B(n7224), .Z(n7218) );
  ANDN U9778 ( .B(n7225), .A(n7226), .Z(n7223) );
  AND U9779 ( .A(a[60]), .B(b[29]), .Z(n7222) );
  XOR U9780 ( .A(n7227), .B(n7048), .Z(n7049) );
  XOR U9781 ( .A(n7228), .B(n7229), .Z(n7048) );
  AND U9782 ( .A(n7230), .B(n7231), .Z(n7228) );
  AND U9783 ( .A(a[61]), .B(b[28]), .Z(n7227) );
  XOR U9784 ( .A(n7232), .B(n7053), .Z(n7055) );
  XOR U9785 ( .A(n7233), .B(n7234), .Z(n7053) );
  AND U9786 ( .A(n7235), .B(n7236), .Z(n7233) );
  AND U9787 ( .A(a[62]), .B(b[27]), .Z(n7232) );
  XOR U9788 ( .A(n7237), .B(n7058), .Z(n7060) );
  XOR U9789 ( .A(n7238), .B(n7239), .Z(n7058) );
  AND U9790 ( .A(n7240), .B(n7241), .Z(n7238) );
  AND U9791 ( .A(a[63]), .B(b[26]), .Z(n7237) );
  XOR U9792 ( .A(n7242), .B(n7063), .Z(n7065) );
  XOR U9793 ( .A(n7243), .B(n7244), .Z(n7063) );
  AND U9794 ( .A(n7245), .B(n7246), .Z(n7243) );
  AND U9795 ( .A(a[64]), .B(b[25]), .Z(n7242) );
  XOR U9796 ( .A(n7247), .B(n7068), .Z(n7070) );
  XOR U9797 ( .A(n7248), .B(n7249), .Z(n7068) );
  AND U9798 ( .A(n7250), .B(n7251), .Z(n7248) );
  AND U9799 ( .A(a[65]), .B(b[24]), .Z(n7247) );
  XOR U9800 ( .A(n7252), .B(n7073), .Z(n7075) );
  XOR U9801 ( .A(n7253), .B(n7254), .Z(n7073) );
  AND U9802 ( .A(n7255), .B(n7256), .Z(n7253) );
  AND U9803 ( .A(a[66]), .B(b[23]), .Z(n7252) );
  XOR U9804 ( .A(n7257), .B(n7258), .Z(n7077) );
  AND U9805 ( .A(n7259), .B(n7260), .Z(n7257) );
  XOR U9806 ( .A(n7261), .B(n7082), .Z(n7084) );
  XOR U9807 ( .A(n7262), .B(n7263), .Z(n7082) );
  AND U9808 ( .A(n7264), .B(n7265), .Z(n7262) );
  AND U9809 ( .A(a[67]), .B(b[22]), .Z(n7261) );
  XOR U9810 ( .A(n7267), .B(n7268), .Z(n7087) );
  AND U9811 ( .A(n7269), .B(n7270), .Z(n7267) );
  AND U9812 ( .A(a[69]), .B(b[20]), .Z(n7266) );
  XOR U9813 ( .A(n7272), .B(n7273), .Z(n7092) );
  AND U9814 ( .A(n7274), .B(n7275), .Z(n7272) );
  AND U9815 ( .A(a[70]), .B(b[19]), .Z(n7271) );
  XOR U9816 ( .A(n7277), .B(n7278), .Z(n7097) );
  AND U9817 ( .A(n7279), .B(n7280), .Z(n7277) );
  AND U9818 ( .A(a[71]), .B(b[18]), .Z(n7276) );
  XOR U9819 ( .A(n7282), .B(n7283), .Z(n7102) );
  AND U9820 ( .A(n7284), .B(n7285), .Z(n7282) );
  AND U9821 ( .A(a[72]), .B(b[17]), .Z(n7281) );
  XOR U9822 ( .A(n7287), .B(n7288), .Z(n7107) );
  AND U9823 ( .A(n7289), .B(n7290), .Z(n7287) );
  AND U9824 ( .A(a[73]), .B(b[16]), .Z(n7286) );
  XOR U9825 ( .A(n7292), .B(n7293), .Z(n7112) );
  AND U9826 ( .A(n7294), .B(n7295), .Z(n7292) );
  AND U9827 ( .A(a[74]), .B(b[15]), .Z(n7291) );
  XOR U9828 ( .A(n7297), .B(n7298), .Z(n7117) );
  AND U9829 ( .A(n7299), .B(n7300), .Z(n7297) );
  AND U9830 ( .A(a[75]), .B(b[14]), .Z(n7296) );
  XOR U9831 ( .A(n7302), .B(n7303), .Z(n7122) );
  AND U9832 ( .A(n7304), .B(n7305), .Z(n7302) );
  AND U9833 ( .A(a[76]), .B(b[13]), .Z(n7301) );
  XOR U9834 ( .A(n7307), .B(n7308), .Z(n7127) );
  AND U9835 ( .A(n7309), .B(n7310), .Z(n7307) );
  AND U9836 ( .A(a[77]), .B(b[12]), .Z(n7306) );
  XOR U9837 ( .A(n7312), .B(n7313), .Z(n7132) );
  AND U9838 ( .A(n7314), .B(n7315), .Z(n7312) );
  AND U9839 ( .A(a[78]), .B(b[11]), .Z(n7311) );
  XOR U9840 ( .A(n7317), .B(n7318), .Z(n7137) );
  AND U9841 ( .A(n7319), .B(n7320), .Z(n7317) );
  AND U9842 ( .A(a[79]), .B(b[10]), .Z(n7316) );
  XOR U9843 ( .A(n7322), .B(n7323), .Z(n7142) );
  AND U9844 ( .A(n7324), .B(n7325), .Z(n7322) );
  AND U9845 ( .A(a[80]), .B(b[9]), .Z(n7321) );
  XOR U9846 ( .A(n7327), .B(n7328), .Z(n7147) );
  AND U9847 ( .A(n7329), .B(n7330), .Z(n7327) );
  AND U9848 ( .A(a[81]), .B(b[8]), .Z(n7326) );
  XOR U9849 ( .A(n7332), .B(n7333), .Z(n7152) );
  AND U9850 ( .A(n7334), .B(n7335), .Z(n7332) );
  AND U9851 ( .A(a[82]), .B(b[7]), .Z(n7331) );
  XOR U9852 ( .A(n7337), .B(n7338), .Z(n7157) );
  AND U9853 ( .A(n7339), .B(n7340), .Z(n7337) );
  AND U9854 ( .A(a[83]), .B(b[6]), .Z(n7336) );
  XOR U9855 ( .A(n7342), .B(n7343), .Z(n7162) );
  AND U9856 ( .A(n7344), .B(n7345), .Z(n7342) );
  AND U9857 ( .A(a[84]), .B(b[5]), .Z(n7341) );
  XOR U9858 ( .A(n7347), .B(n7348), .Z(n7167) );
  AND U9859 ( .A(n7349), .B(n7350), .Z(n7347) );
  AND U9860 ( .A(a[85]), .B(b[4]), .Z(n7346) );
  XOR U9861 ( .A(n7352), .B(n7353), .Z(n7172) );
  AND U9862 ( .A(n7354), .B(n7355), .Z(n7352) );
  AND U9863 ( .A(a[86]), .B(b[3]), .Z(n7351) );
  XOR U9864 ( .A(n7357), .B(n7358), .Z(n7177) );
  OR U9865 ( .A(n7359), .B(n7360), .Z(n7358) );
  AND U9866 ( .A(a[87]), .B(b[2]), .Z(n7356) );
  XNOR U9867 ( .A(n7187), .B(n7361), .Z(n7183) );
  NAND U9868 ( .A(a[88]), .B(b[1]), .Z(n7361) );
  IV U9869 ( .A(n7181), .Z(n7187) );
  ANDN U9870 ( .B(n5112), .A(n5114), .Z(n7181) );
  NAND U9871 ( .A(a[88]), .B(b[0]), .Z(n5114) );
  XOR U9872 ( .A(n7359), .B(n7360), .Z(n5112) );
  XOR U9873 ( .A(n7363), .B(n7354), .Z(n7362) );
  XOR U9874 ( .A(n7349), .B(n7353), .Z(n7364) );
  XOR U9875 ( .A(n7344), .B(n7348), .Z(n7365) );
  XOR U9876 ( .A(n7339), .B(n7343), .Z(n7366) );
  XOR U9877 ( .A(n7334), .B(n7338), .Z(n7367) );
  XOR U9878 ( .A(n7329), .B(n7333), .Z(n7368) );
  XOR U9879 ( .A(n7324), .B(n7328), .Z(n7369) );
  XOR U9880 ( .A(n7319), .B(n7323), .Z(n7370) );
  XOR U9881 ( .A(n7314), .B(n7318), .Z(n7371) );
  XOR U9882 ( .A(n7309), .B(n7313), .Z(n7372) );
  XOR U9883 ( .A(n7304), .B(n7308), .Z(n7373) );
  XOR U9884 ( .A(n7299), .B(n7303), .Z(n7374) );
  XOR U9885 ( .A(n7294), .B(n7298), .Z(n7375) );
  XOR U9886 ( .A(n7289), .B(n7293), .Z(n7376) );
  XOR U9887 ( .A(n7284), .B(n7288), .Z(n7377) );
  XOR U9888 ( .A(n7279), .B(n7283), .Z(n7378) );
  XOR U9889 ( .A(n7274), .B(n7278), .Z(n7379) );
  XOR U9890 ( .A(n7269), .B(n7273), .Z(n7380) );
  XOR U9891 ( .A(n7259), .B(n7268), .Z(n7381) );
  XOR U9892 ( .A(n7382), .B(n7258), .Z(n7259) );
  AND U9893 ( .A(b[20]), .B(a[68]), .Z(n7382) );
  XNOR U9894 ( .A(n7258), .B(n7264), .Z(n7383) );
  XNOR U9895 ( .A(n7263), .B(n7255), .Z(n7384) );
  XNOR U9896 ( .A(n7254), .B(n7250), .Z(n7385) );
  XNOR U9897 ( .A(n7249), .B(n7245), .Z(n7386) );
  XNOR U9898 ( .A(n7244), .B(n7240), .Z(n7387) );
  XNOR U9899 ( .A(n7239), .B(n7235), .Z(n7388) );
  XNOR U9900 ( .A(n7234), .B(n7230), .Z(n7389) );
  XOR U9901 ( .A(n7229), .B(n7226), .Z(n7390) );
  XOR U9902 ( .A(n7391), .B(n7392), .Z(n7226) );
  XOR U9903 ( .A(n7224), .B(n7393), .Z(n7392) );
  XOR U9904 ( .A(n7394), .B(n7395), .Z(n7393) );
  XOR U9905 ( .A(n7396), .B(n7397), .Z(n7395) );
  NAND U9906 ( .A(a[58]), .B(b[30]), .Z(n7397) );
  AND U9907 ( .A(a[57]), .B(b[31]), .Z(n7396) );
  XOR U9908 ( .A(n7398), .B(n7394), .Z(n7391) );
  XOR U9909 ( .A(n7399), .B(n7400), .Z(n7394) );
  ANDN U9910 ( .B(n7401), .A(n7402), .Z(n7399) );
  AND U9911 ( .A(a[59]), .B(b[29]), .Z(n7398) );
  XOR U9912 ( .A(n7403), .B(n7224), .Z(n7225) );
  XOR U9913 ( .A(n7404), .B(n7405), .Z(n7224) );
  AND U9914 ( .A(n7406), .B(n7407), .Z(n7404) );
  AND U9915 ( .A(a[60]), .B(b[28]), .Z(n7403) );
  XOR U9916 ( .A(n7408), .B(n7229), .Z(n7231) );
  XOR U9917 ( .A(n7409), .B(n7410), .Z(n7229) );
  AND U9918 ( .A(n7411), .B(n7412), .Z(n7409) );
  AND U9919 ( .A(a[61]), .B(b[27]), .Z(n7408) );
  XOR U9920 ( .A(n7413), .B(n7234), .Z(n7236) );
  XOR U9921 ( .A(n7414), .B(n7415), .Z(n7234) );
  AND U9922 ( .A(n7416), .B(n7417), .Z(n7414) );
  AND U9923 ( .A(a[62]), .B(b[26]), .Z(n7413) );
  XOR U9924 ( .A(n7418), .B(n7239), .Z(n7241) );
  XOR U9925 ( .A(n7419), .B(n7420), .Z(n7239) );
  AND U9926 ( .A(n7421), .B(n7422), .Z(n7419) );
  AND U9927 ( .A(a[63]), .B(b[25]), .Z(n7418) );
  XOR U9928 ( .A(n7423), .B(n7244), .Z(n7246) );
  XOR U9929 ( .A(n7424), .B(n7425), .Z(n7244) );
  AND U9930 ( .A(n7426), .B(n7427), .Z(n7424) );
  AND U9931 ( .A(a[64]), .B(b[24]), .Z(n7423) );
  XOR U9932 ( .A(n7428), .B(n7249), .Z(n7251) );
  XOR U9933 ( .A(n7429), .B(n7430), .Z(n7249) );
  AND U9934 ( .A(n7431), .B(n7432), .Z(n7429) );
  AND U9935 ( .A(a[65]), .B(b[23]), .Z(n7428) );
  XOR U9936 ( .A(n7433), .B(n7254), .Z(n7256) );
  XOR U9937 ( .A(n7434), .B(n7435), .Z(n7254) );
  AND U9938 ( .A(n7436), .B(n7437), .Z(n7434) );
  AND U9939 ( .A(a[66]), .B(b[22]), .Z(n7433) );
  XOR U9940 ( .A(n7438), .B(n7439), .Z(n7258) );
  AND U9941 ( .A(n7440), .B(n7441), .Z(n7438) );
  XOR U9942 ( .A(n7442), .B(n7263), .Z(n7265) );
  XOR U9943 ( .A(n7443), .B(n7444), .Z(n7263) );
  AND U9944 ( .A(n7445), .B(n7446), .Z(n7443) );
  AND U9945 ( .A(a[67]), .B(b[21]), .Z(n7442) );
  XOR U9946 ( .A(n7448), .B(n7449), .Z(n7268) );
  AND U9947 ( .A(n7450), .B(n7451), .Z(n7448) );
  AND U9948 ( .A(a[69]), .B(b[19]), .Z(n7447) );
  XOR U9949 ( .A(n7453), .B(n7454), .Z(n7273) );
  AND U9950 ( .A(n7455), .B(n7456), .Z(n7453) );
  AND U9951 ( .A(a[70]), .B(b[18]), .Z(n7452) );
  XOR U9952 ( .A(n7458), .B(n7459), .Z(n7278) );
  AND U9953 ( .A(n7460), .B(n7461), .Z(n7458) );
  AND U9954 ( .A(a[71]), .B(b[17]), .Z(n7457) );
  XOR U9955 ( .A(n7463), .B(n7464), .Z(n7283) );
  AND U9956 ( .A(n7465), .B(n7466), .Z(n7463) );
  AND U9957 ( .A(a[72]), .B(b[16]), .Z(n7462) );
  XOR U9958 ( .A(n7468), .B(n7469), .Z(n7288) );
  AND U9959 ( .A(n7470), .B(n7471), .Z(n7468) );
  AND U9960 ( .A(a[73]), .B(b[15]), .Z(n7467) );
  XOR U9961 ( .A(n7473), .B(n7474), .Z(n7293) );
  AND U9962 ( .A(n7475), .B(n7476), .Z(n7473) );
  AND U9963 ( .A(a[74]), .B(b[14]), .Z(n7472) );
  XOR U9964 ( .A(n7478), .B(n7479), .Z(n7298) );
  AND U9965 ( .A(n7480), .B(n7481), .Z(n7478) );
  AND U9966 ( .A(a[75]), .B(b[13]), .Z(n7477) );
  XOR U9967 ( .A(n7483), .B(n7484), .Z(n7303) );
  AND U9968 ( .A(n7485), .B(n7486), .Z(n7483) );
  AND U9969 ( .A(a[76]), .B(b[12]), .Z(n7482) );
  XOR U9970 ( .A(n7488), .B(n7489), .Z(n7308) );
  AND U9971 ( .A(n7490), .B(n7491), .Z(n7488) );
  AND U9972 ( .A(a[77]), .B(b[11]), .Z(n7487) );
  XOR U9973 ( .A(n7493), .B(n7494), .Z(n7313) );
  AND U9974 ( .A(n7495), .B(n7496), .Z(n7493) );
  AND U9975 ( .A(a[78]), .B(b[10]), .Z(n7492) );
  XOR U9976 ( .A(n7498), .B(n7499), .Z(n7318) );
  AND U9977 ( .A(n7500), .B(n7501), .Z(n7498) );
  AND U9978 ( .A(a[79]), .B(b[9]), .Z(n7497) );
  XOR U9979 ( .A(n7503), .B(n7504), .Z(n7323) );
  AND U9980 ( .A(n7505), .B(n7506), .Z(n7503) );
  AND U9981 ( .A(a[80]), .B(b[8]), .Z(n7502) );
  XOR U9982 ( .A(n7508), .B(n7509), .Z(n7328) );
  AND U9983 ( .A(n7510), .B(n7511), .Z(n7508) );
  AND U9984 ( .A(a[81]), .B(b[7]), .Z(n7507) );
  XOR U9985 ( .A(n7513), .B(n7514), .Z(n7333) );
  AND U9986 ( .A(n7515), .B(n7516), .Z(n7513) );
  AND U9987 ( .A(a[82]), .B(b[6]), .Z(n7512) );
  XOR U9988 ( .A(n7518), .B(n7519), .Z(n7338) );
  AND U9989 ( .A(n7520), .B(n7521), .Z(n7518) );
  AND U9990 ( .A(a[83]), .B(b[5]), .Z(n7517) );
  XOR U9991 ( .A(n7523), .B(n7524), .Z(n7343) );
  AND U9992 ( .A(n7525), .B(n7526), .Z(n7523) );
  AND U9993 ( .A(a[84]), .B(b[4]), .Z(n7522) );
  XOR U9994 ( .A(n7528), .B(n7529), .Z(n7348) );
  AND U9995 ( .A(n7530), .B(n7531), .Z(n7528) );
  AND U9996 ( .A(a[85]), .B(b[3]), .Z(n7527) );
  XOR U9997 ( .A(n7533), .B(n7534), .Z(n7353) );
  OR U9998 ( .A(n7535), .B(n7536), .Z(n7534) );
  AND U9999 ( .A(a[86]), .B(b[2]), .Z(n7532) );
  XNOR U10000 ( .A(n7363), .B(n7537), .Z(n7359) );
  NAND U10001 ( .A(a[87]), .B(b[1]), .Z(n7537) );
  IV U10002 ( .A(n7357), .Z(n7363) );
  ANDN U10003 ( .B(n5117), .A(n5119), .Z(n7357) );
  NAND U10004 ( .A(a[87]), .B(b[0]), .Z(n5119) );
  XOR U10005 ( .A(n7535), .B(n7536), .Z(n5117) );
  XOR U10006 ( .A(n7539), .B(n7530), .Z(n7538) );
  XOR U10007 ( .A(n7525), .B(n7529), .Z(n7540) );
  XOR U10008 ( .A(n7520), .B(n7524), .Z(n7541) );
  XOR U10009 ( .A(n7515), .B(n7519), .Z(n7542) );
  XOR U10010 ( .A(n7510), .B(n7514), .Z(n7543) );
  XOR U10011 ( .A(n7505), .B(n7509), .Z(n7544) );
  XOR U10012 ( .A(n7500), .B(n7504), .Z(n7545) );
  XOR U10013 ( .A(n7495), .B(n7499), .Z(n7546) );
  XOR U10014 ( .A(n7490), .B(n7494), .Z(n7547) );
  XOR U10015 ( .A(n7485), .B(n7489), .Z(n7548) );
  XOR U10016 ( .A(n7480), .B(n7484), .Z(n7549) );
  XOR U10017 ( .A(n7475), .B(n7479), .Z(n7550) );
  XOR U10018 ( .A(n7470), .B(n7474), .Z(n7551) );
  XOR U10019 ( .A(n7465), .B(n7469), .Z(n7552) );
  XOR U10020 ( .A(n7460), .B(n7464), .Z(n7553) );
  XOR U10021 ( .A(n7455), .B(n7459), .Z(n7554) );
  XOR U10022 ( .A(n7450), .B(n7454), .Z(n7555) );
  XOR U10023 ( .A(n7440), .B(n7449), .Z(n7556) );
  XOR U10024 ( .A(n7557), .B(n7439), .Z(n7440) );
  AND U10025 ( .A(b[19]), .B(a[68]), .Z(n7557) );
  XNOR U10026 ( .A(n7439), .B(n7445), .Z(n7558) );
  XNOR U10027 ( .A(n7444), .B(n7436), .Z(n7559) );
  XNOR U10028 ( .A(n7435), .B(n7431), .Z(n7560) );
  XNOR U10029 ( .A(n7430), .B(n7426), .Z(n7561) );
  XNOR U10030 ( .A(n7425), .B(n7421), .Z(n7562) );
  XNOR U10031 ( .A(n7420), .B(n7416), .Z(n7563) );
  XNOR U10032 ( .A(n7415), .B(n7411), .Z(n7564) );
  XNOR U10033 ( .A(n7410), .B(n7406), .Z(n7565) );
  XOR U10034 ( .A(n7405), .B(n7402), .Z(n7566) );
  XOR U10035 ( .A(n7567), .B(n7568), .Z(n7402) );
  XOR U10036 ( .A(n7400), .B(n7569), .Z(n7568) );
  XOR U10037 ( .A(n7570), .B(n7571), .Z(n7569) );
  XOR U10038 ( .A(n7572), .B(n7573), .Z(n7571) );
  NAND U10039 ( .A(a[57]), .B(b[30]), .Z(n7573) );
  AND U10040 ( .A(a[56]), .B(b[31]), .Z(n7572) );
  XOR U10041 ( .A(n7574), .B(n7570), .Z(n7567) );
  XOR U10042 ( .A(n7575), .B(n7576), .Z(n7570) );
  ANDN U10043 ( .B(n7577), .A(n7578), .Z(n7575) );
  AND U10044 ( .A(a[58]), .B(b[29]), .Z(n7574) );
  XOR U10045 ( .A(n7579), .B(n7400), .Z(n7401) );
  XOR U10046 ( .A(n7580), .B(n7581), .Z(n7400) );
  AND U10047 ( .A(n7582), .B(n7583), .Z(n7580) );
  AND U10048 ( .A(a[59]), .B(b[28]), .Z(n7579) );
  XOR U10049 ( .A(n7584), .B(n7405), .Z(n7407) );
  XOR U10050 ( .A(n7585), .B(n7586), .Z(n7405) );
  AND U10051 ( .A(n7587), .B(n7588), .Z(n7585) );
  AND U10052 ( .A(a[60]), .B(b[27]), .Z(n7584) );
  XOR U10053 ( .A(n7589), .B(n7410), .Z(n7412) );
  XOR U10054 ( .A(n7590), .B(n7591), .Z(n7410) );
  AND U10055 ( .A(n7592), .B(n7593), .Z(n7590) );
  AND U10056 ( .A(a[61]), .B(b[26]), .Z(n7589) );
  XOR U10057 ( .A(n7594), .B(n7415), .Z(n7417) );
  XOR U10058 ( .A(n7595), .B(n7596), .Z(n7415) );
  AND U10059 ( .A(n7597), .B(n7598), .Z(n7595) );
  AND U10060 ( .A(a[62]), .B(b[25]), .Z(n7594) );
  XOR U10061 ( .A(n7599), .B(n7420), .Z(n7422) );
  XOR U10062 ( .A(n7600), .B(n7601), .Z(n7420) );
  AND U10063 ( .A(n7602), .B(n7603), .Z(n7600) );
  AND U10064 ( .A(a[63]), .B(b[24]), .Z(n7599) );
  XOR U10065 ( .A(n7604), .B(n7425), .Z(n7427) );
  XOR U10066 ( .A(n7605), .B(n7606), .Z(n7425) );
  AND U10067 ( .A(n7607), .B(n7608), .Z(n7605) );
  AND U10068 ( .A(a[64]), .B(b[23]), .Z(n7604) );
  XOR U10069 ( .A(n7609), .B(n7430), .Z(n7432) );
  XOR U10070 ( .A(n7610), .B(n7611), .Z(n7430) );
  AND U10071 ( .A(n7612), .B(n7613), .Z(n7610) );
  AND U10072 ( .A(a[65]), .B(b[22]), .Z(n7609) );
  XOR U10073 ( .A(n7614), .B(n7435), .Z(n7437) );
  XOR U10074 ( .A(n7615), .B(n7616), .Z(n7435) );
  AND U10075 ( .A(n7617), .B(n7618), .Z(n7615) );
  AND U10076 ( .A(a[66]), .B(b[21]), .Z(n7614) );
  XOR U10077 ( .A(n7619), .B(n7620), .Z(n7439) );
  AND U10078 ( .A(n7621), .B(n7622), .Z(n7619) );
  XOR U10079 ( .A(n7623), .B(n7444), .Z(n7446) );
  XOR U10080 ( .A(n7624), .B(n7625), .Z(n7444) );
  AND U10081 ( .A(n7626), .B(n7627), .Z(n7624) );
  AND U10082 ( .A(a[67]), .B(b[20]), .Z(n7623) );
  XOR U10083 ( .A(n7629), .B(n7630), .Z(n7449) );
  AND U10084 ( .A(n7631), .B(n7632), .Z(n7629) );
  AND U10085 ( .A(a[69]), .B(b[18]), .Z(n7628) );
  XOR U10086 ( .A(n7634), .B(n7635), .Z(n7454) );
  AND U10087 ( .A(n7636), .B(n7637), .Z(n7634) );
  AND U10088 ( .A(a[70]), .B(b[17]), .Z(n7633) );
  XOR U10089 ( .A(n7639), .B(n7640), .Z(n7459) );
  AND U10090 ( .A(n7641), .B(n7642), .Z(n7639) );
  AND U10091 ( .A(a[71]), .B(b[16]), .Z(n7638) );
  XOR U10092 ( .A(n7644), .B(n7645), .Z(n7464) );
  AND U10093 ( .A(n7646), .B(n7647), .Z(n7644) );
  AND U10094 ( .A(a[72]), .B(b[15]), .Z(n7643) );
  XOR U10095 ( .A(n7649), .B(n7650), .Z(n7469) );
  AND U10096 ( .A(n7651), .B(n7652), .Z(n7649) );
  AND U10097 ( .A(a[73]), .B(b[14]), .Z(n7648) );
  XOR U10098 ( .A(n7654), .B(n7655), .Z(n7474) );
  AND U10099 ( .A(n7656), .B(n7657), .Z(n7654) );
  AND U10100 ( .A(a[74]), .B(b[13]), .Z(n7653) );
  XOR U10101 ( .A(n7659), .B(n7660), .Z(n7479) );
  AND U10102 ( .A(n7661), .B(n7662), .Z(n7659) );
  AND U10103 ( .A(a[75]), .B(b[12]), .Z(n7658) );
  XOR U10104 ( .A(n7664), .B(n7665), .Z(n7484) );
  AND U10105 ( .A(n7666), .B(n7667), .Z(n7664) );
  AND U10106 ( .A(a[76]), .B(b[11]), .Z(n7663) );
  XOR U10107 ( .A(n7669), .B(n7670), .Z(n7489) );
  AND U10108 ( .A(n7671), .B(n7672), .Z(n7669) );
  AND U10109 ( .A(a[77]), .B(b[10]), .Z(n7668) );
  XOR U10110 ( .A(n7674), .B(n7675), .Z(n7494) );
  AND U10111 ( .A(n7676), .B(n7677), .Z(n7674) );
  AND U10112 ( .A(a[78]), .B(b[9]), .Z(n7673) );
  XOR U10113 ( .A(n7679), .B(n7680), .Z(n7499) );
  AND U10114 ( .A(n7681), .B(n7682), .Z(n7679) );
  AND U10115 ( .A(a[79]), .B(b[8]), .Z(n7678) );
  XOR U10116 ( .A(n7684), .B(n7685), .Z(n7504) );
  AND U10117 ( .A(n7686), .B(n7687), .Z(n7684) );
  AND U10118 ( .A(a[80]), .B(b[7]), .Z(n7683) );
  XOR U10119 ( .A(n7689), .B(n7690), .Z(n7509) );
  AND U10120 ( .A(n7691), .B(n7692), .Z(n7689) );
  AND U10121 ( .A(a[81]), .B(b[6]), .Z(n7688) );
  XOR U10122 ( .A(n7694), .B(n7695), .Z(n7514) );
  AND U10123 ( .A(n7696), .B(n7697), .Z(n7694) );
  AND U10124 ( .A(a[82]), .B(b[5]), .Z(n7693) );
  XOR U10125 ( .A(n7699), .B(n7700), .Z(n7519) );
  AND U10126 ( .A(n7701), .B(n7702), .Z(n7699) );
  AND U10127 ( .A(a[83]), .B(b[4]), .Z(n7698) );
  XOR U10128 ( .A(n7704), .B(n7705), .Z(n7524) );
  AND U10129 ( .A(n7706), .B(n7707), .Z(n7704) );
  AND U10130 ( .A(a[84]), .B(b[3]), .Z(n7703) );
  XOR U10131 ( .A(n7709), .B(n7710), .Z(n7529) );
  OR U10132 ( .A(n7711), .B(n7712), .Z(n7710) );
  AND U10133 ( .A(a[85]), .B(b[2]), .Z(n7708) );
  XNOR U10134 ( .A(n7539), .B(n7713), .Z(n7535) );
  NAND U10135 ( .A(a[86]), .B(b[1]), .Z(n7713) );
  IV U10136 ( .A(n7533), .Z(n7539) );
  ANDN U10137 ( .B(n5122), .A(n5124), .Z(n7533) );
  NAND U10138 ( .A(a[86]), .B(b[0]), .Z(n5124) );
  XOR U10139 ( .A(n7711), .B(n7712), .Z(n5122) );
  XOR U10140 ( .A(n7715), .B(n7706), .Z(n7714) );
  XOR U10141 ( .A(n7701), .B(n7705), .Z(n7716) );
  XOR U10142 ( .A(n7696), .B(n7700), .Z(n7717) );
  XOR U10143 ( .A(n7691), .B(n7695), .Z(n7718) );
  XOR U10144 ( .A(n7686), .B(n7690), .Z(n7719) );
  XOR U10145 ( .A(n7681), .B(n7685), .Z(n7720) );
  XOR U10146 ( .A(n7676), .B(n7680), .Z(n7721) );
  XOR U10147 ( .A(n7671), .B(n7675), .Z(n7722) );
  XOR U10148 ( .A(n7666), .B(n7670), .Z(n7723) );
  XOR U10149 ( .A(n7661), .B(n7665), .Z(n7724) );
  XOR U10150 ( .A(n7656), .B(n7660), .Z(n7725) );
  XOR U10151 ( .A(n7651), .B(n7655), .Z(n7726) );
  XOR U10152 ( .A(n7646), .B(n7650), .Z(n7727) );
  XOR U10153 ( .A(n7641), .B(n7645), .Z(n7728) );
  XOR U10154 ( .A(n7636), .B(n7640), .Z(n7729) );
  XOR U10155 ( .A(n7631), .B(n7635), .Z(n7730) );
  XOR U10156 ( .A(n7621), .B(n7630), .Z(n7731) );
  XOR U10157 ( .A(n7732), .B(n7620), .Z(n7621) );
  AND U10158 ( .A(b[18]), .B(a[68]), .Z(n7732) );
  XNOR U10159 ( .A(n7620), .B(n7626), .Z(n7733) );
  XNOR U10160 ( .A(n7625), .B(n7617), .Z(n7734) );
  XNOR U10161 ( .A(n7616), .B(n7612), .Z(n7735) );
  XNOR U10162 ( .A(n7611), .B(n7607), .Z(n7736) );
  XNOR U10163 ( .A(n7606), .B(n7602), .Z(n7737) );
  XNOR U10164 ( .A(n7601), .B(n7597), .Z(n7738) );
  XNOR U10165 ( .A(n7596), .B(n7592), .Z(n7739) );
  XNOR U10166 ( .A(n7591), .B(n7587), .Z(n7740) );
  XNOR U10167 ( .A(n7586), .B(n7582), .Z(n7741) );
  XOR U10168 ( .A(n7581), .B(n7578), .Z(n7742) );
  XOR U10169 ( .A(n7743), .B(n7744), .Z(n7578) );
  XOR U10170 ( .A(n7576), .B(n7745), .Z(n7744) );
  XOR U10171 ( .A(n7746), .B(n7747), .Z(n7745) );
  XOR U10172 ( .A(n7748), .B(n7749), .Z(n7747) );
  NAND U10173 ( .A(a[56]), .B(b[30]), .Z(n7749) );
  AND U10174 ( .A(a[55]), .B(b[31]), .Z(n7748) );
  XOR U10175 ( .A(n7750), .B(n7746), .Z(n7743) );
  XOR U10176 ( .A(n7751), .B(n7752), .Z(n7746) );
  ANDN U10177 ( .B(n7753), .A(n7754), .Z(n7751) );
  AND U10178 ( .A(a[57]), .B(b[29]), .Z(n7750) );
  XOR U10179 ( .A(n7755), .B(n7576), .Z(n7577) );
  XOR U10180 ( .A(n7756), .B(n7757), .Z(n7576) );
  AND U10181 ( .A(n7758), .B(n7759), .Z(n7756) );
  AND U10182 ( .A(a[58]), .B(b[28]), .Z(n7755) );
  XOR U10183 ( .A(n7760), .B(n7581), .Z(n7583) );
  XOR U10184 ( .A(n7761), .B(n7762), .Z(n7581) );
  AND U10185 ( .A(n7763), .B(n7764), .Z(n7761) );
  AND U10186 ( .A(a[59]), .B(b[27]), .Z(n7760) );
  XOR U10187 ( .A(n7765), .B(n7586), .Z(n7588) );
  XOR U10188 ( .A(n7766), .B(n7767), .Z(n7586) );
  AND U10189 ( .A(n7768), .B(n7769), .Z(n7766) );
  AND U10190 ( .A(a[60]), .B(b[26]), .Z(n7765) );
  XOR U10191 ( .A(n7770), .B(n7591), .Z(n7593) );
  XOR U10192 ( .A(n7771), .B(n7772), .Z(n7591) );
  AND U10193 ( .A(n7773), .B(n7774), .Z(n7771) );
  AND U10194 ( .A(a[61]), .B(b[25]), .Z(n7770) );
  XOR U10195 ( .A(n7775), .B(n7596), .Z(n7598) );
  XOR U10196 ( .A(n7776), .B(n7777), .Z(n7596) );
  AND U10197 ( .A(n7778), .B(n7779), .Z(n7776) );
  AND U10198 ( .A(a[62]), .B(b[24]), .Z(n7775) );
  XOR U10199 ( .A(n7780), .B(n7601), .Z(n7603) );
  XOR U10200 ( .A(n7781), .B(n7782), .Z(n7601) );
  AND U10201 ( .A(n7783), .B(n7784), .Z(n7781) );
  AND U10202 ( .A(a[63]), .B(b[23]), .Z(n7780) );
  XOR U10203 ( .A(n7785), .B(n7606), .Z(n7608) );
  XOR U10204 ( .A(n7786), .B(n7787), .Z(n7606) );
  AND U10205 ( .A(n7788), .B(n7789), .Z(n7786) );
  AND U10206 ( .A(a[64]), .B(b[22]), .Z(n7785) );
  XOR U10207 ( .A(n7790), .B(n7611), .Z(n7613) );
  XOR U10208 ( .A(n7791), .B(n7792), .Z(n7611) );
  AND U10209 ( .A(n7793), .B(n7794), .Z(n7791) );
  AND U10210 ( .A(a[65]), .B(b[21]), .Z(n7790) );
  XOR U10211 ( .A(n7795), .B(n7616), .Z(n7618) );
  XOR U10212 ( .A(n7796), .B(n7797), .Z(n7616) );
  AND U10213 ( .A(n7798), .B(n7799), .Z(n7796) );
  AND U10214 ( .A(a[66]), .B(b[20]), .Z(n7795) );
  XOR U10215 ( .A(n7800), .B(n7801), .Z(n7620) );
  AND U10216 ( .A(n7802), .B(n7803), .Z(n7800) );
  XOR U10217 ( .A(n7804), .B(n7625), .Z(n7627) );
  XOR U10218 ( .A(n7805), .B(n7806), .Z(n7625) );
  AND U10219 ( .A(n7807), .B(n7808), .Z(n7805) );
  AND U10220 ( .A(a[67]), .B(b[19]), .Z(n7804) );
  XOR U10221 ( .A(n7810), .B(n7811), .Z(n7630) );
  AND U10222 ( .A(n7812), .B(n7813), .Z(n7810) );
  AND U10223 ( .A(a[69]), .B(b[17]), .Z(n7809) );
  XOR U10224 ( .A(n7815), .B(n7816), .Z(n7635) );
  AND U10225 ( .A(n7817), .B(n7818), .Z(n7815) );
  AND U10226 ( .A(a[70]), .B(b[16]), .Z(n7814) );
  XOR U10227 ( .A(n7820), .B(n7821), .Z(n7640) );
  AND U10228 ( .A(n7822), .B(n7823), .Z(n7820) );
  AND U10229 ( .A(a[71]), .B(b[15]), .Z(n7819) );
  XOR U10230 ( .A(n7825), .B(n7826), .Z(n7645) );
  AND U10231 ( .A(n7827), .B(n7828), .Z(n7825) );
  AND U10232 ( .A(a[72]), .B(b[14]), .Z(n7824) );
  XOR U10233 ( .A(n7830), .B(n7831), .Z(n7650) );
  AND U10234 ( .A(n7832), .B(n7833), .Z(n7830) );
  AND U10235 ( .A(a[73]), .B(b[13]), .Z(n7829) );
  XOR U10236 ( .A(n7835), .B(n7836), .Z(n7655) );
  AND U10237 ( .A(n7837), .B(n7838), .Z(n7835) );
  AND U10238 ( .A(a[74]), .B(b[12]), .Z(n7834) );
  XOR U10239 ( .A(n7840), .B(n7841), .Z(n7660) );
  AND U10240 ( .A(n7842), .B(n7843), .Z(n7840) );
  AND U10241 ( .A(a[75]), .B(b[11]), .Z(n7839) );
  XOR U10242 ( .A(n7845), .B(n7846), .Z(n7665) );
  AND U10243 ( .A(n7847), .B(n7848), .Z(n7845) );
  AND U10244 ( .A(a[76]), .B(b[10]), .Z(n7844) );
  XOR U10245 ( .A(n7850), .B(n7851), .Z(n7670) );
  AND U10246 ( .A(n7852), .B(n7853), .Z(n7850) );
  AND U10247 ( .A(a[77]), .B(b[9]), .Z(n7849) );
  XOR U10248 ( .A(n7855), .B(n7856), .Z(n7675) );
  AND U10249 ( .A(n7857), .B(n7858), .Z(n7855) );
  AND U10250 ( .A(a[78]), .B(b[8]), .Z(n7854) );
  XOR U10251 ( .A(n7860), .B(n7861), .Z(n7680) );
  AND U10252 ( .A(n7862), .B(n7863), .Z(n7860) );
  AND U10253 ( .A(a[79]), .B(b[7]), .Z(n7859) );
  XOR U10254 ( .A(n7865), .B(n7866), .Z(n7685) );
  AND U10255 ( .A(n7867), .B(n7868), .Z(n7865) );
  AND U10256 ( .A(a[80]), .B(b[6]), .Z(n7864) );
  XOR U10257 ( .A(n7870), .B(n7871), .Z(n7690) );
  AND U10258 ( .A(n7872), .B(n7873), .Z(n7870) );
  AND U10259 ( .A(a[81]), .B(b[5]), .Z(n7869) );
  XOR U10260 ( .A(n7875), .B(n7876), .Z(n7695) );
  AND U10261 ( .A(n7877), .B(n7878), .Z(n7875) );
  AND U10262 ( .A(a[82]), .B(b[4]), .Z(n7874) );
  XOR U10263 ( .A(n7880), .B(n7881), .Z(n7700) );
  AND U10264 ( .A(n7882), .B(n7883), .Z(n7880) );
  AND U10265 ( .A(a[83]), .B(b[3]), .Z(n7879) );
  XOR U10266 ( .A(n7885), .B(n7886), .Z(n7705) );
  OR U10267 ( .A(n7887), .B(n7888), .Z(n7886) );
  AND U10268 ( .A(a[84]), .B(b[2]), .Z(n7884) );
  XNOR U10269 ( .A(n7715), .B(n7889), .Z(n7711) );
  NAND U10270 ( .A(a[85]), .B(b[1]), .Z(n7889) );
  IV U10271 ( .A(n7709), .Z(n7715) );
  ANDN U10272 ( .B(n5127), .A(n5129), .Z(n7709) );
  NAND U10273 ( .A(a[85]), .B(b[0]), .Z(n5129) );
  XOR U10274 ( .A(n7887), .B(n7888), .Z(n5127) );
  XOR U10275 ( .A(n7891), .B(n7882), .Z(n7890) );
  XOR U10276 ( .A(n7877), .B(n7881), .Z(n7892) );
  XOR U10277 ( .A(n7872), .B(n7876), .Z(n7893) );
  XOR U10278 ( .A(n7867), .B(n7871), .Z(n7894) );
  XOR U10279 ( .A(n7862), .B(n7866), .Z(n7895) );
  XOR U10280 ( .A(n7857), .B(n7861), .Z(n7896) );
  XOR U10281 ( .A(n7852), .B(n7856), .Z(n7897) );
  XOR U10282 ( .A(n7847), .B(n7851), .Z(n7898) );
  XOR U10283 ( .A(n7842), .B(n7846), .Z(n7899) );
  XOR U10284 ( .A(n7837), .B(n7841), .Z(n7900) );
  XOR U10285 ( .A(n7832), .B(n7836), .Z(n7901) );
  XOR U10286 ( .A(n7827), .B(n7831), .Z(n7902) );
  XOR U10287 ( .A(n7822), .B(n7826), .Z(n7903) );
  XOR U10288 ( .A(n7817), .B(n7821), .Z(n7904) );
  XOR U10289 ( .A(n7812), .B(n7816), .Z(n7905) );
  XOR U10290 ( .A(n7802), .B(n7811), .Z(n7906) );
  XOR U10291 ( .A(n7907), .B(n7801), .Z(n7802) );
  AND U10292 ( .A(b[17]), .B(a[68]), .Z(n7907) );
  XNOR U10293 ( .A(n7801), .B(n7807), .Z(n7908) );
  XNOR U10294 ( .A(n7806), .B(n7798), .Z(n7909) );
  XNOR U10295 ( .A(n7797), .B(n7793), .Z(n7910) );
  XNOR U10296 ( .A(n7792), .B(n7788), .Z(n7911) );
  XNOR U10297 ( .A(n7787), .B(n7783), .Z(n7912) );
  XNOR U10298 ( .A(n7782), .B(n7778), .Z(n7913) );
  XNOR U10299 ( .A(n7777), .B(n7773), .Z(n7914) );
  XNOR U10300 ( .A(n7772), .B(n7768), .Z(n7915) );
  XNOR U10301 ( .A(n7767), .B(n7763), .Z(n7916) );
  XNOR U10302 ( .A(n7762), .B(n7758), .Z(n7917) );
  XOR U10303 ( .A(n7757), .B(n7754), .Z(n7918) );
  XOR U10304 ( .A(n7919), .B(n7920), .Z(n7754) );
  XOR U10305 ( .A(n7752), .B(n7921), .Z(n7920) );
  XOR U10306 ( .A(n7922), .B(n7923), .Z(n7921) );
  XOR U10307 ( .A(n7924), .B(n7925), .Z(n7923) );
  NAND U10308 ( .A(a[55]), .B(b[30]), .Z(n7925) );
  AND U10309 ( .A(a[54]), .B(b[31]), .Z(n7924) );
  XOR U10310 ( .A(n7926), .B(n7922), .Z(n7919) );
  XOR U10311 ( .A(n7927), .B(n7928), .Z(n7922) );
  ANDN U10312 ( .B(n7929), .A(n7930), .Z(n7927) );
  AND U10313 ( .A(a[56]), .B(b[29]), .Z(n7926) );
  XOR U10314 ( .A(n7931), .B(n7752), .Z(n7753) );
  XOR U10315 ( .A(n7932), .B(n7933), .Z(n7752) );
  AND U10316 ( .A(n7934), .B(n7935), .Z(n7932) );
  AND U10317 ( .A(a[57]), .B(b[28]), .Z(n7931) );
  XOR U10318 ( .A(n7936), .B(n7757), .Z(n7759) );
  XOR U10319 ( .A(n7937), .B(n7938), .Z(n7757) );
  AND U10320 ( .A(n7939), .B(n7940), .Z(n7937) );
  AND U10321 ( .A(a[58]), .B(b[27]), .Z(n7936) );
  XOR U10322 ( .A(n7941), .B(n7762), .Z(n7764) );
  XOR U10323 ( .A(n7942), .B(n7943), .Z(n7762) );
  AND U10324 ( .A(n7944), .B(n7945), .Z(n7942) );
  AND U10325 ( .A(a[59]), .B(b[26]), .Z(n7941) );
  XOR U10326 ( .A(n7946), .B(n7767), .Z(n7769) );
  XOR U10327 ( .A(n7947), .B(n7948), .Z(n7767) );
  AND U10328 ( .A(n7949), .B(n7950), .Z(n7947) );
  AND U10329 ( .A(a[60]), .B(b[25]), .Z(n7946) );
  XOR U10330 ( .A(n7951), .B(n7772), .Z(n7774) );
  XOR U10331 ( .A(n7952), .B(n7953), .Z(n7772) );
  AND U10332 ( .A(n7954), .B(n7955), .Z(n7952) );
  AND U10333 ( .A(a[61]), .B(b[24]), .Z(n7951) );
  XOR U10334 ( .A(n7956), .B(n7777), .Z(n7779) );
  XOR U10335 ( .A(n7957), .B(n7958), .Z(n7777) );
  AND U10336 ( .A(n7959), .B(n7960), .Z(n7957) );
  AND U10337 ( .A(a[62]), .B(b[23]), .Z(n7956) );
  XOR U10338 ( .A(n7961), .B(n7782), .Z(n7784) );
  XOR U10339 ( .A(n7962), .B(n7963), .Z(n7782) );
  AND U10340 ( .A(n7964), .B(n7965), .Z(n7962) );
  AND U10341 ( .A(a[63]), .B(b[22]), .Z(n7961) );
  XOR U10342 ( .A(n7966), .B(n7787), .Z(n7789) );
  XOR U10343 ( .A(n7967), .B(n7968), .Z(n7787) );
  AND U10344 ( .A(n7969), .B(n7970), .Z(n7967) );
  AND U10345 ( .A(a[64]), .B(b[21]), .Z(n7966) );
  XOR U10346 ( .A(n7971), .B(n7792), .Z(n7794) );
  XOR U10347 ( .A(n7972), .B(n7973), .Z(n7792) );
  AND U10348 ( .A(n7974), .B(n7975), .Z(n7972) );
  AND U10349 ( .A(a[65]), .B(b[20]), .Z(n7971) );
  XOR U10350 ( .A(n7976), .B(n7797), .Z(n7799) );
  XOR U10351 ( .A(n7977), .B(n7978), .Z(n7797) );
  AND U10352 ( .A(n7979), .B(n7980), .Z(n7977) );
  AND U10353 ( .A(a[66]), .B(b[19]), .Z(n7976) );
  XOR U10354 ( .A(n7981), .B(n7982), .Z(n7801) );
  AND U10355 ( .A(n7983), .B(n7984), .Z(n7981) );
  XOR U10356 ( .A(n7985), .B(n7806), .Z(n7808) );
  XOR U10357 ( .A(n7986), .B(n7987), .Z(n7806) );
  AND U10358 ( .A(n7988), .B(n7989), .Z(n7986) );
  AND U10359 ( .A(a[67]), .B(b[18]), .Z(n7985) );
  XOR U10360 ( .A(n7991), .B(n7992), .Z(n7811) );
  AND U10361 ( .A(n7993), .B(n7994), .Z(n7991) );
  AND U10362 ( .A(a[69]), .B(b[16]), .Z(n7990) );
  XOR U10363 ( .A(n7996), .B(n7997), .Z(n7816) );
  AND U10364 ( .A(n7998), .B(n7999), .Z(n7996) );
  AND U10365 ( .A(a[70]), .B(b[15]), .Z(n7995) );
  XOR U10366 ( .A(n8001), .B(n8002), .Z(n7821) );
  AND U10367 ( .A(n8003), .B(n8004), .Z(n8001) );
  AND U10368 ( .A(a[71]), .B(b[14]), .Z(n8000) );
  XOR U10369 ( .A(n8006), .B(n8007), .Z(n7826) );
  AND U10370 ( .A(n8008), .B(n8009), .Z(n8006) );
  AND U10371 ( .A(a[72]), .B(b[13]), .Z(n8005) );
  XOR U10372 ( .A(n8011), .B(n8012), .Z(n7831) );
  AND U10373 ( .A(n8013), .B(n8014), .Z(n8011) );
  AND U10374 ( .A(a[73]), .B(b[12]), .Z(n8010) );
  XOR U10375 ( .A(n8016), .B(n8017), .Z(n7836) );
  AND U10376 ( .A(n8018), .B(n8019), .Z(n8016) );
  AND U10377 ( .A(a[74]), .B(b[11]), .Z(n8015) );
  XOR U10378 ( .A(n8021), .B(n8022), .Z(n7841) );
  AND U10379 ( .A(n8023), .B(n8024), .Z(n8021) );
  AND U10380 ( .A(a[75]), .B(b[10]), .Z(n8020) );
  XOR U10381 ( .A(n8026), .B(n8027), .Z(n7846) );
  AND U10382 ( .A(n8028), .B(n8029), .Z(n8026) );
  AND U10383 ( .A(a[76]), .B(b[9]), .Z(n8025) );
  XOR U10384 ( .A(n8031), .B(n8032), .Z(n7851) );
  AND U10385 ( .A(n8033), .B(n8034), .Z(n8031) );
  AND U10386 ( .A(a[77]), .B(b[8]), .Z(n8030) );
  XOR U10387 ( .A(n8036), .B(n8037), .Z(n7856) );
  AND U10388 ( .A(n8038), .B(n8039), .Z(n8036) );
  AND U10389 ( .A(a[78]), .B(b[7]), .Z(n8035) );
  XOR U10390 ( .A(n8041), .B(n8042), .Z(n7861) );
  AND U10391 ( .A(n8043), .B(n8044), .Z(n8041) );
  AND U10392 ( .A(a[79]), .B(b[6]), .Z(n8040) );
  XOR U10393 ( .A(n8046), .B(n8047), .Z(n7866) );
  AND U10394 ( .A(n8048), .B(n8049), .Z(n8046) );
  AND U10395 ( .A(a[80]), .B(b[5]), .Z(n8045) );
  XOR U10396 ( .A(n8051), .B(n8052), .Z(n7871) );
  AND U10397 ( .A(n8053), .B(n8054), .Z(n8051) );
  AND U10398 ( .A(a[81]), .B(b[4]), .Z(n8050) );
  XOR U10399 ( .A(n8056), .B(n8057), .Z(n7876) );
  AND U10400 ( .A(n8058), .B(n8059), .Z(n8056) );
  AND U10401 ( .A(a[82]), .B(b[3]), .Z(n8055) );
  XOR U10402 ( .A(n8061), .B(n8062), .Z(n7881) );
  OR U10403 ( .A(n8063), .B(n8064), .Z(n8062) );
  AND U10404 ( .A(a[83]), .B(b[2]), .Z(n8060) );
  XNOR U10405 ( .A(n7891), .B(n8065), .Z(n7887) );
  NAND U10406 ( .A(a[84]), .B(b[1]), .Z(n8065) );
  IV U10407 ( .A(n7885), .Z(n7891) );
  ANDN U10408 ( .B(n5132), .A(n5134), .Z(n7885) );
  NAND U10409 ( .A(a[84]), .B(b[0]), .Z(n5134) );
  XOR U10410 ( .A(n8063), .B(n8064), .Z(n5132) );
  XOR U10411 ( .A(n8067), .B(n8058), .Z(n8066) );
  XOR U10412 ( .A(n8053), .B(n8057), .Z(n8068) );
  XOR U10413 ( .A(n8048), .B(n8052), .Z(n8069) );
  XOR U10414 ( .A(n8043), .B(n8047), .Z(n8070) );
  XOR U10415 ( .A(n8038), .B(n8042), .Z(n8071) );
  XOR U10416 ( .A(n8033), .B(n8037), .Z(n8072) );
  XOR U10417 ( .A(n8028), .B(n8032), .Z(n8073) );
  XOR U10418 ( .A(n8023), .B(n8027), .Z(n8074) );
  XOR U10419 ( .A(n8018), .B(n8022), .Z(n8075) );
  XOR U10420 ( .A(n8013), .B(n8017), .Z(n8076) );
  XOR U10421 ( .A(n8008), .B(n8012), .Z(n8077) );
  XOR U10422 ( .A(n8003), .B(n8007), .Z(n8078) );
  XOR U10423 ( .A(n7998), .B(n8002), .Z(n8079) );
  XOR U10424 ( .A(n7993), .B(n7997), .Z(n8080) );
  XOR U10425 ( .A(n7983), .B(n7992), .Z(n8081) );
  XOR U10426 ( .A(n8082), .B(n7982), .Z(n7983) );
  AND U10427 ( .A(b[16]), .B(a[68]), .Z(n8082) );
  XNOR U10428 ( .A(n7982), .B(n7988), .Z(n8083) );
  XNOR U10429 ( .A(n7987), .B(n7979), .Z(n8084) );
  XNOR U10430 ( .A(n7978), .B(n7974), .Z(n8085) );
  XNOR U10431 ( .A(n7973), .B(n7969), .Z(n8086) );
  XNOR U10432 ( .A(n7968), .B(n7964), .Z(n8087) );
  XNOR U10433 ( .A(n7963), .B(n7959), .Z(n8088) );
  XNOR U10434 ( .A(n7958), .B(n7954), .Z(n8089) );
  XNOR U10435 ( .A(n7953), .B(n7949), .Z(n8090) );
  XNOR U10436 ( .A(n7948), .B(n7944), .Z(n8091) );
  XNOR U10437 ( .A(n7943), .B(n7939), .Z(n8092) );
  XNOR U10438 ( .A(n7938), .B(n7934), .Z(n8093) );
  XOR U10439 ( .A(n7933), .B(n7930), .Z(n8094) );
  XOR U10440 ( .A(n8095), .B(n8096), .Z(n7930) );
  XOR U10441 ( .A(n7928), .B(n8097), .Z(n8096) );
  XOR U10442 ( .A(n8098), .B(n8099), .Z(n8097) );
  XOR U10443 ( .A(n8100), .B(n8101), .Z(n8099) );
  NAND U10444 ( .A(a[54]), .B(b[30]), .Z(n8101) );
  AND U10445 ( .A(a[53]), .B(b[31]), .Z(n8100) );
  XOR U10446 ( .A(n8102), .B(n8098), .Z(n8095) );
  XOR U10447 ( .A(n8103), .B(n8104), .Z(n8098) );
  ANDN U10448 ( .B(n8105), .A(n8106), .Z(n8103) );
  AND U10449 ( .A(a[55]), .B(b[29]), .Z(n8102) );
  XOR U10450 ( .A(n8107), .B(n7928), .Z(n7929) );
  XOR U10451 ( .A(n8108), .B(n8109), .Z(n7928) );
  AND U10452 ( .A(n8110), .B(n8111), .Z(n8108) );
  AND U10453 ( .A(a[56]), .B(b[28]), .Z(n8107) );
  XOR U10454 ( .A(n8112), .B(n7933), .Z(n7935) );
  XOR U10455 ( .A(n8113), .B(n8114), .Z(n7933) );
  AND U10456 ( .A(n8115), .B(n8116), .Z(n8113) );
  AND U10457 ( .A(a[57]), .B(b[27]), .Z(n8112) );
  XOR U10458 ( .A(n8117), .B(n7938), .Z(n7940) );
  XOR U10459 ( .A(n8118), .B(n8119), .Z(n7938) );
  AND U10460 ( .A(n8120), .B(n8121), .Z(n8118) );
  AND U10461 ( .A(a[58]), .B(b[26]), .Z(n8117) );
  XOR U10462 ( .A(n8122), .B(n7943), .Z(n7945) );
  XOR U10463 ( .A(n8123), .B(n8124), .Z(n7943) );
  AND U10464 ( .A(n8125), .B(n8126), .Z(n8123) );
  AND U10465 ( .A(a[59]), .B(b[25]), .Z(n8122) );
  XOR U10466 ( .A(n8127), .B(n7948), .Z(n7950) );
  XOR U10467 ( .A(n8128), .B(n8129), .Z(n7948) );
  AND U10468 ( .A(n8130), .B(n8131), .Z(n8128) );
  AND U10469 ( .A(a[60]), .B(b[24]), .Z(n8127) );
  XOR U10470 ( .A(n8132), .B(n7953), .Z(n7955) );
  XOR U10471 ( .A(n8133), .B(n8134), .Z(n7953) );
  AND U10472 ( .A(n8135), .B(n8136), .Z(n8133) );
  AND U10473 ( .A(a[61]), .B(b[23]), .Z(n8132) );
  XOR U10474 ( .A(n8137), .B(n7958), .Z(n7960) );
  XOR U10475 ( .A(n8138), .B(n8139), .Z(n7958) );
  AND U10476 ( .A(n8140), .B(n8141), .Z(n8138) );
  AND U10477 ( .A(a[62]), .B(b[22]), .Z(n8137) );
  XOR U10478 ( .A(n8142), .B(n7963), .Z(n7965) );
  XOR U10479 ( .A(n8143), .B(n8144), .Z(n7963) );
  AND U10480 ( .A(n8145), .B(n8146), .Z(n8143) );
  AND U10481 ( .A(a[63]), .B(b[21]), .Z(n8142) );
  XOR U10482 ( .A(n8147), .B(n7968), .Z(n7970) );
  XOR U10483 ( .A(n8148), .B(n8149), .Z(n7968) );
  AND U10484 ( .A(n8150), .B(n8151), .Z(n8148) );
  AND U10485 ( .A(a[64]), .B(b[20]), .Z(n8147) );
  XOR U10486 ( .A(n8152), .B(n7973), .Z(n7975) );
  XOR U10487 ( .A(n8153), .B(n8154), .Z(n7973) );
  AND U10488 ( .A(n8155), .B(n8156), .Z(n8153) );
  AND U10489 ( .A(a[65]), .B(b[19]), .Z(n8152) );
  XOR U10490 ( .A(n8157), .B(n7978), .Z(n7980) );
  XOR U10491 ( .A(n8158), .B(n8159), .Z(n7978) );
  AND U10492 ( .A(n8160), .B(n8161), .Z(n8158) );
  AND U10493 ( .A(a[66]), .B(b[18]), .Z(n8157) );
  XOR U10494 ( .A(n8162), .B(n8163), .Z(n7982) );
  AND U10495 ( .A(n8164), .B(n8165), .Z(n8162) );
  XOR U10496 ( .A(n8166), .B(n7987), .Z(n7989) );
  XOR U10497 ( .A(n8167), .B(n8168), .Z(n7987) );
  AND U10498 ( .A(n8169), .B(n8170), .Z(n8167) );
  AND U10499 ( .A(a[67]), .B(b[17]), .Z(n8166) );
  XOR U10500 ( .A(n8172), .B(n8173), .Z(n7992) );
  AND U10501 ( .A(n8174), .B(n8175), .Z(n8172) );
  AND U10502 ( .A(a[69]), .B(b[15]), .Z(n8171) );
  XOR U10503 ( .A(n8177), .B(n8178), .Z(n7997) );
  AND U10504 ( .A(n8179), .B(n8180), .Z(n8177) );
  AND U10505 ( .A(a[70]), .B(b[14]), .Z(n8176) );
  XOR U10506 ( .A(n8182), .B(n8183), .Z(n8002) );
  AND U10507 ( .A(n8184), .B(n8185), .Z(n8182) );
  AND U10508 ( .A(a[71]), .B(b[13]), .Z(n8181) );
  XOR U10509 ( .A(n8187), .B(n8188), .Z(n8007) );
  AND U10510 ( .A(n8189), .B(n8190), .Z(n8187) );
  AND U10511 ( .A(a[72]), .B(b[12]), .Z(n8186) );
  XOR U10512 ( .A(n8192), .B(n8193), .Z(n8012) );
  AND U10513 ( .A(n8194), .B(n8195), .Z(n8192) );
  AND U10514 ( .A(a[73]), .B(b[11]), .Z(n8191) );
  XOR U10515 ( .A(n8197), .B(n8198), .Z(n8017) );
  AND U10516 ( .A(n8199), .B(n8200), .Z(n8197) );
  AND U10517 ( .A(a[74]), .B(b[10]), .Z(n8196) );
  XOR U10518 ( .A(n8202), .B(n8203), .Z(n8022) );
  AND U10519 ( .A(n8204), .B(n8205), .Z(n8202) );
  AND U10520 ( .A(a[75]), .B(b[9]), .Z(n8201) );
  XOR U10521 ( .A(n8207), .B(n8208), .Z(n8027) );
  AND U10522 ( .A(n8209), .B(n8210), .Z(n8207) );
  AND U10523 ( .A(a[76]), .B(b[8]), .Z(n8206) );
  XOR U10524 ( .A(n8212), .B(n8213), .Z(n8032) );
  AND U10525 ( .A(n8214), .B(n8215), .Z(n8212) );
  AND U10526 ( .A(a[77]), .B(b[7]), .Z(n8211) );
  XOR U10527 ( .A(n8217), .B(n8218), .Z(n8037) );
  AND U10528 ( .A(n8219), .B(n8220), .Z(n8217) );
  AND U10529 ( .A(a[78]), .B(b[6]), .Z(n8216) );
  XOR U10530 ( .A(n8222), .B(n8223), .Z(n8042) );
  AND U10531 ( .A(n8224), .B(n8225), .Z(n8222) );
  AND U10532 ( .A(a[79]), .B(b[5]), .Z(n8221) );
  XOR U10533 ( .A(n8227), .B(n8228), .Z(n8047) );
  AND U10534 ( .A(n8229), .B(n8230), .Z(n8227) );
  AND U10535 ( .A(a[80]), .B(b[4]), .Z(n8226) );
  XOR U10536 ( .A(n8232), .B(n8233), .Z(n8052) );
  AND U10537 ( .A(n8234), .B(n8235), .Z(n8232) );
  AND U10538 ( .A(a[81]), .B(b[3]), .Z(n8231) );
  XOR U10539 ( .A(n8237), .B(n8238), .Z(n8057) );
  OR U10540 ( .A(n8239), .B(n8240), .Z(n8238) );
  AND U10541 ( .A(a[82]), .B(b[2]), .Z(n8236) );
  XNOR U10542 ( .A(n8067), .B(n8241), .Z(n8063) );
  NAND U10543 ( .A(a[83]), .B(b[1]), .Z(n8241) );
  IV U10544 ( .A(n8061), .Z(n8067) );
  ANDN U10545 ( .B(n5137), .A(n5139), .Z(n8061) );
  NAND U10546 ( .A(a[83]), .B(b[0]), .Z(n5139) );
  XOR U10547 ( .A(n8239), .B(n8240), .Z(n5137) );
  XOR U10548 ( .A(n8243), .B(n8234), .Z(n8242) );
  XOR U10549 ( .A(n8229), .B(n8233), .Z(n8244) );
  XOR U10550 ( .A(n8224), .B(n8228), .Z(n8245) );
  XOR U10551 ( .A(n8219), .B(n8223), .Z(n8246) );
  XOR U10552 ( .A(n8214), .B(n8218), .Z(n8247) );
  XOR U10553 ( .A(n8209), .B(n8213), .Z(n8248) );
  XOR U10554 ( .A(n8204), .B(n8208), .Z(n8249) );
  XOR U10555 ( .A(n8199), .B(n8203), .Z(n8250) );
  XOR U10556 ( .A(n8194), .B(n8198), .Z(n8251) );
  XOR U10557 ( .A(n8189), .B(n8193), .Z(n8252) );
  XOR U10558 ( .A(n8184), .B(n8188), .Z(n8253) );
  XOR U10559 ( .A(n8179), .B(n8183), .Z(n8254) );
  XOR U10560 ( .A(n8174), .B(n8178), .Z(n8255) );
  XOR U10561 ( .A(n8164), .B(n8173), .Z(n8256) );
  XOR U10562 ( .A(n8257), .B(n8163), .Z(n8164) );
  AND U10563 ( .A(b[15]), .B(a[68]), .Z(n8257) );
  XNOR U10564 ( .A(n8163), .B(n8169), .Z(n8258) );
  XNOR U10565 ( .A(n8168), .B(n8160), .Z(n8259) );
  XNOR U10566 ( .A(n8159), .B(n8155), .Z(n8260) );
  XNOR U10567 ( .A(n8154), .B(n8150), .Z(n8261) );
  XNOR U10568 ( .A(n8149), .B(n8145), .Z(n8262) );
  XNOR U10569 ( .A(n8144), .B(n8140), .Z(n8263) );
  XNOR U10570 ( .A(n8139), .B(n8135), .Z(n8264) );
  XNOR U10571 ( .A(n8134), .B(n8130), .Z(n8265) );
  XNOR U10572 ( .A(n8129), .B(n8125), .Z(n8266) );
  XNOR U10573 ( .A(n8124), .B(n8120), .Z(n8267) );
  XNOR U10574 ( .A(n8119), .B(n8115), .Z(n8268) );
  XNOR U10575 ( .A(n8114), .B(n8110), .Z(n8269) );
  XOR U10576 ( .A(n8109), .B(n8106), .Z(n8270) );
  XOR U10577 ( .A(n8271), .B(n8272), .Z(n8106) );
  XOR U10578 ( .A(n8104), .B(n8273), .Z(n8272) );
  XOR U10579 ( .A(n8274), .B(n8275), .Z(n8273) );
  XOR U10580 ( .A(n8276), .B(n8277), .Z(n8275) );
  NAND U10581 ( .A(a[53]), .B(b[30]), .Z(n8277) );
  AND U10582 ( .A(a[52]), .B(b[31]), .Z(n8276) );
  XOR U10583 ( .A(n8278), .B(n8274), .Z(n8271) );
  XOR U10584 ( .A(n8279), .B(n8280), .Z(n8274) );
  ANDN U10585 ( .B(n8281), .A(n8282), .Z(n8279) );
  AND U10586 ( .A(a[54]), .B(b[29]), .Z(n8278) );
  XOR U10587 ( .A(n8283), .B(n8104), .Z(n8105) );
  XOR U10588 ( .A(n8284), .B(n8285), .Z(n8104) );
  AND U10589 ( .A(n8286), .B(n8287), .Z(n8284) );
  AND U10590 ( .A(a[55]), .B(b[28]), .Z(n8283) );
  XOR U10591 ( .A(n8288), .B(n8109), .Z(n8111) );
  XOR U10592 ( .A(n8289), .B(n8290), .Z(n8109) );
  AND U10593 ( .A(n8291), .B(n8292), .Z(n8289) );
  AND U10594 ( .A(a[56]), .B(b[27]), .Z(n8288) );
  XOR U10595 ( .A(n8293), .B(n8114), .Z(n8116) );
  XOR U10596 ( .A(n8294), .B(n8295), .Z(n8114) );
  AND U10597 ( .A(n8296), .B(n8297), .Z(n8294) );
  AND U10598 ( .A(a[57]), .B(b[26]), .Z(n8293) );
  XOR U10599 ( .A(n8298), .B(n8119), .Z(n8121) );
  XOR U10600 ( .A(n8299), .B(n8300), .Z(n8119) );
  AND U10601 ( .A(n8301), .B(n8302), .Z(n8299) );
  AND U10602 ( .A(a[58]), .B(b[25]), .Z(n8298) );
  XOR U10603 ( .A(n8303), .B(n8124), .Z(n8126) );
  XOR U10604 ( .A(n8304), .B(n8305), .Z(n8124) );
  AND U10605 ( .A(n8306), .B(n8307), .Z(n8304) );
  AND U10606 ( .A(a[59]), .B(b[24]), .Z(n8303) );
  XOR U10607 ( .A(n8308), .B(n8129), .Z(n8131) );
  XOR U10608 ( .A(n8309), .B(n8310), .Z(n8129) );
  AND U10609 ( .A(n8311), .B(n8312), .Z(n8309) );
  AND U10610 ( .A(a[60]), .B(b[23]), .Z(n8308) );
  XOR U10611 ( .A(n8313), .B(n8134), .Z(n8136) );
  XOR U10612 ( .A(n8314), .B(n8315), .Z(n8134) );
  AND U10613 ( .A(n8316), .B(n8317), .Z(n8314) );
  AND U10614 ( .A(a[61]), .B(b[22]), .Z(n8313) );
  XOR U10615 ( .A(n8318), .B(n8139), .Z(n8141) );
  XOR U10616 ( .A(n8319), .B(n8320), .Z(n8139) );
  AND U10617 ( .A(n8321), .B(n8322), .Z(n8319) );
  AND U10618 ( .A(a[62]), .B(b[21]), .Z(n8318) );
  XOR U10619 ( .A(n8323), .B(n8144), .Z(n8146) );
  XOR U10620 ( .A(n8324), .B(n8325), .Z(n8144) );
  AND U10621 ( .A(n8326), .B(n8327), .Z(n8324) );
  AND U10622 ( .A(a[63]), .B(b[20]), .Z(n8323) );
  XOR U10623 ( .A(n8328), .B(n8149), .Z(n8151) );
  XOR U10624 ( .A(n8329), .B(n8330), .Z(n8149) );
  AND U10625 ( .A(n8331), .B(n8332), .Z(n8329) );
  AND U10626 ( .A(a[64]), .B(b[19]), .Z(n8328) );
  XOR U10627 ( .A(n8333), .B(n8154), .Z(n8156) );
  XOR U10628 ( .A(n8334), .B(n8335), .Z(n8154) );
  AND U10629 ( .A(n8336), .B(n8337), .Z(n8334) );
  AND U10630 ( .A(a[65]), .B(b[18]), .Z(n8333) );
  XOR U10631 ( .A(n8338), .B(n8159), .Z(n8161) );
  XOR U10632 ( .A(n8339), .B(n8340), .Z(n8159) );
  AND U10633 ( .A(n8341), .B(n8342), .Z(n8339) );
  AND U10634 ( .A(a[66]), .B(b[17]), .Z(n8338) );
  XOR U10635 ( .A(n8343), .B(n8344), .Z(n8163) );
  AND U10636 ( .A(n8345), .B(n8346), .Z(n8343) );
  XOR U10637 ( .A(n8347), .B(n8168), .Z(n8170) );
  XOR U10638 ( .A(n8348), .B(n8349), .Z(n8168) );
  AND U10639 ( .A(n8350), .B(n8351), .Z(n8348) );
  AND U10640 ( .A(a[67]), .B(b[16]), .Z(n8347) );
  XOR U10641 ( .A(n8353), .B(n8354), .Z(n8173) );
  AND U10642 ( .A(n8355), .B(n8356), .Z(n8353) );
  AND U10643 ( .A(a[69]), .B(b[14]), .Z(n8352) );
  XOR U10644 ( .A(n8358), .B(n8359), .Z(n8178) );
  AND U10645 ( .A(n8360), .B(n8361), .Z(n8358) );
  AND U10646 ( .A(a[70]), .B(b[13]), .Z(n8357) );
  XOR U10647 ( .A(n8363), .B(n8364), .Z(n8183) );
  AND U10648 ( .A(n8365), .B(n8366), .Z(n8363) );
  AND U10649 ( .A(a[71]), .B(b[12]), .Z(n8362) );
  XOR U10650 ( .A(n8368), .B(n8369), .Z(n8188) );
  AND U10651 ( .A(n8370), .B(n8371), .Z(n8368) );
  AND U10652 ( .A(a[72]), .B(b[11]), .Z(n8367) );
  XOR U10653 ( .A(n8373), .B(n8374), .Z(n8193) );
  AND U10654 ( .A(n8375), .B(n8376), .Z(n8373) );
  AND U10655 ( .A(a[73]), .B(b[10]), .Z(n8372) );
  XOR U10656 ( .A(n8378), .B(n8379), .Z(n8198) );
  AND U10657 ( .A(n8380), .B(n8381), .Z(n8378) );
  AND U10658 ( .A(a[74]), .B(b[9]), .Z(n8377) );
  XOR U10659 ( .A(n8383), .B(n8384), .Z(n8203) );
  AND U10660 ( .A(n8385), .B(n8386), .Z(n8383) );
  AND U10661 ( .A(a[75]), .B(b[8]), .Z(n8382) );
  XOR U10662 ( .A(n8388), .B(n8389), .Z(n8208) );
  AND U10663 ( .A(n8390), .B(n8391), .Z(n8388) );
  AND U10664 ( .A(a[76]), .B(b[7]), .Z(n8387) );
  XOR U10665 ( .A(n8393), .B(n8394), .Z(n8213) );
  AND U10666 ( .A(n8395), .B(n8396), .Z(n8393) );
  AND U10667 ( .A(a[77]), .B(b[6]), .Z(n8392) );
  XOR U10668 ( .A(n8398), .B(n8399), .Z(n8218) );
  AND U10669 ( .A(n8400), .B(n8401), .Z(n8398) );
  AND U10670 ( .A(a[78]), .B(b[5]), .Z(n8397) );
  XOR U10671 ( .A(n8403), .B(n8404), .Z(n8223) );
  AND U10672 ( .A(n8405), .B(n8406), .Z(n8403) );
  AND U10673 ( .A(a[79]), .B(b[4]), .Z(n8402) );
  XOR U10674 ( .A(n8408), .B(n8409), .Z(n8228) );
  AND U10675 ( .A(n8410), .B(n8411), .Z(n8408) );
  AND U10676 ( .A(a[80]), .B(b[3]), .Z(n8407) );
  XOR U10677 ( .A(n8413), .B(n8414), .Z(n8233) );
  OR U10678 ( .A(n8415), .B(n8416), .Z(n8414) );
  AND U10679 ( .A(a[81]), .B(b[2]), .Z(n8412) );
  XNOR U10680 ( .A(n8243), .B(n8417), .Z(n8239) );
  NAND U10681 ( .A(a[82]), .B(b[1]), .Z(n8417) );
  IV U10682 ( .A(n8237), .Z(n8243) );
  ANDN U10683 ( .B(n5142), .A(n5144), .Z(n8237) );
  NAND U10684 ( .A(a[82]), .B(b[0]), .Z(n5144) );
  XOR U10685 ( .A(n8415), .B(n8416), .Z(n5142) );
  XOR U10686 ( .A(n8419), .B(n8410), .Z(n8418) );
  XOR U10687 ( .A(n8405), .B(n8409), .Z(n8420) );
  XOR U10688 ( .A(n8400), .B(n8404), .Z(n8421) );
  XOR U10689 ( .A(n8395), .B(n8399), .Z(n8422) );
  XOR U10690 ( .A(n8390), .B(n8394), .Z(n8423) );
  XOR U10691 ( .A(n8385), .B(n8389), .Z(n8424) );
  XOR U10692 ( .A(n8380), .B(n8384), .Z(n8425) );
  XOR U10693 ( .A(n8375), .B(n8379), .Z(n8426) );
  XOR U10694 ( .A(n8370), .B(n8374), .Z(n8427) );
  XOR U10695 ( .A(n8365), .B(n8369), .Z(n8428) );
  XOR U10696 ( .A(n8360), .B(n8364), .Z(n8429) );
  XOR U10697 ( .A(n8355), .B(n8359), .Z(n8430) );
  XOR U10698 ( .A(n8345), .B(n8354), .Z(n8431) );
  XOR U10699 ( .A(n8432), .B(n8344), .Z(n8345) );
  AND U10700 ( .A(b[14]), .B(a[68]), .Z(n8432) );
  XNOR U10701 ( .A(n8344), .B(n8350), .Z(n8433) );
  XNOR U10702 ( .A(n8349), .B(n8341), .Z(n8434) );
  XNOR U10703 ( .A(n8340), .B(n8336), .Z(n8435) );
  XNOR U10704 ( .A(n8335), .B(n8331), .Z(n8436) );
  XNOR U10705 ( .A(n8330), .B(n8326), .Z(n8437) );
  XNOR U10706 ( .A(n8325), .B(n8321), .Z(n8438) );
  XNOR U10707 ( .A(n8320), .B(n8316), .Z(n8439) );
  XNOR U10708 ( .A(n8315), .B(n8311), .Z(n8440) );
  XNOR U10709 ( .A(n8310), .B(n8306), .Z(n8441) );
  XNOR U10710 ( .A(n8305), .B(n8301), .Z(n8442) );
  XNOR U10711 ( .A(n8300), .B(n8296), .Z(n8443) );
  XNOR U10712 ( .A(n8295), .B(n8291), .Z(n8444) );
  XNOR U10713 ( .A(n8290), .B(n8286), .Z(n8445) );
  XOR U10714 ( .A(n8285), .B(n8282), .Z(n8446) );
  XOR U10715 ( .A(n8447), .B(n8448), .Z(n8282) );
  XOR U10716 ( .A(n8280), .B(n8449), .Z(n8448) );
  XOR U10717 ( .A(n8450), .B(n8451), .Z(n8449) );
  XOR U10718 ( .A(n8452), .B(n8453), .Z(n8451) );
  NAND U10719 ( .A(a[52]), .B(b[30]), .Z(n8453) );
  AND U10720 ( .A(a[51]), .B(b[31]), .Z(n8452) );
  XOR U10721 ( .A(n8454), .B(n8450), .Z(n8447) );
  XOR U10722 ( .A(n8455), .B(n8456), .Z(n8450) );
  ANDN U10723 ( .B(n8457), .A(n8458), .Z(n8455) );
  AND U10724 ( .A(a[53]), .B(b[29]), .Z(n8454) );
  XOR U10725 ( .A(n8459), .B(n8280), .Z(n8281) );
  XOR U10726 ( .A(n8460), .B(n8461), .Z(n8280) );
  AND U10727 ( .A(n8462), .B(n8463), .Z(n8460) );
  AND U10728 ( .A(a[54]), .B(b[28]), .Z(n8459) );
  XOR U10729 ( .A(n8464), .B(n8285), .Z(n8287) );
  XOR U10730 ( .A(n8465), .B(n8466), .Z(n8285) );
  AND U10731 ( .A(n8467), .B(n8468), .Z(n8465) );
  AND U10732 ( .A(a[55]), .B(b[27]), .Z(n8464) );
  XOR U10733 ( .A(n8469), .B(n8290), .Z(n8292) );
  XOR U10734 ( .A(n8470), .B(n8471), .Z(n8290) );
  AND U10735 ( .A(n8472), .B(n8473), .Z(n8470) );
  AND U10736 ( .A(a[56]), .B(b[26]), .Z(n8469) );
  XOR U10737 ( .A(n8474), .B(n8295), .Z(n8297) );
  XOR U10738 ( .A(n8475), .B(n8476), .Z(n8295) );
  AND U10739 ( .A(n8477), .B(n8478), .Z(n8475) );
  AND U10740 ( .A(a[57]), .B(b[25]), .Z(n8474) );
  XOR U10741 ( .A(n8479), .B(n8300), .Z(n8302) );
  XOR U10742 ( .A(n8480), .B(n8481), .Z(n8300) );
  AND U10743 ( .A(n8482), .B(n8483), .Z(n8480) );
  AND U10744 ( .A(a[58]), .B(b[24]), .Z(n8479) );
  XOR U10745 ( .A(n8484), .B(n8305), .Z(n8307) );
  XOR U10746 ( .A(n8485), .B(n8486), .Z(n8305) );
  AND U10747 ( .A(n8487), .B(n8488), .Z(n8485) );
  AND U10748 ( .A(a[59]), .B(b[23]), .Z(n8484) );
  XOR U10749 ( .A(n8489), .B(n8310), .Z(n8312) );
  XOR U10750 ( .A(n8490), .B(n8491), .Z(n8310) );
  AND U10751 ( .A(n8492), .B(n8493), .Z(n8490) );
  AND U10752 ( .A(a[60]), .B(b[22]), .Z(n8489) );
  XOR U10753 ( .A(n8494), .B(n8315), .Z(n8317) );
  XOR U10754 ( .A(n8495), .B(n8496), .Z(n8315) );
  AND U10755 ( .A(n8497), .B(n8498), .Z(n8495) );
  AND U10756 ( .A(a[61]), .B(b[21]), .Z(n8494) );
  XOR U10757 ( .A(n8499), .B(n8320), .Z(n8322) );
  XOR U10758 ( .A(n8500), .B(n8501), .Z(n8320) );
  AND U10759 ( .A(n8502), .B(n8503), .Z(n8500) );
  AND U10760 ( .A(a[62]), .B(b[20]), .Z(n8499) );
  XOR U10761 ( .A(n8504), .B(n8325), .Z(n8327) );
  XOR U10762 ( .A(n8505), .B(n8506), .Z(n8325) );
  AND U10763 ( .A(n8507), .B(n8508), .Z(n8505) );
  AND U10764 ( .A(a[63]), .B(b[19]), .Z(n8504) );
  XOR U10765 ( .A(n8509), .B(n8330), .Z(n8332) );
  XOR U10766 ( .A(n8510), .B(n8511), .Z(n8330) );
  AND U10767 ( .A(n8512), .B(n8513), .Z(n8510) );
  AND U10768 ( .A(a[64]), .B(b[18]), .Z(n8509) );
  XOR U10769 ( .A(n8514), .B(n8335), .Z(n8337) );
  XOR U10770 ( .A(n8515), .B(n8516), .Z(n8335) );
  AND U10771 ( .A(n8517), .B(n8518), .Z(n8515) );
  AND U10772 ( .A(a[65]), .B(b[17]), .Z(n8514) );
  XOR U10773 ( .A(n8519), .B(n8340), .Z(n8342) );
  XOR U10774 ( .A(n8520), .B(n8521), .Z(n8340) );
  AND U10775 ( .A(n8522), .B(n8523), .Z(n8520) );
  AND U10776 ( .A(a[66]), .B(b[16]), .Z(n8519) );
  XOR U10777 ( .A(n8524), .B(n8525), .Z(n8344) );
  AND U10778 ( .A(n8526), .B(n8527), .Z(n8524) );
  XOR U10779 ( .A(n8528), .B(n8349), .Z(n8351) );
  XOR U10780 ( .A(n8529), .B(n8530), .Z(n8349) );
  AND U10781 ( .A(n8531), .B(n8532), .Z(n8529) );
  AND U10782 ( .A(a[67]), .B(b[15]), .Z(n8528) );
  XOR U10783 ( .A(n8534), .B(n8535), .Z(n8354) );
  AND U10784 ( .A(n8536), .B(n8537), .Z(n8534) );
  AND U10785 ( .A(a[69]), .B(b[13]), .Z(n8533) );
  XOR U10786 ( .A(n8539), .B(n8540), .Z(n8359) );
  AND U10787 ( .A(n8541), .B(n8542), .Z(n8539) );
  AND U10788 ( .A(a[70]), .B(b[12]), .Z(n8538) );
  XOR U10789 ( .A(n8544), .B(n8545), .Z(n8364) );
  AND U10790 ( .A(n8546), .B(n8547), .Z(n8544) );
  AND U10791 ( .A(a[71]), .B(b[11]), .Z(n8543) );
  XOR U10792 ( .A(n8549), .B(n8550), .Z(n8369) );
  AND U10793 ( .A(n8551), .B(n8552), .Z(n8549) );
  AND U10794 ( .A(a[72]), .B(b[10]), .Z(n8548) );
  XOR U10795 ( .A(n8554), .B(n8555), .Z(n8374) );
  AND U10796 ( .A(n8556), .B(n8557), .Z(n8554) );
  AND U10797 ( .A(a[73]), .B(b[9]), .Z(n8553) );
  XOR U10798 ( .A(n8559), .B(n8560), .Z(n8379) );
  AND U10799 ( .A(n8561), .B(n8562), .Z(n8559) );
  AND U10800 ( .A(a[74]), .B(b[8]), .Z(n8558) );
  XOR U10801 ( .A(n8564), .B(n8565), .Z(n8384) );
  AND U10802 ( .A(n8566), .B(n8567), .Z(n8564) );
  AND U10803 ( .A(a[75]), .B(b[7]), .Z(n8563) );
  XOR U10804 ( .A(n8569), .B(n8570), .Z(n8389) );
  AND U10805 ( .A(n8571), .B(n8572), .Z(n8569) );
  AND U10806 ( .A(a[76]), .B(b[6]), .Z(n8568) );
  XOR U10807 ( .A(n8574), .B(n8575), .Z(n8394) );
  AND U10808 ( .A(n8576), .B(n8577), .Z(n8574) );
  AND U10809 ( .A(a[77]), .B(b[5]), .Z(n8573) );
  XOR U10810 ( .A(n8579), .B(n8580), .Z(n8399) );
  AND U10811 ( .A(n8581), .B(n8582), .Z(n8579) );
  AND U10812 ( .A(a[78]), .B(b[4]), .Z(n8578) );
  XOR U10813 ( .A(n8584), .B(n8585), .Z(n8404) );
  AND U10814 ( .A(n8586), .B(n8587), .Z(n8584) );
  AND U10815 ( .A(a[79]), .B(b[3]), .Z(n8583) );
  XOR U10816 ( .A(n8589), .B(n8590), .Z(n8409) );
  OR U10817 ( .A(n8591), .B(n8592), .Z(n8590) );
  AND U10818 ( .A(a[80]), .B(b[2]), .Z(n8588) );
  XNOR U10819 ( .A(n8419), .B(n8593), .Z(n8415) );
  NAND U10820 ( .A(a[81]), .B(b[1]), .Z(n8593) );
  IV U10821 ( .A(n8413), .Z(n8419) );
  ANDN U10822 ( .B(n5147), .A(n5149), .Z(n8413) );
  NAND U10823 ( .A(a[81]), .B(b[0]), .Z(n5149) );
  XOR U10824 ( .A(n8591), .B(n8592), .Z(n5147) );
  XOR U10825 ( .A(n8595), .B(n8586), .Z(n8594) );
  XOR U10826 ( .A(n8581), .B(n8585), .Z(n8596) );
  XOR U10827 ( .A(n8576), .B(n8580), .Z(n8597) );
  XOR U10828 ( .A(n8571), .B(n8575), .Z(n8598) );
  XOR U10829 ( .A(n8566), .B(n8570), .Z(n8599) );
  XOR U10830 ( .A(n8561), .B(n8565), .Z(n8600) );
  XOR U10831 ( .A(n8556), .B(n8560), .Z(n8601) );
  XOR U10832 ( .A(n8551), .B(n8555), .Z(n8602) );
  XOR U10833 ( .A(n8546), .B(n8550), .Z(n8603) );
  XOR U10834 ( .A(n8541), .B(n8545), .Z(n8604) );
  XOR U10835 ( .A(n8536), .B(n8540), .Z(n8605) );
  XOR U10836 ( .A(n8526), .B(n8535), .Z(n8606) );
  XOR U10837 ( .A(n8607), .B(n8525), .Z(n8526) );
  AND U10838 ( .A(b[13]), .B(a[68]), .Z(n8607) );
  XNOR U10839 ( .A(n8525), .B(n8531), .Z(n8608) );
  XNOR U10840 ( .A(n8530), .B(n8522), .Z(n8609) );
  XNOR U10841 ( .A(n8521), .B(n8517), .Z(n8610) );
  XNOR U10842 ( .A(n8516), .B(n8512), .Z(n8611) );
  XNOR U10843 ( .A(n8511), .B(n8507), .Z(n8612) );
  XNOR U10844 ( .A(n8506), .B(n8502), .Z(n8613) );
  XNOR U10845 ( .A(n8501), .B(n8497), .Z(n8614) );
  XNOR U10846 ( .A(n8496), .B(n8492), .Z(n8615) );
  XNOR U10847 ( .A(n8491), .B(n8487), .Z(n8616) );
  XNOR U10848 ( .A(n8486), .B(n8482), .Z(n8617) );
  XNOR U10849 ( .A(n8481), .B(n8477), .Z(n8618) );
  XNOR U10850 ( .A(n8476), .B(n8472), .Z(n8619) );
  XNOR U10851 ( .A(n8471), .B(n8467), .Z(n8620) );
  XNOR U10852 ( .A(n8466), .B(n8462), .Z(n8621) );
  XOR U10853 ( .A(n8461), .B(n8458), .Z(n8622) );
  XOR U10854 ( .A(n8623), .B(n8624), .Z(n8458) );
  XOR U10855 ( .A(n8456), .B(n8625), .Z(n8624) );
  XOR U10856 ( .A(n8626), .B(n8627), .Z(n8625) );
  XOR U10857 ( .A(n8628), .B(n8629), .Z(n8627) );
  NAND U10858 ( .A(a[51]), .B(b[30]), .Z(n8629) );
  AND U10859 ( .A(a[50]), .B(b[31]), .Z(n8628) );
  XOR U10860 ( .A(n8630), .B(n8626), .Z(n8623) );
  XOR U10861 ( .A(n8631), .B(n8632), .Z(n8626) );
  ANDN U10862 ( .B(n8633), .A(n8634), .Z(n8631) );
  AND U10863 ( .A(a[52]), .B(b[29]), .Z(n8630) );
  XOR U10864 ( .A(n8635), .B(n8456), .Z(n8457) );
  XOR U10865 ( .A(n8636), .B(n8637), .Z(n8456) );
  AND U10866 ( .A(n8638), .B(n8639), .Z(n8636) );
  AND U10867 ( .A(a[53]), .B(b[28]), .Z(n8635) );
  XOR U10868 ( .A(n8640), .B(n8461), .Z(n8463) );
  XOR U10869 ( .A(n8641), .B(n8642), .Z(n8461) );
  AND U10870 ( .A(n8643), .B(n8644), .Z(n8641) );
  AND U10871 ( .A(a[54]), .B(b[27]), .Z(n8640) );
  XOR U10872 ( .A(n8645), .B(n8466), .Z(n8468) );
  XOR U10873 ( .A(n8646), .B(n8647), .Z(n8466) );
  AND U10874 ( .A(n8648), .B(n8649), .Z(n8646) );
  AND U10875 ( .A(a[55]), .B(b[26]), .Z(n8645) );
  XOR U10876 ( .A(n8650), .B(n8471), .Z(n8473) );
  XOR U10877 ( .A(n8651), .B(n8652), .Z(n8471) );
  AND U10878 ( .A(n8653), .B(n8654), .Z(n8651) );
  AND U10879 ( .A(a[56]), .B(b[25]), .Z(n8650) );
  XOR U10880 ( .A(n8655), .B(n8476), .Z(n8478) );
  XOR U10881 ( .A(n8656), .B(n8657), .Z(n8476) );
  AND U10882 ( .A(n8658), .B(n8659), .Z(n8656) );
  AND U10883 ( .A(a[57]), .B(b[24]), .Z(n8655) );
  XOR U10884 ( .A(n8660), .B(n8481), .Z(n8483) );
  XOR U10885 ( .A(n8661), .B(n8662), .Z(n8481) );
  AND U10886 ( .A(n8663), .B(n8664), .Z(n8661) );
  AND U10887 ( .A(a[58]), .B(b[23]), .Z(n8660) );
  XOR U10888 ( .A(n8665), .B(n8486), .Z(n8488) );
  XOR U10889 ( .A(n8666), .B(n8667), .Z(n8486) );
  AND U10890 ( .A(n8668), .B(n8669), .Z(n8666) );
  AND U10891 ( .A(a[59]), .B(b[22]), .Z(n8665) );
  XOR U10892 ( .A(n8670), .B(n8491), .Z(n8493) );
  XOR U10893 ( .A(n8671), .B(n8672), .Z(n8491) );
  AND U10894 ( .A(n8673), .B(n8674), .Z(n8671) );
  AND U10895 ( .A(a[60]), .B(b[21]), .Z(n8670) );
  XOR U10896 ( .A(n8675), .B(n8496), .Z(n8498) );
  XOR U10897 ( .A(n8676), .B(n8677), .Z(n8496) );
  AND U10898 ( .A(n8678), .B(n8679), .Z(n8676) );
  AND U10899 ( .A(a[61]), .B(b[20]), .Z(n8675) );
  XOR U10900 ( .A(n8680), .B(n8501), .Z(n8503) );
  XOR U10901 ( .A(n8681), .B(n8682), .Z(n8501) );
  AND U10902 ( .A(n8683), .B(n8684), .Z(n8681) );
  AND U10903 ( .A(a[62]), .B(b[19]), .Z(n8680) );
  XOR U10904 ( .A(n8685), .B(n8506), .Z(n8508) );
  XOR U10905 ( .A(n8686), .B(n8687), .Z(n8506) );
  AND U10906 ( .A(n8688), .B(n8689), .Z(n8686) );
  AND U10907 ( .A(a[63]), .B(b[18]), .Z(n8685) );
  XOR U10908 ( .A(n8690), .B(n8511), .Z(n8513) );
  XOR U10909 ( .A(n8691), .B(n8692), .Z(n8511) );
  AND U10910 ( .A(n8693), .B(n8694), .Z(n8691) );
  AND U10911 ( .A(a[64]), .B(b[17]), .Z(n8690) );
  XOR U10912 ( .A(n8695), .B(n8516), .Z(n8518) );
  XOR U10913 ( .A(n8696), .B(n8697), .Z(n8516) );
  AND U10914 ( .A(n8698), .B(n8699), .Z(n8696) );
  AND U10915 ( .A(a[65]), .B(b[16]), .Z(n8695) );
  XOR U10916 ( .A(n8700), .B(n8521), .Z(n8523) );
  XOR U10917 ( .A(n8701), .B(n8702), .Z(n8521) );
  AND U10918 ( .A(n8703), .B(n8704), .Z(n8701) );
  AND U10919 ( .A(a[66]), .B(b[15]), .Z(n8700) );
  XOR U10920 ( .A(n8705), .B(n8706), .Z(n8525) );
  AND U10921 ( .A(n8707), .B(n8708), .Z(n8705) );
  XOR U10922 ( .A(n8709), .B(n8530), .Z(n8532) );
  XOR U10923 ( .A(n8710), .B(n8711), .Z(n8530) );
  AND U10924 ( .A(n8712), .B(n8713), .Z(n8710) );
  AND U10925 ( .A(a[67]), .B(b[14]), .Z(n8709) );
  XOR U10926 ( .A(n8715), .B(n8716), .Z(n8535) );
  AND U10927 ( .A(n8717), .B(n8718), .Z(n8715) );
  AND U10928 ( .A(a[69]), .B(b[12]), .Z(n8714) );
  XOR U10929 ( .A(n8720), .B(n8721), .Z(n8540) );
  AND U10930 ( .A(n8722), .B(n8723), .Z(n8720) );
  AND U10931 ( .A(a[70]), .B(b[11]), .Z(n8719) );
  XOR U10932 ( .A(n8725), .B(n8726), .Z(n8545) );
  AND U10933 ( .A(n8727), .B(n8728), .Z(n8725) );
  AND U10934 ( .A(a[71]), .B(b[10]), .Z(n8724) );
  XOR U10935 ( .A(n8730), .B(n8731), .Z(n8550) );
  AND U10936 ( .A(n8732), .B(n8733), .Z(n8730) );
  AND U10937 ( .A(a[72]), .B(b[9]), .Z(n8729) );
  XOR U10938 ( .A(n8735), .B(n8736), .Z(n8555) );
  AND U10939 ( .A(n8737), .B(n8738), .Z(n8735) );
  AND U10940 ( .A(a[73]), .B(b[8]), .Z(n8734) );
  XOR U10941 ( .A(n8740), .B(n8741), .Z(n8560) );
  AND U10942 ( .A(n8742), .B(n8743), .Z(n8740) );
  AND U10943 ( .A(a[74]), .B(b[7]), .Z(n8739) );
  XOR U10944 ( .A(n8745), .B(n8746), .Z(n8565) );
  AND U10945 ( .A(n8747), .B(n8748), .Z(n8745) );
  AND U10946 ( .A(a[75]), .B(b[6]), .Z(n8744) );
  XOR U10947 ( .A(n8750), .B(n8751), .Z(n8570) );
  AND U10948 ( .A(n8752), .B(n8753), .Z(n8750) );
  AND U10949 ( .A(a[76]), .B(b[5]), .Z(n8749) );
  XOR U10950 ( .A(n8755), .B(n8756), .Z(n8575) );
  AND U10951 ( .A(n8757), .B(n8758), .Z(n8755) );
  AND U10952 ( .A(a[77]), .B(b[4]), .Z(n8754) );
  XOR U10953 ( .A(n8760), .B(n8761), .Z(n8580) );
  AND U10954 ( .A(n8762), .B(n8763), .Z(n8760) );
  AND U10955 ( .A(a[78]), .B(b[3]), .Z(n8759) );
  XOR U10956 ( .A(n8765), .B(n8766), .Z(n8585) );
  OR U10957 ( .A(n8767), .B(n8768), .Z(n8766) );
  AND U10958 ( .A(a[79]), .B(b[2]), .Z(n8764) );
  XNOR U10959 ( .A(n8595), .B(n8769), .Z(n8591) );
  NAND U10960 ( .A(a[80]), .B(b[1]), .Z(n8769) );
  IV U10961 ( .A(n8589), .Z(n8595) );
  ANDN U10962 ( .B(n5152), .A(n5154), .Z(n8589) );
  NAND U10963 ( .A(a[80]), .B(b[0]), .Z(n5154) );
  XOR U10964 ( .A(n8767), .B(n8768), .Z(n5152) );
  XOR U10965 ( .A(n8771), .B(n8762), .Z(n8770) );
  XOR U10966 ( .A(n8757), .B(n8761), .Z(n8772) );
  XOR U10967 ( .A(n8752), .B(n8756), .Z(n8773) );
  XOR U10968 ( .A(n8747), .B(n8751), .Z(n8774) );
  XOR U10969 ( .A(n8742), .B(n8746), .Z(n8775) );
  XOR U10970 ( .A(n8737), .B(n8741), .Z(n8776) );
  XOR U10971 ( .A(n8732), .B(n8736), .Z(n8777) );
  XOR U10972 ( .A(n8727), .B(n8731), .Z(n8778) );
  XOR U10973 ( .A(n8722), .B(n8726), .Z(n8779) );
  XOR U10974 ( .A(n8717), .B(n8721), .Z(n8780) );
  XOR U10975 ( .A(n8707), .B(n8716), .Z(n8781) );
  XOR U10976 ( .A(n8782), .B(n8706), .Z(n8707) );
  AND U10977 ( .A(b[12]), .B(a[68]), .Z(n8782) );
  XNOR U10978 ( .A(n8706), .B(n8712), .Z(n8783) );
  XNOR U10979 ( .A(n8711), .B(n8703), .Z(n8784) );
  XNOR U10980 ( .A(n8702), .B(n8698), .Z(n8785) );
  XNOR U10981 ( .A(n8697), .B(n8693), .Z(n8786) );
  XNOR U10982 ( .A(n8692), .B(n8688), .Z(n8787) );
  XNOR U10983 ( .A(n8687), .B(n8683), .Z(n8788) );
  XNOR U10984 ( .A(n8682), .B(n8678), .Z(n8789) );
  XNOR U10985 ( .A(n8677), .B(n8673), .Z(n8790) );
  XNOR U10986 ( .A(n8672), .B(n8668), .Z(n8791) );
  XNOR U10987 ( .A(n8667), .B(n8663), .Z(n8792) );
  XNOR U10988 ( .A(n8662), .B(n8658), .Z(n8793) );
  XNOR U10989 ( .A(n8657), .B(n8653), .Z(n8794) );
  XNOR U10990 ( .A(n8652), .B(n8648), .Z(n8795) );
  XNOR U10991 ( .A(n8647), .B(n8643), .Z(n8796) );
  XNOR U10992 ( .A(n8642), .B(n8638), .Z(n8797) );
  XOR U10993 ( .A(n8637), .B(n8634), .Z(n8798) );
  XOR U10994 ( .A(n8799), .B(n8800), .Z(n8634) );
  XOR U10995 ( .A(n8632), .B(n8801), .Z(n8800) );
  XOR U10996 ( .A(n8802), .B(n8803), .Z(n8801) );
  XOR U10997 ( .A(n8804), .B(n8805), .Z(n8803) );
  NAND U10998 ( .A(a[50]), .B(b[30]), .Z(n8805) );
  AND U10999 ( .A(a[49]), .B(b[31]), .Z(n8804) );
  XOR U11000 ( .A(n8806), .B(n8802), .Z(n8799) );
  XOR U11001 ( .A(n8807), .B(n8808), .Z(n8802) );
  ANDN U11002 ( .B(n8809), .A(n8810), .Z(n8807) );
  AND U11003 ( .A(a[51]), .B(b[29]), .Z(n8806) );
  XOR U11004 ( .A(n8811), .B(n8632), .Z(n8633) );
  XOR U11005 ( .A(n8812), .B(n8813), .Z(n8632) );
  AND U11006 ( .A(n8814), .B(n8815), .Z(n8812) );
  AND U11007 ( .A(a[52]), .B(b[28]), .Z(n8811) );
  XOR U11008 ( .A(n8816), .B(n8637), .Z(n8639) );
  XOR U11009 ( .A(n8817), .B(n8818), .Z(n8637) );
  AND U11010 ( .A(n8819), .B(n8820), .Z(n8817) );
  AND U11011 ( .A(a[53]), .B(b[27]), .Z(n8816) );
  XOR U11012 ( .A(n8821), .B(n8642), .Z(n8644) );
  XOR U11013 ( .A(n8822), .B(n8823), .Z(n8642) );
  AND U11014 ( .A(n8824), .B(n8825), .Z(n8822) );
  AND U11015 ( .A(a[54]), .B(b[26]), .Z(n8821) );
  XOR U11016 ( .A(n8826), .B(n8647), .Z(n8649) );
  XOR U11017 ( .A(n8827), .B(n8828), .Z(n8647) );
  AND U11018 ( .A(n8829), .B(n8830), .Z(n8827) );
  AND U11019 ( .A(a[55]), .B(b[25]), .Z(n8826) );
  XOR U11020 ( .A(n8831), .B(n8652), .Z(n8654) );
  XOR U11021 ( .A(n8832), .B(n8833), .Z(n8652) );
  AND U11022 ( .A(n8834), .B(n8835), .Z(n8832) );
  AND U11023 ( .A(a[56]), .B(b[24]), .Z(n8831) );
  XOR U11024 ( .A(n8836), .B(n8657), .Z(n8659) );
  XOR U11025 ( .A(n8837), .B(n8838), .Z(n8657) );
  AND U11026 ( .A(n8839), .B(n8840), .Z(n8837) );
  AND U11027 ( .A(a[57]), .B(b[23]), .Z(n8836) );
  XOR U11028 ( .A(n8841), .B(n8662), .Z(n8664) );
  XOR U11029 ( .A(n8842), .B(n8843), .Z(n8662) );
  AND U11030 ( .A(n8844), .B(n8845), .Z(n8842) );
  AND U11031 ( .A(a[58]), .B(b[22]), .Z(n8841) );
  XOR U11032 ( .A(n8846), .B(n8667), .Z(n8669) );
  XOR U11033 ( .A(n8847), .B(n8848), .Z(n8667) );
  AND U11034 ( .A(n8849), .B(n8850), .Z(n8847) );
  AND U11035 ( .A(a[59]), .B(b[21]), .Z(n8846) );
  XOR U11036 ( .A(n8851), .B(n8672), .Z(n8674) );
  XOR U11037 ( .A(n8852), .B(n8853), .Z(n8672) );
  AND U11038 ( .A(n8854), .B(n8855), .Z(n8852) );
  AND U11039 ( .A(a[60]), .B(b[20]), .Z(n8851) );
  XOR U11040 ( .A(n8856), .B(n8677), .Z(n8679) );
  XOR U11041 ( .A(n8857), .B(n8858), .Z(n8677) );
  AND U11042 ( .A(n8859), .B(n8860), .Z(n8857) );
  AND U11043 ( .A(a[61]), .B(b[19]), .Z(n8856) );
  XOR U11044 ( .A(n8861), .B(n8682), .Z(n8684) );
  XOR U11045 ( .A(n8862), .B(n8863), .Z(n8682) );
  AND U11046 ( .A(n8864), .B(n8865), .Z(n8862) );
  AND U11047 ( .A(a[62]), .B(b[18]), .Z(n8861) );
  XOR U11048 ( .A(n8866), .B(n8687), .Z(n8689) );
  XOR U11049 ( .A(n8867), .B(n8868), .Z(n8687) );
  AND U11050 ( .A(n8869), .B(n8870), .Z(n8867) );
  AND U11051 ( .A(a[63]), .B(b[17]), .Z(n8866) );
  XOR U11052 ( .A(n8871), .B(n8692), .Z(n8694) );
  XOR U11053 ( .A(n8872), .B(n8873), .Z(n8692) );
  AND U11054 ( .A(n8874), .B(n8875), .Z(n8872) );
  AND U11055 ( .A(a[64]), .B(b[16]), .Z(n8871) );
  XOR U11056 ( .A(n8876), .B(n8697), .Z(n8699) );
  XOR U11057 ( .A(n8877), .B(n8878), .Z(n8697) );
  AND U11058 ( .A(n8879), .B(n8880), .Z(n8877) );
  AND U11059 ( .A(a[65]), .B(b[15]), .Z(n8876) );
  XOR U11060 ( .A(n8881), .B(n8702), .Z(n8704) );
  XOR U11061 ( .A(n8882), .B(n8883), .Z(n8702) );
  AND U11062 ( .A(n8884), .B(n8885), .Z(n8882) );
  AND U11063 ( .A(a[66]), .B(b[14]), .Z(n8881) );
  XOR U11064 ( .A(n8886), .B(n8887), .Z(n8706) );
  AND U11065 ( .A(n8888), .B(n8889), .Z(n8886) );
  XOR U11066 ( .A(n8890), .B(n8711), .Z(n8713) );
  XOR U11067 ( .A(n8891), .B(n8892), .Z(n8711) );
  AND U11068 ( .A(n8893), .B(n8894), .Z(n8891) );
  AND U11069 ( .A(a[67]), .B(b[13]), .Z(n8890) );
  XOR U11070 ( .A(n8896), .B(n8897), .Z(n8716) );
  AND U11071 ( .A(n8898), .B(n8899), .Z(n8896) );
  AND U11072 ( .A(a[69]), .B(b[11]), .Z(n8895) );
  XOR U11073 ( .A(n8901), .B(n8902), .Z(n8721) );
  AND U11074 ( .A(n8903), .B(n8904), .Z(n8901) );
  AND U11075 ( .A(a[70]), .B(b[10]), .Z(n8900) );
  XOR U11076 ( .A(n8906), .B(n8907), .Z(n8726) );
  AND U11077 ( .A(n8908), .B(n8909), .Z(n8906) );
  AND U11078 ( .A(a[71]), .B(b[9]), .Z(n8905) );
  XOR U11079 ( .A(n8911), .B(n8912), .Z(n8731) );
  AND U11080 ( .A(n8913), .B(n8914), .Z(n8911) );
  AND U11081 ( .A(a[72]), .B(b[8]), .Z(n8910) );
  XOR U11082 ( .A(n8916), .B(n8917), .Z(n8736) );
  AND U11083 ( .A(n8918), .B(n8919), .Z(n8916) );
  AND U11084 ( .A(a[73]), .B(b[7]), .Z(n8915) );
  XOR U11085 ( .A(n8921), .B(n8922), .Z(n8741) );
  AND U11086 ( .A(n8923), .B(n8924), .Z(n8921) );
  AND U11087 ( .A(a[74]), .B(b[6]), .Z(n8920) );
  XOR U11088 ( .A(n8926), .B(n8927), .Z(n8746) );
  AND U11089 ( .A(n8928), .B(n8929), .Z(n8926) );
  AND U11090 ( .A(a[75]), .B(b[5]), .Z(n8925) );
  XOR U11091 ( .A(n8931), .B(n8932), .Z(n8751) );
  AND U11092 ( .A(n8933), .B(n8934), .Z(n8931) );
  AND U11093 ( .A(a[76]), .B(b[4]), .Z(n8930) );
  XOR U11094 ( .A(n8936), .B(n8937), .Z(n8756) );
  AND U11095 ( .A(n8938), .B(n8939), .Z(n8936) );
  AND U11096 ( .A(a[77]), .B(b[3]), .Z(n8935) );
  XOR U11097 ( .A(n8941), .B(n8942), .Z(n8761) );
  OR U11098 ( .A(n8943), .B(n8944), .Z(n8942) );
  AND U11099 ( .A(a[78]), .B(b[2]), .Z(n8940) );
  XNOR U11100 ( .A(n8771), .B(n8945), .Z(n8767) );
  NAND U11101 ( .A(a[79]), .B(b[1]), .Z(n8945) );
  IV U11102 ( .A(n8765), .Z(n8771) );
  ANDN U11103 ( .B(n5157), .A(n5159), .Z(n8765) );
  NAND U11104 ( .A(a[79]), .B(b[0]), .Z(n5159) );
  XOR U11105 ( .A(n8943), .B(n8944), .Z(n5157) );
  XOR U11106 ( .A(n8947), .B(n8938), .Z(n8946) );
  XOR U11107 ( .A(n8933), .B(n8937), .Z(n8948) );
  XOR U11108 ( .A(n8928), .B(n8932), .Z(n8949) );
  XOR U11109 ( .A(n8923), .B(n8927), .Z(n8950) );
  XOR U11110 ( .A(n8918), .B(n8922), .Z(n8951) );
  XOR U11111 ( .A(n8913), .B(n8917), .Z(n8952) );
  XOR U11112 ( .A(n8908), .B(n8912), .Z(n8953) );
  XOR U11113 ( .A(n8903), .B(n8907), .Z(n8954) );
  XOR U11114 ( .A(n8898), .B(n8902), .Z(n8955) );
  XOR U11115 ( .A(n8888), .B(n8897), .Z(n8956) );
  XOR U11116 ( .A(n8957), .B(n8887), .Z(n8888) );
  AND U11117 ( .A(b[11]), .B(a[68]), .Z(n8957) );
  XNOR U11118 ( .A(n8887), .B(n8893), .Z(n8958) );
  XNOR U11119 ( .A(n8892), .B(n8884), .Z(n8959) );
  XNOR U11120 ( .A(n8883), .B(n8879), .Z(n8960) );
  XNOR U11121 ( .A(n8878), .B(n8874), .Z(n8961) );
  XNOR U11122 ( .A(n8873), .B(n8869), .Z(n8962) );
  XNOR U11123 ( .A(n8868), .B(n8864), .Z(n8963) );
  XNOR U11124 ( .A(n8863), .B(n8859), .Z(n8964) );
  XNOR U11125 ( .A(n8858), .B(n8854), .Z(n8965) );
  XNOR U11126 ( .A(n8853), .B(n8849), .Z(n8966) );
  XNOR U11127 ( .A(n8848), .B(n8844), .Z(n8967) );
  XNOR U11128 ( .A(n8843), .B(n8839), .Z(n8968) );
  XNOR U11129 ( .A(n8838), .B(n8834), .Z(n8969) );
  XNOR U11130 ( .A(n8833), .B(n8829), .Z(n8970) );
  XNOR U11131 ( .A(n8828), .B(n8824), .Z(n8971) );
  XNOR U11132 ( .A(n8823), .B(n8819), .Z(n8972) );
  XNOR U11133 ( .A(n8818), .B(n8814), .Z(n8973) );
  XOR U11134 ( .A(n8813), .B(n8810), .Z(n8974) );
  XOR U11135 ( .A(n8975), .B(n8976), .Z(n8810) );
  XOR U11136 ( .A(n8808), .B(n8977), .Z(n8976) );
  XOR U11137 ( .A(n8978), .B(n8979), .Z(n8977) );
  XOR U11138 ( .A(n8980), .B(n8981), .Z(n8979) );
  NAND U11139 ( .A(a[49]), .B(b[30]), .Z(n8981) );
  AND U11140 ( .A(a[48]), .B(b[31]), .Z(n8980) );
  XOR U11141 ( .A(n8982), .B(n8978), .Z(n8975) );
  XOR U11142 ( .A(n8983), .B(n8984), .Z(n8978) );
  ANDN U11143 ( .B(n8985), .A(n8986), .Z(n8983) );
  AND U11144 ( .A(a[50]), .B(b[29]), .Z(n8982) );
  XOR U11145 ( .A(n8987), .B(n8808), .Z(n8809) );
  XOR U11146 ( .A(n8988), .B(n8989), .Z(n8808) );
  AND U11147 ( .A(n8990), .B(n8991), .Z(n8988) );
  AND U11148 ( .A(a[51]), .B(b[28]), .Z(n8987) );
  XOR U11149 ( .A(n8992), .B(n8813), .Z(n8815) );
  XOR U11150 ( .A(n8993), .B(n8994), .Z(n8813) );
  AND U11151 ( .A(n8995), .B(n8996), .Z(n8993) );
  AND U11152 ( .A(a[52]), .B(b[27]), .Z(n8992) );
  XOR U11153 ( .A(n8997), .B(n8818), .Z(n8820) );
  XOR U11154 ( .A(n8998), .B(n8999), .Z(n8818) );
  AND U11155 ( .A(n9000), .B(n9001), .Z(n8998) );
  AND U11156 ( .A(a[53]), .B(b[26]), .Z(n8997) );
  XOR U11157 ( .A(n9002), .B(n8823), .Z(n8825) );
  XOR U11158 ( .A(n9003), .B(n9004), .Z(n8823) );
  AND U11159 ( .A(n9005), .B(n9006), .Z(n9003) );
  AND U11160 ( .A(a[54]), .B(b[25]), .Z(n9002) );
  XOR U11161 ( .A(n9007), .B(n8828), .Z(n8830) );
  XOR U11162 ( .A(n9008), .B(n9009), .Z(n8828) );
  AND U11163 ( .A(n9010), .B(n9011), .Z(n9008) );
  AND U11164 ( .A(a[55]), .B(b[24]), .Z(n9007) );
  XOR U11165 ( .A(n9012), .B(n8833), .Z(n8835) );
  XOR U11166 ( .A(n9013), .B(n9014), .Z(n8833) );
  AND U11167 ( .A(n9015), .B(n9016), .Z(n9013) );
  AND U11168 ( .A(a[56]), .B(b[23]), .Z(n9012) );
  XOR U11169 ( .A(n9017), .B(n8838), .Z(n8840) );
  XOR U11170 ( .A(n9018), .B(n9019), .Z(n8838) );
  AND U11171 ( .A(n9020), .B(n9021), .Z(n9018) );
  AND U11172 ( .A(a[57]), .B(b[22]), .Z(n9017) );
  XOR U11173 ( .A(n9022), .B(n8843), .Z(n8845) );
  XOR U11174 ( .A(n9023), .B(n9024), .Z(n8843) );
  AND U11175 ( .A(n9025), .B(n9026), .Z(n9023) );
  AND U11176 ( .A(a[58]), .B(b[21]), .Z(n9022) );
  XOR U11177 ( .A(n9027), .B(n8848), .Z(n8850) );
  XOR U11178 ( .A(n9028), .B(n9029), .Z(n8848) );
  AND U11179 ( .A(n9030), .B(n9031), .Z(n9028) );
  AND U11180 ( .A(a[59]), .B(b[20]), .Z(n9027) );
  XOR U11181 ( .A(n9032), .B(n8853), .Z(n8855) );
  XOR U11182 ( .A(n9033), .B(n9034), .Z(n8853) );
  AND U11183 ( .A(n9035), .B(n9036), .Z(n9033) );
  AND U11184 ( .A(a[60]), .B(b[19]), .Z(n9032) );
  XOR U11185 ( .A(n9037), .B(n8858), .Z(n8860) );
  XOR U11186 ( .A(n9038), .B(n9039), .Z(n8858) );
  AND U11187 ( .A(n9040), .B(n9041), .Z(n9038) );
  AND U11188 ( .A(a[61]), .B(b[18]), .Z(n9037) );
  XOR U11189 ( .A(n9042), .B(n8863), .Z(n8865) );
  XOR U11190 ( .A(n9043), .B(n9044), .Z(n8863) );
  AND U11191 ( .A(n9045), .B(n9046), .Z(n9043) );
  AND U11192 ( .A(a[62]), .B(b[17]), .Z(n9042) );
  XOR U11193 ( .A(n9047), .B(n8868), .Z(n8870) );
  XOR U11194 ( .A(n9048), .B(n9049), .Z(n8868) );
  AND U11195 ( .A(n9050), .B(n9051), .Z(n9048) );
  AND U11196 ( .A(a[63]), .B(b[16]), .Z(n9047) );
  XOR U11197 ( .A(n9052), .B(n8873), .Z(n8875) );
  XOR U11198 ( .A(n9053), .B(n9054), .Z(n8873) );
  AND U11199 ( .A(n9055), .B(n9056), .Z(n9053) );
  AND U11200 ( .A(a[64]), .B(b[15]), .Z(n9052) );
  XOR U11201 ( .A(n9057), .B(n8878), .Z(n8880) );
  XOR U11202 ( .A(n9058), .B(n9059), .Z(n8878) );
  AND U11203 ( .A(n9060), .B(n9061), .Z(n9058) );
  AND U11204 ( .A(a[65]), .B(b[14]), .Z(n9057) );
  XOR U11205 ( .A(n9062), .B(n8883), .Z(n8885) );
  XOR U11206 ( .A(n9063), .B(n9064), .Z(n8883) );
  AND U11207 ( .A(n9065), .B(n9066), .Z(n9063) );
  AND U11208 ( .A(a[66]), .B(b[13]), .Z(n9062) );
  XOR U11209 ( .A(n9067), .B(n9068), .Z(n8887) );
  AND U11210 ( .A(n9069), .B(n9070), .Z(n9067) );
  XOR U11211 ( .A(n9071), .B(n8892), .Z(n8894) );
  XOR U11212 ( .A(n9072), .B(n9073), .Z(n8892) );
  AND U11213 ( .A(n9074), .B(n9075), .Z(n9072) );
  AND U11214 ( .A(a[67]), .B(b[12]), .Z(n9071) );
  XOR U11215 ( .A(n9077), .B(n9078), .Z(n8897) );
  AND U11216 ( .A(n9079), .B(n9080), .Z(n9077) );
  AND U11217 ( .A(a[69]), .B(b[10]), .Z(n9076) );
  XOR U11218 ( .A(n9082), .B(n9083), .Z(n8902) );
  AND U11219 ( .A(n9084), .B(n9085), .Z(n9082) );
  AND U11220 ( .A(a[70]), .B(b[9]), .Z(n9081) );
  XOR U11221 ( .A(n9087), .B(n9088), .Z(n8907) );
  AND U11222 ( .A(n9089), .B(n9090), .Z(n9087) );
  AND U11223 ( .A(a[71]), .B(b[8]), .Z(n9086) );
  XOR U11224 ( .A(n9092), .B(n9093), .Z(n8912) );
  AND U11225 ( .A(n9094), .B(n9095), .Z(n9092) );
  AND U11226 ( .A(a[72]), .B(b[7]), .Z(n9091) );
  XOR U11227 ( .A(n9097), .B(n9098), .Z(n8917) );
  AND U11228 ( .A(n9099), .B(n9100), .Z(n9097) );
  AND U11229 ( .A(a[73]), .B(b[6]), .Z(n9096) );
  XOR U11230 ( .A(n9102), .B(n9103), .Z(n8922) );
  AND U11231 ( .A(n9104), .B(n9105), .Z(n9102) );
  AND U11232 ( .A(a[74]), .B(b[5]), .Z(n9101) );
  XOR U11233 ( .A(n9107), .B(n9108), .Z(n8927) );
  AND U11234 ( .A(n9109), .B(n9110), .Z(n9107) );
  AND U11235 ( .A(a[75]), .B(b[4]), .Z(n9106) );
  XOR U11236 ( .A(n9112), .B(n9113), .Z(n8932) );
  AND U11237 ( .A(n9114), .B(n9115), .Z(n9112) );
  AND U11238 ( .A(a[76]), .B(b[3]), .Z(n9111) );
  XOR U11239 ( .A(n9117), .B(n9118), .Z(n8937) );
  OR U11240 ( .A(n9119), .B(n9120), .Z(n9118) );
  AND U11241 ( .A(a[77]), .B(b[2]), .Z(n9116) );
  XNOR U11242 ( .A(n8947), .B(n9121), .Z(n8943) );
  NAND U11243 ( .A(a[78]), .B(b[1]), .Z(n9121) );
  IV U11244 ( .A(n8941), .Z(n8947) );
  ANDN U11245 ( .B(n5162), .A(n5164), .Z(n8941) );
  NAND U11246 ( .A(a[78]), .B(b[0]), .Z(n5164) );
  XOR U11247 ( .A(n9119), .B(n9120), .Z(n5162) );
  XOR U11248 ( .A(n9123), .B(n9114), .Z(n9122) );
  XOR U11249 ( .A(n9109), .B(n9113), .Z(n9124) );
  XOR U11250 ( .A(n9104), .B(n9108), .Z(n9125) );
  XOR U11251 ( .A(n9099), .B(n9103), .Z(n9126) );
  XOR U11252 ( .A(n9094), .B(n9098), .Z(n9127) );
  XOR U11253 ( .A(n9089), .B(n9093), .Z(n9128) );
  XOR U11254 ( .A(n9084), .B(n9088), .Z(n9129) );
  XOR U11255 ( .A(n9079), .B(n9083), .Z(n9130) );
  XOR U11256 ( .A(n9069), .B(n9078), .Z(n9131) );
  XOR U11257 ( .A(n9132), .B(n9068), .Z(n9069) );
  AND U11258 ( .A(b[10]), .B(a[68]), .Z(n9132) );
  XNOR U11259 ( .A(n9068), .B(n9074), .Z(n9133) );
  XNOR U11260 ( .A(n9073), .B(n9065), .Z(n9134) );
  XNOR U11261 ( .A(n9064), .B(n9060), .Z(n9135) );
  XNOR U11262 ( .A(n9059), .B(n9055), .Z(n9136) );
  XNOR U11263 ( .A(n9054), .B(n9050), .Z(n9137) );
  XNOR U11264 ( .A(n9049), .B(n9045), .Z(n9138) );
  XNOR U11265 ( .A(n9044), .B(n9040), .Z(n9139) );
  XNOR U11266 ( .A(n9039), .B(n9035), .Z(n9140) );
  XNOR U11267 ( .A(n9034), .B(n9030), .Z(n9141) );
  XNOR U11268 ( .A(n9029), .B(n9025), .Z(n9142) );
  XNOR U11269 ( .A(n9024), .B(n9020), .Z(n9143) );
  XNOR U11270 ( .A(n9019), .B(n9015), .Z(n9144) );
  XNOR U11271 ( .A(n9014), .B(n9010), .Z(n9145) );
  XNOR U11272 ( .A(n9009), .B(n9005), .Z(n9146) );
  XNOR U11273 ( .A(n9004), .B(n9000), .Z(n9147) );
  XNOR U11274 ( .A(n8999), .B(n8995), .Z(n9148) );
  XNOR U11275 ( .A(n8994), .B(n8990), .Z(n9149) );
  XOR U11276 ( .A(n8989), .B(n8986), .Z(n9150) );
  XOR U11277 ( .A(n9151), .B(n9152), .Z(n8986) );
  XOR U11278 ( .A(n8984), .B(n9153), .Z(n9152) );
  XOR U11279 ( .A(n9154), .B(n9155), .Z(n9153) );
  XOR U11280 ( .A(n9156), .B(n9157), .Z(n9155) );
  NAND U11281 ( .A(a[48]), .B(b[30]), .Z(n9157) );
  AND U11282 ( .A(a[47]), .B(b[31]), .Z(n9156) );
  XOR U11283 ( .A(n9158), .B(n9154), .Z(n9151) );
  XOR U11284 ( .A(n9159), .B(n9160), .Z(n9154) );
  ANDN U11285 ( .B(n9161), .A(n9162), .Z(n9159) );
  AND U11286 ( .A(a[49]), .B(b[29]), .Z(n9158) );
  XOR U11287 ( .A(n9163), .B(n8984), .Z(n8985) );
  XOR U11288 ( .A(n9164), .B(n9165), .Z(n8984) );
  AND U11289 ( .A(n9166), .B(n9167), .Z(n9164) );
  AND U11290 ( .A(a[50]), .B(b[28]), .Z(n9163) );
  XOR U11291 ( .A(n9168), .B(n8989), .Z(n8991) );
  XOR U11292 ( .A(n9169), .B(n9170), .Z(n8989) );
  AND U11293 ( .A(n9171), .B(n9172), .Z(n9169) );
  AND U11294 ( .A(a[51]), .B(b[27]), .Z(n9168) );
  XOR U11295 ( .A(n9173), .B(n8994), .Z(n8996) );
  XOR U11296 ( .A(n9174), .B(n9175), .Z(n8994) );
  AND U11297 ( .A(n9176), .B(n9177), .Z(n9174) );
  AND U11298 ( .A(a[52]), .B(b[26]), .Z(n9173) );
  XOR U11299 ( .A(n9178), .B(n8999), .Z(n9001) );
  XOR U11300 ( .A(n9179), .B(n9180), .Z(n8999) );
  AND U11301 ( .A(n9181), .B(n9182), .Z(n9179) );
  AND U11302 ( .A(a[53]), .B(b[25]), .Z(n9178) );
  XOR U11303 ( .A(n9183), .B(n9004), .Z(n9006) );
  XOR U11304 ( .A(n9184), .B(n9185), .Z(n9004) );
  AND U11305 ( .A(n9186), .B(n9187), .Z(n9184) );
  AND U11306 ( .A(a[54]), .B(b[24]), .Z(n9183) );
  XOR U11307 ( .A(n9188), .B(n9009), .Z(n9011) );
  XOR U11308 ( .A(n9189), .B(n9190), .Z(n9009) );
  AND U11309 ( .A(n9191), .B(n9192), .Z(n9189) );
  AND U11310 ( .A(a[55]), .B(b[23]), .Z(n9188) );
  XOR U11311 ( .A(n9193), .B(n9014), .Z(n9016) );
  XOR U11312 ( .A(n9194), .B(n9195), .Z(n9014) );
  AND U11313 ( .A(n9196), .B(n9197), .Z(n9194) );
  AND U11314 ( .A(a[56]), .B(b[22]), .Z(n9193) );
  XOR U11315 ( .A(n9198), .B(n9019), .Z(n9021) );
  XOR U11316 ( .A(n9199), .B(n9200), .Z(n9019) );
  AND U11317 ( .A(n9201), .B(n9202), .Z(n9199) );
  AND U11318 ( .A(a[57]), .B(b[21]), .Z(n9198) );
  XOR U11319 ( .A(n9203), .B(n9024), .Z(n9026) );
  XOR U11320 ( .A(n9204), .B(n9205), .Z(n9024) );
  AND U11321 ( .A(n9206), .B(n9207), .Z(n9204) );
  AND U11322 ( .A(a[58]), .B(b[20]), .Z(n9203) );
  XOR U11323 ( .A(n9208), .B(n9029), .Z(n9031) );
  XOR U11324 ( .A(n9209), .B(n9210), .Z(n9029) );
  AND U11325 ( .A(n9211), .B(n9212), .Z(n9209) );
  AND U11326 ( .A(a[59]), .B(b[19]), .Z(n9208) );
  XOR U11327 ( .A(n9213), .B(n9034), .Z(n9036) );
  XOR U11328 ( .A(n9214), .B(n9215), .Z(n9034) );
  AND U11329 ( .A(n9216), .B(n9217), .Z(n9214) );
  AND U11330 ( .A(a[60]), .B(b[18]), .Z(n9213) );
  XOR U11331 ( .A(n9218), .B(n9039), .Z(n9041) );
  XOR U11332 ( .A(n9219), .B(n9220), .Z(n9039) );
  AND U11333 ( .A(n9221), .B(n9222), .Z(n9219) );
  AND U11334 ( .A(a[61]), .B(b[17]), .Z(n9218) );
  XOR U11335 ( .A(n9223), .B(n9044), .Z(n9046) );
  XOR U11336 ( .A(n9224), .B(n9225), .Z(n9044) );
  AND U11337 ( .A(n9226), .B(n9227), .Z(n9224) );
  AND U11338 ( .A(a[62]), .B(b[16]), .Z(n9223) );
  XOR U11339 ( .A(n9228), .B(n9049), .Z(n9051) );
  XOR U11340 ( .A(n9229), .B(n9230), .Z(n9049) );
  AND U11341 ( .A(n9231), .B(n9232), .Z(n9229) );
  AND U11342 ( .A(a[63]), .B(b[15]), .Z(n9228) );
  XOR U11343 ( .A(n9233), .B(n9054), .Z(n9056) );
  XOR U11344 ( .A(n9234), .B(n9235), .Z(n9054) );
  AND U11345 ( .A(n9236), .B(n9237), .Z(n9234) );
  AND U11346 ( .A(a[64]), .B(b[14]), .Z(n9233) );
  XOR U11347 ( .A(n9238), .B(n9059), .Z(n9061) );
  XOR U11348 ( .A(n9239), .B(n9240), .Z(n9059) );
  AND U11349 ( .A(n9241), .B(n9242), .Z(n9239) );
  AND U11350 ( .A(a[65]), .B(b[13]), .Z(n9238) );
  XOR U11351 ( .A(n9243), .B(n9064), .Z(n9066) );
  XOR U11352 ( .A(n9244), .B(n9245), .Z(n9064) );
  AND U11353 ( .A(n9246), .B(n9247), .Z(n9244) );
  AND U11354 ( .A(a[66]), .B(b[12]), .Z(n9243) );
  XOR U11355 ( .A(n9248), .B(n9249), .Z(n9068) );
  AND U11356 ( .A(n9250), .B(n9251), .Z(n9248) );
  XOR U11357 ( .A(n9252), .B(n9073), .Z(n9075) );
  XOR U11358 ( .A(n9253), .B(n9254), .Z(n9073) );
  AND U11359 ( .A(n9255), .B(n9256), .Z(n9253) );
  AND U11360 ( .A(a[67]), .B(b[11]), .Z(n9252) );
  XOR U11361 ( .A(n9258), .B(n9259), .Z(n9078) );
  AND U11362 ( .A(n9260), .B(n9261), .Z(n9258) );
  AND U11363 ( .A(a[69]), .B(b[9]), .Z(n9257) );
  XOR U11364 ( .A(n9263), .B(n9264), .Z(n9083) );
  AND U11365 ( .A(n9265), .B(n9266), .Z(n9263) );
  AND U11366 ( .A(a[70]), .B(b[8]), .Z(n9262) );
  XOR U11367 ( .A(n9268), .B(n9269), .Z(n9088) );
  AND U11368 ( .A(n9270), .B(n9271), .Z(n9268) );
  AND U11369 ( .A(a[71]), .B(b[7]), .Z(n9267) );
  XOR U11370 ( .A(n9273), .B(n9274), .Z(n9093) );
  AND U11371 ( .A(n9275), .B(n9276), .Z(n9273) );
  AND U11372 ( .A(a[72]), .B(b[6]), .Z(n9272) );
  XOR U11373 ( .A(n9278), .B(n9279), .Z(n9098) );
  AND U11374 ( .A(n9280), .B(n9281), .Z(n9278) );
  AND U11375 ( .A(a[73]), .B(b[5]), .Z(n9277) );
  XOR U11376 ( .A(n9283), .B(n9284), .Z(n9103) );
  AND U11377 ( .A(n9285), .B(n9286), .Z(n9283) );
  AND U11378 ( .A(a[74]), .B(b[4]), .Z(n9282) );
  XOR U11379 ( .A(n9288), .B(n9289), .Z(n9108) );
  AND U11380 ( .A(n9290), .B(n9291), .Z(n9288) );
  AND U11381 ( .A(a[75]), .B(b[3]), .Z(n9287) );
  XOR U11382 ( .A(n9293), .B(n9294), .Z(n9113) );
  OR U11383 ( .A(n9295), .B(n9296), .Z(n9294) );
  AND U11384 ( .A(a[76]), .B(b[2]), .Z(n9292) );
  XNOR U11385 ( .A(n9123), .B(n9297), .Z(n9119) );
  NAND U11386 ( .A(a[77]), .B(b[1]), .Z(n9297) );
  IV U11387 ( .A(n9117), .Z(n9123) );
  ANDN U11388 ( .B(n5167), .A(n5169), .Z(n9117) );
  NAND U11389 ( .A(a[77]), .B(b[0]), .Z(n5169) );
  XOR U11390 ( .A(n9295), .B(n9296), .Z(n5167) );
  XOR U11391 ( .A(n9299), .B(n9290), .Z(n9298) );
  XOR U11392 ( .A(n9285), .B(n9289), .Z(n9300) );
  XOR U11393 ( .A(n9280), .B(n9284), .Z(n9301) );
  XOR U11394 ( .A(n9275), .B(n9279), .Z(n9302) );
  XOR U11395 ( .A(n9270), .B(n9274), .Z(n9303) );
  XOR U11396 ( .A(n9265), .B(n9269), .Z(n9304) );
  XOR U11397 ( .A(n9260), .B(n9264), .Z(n9305) );
  XOR U11398 ( .A(n9250), .B(n9259), .Z(n9306) );
  XOR U11399 ( .A(n9307), .B(n9249), .Z(n9250) );
  AND U11400 ( .A(b[9]), .B(a[68]), .Z(n9307) );
  XNOR U11401 ( .A(n9249), .B(n9255), .Z(n9308) );
  XNOR U11402 ( .A(n9254), .B(n9246), .Z(n9309) );
  XNOR U11403 ( .A(n9245), .B(n9241), .Z(n9310) );
  XNOR U11404 ( .A(n9240), .B(n9236), .Z(n9311) );
  XNOR U11405 ( .A(n9235), .B(n9231), .Z(n9312) );
  XNOR U11406 ( .A(n9230), .B(n9226), .Z(n9313) );
  XNOR U11407 ( .A(n9225), .B(n9221), .Z(n9314) );
  XNOR U11408 ( .A(n9220), .B(n9216), .Z(n9315) );
  XNOR U11409 ( .A(n9215), .B(n9211), .Z(n9316) );
  XNOR U11410 ( .A(n9210), .B(n9206), .Z(n9317) );
  XNOR U11411 ( .A(n9205), .B(n9201), .Z(n9318) );
  XNOR U11412 ( .A(n9200), .B(n9196), .Z(n9319) );
  XNOR U11413 ( .A(n9195), .B(n9191), .Z(n9320) );
  XNOR U11414 ( .A(n9190), .B(n9186), .Z(n9321) );
  XNOR U11415 ( .A(n9185), .B(n9181), .Z(n9322) );
  XNOR U11416 ( .A(n9180), .B(n9176), .Z(n9323) );
  XNOR U11417 ( .A(n9175), .B(n9171), .Z(n9324) );
  XNOR U11418 ( .A(n9170), .B(n9166), .Z(n9325) );
  XOR U11419 ( .A(n9165), .B(n9162), .Z(n9326) );
  XOR U11420 ( .A(n9327), .B(n9328), .Z(n9162) );
  XOR U11421 ( .A(n9160), .B(n9329), .Z(n9328) );
  XOR U11422 ( .A(n9330), .B(n9331), .Z(n9329) );
  XOR U11423 ( .A(n9332), .B(n9333), .Z(n9331) );
  NAND U11424 ( .A(a[47]), .B(b[30]), .Z(n9333) );
  AND U11425 ( .A(a[46]), .B(b[31]), .Z(n9332) );
  XOR U11426 ( .A(n9334), .B(n9330), .Z(n9327) );
  XOR U11427 ( .A(n9335), .B(n9336), .Z(n9330) );
  ANDN U11428 ( .B(n9337), .A(n9338), .Z(n9335) );
  AND U11429 ( .A(a[48]), .B(b[29]), .Z(n9334) );
  XOR U11430 ( .A(n9339), .B(n9160), .Z(n9161) );
  XOR U11431 ( .A(n9340), .B(n9341), .Z(n9160) );
  AND U11432 ( .A(n9342), .B(n9343), .Z(n9340) );
  AND U11433 ( .A(a[49]), .B(b[28]), .Z(n9339) );
  XOR U11434 ( .A(n9344), .B(n9165), .Z(n9167) );
  XOR U11435 ( .A(n9345), .B(n9346), .Z(n9165) );
  AND U11436 ( .A(n9347), .B(n9348), .Z(n9345) );
  AND U11437 ( .A(a[50]), .B(b[27]), .Z(n9344) );
  XOR U11438 ( .A(n9349), .B(n9170), .Z(n9172) );
  XOR U11439 ( .A(n9350), .B(n9351), .Z(n9170) );
  AND U11440 ( .A(n9352), .B(n9353), .Z(n9350) );
  AND U11441 ( .A(a[51]), .B(b[26]), .Z(n9349) );
  XOR U11442 ( .A(n9354), .B(n9175), .Z(n9177) );
  XOR U11443 ( .A(n9355), .B(n9356), .Z(n9175) );
  AND U11444 ( .A(n9357), .B(n9358), .Z(n9355) );
  AND U11445 ( .A(a[52]), .B(b[25]), .Z(n9354) );
  XOR U11446 ( .A(n9359), .B(n9180), .Z(n9182) );
  XOR U11447 ( .A(n9360), .B(n9361), .Z(n9180) );
  AND U11448 ( .A(n9362), .B(n9363), .Z(n9360) );
  AND U11449 ( .A(a[53]), .B(b[24]), .Z(n9359) );
  XOR U11450 ( .A(n9364), .B(n9185), .Z(n9187) );
  XOR U11451 ( .A(n9365), .B(n9366), .Z(n9185) );
  AND U11452 ( .A(n9367), .B(n9368), .Z(n9365) );
  AND U11453 ( .A(a[54]), .B(b[23]), .Z(n9364) );
  XOR U11454 ( .A(n9369), .B(n9190), .Z(n9192) );
  XOR U11455 ( .A(n9370), .B(n9371), .Z(n9190) );
  AND U11456 ( .A(n9372), .B(n9373), .Z(n9370) );
  AND U11457 ( .A(a[55]), .B(b[22]), .Z(n9369) );
  XOR U11458 ( .A(n9374), .B(n9195), .Z(n9197) );
  XOR U11459 ( .A(n9375), .B(n9376), .Z(n9195) );
  AND U11460 ( .A(n9377), .B(n9378), .Z(n9375) );
  AND U11461 ( .A(a[56]), .B(b[21]), .Z(n9374) );
  XOR U11462 ( .A(n9379), .B(n9200), .Z(n9202) );
  XOR U11463 ( .A(n9380), .B(n9381), .Z(n9200) );
  AND U11464 ( .A(n9382), .B(n9383), .Z(n9380) );
  AND U11465 ( .A(a[57]), .B(b[20]), .Z(n9379) );
  XOR U11466 ( .A(n9384), .B(n9205), .Z(n9207) );
  XOR U11467 ( .A(n9385), .B(n9386), .Z(n9205) );
  AND U11468 ( .A(n9387), .B(n9388), .Z(n9385) );
  AND U11469 ( .A(a[58]), .B(b[19]), .Z(n9384) );
  XOR U11470 ( .A(n9389), .B(n9210), .Z(n9212) );
  XOR U11471 ( .A(n9390), .B(n9391), .Z(n9210) );
  AND U11472 ( .A(n9392), .B(n9393), .Z(n9390) );
  AND U11473 ( .A(a[59]), .B(b[18]), .Z(n9389) );
  XOR U11474 ( .A(n9394), .B(n9215), .Z(n9217) );
  XOR U11475 ( .A(n9395), .B(n9396), .Z(n9215) );
  AND U11476 ( .A(n9397), .B(n9398), .Z(n9395) );
  AND U11477 ( .A(a[60]), .B(b[17]), .Z(n9394) );
  XOR U11478 ( .A(n9399), .B(n9220), .Z(n9222) );
  XOR U11479 ( .A(n9400), .B(n9401), .Z(n9220) );
  AND U11480 ( .A(n9402), .B(n9403), .Z(n9400) );
  AND U11481 ( .A(a[61]), .B(b[16]), .Z(n9399) );
  XOR U11482 ( .A(n9404), .B(n9225), .Z(n9227) );
  XOR U11483 ( .A(n9405), .B(n9406), .Z(n9225) );
  AND U11484 ( .A(n9407), .B(n9408), .Z(n9405) );
  AND U11485 ( .A(a[62]), .B(b[15]), .Z(n9404) );
  XOR U11486 ( .A(n9409), .B(n9230), .Z(n9232) );
  XOR U11487 ( .A(n9410), .B(n9411), .Z(n9230) );
  AND U11488 ( .A(n9412), .B(n9413), .Z(n9410) );
  AND U11489 ( .A(a[63]), .B(b[14]), .Z(n9409) );
  XOR U11490 ( .A(n9414), .B(n9235), .Z(n9237) );
  XOR U11491 ( .A(n9415), .B(n9416), .Z(n9235) );
  AND U11492 ( .A(n9417), .B(n9418), .Z(n9415) );
  AND U11493 ( .A(a[64]), .B(b[13]), .Z(n9414) );
  XOR U11494 ( .A(n9419), .B(n9240), .Z(n9242) );
  XOR U11495 ( .A(n9420), .B(n9421), .Z(n9240) );
  AND U11496 ( .A(n9422), .B(n9423), .Z(n9420) );
  AND U11497 ( .A(a[65]), .B(b[12]), .Z(n9419) );
  XOR U11498 ( .A(n9424), .B(n9245), .Z(n9247) );
  XOR U11499 ( .A(n9425), .B(n9426), .Z(n9245) );
  AND U11500 ( .A(n9427), .B(n9428), .Z(n9425) );
  AND U11501 ( .A(a[66]), .B(b[11]), .Z(n9424) );
  XOR U11502 ( .A(n9429), .B(n9430), .Z(n9249) );
  AND U11503 ( .A(n9431), .B(n9432), .Z(n9429) );
  XOR U11504 ( .A(n9433), .B(n9254), .Z(n9256) );
  XOR U11505 ( .A(n9434), .B(n9435), .Z(n9254) );
  AND U11506 ( .A(n9436), .B(n9437), .Z(n9434) );
  AND U11507 ( .A(a[67]), .B(b[10]), .Z(n9433) );
  XOR U11508 ( .A(n9439), .B(n9440), .Z(n9259) );
  AND U11509 ( .A(n9441), .B(n9442), .Z(n9439) );
  AND U11510 ( .A(a[69]), .B(b[8]), .Z(n9438) );
  XOR U11511 ( .A(n9444), .B(n9445), .Z(n9264) );
  AND U11512 ( .A(n9446), .B(n9447), .Z(n9444) );
  AND U11513 ( .A(a[70]), .B(b[7]), .Z(n9443) );
  XOR U11514 ( .A(n9449), .B(n9450), .Z(n9269) );
  AND U11515 ( .A(n9451), .B(n9452), .Z(n9449) );
  AND U11516 ( .A(a[71]), .B(b[6]), .Z(n9448) );
  XOR U11517 ( .A(n9454), .B(n9455), .Z(n9274) );
  AND U11518 ( .A(n9456), .B(n9457), .Z(n9454) );
  AND U11519 ( .A(a[72]), .B(b[5]), .Z(n9453) );
  XOR U11520 ( .A(n9459), .B(n9460), .Z(n9279) );
  AND U11521 ( .A(n9461), .B(n9462), .Z(n9459) );
  AND U11522 ( .A(a[73]), .B(b[4]), .Z(n9458) );
  XOR U11523 ( .A(n9464), .B(n9465), .Z(n9284) );
  AND U11524 ( .A(n9466), .B(n9467), .Z(n9464) );
  AND U11525 ( .A(a[74]), .B(b[3]), .Z(n9463) );
  XOR U11526 ( .A(n9469), .B(n9470), .Z(n9289) );
  OR U11527 ( .A(n9471), .B(n9472), .Z(n9470) );
  AND U11528 ( .A(a[75]), .B(b[2]), .Z(n9468) );
  XNOR U11529 ( .A(n9299), .B(n9473), .Z(n9295) );
  NAND U11530 ( .A(a[76]), .B(b[1]), .Z(n9473) );
  IV U11531 ( .A(n9293), .Z(n9299) );
  ANDN U11532 ( .B(n5172), .A(n5174), .Z(n9293) );
  NAND U11533 ( .A(a[76]), .B(b[0]), .Z(n5174) );
  XOR U11534 ( .A(n9471), .B(n9472), .Z(n5172) );
  XOR U11535 ( .A(n9475), .B(n9466), .Z(n9474) );
  XOR U11536 ( .A(n9461), .B(n9465), .Z(n9476) );
  XOR U11537 ( .A(n9456), .B(n9460), .Z(n9477) );
  XOR U11538 ( .A(n9451), .B(n9455), .Z(n9478) );
  XOR U11539 ( .A(n9446), .B(n9450), .Z(n9479) );
  XOR U11540 ( .A(n9441), .B(n9445), .Z(n9480) );
  XOR U11541 ( .A(n9431), .B(n9440), .Z(n9481) );
  XOR U11542 ( .A(n9482), .B(n9430), .Z(n9431) );
  AND U11543 ( .A(b[8]), .B(a[68]), .Z(n9482) );
  XNOR U11544 ( .A(n9430), .B(n9436), .Z(n9483) );
  XNOR U11545 ( .A(n9435), .B(n9427), .Z(n9484) );
  XNOR U11546 ( .A(n9426), .B(n9422), .Z(n9485) );
  XNOR U11547 ( .A(n9421), .B(n9417), .Z(n9486) );
  XNOR U11548 ( .A(n9416), .B(n9412), .Z(n9487) );
  XNOR U11549 ( .A(n9411), .B(n9407), .Z(n9488) );
  XNOR U11550 ( .A(n9406), .B(n9402), .Z(n9489) );
  XNOR U11551 ( .A(n9401), .B(n9397), .Z(n9490) );
  XNOR U11552 ( .A(n9396), .B(n9392), .Z(n9491) );
  XNOR U11553 ( .A(n9391), .B(n9387), .Z(n9492) );
  XNOR U11554 ( .A(n9386), .B(n9382), .Z(n9493) );
  XNOR U11555 ( .A(n9381), .B(n9377), .Z(n9494) );
  XNOR U11556 ( .A(n9376), .B(n9372), .Z(n9495) );
  XNOR U11557 ( .A(n9371), .B(n9367), .Z(n9496) );
  XNOR U11558 ( .A(n9366), .B(n9362), .Z(n9497) );
  XNOR U11559 ( .A(n9361), .B(n9357), .Z(n9498) );
  XNOR U11560 ( .A(n9356), .B(n9352), .Z(n9499) );
  XNOR U11561 ( .A(n9351), .B(n9347), .Z(n9500) );
  XNOR U11562 ( .A(n9346), .B(n9342), .Z(n9501) );
  XOR U11563 ( .A(n9341), .B(n9338), .Z(n9502) );
  XOR U11564 ( .A(n9503), .B(n9504), .Z(n9338) );
  XOR U11565 ( .A(n9336), .B(n9505), .Z(n9504) );
  XOR U11566 ( .A(n9506), .B(n9507), .Z(n9505) );
  XOR U11567 ( .A(n9508), .B(n9509), .Z(n9507) );
  NAND U11568 ( .A(a[46]), .B(b[30]), .Z(n9509) );
  AND U11569 ( .A(a[45]), .B(b[31]), .Z(n9508) );
  XOR U11570 ( .A(n9510), .B(n9506), .Z(n9503) );
  XOR U11571 ( .A(n9511), .B(n9512), .Z(n9506) );
  ANDN U11572 ( .B(n9513), .A(n9514), .Z(n9511) );
  AND U11573 ( .A(a[47]), .B(b[29]), .Z(n9510) );
  XOR U11574 ( .A(n9515), .B(n9336), .Z(n9337) );
  XOR U11575 ( .A(n9516), .B(n9517), .Z(n9336) );
  AND U11576 ( .A(n9518), .B(n9519), .Z(n9516) );
  AND U11577 ( .A(a[48]), .B(b[28]), .Z(n9515) );
  XOR U11578 ( .A(n9520), .B(n9341), .Z(n9343) );
  XOR U11579 ( .A(n9521), .B(n9522), .Z(n9341) );
  AND U11580 ( .A(n9523), .B(n9524), .Z(n9521) );
  AND U11581 ( .A(a[49]), .B(b[27]), .Z(n9520) );
  XOR U11582 ( .A(n9525), .B(n9346), .Z(n9348) );
  XOR U11583 ( .A(n9526), .B(n9527), .Z(n9346) );
  AND U11584 ( .A(n9528), .B(n9529), .Z(n9526) );
  AND U11585 ( .A(a[50]), .B(b[26]), .Z(n9525) );
  XOR U11586 ( .A(n9530), .B(n9351), .Z(n9353) );
  XOR U11587 ( .A(n9531), .B(n9532), .Z(n9351) );
  AND U11588 ( .A(n9533), .B(n9534), .Z(n9531) );
  AND U11589 ( .A(a[51]), .B(b[25]), .Z(n9530) );
  XOR U11590 ( .A(n9535), .B(n9356), .Z(n9358) );
  XOR U11591 ( .A(n9536), .B(n9537), .Z(n9356) );
  AND U11592 ( .A(n9538), .B(n9539), .Z(n9536) );
  AND U11593 ( .A(a[52]), .B(b[24]), .Z(n9535) );
  XOR U11594 ( .A(n9540), .B(n9361), .Z(n9363) );
  XOR U11595 ( .A(n9541), .B(n9542), .Z(n9361) );
  AND U11596 ( .A(n9543), .B(n9544), .Z(n9541) );
  AND U11597 ( .A(a[53]), .B(b[23]), .Z(n9540) );
  XOR U11598 ( .A(n9545), .B(n9366), .Z(n9368) );
  XOR U11599 ( .A(n9546), .B(n9547), .Z(n9366) );
  AND U11600 ( .A(n9548), .B(n9549), .Z(n9546) );
  AND U11601 ( .A(a[54]), .B(b[22]), .Z(n9545) );
  XOR U11602 ( .A(n9550), .B(n9371), .Z(n9373) );
  XOR U11603 ( .A(n9551), .B(n9552), .Z(n9371) );
  AND U11604 ( .A(n9553), .B(n9554), .Z(n9551) );
  AND U11605 ( .A(a[55]), .B(b[21]), .Z(n9550) );
  XOR U11606 ( .A(n9555), .B(n9376), .Z(n9378) );
  XOR U11607 ( .A(n9556), .B(n9557), .Z(n9376) );
  AND U11608 ( .A(n9558), .B(n9559), .Z(n9556) );
  AND U11609 ( .A(a[56]), .B(b[20]), .Z(n9555) );
  XOR U11610 ( .A(n9560), .B(n9381), .Z(n9383) );
  XOR U11611 ( .A(n9561), .B(n9562), .Z(n9381) );
  AND U11612 ( .A(n9563), .B(n9564), .Z(n9561) );
  AND U11613 ( .A(a[57]), .B(b[19]), .Z(n9560) );
  XOR U11614 ( .A(n9565), .B(n9386), .Z(n9388) );
  XOR U11615 ( .A(n9566), .B(n9567), .Z(n9386) );
  AND U11616 ( .A(n9568), .B(n9569), .Z(n9566) );
  AND U11617 ( .A(a[58]), .B(b[18]), .Z(n9565) );
  XOR U11618 ( .A(n9570), .B(n9391), .Z(n9393) );
  XOR U11619 ( .A(n9571), .B(n9572), .Z(n9391) );
  AND U11620 ( .A(n9573), .B(n9574), .Z(n9571) );
  AND U11621 ( .A(a[59]), .B(b[17]), .Z(n9570) );
  XOR U11622 ( .A(n9575), .B(n9396), .Z(n9398) );
  XOR U11623 ( .A(n9576), .B(n9577), .Z(n9396) );
  AND U11624 ( .A(n9578), .B(n9579), .Z(n9576) );
  AND U11625 ( .A(a[60]), .B(b[16]), .Z(n9575) );
  XOR U11626 ( .A(n9580), .B(n9401), .Z(n9403) );
  XOR U11627 ( .A(n9581), .B(n9582), .Z(n9401) );
  AND U11628 ( .A(n9583), .B(n9584), .Z(n9581) );
  AND U11629 ( .A(a[61]), .B(b[15]), .Z(n9580) );
  XOR U11630 ( .A(n9585), .B(n9406), .Z(n9408) );
  XOR U11631 ( .A(n9586), .B(n9587), .Z(n9406) );
  AND U11632 ( .A(n9588), .B(n9589), .Z(n9586) );
  AND U11633 ( .A(a[62]), .B(b[14]), .Z(n9585) );
  XOR U11634 ( .A(n9590), .B(n9411), .Z(n9413) );
  XOR U11635 ( .A(n9591), .B(n9592), .Z(n9411) );
  AND U11636 ( .A(n9593), .B(n9594), .Z(n9591) );
  AND U11637 ( .A(a[63]), .B(b[13]), .Z(n9590) );
  XOR U11638 ( .A(n9595), .B(n9416), .Z(n9418) );
  XOR U11639 ( .A(n9596), .B(n9597), .Z(n9416) );
  AND U11640 ( .A(n9598), .B(n9599), .Z(n9596) );
  AND U11641 ( .A(a[64]), .B(b[12]), .Z(n9595) );
  XOR U11642 ( .A(n9600), .B(n9421), .Z(n9423) );
  XOR U11643 ( .A(n9601), .B(n9602), .Z(n9421) );
  AND U11644 ( .A(n9603), .B(n9604), .Z(n9601) );
  AND U11645 ( .A(a[65]), .B(b[11]), .Z(n9600) );
  XOR U11646 ( .A(n9605), .B(n9426), .Z(n9428) );
  XOR U11647 ( .A(n9606), .B(n9607), .Z(n9426) );
  AND U11648 ( .A(n9608), .B(n9609), .Z(n9606) );
  AND U11649 ( .A(a[66]), .B(b[10]), .Z(n9605) );
  XOR U11650 ( .A(n9610), .B(n9611), .Z(n9430) );
  AND U11651 ( .A(n9612), .B(n9613), .Z(n9610) );
  XOR U11652 ( .A(n9614), .B(n9435), .Z(n9437) );
  XOR U11653 ( .A(n9615), .B(n9616), .Z(n9435) );
  AND U11654 ( .A(n9617), .B(n9618), .Z(n9615) );
  AND U11655 ( .A(a[67]), .B(b[9]), .Z(n9614) );
  XOR U11656 ( .A(n9620), .B(n9621), .Z(n9440) );
  AND U11657 ( .A(n9622), .B(n9623), .Z(n9620) );
  AND U11658 ( .A(a[69]), .B(b[7]), .Z(n9619) );
  XOR U11659 ( .A(n9625), .B(n9626), .Z(n9445) );
  AND U11660 ( .A(n9627), .B(n9628), .Z(n9625) );
  AND U11661 ( .A(a[70]), .B(b[6]), .Z(n9624) );
  XOR U11662 ( .A(n9630), .B(n9631), .Z(n9450) );
  AND U11663 ( .A(n9632), .B(n9633), .Z(n9630) );
  AND U11664 ( .A(a[71]), .B(b[5]), .Z(n9629) );
  XOR U11665 ( .A(n9635), .B(n9636), .Z(n9455) );
  AND U11666 ( .A(n9637), .B(n9638), .Z(n9635) );
  AND U11667 ( .A(a[72]), .B(b[4]), .Z(n9634) );
  XOR U11668 ( .A(n9640), .B(n9641), .Z(n9460) );
  AND U11669 ( .A(n9642), .B(n9643), .Z(n9640) );
  AND U11670 ( .A(a[73]), .B(b[3]), .Z(n9639) );
  XOR U11671 ( .A(n9645), .B(n9646), .Z(n9465) );
  OR U11672 ( .A(n9647), .B(n9648), .Z(n9646) );
  AND U11673 ( .A(a[74]), .B(b[2]), .Z(n9644) );
  XNOR U11674 ( .A(n9475), .B(n9649), .Z(n9471) );
  NAND U11675 ( .A(a[75]), .B(b[1]), .Z(n9649) );
  IV U11676 ( .A(n9469), .Z(n9475) );
  ANDN U11677 ( .B(n5177), .A(n5179), .Z(n9469) );
  NAND U11678 ( .A(a[75]), .B(b[0]), .Z(n5179) );
  XOR U11679 ( .A(n9647), .B(n9648), .Z(n5177) );
  XOR U11680 ( .A(n9651), .B(n9642), .Z(n9650) );
  XOR U11681 ( .A(n9637), .B(n9641), .Z(n9652) );
  XOR U11682 ( .A(n9632), .B(n9636), .Z(n9653) );
  XOR U11683 ( .A(n9627), .B(n9631), .Z(n9654) );
  XOR U11684 ( .A(n9622), .B(n9626), .Z(n9655) );
  XOR U11685 ( .A(n9612), .B(n9621), .Z(n9656) );
  XOR U11686 ( .A(n9657), .B(n9611), .Z(n9612) );
  AND U11687 ( .A(b[7]), .B(a[68]), .Z(n9657) );
  XNOR U11688 ( .A(n9611), .B(n9617), .Z(n9658) );
  XNOR U11689 ( .A(n9616), .B(n9608), .Z(n9659) );
  XNOR U11690 ( .A(n9607), .B(n9603), .Z(n9660) );
  XNOR U11691 ( .A(n9602), .B(n9598), .Z(n9661) );
  XNOR U11692 ( .A(n9597), .B(n9593), .Z(n9662) );
  XNOR U11693 ( .A(n9592), .B(n9588), .Z(n9663) );
  XNOR U11694 ( .A(n9587), .B(n9583), .Z(n9664) );
  XNOR U11695 ( .A(n9582), .B(n9578), .Z(n9665) );
  XNOR U11696 ( .A(n9577), .B(n9573), .Z(n9666) );
  XNOR U11697 ( .A(n9572), .B(n9568), .Z(n9667) );
  XNOR U11698 ( .A(n9567), .B(n9563), .Z(n9668) );
  XNOR U11699 ( .A(n9562), .B(n9558), .Z(n9669) );
  XNOR U11700 ( .A(n9557), .B(n9553), .Z(n9670) );
  XNOR U11701 ( .A(n9552), .B(n9548), .Z(n9671) );
  XNOR U11702 ( .A(n9547), .B(n9543), .Z(n9672) );
  XNOR U11703 ( .A(n9542), .B(n9538), .Z(n9673) );
  XNOR U11704 ( .A(n9537), .B(n9533), .Z(n9674) );
  XNOR U11705 ( .A(n9532), .B(n9528), .Z(n9675) );
  XNOR U11706 ( .A(n9527), .B(n9523), .Z(n9676) );
  XNOR U11707 ( .A(n9522), .B(n9518), .Z(n9677) );
  XOR U11708 ( .A(n9517), .B(n9514), .Z(n9678) );
  XOR U11709 ( .A(n9679), .B(n9680), .Z(n9514) );
  XOR U11710 ( .A(n9512), .B(n9681), .Z(n9680) );
  XOR U11711 ( .A(n9682), .B(n9683), .Z(n9681) );
  XOR U11712 ( .A(n9684), .B(n9685), .Z(n9683) );
  NAND U11713 ( .A(a[45]), .B(b[30]), .Z(n9685) );
  AND U11714 ( .A(a[44]), .B(b[31]), .Z(n9684) );
  XOR U11715 ( .A(n9686), .B(n9682), .Z(n9679) );
  XOR U11716 ( .A(n9687), .B(n9688), .Z(n9682) );
  ANDN U11717 ( .B(n9689), .A(n9690), .Z(n9687) );
  AND U11718 ( .A(a[46]), .B(b[29]), .Z(n9686) );
  XOR U11719 ( .A(n9691), .B(n9512), .Z(n9513) );
  XOR U11720 ( .A(n9692), .B(n9693), .Z(n9512) );
  AND U11721 ( .A(n9694), .B(n9695), .Z(n9692) );
  AND U11722 ( .A(a[47]), .B(b[28]), .Z(n9691) );
  XOR U11723 ( .A(n9696), .B(n9517), .Z(n9519) );
  XOR U11724 ( .A(n9697), .B(n9698), .Z(n9517) );
  AND U11725 ( .A(n9699), .B(n9700), .Z(n9697) );
  AND U11726 ( .A(a[48]), .B(b[27]), .Z(n9696) );
  XOR U11727 ( .A(n9701), .B(n9522), .Z(n9524) );
  XOR U11728 ( .A(n9702), .B(n9703), .Z(n9522) );
  AND U11729 ( .A(n9704), .B(n9705), .Z(n9702) );
  AND U11730 ( .A(a[49]), .B(b[26]), .Z(n9701) );
  XOR U11731 ( .A(n9706), .B(n9527), .Z(n9529) );
  XOR U11732 ( .A(n9707), .B(n9708), .Z(n9527) );
  AND U11733 ( .A(n9709), .B(n9710), .Z(n9707) );
  AND U11734 ( .A(a[50]), .B(b[25]), .Z(n9706) );
  XOR U11735 ( .A(n9711), .B(n9532), .Z(n9534) );
  XOR U11736 ( .A(n9712), .B(n9713), .Z(n9532) );
  AND U11737 ( .A(n9714), .B(n9715), .Z(n9712) );
  AND U11738 ( .A(a[51]), .B(b[24]), .Z(n9711) );
  XOR U11739 ( .A(n9716), .B(n9537), .Z(n9539) );
  XOR U11740 ( .A(n9717), .B(n9718), .Z(n9537) );
  AND U11741 ( .A(n9719), .B(n9720), .Z(n9717) );
  AND U11742 ( .A(a[52]), .B(b[23]), .Z(n9716) );
  XOR U11743 ( .A(n9721), .B(n9542), .Z(n9544) );
  XOR U11744 ( .A(n9722), .B(n9723), .Z(n9542) );
  AND U11745 ( .A(n9724), .B(n9725), .Z(n9722) );
  AND U11746 ( .A(a[53]), .B(b[22]), .Z(n9721) );
  XOR U11747 ( .A(n9726), .B(n9547), .Z(n9549) );
  XOR U11748 ( .A(n9727), .B(n9728), .Z(n9547) );
  AND U11749 ( .A(n9729), .B(n9730), .Z(n9727) );
  AND U11750 ( .A(a[54]), .B(b[21]), .Z(n9726) );
  XOR U11751 ( .A(n9731), .B(n9552), .Z(n9554) );
  XOR U11752 ( .A(n9732), .B(n9733), .Z(n9552) );
  AND U11753 ( .A(n9734), .B(n9735), .Z(n9732) );
  AND U11754 ( .A(a[55]), .B(b[20]), .Z(n9731) );
  XOR U11755 ( .A(n9736), .B(n9557), .Z(n9559) );
  XOR U11756 ( .A(n9737), .B(n9738), .Z(n9557) );
  AND U11757 ( .A(n9739), .B(n9740), .Z(n9737) );
  AND U11758 ( .A(a[56]), .B(b[19]), .Z(n9736) );
  XOR U11759 ( .A(n9741), .B(n9562), .Z(n9564) );
  XOR U11760 ( .A(n9742), .B(n9743), .Z(n9562) );
  AND U11761 ( .A(n9744), .B(n9745), .Z(n9742) );
  AND U11762 ( .A(a[57]), .B(b[18]), .Z(n9741) );
  XOR U11763 ( .A(n9746), .B(n9567), .Z(n9569) );
  XOR U11764 ( .A(n9747), .B(n9748), .Z(n9567) );
  AND U11765 ( .A(n9749), .B(n9750), .Z(n9747) );
  AND U11766 ( .A(a[58]), .B(b[17]), .Z(n9746) );
  XOR U11767 ( .A(n9751), .B(n9572), .Z(n9574) );
  XOR U11768 ( .A(n9752), .B(n9753), .Z(n9572) );
  AND U11769 ( .A(n9754), .B(n9755), .Z(n9752) );
  AND U11770 ( .A(a[59]), .B(b[16]), .Z(n9751) );
  XOR U11771 ( .A(n9756), .B(n9577), .Z(n9579) );
  XOR U11772 ( .A(n9757), .B(n9758), .Z(n9577) );
  AND U11773 ( .A(n9759), .B(n9760), .Z(n9757) );
  AND U11774 ( .A(a[60]), .B(b[15]), .Z(n9756) );
  XOR U11775 ( .A(n9761), .B(n9582), .Z(n9584) );
  XOR U11776 ( .A(n9762), .B(n9763), .Z(n9582) );
  AND U11777 ( .A(n9764), .B(n9765), .Z(n9762) );
  AND U11778 ( .A(a[61]), .B(b[14]), .Z(n9761) );
  XOR U11779 ( .A(n9766), .B(n9587), .Z(n9589) );
  XOR U11780 ( .A(n9767), .B(n9768), .Z(n9587) );
  AND U11781 ( .A(n9769), .B(n9770), .Z(n9767) );
  AND U11782 ( .A(a[62]), .B(b[13]), .Z(n9766) );
  XOR U11783 ( .A(n9771), .B(n9592), .Z(n9594) );
  XOR U11784 ( .A(n9772), .B(n9773), .Z(n9592) );
  AND U11785 ( .A(n9774), .B(n9775), .Z(n9772) );
  AND U11786 ( .A(a[63]), .B(b[12]), .Z(n9771) );
  XOR U11787 ( .A(n9776), .B(n9597), .Z(n9599) );
  XOR U11788 ( .A(n9777), .B(n9778), .Z(n9597) );
  AND U11789 ( .A(n9779), .B(n9780), .Z(n9777) );
  AND U11790 ( .A(a[64]), .B(b[11]), .Z(n9776) );
  XOR U11791 ( .A(n9781), .B(n9602), .Z(n9604) );
  XOR U11792 ( .A(n9782), .B(n9783), .Z(n9602) );
  AND U11793 ( .A(n9784), .B(n9785), .Z(n9782) );
  AND U11794 ( .A(a[65]), .B(b[10]), .Z(n9781) );
  XOR U11795 ( .A(n9786), .B(n9607), .Z(n9609) );
  XOR U11796 ( .A(n9787), .B(n9788), .Z(n9607) );
  AND U11797 ( .A(n9789), .B(n9790), .Z(n9787) );
  AND U11798 ( .A(a[66]), .B(b[9]), .Z(n9786) );
  XOR U11799 ( .A(n9791), .B(n9792), .Z(n9611) );
  AND U11800 ( .A(n9793), .B(n9794), .Z(n9791) );
  XOR U11801 ( .A(n9795), .B(n9616), .Z(n9618) );
  XOR U11802 ( .A(n9796), .B(n9797), .Z(n9616) );
  AND U11803 ( .A(n9798), .B(n9799), .Z(n9796) );
  AND U11804 ( .A(a[67]), .B(b[8]), .Z(n9795) );
  XOR U11805 ( .A(n9801), .B(n9802), .Z(n9621) );
  AND U11806 ( .A(n9803), .B(n9804), .Z(n9801) );
  AND U11807 ( .A(a[69]), .B(b[6]), .Z(n9800) );
  XOR U11808 ( .A(n9806), .B(n9807), .Z(n9626) );
  AND U11809 ( .A(n9808), .B(n9809), .Z(n9806) );
  AND U11810 ( .A(a[70]), .B(b[5]), .Z(n9805) );
  XOR U11811 ( .A(n9811), .B(n9812), .Z(n9631) );
  AND U11812 ( .A(n9813), .B(n9814), .Z(n9811) );
  AND U11813 ( .A(a[71]), .B(b[4]), .Z(n9810) );
  XOR U11814 ( .A(n9816), .B(n9817), .Z(n9636) );
  AND U11815 ( .A(n9818), .B(n9819), .Z(n9816) );
  AND U11816 ( .A(a[72]), .B(b[3]), .Z(n9815) );
  XOR U11817 ( .A(n9821), .B(n9822), .Z(n9641) );
  OR U11818 ( .A(n9823), .B(n9824), .Z(n9822) );
  AND U11819 ( .A(a[73]), .B(b[2]), .Z(n9820) );
  XNOR U11820 ( .A(n9651), .B(n9825), .Z(n9647) );
  NAND U11821 ( .A(a[74]), .B(b[1]), .Z(n9825) );
  IV U11822 ( .A(n9645), .Z(n9651) );
  ANDN U11823 ( .B(n5182), .A(n5184), .Z(n9645) );
  NAND U11824 ( .A(a[74]), .B(b[0]), .Z(n5184) );
  XOR U11825 ( .A(n9823), .B(n9824), .Z(n5182) );
  XOR U11826 ( .A(n9827), .B(n9818), .Z(n9826) );
  XOR U11827 ( .A(n9813), .B(n9817), .Z(n9828) );
  XOR U11828 ( .A(n9808), .B(n9812), .Z(n9829) );
  XOR U11829 ( .A(n9803), .B(n9807), .Z(n9830) );
  XOR U11830 ( .A(n9793), .B(n9802), .Z(n9831) );
  XOR U11831 ( .A(n9832), .B(n9792), .Z(n9793) );
  AND U11832 ( .A(b[6]), .B(a[68]), .Z(n9832) );
  XNOR U11833 ( .A(n9792), .B(n9798), .Z(n9833) );
  XNOR U11834 ( .A(n9797), .B(n9789), .Z(n9834) );
  XNOR U11835 ( .A(n9788), .B(n9784), .Z(n9835) );
  XNOR U11836 ( .A(n9783), .B(n9779), .Z(n9836) );
  XNOR U11837 ( .A(n9778), .B(n9774), .Z(n9837) );
  XNOR U11838 ( .A(n9773), .B(n9769), .Z(n9838) );
  XNOR U11839 ( .A(n9768), .B(n9764), .Z(n9839) );
  XNOR U11840 ( .A(n9763), .B(n9759), .Z(n9840) );
  XNOR U11841 ( .A(n9758), .B(n9754), .Z(n9841) );
  XNOR U11842 ( .A(n9753), .B(n9749), .Z(n9842) );
  XNOR U11843 ( .A(n9748), .B(n9744), .Z(n9843) );
  XNOR U11844 ( .A(n9743), .B(n9739), .Z(n9844) );
  XNOR U11845 ( .A(n9738), .B(n9734), .Z(n9845) );
  XNOR U11846 ( .A(n9733), .B(n9729), .Z(n9846) );
  XNOR U11847 ( .A(n9728), .B(n9724), .Z(n9847) );
  XNOR U11848 ( .A(n9723), .B(n9719), .Z(n9848) );
  XNOR U11849 ( .A(n9718), .B(n9714), .Z(n9849) );
  XNOR U11850 ( .A(n9713), .B(n9709), .Z(n9850) );
  XNOR U11851 ( .A(n9708), .B(n9704), .Z(n9851) );
  XNOR U11852 ( .A(n9703), .B(n9699), .Z(n9852) );
  XNOR U11853 ( .A(n9698), .B(n9694), .Z(n9853) );
  XOR U11854 ( .A(n9693), .B(n9690), .Z(n9854) );
  XOR U11855 ( .A(n9855), .B(n9856), .Z(n9690) );
  XOR U11856 ( .A(n9688), .B(n9857), .Z(n9856) );
  XOR U11857 ( .A(n9858), .B(n9859), .Z(n9857) );
  XOR U11858 ( .A(n9860), .B(n9861), .Z(n9859) );
  NAND U11859 ( .A(a[44]), .B(b[30]), .Z(n9861) );
  AND U11860 ( .A(a[43]), .B(b[31]), .Z(n9860) );
  XOR U11861 ( .A(n9862), .B(n9858), .Z(n9855) );
  XOR U11862 ( .A(n9863), .B(n9864), .Z(n9858) );
  ANDN U11863 ( .B(n9865), .A(n9866), .Z(n9863) );
  AND U11864 ( .A(a[45]), .B(b[29]), .Z(n9862) );
  XOR U11865 ( .A(n9867), .B(n9688), .Z(n9689) );
  XOR U11866 ( .A(n9868), .B(n9869), .Z(n9688) );
  AND U11867 ( .A(n9870), .B(n9871), .Z(n9868) );
  AND U11868 ( .A(a[46]), .B(b[28]), .Z(n9867) );
  XOR U11869 ( .A(n9872), .B(n9693), .Z(n9695) );
  XOR U11870 ( .A(n9873), .B(n9874), .Z(n9693) );
  AND U11871 ( .A(n9875), .B(n9876), .Z(n9873) );
  AND U11872 ( .A(a[47]), .B(b[27]), .Z(n9872) );
  XOR U11873 ( .A(n9877), .B(n9698), .Z(n9700) );
  XOR U11874 ( .A(n9878), .B(n9879), .Z(n9698) );
  AND U11875 ( .A(n9880), .B(n9881), .Z(n9878) );
  AND U11876 ( .A(a[48]), .B(b[26]), .Z(n9877) );
  XOR U11877 ( .A(n9882), .B(n9703), .Z(n9705) );
  XOR U11878 ( .A(n9883), .B(n9884), .Z(n9703) );
  AND U11879 ( .A(n9885), .B(n9886), .Z(n9883) );
  AND U11880 ( .A(a[49]), .B(b[25]), .Z(n9882) );
  XOR U11881 ( .A(n9887), .B(n9708), .Z(n9710) );
  XOR U11882 ( .A(n9888), .B(n9889), .Z(n9708) );
  AND U11883 ( .A(n9890), .B(n9891), .Z(n9888) );
  AND U11884 ( .A(a[50]), .B(b[24]), .Z(n9887) );
  XOR U11885 ( .A(n9892), .B(n9713), .Z(n9715) );
  XOR U11886 ( .A(n9893), .B(n9894), .Z(n9713) );
  AND U11887 ( .A(n9895), .B(n9896), .Z(n9893) );
  AND U11888 ( .A(a[51]), .B(b[23]), .Z(n9892) );
  XOR U11889 ( .A(n9897), .B(n9718), .Z(n9720) );
  XOR U11890 ( .A(n9898), .B(n9899), .Z(n9718) );
  AND U11891 ( .A(n9900), .B(n9901), .Z(n9898) );
  AND U11892 ( .A(a[52]), .B(b[22]), .Z(n9897) );
  XOR U11893 ( .A(n9902), .B(n9723), .Z(n9725) );
  XOR U11894 ( .A(n9903), .B(n9904), .Z(n9723) );
  AND U11895 ( .A(n9905), .B(n9906), .Z(n9903) );
  AND U11896 ( .A(a[53]), .B(b[21]), .Z(n9902) );
  XOR U11897 ( .A(n9907), .B(n9728), .Z(n9730) );
  XOR U11898 ( .A(n9908), .B(n9909), .Z(n9728) );
  AND U11899 ( .A(n9910), .B(n9911), .Z(n9908) );
  AND U11900 ( .A(a[54]), .B(b[20]), .Z(n9907) );
  XOR U11901 ( .A(n9912), .B(n9733), .Z(n9735) );
  XOR U11902 ( .A(n9913), .B(n9914), .Z(n9733) );
  AND U11903 ( .A(n9915), .B(n9916), .Z(n9913) );
  AND U11904 ( .A(a[55]), .B(b[19]), .Z(n9912) );
  XOR U11905 ( .A(n9917), .B(n9738), .Z(n9740) );
  XOR U11906 ( .A(n9918), .B(n9919), .Z(n9738) );
  AND U11907 ( .A(n9920), .B(n9921), .Z(n9918) );
  AND U11908 ( .A(a[56]), .B(b[18]), .Z(n9917) );
  XOR U11909 ( .A(n9922), .B(n9743), .Z(n9745) );
  XOR U11910 ( .A(n9923), .B(n9924), .Z(n9743) );
  AND U11911 ( .A(n9925), .B(n9926), .Z(n9923) );
  AND U11912 ( .A(a[57]), .B(b[17]), .Z(n9922) );
  XOR U11913 ( .A(n9927), .B(n9748), .Z(n9750) );
  XOR U11914 ( .A(n9928), .B(n9929), .Z(n9748) );
  AND U11915 ( .A(n9930), .B(n9931), .Z(n9928) );
  AND U11916 ( .A(a[58]), .B(b[16]), .Z(n9927) );
  XOR U11917 ( .A(n9932), .B(n9753), .Z(n9755) );
  XOR U11918 ( .A(n9933), .B(n9934), .Z(n9753) );
  AND U11919 ( .A(n9935), .B(n9936), .Z(n9933) );
  AND U11920 ( .A(a[59]), .B(b[15]), .Z(n9932) );
  XOR U11921 ( .A(n9937), .B(n9758), .Z(n9760) );
  XOR U11922 ( .A(n9938), .B(n9939), .Z(n9758) );
  AND U11923 ( .A(n9940), .B(n9941), .Z(n9938) );
  AND U11924 ( .A(a[60]), .B(b[14]), .Z(n9937) );
  XOR U11925 ( .A(n9942), .B(n9763), .Z(n9765) );
  XOR U11926 ( .A(n9943), .B(n9944), .Z(n9763) );
  AND U11927 ( .A(n9945), .B(n9946), .Z(n9943) );
  AND U11928 ( .A(a[61]), .B(b[13]), .Z(n9942) );
  XOR U11929 ( .A(n9947), .B(n9768), .Z(n9770) );
  XOR U11930 ( .A(n9948), .B(n9949), .Z(n9768) );
  AND U11931 ( .A(n9950), .B(n9951), .Z(n9948) );
  AND U11932 ( .A(a[62]), .B(b[12]), .Z(n9947) );
  XOR U11933 ( .A(n9952), .B(n9773), .Z(n9775) );
  XOR U11934 ( .A(n9953), .B(n9954), .Z(n9773) );
  AND U11935 ( .A(n9955), .B(n9956), .Z(n9953) );
  AND U11936 ( .A(a[63]), .B(b[11]), .Z(n9952) );
  XOR U11937 ( .A(n9957), .B(n9778), .Z(n9780) );
  XOR U11938 ( .A(n9958), .B(n9959), .Z(n9778) );
  AND U11939 ( .A(n9960), .B(n9961), .Z(n9958) );
  AND U11940 ( .A(a[64]), .B(b[10]), .Z(n9957) );
  XOR U11941 ( .A(n9962), .B(n9783), .Z(n9785) );
  XOR U11942 ( .A(n9963), .B(n9964), .Z(n9783) );
  AND U11943 ( .A(n9965), .B(n9966), .Z(n9963) );
  AND U11944 ( .A(a[65]), .B(b[9]), .Z(n9962) );
  XOR U11945 ( .A(n9967), .B(n9788), .Z(n9790) );
  XOR U11946 ( .A(n9968), .B(n9969), .Z(n9788) );
  AND U11947 ( .A(n9970), .B(n9971), .Z(n9968) );
  AND U11948 ( .A(a[66]), .B(b[8]), .Z(n9967) );
  XOR U11949 ( .A(n9972), .B(n9973), .Z(n9792) );
  AND U11950 ( .A(n9974), .B(n9975), .Z(n9972) );
  XOR U11951 ( .A(n9976), .B(n9797), .Z(n9799) );
  XOR U11952 ( .A(n9977), .B(n9978), .Z(n9797) );
  AND U11953 ( .A(n9979), .B(n9980), .Z(n9977) );
  AND U11954 ( .A(a[67]), .B(b[7]), .Z(n9976) );
  XOR U11955 ( .A(n9982), .B(n9983), .Z(n9802) );
  AND U11956 ( .A(n9984), .B(n9985), .Z(n9982) );
  AND U11957 ( .A(a[69]), .B(b[5]), .Z(n9981) );
  XOR U11958 ( .A(n9987), .B(n9988), .Z(n9807) );
  AND U11959 ( .A(n9989), .B(n9990), .Z(n9987) );
  AND U11960 ( .A(a[70]), .B(b[4]), .Z(n9986) );
  XOR U11961 ( .A(n9992), .B(n9993), .Z(n9812) );
  AND U11962 ( .A(n9994), .B(n9995), .Z(n9992) );
  AND U11963 ( .A(a[71]), .B(b[3]), .Z(n9991) );
  XOR U11964 ( .A(n9997), .B(n9998), .Z(n9817) );
  OR U11965 ( .A(n9999), .B(n10000), .Z(n9998) );
  AND U11966 ( .A(a[72]), .B(b[2]), .Z(n9996) );
  XNOR U11967 ( .A(n9827), .B(n10001), .Z(n9823) );
  NAND U11968 ( .A(a[73]), .B(b[1]), .Z(n10001) );
  IV U11969 ( .A(n9821), .Z(n9827) );
  ANDN U11970 ( .B(n5187), .A(n5189), .Z(n9821) );
  NAND U11971 ( .A(a[73]), .B(b[0]), .Z(n5189) );
  XOR U11972 ( .A(n9999), .B(n10000), .Z(n5187) );
  XOR U11973 ( .A(n10003), .B(n9994), .Z(n10002) );
  XOR U11974 ( .A(n9989), .B(n9993), .Z(n10004) );
  XOR U11975 ( .A(n9984), .B(n9988), .Z(n10005) );
  XOR U11976 ( .A(n9974), .B(n9983), .Z(n10006) );
  XOR U11977 ( .A(n10007), .B(n9973), .Z(n9974) );
  AND U11978 ( .A(b[5]), .B(a[68]), .Z(n10007) );
  XNOR U11979 ( .A(n9973), .B(n9979), .Z(n10008) );
  XNOR U11980 ( .A(n9978), .B(n9970), .Z(n10009) );
  XNOR U11981 ( .A(n9969), .B(n9965), .Z(n10010) );
  XNOR U11982 ( .A(n9964), .B(n9960), .Z(n10011) );
  XNOR U11983 ( .A(n9959), .B(n9955), .Z(n10012) );
  XNOR U11984 ( .A(n9954), .B(n9950), .Z(n10013) );
  XNOR U11985 ( .A(n9949), .B(n9945), .Z(n10014) );
  XNOR U11986 ( .A(n9944), .B(n9940), .Z(n10015) );
  XNOR U11987 ( .A(n9939), .B(n9935), .Z(n10016) );
  XNOR U11988 ( .A(n9934), .B(n9930), .Z(n10017) );
  XNOR U11989 ( .A(n9929), .B(n9925), .Z(n10018) );
  XNOR U11990 ( .A(n9924), .B(n9920), .Z(n10019) );
  XNOR U11991 ( .A(n9919), .B(n9915), .Z(n10020) );
  XNOR U11992 ( .A(n9914), .B(n9910), .Z(n10021) );
  XNOR U11993 ( .A(n9909), .B(n9905), .Z(n10022) );
  XNOR U11994 ( .A(n9904), .B(n9900), .Z(n10023) );
  XNOR U11995 ( .A(n9899), .B(n9895), .Z(n10024) );
  XNOR U11996 ( .A(n9894), .B(n9890), .Z(n10025) );
  XNOR U11997 ( .A(n9889), .B(n9885), .Z(n10026) );
  XNOR U11998 ( .A(n9884), .B(n9880), .Z(n10027) );
  XNOR U11999 ( .A(n9879), .B(n9875), .Z(n10028) );
  XNOR U12000 ( .A(n9874), .B(n9870), .Z(n10029) );
  XOR U12001 ( .A(n9869), .B(n9866), .Z(n10030) );
  XOR U12002 ( .A(n10031), .B(n10032), .Z(n9866) );
  XOR U12003 ( .A(n9864), .B(n10033), .Z(n10032) );
  XOR U12004 ( .A(n10034), .B(n10035), .Z(n10033) );
  XOR U12005 ( .A(n10036), .B(n10037), .Z(n10035) );
  NAND U12006 ( .A(a[43]), .B(b[30]), .Z(n10037) );
  AND U12007 ( .A(a[42]), .B(b[31]), .Z(n10036) );
  XOR U12008 ( .A(n10038), .B(n10034), .Z(n10031) );
  XOR U12009 ( .A(n10039), .B(n10040), .Z(n10034) );
  ANDN U12010 ( .B(n10041), .A(n10042), .Z(n10039) );
  AND U12011 ( .A(a[44]), .B(b[29]), .Z(n10038) );
  XOR U12012 ( .A(n10043), .B(n9864), .Z(n9865) );
  XOR U12013 ( .A(n10044), .B(n10045), .Z(n9864) );
  AND U12014 ( .A(n10046), .B(n10047), .Z(n10044) );
  AND U12015 ( .A(a[45]), .B(b[28]), .Z(n10043) );
  XOR U12016 ( .A(n10048), .B(n9869), .Z(n9871) );
  XOR U12017 ( .A(n10049), .B(n10050), .Z(n9869) );
  AND U12018 ( .A(n10051), .B(n10052), .Z(n10049) );
  AND U12019 ( .A(a[46]), .B(b[27]), .Z(n10048) );
  XOR U12020 ( .A(n10053), .B(n9874), .Z(n9876) );
  XOR U12021 ( .A(n10054), .B(n10055), .Z(n9874) );
  AND U12022 ( .A(n10056), .B(n10057), .Z(n10054) );
  AND U12023 ( .A(a[47]), .B(b[26]), .Z(n10053) );
  XOR U12024 ( .A(n10058), .B(n9879), .Z(n9881) );
  XOR U12025 ( .A(n10059), .B(n10060), .Z(n9879) );
  AND U12026 ( .A(n10061), .B(n10062), .Z(n10059) );
  AND U12027 ( .A(a[48]), .B(b[25]), .Z(n10058) );
  XOR U12028 ( .A(n10063), .B(n9884), .Z(n9886) );
  XOR U12029 ( .A(n10064), .B(n10065), .Z(n9884) );
  AND U12030 ( .A(n10066), .B(n10067), .Z(n10064) );
  AND U12031 ( .A(a[49]), .B(b[24]), .Z(n10063) );
  XOR U12032 ( .A(n10068), .B(n9889), .Z(n9891) );
  XOR U12033 ( .A(n10069), .B(n10070), .Z(n9889) );
  AND U12034 ( .A(n10071), .B(n10072), .Z(n10069) );
  AND U12035 ( .A(a[50]), .B(b[23]), .Z(n10068) );
  XOR U12036 ( .A(n10073), .B(n9894), .Z(n9896) );
  XOR U12037 ( .A(n10074), .B(n10075), .Z(n9894) );
  AND U12038 ( .A(n10076), .B(n10077), .Z(n10074) );
  AND U12039 ( .A(a[51]), .B(b[22]), .Z(n10073) );
  XOR U12040 ( .A(n10078), .B(n9899), .Z(n9901) );
  XOR U12041 ( .A(n10079), .B(n10080), .Z(n9899) );
  AND U12042 ( .A(n10081), .B(n10082), .Z(n10079) );
  AND U12043 ( .A(a[52]), .B(b[21]), .Z(n10078) );
  XOR U12044 ( .A(n10083), .B(n9904), .Z(n9906) );
  XOR U12045 ( .A(n10084), .B(n10085), .Z(n9904) );
  AND U12046 ( .A(n10086), .B(n10087), .Z(n10084) );
  AND U12047 ( .A(a[53]), .B(b[20]), .Z(n10083) );
  XOR U12048 ( .A(n10088), .B(n9909), .Z(n9911) );
  XOR U12049 ( .A(n10089), .B(n10090), .Z(n9909) );
  AND U12050 ( .A(n10091), .B(n10092), .Z(n10089) );
  AND U12051 ( .A(a[54]), .B(b[19]), .Z(n10088) );
  XOR U12052 ( .A(n10093), .B(n9914), .Z(n9916) );
  XOR U12053 ( .A(n10094), .B(n10095), .Z(n9914) );
  AND U12054 ( .A(n10096), .B(n10097), .Z(n10094) );
  AND U12055 ( .A(a[55]), .B(b[18]), .Z(n10093) );
  XOR U12056 ( .A(n10098), .B(n9919), .Z(n9921) );
  XOR U12057 ( .A(n10099), .B(n10100), .Z(n9919) );
  AND U12058 ( .A(n10101), .B(n10102), .Z(n10099) );
  AND U12059 ( .A(a[56]), .B(b[17]), .Z(n10098) );
  XOR U12060 ( .A(n10103), .B(n9924), .Z(n9926) );
  XOR U12061 ( .A(n10104), .B(n10105), .Z(n9924) );
  AND U12062 ( .A(n10106), .B(n10107), .Z(n10104) );
  AND U12063 ( .A(a[57]), .B(b[16]), .Z(n10103) );
  XOR U12064 ( .A(n10108), .B(n9929), .Z(n9931) );
  XOR U12065 ( .A(n10109), .B(n10110), .Z(n9929) );
  AND U12066 ( .A(n10111), .B(n10112), .Z(n10109) );
  AND U12067 ( .A(a[58]), .B(b[15]), .Z(n10108) );
  XOR U12068 ( .A(n10113), .B(n9934), .Z(n9936) );
  XOR U12069 ( .A(n10114), .B(n10115), .Z(n9934) );
  AND U12070 ( .A(n10116), .B(n10117), .Z(n10114) );
  AND U12071 ( .A(a[59]), .B(b[14]), .Z(n10113) );
  XOR U12072 ( .A(n10118), .B(n9939), .Z(n9941) );
  XOR U12073 ( .A(n10119), .B(n10120), .Z(n9939) );
  AND U12074 ( .A(n10121), .B(n10122), .Z(n10119) );
  AND U12075 ( .A(a[60]), .B(b[13]), .Z(n10118) );
  XOR U12076 ( .A(n10123), .B(n9944), .Z(n9946) );
  XOR U12077 ( .A(n10124), .B(n10125), .Z(n9944) );
  AND U12078 ( .A(n10126), .B(n10127), .Z(n10124) );
  AND U12079 ( .A(a[61]), .B(b[12]), .Z(n10123) );
  XOR U12080 ( .A(n10128), .B(n9949), .Z(n9951) );
  XOR U12081 ( .A(n10129), .B(n10130), .Z(n9949) );
  AND U12082 ( .A(n10131), .B(n10132), .Z(n10129) );
  AND U12083 ( .A(a[62]), .B(b[11]), .Z(n10128) );
  XOR U12084 ( .A(n10133), .B(n9954), .Z(n9956) );
  XOR U12085 ( .A(n10134), .B(n10135), .Z(n9954) );
  AND U12086 ( .A(n10136), .B(n10137), .Z(n10134) );
  AND U12087 ( .A(a[63]), .B(b[10]), .Z(n10133) );
  XOR U12088 ( .A(n10138), .B(n9959), .Z(n9961) );
  XOR U12089 ( .A(n10139), .B(n10140), .Z(n9959) );
  AND U12090 ( .A(n10141), .B(n10142), .Z(n10139) );
  AND U12091 ( .A(a[64]), .B(b[9]), .Z(n10138) );
  XOR U12092 ( .A(n10143), .B(n9964), .Z(n9966) );
  XOR U12093 ( .A(n10144), .B(n10145), .Z(n9964) );
  AND U12094 ( .A(n10146), .B(n10147), .Z(n10144) );
  AND U12095 ( .A(a[65]), .B(b[8]), .Z(n10143) );
  XOR U12096 ( .A(n10148), .B(n9969), .Z(n9971) );
  XOR U12097 ( .A(n10149), .B(n10150), .Z(n9969) );
  AND U12098 ( .A(n10151), .B(n10152), .Z(n10149) );
  AND U12099 ( .A(a[66]), .B(b[7]), .Z(n10148) );
  XOR U12100 ( .A(n10153), .B(n10154), .Z(n9973) );
  AND U12101 ( .A(n10155), .B(n10156), .Z(n10153) );
  XOR U12102 ( .A(n10157), .B(n9978), .Z(n9980) );
  XOR U12103 ( .A(n10158), .B(n10159), .Z(n9978) );
  AND U12104 ( .A(n10160), .B(n10161), .Z(n10158) );
  AND U12105 ( .A(a[67]), .B(b[6]), .Z(n10157) );
  XOR U12106 ( .A(n10163), .B(n10164), .Z(n9983) );
  AND U12107 ( .A(n10165), .B(n10166), .Z(n10163) );
  AND U12108 ( .A(a[69]), .B(b[4]), .Z(n10162) );
  XOR U12109 ( .A(n10168), .B(n10169), .Z(n9988) );
  AND U12110 ( .A(n10170), .B(n10171), .Z(n10168) );
  AND U12111 ( .A(a[70]), .B(b[3]), .Z(n10167) );
  XOR U12112 ( .A(n10173), .B(n10174), .Z(n9993) );
  OR U12113 ( .A(n10175), .B(n10176), .Z(n10174) );
  AND U12114 ( .A(a[71]), .B(b[2]), .Z(n10172) );
  XNOR U12115 ( .A(n10003), .B(n10177), .Z(n9999) );
  NAND U12116 ( .A(a[72]), .B(b[1]), .Z(n10177) );
  IV U12117 ( .A(n9997), .Z(n10003) );
  ANDN U12118 ( .B(n5192), .A(n5194), .Z(n9997) );
  NAND U12119 ( .A(a[72]), .B(b[0]), .Z(n5194) );
  XOR U12120 ( .A(n10175), .B(n10176), .Z(n5192) );
  XOR U12121 ( .A(n10179), .B(n10170), .Z(n10178) );
  XOR U12122 ( .A(n10165), .B(n10169), .Z(n10180) );
  XOR U12123 ( .A(n10155), .B(n10164), .Z(n10181) );
  XOR U12124 ( .A(n10182), .B(n10154), .Z(n10155) );
  AND U12125 ( .A(b[4]), .B(a[68]), .Z(n10182) );
  XNOR U12126 ( .A(n10154), .B(n10160), .Z(n10183) );
  XNOR U12127 ( .A(n10159), .B(n10151), .Z(n10184) );
  XNOR U12128 ( .A(n10150), .B(n10146), .Z(n10185) );
  XNOR U12129 ( .A(n10145), .B(n10141), .Z(n10186) );
  XNOR U12130 ( .A(n10140), .B(n10136), .Z(n10187) );
  XNOR U12131 ( .A(n10135), .B(n10131), .Z(n10188) );
  XNOR U12132 ( .A(n10130), .B(n10126), .Z(n10189) );
  XNOR U12133 ( .A(n10125), .B(n10121), .Z(n10190) );
  XNOR U12134 ( .A(n10120), .B(n10116), .Z(n10191) );
  XNOR U12135 ( .A(n10115), .B(n10111), .Z(n10192) );
  XNOR U12136 ( .A(n10110), .B(n10106), .Z(n10193) );
  XNOR U12137 ( .A(n10105), .B(n10101), .Z(n10194) );
  XNOR U12138 ( .A(n10100), .B(n10096), .Z(n10195) );
  XNOR U12139 ( .A(n10095), .B(n10091), .Z(n10196) );
  XNOR U12140 ( .A(n10090), .B(n10086), .Z(n10197) );
  XNOR U12141 ( .A(n10085), .B(n10081), .Z(n10198) );
  XNOR U12142 ( .A(n10080), .B(n10076), .Z(n10199) );
  XNOR U12143 ( .A(n10075), .B(n10071), .Z(n10200) );
  XNOR U12144 ( .A(n10070), .B(n10066), .Z(n10201) );
  XNOR U12145 ( .A(n10065), .B(n10061), .Z(n10202) );
  XNOR U12146 ( .A(n10060), .B(n10056), .Z(n10203) );
  XNOR U12147 ( .A(n10055), .B(n10051), .Z(n10204) );
  XNOR U12148 ( .A(n10050), .B(n10046), .Z(n10205) );
  XOR U12149 ( .A(n10045), .B(n10042), .Z(n10206) );
  XOR U12150 ( .A(n10207), .B(n10208), .Z(n10042) );
  XOR U12151 ( .A(n10040), .B(n10209), .Z(n10208) );
  XOR U12152 ( .A(n10210), .B(n10211), .Z(n10209) );
  XOR U12153 ( .A(n10212), .B(n10213), .Z(n10211) );
  NAND U12154 ( .A(a[42]), .B(b[30]), .Z(n10213) );
  AND U12155 ( .A(a[41]), .B(b[31]), .Z(n10212) );
  XOR U12156 ( .A(n10214), .B(n10210), .Z(n10207) );
  XOR U12157 ( .A(n10215), .B(n10216), .Z(n10210) );
  ANDN U12158 ( .B(n10217), .A(n10218), .Z(n10215) );
  AND U12159 ( .A(a[43]), .B(b[29]), .Z(n10214) );
  XOR U12160 ( .A(n10219), .B(n10040), .Z(n10041) );
  XOR U12161 ( .A(n10220), .B(n10221), .Z(n10040) );
  AND U12162 ( .A(n10222), .B(n10223), .Z(n10220) );
  AND U12163 ( .A(a[44]), .B(b[28]), .Z(n10219) );
  XOR U12164 ( .A(n10224), .B(n10045), .Z(n10047) );
  XOR U12165 ( .A(n10225), .B(n10226), .Z(n10045) );
  AND U12166 ( .A(n10227), .B(n10228), .Z(n10225) );
  AND U12167 ( .A(a[45]), .B(b[27]), .Z(n10224) );
  XOR U12168 ( .A(n10229), .B(n10050), .Z(n10052) );
  XOR U12169 ( .A(n10230), .B(n10231), .Z(n10050) );
  AND U12170 ( .A(n10232), .B(n10233), .Z(n10230) );
  AND U12171 ( .A(a[46]), .B(b[26]), .Z(n10229) );
  XOR U12172 ( .A(n10234), .B(n10055), .Z(n10057) );
  XOR U12173 ( .A(n10235), .B(n10236), .Z(n10055) );
  AND U12174 ( .A(n10237), .B(n10238), .Z(n10235) );
  AND U12175 ( .A(a[47]), .B(b[25]), .Z(n10234) );
  XOR U12176 ( .A(n10239), .B(n10060), .Z(n10062) );
  XOR U12177 ( .A(n10240), .B(n10241), .Z(n10060) );
  AND U12178 ( .A(n10242), .B(n10243), .Z(n10240) );
  AND U12179 ( .A(a[48]), .B(b[24]), .Z(n10239) );
  XOR U12180 ( .A(n10244), .B(n10065), .Z(n10067) );
  XOR U12181 ( .A(n10245), .B(n10246), .Z(n10065) );
  AND U12182 ( .A(n10247), .B(n10248), .Z(n10245) );
  AND U12183 ( .A(a[49]), .B(b[23]), .Z(n10244) );
  XOR U12184 ( .A(n10249), .B(n10070), .Z(n10072) );
  XOR U12185 ( .A(n10250), .B(n10251), .Z(n10070) );
  AND U12186 ( .A(n10252), .B(n10253), .Z(n10250) );
  AND U12187 ( .A(a[50]), .B(b[22]), .Z(n10249) );
  XOR U12188 ( .A(n10254), .B(n10075), .Z(n10077) );
  XOR U12189 ( .A(n10255), .B(n10256), .Z(n10075) );
  AND U12190 ( .A(n10257), .B(n10258), .Z(n10255) );
  AND U12191 ( .A(a[51]), .B(b[21]), .Z(n10254) );
  XOR U12192 ( .A(n10259), .B(n10080), .Z(n10082) );
  XOR U12193 ( .A(n10260), .B(n10261), .Z(n10080) );
  AND U12194 ( .A(n10262), .B(n10263), .Z(n10260) );
  AND U12195 ( .A(a[52]), .B(b[20]), .Z(n10259) );
  XOR U12196 ( .A(n10264), .B(n10085), .Z(n10087) );
  XOR U12197 ( .A(n10265), .B(n10266), .Z(n10085) );
  AND U12198 ( .A(n10267), .B(n10268), .Z(n10265) );
  AND U12199 ( .A(a[53]), .B(b[19]), .Z(n10264) );
  XOR U12200 ( .A(n10269), .B(n10090), .Z(n10092) );
  XOR U12201 ( .A(n10270), .B(n10271), .Z(n10090) );
  AND U12202 ( .A(n10272), .B(n10273), .Z(n10270) );
  AND U12203 ( .A(a[54]), .B(b[18]), .Z(n10269) );
  XOR U12204 ( .A(n10274), .B(n10095), .Z(n10097) );
  XOR U12205 ( .A(n10275), .B(n10276), .Z(n10095) );
  AND U12206 ( .A(n10277), .B(n10278), .Z(n10275) );
  AND U12207 ( .A(a[55]), .B(b[17]), .Z(n10274) );
  XOR U12208 ( .A(n10279), .B(n10100), .Z(n10102) );
  XOR U12209 ( .A(n10280), .B(n10281), .Z(n10100) );
  AND U12210 ( .A(n10282), .B(n10283), .Z(n10280) );
  AND U12211 ( .A(a[56]), .B(b[16]), .Z(n10279) );
  XOR U12212 ( .A(n10284), .B(n10105), .Z(n10107) );
  XOR U12213 ( .A(n10285), .B(n10286), .Z(n10105) );
  AND U12214 ( .A(n10287), .B(n10288), .Z(n10285) );
  AND U12215 ( .A(a[57]), .B(b[15]), .Z(n10284) );
  XOR U12216 ( .A(n10289), .B(n10110), .Z(n10112) );
  XOR U12217 ( .A(n10290), .B(n10291), .Z(n10110) );
  AND U12218 ( .A(n10292), .B(n10293), .Z(n10290) );
  AND U12219 ( .A(a[58]), .B(b[14]), .Z(n10289) );
  XOR U12220 ( .A(n10294), .B(n10115), .Z(n10117) );
  XOR U12221 ( .A(n10295), .B(n10296), .Z(n10115) );
  AND U12222 ( .A(n10297), .B(n10298), .Z(n10295) );
  AND U12223 ( .A(a[59]), .B(b[13]), .Z(n10294) );
  XOR U12224 ( .A(n10299), .B(n10120), .Z(n10122) );
  XOR U12225 ( .A(n10300), .B(n10301), .Z(n10120) );
  AND U12226 ( .A(n10302), .B(n10303), .Z(n10300) );
  AND U12227 ( .A(a[60]), .B(b[12]), .Z(n10299) );
  XOR U12228 ( .A(n10304), .B(n10125), .Z(n10127) );
  XOR U12229 ( .A(n10305), .B(n10306), .Z(n10125) );
  AND U12230 ( .A(n10307), .B(n10308), .Z(n10305) );
  AND U12231 ( .A(a[61]), .B(b[11]), .Z(n10304) );
  XOR U12232 ( .A(n10309), .B(n10130), .Z(n10132) );
  XOR U12233 ( .A(n10310), .B(n10311), .Z(n10130) );
  AND U12234 ( .A(n10312), .B(n10313), .Z(n10310) );
  AND U12235 ( .A(a[62]), .B(b[10]), .Z(n10309) );
  XOR U12236 ( .A(n10314), .B(n10135), .Z(n10137) );
  XOR U12237 ( .A(n10315), .B(n10316), .Z(n10135) );
  AND U12238 ( .A(n10317), .B(n10318), .Z(n10315) );
  AND U12239 ( .A(a[63]), .B(b[9]), .Z(n10314) );
  XOR U12240 ( .A(n10319), .B(n10140), .Z(n10142) );
  XOR U12241 ( .A(n10320), .B(n10321), .Z(n10140) );
  AND U12242 ( .A(n10322), .B(n10323), .Z(n10320) );
  AND U12243 ( .A(a[64]), .B(b[8]), .Z(n10319) );
  XOR U12244 ( .A(n10324), .B(n10145), .Z(n10147) );
  XOR U12245 ( .A(n10325), .B(n10326), .Z(n10145) );
  AND U12246 ( .A(n10327), .B(n10328), .Z(n10325) );
  AND U12247 ( .A(a[65]), .B(b[7]), .Z(n10324) );
  XOR U12248 ( .A(n10329), .B(n10150), .Z(n10152) );
  XOR U12249 ( .A(n10330), .B(n10331), .Z(n10150) );
  AND U12250 ( .A(n10332), .B(n10333), .Z(n10330) );
  AND U12251 ( .A(a[66]), .B(b[6]), .Z(n10329) );
  XOR U12252 ( .A(n10334), .B(n10335), .Z(n10154) );
  AND U12253 ( .A(n10336), .B(n10337), .Z(n10334) );
  XOR U12254 ( .A(n10338), .B(n10159), .Z(n10161) );
  XOR U12255 ( .A(n10339), .B(n10340), .Z(n10159) );
  AND U12256 ( .A(n10341), .B(n10342), .Z(n10339) );
  AND U12257 ( .A(a[67]), .B(b[5]), .Z(n10338) );
  XOR U12258 ( .A(n10344), .B(n10345), .Z(n10164) );
  AND U12259 ( .A(n10346), .B(n10347), .Z(n10344) );
  AND U12260 ( .A(a[69]), .B(b[3]), .Z(n10343) );
  XOR U12261 ( .A(n10349), .B(n10350), .Z(n10169) );
  OR U12262 ( .A(n10351), .B(n10352), .Z(n10350) );
  AND U12263 ( .A(a[70]), .B(b[2]), .Z(n10348) );
  XNOR U12264 ( .A(n10179), .B(n10353), .Z(n10175) );
  NAND U12265 ( .A(a[71]), .B(b[1]), .Z(n10353) );
  IV U12266 ( .A(n10173), .Z(n10179) );
  ANDN U12267 ( .B(n5197), .A(n5199), .Z(n10173) );
  NAND U12268 ( .A(a[71]), .B(b[0]), .Z(n5199) );
  XOR U12269 ( .A(n10351), .B(n10352), .Z(n5197) );
  XOR U12270 ( .A(n10355), .B(n10346), .Z(n10354) );
  XOR U12271 ( .A(n10336), .B(n10345), .Z(n10356) );
  XOR U12272 ( .A(n10357), .B(n10335), .Z(n10336) );
  AND U12273 ( .A(b[3]), .B(a[68]), .Z(n10357) );
  XNOR U12274 ( .A(n10335), .B(n10341), .Z(n10358) );
  XNOR U12275 ( .A(n10340), .B(n10332), .Z(n10359) );
  XNOR U12276 ( .A(n10331), .B(n10327), .Z(n10360) );
  XNOR U12277 ( .A(n10326), .B(n10322), .Z(n10361) );
  XNOR U12278 ( .A(n10321), .B(n10317), .Z(n10362) );
  XNOR U12279 ( .A(n10316), .B(n10312), .Z(n10363) );
  XNOR U12280 ( .A(n10311), .B(n10307), .Z(n10364) );
  XNOR U12281 ( .A(n10306), .B(n10302), .Z(n10365) );
  XNOR U12282 ( .A(n10301), .B(n10297), .Z(n10366) );
  XNOR U12283 ( .A(n10296), .B(n10292), .Z(n10367) );
  XNOR U12284 ( .A(n10291), .B(n10287), .Z(n10368) );
  XNOR U12285 ( .A(n10286), .B(n10282), .Z(n10369) );
  XNOR U12286 ( .A(n10281), .B(n10277), .Z(n10370) );
  XNOR U12287 ( .A(n10276), .B(n10272), .Z(n10371) );
  XNOR U12288 ( .A(n10271), .B(n10267), .Z(n10372) );
  XNOR U12289 ( .A(n10266), .B(n10262), .Z(n10373) );
  XNOR U12290 ( .A(n10261), .B(n10257), .Z(n10374) );
  XNOR U12291 ( .A(n10256), .B(n10252), .Z(n10375) );
  XNOR U12292 ( .A(n10251), .B(n10247), .Z(n10376) );
  XNOR U12293 ( .A(n10246), .B(n10242), .Z(n10377) );
  XNOR U12294 ( .A(n10241), .B(n10237), .Z(n10378) );
  XNOR U12295 ( .A(n10236), .B(n10232), .Z(n10379) );
  XNOR U12296 ( .A(n10231), .B(n10227), .Z(n10380) );
  XNOR U12297 ( .A(n10226), .B(n10222), .Z(n10381) );
  XOR U12298 ( .A(n10221), .B(n10218), .Z(n10382) );
  XOR U12299 ( .A(n10383), .B(n10384), .Z(n10218) );
  XOR U12300 ( .A(n10216), .B(n10385), .Z(n10384) );
  XOR U12301 ( .A(n10386), .B(n10387), .Z(n10385) );
  XOR U12302 ( .A(n10388), .B(n10389), .Z(n10387) );
  NAND U12303 ( .A(a[41]), .B(b[30]), .Z(n10389) );
  AND U12304 ( .A(a[40]), .B(b[31]), .Z(n10388) );
  XOR U12305 ( .A(n10390), .B(n10386), .Z(n10383) );
  XOR U12306 ( .A(n10391), .B(n10392), .Z(n10386) );
  ANDN U12307 ( .B(n10393), .A(n10394), .Z(n10391) );
  AND U12308 ( .A(a[42]), .B(b[29]), .Z(n10390) );
  XOR U12309 ( .A(n10395), .B(n10216), .Z(n10217) );
  XOR U12310 ( .A(n10396), .B(n10397), .Z(n10216) );
  AND U12311 ( .A(n10398), .B(n10399), .Z(n10396) );
  AND U12312 ( .A(a[43]), .B(b[28]), .Z(n10395) );
  XOR U12313 ( .A(n10400), .B(n10221), .Z(n10223) );
  XOR U12314 ( .A(n10401), .B(n10402), .Z(n10221) );
  AND U12315 ( .A(n10403), .B(n10404), .Z(n10401) );
  AND U12316 ( .A(a[44]), .B(b[27]), .Z(n10400) );
  XOR U12317 ( .A(n10405), .B(n10226), .Z(n10228) );
  XOR U12318 ( .A(n10406), .B(n10407), .Z(n10226) );
  AND U12319 ( .A(n10408), .B(n10409), .Z(n10406) );
  AND U12320 ( .A(a[45]), .B(b[26]), .Z(n10405) );
  XOR U12321 ( .A(n10410), .B(n10231), .Z(n10233) );
  XOR U12322 ( .A(n10411), .B(n10412), .Z(n10231) );
  AND U12323 ( .A(n10413), .B(n10414), .Z(n10411) );
  AND U12324 ( .A(a[46]), .B(b[25]), .Z(n10410) );
  XOR U12325 ( .A(n10415), .B(n10236), .Z(n10238) );
  XOR U12326 ( .A(n10416), .B(n10417), .Z(n10236) );
  AND U12327 ( .A(n10418), .B(n10419), .Z(n10416) );
  AND U12328 ( .A(a[47]), .B(b[24]), .Z(n10415) );
  XOR U12329 ( .A(n10420), .B(n10241), .Z(n10243) );
  XOR U12330 ( .A(n10421), .B(n10422), .Z(n10241) );
  AND U12331 ( .A(n10423), .B(n10424), .Z(n10421) );
  AND U12332 ( .A(a[48]), .B(b[23]), .Z(n10420) );
  XOR U12333 ( .A(n10425), .B(n10246), .Z(n10248) );
  XOR U12334 ( .A(n10426), .B(n10427), .Z(n10246) );
  AND U12335 ( .A(n10428), .B(n10429), .Z(n10426) );
  AND U12336 ( .A(a[49]), .B(b[22]), .Z(n10425) );
  XOR U12337 ( .A(n10430), .B(n10251), .Z(n10253) );
  XOR U12338 ( .A(n10431), .B(n10432), .Z(n10251) );
  AND U12339 ( .A(n10433), .B(n10434), .Z(n10431) );
  AND U12340 ( .A(a[50]), .B(b[21]), .Z(n10430) );
  XOR U12341 ( .A(n10435), .B(n10256), .Z(n10258) );
  XOR U12342 ( .A(n10436), .B(n10437), .Z(n10256) );
  AND U12343 ( .A(n10438), .B(n10439), .Z(n10436) );
  AND U12344 ( .A(a[51]), .B(b[20]), .Z(n10435) );
  XOR U12345 ( .A(n10440), .B(n10261), .Z(n10263) );
  XOR U12346 ( .A(n10441), .B(n10442), .Z(n10261) );
  AND U12347 ( .A(n10443), .B(n10444), .Z(n10441) );
  AND U12348 ( .A(a[52]), .B(b[19]), .Z(n10440) );
  XOR U12349 ( .A(n10445), .B(n10266), .Z(n10268) );
  XOR U12350 ( .A(n10446), .B(n10447), .Z(n10266) );
  AND U12351 ( .A(n10448), .B(n10449), .Z(n10446) );
  AND U12352 ( .A(a[53]), .B(b[18]), .Z(n10445) );
  XOR U12353 ( .A(n10450), .B(n10271), .Z(n10273) );
  XOR U12354 ( .A(n10451), .B(n10452), .Z(n10271) );
  AND U12355 ( .A(n10453), .B(n10454), .Z(n10451) );
  AND U12356 ( .A(a[54]), .B(b[17]), .Z(n10450) );
  XOR U12357 ( .A(n10455), .B(n10276), .Z(n10278) );
  XOR U12358 ( .A(n10456), .B(n10457), .Z(n10276) );
  AND U12359 ( .A(n10458), .B(n10459), .Z(n10456) );
  AND U12360 ( .A(a[55]), .B(b[16]), .Z(n10455) );
  XOR U12361 ( .A(n10460), .B(n10281), .Z(n10283) );
  XOR U12362 ( .A(n10461), .B(n10462), .Z(n10281) );
  AND U12363 ( .A(n10463), .B(n10464), .Z(n10461) );
  AND U12364 ( .A(a[56]), .B(b[15]), .Z(n10460) );
  XOR U12365 ( .A(n10465), .B(n10286), .Z(n10288) );
  XOR U12366 ( .A(n10466), .B(n10467), .Z(n10286) );
  AND U12367 ( .A(n10468), .B(n10469), .Z(n10466) );
  AND U12368 ( .A(a[57]), .B(b[14]), .Z(n10465) );
  XOR U12369 ( .A(n10470), .B(n10291), .Z(n10293) );
  XOR U12370 ( .A(n10471), .B(n10472), .Z(n10291) );
  AND U12371 ( .A(n10473), .B(n10474), .Z(n10471) );
  AND U12372 ( .A(a[58]), .B(b[13]), .Z(n10470) );
  XOR U12373 ( .A(n10475), .B(n10296), .Z(n10298) );
  XOR U12374 ( .A(n10476), .B(n10477), .Z(n10296) );
  AND U12375 ( .A(n10478), .B(n10479), .Z(n10476) );
  AND U12376 ( .A(a[59]), .B(b[12]), .Z(n10475) );
  XOR U12377 ( .A(n10480), .B(n10301), .Z(n10303) );
  XOR U12378 ( .A(n10481), .B(n10482), .Z(n10301) );
  AND U12379 ( .A(n10483), .B(n10484), .Z(n10481) );
  AND U12380 ( .A(a[60]), .B(b[11]), .Z(n10480) );
  XOR U12381 ( .A(n10485), .B(n10306), .Z(n10308) );
  XOR U12382 ( .A(n10486), .B(n10487), .Z(n10306) );
  AND U12383 ( .A(n10488), .B(n10489), .Z(n10486) );
  AND U12384 ( .A(a[61]), .B(b[10]), .Z(n10485) );
  XOR U12385 ( .A(n10490), .B(n10311), .Z(n10313) );
  XOR U12386 ( .A(n10491), .B(n10492), .Z(n10311) );
  AND U12387 ( .A(n10493), .B(n10494), .Z(n10491) );
  AND U12388 ( .A(a[62]), .B(b[9]), .Z(n10490) );
  XOR U12389 ( .A(n10495), .B(n10316), .Z(n10318) );
  XOR U12390 ( .A(n10496), .B(n10497), .Z(n10316) );
  AND U12391 ( .A(n10498), .B(n10499), .Z(n10496) );
  AND U12392 ( .A(a[63]), .B(b[8]), .Z(n10495) );
  XOR U12393 ( .A(n10500), .B(n10321), .Z(n10323) );
  XOR U12394 ( .A(n10501), .B(n10502), .Z(n10321) );
  AND U12395 ( .A(n10503), .B(n10504), .Z(n10501) );
  AND U12396 ( .A(a[64]), .B(b[7]), .Z(n10500) );
  XOR U12397 ( .A(n10505), .B(n10326), .Z(n10328) );
  XOR U12398 ( .A(n10506), .B(n10507), .Z(n10326) );
  AND U12399 ( .A(n10508), .B(n10509), .Z(n10506) );
  AND U12400 ( .A(a[65]), .B(b[6]), .Z(n10505) );
  XOR U12401 ( .A(n10510), .B(n10331), .Z(n10333) );
  XOR U12402 ( .A(n10511), .B(n10512), .Z(n10331) );
  AND U12403 ( .A(n10513), .B(n10514), .Z(n10511) );
  AND U12404 ( .A(a[66]), .B(b[5]), .Z(n10510) );
  XNOR U12405 ( .A(n10515), .B(n10516), .Z(n10335) );
  ANDN U12406 ( .B(n10517), .A(n10518), .Z(n10515) );
  XOR U12407 ( .A(n10519), .B(n10340), .Z(n10342) );
  XOR U12408 ( .A(n10520), .B(n10521), .Z(n10340) );
  AND U12409 ( .A(n10522), .B(n10523), .Z(n10520) );
  AND U12410 ( .A(a[67]), .B(b[4]), .Z(n10519) );
  XOR U12411 ( .A(n10525), .B(n10526), .Z(n10345) );
  OR U12412 ( .A(n10527), .B(n10528), .Z(n10526) );
  AND U12413 ( .A(a[69]), .B(b[2]), .Z(n10524) );
  XNOR U12414 ( .A(n10355), .B(n10529), .Z(n10351) );
  NAND U12415 ( .A(a[70]), .B(b[1]), .Z(n10529) );
  IV U12416 ( .A(n10349), .Z(n10355) );
  ANDN U12417 ( .B(n5202), .A(n5204), .Z(n10349) );
  NAND U12418 ( .A(a[70]), .B(b[0]), .Z(n5204) );
  XOR U12419 ( .A(n10527), .B(n10528), .Z(n5202) );
  XNOR U12420 ( .A(n10531), .B(n10518), .Z(n10530) );
  XOR U12421 ( .A(n10532), .B(n10516), .Z(n10518) );
  AND U12422 ( .A(b[2]), .B(a[68]), .Z(n10532) );
  XOR U12423 ( .A(n10516), .B(n10522), .Z(n10533) );
  XNOR U12424 ( .A(n10521), .B(n10513), .Z(n10534) );
  XNOR U12425 ( .A(n10512), .B(n10508), .Z(n10535) );
  XNOR U12426 ( .A(n10507), .B(n10503), .Z(n10536) );
  XNOR U12427 ( .A(n10502), .B(n10498), .Z(n10537) );
  XNOR U12428 ( .A(n10497), .B(n10493), .Z(n10538) );
  XNOR U12429 ( .A(n10492), .B(n10488), .Z(n10539) );
  XNOR U12430 ( .A(n10487), .B(n10483), .Z(n10540) );
  XNOR U12431 ( .A(n10482), .B(n10478), .Z(n10541) );
  XNOR U12432 ( .A(n10477), .B(n10473), .Z(n10542) );
  XNOR U12433 ( .A(n10472), .B(n10468), .Z(n10543) );
  XNOR U12434 ( .A(n10467), .B(n10463), .Z(n10544) );
  XNOR U12435 ( .A(n10462), .B(n10458), .Z(n10545) );
  XNOR U12436 ( .A(n10457), .B(n10453), .Z(n10546) );
  XNOR U12437 ( .A(n10452), .B(n10448), .Z(n10547) );
  XNOR U12438 ( .A(n10447), .B(n10443), .Z(n10548) );
  XNOR U12439 ( .A(n10442), .B(n10438), .Z(n10549) );
  XNOR U12440 ( .A(n10437), .B(n10433), .Z(n10550) );
  XNOR U12441 ( .A(n10432), .B(n10428), .Z(n10551) );
  XNOR U12442 ( .A(n10427), .B(n10423), .Z(n10552) );
  XNOR U12443 ( .A(n10422), .B(n10418), .Z(n10553) );
  XNOR U12444 ( .A(n10417), .B(n10413), .Z(n10554) );
  XNOR U12445 ( .A(n10412), .B(n10408), .Z(n10555) );
  XNOR U12446 ( .A(n10407), .B(n10403), .Z(n10556) );
  XNOR U12447 ( .A(n10402), .B(n10398), .Z(n10557) );
  XOR U12448 ( .A(n10397), .B(n10394), .Z(n10558) );
  XOR U12449 ( .A(n10559), .B(n10560), .Z(n10394) );
  XOR U12450 ( .A(n10392), .B(n10561), .Z(n10560) );
  XOR U12451 ( .A(n10562), .B(n10563), .Z(n10561) );
  XOR U12452 ( .A(n10564), .B(n10565), .Z(n10563) );
  NAND U12453 ( .A(a[40]), .B(b[30]), .Z(n10565) );
  AND U12454 ( .A(a[39]), .B(b[31]), .Z(n10564) );
  XOR U12455 ( .A(n10566), .B(n10562), .Z(n10559) );
  XOR U12456 ( .A(n10567), .B(n10568), .Z(n10562) );
  ANDN U12457 ( .B(n10569), .A(n10570), .Z(n10567) );
  AND U12458 ( .A(a[41]), .B(b[29]), .Z(n10566) );
  XOR U12459 ( .A(n10571), .B(n10392), .Z(n10393) );
  XOR U12460 ( .A(n10572), .B(n10573), .Z(n10392) );
  AND U12461 ( .A(n10574), .B(n10575), .Z(n10572) );
  AND U12462 ( .A(a[42]), .B(b[28]), .Z(n10571) );
  XOR U12463 ( .A(n10576), .B(n10397), .Z(n10399) );
  XOR U12464 ( .A(n10577), .B(n10578), .Z(n10397) );
  AND U12465 ( .A(n10579), .B(n10580), .Z(n10577) );
  AND U12466 ( .A(a[43]), .B(b[27]), .Z(n10576) );
  XOR U12467 ( .A(n10581), .B(n10402), .Z(n10404) );
  XOR U12468 ( .A(n10582), .B(n10583), .Z(n10402) );
  AND U12469 ( .A(n10584), .B(n10585), .Z(n10582) );
  AND U12470 ( .A(a[44]), .B(b[26]), .Z(n10581) );
  XOR U12471 ( .A(n10586), .B(n10407), .Z(n10409) );
  XOR U12472 ( .A(n10587), .B(n10588), .Z(n10407) );
  AND U12473 ( .A(n10589), .B(n10590), .Z(n10587) );
  AND U12474 ( .A(a[45]), .B(b[25]), .Z(n10586) );
  XOR U12475 ( .A(n10591), .B(n10412), .Z(n10414) );
  XOR U12476 ( .A(n10592), .B(n10593), .Z(n10412) );
  AND U12477 ( .A(n10594), .B(n10595), .Z(n10592) );
  AND U12478 ( .A(a[46]), .B(b[24]), .Z(n10591) );
  XOR U12479 ( .A(n10596), .B(n10417), .Z(n10419) );
  XOR U12480 ( .A(n10597), .B(n10598), .Z(n10417) );
  AND U12481 ( .A(n10599), .B(n10600), .Z(n10597) );
  AND U12482 ( .A(a[47]), .B(b[23]), .Z(n10596) );
  XOR U12483 ( .A(n10601), .B(n10422), .Z(n10424) );
  XOR U12484 ( .A(n10602), .B(n10603), .Z(n10422) );
  AND U12485 ( .A(n10604), .B(n10605), .Z(n10602) );
  AND U12486 ( .A(a[48]), .B(b[22]), .Z(n10601) );
  XOR U12487 ( .A(n10606), .B(n10427), .Z(n10429) );
  XOR U12488 ( .A(n10607), .B(n10608), .Z(n10427) );
  AND U12489 ( .A(n10609), .B(n10610), .Z(n10607) );
  AND U12490 ( .A(a[49]), .B(b[21]), .Z(n10606) );
  XOR U12491 ( .A(n10611), .B(n10432), .Z(n10434) );
  XOR U12492 ( .A(n10612), .B(n10613), .Z(n10432) );
  AND U12493 ( .A(n10614), .B(n10615), .Z(n10612) );
  AND U12494 ( .A(a[50]), .B(b[20]), .Z(n10611) );
  XOR U12495 ( .A(n10616), .B(n10437), .Z(n10439) );
  XOR U12496 ( .A(n10617), .B(n10618), .Z(n10437) );
  AND U12497 ( .A(n10619), .B(n10620), .Z(n10617) );
  AND U12498 ( .A(a[51]), .B(b[19]), .Z(n10616) );
  XOR U12499 ( .A(n10621), .B(n10442), .Z(n10444) );
  XOR U12500 ( .A(n10622), .B(n10623), .Z(n10442) );
  AND U12501 ( .A(n10624), .B(n10625), .Z(n10622) );
  AND U12502 ( .A(a[52]), .B(b[18]), .Z(n10621) );
  XOR U12503 ( .A(n10626), .B(n10447), .Z(n10449) );
  XOR U12504 ( .A(n10627), .B(n10628), .Z(n10447) );
  AND U12505 ( .A(n10629), .B(n10630), .Z(n10627) );
  AND U12506 ( .A(a[53]), .B(b[17]), .Z(n10626) );
  XOR U12507 ( .A(n10631), .B(n10452), .Z(n10454) );
  XOR U12508 ( .A(n10632), .B(n10633), .Z(n10452) );
  AND U12509 ( .A(n10634), .B(n10635), .Z(n10632) );
  AND U12510 ( .A(a[54]), .B(b[16]), .Z(n10631) );
  XOR U12511 ( .A(n10636), .B(n10457), .Z(n10459) );
  XOR U12512 ( .A(n10637), .B(n10638), .Z(n10457) );
  AND U12513 ( .A(n10639), .B(n10640), .Z(n10637) );
  AND U12514 ( .A(a[55]), .B(b[15]), .Z(n10636) );
  XOR U12515 ( .A(n10641), .B(n10462), .Z(n10464) );
  XOR U12516 ( .A(n10642), .B(n10643), .Z(n10462) );
  AND U12517 ( .A(n10644), .B(n10645), .Z(n10642) );
  AND U12518 ( .A(a[56]), .B(b[14]), .Z(n10641) );
  XOR U12519 ( .A(n10646), .B(n10467), .Z(n10469) );
  XOR U12520 ( .A(n10647), .B(n10648), .Z(n10467) );
  AND U12521 ( .A(n10649), .B(n10650), .Z(n10647) );
  AND U12522 ( .A(a[57]), .B(b[13]), .Z(n10646) );
  XOR U12523 ( .A(n10651), .B(n10472), .Z(n10474) );
  XOR U12524 ( .A(n10652), .B(n10653), .Z(n10472) );
  AND U12525 ( .A(n10654), .B(n10655), .Z(n10652) );
  AND U12526 ( .A(a[58]), .B(b[12]), .Z(n10651) );
  XOR U12527 ( .A(n10656), .B(n10477), .Z(n10479) );
  XOR U12528 ( .A(n10657), .B(n10658), .Z(n10477) );
  AND U12529 ( .A(n10659), .B(n10660), .Z(n10657) );
  AND U12530 ( .A(a[59]), .B(b[11]), .Z(n10656) );
  XOR U12531 ( .A(n10661), .B(n10482), .Z(n10484) );
  XOR U12532 ( .A(n10662), .B(n10663), .Z(n10482) );
  AND U12533 ( .A(n10664), .B(n10665), .Z(n10662) );
  AND U12534 ( .A(a[60]), .B(b[10]), .Z(n10661) );
  XOR U12535 ( .A(n10666), .B(n10487), .Z(n10489) );
  XOR U12536 ( .A(n10667), .B(n10668), .Z(n10487) );
  AND U12537 ( .A(n10669), .B(n10670), .Z(n10667) );
  AND U12538 ( .A(a[61]), .B(b[9]), .Z(n10666) );
  XOR U12539 ( .A(n10671), .B(n10492), .Z(n10494) );
  XOR U12540 ( .A(n10672), .B(n10673), .Z(n10492) );
  AND U12541 ( .A(n10674), .B(n10675), .Z(n10672) );
  AND U12542 ( .A(a[62]), .B(b[8]), .Z(n10671) );
  XOR U12543 ( .A(n10676), .B(n10497), .Z(n10499) );
  XOR U12544 ( .A(n10677), .B(n10678), .Z(n10497) );
  AND U12545 ( .A(n10679), .B(n10680), .Z(n10677) );
  AND U12546 ( .A(a[63]), .B(b[7]), .Z(n10676) );
  XOR U12547 ( .A(n10681), .B(n10502), .Z(n10504) );
  XOR U12548 ( .A(n10682), .B(n10683), .Z(n10502) );
  AND U12549 ( .A(n10684), .B(n10685), .Z(n10682) );
  AND U12550 ( .A(a[64]), .B(b[6]), .Z(n10681) );
  XOR U12551 ( .A(n10686), .B(n10507), .Z(n10509) );
  XOR U12552 ( .A(n10687), .B(n10688), .Z(n10507) );
  AND U12553 ( .A(n10689), .B(n10690), .Z(n10687) );
  AND U12554 ( .A(a[65]), .B(b[5]), .Z(n10686) );
  XOR U12555 ( .A(n10691), .B(n10512), .Z(n10514) );
  XOR U12556 ( .A(n10692), .B(n10693), .Z(n10512) );
  AND U12557 ( .A(n10694), .B(n10695), .Z(n10692) );
  AND U12558 ( .A(a[66]), .B(b[4]), .Z(n10691) );
  XOR U12559 ( .A(n10696), .B(n10697), .Z(n10516) );
  OR U12560 ( .A(n10698), .B(n10699), .Z(n10697) );
  XOR U12561 ( .A(n10700), .B(n10521), .Z(n10523) );
  XNOR U12562 ( .A(n10701), .B(n10702), .Z(n10521) );
  ANDN U12563 ( .B(n10703), .A(n10704), .Z(n10701) );
  AND U12564 ( .A(a[67]), .B(b[3]), .Z(n10700) );
  XNOR U12565 ( .A(n10531), .B(n10705), .Z(n10527) );
  NAND U12566 ( .A(a[69]), .B(b[1]), .Z(n10705) );
  IV U12567 ( .A(n10525), .Z(n10531) );
  ANDN U12568 ( .B(n5207), .A(n5209), .Z(n10525) );
  NAND U12569 ( .A(a[69]), .B(b[0]), .Z(n5209) );
  XOR U12570 ( .A(n10699), .B(n10698), .Z(n5207) );
  XOR U12571 ( .A(n10696), .B(n10706), .Z(n10698) );
  NAND U12572 ( .A(b[1]), .B(a[68]), .Z(n10706) );
  XOR U12573 ( .A(n10696), .B(n10704), .Z(n10707) );
  XOR U12574 ( .A(n10708), .B(n10702), .Z(n10704) );
  AND U12575 ( .A(a[67]), .B(b[2]), .Z(n10708) );
  ANDN U12576 ( .B(n5212), .A(n5214), .Z(n10696) );
  NAND U12577 ( .A(a[68]), .B(b[0]), .Z(n5214) );
  XOR U12578 ( .A(n10709), .B(n10710), .Z(n5212) );
  XOR U12579 ( .A(n10702), .B(n10694), .Z(n10711) );
  XNOR U12580 ( .A(n10693), .B(n10689), .Z(n10712) );
  XNOR U12581 ( .A(n10688), .B(n10684), .Z(n10713) );
  XNOR U12582 ( .A(n10683), .B(n10679), .Z(n10714) );
  XNOR U12583 ( .A(n10678), .B(n10674), .Z(n10715) );
  XNOR U12584 ( .A(n10673), .B(n10669), .Z(n10716) );
  XNOR U12585 ( .A(n10668), .B(n10664), .Z(n10717) );
  XNOR U12586 ( .A(n10663), .B(n10659), .Z(n10718) );
  XNOR U12587 ( .A(n10658), .B(n10654), .Z(n10719) );
  XNOR U12588 ( .A(n10653), .B(n10649), .Z(n10720) );
  XNOR U12589 ( .A(n10648), .B(n10644), .Z(n10721) );
  XNOR U12590 ( .A(n10643), .B(n10639), .Z(n10722) );
  XNOR U12591 ( .A(n10638), .B(n10634), .Z(n10723) );
  XNOR U12592 ( .A(n10633), .B(n10629), .Z(n10724) );
  XNOR U12593 ( .A(n10628), .B(n10624), .Z(n10725) );
  XNOR U12594 ( .A(n10623), .B(n10619), .Z(n10726) );
  XNOR U12595 ( .A(n10618), .B(n10614), .Z(n10727) );
  XNOR U12596 ( .A(n10613), .B(n10609), .Z(n10728) );
  XNOR U12597 ( .A(n10608), .B(n10604), .Z(n10729) );
  XNOR U12598 ( .A(n10603), .B(n10599), .Z(n10730) );
  XNOR U12599 ( .A(n10598), .B(n10594), .Z(n10731) );
  XNOR U12600 ( .A(n10593), .B(n10589), .Z(n10732) );
  XNOR U12601 ( .A(n10588), .B(n10584), .Z(n10733) );
  XNOR U12602 ( .A(n10583), .B(n10579), .Z(n10734) );
  XNOR U12603 ( .A(n10578), .B(n10574), .Z(n10735) );
  XOR U12604 ( .A(n10573), .B(n10570), .Z(n10736) );
  XOR U12605 ( .A(n10737), .B(n10738), .Z(n10570) );
  XOR U12606 ( .A(n10568), .B(n10739), .Z(n10738) );
  XNOR U12607 ( .A(n10740), .B(n10741), .Z(n10739) );
  XOR U12608 ( .A(n10742), .B(n10743), .Z(n10741) );
  NAND U12609 ( .A(a[39]), .B(b[30]), .Z(n10743) );
  AND U12610 ( .A(a[38]), .B(b[31]), .Z(n10742) );
  XNOR U12611 ( .A(n10744), .B(n10740), .Z(n10737) );
  XNOR U12612 ( .A(n10745), .B(n10746), .Z(n10740) );
  ANDN U12613 ( .B(n10747), .A(n10748), .Z(n10745) );
  AND U12614 ( .A(a[40]), .B(b[29]), .Z(n10744) );
  XOR U12615 ( .A(n10749), .B(n10568), .Z(n10569) );
  XOR U12616 ( .A(n10750), .B(n10751), .Z(n10568) );
  AND U12617 ( .A(n10752), .B(n10753), .Z(n10750) );
  AND U12618 ( .A(a[41]), .B(b[28]), .Z(n10749) );
  XOR U12619 ( .A(n10754), .B(n10573), .Z(n10575) );
  XOR U12620 ( .A(n10755), .B(n10756), .Z(n10573) );
  AND U12621 ( .A(n10757), .B(n10758), .Z(n10755) );
  AND U12622 ( .A(a[42]), .B(b[27]), .Z(n10754) );
  XOR U12623 ( .A(n10759), .B(n10578), .Z(n10580) );
  XOR U12624 ( .A(n10760), .B(n10761), .Z(n10578) );
  AND U12625 ( .A(n10762), .B(n10763), .Z(n10760) );
  AND U12626 ( .A(a[43]), .B(b[26]), .Z(n10759) );
  XOR U12627 ( .A(n10764), .B(n10583), .Z(n10585) );
  XOR U12628 ( .A(n10765), .B(n10766), .Z(n10583) );
  AND U12629 ( .A(n10767), .B(n10768), .Z(n10765) );
  AND U12630 ( .A(a[44]), .B(b[25]), .Z(n10764) );
  XOR U12631 ( .A(n10769), .B(n10588), .Z(n10590) );
  XOR U12632 ( .A(n10770), .B(n10771), .Z(n10588) );
  AND U12633 ( .A(n10772), .B(n10773), .Z(n10770) );
  AND U12634 ( .A(a[45]), .B(b[24]), .Z(n10769) );
  XOR U12635 ( .A(n10774), .B(n10593), .Z(n10595) );
  XOR U12636 ( .A(n10775), .B(n10776), .Z(n10593) );
  AND U12637 ( .A(n10777), .B(n10778), .Z(n10775) );
  AND U12638 ( .A(a[46]), .B(b[23]), .Z(n10774) );
  XOR U12639 ( .A(n10779), .B(n10598), .Z(n10600) );
  XOR U12640 ( .A(n10780), .B(n10781), .Z(n10598) );
  AND U12641 ( .A(n10782), .B(n10783), .Z(n10780) );
  AND U12642 ( .A(a[47]), .B(b[22]), .Z(n10779) );
  XOR U12643 ( .A(n10784), .B(n10603), .Z(n10605) );
  XOR U12644 ( .A(n10785), .B(n10786), .Z(n10603) );
  AND U12645 ( .A(n10787), .B(n10788), .Z(n10785) );
  AND U12646 ( .A(a[48]), .B(b[21]), .Z(n10784) );
  XOR U12647 ( .A(n10789), .B(n10608), .Z(n10610) );
  XOR U12648 ( .A(n10790), .B(n10791), .Z(n10608) );
  AND U12649 ( .A(n10792), .B(n10793), .Z(n10790) );
  AND U12650 ( .A(a[49]), .B(b[20]), .Z(n10789) );
  XOR U12651 ( .A(n10794), .B(n10613), .Z(n10615) );
  XOR U12652 ( .A(n10795), .B(n10796), .Z(n10613) );
  AND U12653 ( .A(n10797), .B(n10798), .Z(n10795) );
  AND U12654 ( .A(a[50]), .B(b[19]), .Z(n10794) );
  XOR U12655 ( .A(n10799), .B(n10618), .Z(n10620) );
  XOR U12656 ( .A(n10800), .B(n10801), .Z(n10618) );
  AND U12657 ( .A(n10802), .B(n10803), .Z(n10800) );
  AND U12658 ( .A(a[51]), .B(b[18]), .Z(n10799) );
  XOR U12659 ( .A(n10804), .B(n10623), .Z(n10625) );
  XOR U12660 ( .A(n10805), .B(n10806), .Z(n10623) );
  AND U12661 ( .A(n10807), .B(n10808), .Z(n10805) );
  AND U12662 ( .A(a[52]), .B(b[17]), .Z(n10804) );
  XOR U12663 ( .A(n10809), .B(n10628), .Z(n10630) );
  XOR U12664 ( .A(n10810), .B(n10811), .Z(n10628) );
  AND U12665 ( .A(n10812), .B(n10813), .Z(n10810) );
  AND U12666 ( .A(a[53]), .B(b[16]), .Z(n10809) );
  XOR U12667 ( .A(n10814), .B(n10633), .Z(n10635) );
  XOR U12668 ( .A(n10815), .B(n10816), .Z(n10633) );
  AND U12669 ( .A(n10817), .B(n10818), .Z(n10815) );
  AND U12670 ( .A(a[54]), .B(b[15]), .Z(n10814) );
  XOR U12671 ( .A(n10819), .B(n10638), .Z(n10640) );
  XOR U12672 ( .A(n10820), .B(n10821), .Z(n10638) );
  AND U12673 ( .A(n10822), .B(n10823), .Z(n10820) );
  AND U12674 ( .A(a[55]), .B(b[14]), .Z(n10819) );
  XOR U12675 ( .A(n10824), .B(n10643), .Z(n10645) );
  XOR U12676 ( .A(n10825), .B(n10826), .Z(n10643) );
  AND U12677 ( .A(n10827), .B(n10828), .Z(n10825) );
  AND U12678 ( .A(a[56]), .B(b[13]), .Z(n10824) );
  XOR U12679 ( .A(n10829), .B(n10648), .Z(n10650) );
  XOR U12680 ( .A(n10830), .B(n10831), .Z(n10648) );
  AND U12681 ( .A(n10832), .B(n10833), .Z(n10830) );
  AND U12682 ( .A(a[57]), .B(b[12]), .Z(n10829) );
  XOR U12683 ( .A(n10834), .B(n10653), .Z(n10655) );
  XOR U12684 ( .A(n10835), .B(n10836), .Z(n10653) );
  AND U12685 ( .A(n10837), .B(n10838), .Z(n10835) );
  AND U12686 ( .A(a[58]), .B(b[11]), .Z(n10834) );
  XOR U12687 ( .A(n10839), .B(n10658), .Z(n10660) );
  XOR U12688 ( .A(n10840), .B(n10841), .Z(n10658) );
  AND U12689 ( .A(n10842), .B(n10843), .Z(n10840) );
  AND U12690 ( .A(a[59]), .B(b[10]), .Z(n10839) );
  XOR U12691 ( .A(n10844), .B(n10663), .Z(n10665) );
  XOR U12692 ( .A(n10845), .B(n10846), .Z(n10663) );
  AND U12693 ( .A(n10847), .B(n10848), .Z(n10845) );
  AND U12694 ( .A(a[60]), .B(b[9]), .Z(n10844) );
  XOR U12695 ( .A(n10849), .B(n10668), .Z(n10670) );
  XOR U12696 ( .A(n10850), .B(n10851), .Z(n10668) );
  AND U12697 ( .A(n10852), .B(n10853), .Z(n10850) );
  AND U12698 ( .A(a[61]), .B(b[8]), .Z(n10849) );
  XOR U12699 ( .A(n10854), .B(n10673), .Z(n10675) );
  XOR U12700 ( .A(n10855), .B(n10856), .Z(n10673) );
  AND U12701 ( .A(n10857), .B(n10858), .Z(n10855) );
  AND U12702 ( .A(a[62]), .B(b[7]), .Z(n10854) );
  XOR U12703 ( .A(n10859), .B(n10678), .Z(n10680) );
  XOR U12704 ( .A(n10860), .B(n10861), .Z(n10678) );
  AND U12705 ( .A(n10862), .B(n10863), .Z(n10860) );
  AND U12706 ( .A(a[63]), .B(b[6]), .Z(n10859) );
  XOR U12707 ( .A(n10864), .B(n10683), .Z(n10685) );
  XOR U12708 ( .A(n10865), .B(n10866), .Z(n10683) );
  AND U12709 ( .A(n10867), .B(n10868), .Z(n10865) );
  AND U12710 ( .A(a[64]), .B(b[5]), .Z(n10864) );
  XOR U12711 ( .A(n10869), .B(n10688), .Z(n10690) );
  XOR U12712 ( .A(n10870), .B(n10871), .Z(n10688) );
  AND U12713 ( .A(n10872), .B(n10873), .Z(n10870) );
  AND U12714 ( .A(a[65]), .B(b[4]), .Z(n10869) );
  XNOR U12715 ( .A(n10874), .B(n10875), .Z(n10702) );
  OR U12716 ( .A(n10710), .B(n10709), .Z(n10875) );
  XNOR U12717 ( .A(n10874), .B(n10876), .Z(n10709) );
  NAND U12718 ( .A(a[67]), .B(b[1]), .Z(n10876) );
  XOR U12719 ( .A(n10877), .B(n10878), .Z(n10710) );
  XOR U12720 ( .A(n10874), .B(n10879), .Z(n10878) );
  NANDN U12721 ( .A(n5219), .B(n5217), .Z(n10874) );
  XNOR U12722 ( .A(n10880), .B(n10881), .Z(n5217) );
  NAND U12723 ( .A(a[67]), .B(b[0]), .Z(n5219) );
  XOR U12724 ( .A(n10882), .B(n10693), .Z(n10695) );
  XNOR U12725 ( .A(n10883), .B(n10884), .Z(n10693) );
  AND U12726 ( .A(n10879), .B(n10877), .Z(n10883) );
  XNOR U12727 ( .A(n10885), .B(n10884), .Z(n10877) );
  AND U12728 ( .A(b[2]), .B(a[66]), .Z(n10885) );
  XOR U12729 ( .A(n10872), .B(n10884), .Z(n10886) );
  XOR U12730 ( .A(n10887), .B(n10888), .Z(n10884) );
  NANDN U12731 ( .A(n10880), .B(n10881), .Z(n10888) );
  XNOR U12732 ( .A(n10889), .B(n10890), .Z(n10881) );
  XNOR U12733 ( .A(n10887), .B(n10891), .Z(n10890) );
  NAND U12734 ( .A(a[66]), .B(b[1]), .Z(n10892) );
  ANDN U12735 ( .B(n5222), .A(n5224), .Z(n10887) );
  NAND U12736 ( .A(a[66]), .B(b[0]), .Z(n5224) );
  XNOR U12737 ( .A(n10893), .B(n10894), .Z(n5222) );
  XOR U12738 ( .A(n10867), .B(n10896), .Z(n10895) );
  XOR U12739 ( .A(n10862), .B(n10898), .Z(n10897) );
  XOR U12740 ( .A(n10857), .B(n10900), .Z(n10899) );
  XOR U12741 ( .A(n10852), .B(n10902), .Z(n10901) );
  XOR U12742 ( .A(n10847), .B(n10904), .Z(n10903) );
  XOR U12743 ( .A(n10842), .B(n10906), .Z(n10905) );
  XOR U12744 ( .A(n10837), .B(n10908), .Z(n10907) );
  XOR U12745 ( .A(n10832), .B(n10910), .Z(n10909) );
  XOR U12746 ( .A(n10827), .B(n10912), .Z(n10911) );
  XOR U12747 ( .A(n10822), .B(n10914), .Z(n10913) );
  XOR U12748 ( .A(n10817), .B(n10916), .Z(n10915) );
  XOR U12749 ( .A(n10812), .B(n10918), .Z(n10917) );
  XOR U12750 ( .A(n10807), .B(n10920), .Z(n10919) );
  XOR U12751 ( .A(n10802), .B(n10922), .Z(n10921) );
  XOR U12752 ( .A(n10797), .B(n10924), .Z(n10923) );
  XOR U12753 ( .A(n10792), .B(n10926), .Z(n10925) );
  XOR U12754 ( .A(n10787), .B(n10928), .Z(n10927) );
  XOR U12755 ( .A(n10782), .B(n10930), .Z(n10929) );
  XOR U12756 ( .A(n10777), .B(n10932), .Z(n10931) );
  XOR U12757 ( .A(n10772), .B(n10934), .Z(n10933) );
  XOR U12758 ( .A(n10767), .B(n10936), .Z(n10935) );
  XOR U12759 ( .A(n10762), .B(n10938), .Z(n10937) );
  XOR U12760 ( .A(n10757), .B(n10940), .Z(n10939) );
  XOR U12761 ( .A(n10752), .B(n10942), .Z(n10941) );
  XNOR U12762 ( .A(n10748), .B(n10944), .Z(n10943) );
  XOR U12763 ( .A(n10945), .B(n10946), .Z(n10748) );
  XOR U12764 ( .A(n10947), .B(n10948), .Z(n10946) );
  XNOR U12765 ( .A(n10949), .B(n10950), .Z(n10947) );
  XOR U12766 ( .A(n10951), .B(n10952), .Z(n10950) );
  AND U12767 ( .A(b[31]), .B(a[37]), .Z(n10952) );
  AND U12768 ( .A(a[38]), .B(b[30]), .Z(n10951) );
  XNOR U12769 ( .A(n10953), .B(n10949), .Z(n10945) );
  XNOR U12770 ( .A(n10954), .B(n10955), .Z(n10949) );
  ANDN U12771 ( .B(n10956), .A(n10957), .Z(n10954) );
  AND U12772 ( .A(a[39]), .B(b[29]), .Z(n10953) );
  XOR U12773 ( .A(n10958), .B(n10746), .Z(n10747) );
  IV U12774 ( .A(n10948), .Z(n10746) );
  XOR U12775 ( .A(n10959), .B(n10960), .Z(n10948) );
  AND U12776 ( .A(n10961), .B(n10962), .Z(n10959) );
  AND U12777 ( .A(a[40]), .B(b[28]), .Z(n10958) );
  XOR U12778 ( .A(n10963), .B(n10751), .Z(n10753) );
  IV U12779 ( .A(n10944), .Z(n10751) );
  XOR U12780 ( .A(n10964), .B(n10965), .Z(n10944) );
  AND U12781 ( .A(n10966), .B(n10967), .Z(n10964) );
  AND U12782 ( .A(a[41]), .B(b[27]), .Z(n10963) );
  XOR U12783 ( .A(n10968), .B(n10756), .Z(n10758) );
  IV U12784 ( .A(n10942), .Z(n10756) );
  XOR U12785 ( .A(n10969), .B(n10970), .Z(n10942) );
  AND U12786 ( .A(n10971), .B(n10972), .Z(n10969) );
  AND U12787 ( .A(a[42]), .B(b[26]), .Z(n10968) );
  XOR U12788 ( .A(n10973), .B(n10761), .Z(n10763) );
  IV U12789 ( .A(n10940), .Z(n10761) );
  XOR U12790 ( .A(n10974), .B(n10975), .Z(n10940) );
  AND U12791 ( .A(n10976), .B(n10977), .Z(n10974) );
  AND U12792 ( .A(a[43]), .B(b[25]), .Z(n10973) );
  XOR U12793 ( .A(n10978), .B(n10766), .Z(n10768) );
  IV U12794 ( .A(n10938), .Z(n10766) );
  XOR U12795 ( .A(n10979), .B(n10980), .Z(n10938) );
  AND U12796 ( .A(n10981), .B(n10982), .Z(n10979) );
  AND U12797 ( .A(a[44]), .B(b[24]), .Z(n10978) );
  XOR U12798 ( .A(n10983), .B(n10771), .Z(n10773) );
  IV U12799 ( .A(n10936), .Z(n10771) );
  XOR U12800 ( .A(n10984), .B(n10985), .Z(n10936) );
  AND U12801 ( .A(n10986), .B(n10987), .Z(n10984) );
  AND U12802 ( .A(a[45]), .B(b[23]), .Z(n10983) );
  XOR U12803 ( .A(n10988), .B(n10776), .Z(n10778) );
  IV U12804 ( .A(n10934), .Z(n10776) );
  XOR U12805 ( .A(n10989), .B(n10990), .Z(n10934) );
  AND U12806 ( .A(n10991), .B(n10992), .Z(n10989) );
  AND U12807 ( .A(a[46]), .B(b[22]), .Z(n10988) );
  XOR U12808 ( .A(n10993), .B(n10781), .Z(n10783) );
  IV U12809 ( .A(n10932), .Z(n10781) );
  XOR U12810 ( .A(n10994), .B(n10995), .Z(n10932) );
  AND U12811 ( .A(n10996), .B(n10997), .Z(n10994) );
  AND U12812 ( .A(a[47]), .B(b[21]), .Z(n10993) );
  XOR U12813 ( .A(n10998), .B(n10786), .Z(n10788) );
  IV U12814 ( .A(n10930), .Z(n10786) );
  XOR U12815 ( .A(n10999), .B(n11000), .Z(n10930) );
  AND U12816 ( .A(n11001), .B(n11002), .Z(n10999) );
  AND U12817 ( .A(a[48]), .B(b[20]), .Z(n10998) );
  XOR U12818 ( .A(n11003), .B(n10791), .Z(n10793) );
  IV U12819 ( .A(n10928), .Z(n10791) );
  XOR U12820 ( .A(n11004), .B(n11005), .Z(n10928) );
  AND U12821 ( .A(n11006), .B(n11007), .Z(n11004) );
  AND U12822 ( .A(a[49]), .B(b[19]), .Z(n11003) );
  XOR U12823 ( .A(n11008), .B(n10796), .Z(n10798) );
  IV U12824 ( .A(n10926), .Z(n10796) );
  XOR U12825 ( .A(n11009), .B(n11010), .Z(n10926) );
  AND U12826 ( .A(n11011), .B(n11012), .Z(n11009) );
  AND U12827 ( .A(a[50]), .B(b[18]), .Z(n11008) );
  XOR U12828 ( .A(n11013), .B(n10801), .Z(n10803) );
  IV U12829 ( .A(n10924), .Z(n10801) );
  XOR U12830 ( .A(n11014), .B(n11015), .Z(n10924) );
  AND U12831 ( .A(n11016), .B(n11017), .Z(n11014) );
  AND U12832 ( .A(a[51]), .B(b[17]), .Z(n11013) );
  XOR U12833 ( .A(n11018), .B(n10806), .Z(n10808) );
  IV U12834 ( .A(n10922), .Z(n10806) );
  XOR U12835 ( .A(n11019), .B(n11020), .Z(n10922) );
  AND U12836 ( .A(n11021), .B(n11022), .Z(n11019) );
  AND U12837 ( .A(a[52]), .B(b[16]), .Z(n11018) );
  XOR U12838 ( .A(n11023), .B(n10811), .Z(n10813) );
  IV U12839 ( .A(n10920), .Z(n10811) );
  XOR U12840 ( .A(n11024), .B(n11025), .Z(n10920) );
  AND U12841 ( .A(n11026), .B(n11027), .Z(n11024) );
  AND U12842 ( .A(a[53]), .B(b[15]), .Z(n11023) );
  XOR U12843 ( .A(n11028), .B(n10816), .Z(n10818) );
  IV U12844 ( .A(n10918), .Z(n10816) );
  XOR U12845 ( .A(n11029), .B(n11030), .Z(n10918) );
  AND U12846 ( .A(n11031), .B(n11032), .Z(n11029) );
  AND U12847 ( .A(a[54]), .B(b[14]), .Z(n11028) );
  XOR U12848 ( .A(n11033), .B(n10821), .Z(n10823) );
  IV U12849 ( .A(n10916), .Z(n10821) );
  XOR U12850 ( .A(n11034), .B(n11035), .Z(n10916) );
  AND U12851 ( .A(n11036), .B(n11037), .Z(n11034) );
  AND U12852 ( .A(a[55]), .B(b[13]), .Z(n11033) );
  XOR U12853 ( .A(n11038), .B(n10826), .Z(n10828) );
  IV U12854 ( .A(n10914), .Z(n10826) );
  XOR U12855 ( .A(n11039), .B(n11040), .Z(n10914) );
  AND U12856 ( .A(n11041), .B(n11042), .Z(n11039) );
  AND U12857 ( .A(a[56]), .B(b[12]), .Z(n11038) );
  XOR U12858 ( .A(n11043), .B(n10831), .Z(n10833) );
  IV U12859 ( .A(n10912), .Z(n10831) );
  XOR U12860 ( .A(n11044), .B(n11045), .Z(n10912) );
  AND U12861 ( .A(n11046), .B(n11047), .Z(n11044) );
  AND U12862 ( .A(a[57]), .B(b[11]), .Z(n11043) );
  XOR U12863 ( .A(n11048), .B(n10836), .Z(n10838) );
  IV U12864 ( .A(n10910), .Z(n10836) );
  XOR U12865 ( .A(n11049), .B(n11050), .Z(n10910) );
  AND U12866 ( .A(n11051), .B(n11052), .Z(n11049) );
  AND U12867 ( .A(a[58]), .B(b[10]), .Z(n11048) );
  XOR U12868 ( .A(n11053), .B(n10841), .Z(n10843) );
  IV U12869 ( .A(n10908), .Z(n10841) );
  XOR U12870 ( .A(n11054), .B(n11055), .Z(n10908) );
  AND U12871 ( .A(n11056), .B(n11057), .Z(n11054) );
  AND U12872 ( .A(a[59]), .B(b[9]), .Z(n11053) );
  XOR U12873 ( .A(n11058), .B(n10846), .Z(n10848) );
  IV U12874 ( .A(n10906), .Z(n10846) );
  XOR U12875 ( .A(n11059), .B(n11060), .Z(n10906) );
  AND U12876 ( .A(n11061), .B(n11062), .Z(n11059) );
  AND U12877 ( .A(a[60]), .B(b[8]), .Z(n11058) );
  XOR U12878 ( .A(n11063), .B(n10851), .Z(n10853) );
  IV U12879 ( .A(n10904), .Z(n10851) );
  XOR U12880 ( .A(n11064), .B(n11065), .Z(n10904) );
  AND U12881 ( .A(n11066), .B(n11067), .Z(n11064) );
  AND U12882 ( .A(a[61]), .B(b[7]), .Z(n11063) );
  XOR U12883 ( .A(n11068), .B(n10856), .Z(n10858) );
  IV U12884 ( .A(n10902), .Z(n10856) );
  XOR U12885 ( .A(n11069), .B(n11070), .Z(n10902) );
  AND U12886 ( .A(n11071), .B(n11072), .Z(n11069) );
  AND U12887 ( .A(a[62]), .B(b[6]), .Z(n11068) );
  XOR U12888 ( .A(n11073), .B(n10861), .Z(n10863) );
  IV U12889 ( .A(n10900), .Z(n10861) );
  XOR U12890 ( .A(n11074), .B(n11075), .Z(n10900) );
  AND U12891 ( .A(n11076), .B(n11077), .Z(n11074) );
  AND U12892 ( .A(a[63]), .B(b[5]), .Z(n11073) );
  XOR U12893 ( .A(n11078), .B(n10866), .Z(n10868) );
  IV U12894 ( .A(n10898), .Z(n10866) );
  XOR U12895 ( .A(n11079), .B(n11080), .Z(n10898) );
  AND U12896 ( .A(n11081), .B(n11082), .Z(n11079) );
  AND U12897 ( .A(a[64]), .B(b[4]), .Z(n11078) );
  XOR U12898 ( .A(n11083), .B(n10871), .Z(n10873) );
  IV U12899 ( .A(n10896), .Z(n10871) );
  XOR U12900 ( .A(n11084), .B(n11085), .Z(n10896) );
  AND U12901 ( .A(n10891), .B(n10889), .Z(n11084) );
  AND U12902 ( .A(b[2]), .B(a[65]), .Z(n11086) );
  XOR U12903 ( .A(n11081), .B(n11085), .Z(n11087) );
  XOR U12904 ( .A(n11088), .B(n11089), .Z(n11085) );
  NANDN U12905 ( .A(n10894), .B(n10893), .Z(n11089) );
  XOR U12906 ( .A(n11090), .B(n11091), .Z(n10893) );
  NAND U12907 ( .A(a[65]), .B(b[1]), .Z(n11091) );
  XOR U12908 ( .A(n11092), .B(n11093), .Z(n10894) );
  XOR U12909 ( .A(n11090), .B(n11094), .Z(n11093) );
  IV U12910 ( .A(n11088), .Z(n11090) );
  ANDN U12911 ( .B(n5227), .A(n5229), .Z(n11088) );
  NAND U12912 ( .A(a[65]), .B(b[0]), .Z(n5229) );
  XNOR U12913 ( .A(n11095), .B(n11096), .Z(n5227) );
  XOR U12914 ( .A(n11076), .B(n11080), .Z(n11097) );
  XOR U12915 ( .A(n11071), .B(n11075), .Z(n11098) );
  XOR U12916 ( .A(n11066), .B(n11070), .Z(n11099) );
  XOR U12917 ( .A(n11061), .B(n11065), .Z(n11100) );
  XOR U12918 ( .A(n11056), .B(n11060), .Z(n11101) );
  XOR U12919 ( .A(n11051), .B(n11055), .Z(n11102) );
  XOR U12920 ( .A(n11046), .B(n11050), .Z(n11103) );
  XOR U12921 ( .A(n11041), .B(n11045), .Z(n11104) );
  XOR U12922 ( .A(n11036), .B(n11040), .Z(n11105) );
  XOR U12923 ( .A(n11031), .B(n11035), .Z(n11106) );
  XOR U12924 ( .A(n11026), .B(n11030), .Z(n11107) );
  XOR U12925 ( .A(n11021), .B(n11025), .Z(n11108) );
  XOR U12926 ( .A(n11016), .B(n11020), .Z(n11109) );
  XOR U12927 ( .A(n11011), .B(n11015), .Z(n11110) );
  XOR U12928 ( .A(n11006), .B(n11010), .Z(n11111) );
  XOR U12929 ( .A(n11001), .B(n11005), .Z(n11112) );
  XOR U12930 ( .A(n10996), .B(n11000), .Z(n11113) );
  XOR U12931 ( .A(n10991), .B(n10995), .Z(n11114) );
  XOR U12932 ( .A(n10986), .B(n10990), .Z(n11115) );
  XOR U12933 ( .A(n10981), .B(n10985), .Z(n11116) );
  XOR U12934 ( .A(n10976), .B(n10980), .Z(n11117) );
  XOR U12935 ( .A(n10971), .B(n10975), .Z(n11118) );
  XOR U12936 ( .A(n10966), .B(n10970), .Z(n11119) );
  XOR U12937 ( .A(n10961), .B(n10965), .Z(n11120) );
  XNOR U12938 ( .A(n10957), .B(n10960), .Z(n11121) );
  XOR U12939 ( .A(n11122), .B(n11123), .Z(n10957) );
  XOR U12940 ( .A(n11124), .B(n11125), .Z(n11123) );
  XNOR U12941 ( .A(n11126), .B(n11127), .Z(n11124) );
  XOR U12942 ( .A(n11128), .B(n11129), .Z(n11127) );
  AND U12943 ( .A(b[30]), .B(a[37]), .Z(n11129) );
  AND U12944 ( .A(a[36]), .B(b[31]), .Z(n11128) );
  XNOR U12945 ( .A(n11130), .B(n11126), .Z(n11122) );
  XNOR U12946 ( .A(n11131), .B(n11132), .Z(n11126) );
  ANDN U12947 ( .B(n11133), .A(n11134), .Z(n11131) );
  AND U12948 ( .A(a[38]), .B(b[29]), .Z(n11130) );
  XOR U12949 ( .A(n11135), .B(n10955), .Z(n10956) );
  IV U12950 ( .A(n11125), .Z(n10955) );
  XOR U12951 ( .A(n11136), .B(n11137), .Z(n11125) );
  AND U12952 ( .A(n11138), .B(n11139), .Z(n11136) );
  AND U12953 ( .A(a[39]), .B(b[28]), .Z(n11135) );
  XOR U12954 ( .A(n11141), .B(n11142), .Z(n10960) );
  AND U12955 ( .A(n11143), .B(n11144), .Z(n11141) );
  AND U12956 ( .A(a[40]), .B(b[27]), .Z(n11140) );
  XOR U12957 ( .A(n11146), .B(n11147), .Z(n10965) );
  AND U12958 ( .A(n11148), .B(n11149), .Z(n11146) );
  AND U12959 ( .A(a[41]), .B(b[26]), .Z(n11145) );
  XOR U12960 ( .A(n11151), .B(n11152), .Z(n10970) );
  AND U12961 ( .A(n11153), .B(n11154), .Z(n11151) );
  AND U12962 ( .A(a[42]), .B(b[25]), .Z(n11150) );
  XOR U12963 ( .A(n11156), .B(n11157), .Z(n10975) );
  AND U12964 ( .A(n11158), .B(n11159), .Z(n11156) );
  AND U12965 ( .A(a[43]), .B(b[24]), .Z(n11155) );
  XOR U12966 ( .A(n11161), .B(n11162), .Z(n10980) );
  AND U12967 ( .A(n11163), .B(n11164), .Z(n11161) );
  AND U12968 ( .A(a[44]), .B(b[23]), .Z(n11160) );
  XOR U12969 ( .A(n11166), .B(n11167), .Z(n10985) );
  AND U12970 ( .A(n11168), .B(n11169), .Z(n11166) );
  AND U12971 ( .A(a[45]), .B(b[22]), .Z(n11165) );
  XOR U12972 ( .A(n11171), .B(n11172), .Z(n10990) );
  AND U12973 ( .A(n11173), .B(n11174), .Z(n11171) );
  AND U12974 ( .A(a[46]), .B(b[21]), .Z(n11170) );
  XOR U12975 ( .A(n11176), .B(n11177), .Z(n10995) );
  AND U12976 ( .A(n11178), .B(n11179), .Z(n11176) );
  AND U12977 ( .A(a[47]), .B(b[20]), .Z(n11175) );
  XOR U12978 ( .A(n11181), .B(n11182), .Z(n11000) );
  AND U12979 ( .A(n11183), .B(n11184), .Z(n11181) );
  AND U12980 ( .A(a[48]), .B(b[19]), .Z(n11180) );
  XOR U12981 ( .A(n11186), .B(n11187), .Z(n11005) );
  AND U12982 ( .A(n11188), .B(n11189), .Z(n11186) );
  AND U12983 ( .A(a[49]), .B(b[18]), .Z(n11185) );
  XOR U12984 ( .A(n11191), .B(n11192), .Z(n11010) );
  AND U12985 ( .A(n11193), .B(n11194), .Z(n11191) );
  AND U12986 ( .A(a[50]), .B(b[17]), .Z(n11190) );
  XOR U12987 ( .A(n11196), .B(n11197), .Z(n11015) );
  AND U12988 ( .A(n11198), .B(n11199), .Z(n11196) );
  AND U12989 ( .A(a[51]), .B(b[16]), .Z(n11195) );
  XOR U12990 ( .A(n11201), .B(n11202), .Z(n11020) );
  AND U12991 ( .A(n11203), .B(n11204), .Z(n11201) );
  AND U12992 ( .A(a[52]), .B(b[15]), .Z(n11200) );
  XOR U12993 ( .A(n11206), .B(n11207), .Z(n11025) );
  AND U12994 ( .A(n11208), .B(n11209), .Z(n11206) );
  AND U12995 ( .A(a[53]), .B(b[14]), .Z(n11205) );
  XOR U12996 ( .A(n11211), .B(n11212), .Z(n11030) );
  AND U12997 ( .A(n11213), .B(n11214), .Z(n11211) );
  AND U12998 ( .A(a[54]), .B(b[13]), .Z(n11210) );
  XOR U12999 ( .A(n11216), .B(n11217), .Z(n11035) );
  AND U13000 ( .A(n11218), .B(n11219), .Z(n11216) );
  AND U13001 ( .A(a[55]), .B(b[12]), .Z(n11215) );
  XOR U13002 ( .A(n11221), .B(n11222), .Z(n11040) );
  AND U13003 ( .A(n11223), .B(n11224), .Z(n11221) );
  AND U13004 ( .A(a[56]), .B(b[11]), .Z(n11220) );
  XOR U13005 ( .A(n11226), .B(n11227), .Z(n11045) );
  AND U13006 ( .A(n11228), .B(n11229), .Z(n11226) );
  AND U13007 ( .A(a[57]), .B(b[10]), .Z(n11225) );
  XOR U13008 ( .A(n11231), .B(n11232), .Z(n11050) );
  AND U13009 ( .A(n11233), .B(n11234), .Z(n11231) );
  AND U13010 ( .A(a[58]), .B(b[9]), .Z(n11230) );
  XOR U13011 ( .A(n11236), .B(n11237), .Z(n11055) );
  AND U13012 ( .A(n11238), .B(n11239), .Z(n11236) );
  AND U13013 ( .A(a[59]), .B(b[8]), .Z(n11235) );
  XOR U13014 ( .A(n11241), .B(n11242), .Z(n11060) );
  AND U13015 ( .A(n11243), .B(n11244), .Z(n11241) );
  AND U13016 ( .A(a[60]), .B(b[7]), .Z(n11240) );
  XOR U13017 ( .A(n11246), .B(n11247), .Z(n11065) );
  AND U13018 ( .A(n11248), .B(n11249), .Z(n11246) );
  AND U13019 ( .A(a[61]), .B(b[6]), .Z(n11245) );
  XOR U13020 ( .A(n11251), .B(n11252), .Z(n11070) );
  AND U13021 ( .A(n11253), .B(n11254), .Z(n11251) );
  AND U13022 ( .A(a[62]), .B(b[5]), .Z(n11250) );
  XOR U13023 ( .A(n11256), .B(n11257), .Z(n11075) );
  AND U13024 ( .A(n11258), .B(n11259), .Z(n11256) );
  AND U13025 ( .A(a[63]), .B(b[4]), .Z(n11255) );
  XOR U13026 ( .A(n11261), .B(n11262), .Z(n11080) );
  AND U13027 ( .A(n11094), .B(n11092), .Z(n11261) );
  AND U13028 ( .A(b[2]), .B(a[64]), .Z(n11263) );
  XOR U13029 ( .A(n11258), .B(n11262), .Z(n11264) );
  XOR U13030 ( .A(n11265), .B(n11266), .Z(n11262) );
  NANDN U13031 ( .A(n11096), .B(n11095), .Z(n11266) );
  XOR U13032 ( .A(n11267), .B(n11268), .Z(n11095) );
  NAND U13033 ( .A(a[64]), .B(b[1]), .Z(n11268) );
  XOR U13034 ( .A(n11269), .B(n11270), .Z(n11096) );
  XOR U13035 ( .A(n11267), .B(n11271), .Z(n11270) );
  IV U13036 ( .A(n11265), .Z(n11267) );
  ANDN U13037 ( .B(n5232), .A(n5234), .Z(n11265) );
  NAND U13038 ( .A(a[64]), .B(b[0]), .Z(n5234) );
  XNOR U13039 ( .A(n11272), .B(n11273), .Z(n5232) );
  XOR U13040 ( .A(n11253), .B(n11257), .Z(n11274) );
  XOR U13041 ( .A(n11248), .B(n11252), .Z(n11275) );
  XOR U13042 ( .A(n11243), .B(n11247), .Z(n11276) );
  XOR U13043 ( .A(n11238), .B(n11242), .Z(n11277) );
  XOR U13044 ( .A(n11233), .B(n11237), .Z(n11278) );
  XOR U13045 ( .A(n11228), .B(n11232), .Z(n11279) );
  XOR U13046 ( .A(n11223), .B(n11227), .Z(n11280) );
  XOR U13047 ( .A(n11218), .B(n11222), .Z(n11281) );
  XOR U13048 ( .A(n11213), .B(n11217), .Z(n11282) );
  XOR U13049 ( .A(n11208), .B(n11212), .Z(n11283) );
  XOR U13050 ( .A(n11203), .B(n11207), .Z(n11284) );
  XOR U13051 ( .A(n11198), .B(n11202), .Z(n11285) );
  XOR U13052 ( .A(n11193), .B(n11197), .Z(n11286) );
  XOR U13053 ( .A(n11188), .B(n11192), .Z(n11287) );
  XOR U13054 ( .A(n11183), .B(n11187), .Z(n11288) );
  XOR U13055 ( .A(n11178), .B(n11182), .Z(n11289) );
  XOR U13056 ( .A(n11173), .B(n11177), .Z(n11290) );
  XOR U13057 ( .A(n11168), .B(n11172), .Z(n11291) );
  XOR U13058 ( .A(n11163), .B(n11167), .Z(n11292) );
  XOR U13059 ( .A(n11158), .B(n11162), .Z(n11293) );
  XOR U13060 ( .A(n11153), .B(n11157), .Z(n11294) );
  XOR U13061 ( .A(n11148), .B(n11152), .Z(n11295) );
  XOR U13062 ( .A(n11143), .B(n11147), .Z(n11296) );
  XOR U13063 ( .A(n11138), .B(n11142), .Z(n11297) );
  XNOR U13064 ( .A(n11134), .B(n11137), .Z(n11298) );
  XOR U13065 ( .A(n11299), .B(n11300), .Z(n11134) );
  XOR U13066 ( .A(n11301), .B(n11302), .Z(n11300) );
  XOR U13067 ( .A(n11303), .B(n11304), .Z(n11301) );
  AND U13068 ( .A(b[29]), .B(a[37]), .Z(n11303) );
  XOR U13069 ( .A(n11304), .B(n11305), .Z(n11299) );
  XOR U13070 ( .A(n11306), .B(n11307), .Z(n11305) );
  AND U13071 ( .A(a[36]), .B(b[30]), .Z(n11307) );
  AND U13072 ( .A(a[35]), .B(b[31]), .Z(n11306) );
  XOR U13073 ( .A(n11308), .B(n11309), .Z(n11304) );
  ANDN U13074 ( .B(n11310), .A(n11311), .Z(n11308) );
  XOR U13075 ( .A(n11312), .B(n11132), .Z(n11133) );
  IV U13076 ( .A(n11302), .Z(n11132) );
  XOR U13077 ( .A(n11313), .B(n11314), .Z(n11302) );
  ANDN U13078 ( .B(n11315), .A(n11316), .Z(n11313) );
  AND U13079 ( .A(a[38]), .B(b[28]), .Z(n11312) );
  XOR U13080 ( .A(n11318), .B(n11319), .Z(n11137) );
  AND U13081 ( .A(n11320), .B(n11321), .Z(n11318) );
  AND U13082 ( .A(a[39]), .B(b[27]), .Z(n11317) );
  XOR U13083 ( .A(n11323), .B(n11324), .Z(n11142) );
  AND U13084 ( .A(n11325), .B(n11326), .Z(n11323) );
  AND U13085 ( .A(a[40]), .B(b[26]), .Z(n11322) );
  XOR U13086 ( .A(n11328), .B(n11329), .Z(n11147) );
  AND U13087 ( .A(n11330), .B(n11331), .Z(n11328) );
  AND U13088 ( .A(a[41]), .B(b[25]), .Z(n11327) );
  XOR U13089 ( .A(n11333), .B(n11334), .Z(n11152) );
  AND U13090 ( .A(n11335), .B(n11336), .Z(n11333) );
  AND U13091 ( .A(a[42]), .B(b[24]), .Z(n11332) );
  XOR U13092 ( .A(n11338), .B(n11339), .Z(n11157) );
  AND U13093 ( .A(n11340), .B(n11341), .Z(n11338) );
  AND U13094 ( .A(a[43]), .B(b[23]), .Z(n11337) );
  XOR U13095 ( .A(n11343), .B(n11344), .Z(n11162) );
  AND U13096 ( .A(n11345), .B(n11346), .Z(n11343) );
  AND U13097 ( .A(a[44]), .B(b[22]), .Z(n11342) );
  XOR U13098 ( .A(n11348), .B(n11349), .Z(n11167) );
  AND U13099 ( .A(n11350), .B(n11351), .Z(n11348) );
  AND U13100 ( .A(a[45]), .B(b[21]), .Z(n11347) );
  XOR U13101 ( .A(n11353), .B(n11354), .Z(n11172) );
  AND U13102 ( .A(n11355), .B(n11356), .Z(n11353) );
  AND U13103 ( .A(a[46]), .B(b[20]), .Z(n11352) );
  XOR U13104 ( .A(n11358), .B(n11359), .Z(n11177) );
  AND U13105 ( .A(n11360), .B(n11361), .Z(n11358) );
  AND U13106 ( .A(a[47]), .B(b[19]), .Z(n11357) );
  XOR U13107 ( .A(n11363), .B(n11364), .Z(n11182) );
  AND U13108 ( .A(n11365), .B(n11366), .Z(n11363) );
  AND U13109 ( .A(a[48]), .B(b[18]), .Z(n11362) );
  XOR U13110 ( .A(n11368), .B(n11369), .Z(n11187) );
  AND U13111 ( .A(n11370), .B(n11371), .Z(n11368) );
  AND U13112 ( .A(a[49]), .B(b[17]), .Z(n11367) );
  XOR U13113 ( .A(n11373), .B(n11374), .Z(n11192) );
  AND U13114 ( .A(n11375), .B(n11376), .Z(n11373) );
  AND U13115 ( .A(a[50]), .B(b[16]), .Z(n11372) );
  XOR U13116 ( .A(n11378), .B(n11379), .Z(n11197) );
  AND U13117 ( .A(n11380), .B(n11381), .Z(n11378) );
  AND U13118 ( .A(a[51]), .B(b[15]), .Z(n11377) );
  XOR U13119 ( .A(n11383), .B(n11384), .Z(n11202) );
  AND U13120 ( .A(n11385), .B(n11386), .Z(n11383) );
  AND U13121 ( .A(a[52]), .B(b[14]), .Z(n11382) );
  XOR U13122 ( .A(n11388), .B(n11389), .Z(n11207) );
  AND U13123 ( .A(n11390), .B(n11391), .Z(n11388) );
  AND U13124 ( .A(a[53]), .B(b[13]), .Z(n11387) );
  XOR U13125 ( .A(n11393), .B(n11394), .Z(n11212) );
  AND U13126 ( .A(n11395), .B(n11396), .Z(n11393) );
  AND U13127 ( .A(a[54]), .B(b[12]), .Z(n11392) );
  XOR U13128 ( .A(n11398), .B(n11399), .Z(n11217) );
  AND U13129 ( .A(n11400), .B(n11401), .Z(n11398) );
  AND U13130 ( .A(a[55]), .B(b[11]), .Z(n11397) );
  XOR U13131 ( .A(n11403), .B(n11404), .Z(n11222) );
  AND U13132 ( .A(n11405), .B(n11406), .Z(n11403) );
  AND U13133 ( .A(a[56]), .B(b[10]), .Z(n11402) );
  XOR U13134 ( .A(n11408), .B(n11409), .Z(n11227) );
  AND U13135 ( .A(n11410), .B(n11411), .Z(n11408) );
  AND U13136 ( .A(a[57]), .B(b[9]), .Z(n11407) );
  XOR U13137 ( .A(n11413), .B(n11414), .Z(n11232) );
  AND U13138 ( .A(n11415), .B(n11416), .Z(n11413) );
  AND U13139 ( .A(a[58]), .B(b[8]), .Z(n11412) );
  XOR U13140 ( .A(n11418), .B(n11419), .Z(n11237) );
  AND U13141 ( .A(n11420), .B(n11421), .Z(n11418) );
  AND U13142 ( .A(a[59]), .B(b[7]), .Z(n11417) );
  XOR U13143 ( .A(n11423), .B(n11424), .Z(n11242) );
  AND U13144 ( .A(n11425), .B(n11426), .Z(n11423) );
  AND U13145 ( .A(a[60]), .B(b[6]), .Z(n11422) );
  XOR U13146 ( .A(n11428), .B(n11429), .Z(n11247) );
  AND U13147 ( .A(n11430), .B(n11431), .Z(n11428) );
  AND U13148 ( .A(a[61]), .B(b[5]), .Z(n11427) );
  XOR U13149 ( .A(n11433), .B(n11434), .Z(n11252) );
  AND U13150 ( .A(n11435), .B(n11436), .Z(n11433) );
  AND U13151 ( .A(a[62]), .B(b[4]), .Z(n11432) );
  XOR U13152 ( .A(n11438), .B(n11439), .Z(n11257) );
  AND U13153 ( .A(n11271), .B(n11269), .Z(n11438) );
  AND U13154 ( .A(b[2]), .B(a[63]), .Z(n11440) );
  XOR U13155 ( .A(n11435), .B(n11439), .Z(n11441) );
  XOR U13156 ( .A(n11442), .B(n11443), .Z(n11439) );
  NANDN U13157 ( .A(n11273), .B(n11272), .Z(n11443) );
  XOR U13158 ( .A(n11444), .B(n11445), .Z(n11272) );
  NAND U13159 ( .A(a[63]), .B(b[1]), .Z(n11445) );
  XOR U13160 ( .A(n11446), .B(n11447), .Z(n11273) );
  XOR U13161 ( .A(n11444), .B(n11448), .Z(n11447) );
  IV U13162 ( .A(n11442), .Z(n11444) );
  ANDN U13163 ( .B(n5237), .A(n5239), .Z(n11442) );
  NAND U13164 ( .A(a[63]), .B(b[0]), .Z(n5239) );
  XNOR U13165 ( .A(n11449), .B(n11450), .Z(n5237) );
  XOR U13166 ( .A(n11430), .B(n11434), .Z(n11451) );
  XOR U13167 ( .A(n11425), .B(n11429), .Z(n11452) );
  XOR U13168 ( .A(n11420), .B(n11424), .Z(n11453) );
  XOR U13169 ( .A(n11415), .B(n11419), .Z(n11454) );
  XOR U13170 ( .A(n11410), .B(n11414), .Z(n11455) );
  XOR U13171 ( .A(n11405), .B(n11409), .Z(n11456) );
  XOR U13172 ( .A(n11400), .B(n11404), .Z(n11457) );
  XOR U13173 ( .A(n11395), .B(n11399), .Z(n11458) );
  XOR U13174 ( .A(n11390), .B(n11394), .Z(n11459) );
  XOR U13175 ( .A(n11385), .B(n11389), .Z(n11460) );
  XOR U13176 ( .A(n11380), .B(n11384), .Z(n11461) );
  XOR U13177 ( .A(n11375), .B(n11379), .Z(n11462) );
  XOR U13178 ( .A(n11370), .B(n11374), .Z(n11463) );
  XOR U13179 ( .A(n11365), .B(n11369), .Z(n11464) );
  XOR U13180 ( .A(n11360), .B(n11364), .Z(n11465) );
  XOR U13181 ( .A(n11355), .B(n11359), .Z(n11466) );
  XOR U13182 ( .A(n11350), .B(n11354), .Z(n11467) );
  XOR U13183 ( .A(n11345), .B(n11349), .Z(n11468) );
  XOR U13184 ( .A(n11340), .B(n11344), .Z(n11469) );
  XOR U13185 ( .A(n11335), .B(n11339), .Z(n11470) );
  XOR U13186 ( .A(n11330), .B(n11334), .Z(n11471) );
  XOR U13187 ( .A(n11325), .B(n11329), .Z(n11472) );
  XOR U13188 ( .A(n11320), .B(n11324), .Z(n11473) );
  XNOR U13189 ( .A(n11316), .B(n11319), .Z(n11474) );
  XNOR U13190 ( .A(n11311), .B(n11475), .Z(n11316) );
  XOR U13191 ( .A(n11310), .B(n11314), .Z(n11475) );
  XOR U13192 ( .A(n11476), .B(n11309), .Z(n11310) );
  AND U13193 ( .A(b[28]), .B(a[37]), .Z(n11476) );
  XOR U13194 ( .A(n11477), .B(n11478), .Z(n11311) );
  XOR U13195 ( .A(n11309), .B(n11479), .Z(n11478) );
  XOR U13196 ( .A(n11480), .B(n11481), .Z(n11479) );
  XOR U13197 ( .A(n11482), .B(n11483), .Z(n11481) );
  NAND U13198 ( .A(a[35]), .B(b[30]), .Z(n11483) );
  AND U13199 ( .A(a[34]), .B(b[31]), .Z(n11482) );
  XOR U13200 ( .A(n11484), .B(n11485), .Z(n11309) );
  AND U13201 ( .A(n11486), .B(n11487), .Z(n11484) );
  XOR U13202 ( .A(n11488), .B(n11480), .Z(n11477) );
  XOR U13203 ( .A(n11489), .B(n11490), .Z(n11480) );
  ANDN U13204 ( .B(n11491), .A(n11492), .Z(n11489) );
  AND U13205 ( .A(a[36]), .B(b[29]), .Z(n11488) );
  XOR U13206 ( .A(n11494), .B(n11495), .Z(n11314) );
  AND U13207 ( .A(n11496), .B(n11497), .Z(n11494) );
  AND U13208 ( .A(a[38]), .B(b[27]), .Z(n11493) );
  XOR U13209 ( .A(n11499), .B(n11500), .Z(n11319) );
  AND U13210 ( .A(n11501), .B(n11502), .Z(n11499) );
  AND U13211 ( .A(a[39]), .B(b[26]), .Z(n11498) );
  XOR U13212 ( .A(n11504), .B(n11505), .Z(n11324) );
  AND U13213 ( .A(n11506), .B(n11507), .Z(n11504) );
  AND U13214 ( .A(a[40]), .B(b[25]), .Z(n11503) );
  XOR U13215 ( .A(n11509), .B(n11510), .Z(n11329) );
  AND U13216 ( .A(n11511), .B(n11512), .Z(n11509) );
  AND U13217 ( .A(a[41]), .B(b[24]), .Z(n11508) );
  XOR U13218 ( .A(n11514), .B(n11515), .Z(n11334) );
  AND U13219 ( .A(n11516), .B(n11517), .Z(n11514) );
  AND U13220 ( .A(a[42]), .B(b[23]), .Z(n11513) );
  XOR U13221 ( .A(n11519), .B(n11520), .Z(n11339) );
  AND U13222 ( .A(n11521), .B(n11522), .Z(n11519) );
  AND U13223 ( .A(a[43]), .B(b[22]), .Z(n11518) );
  XOR U13224 ( .A(n11524), .B(n11525), .Z(n11344) );
  AND U13225 ( .A(n11526), .B(n11527), .Z(n11524) );
  AND U13226 ( .A(a[44]), .B(b[21]), .Z(n11523) );
  XOR U13227 ( .A(n11529), .B(n11530), .Z(n11349) );
  AND U13228 ( .A(n11531), .B(n11532), .Z(n11529) );
  AND U13229 ( .A(a[45]), .B(b[20]), .Z(n11528) );
  XOR U13230 ( .A(n11534), .B(n11535), .Z(n11354) );
  AND U13231 ( .A(n11536), .B(n11537), .Z(n11534) );
  AND U13232 ( .A(a[46]), .B(b[19]), .Z(n11533) );
  XOR U13233 ( .A(n11539), .B(n11540), .Z(n11359) );
  AND U13234 ( .A(n11541), .B(n11542), .Z(n11539) );
  AND U13235 ( .A(a[47]), .B(b[18]), .Z(n11538) );
  XOR U13236 ( .A(n11544), .B(n11545), .Z(n11364) );
  AND U13237 ( .A(n11546), .B(n11547), .Z(n11544) );
  AND U13238 ( .A(a[48]), .B(b[17]), .Z(n11543) );
  XOR U13239 ( .A(n11549), .B(n11550), .Z(n11369) );
  AND U13240 ( .A(n11551), .B(n11552), .Z(n11549) );
  AND U13241 ( .A(a[49]), .B(b[16]), .Z(n11548) );
  XOR U13242 ( .A(n11554), .B(n11555), .Z(n11374) );
  AND U13243 ( .A(n11556), .B(n11557), .Z(n11554) );
  AND U13244 ( .A(a[50]), .B(b[15]), .Z(n11553) );
  XOR U13245 ( .A(n11559), .B(n11560), .Z(n11379) );
  AND U13246 ( .A(n11561), .B(n11562), .Z(n11559) );
  AND U13247 ( .A(a[51]), .B(b[14]), .Z(n11558) );
  XOR U13248 ( .A(n11564), .B(n11565), .Z(n11384) );
  AND U13249 ( .A(n11566), .B(n11567), .Z(n11564) );
  AND U13250 ( .A(a[52]), .B(b[13]), .Z(n11563) );
  XOR U13251 ( .A(n11569), .B(n11570), .Z(n11389) );
  AND U13252 ( .A(n11571), .B(n11572), .Z(n11569) );
  AND U13253 ( .A(a[53]), .B(b[12]), .Z(n11568) );
  XOR U13254 ( .A(n11574), .B(n11575), .Z(n11394) );
  AND U13255 ( .A(n11576), .B(n11577), .Z(n11574) );
  AND U13256 ( .A(a[54]), .B(b[11]), .Z(n11573) );
  XOR U13257 ( .A(n11579), .B(n11580), .Z(n11399) );
  AND U13258 ( .A(n11581), .B(n11582), .Z(n11579) );
  AND U13259 ( .A(a[55]), .B(b[10]), .Z(n11578) );
  XOR U13260 ( .A(n11584), .B(n11585), .Z(n11404) );
  AND U13261 ( .A(n11586), .B(n11587), .Z(n11584) );
  AND U13262 ( .A(a[56]), .B(b[9]), .Z(n11583) );
  XOR U13263 ( .A(n11589), .B(n11590), .Z(n11409) );
  AND U13264 ( .A(n11591), .B(n11592), .Z(n11589) );
  AND U13265 ( .A(a[57]), .B(b[8]), .Z(n11588) );
  XOR U13266 ( .A(n11594), .B(n11595), .Z(n11414) );
  AND U13267 ( .A(n11596), .B(n11597), .Z(n11594) );
  AND U13268 ( .A(a[58]), .B(b[7]), .Z(n11593) );
  XOR U13269 ( .A(n11599), .B(n11600), .Z(n11419) );
  AND U13270 ( .A(n11601), .B(n11602), .Z(n11599) );
  AND U13271 ( .A(a[59]), .B(b[6]), .Z(n11598) );
  XOR U13272 ( .A(n11604), .B(n11605), .Z(n11424) );
  AND U13273 ( .A(n11606), .B(n11607), .Z(n11604) );
  AND U13274 ( .A(a[60]), .B(b[5]), .Z(n11603) );
  XOR U13275 ( .A(n11609), .B(n11610), .Z(n11429) );
  AND U13276 ( .A(n11611), .B(n11612), .Z(n11609) );
  AND U13277 ( .A(a[61]), .B(b[4]), .Z(n11608) );
  XOR U13278 ( .A(n11614), .B(n11615), .Z(n11434) );
  AND U13279 ( .A(n11448), .B(n11446), .Z(n11614) );
  AND U13280 ( .A(b[2]), .B(a[62]), .Z(n11616) );
  XOR U13281 ( .A(n11611), .B(n11615), .Z(n11617) );
  XOR U13282 ( .A(n11618), .B(n11619), .Z(n11615) );
  NANDN U13283 ( .A(n11450), .B(n11449), .Z(n11619) );
  XOR U13284 ( .A(n11620), .B(n11621), .Z(n11449) );
  NAND U13285 ( .A(a[62]), .B(b[1]), .Z(n11621) );
  XOR U13286 ( .A(n11622), .B(n11623), .Z(n11450) );
  XOR U13287 ( .A(n11620), .B(n11624), .Z(n11623) );
  IV U13288 ( .A(n11618), .Z(n11620) );
  ANDN U13289 ( .B(n5242), .A(n5244), .Z(n11618) );
  NAND U13290 ( .A(a[62]), .B(b[0]), .Z(n5244) );
  XNOR U13291 ( .A(n11625), .B(n11626), .Z(n5242) );
  XOR U13292 ( .A(n11606), .B(n11610), .Z(n11627) );
  XOR U13293 ( .A(n11601), .B(n11605), .Z(n11628) );
  XOR U13294 ( .A(n11596), .B(n11600), .Z(n11629) );
  XOR U13295 ( .A(n11591), .B(n11595), .Z(n11630) );
  XOR U13296 ( .A(n11586), .B(n11590), .Z(n11631) );
  XOR U13297 ( .A(n11581), .B(n11585), .Z(n11632) );
  XOR U13298 ( .A(n11576), .B(n11580), .Z(n11633) );
  XOR U13299 ( .A(n11571), .B(n11575), .Z(n11634) );
  XOR U13300 ( .A(n11566), .B(n11570), .Z(n11635) );
  XOR U13301 ( .A(n11561), .B(n11565), .Z(n11636) );
  XOR U13302 ( .A(n11556), .B(n11560), .Z(n11637) );
  XOR U13303 ( .A(n11551), .B(n11555), .Z(n11638) );
  XOR U13304 ( .A(n11546), .B(n11550), .Z(n11639) );
  XOR U13305 ( .A(n11541), .B(n11545), .Z(n11640) );
  XOR U13306 ( .A(n11536), .B(n11540), .Z(n11641) );
  XOR U13307 ( .A(n11531), .B(n11535), .Z(n11642) );
  XOR U13308 ( .A(n11526), .B(n11530), .Z(n11643) );
  XOR U13309 ( .A(n11521), .B(n11525), .Z(n11644) );
  XOR U13310 ( .A(n11516), .B(n11520), .Z(n11645) );
  XOR U13311 ( .A(n11511), .B(n11515), .Z(n11646) );
  XOR U13312 ( .A(n11506), .B(n11510), .Z(n11647) );
  XOR U13313 ( .A(n11501), .B(n11505), .Z(n11648) );
  XOR U13314 ( .A(n11496), .B(n11500), .Z(n11649) );
  XOR U13315 ( .A(n11486), .B(n11495), .Z(n11650) );
  XOR U13316 ( .A(n11651), .B(n11485), .Z(n11486) );
  AND U13317 ( .A(b[27]), .B(a[37]), .Z(n11651) );
  XOR U13318 ( .A(n11485), .B(n11492), .Z(n11652) );
  XOR U13319 ( .A(n11653), .B(n11654), .Z(n11492) );
  XOR U13320 ( .A(n11490), .B(n11655), .Z(n11654) );
  XOR U13321 ( .A(n11656), .B(n11657), .Z(n11655) );
  XOR U13322 ( .A(n11658), .B(n11659), .Z(n11657) );
  NAND U13323 ( .A(a[34]), .B(b[30]), .Z(n11659) );
  AND U13324 ( .A(a[33]), .B(b[31]), .Z(n11658) );
  XOR U13325 ( .A(n11660), .B(n11656), .Z(n11653) );
  XOR U13326 ( .A(n11661), .B(n11662), .Z(n11656) );
  ANDN U13327 ( .B(n11663), .A(n11664), .Z(n11661) );
  AND U13328 ( .A(a[35]), .B(b[29]), .Z(n11660) );
  XOR U13329 ( .A(n11665), .B(n11666), .Z(n11485) );
  AND U13330 ( .A(n11667), .B(n11668), .Z(n11665) );
  XOR U13331 ( .A(n11669), .B(n11490), .Z(n11491) );
  XOR U13332 ( .A(n11670), .B(n11671), .Z(n11490) );
  AND U13333 ( .A(n11672), .B(n11673), .Z(n11670) );
  AND U13334 ( .A(a[36]), .B(b[28]), .Z(n11669) );
  XOR U13335 ( .A(n11675), .B(n11676), .Z(n11495) );
  AND U13336 ( .A(n11677), .B(n11678), .Z(n11675) );
  AND U13337 ( .A(a[38]), .B(b[26]), .Z(n11674) );
  XOR U13338 ( .A(n11680), .B(n11681), .Z(n11500) );
  AND U13339 ( .A(n11682), .B(n11683), .Z(n11680) );
  AND U13340 ( .A(a[39]), .B(b[25]), .Z(n11679) );
  XOR U13341 ( .A(n11685), .B(n11686), .Z(n11505) );
  AND U13342 ( .A(n11687), .B(n11688), .Z(n11685) );
  AND U13343 ( .A(a[40]), .B(b[24]), .Z(n11684) );
  XOR U13344 ( .A(n11690), .B(n11691), .Z(n11510) );
  AND U13345 ( .A(n11692), .B(n11693), .Z(n11690) );
  AND U13346 ( .A(a[41]), .B(b[23]), .Z(n11689) );
  XOR U13347 ( .A(n11695), .B(n11696), .Z(n11515) );
  AND U13348 ( .A(n11697), .B(n11698), .Z(n11695) );
  AND U13349 ( .A(a[42]), .B(b[22]), .Z(n11694) );
  XOR U13350 ( .A(n11700), .B(n11701), .Z(n11520) );
  AND U13351 ( .A(n11702), .B(n11703), .Z(n11700) );
  AND U13352 ( .A(a[43]), .B(b[21]), .Z(n11699) );
  XOR U13353 ( .A(n11705), .B(n11706), .Z(n11525) );
  AND U13354 ( .A(n11707), .B(n11708), .Z(n11705) );
  AND U13355 ( .A(a[44]), .B(b[20]), .Z(n11704) );
  XOR U13356 ( .A(n11710), .B(n11711), .Z(n11530) );
  AND U13357 ( .A(n11712), .B(n11713), .Z(n11710) );
  AND U13358 ( .A(a[45]), .B(b[19]), .Z(n11709) );
  XOR U13359 ( .A(n11715), .B(n11716), .Z(n11535) );
  AND U13360 ( .A(n11717), .B(n11718), .Z(n11715) );
  AND U13361 ( .A(a[46]), .B(b[18]), .Z(n11714) );
  XOR U13362 ( .A(n11720), .B(n11721), .Z(n11540) );
  AND U13363 ( .A(n11722), .B(n11723), .Z(n11720) );
  AND U13364 ( .A(a[47]), .B(b[17]), .Z(n11719) );
  XOR U13365 ( .A(n11725), .B(n11726), .Z(n11545) );
  AND U13366 ( .A(n11727), .B(n11728), .Z(n11725) );
  AND U13367 ( .A(a[48]), .B(b[16]), .Z(n11724) );
  XOR U13368 ( .A(n11730), .B(n11731), .Z(n11550) );
  AND U13369 ( .A(n11732), .B(n11733), .Z(n11730) );
  AND U13370 ( .A(a[49]), .B(b[15]), .Z(n11729) );
  XOR U13371 ( .A(n11735), .B(n11736), .Z(n11555) );
  AND U13372 ( .A(n11737), .B(n11738), .Z(n11735) );
  AND U13373 ( .A(a[50]), .B(b[14]), .Z(n11734) );
  XOR U13374 ( .A(n11740), .B(n11741), .Z(n11560) );
  AND U13375 ( .A(n11742), .B(n11743), .Z(n11740) );
  AND U13376 ( .A(a[51]), .B(b[13]), .Z(n11739) );
  XOR U13377 ( .A(n11745), .B(n11746), .Z(n11565) );
  AND U13378 ( .A(n11747), .B(n11748), .Z(n11745) );
  AND U13379 ( .A(a[52]), .B(b[12]), .Z(n11744) );
  XOR U13380 ( .A(n11750), .B(n11751), .Z(n11570) );
  AND U13381 ( .A(n11752), .B(n11753), .Z(n11750) );
  AND U13382 ( .A(a[53]), .B(b[11]), .Z(n11749) );
  XOR U13383 ( .A(n11755), .B(n11756), .Z(n11575) );
  AND U13384 ( .A(n11757), .B(n11758), .Z(n11755) );
  AND U13385 ( .A(a[54]), .B(b[10]), .Z(n11754) );
  XOR U13386 ( .A(n11760), .B(n11761), .Z(n11580) );
  AND U13387 ( .A(n11762), .B(n11763), .Z(n11760) );
  AND U13388 ( .A(a[55]), .B(b[9]), .Z(n11759) );
  XOR U13389 ( .A(n11765), .B(n11766), .Z(n11585) );
  AND U13390 ( .A(n11767), .B(n11768), .Z(n11765) );
  AND U13391 ( .A(a[56]), .B(b[8]), .Z(n11764) );
  XOR U13392 ( .A(n11770), .B(n11771), .Z(n11590) );
  AND U13393 ( .A(n11772), .B(n11773), .Z(n11770) );
  AND U13394 ( .A(a[57]), .B(b[7]), .Z(n11769) );
  XOR U13395 ( .A(n11775), .B(n11776), .Z(n11595) );
  AND U13396 ( .A(n11777), .B(n11778), .Z(n11775) );
  AND U13397 ( .A(a[58]), .B(b[6]), .Z(n11774) );
  XOR U13398 ( .A(n11780), .B(n11781), .Z(n11600) );
  AND U13399 ( .A(n11782), .B(n11783), .Z(n11780) );
  AND U13400 ( .A(a[59]), .B(b[5]), .Z(n11779) );
  XOR U13401 ( .A(n11785), .B(n11786), .Z(n11605) );
  AND U13402 ( .A(n11787), .B(n11788), .Z(n11785) );
  AND U13403 ( .A(a[60]), .B(b[4]), .Z(n11784) );
  XOR U13404 ( .A(n11790), .B(n11791), .Z(n11610) );
  AND U13405 ( .A(n11624), .B(n11622), .Z(n11790) );
  AND U13406 ( .A(b[2]), .B(a[61]), .Z(n11792) );
  XOR U13407 ( .A(n11787), .B(n11791), .Z(n11793) );
  XOR U13408 ( .A(n11794), .B(n11795), .Z(n11791) );
  NANDN U13409 ( .A(n11626), .B(n11625), .Z(n11795) );
  XOR U13410 ( .A(n11796), .B(n11797), .Z(n11625) );
  NAND U13411 ( .A(a[61]), .B(b[1]), .Z(n11797) );
  XOR U13412 ( .A(n11798), .B(n11799), .Z(n11626) );
  XOR U13413 ( .A(n11796), .B(n11800), .Z(n11799) );
  IV U13414 ( .A(n11794), .Z(n11796) );
  ANDN U13415 ( .B(n5247), .A(n5249), .Z(n11794) );
  NAND U13416 ( .A(a[61]), .B(b[0]), .Z(n5249) );
  XNOR U13417 ( .A(n11801), .B(n11802), .Z(n5247) );
  XOR U13418 ( .A(n11782), .B(n11786), .Z(n11803) );
  XOR U13419 ( .A(n11777), .B(n11781), .Z(n11804) );
  XOR U13420 ( .A(n11772), .B(n11776), .Z(n11805) );
  XOR U13421 ( .A(n11767), .B(n11771), .Z(n11806) );
  XOR U13422 ( .A(n11762), .B(n11766), .Z(n11807) );
  XOR U13423 ( .A(n11757), .B(n11761), .Z(n11808) );
  XOR U13424 ( .A(n11752), .B(n11756), .Z(n11809) );
  XOR U13425 ( .A(n11747), .B(n11751), .Z(n11810) );
  XOR U13426 ( .A(n11742), .B(n11746), .Z(n11811) );
  XOR U13427 ( .A(n11737), .B(n11741), .Z(n11812) );
  XOR U13428 ( .A(n11732), .B(n11736), .Z(n11813) );
  XOR U13429 ( .A(n11727), .B(n11731), .Z(n11814) );
  XOR U13430 ( .A(n11722), .B(n11726), .Z(n11815) );
  XOR U13431 ( .A(n11717), .B(n11721), .Z(n11816) );
  XOR U13432 ( .A(n11712), .B(n11716), .Z(n11817) );
  XOR U13433 ( .A(n11707), .B(n11711), .Z(n11818) );
  XOR U13434 ( .A(n11702), .B(n11706), .Z(n11819) );
  XOR U13435 ( .A(n11697), .B(n11701), .Z(n11820) );
  XOR U13436 ( .A(n11692), .B(n11696), .Z(n11821) );
  XOR U13437 ( .A(n11687), .B(n11691), .Z(n11822) );
  XOR U13438 ( .A(n11682), .B(n11686), .Z(n11823) );
  XOR U13439 ( .A(n11677), .B(n11681), .Z(n11824) );
  XOR U13440 ( .A(n11667), .B(n11676), .Z(n11825) );
  XOR U13441 ( .A(n11826), .B(n11666), .Z(n11667) );
  AND U13442 ( .A(b[26]), .B(a[37]), .Z(n11826) );
  XNOR U13443 ( .A(n11666), .B(n11672), .Z(n11827) );
  XOR U13444 ( .A(n11671), .B(n11664), .Z(n11828) );
  XOR U13445 ( .A(n11829), .B(n11830), .Z(n11664) );
  XOR U13446 ( .A(n11662), .B(n11831), .Z(n11830) );
  XOR U13447 ( .A(n11832), .B(n11833), .Z(n11831) );
  XOR U13448 ( .A(n11834), .B(n11835), .Z(n11833) );
  NAND U13449 ( .A(a[33]), .B(b[30]), .Z(n11835) );
  AND U13450 ( .A(a[32]), .B(b[31]), .Z(n11834) );
  XOR U13451 ( .A(n11836), .B(n11832), .Z(n11829) );
  XOR U13452 ( .A(n11837), .B(n11838), .Z(n11832) );
  ANDN U13453 ( .B(n11839), .A(n11840), .Z(n11837) );
  AND U13454 ( .A(a[34]), .B(b[29]), .Z(n11836) );
  XOR U13455 ( .A(n11841), .B(n11662), .Z(n11663) );
  XOR U13456 ( .A(n11842), .B(n11843), .Z(n11662) );
  AND U13457 ( .A(n11844), .B(n11845), .Z(n11842) );
  AND U13458 ( .A(a[35]), .B(b[28]), .Z(n11841) );
  XOR U13459 ( .A(n11846), .B(n11847), .Z(n11666) );
  AND U13460 ( .A(n11848), .B(n11849), .Z(n11846) );
  XOR U13461 ( .A(n11850), .B(n11671), .Z(n11673) );
  XOR U13462 ( .A(n11851), .B(n11852), .Z(n11671) );
  AND U13463 ( .A(n11853), .B(n11854), .Z(n11851) );
  AND U13464 ( .A(a[36]), .B(b[27]), .Z(n11850) );
  XOR U13465 ( .A(n11856), .B(n11857), .Z(n11676) );
  AND U13466 ( .A(n11858), .B(n11859), .Z(n11856) );
  AND U13467 ( .A(a[38]), .B(b[25]), .Z(n11855) );
  XOR U13468 ( .A(n11861), .B(n11862), .Z(n11681) );
  AND U13469 ( .A(n11863), .B(n11864), .Z(n11861) );
  AND U13470 ( .A(a[39]), .B(b[24]), .Z(n11860) );
  XOR U13471 ( .A(n11866), .B(n11867), .Z(n11686) );
  AND U13472 ( .A(n11868), .B(n11869), .Z(n11866) );
  AND U13473 ( .A(a[40]), .B(b[23]), .Z(n11865) );
  XOR U13474 ( .A(n11871), .B(n11872), .Z(n11691) );
  AND U13475 ( .A(n11873), .B(n11874), .Z(n11871) );
  AND U13476 ( .A(a[41]), .B(b[22]), .Z(n11870) );
  XOR U13477 ( .A(n11876), .B(n11877), .Z(n11696) );
  AND U13478 ( .A(n11878), .B(n11879), .Z(n11876) );
  AND U13479 ( .A(a[42]), .B(b[21]), .Z(n11875) );
  XOR U13480 ( .A(n11881), .B(n11882), .Z(n11701) );
  AND U13481 ( .A(n11883), .B(n11884), .Z(n11881) );
  AND U13482 ( .A(a[43]), .B(b[20]), .Z(n11880) );
  XOR U13483 ( .A(n11886), .B(n11887), .Z(n11706) );
  AND U13484 ( .A(n11888), .B(n11889), .Z(n11886) );
  AND U13485 ( .A(a[44]), .B(b[19]), .Z(n11885) );
  XOR U13486 ( .A(n11891), .B(n11892), .Z(n11711) );
  AND U13487 ( .A(n11893), .B(n11894), .Z(n11891) );
  AND U13488 ( .A(a[45]), .B(b[18]), .Z(n11890) );
  XOR U13489 ( .A(n11896), .B(n11897), .Z(n11716) );
  AND U13490 ( .A(n11898), .B(n11899), .Z(n11896) );
  AND U13491 ( .A(a[46]), .B(b[17]), .Z(n11895) );
  XOR U13492 ( .A(n11901), .B(n11902), .Z(n11721) );
  AND U13493 ( .A(n11903), .B(n11904), .Z(n11901) );
  AND U13494 ( .A(a[47]), .B(b[16]), .Z(n11900) );
  XOR U13495 ( .A(n11906), .B(n11907), .Z(n11726) );
  AND U13496 ( .A(n11908), .B(n11909), .Z(n11906) );
  AND U13497 ( .A(a[48]), .B(b[15]), .Z(n11905) );
  XOR U13498 ( .A(n11911), .B(n11912), .Z(n11731) );
  AND U13499 ( .A(n11913), .B(n11914), .Z(n11911) );
  AND U13500 ( .A(a[49]), .B(b[14]), .Z(n11910) );
  XOR U13501 ( .A(n11916), .B(n11917), .Z(n11736) );
  AND U13502 ( .A(n11918), .B(n11919), .Z(n11916) );
  AND U13503 ( .A(a[50]), .B(b[13]), .Z(n11915) );
  XOR U13504 ( .A(n11921), .B(n11922), .Z(n11741) );
  AND U13505 ( .A(n11923), .B(n11924), .Z(n11921) );
  AND U13506 ( .A(a[51]), .B(b[12]), .Z(n11920) );
  XOR U13507 ( .A(n11926), .B(n11927), .Z(n11746) );
  AND U13508 ( .A(n11928), .B(n11929), .Z(n11926) );
  AND U13509 ( .A(a[52]), .B(b[11]), .Z(n11925) );
  XOR U13510 ( .A(n11931), .B(n11932), .Z(n11751) );
  AND U13511 ( .A(n11933), .B(n11934), .Z(n11931) );
  AND U13512 ( .A(a[53]), .B(b[10]), .Z(n11930) );
  XOR U13513 ( .A(n11936), .B(n11937), .Z(n11756) );
  AND U13514 ( .A(n11938), .B(n11939), .Z(n11936) );
  AND U13515 ( .A(a[54]), .B(b[9]), .Z(n11935) );
  XOR U13516 ( .A(n11941), .B(n11942), .Z(n11761) );
  AND U13517 ( .A(n11943), .B(n11944), .Z(n11941) );
  AND U13518 ( .A(a[55]), .B(b[8]), .Z(n11940) );
  XOR U13519 ( .A(n11946), .B(n11947), .Z(n11766) );
  AND U13520 ( .A(n11948), .B(n11949), .Z(n11946) );
  AND U13521 ( .A(a[56]), .B(b[7]), .Z(n11945) );
  XOR U13522 ( .A(n11951), .B(n11952), .Z(n11771) );
  AND U13523 ( .A(n11953), .B(n11954), .Z(n11951) );
  AND U13524 ( .A(a[57]), .B(b[6]), .Z(n11950) );
  XOR U13525 ( .A(n11956), .B(n11957), .Z(n11776) );
  AND U13526 ( .A(n11958), .B(n11959), .Z(n11956) );
  AND U13527 ( .A(a[58]), .B(b[5]), .Z(n11955) );
  XOR U13528 ( .A(n11961), .B(n11962), .Z(n11781) );
  AND U13529 ( .A(n11963), .B(n11964), .Z(n11961) );
  AND U13530 ( .A(a[59]), .B(b[4]), .Z(n11960) );
  XOR U13531 ( .A(n11966), .B(n11967), .Z(n11786) );
  AND U13532 ( .A(n11800), .B(n11798), .Z(n11966) );
  AND U13533 ( .A(b[2]), .B(a[60]), .Z(n11968) );
  XOR U13534 ( .A(n11963), .B(n11967), .Z(n11969) );
  XOR U13535 ( .A(n11970), .B(n11971), .Z(n11967) );
  NANDN U13536 ( .A(n11802), .B(n11801), .Z(n11971) );
  XOR U13537 ( .A(n11972), .B(n11973), .Z(n11801) );
  NAND U13538 ( .A(a[60]), .B(b[1]), .Z(n11973) );
  XOR U13539 ( .A(n11974), .B(n11975), .Z(n11802) );
  XOR U13540 ( .A(n11972), .B(n11976), .Z(n11975) );
  IV U13541 ( .A(n11970), .Z(n11972) );
  ANDN U13542 ( .B(n5252), .A(n5254), .Z(n11970) );
  NAND U13543 ( .A(a[60]), .B(b[0]), .Z(n5254) );
  XNOR U13544 ( .A(n11977), .B(n11978), .Z(n5252) );
  XOR U13545 ( .A(n11958), .B(n11962), .Z(n11979) );
  XOR U13546 ( .A(n11953), .B(n11957), .Z(n11980) );
  XOR U13547 ( .A(n11948), .B(n11952), .Z(n11981) );
  XOR U13548 ( .A(n11943), .B(n11947), .Z(n11982) );
  XOR U13549 ( .A(n11938), .B(n11942), .Z(n11983) );
  XOR U13550 ( .A(n11933), .B(n11937), .Z(n11984) );
  XOR U13551 ( .A(n11928), .B(n11932), .Z(n11985) );
  XOR U13552 ( .A(n11923), .B(n11927), .Z(n11986) );
  XOR U13553 ( .A(n11918), .B(n11922), .Z(n11987) );
  XOR U13554 ( .A(n11913), .B(n11917), .Z(n11988) );
  XOR U13555 ( .A(n11908), .B(n11912), .Z(n11989) );
  XOR U13556 ( .A(n11903), .B(n11907), .Z(n11990) );
  XOR U13557 ( .A(n11898), .B(n11902), .Z(n11991) );
  XOR U13558 ( .A(n11893), .B(n11897), .Z(n11992) );
  XOR U13559 ( .A(n11888), .B(n11892), .Z(n11993) );
  XOR U13560 ( .A(n11883), .B(n11887), .Z(n11994) );
  XOR U13561 ( .A(n11878), .B(n11882), .Z(n11995) );
  XOR U13562 ( .A(n11873), .B(n11877), .Z(n11996) );
  XOR U13563 ( .A(n11868), .B(n11872), .Z(n11997) );
  XOR U13564 ( .A(n11863), .B(n11867), .Z(n11998) );
  XOR U13565 ( .A(n11858), .B(n11862), .Z(n11999) );
  XOR U13566 ( .A(n11848), .B(n11857), .Z(n12000) );
  XOR U13567 ( .A(n12001), .B(n11847), .Z(n11848) );
  AND U13568 ( .A(b[25]), .B(a[37]), .Z(n12001) );
  XNOR U13569 ( .A(n11847), .B(n11853), .Z(n12002) );
  XNOR U13570 ( .A(n11852), .B(n11844), .Z(n12003) );
  XOR U13571 ( .A(n11843), .B(n11840), .Z(n12004) );
  XOR U13572 ( .A(n12005), .B(n12006), .Z(n11840) );
  XOR U13573 ( .A(n11838), .B(n12007), .Z(n12006) );
  XOR U13574 ( .A(n12008), .B(n12009), .Z(n12007) );
  XOR U13575 ( .A(n12010), .B(n12011), .Z(n12009) );
  NAND U13576 ( .A(a[32]), .B(b[30]), .Z(n12011) );
  AND U13577 ( .A(a[31]), .B(b[31]), .Z(n12010) );
  XOR U13578 ( .A(n12012), .B(n12008), .Z(n12005) );
  XOR U13579 ( .A(n12013), .B(n12014), .Z(n12008) );
  ANDN U13580 ( .B(n12015), .A(n12016), .Z(n12013) );
  AND U13581 ( .A(a[33]), .B(b[29]), .Z(n12012) );
  XOR U13582 ( .A(n12017), .B(n11838), .Z(n11839) );
  XOR U13583 ( .A(n12018), .B(n12019), .Z(n11838) );
  AND U13584 ( .A(n12020), .B(n12021), .Z(n12018) );
  AND U13585 ( .A(a[34]), .B(b[28]), .Z(n12017) );
  XOR U13586 ( .A(n12022), .B(n11843), .Z(n11845) );
  XOR U13587 ( .A(n12023), .B(n12024), .Z(n11843) );
  AND U13588 ( .A(n12025), .B(n12026), .Z(n12023) );
  AND U13589 ( .A(a[35]), .B(b[27]), .Z(n12022) );
  XOR U13590 ( .A(n12027), .B(n12028), .Z(n11847) );
  AND U13591 ( .A(n12029), .B(n12030), .Z(n12027) );
  XOR U13592 ( .A(n12031), .B(n11852), .Z(n11854) );
  XOR U13593 ( .A(n12032), .B(n12033), .Z(n11852) );
  AND U13594 ( .A(n12034), .B(n12035), .Z(n12032) );
  AND U13595 ( .A(a[36]), .B(b[26]), .Z(n12031) );
  XOR U13596 ( .A(n12037), .B(n12038), .Z(n11857) );
  AND U13597 ( .A(n12039), .B(n12040), .Z(n12037) );
  AND U13598 ( .A(a[38]), .B(b[24]), .Z(n12036) );
  XOR U13599 ( .A(n12042), .B(n12043), .Z(n11862) );
  AND U13600 ( .A(n12044), .B(n12045), .Z(n12042) );
  AND U13601 ( .A(a[39]), .B(b[23]), .Z(n12041) );
  XOR U13602 ( .A(n12047), .B(n12048), .Z(n11867) );
  AND U13603 ( .A(n12049), .B(n12050), .Z(n12047) );
  AND U13604 ( .A(a[40]), .B(b[22]), .Z(n12046) );
  XOR U13605 ( .A(n12052), .B(n12053), .Z(n11872) );
  AND U13606 ( .A(n12054), .B(n12055), .Z(n12052) );
  AND U13607 ( .A(a[41]), .B(b[21]), .Z(n12051) );
  XOR U13608 ( .A(n12057), .B(n12058), .Z(n11877) );
  AND U13609 ( .A(n12059), .B(n12060), .Z(n12057) );
  AND U13610 ( .A(a[42]), .B(b[20]), .Z(n12056) );
  XOR U13611 ( .A(n12062), .B(n12063), .Z(n11882) );
  AND U13612 ( .A(n12064), .B(n12065), .Z(n12062) );
  AND U13613 ( .A(a[43]), .B(b[19]), .Z(n12061) );
  XOR U13614 ( .A(n12067), .B(n12068), .Z(n11887) );
  AND U13615 ( .A(n12069), .B(n12070), .Z(n12067) );
  AND U13616 ( .A(a[44]), .B(b[18]), .Z(n12066) );
  XOR U13617 ( .A(n12072), .B(n12073), .Z(n11892) );
  AND U13618 ( .A(n12074), .B(n12075), .Z(n12072) );
  AND U13619 ( .A(a[45]), .B(b[17]), .Z(n12071) );
  XOR U13620 ( .A(n12077), .B(n12078), .Z(n11897) );
  AND U13621 ( .A(n12079), .B(n12080), .Z(n12077) );
  AND U13622 ( .A(a[46]), .B(b[16]), .Z(n12076) );
  XOR U13623 ( .A(n12082), .B(n12083), .Z(n11902) );
  AND U13624 ( .A(n12084), .B(n12085), .Z(n12082) );
  AND U13625 ( .A(a[47]), .B(b[15]), .Z(n12081) );
  XOR U13626 ( .A(n12087), .B(n12088), .Z(n11907) );
  AND U13627 ( .A(n12089), .B(n12090), .Z(n12087) );
  AND U13628 ( .A(a[48]), .B(b[14]), .Z(n12086) );
  XOR U13629 ( .A(n12092), .B(n12093), .Z(n11912) );
  AND U13630 ( .A(n12094), .B(n12095), .Z(n12092) );
  AND U13631 ( .A(a[49]), .B(b[13]), .Z(n12091) );
  XOR U13632 ( .A(n12097), .B(n12098), .Z(n11917) );
  AND U13633 ( .A(n12099), .B(n12100), .Z(n12097) );
  AND U13634 ( .A(a[50]), .B(b[12]), .Z(n12096) );
  XOR U13635 ( .A(n12102), .B(n12103), .Z(n11922) );
  AND U13636 ( .A(n12104), .B(n12105), .Z(n12102) );
  AND U13637 ( .A(a[51]), .B(b[11]), .Z(n12101) );
  XOR U13638 ( .A(n12107), .B(n12108), .Z(n11927) );
  AND U13639 ( .A(n12109), .B(n12110), .Z(n12107) );
  AND U13640 ( .A(a[52]), .B(b[10]), .Z(n12106) );
  XOR U13641 ( .A(n12112), .B(n12113), .Z(n11932) );
  AND U13642 ( .A(n12114), .B(n12115), .Z(n12112) );
  AND U13643 ( .A(a[53]), .B(b[9]), .Z(n12111) );
  XOR U13644 ( .A(n12117), .B(n12118), .Z(n11937) );
  AND U13645 ( .A(n12119), .B(n12120), .Z(n12117) );
  AND U13646 ( .A(a[54]), .B(b[8]), .Z(n12116) );
  XOR U13647 ( .A(n12122), .B(n12123), .Z(n11942) );
  AND U13648 ( .A(n12124), .B(n12125), .Z(n12122) );
  AND U13649 ( .A(a[55]), .B(b[7]), .Z(n12121) );
  XOR U13650 ( .A(n12127), .B(n12128), .Z(n11947) );
  AND U13651 ( .A(n12129), .B(n12130), .Z(n12127) );
  AND U13652 ( .A(a[56]), .B(b[6]), .Z(n12126) );
  XOR U13653 ( .A(n12132), .B(n12133), .Z(n11952) );
  AND U13654 ( .A(n12134), .B(n12135), .Z(n12132) );
  AND U13655 ( .A(a[57]), .B(b[5]), .Z(n12131) );
  XOR U13656 ( .A(n12137), .B(n12138), .Z(n11957) );
  AND U13657 ( .A(n12139), .B(n12140), .Z(n12137) );
  AND U13658 ( .A(a[58]), .B(b[4]), .Z(n12136) );
  XOR U13659 ( .A(n12142), .B(n12143), .Z(n11962) );
  AND U13660 ( .A(n11976), .B(n11974), .Z(n12142) );
  AND U13661 ( .A(b[2]), .B(a[59]), .Z(n12144) );
  XOR U13662 ( .A(n12139), .B(n12143), .Z(n12145) );
  XOR U13663 ( .A(n12146), .B(n12147), .Z(n12143) );
  NANDN U13664 ( .A(n11978), .B(n11977), .Z(n12147) );
  XOR U13665 ( .A(n12148), .B(n12149), .Z(n11977) );
  NAND U13666 ( .A(a[59]), .B(b[1]), .Z(n12149) );
  XOR U13667 ( .A(n12150), .B(n12151), .Z(n11978) );
  XOR U13668 ( .A(n12148), .B(n12152), .Z(n12151) );
  IV U13669 ( .A(n12146), .Z(n12148) );
  ANDN U13670 ( .B(n5257), .A(n5259), .Z(n12146) );
  NAND U13671 ( .A(a[59]), .B(b[0]), .Z(n5259) );
  XNOR U13672 ( .A(n12153), .B(n12154), .Z(n5257) );
  XOR U13673 ( .A(n12134), .B(n12138), .Z(n12155) );
  XOR U13674 ( .A(n12129), .B(n12133), .Z(n12156) );
  XOR U13675 ( .A(n12124), .B(n12128), .Z(n12157) );
  XOR U13676 ( .A(n12119), .B(n12123), .Z(n12158) );
  XOR U13677 ( .A(n12114), .B(n12118), .Z(n12159) );
  XOR U13678 ( .A(n12109), .B(n12113), .Z(n12160) );
  XOR U13679 ( .A(n12104), .B(n12108), .Z(n12161) );
  XOR U13680 ( .A(n12099), .B(n12103), .Z(n12162) );
  XOR U13681 ( .A(n12094), .B(n12098), .Z(n12163) );
  XOR U13682 ( .A(n12089), .B(n12093), .Z(n12164) );
  XOR U13683 ( .A(n12084), .B(n12088), .Z(n12165) );
  XOR U13684 ( .A(n12079), .B(n12083), .Z(n12166) );
  XOR U13685 ( .A(n12074), .B(n12078), .Z(n12167) );
  XOR U13686 ( .A(n12069), .B(n12073), .Z(n12168) );
  XOR U13687 ( .A(n12064), .B(n12068), .Z(n12169) );
  XOR U13688 ( .A(n12059), .B(n12063), .Z(n12170) );
  XOR U13689 ( .A(n12054), .B(n12058), .Z(n12171) );
  XOR U13690 ( .A(n12049), .B(n12053), .Z(n12172) );
  XOR U13691 ( .A(n12044), .B(n12048), .Z(n12173) );
  XOR U13692 ( .A(n12039), .B(n12043), .Z(n12174) );
  XOR U13693 ( .A(n12029), .B(n12038), .Z(n12175) );
  XOR U13694 ( .A(n12176), .B(n12028), .Z(n12029) );
  AND U13695 ( .A(b[24]), .B(a[37]), .Z(n12176) );
  XNOR U13696 ( .A(n12028), .B(n12034), .Z(n12177) );
  XNOR U13697 ( .A(n12033), .B(n12025), .Z(n12178) );
  XNOR U13698 ( .A(n12024), .B(n12020), .Z(n12179) );
  XOR U13699 ( .A(n12019), .B(n12016), .Z(n12180) );
  XOR U13700 ( .A(n12181), .B(n12182), .Z(n12016) );
  XOR U13701 ( .A(n12014), .B(n12183), .Z(n12182) );
  XOR U13702 ( .A(n12184), .B(n12185), .Z(n12183) );
  XOR U13703 ( .A(n12186), .B(n12187), .Z(n12185) );
  NAND U13704 ( .A(a[31]), .B(b[30]), .Z(n12187) );
  AND U13705 ( .A(a[30]), .B(b[31]), .Z(n12186) );
  XOR U13706 ( .A(n12188), .B(n12184), .Z(n12181) );
  XOR U13707 ( .A(n12189), .B(n12190), .Z(n12184) );
  ANDN U13708 ( .B(n12191), .A(n12192), .Z(n12189) );
  AND U13709 ( .A(a[32]), .B(b[29]), .Z(n12188) );
  XOR U13710 ( .A(n12193), .B(n12014), .Z(n12015) );
  XOR U13711 ( .A(n12194), .B(n12195), .Z(n12014) );
  AND U13712 ( .A(n12196), .B(n12197), .Z(n12194) );
  AND U13713 ( .A(a[33]), .B(b[28]), .Z(n12193) );
  XOR U13714 ( .A(n12198), .B(n12019), .Z(n12021) );
  XOR U13715 ( .A(n12199), .B(n12200), .Z(n12019) );
  AND U13716 ( .A(n12201), .B(n12202), .Z(n12199) );
  AND U13717 ( .A(a[34]), .B(b[27]), .Z(n12198) );
  XOR U13718 ( .A(n12203), .B(n12024), .Z(n12026) );
  XOR U13719 ( .A(n12204), .B(n12205), .Z(n12024) );
  AND U13720 ( .A(n12206), .B(n12207), .Z(n12204) );
  AND U13721 ( .A(a[35]), .B(b[26]), .Z(n12203) );
  XOR U13722 ( .A(n12208), .B(n12209), .Z(n12028) );
  AND U13723 ( .A(n12210), .B(n12211), .Z(n12208) );
  XOR U13724 ( .A(n12212), .B(n12033), .Z(n12035) );
  XOR U13725 ( .A(n12213), .B(n12214), .Z(n12033) );
  AND U13726 ( .A(n12215), .B(n12216), .Z(n12213) );
  AND U13727 ( .A(a[36]), .B(b[25]), .Z(n12212) );
  XOR U13728 ( .A(n12218), .B(n12219), .Z(n12038) );
  AND U13729 ( .A(n12220), .B(n12221), .Z(n12218) );
  AND U13730 ( .A(a[38]), .B(b[23]), .Z(n12217) );
  XOR U13731 ( .A(n12223), .B(n12224), .Z(n12043) );
  AND U13732 ( .A(n12225), .B(n12226), .Z(n12223) );
  AND U13733 ( .A(a[39]), .B(b[22]), .Z(n12222) );
  XOR U13734 ( .A(n12228), .B(n12229), .Z(n12048) );
  AND U13735 ( .A(n12230), .B(n12231), .Z(n12228) );
  AND U13736 ( .A(a[40]), .B(b[21]), .Z(n12227) );
  XOR U13737 ( .A(n12233), .B(n12234), .Z(n12053) );
  AND U13738 ( .A(n12235), .B(n12236), .Z(n12233) );
  AND U13739 ( .A(a[41]), .B(b[20]), .Z(n12232) );
  XOR U13740 ( .A(n12238), .B(n12239), .Z(n12058) );
  AND U13741 ( .A(n12240), .B(n12241), .Z(n12238) );
  AND U13742 ( .A(a[42]), .B(b[19]), .Z(n12237) );
  XOR U13743 ( .A(n12243), .B(n12244), .Z(n12063) );
  AND U13744 ( .A(n12245), .B(n12246), .Z(n12243) );
  AND U13745 ( .A(a[43]), .B(b[18]), .Z(n12242) );
  XOR U13746 ( .A(n12248), .B(n12249), .Z(n12068) );
  AND U13747 ( .A(n12250), .B(n12251), .Z(n12248) );
  AND U13748 ( .A(a[44]), .B(b[17]), .Z(n12247) );
  XOR U13749 ( .A(n12253), .B(n12254), .Z(n12073) );
  AND U13750 ( .A(n12255), .B(n12256), .Z(n12253) );
  AND U13751 ( .A(a[45]), .B(b[16]), .Z(n12252) );
  XOR U13752 ( .A(n12258), .B(n12259), .Z(n12078) );
  AND U13753 ( .A(n12260), .B(n12261), .Z(n12258) );
  AND U13754 ( .A(a[46]), .B(b[15]), .Z(n12257) );
  XOR U13755 ( .A(n12263), .B(n12264), .Z(n12083) );
  AND U13756 ( .A(n12265), .B(n12266), .Z(n12263) );
  AND U13757 ( .A(a[47]), .B(b[14]), .Z(n12262) );
  XOR U13758 ( .A(n12268), .B(n12269), .Z(n12088) );
  AND U13759 ( .A(n12270), .B(n12271), .Z(n12268) );
  AND U13760 ( .A(a[48]), .B(b[13]), .Z(n12267) );
  XOR U13761 ( .A(n12273), .B(n12274), .Z(n12093) );
  AND U13762 ( .A(n12275), .B(n12276), .Z(n12273) );
  AND U13763 ( .A(a[49]), .B(b[12]), .Z(n12272) );
  XOR U13764 ( .A(n12278), .B(n12279), .Z(n12098) );
  AND U13765 ( .A(n12280), .B(n12281), .Z(n12278) );
  AND U13766 ( .A(a[50]), .B(b[11]), .Z(n12277) );
  XOR U13767 ( .A(n12283), .B(n12284), .Z(n12103) );
  AND U13768 ( .A(n12285), .B(n12286), .Z(n12283) );
  AND U13769 ( .A(a[51]), .B(b[10]), .Z(n12282) );
  XOR U13770 ( .A(n12288), .B(n12289), .Z(n12108) );
  AND U13771 ( .A(n12290), .B(n12291), .Z(n12288) );
  AND U13772 ( .A(a[52]), .B(b[9]), .Z(n12287) );
  XOR U13773 ( .A(n12293), .B(n12294), .Z(n12113) );
  AND U13774 ( .A(n12295), .B(n12296), .Z(n12293) );
  AND U13775 ( .A(a[53]), .B(b[8]), .Z(n12292) );
  XOR U13776 ( .A(n12298), .B(n12299), .Z(n12118) );
  AND U13777 ( .A(n12300), .B(n12301), .Z(n12298) );
  AND U13778 ( .A(a[54]), .B(b[7]), .Z(n12297) );
  XOR U13779 ( .A(n12303), .B(n12304), .Z(n12123) );
  AND U13780 ( .A(n12305), .B(n12306), .Z(n12303) );
  AND U13781 ( .A(a[55]), .B(b[6]), .Z(n12302) );
  XOR U13782 ( .A(n12308), .B(n12309), .Z(n12128) );
  AND U13783 ( .A(n12310), .B(n12311), .Z(n12308) );
  AND U13784 ( .A(a[56]), .B(b[5]), .Z(n12307) );
  XOR U13785 ( .A(n12313), .B(n12314), .Z(n12133) );
  AND U13786 ( .A(n12315), .B(n12316), .Z(n12313) );
  AND U13787 ( .A(a[57]), .B(b[4]), .Z(n12312) );
  XOR U13788 ( .A(n12318), .B(n12319), .Z(n12138) );
  AND U13789 ( .A(n12152), .B(n12150), .Z(n12318) );
  AND U13790 ( .A(b[2]), .B(a[58]), .Z(n12320) );
  XOR U13791 ( .A(n12315), .B(n12319), .Z(n12321) );
  XOR U13792 ( .A(n12322), .B(n12323), .Z(n12319) );
  NANDN U13793 ( .A(n12154), .B(n12153), .Z(n12323) );
  XOR U13794 ( .A(n12324), .B(n12325), .Z(n12153) );
  NAND U13795 ( .A(a[58]), .B(b[1]), .Z(n12325) );
  XOR U13796 ( .A(n12326), .B(n12327), .Z(n12154) );
  XOR U13797 ( .A(n12324), .B(n12328), .Z(n12327) );
  IV U13798 ( .A(n12322), .Z(n12324) );
  ANDN U13799 ( .B(n5262), .A(n5264), .Z(n12322) );
  NAND U13800 ( .A(a[58]), .B(b[0]), .Z(n5264) );
  XNOR U13801 ( .A(n12329), .B(n12330), .Z(n5262) );
  XOR U13802 ( .A(n12310), .B(n12314), .Z(n12331) );
  XOR U13803 ( .A(n12305), .B(n12309), .Z(n12332) );
  XOR U13804 ( .A(n12300), .B(n12304), .Z(n12333) );
  XOR U13805 ( .A(n12295), .B(n12299), .Z(n12334) );
  XOR U13806 ( .A(n12290), .B(n12294), .Z(n12335) );
  XOR U13807 ( .A(n12285), .B(n12289), .Z(n12336) );
  XOR U13808 ( .A(n12280), .B(n12284), .Z(n12337) );
  XOR U13809 ( .A(n12275), .B(n12279), .Z(n12338) );
  XOR U13810 ( .A(n12270), .B(n12274), .Z(n12339) );
  XOR U13811 ( .A(n12265), .B(n12269), .Z(n12340) );
  XOR U13812 ( .A(n12260), .B(n12264), .Z(n12341) );
  XOR U13813 ( .A(n12255), .B(n12259), .Z(n12342) );
  XOR U13814 ( .A(n12250), .B(n12254), .Z(n12343) );
  XOR U13815 ( .A(n12245), .B(n12249), .Z(n12344) );
  XOR U13816 ( .A(n12240), .B(n12244), .Z(n12345) );
  XOR U13817 ( .A(n12235), .B(n12239), .Z(n12346) );
  XOR U13818 ( .A(n12230), .B(n12234), .Z(n12347) );
  XOR U13819 ( .A(n12225), .B(n12229), .Z(n12348) );
  XOR U13820 ( .A(n12220), .B(n12224), .Z(n12349) );
  XOR U13821 ( .A(n12210), .B(n12219), .Z(n12350) );
  XOR U13822 ( .A(n12351), .B(n12209), .Z(n12210) );
  AND U13823 ( .A(b[23]), .B(a[37]), .Z(n12351) );
  XNOR U13824 ( .A(n12209), .B(n12215), .Z(n12352) );
  XNOR U13825 ( .A(n12214), .B(n12206), .Z(n12353) );
  XNOR U13826 ( .A(n12205), .B(n12201), .Z(n12354) );
  XNOR U13827 ( .A(n12200), .B(n12196), .Z(n12355) );
  XOR U13828 ( .A(n12195), .B(n12192), .Z(n12356) );
  XOR U13829 ( .A(n12357), .B(n12358), .Z(n12192) );
  XOR U13830 ( .A(n12190), .B(n12359), .Z(n12358) );
  XOR U13831 ( .A(n12360), .B(n12361), .Z(n12359) );
  XOR U13832 ( .A(n12362), .B(n12363), .Z(n12361) );
  NAND U13833 ( .A(b[30]), .B(a[30]), .Z(n12363) );
  AND U13834 ( .A(a[29]), .B(b[31]), .Z(n12362) );
  XOR U13835 ( .A(n12364), .B(n12360), .Z(n12357) );
  XOR U13836 ( .A(n12365), .B(n12366), .Z(n12360) );
  ANDN U13837 ( .B(n12367), .A(n12368), .Z(n12365) );
  AND U13838 ( .A(a[31]), .B(b[29]), .Z(n12364) );
  XOR U13839 ( .A(n12369), .B(n12190), .Z(n12191) );
  XOR U13840 ( .A(n12370), .B(n12371), .Z(n12190) );
  AND U13841 ( .A(n12372), .B(n12373), .Z(n12370) );
  AND U13842 ( .A(a[32]), .B(b[28]), .Z(n12369) );
  XOR U13843 ( .A(n12374), .B(n12195), .Z(n12197) );
  XOR U13844 ( .A(n12375), .B(n12376), .Z(n12195) );
  AND U13845 ( .A(n12377), .B(n12378), .Z(n12375) );
  AND U13846 ( .A(a[33]), .B(b[27]), .Z(n12374) );
  XOR U13847 ( .A(n12379), .B(n12200), .Z(n12202) );
  XOR U13848 ( .A(n12380), .B(n12381), .Z(n12200) );
  AND U13849 ( .A(n12382), .B(n12383), .Z(n12380) );
  AND U13850 ( .A(a[34]), .B(b[26]), .Z(n12379) );
  XOR U13851 ( .A(n12384), .B(n12205), .Z(n12207) );
  XOR U13852 ( .A(n12385), .B(n12386), .Z(n12205) );
  AND U13853 ( .A(n12387), .B(n12388), .Z(n12385) );
  AND U13854 ( .A(a[35]), .B(b[25]), .Z(n12384) );
  XOR U13855 ( .A(n12389), .B(n12390), .Z(n12209) );
  AND U13856 ( .A(n12391), .B(n12392), .Z(n12389) );
  XOR U13857 ( .A(n12393), .B(n12214), .Z(n12216) );
  XOR U13858 ( .A(n12394), .B(n12395), .Z(n12214) );
  AND U13859 ( .A(n12396), .B(n12397), .Z(n12394) );
  AND U13860 ( .A(a[36]), .B(b[24]), .Z(n12393) );
  XOR U13861 ( .A(n12399), .B(n12400), .Z(n12219) );
  AND U13862 ( .A(n12401), .B(n12402), .Z(n12399) );
  AND U13863 ( .A(a[38]), .B(b[22]), .Z(n12398) );
  XOR U13864 ( .A(n12404), .B(n12405), .Z(n12224) );
  AND U13865 ( .A(n12406), .B(n12407), .Z(n12404) );
  AND U13866 ( .A(a[39]), .B(b[21]), .Z(n12403) );
  XOR U13867 ( .A(n12409), .B(n12410), .Z(n12229) );
  AND U13868 ( .A(n12411), .B(n12412), .Z(n12409) );
  AND U13869 ( .A(a[40]), .B(b[20]), .Z(n12408) );
  XOR U13870 ( .A(n12414), .B(n12415), .Z(n12234) );
  AND U13871 ( .A(n12416), .B(n12417), .Z(n12414) );
  AND U13872 ( .A(a[41]), .B(b[19]), .Z(n12413) );
  XOR U13873 ( .A(n12419), .B(n12420), .Z(n12239) );
  AND U13874 ( .A(n12421), .B(n12422), .Z(n12419) );
  AND U13875 ( .A(a[42]), .B(b[18]), .Z(n12418) );
  XOR U13876 ( .A(n12424), .B(n12425), .Z(n12244) );
  AND U13877 ( .A(n12426), .B(n12427), .Z(n12424) );
  AND U13878 ( .A(a[43]), .B(b[17]), .Z(n12423) );
  XOR U13879 ( .A(n12429), .B(n12430), .Z(n12249) );
  AND U13880 ( .A(n12431), .B(n12432), .Z(n12429) );
  AND U13881 ( .A(a[44]), .B(b[16]), .Z(n12428) );
  XOR U13882 ( .A(n12434), .B(n12435), .Z(n12254) );
  AND U13883 ( .A(n12436), .B(n12437), .Z(n12434) );
  AND U13884 ( .A(a[45]), .B(b[15]), .Z(n12433) );
  XOR U13885 ( .A(n12439), .B(n12440), .Z(n12259) );
  AND U13886 ( .A(n12441), .B(n12442), .Z(n12439) );
  AND U13887 ( .A(a[46]), .B(b[14]), .Z(n12438) );
  XOR U13888 ( .A(n12444), .B(n12445), .Z(n12264) );
  AND U13889 ( .A(n12446), .B(n12447), .Z(n12444) );
  AND U13890 ( .A(a[47]), .B(b[13]), .Z(n12443) );
  XOR U13891 ( .A(n12449), .B(n12450), .Z(n12269) );
  AND U13892 ( .A(n12451), .B(n12452), .Z(n12449) );
  AND U13893 ( .A(a[48]), .B(b[12]), .Z(n12448) );
  XOR U13894 ( .A(n12454), .B(n12455), .Z(n12274) );
  AND U13895 ( .A(n12456), .B(n12457), .Z(n12454) );
  AND U13896 ( .A(a[49]), .B(b[11]), .Z(n12453) );
  XOR U13897 ( .A(n12459), .B(n12460), .Z(n12279) );
  AND U13898 ( .A(n12461), .B(n12462), .Z(n12459) );
  AND U13899 ( .A(a[50]), .B(b[10]), .Z(n12458) );
  XOR U13900 ( .A(n12464), .B(n12465), .Z(n12284) );
  AND U13901 ( .A(n12466), .B(n12467), .Z(n12464) );
  AND U13902 ( .A(a[51]), .B(b[9]), .Z(n12463) );
  XOR U13903 ( .A(n12469), .B(n12470), .Z(n12289) );
  AND U13904 ( .A(n12471), .B(n12472), .Z(n12469) );
  AND U13905 ( .A(a[52]), .B(b[8]), .Z(n12468) );
  XOR U13906 ( .A(n12474), .B(n12475), .Z(n12294) );
  AND U13907 ( .A(n12476), .B(n12477), .Z(n12474) );
  AND U13908 ( .A(a[53]), .B(b[7]), .Z(n12473) );
  XOR U13909 ( .A(n12479), .B(n12480), .Z(n12299) );
  AND U13910 ( .A(n12481), .B(n12482), .Z(n12479) );
  AND U13911 ( .A(a[54]), .B(b[6]), .Z(n12478) );
  XOR U13912 ( .A(n12484), .B(n12485), .Z(n12304) );
  AND U13913 ( .A(n12486), .B(n12487), .Z(n12484) );
  AND U13914 ( .A(a[55]), .B(b[5]), .Z(n12483) );
  XOR U13915 ( .A(n12489), .B(n12490), .Z(n12309) );
  AND U13916 ( .A(n12491), .B(n12492), .Z(n12489) );
  AND U13917 ( .A(a[56]), .B(b[4]), .Z(n12488) );
  XOR U13918 ( .A(n12494), .B(n12495), .Z(n12314) );
  AND U13919 ( .A(n12328), .B(n12326), .Z(n12494) );
  AND U13920 ( .A(b[2]), .B(a[57]), .Z(n12496) );
  XOR U13921 ( .A(n12491), .B(n12495), .Z(n12497) );
  XOR U13922 ( .A(n12498), .B(n12499), .Z(n12495) );
  NANDN U13923 ( .A(n12330), .B(n12329), .Z(n12499) );
  XOR U13924 ( .A(n12500), .B(n12501), .Z(n12329) );
  NAND U13925 ( .A(a[57]), .B(b[1]), .Z(n12501) );
  XOR U13926 ( .A(n12502), .B(n12503), .Z(n12330) );
  XOR U13927 ( .A(n12500), .B(n12504), .Z(n12503) );
  IV U13928 ( .A(n12498), .Z(n12500) );
  ANDN U13929 ( .B(n5267), .A(n5269), .Z(n12498) );
  NAND U13930 ( .A(a[57]), .B(b[0]), .Z(n5269) );
  XNOR U13931 ( .A(n12505), .B(n12506), .Z(n5267) );
  XOR U13932 ( .A(n12486), .B(n12490), .Z(n12507) );
  XOR U13933 ( .A(n12481), .B(n12485), .Z(n12508) );
  XOR U13934 ( .A(n12476), .B(n12480), .Z(n12509) );
  XOR U13935 ( .A(n12471), .B(n12475), .Z(n12510) );
  XOR U13936 ( .A(n12466), .B(n12470), .Z(n12511) );
  XOR U13937 ( .A(n12461), .B(n12465), .Z(n12512) );
  XOR U13938 ( .A(n12456), .B(n12460), .Z(n12513) );
  XOR U13939 ( .A(n12451), .B(n12455), .Z(n12514) );
  XOR U13940 ( .A(n12446), .B(n12450), .Z(n12515) );
  XOR U13941 ( .A(n12441), .B(n12445), .Z(n12516) );
  XOR U13942 ( .A(n12436), .B(n12440), .Z(n12517) );
  XOR U13943 ( .A(n12431), .B(n12435), .Z(n12518) );
  XOR U13944 ( .A(n12426), .B(n12430), .Z(n12519) );
  XOR U13945 ( .A(n12421), .B(n12425), .Z(n12520) );
  XOR U13946 ( .A(n12416), .B(n12420), .Z(n12521) );
  XOR U13947 ( .A(n12411), .B(n12415), .Z(n12522) );
  XOR U13948 ( .A(n12406), .B(n12410), .Z(n12523) );
  XOR U13949 ( .A(n12401), .B(n12405), .Z(n12524) );
  XOR U13950 ( .A(n12391), .B(n12400), .Z(n12525) );
  XOR U13951 ( .A(n12526), .B(n12390), .Z(n12391) );
  AND U13952 ( .A(b[22]), .B(a[37]), .Z(n12526) );
  XNOR U13953 ( .A(n12390), .B(n12396), .Z(n12527) );
  XNOR U13954 ( .A(n12395), .B(n12387), .Z(n12528) );
  XNOR U13955 ( .A(n12386), .B(n12382), .Z(n12529) );
  XNOR U13956 ( .A(n12381), .B(n12377), .Z(n12530) );
  XNOR U13957 ( .A(n12376), .B(n12372), .Z(n12531) );
  XOR U13958 ( .A(n12371), .B(n12368), .Z(n12532) );
  XOR U13959 ( .A(n12533), .B(n12534), .Z(n12368) );
  XOR U13960 ( .A(n12366), .B(n12535), .Z(n12534) );
  XOR U13961 ( .A(n12536), .B(n12537), .Z(n12535) );
  XOR U13962 ( .A(n12538), .B(n12539), .Z(n12537) );
  NAND U13963 ( .A(a[29]), .B(b[30]), .Z(n12539) );
  AND U13964 ( .A(a[28]), .B(b[31]), .Z(n12538) );
  XOR U13965 ( .A(n12540), .B(n12536), .Z(n12533) );
  XOR U13966 ( .A(n12541), .B(n12542), .Z(n12536) );
  ANDN U13967 ( .B(n12543), .A(n12544), .Z(n12541) );
  AND U13968 ( .A(b[29]), .B(a[30]), .Z(n12540) );
  XOR U13969 ( .A(n12545), .B(n12366), .Z(n12367) );
  XOR U13970 ( .A(n12546), .B(n12547), .Z(n12366) );
  AND U13971 ( .A(n12548), .B(n12549), .Z(n12546) );
  AND U13972 ( .A(a[31]), .B(b[28]), .Z(n12545) );
  XOR U13973 ( .A(n12550), .B(n12371), .Z(n12373) );
  XOR U13974 ( .A(n12551), .B(n12552), .Z(n12371) );
  AND U13975 ( .A(n12553), .B(n12554), .Z(n12551) );
  AND U13976 ( .A(a[32]), .B(b[27]), .Z(n12550) );
  XOR U13977 ( .A(n12555), .B(n12376), .Z(n12378) );
  XOR U13978 ( .A(n12556), .B(n12557), .Z(n12376) );
  AND U13979 ( .A(n12558), .B(n12559), .Z(n12556) );
  AND U13980 ( .A(a[33]), .B(b[26]), .Z(n12555) );
  XOR U13981 ( .A(n12560), .B(n12381), .Z(n12383) );
  XOR U13982 ( .A(n12561), .B(n12562), .Z(n12381) );
  AND U13983 ( .A(n12563), .B(n12564), .Z(n12561) );
  AND U13984 ( .A(a[34]), .B(b[25]), .Z(n12560) );
  XOR U13985 ( .A(n12565), .B(n12386), .Z(n12388) );
  XOR U13986 ( .A(n12566), .B(n12567), .Z(n12386) );
  AND U13987 ( .A(n12568), .B(n12569), .Z(n12566) );
  AND U13988 ( .A(a[35]), .B(b[24]), .Z(n12565) );
  XOR U13989 ( .A(n12570), .B(n12571), .Z(n12390) );
  AND U13990 ( .A(n12572), .B(n12573), .Z(n12570) );
  XOR U13991 ( .A(n12574), .B(n12395), .Z(n12397) );
  XOR U13992 ( .A(n12575), .B(n12576), .Z(n12395) );
  AND U13993 ( .A(n12577), .B(n12578), .Z(n12575) );
  AND U13994 ( .A(a[36]), .B(b[23]), .Z(n12574) );
  XOR U13995 ( .A(n12580), .B(n12581), .Z(n12400) );
  AND U13996 ( .A(n12582), .B(n12583), .Z(n12580) );
  AND U13997 ( .A(a[38]), .B(b[21]), .Z(n12579) );
  XOR U13998 ( .A(n12585), .B(n12586), .Z(n12405) );
  AND U13999 ( .A(n12587), .B(n12588), .Z(n12585) );
  AND U14000 ( .A(a[39]), .B(b[20]), .Z(n12584) );
  XOR U14001 ( .A(n12590), .B(n12591), .Z(n12410) );
  AND U14002 ( .A(n12592), .B(n12593), .Z(n12590) );
  AND U14003 ( .A(a[40]), .B(b[19]), .Z(n12589) );
  XOR U14004 ( .A(n12595), .B(n12596), .Z(n12415) );
  AND U14005 ( .A(n12597), .B(n12598), .Z(n12595) );
  AND U14006 ( .A(a[41]), .B(b[18]), .Z(n12594) );
  XOR U14007 ( .A(n12600), .B(n12601), .Z(n12420) );
  AND U14008 ( .A(n12602), .B(n12603), .Z(n12600) );
  AND U14009 ( .A(a[42]), .B(b[17]), .Z(n12599) );
  XOR U14010 ( .A(n12605), .B(n12606), .Z(n12425) );
  AND U14011 ( .A(n12607), .B(n12608), .Z(n12605) );
  AND U14012 ( .A(a[43]), .B(b[16]), .Z(n12604) );
  XOR U14013 ( .A(n12610), .B(n12611), .Z(n12430) );
  AND U14014 ( .A(n12612), .B(n12613), .Z(n12610) );
  AND U14015 ( .A(a[44]), .B(b[15]), .Z(n12609) );
  XOR U14016 ( .A(n12615), .B(n12616), .Z(n12435) );
  AND U14017 ( .A(n12617), .B(n12618), .Z(n12615) );
  AND U14018 ( .A(a[45]), .B(b[14]), .Z(n12614) );
  XOR U14019 ( .A(n12620), .B(n12621), .Z(n12440) );
  AND U14020 ( .A(n12622), .B(n12623), .Z(n12620) );
  AND U14021 ( .A(a[46]), .B(b[13]), .Z(n12619) );
  XOR U14022 ( .A(n12625), .B(n12626), .Z(n12445) );
  AND U14023 ( .A(n12627), .B(n12628), .Z(n12625) );
  AND U14024 ( .A(a[47]), .B(b[12]), .Z(n12624) );
  XOR U14025 ( .A(n12630), .B(n12631), .Z(n12450) );
  AND U14026 ( .A(n12632), .B(n12633), .Z(n12630) );
  AND U14027 ( .A(a[48]), .B(b[11]), .Z(n12629) );
  XOR U14028 ( .A(n12635), .B(n12636), .Z(n12455) );
  AND U14029 ( .A(n12637), .B(n12638), .Z(n12635) );
  AND U14030 ( .A(a[49]), .B(b[10]), .Z(n12634) );
  XOR U14031 ( .A(n12640), .B(n12641), .Z(n12460) );
  AND U14032 ( .A(n12642), .B(n12643), .Z(n12640) );
  AND U14033 ( .A(a[50]), .B(b[9]), .Z(n12639) );
  XOR U14034 ( .A(n12645), .B(n12646), .Z(n12465) );
  AND U14035 ( .A(n12647), .B(n12648), .Z(n12645) );
  AND U14036 ( .A(a[51]), .B(b[8]), .Z(n12644) );
  XOR U14037 ( .A(n12650), .B(n12651), .Z(n12470) );
  AND U14038 ( .A(n12652), .B(n12653), .Z(n12650) );
  AND U14039 ( .A(a[52]), .B(b[7]), .Z(n12649) );
  XOR U14040 ( .A(n12655), .B(n12656), .Z(n12475) );
  AND U14041 ( .A(n12657), .B(n12658), .Z(n12655) );
  AND U14042 ( .A(a[53]), .B(b[6]), .Z(n12654) );
  XOR U14043 ( .A(n12660), .B(n12661), .Z(n12480) );
  AND U14044 ( .A(n12662), .B(n12663), .Z(n12660) );
  AND U14045 ( .A(a[54]), .B(b[5]), .Z(n12659) );
  XOR U14046 ( .A(n12665), .B(n12666), .Z(n12485) );
  AND U14047 ( .A(n12667), .B(n12668), .Z(n12665) );
  AND U14048 ( .A(a[55]), .B(b[4]), .Z(n12664) );
  XOR U14049 ( .A(n12670), .B(n12671), .Z(n12490) );
  AND U14050 ( .A(n12504), .B(n12502), .Z(n12670) );
  AND U14051 ( .A(b[2]), .B(a[56]), .Z(n12672) );
  XOR U14052 ( .A(n12667), .B(n12671), .Z(n12673) );
  XOR U14053 ( .A(n12674), .B(n12675), .Z(n12671) );
  NANDN U14054 ( .A(n12506), .B(n12505), .Z(n12675) );
  XOR U14055 ( .A(n12676), .B(n12677), .Z(n12505) );
  NAND U14056 ( .A(a[56]), .B(b[1]), .Z(n12677) );
  XOR U14057 ( .A(n12678), .B(n12679), .Z(n12506) );
  XOR U14058 ( .A(n12676), .B(n12680), .Z(n12679) );
  IV U14059 ( .A(n12674), .Z(n12676) );
  ANDN U14060 ( .B(n5272), .A(n5274), .Z(n12674) );
  NAND U14061 ( .A(a[56]), .B(b[0]), .Z(n5274) );
  XNOR U14062 ( .A(n12681), .B(n12682), .Z(n5272) );
  XOR U14063 ( .A(n12662), .B(n12666), .Z(n12683) );
  XOR U14064 ( .A(n12657), .B(n12661), .Z(n12684) );
  XOR U14065 ( .A(n12652), .B(n12656), .Z(n12685) );
  XOR U14066 ( .A(n12647), .B(n12651), .Z(n12686) );
  XOR U14067 ( .A(n12642), .B(n12646), .Z(n12687) );
  XOR U14068 ( .A(n12637), .B(n12641), .Z(n12688) );
  XOR U14069 ( .A(n12632), .B(n12636), .Z(n12689) );
  XOR U14070 ( .A(n12627), .B(n12631), .Z(n12690) );
  XOR U14071 ( .A(n12622), .B(n12626), .Z(n12691) );
  XOR U14072 ( .A(n12617), .B(n12621), .Z(n12692) );
  XOR U14073 ( .A(n12612), .B(n12616), .Z(n12693) );
  XOR U14074 ( .A(n12607), .B(n12611), .Z(n12694) );
  XOR U14075 ( .A(n12602), .B(n12606), .Z(n12695) );
  XOR U14076 ( .A(n12597), .B(n12601), .Z(n12696) );
  XOR U14077 ( .A(n12592), .B(n12596), .Z(n12697) );
  XOR U14078 ( .A(n12587), .B(n12591), .Z(n12698) );
  XOR U14079 ( .A(n12582), .B(n12586), .Z(n12699) );
  XOR U14080 ( .A(n12572), .B(n12581), .Z(n12700) );
  XOR U14081 ( .A(n12701), .B(n12571), .Z(n12572) );
  AND U14082 ( .A(b[21]), .B(a[37]), .Z(n12701) );
  XNOR U14083 ( .A(n12571), .B(n12577), .Z(n12702) );
  XNOR U14084 ( .A(n12576), .B(n12568), .Z(n12703) );
  XNOR U14085 ( .A(n12567), .B(n12563), .Z(n12704) );
  XNOR U14086 ( .A(n12562), .B(n12558), .Z(n12705) );
  XNOR U14087 ( .A(n12557), .B(n12553), .Z(n12706) );
  XNOR U14088 ( .A(n12552), .B(n12548), .Z(n12707) );
  XOR U14089 ( .A(n12547), .B(n12544), .Z(n12708) );
  XOR U14090 ( .A(n12709), .B(n12710), .Z(n12544) );
  XOR U14091 ( .A(n12542), .B(n12711), .Z(n12710) );
  XOR U14092 ( .A(n12712), .B(n12713), .Z(n12711) );
  XOR U14093 ( .A(n12714), .B(n12715), .Z(n12713) );
  NAND U14094 ( .A(a[28]), .B(b[30]), .Z(n12715) );
  AND U14095 ( .A(a[27]), .B(b[31]), .Z(n12714) );
  XOR U14096 ( .A(n12716), .B(n12712), .Z(n12709) );
  XOR U14097 ( .A(n12717), .B(n12718), .Z(n12712) );
  ANDN U14098 ( .B(n12719), .A(n12720), .Z(n12717) );
  AND U14099 ( .A(a[29]), .B(b[29]), .Z(n12716) );
  XOR U14100 ( .A(n12721), .B(n12542), .Z(n12543) );
  XOR U14101 ( .A(n12722), .B(n12723), .Z(n12542) );
  AND U14102 ( .A(n12724), .B(n12725), .Z(n12722) );
  AND U14103 ( .A(b[28]), .B(a[30]), .Z(n12721) );
  XOR U14104 ( .A(n12726), .B(n12547), .Z(n12549) );
  XOR U14105 ( .A(n12727), .B(n12728), .Z(n12547) );
  AND U14106 ( .A(n12729), .B(n12730), .Z(n12727) );
  AND U14107 ( .A(a[31]), .B(b[27]), .Z(n12726) );
  XOR U14108 ( .A(n12731), .B(n12552), .Z(n12554) );
  XOR U14109 ( .A(n12732), .B(n12733), .Z(n12552) );
  AND U14110 ( .A(n12734), .B(n12735), .Z(n12732) );
  AND U14111 ( .A(a[32]), .B(b[26]), .Z(n12731) );
  XOR U14112 ( .A(n12736), .B(n12557), .Z(n12559) );
  XOR U14113 ( .A(n12737), .B(n12738), .Z(n12557) );
  AND U14114 ( .A(n12739), .B(n12740), .Z(n12737) );
  AND U14115 ( .A(a[33]), .B(b[25]), .Z(n12736) );
  XOR U14116 ( .A(n12741), .B(n12562), .Z(n12564) );
  XOR U14117 ( .A(n12742), .B(n12743), .Z(n12562) );
  AND U14118 ( .A(n12744), .B(n12745), .Z(n12742) );
  AND U14119 ( .A(a[34]), .B(b[24]), .Z(n12741) );
  XOR U14120 ( .A(n12746), .B(n12567), .Z(n12569) );
  XOR U14121 ( .A(n12747), .B(n12748), .Z(n12567) );
  AND U14122 ( .A(n12749), .B(n12750), .Z(n12747) );
  AND U14123 ( .A(a[35]), .B(b[23]), .Z(n12746) );
  XOR U14124 ( .A(n12751), .B(n12752), .Z(n12571) );
  AND U14125 ( .A(n12753), .B(n12754), .Z(n12751) );
  XOR U14126 ( .A(n12755), .B(n12576), .Z(n12578) );
  XOR U14127 ( .A(n12756), .B(n12757), .Z(n12576) );
  AND U14128 ( .A(n12758), .B(n12759), .Z(n12756) );
  AND U14129 ( .A(a[36]), .B(b[22]), .Z(n12755) );
  XOR U14130 ( .A(n12761), .B(n12762), .Z(n12581) );
  AND U14131 ( .A(n12763), .B(n12764), .Z(n12761) );
  AND U14132 ( .A(a[38]), .B(b[20]), .Z(n12760) );
  XOR U14133 ( .A(n12766), .B(n12767), .Z(n12586) );
  AND U14134 ( .A(n12768), .B(n12769), .Z(n12766) );
  AND U14135 ( .A(a[39]), .B(b[19]), .Z(n12765) );
  XOR U14136 ( .A(n12771), .B(n12772), .Z(n12591) );
  AND U14137 ( .A(n12773), .B(n12774), .Z(n12771) );
  AND U14138 ( .A(a[40]), .B(b[18]), .Z(n12770) );
  XOR U14139 ( .A(n12776), .B(n12777), .Z(n12596) );
  AND U14140 ( .A(n12778), .B(n12779), .Z(n12776) );
  AND U14141 ( .A(a[41]), .B(b[17]), .Z(n12775) );
  XOR U14142 ( .A(n12781), .B(n12782), .Z(n12601) );
  AND U14143 ( .A(n12783), .B(n12784), .Z(n12781) );
  AND U14144 ( .A(a[42]), .B(b[16]), .Z(n12780) );
  XOR U14145 ( .A(n12786), .B(n12787), .Z(n12606) );
  AND U14146 ( .A(n12788), .B(n12789), .Z(n12786) );
  AND U14147 ( .A(a[43]), .B(b[15]), .Z(n12785) );
  XOR U14148 ( .A(n12791), .B(n12792), .Z(n12611) );
  AND U14149 ( .A(n12793), .B(n12794), .Z(n12791) );
  AND U14150 ( .A(a[44]), .B(b[14]), .Z(n12790) );
  XOR U14151 ( .A(n12796), .B(n12797), .Z(n12616) );
  AND U14152 ( .A(n12798), .B(n12799), .Z(n12796) );
  AND U14153 ( .A(a[45]), .B(b[13]), .Z(n12795) );
  XOR U14154 ( .A(n12801), .B(n12802), .Z(n12621) );
  AND U14155 ( .A(n12803), .B(n12804), .Z(n12801) );
  AND U14156 ( .A(a[46]), .B(b[12]), .Z(n12800) );
  XOR U14157 ( .A(n12806), .B(n12807), .Z(n12626) );
  AND U14158 ( .A(n12808), .B(n12809), .Z(n12806) );
  AND U14159 ( .A(a[47]), .B(b[11]), .Z(n12805) );
  XOR U14160 ( .A(n12811), .B(n12812), .Z(n12631) );
  AND U14161 ( .A(n12813), .B(n12814), .Z(n12811) );
  AND U14162 ( .A(a[48]), .B(b[10]), .Z(n12810) );
  XOR U14163 ( .A(n12816), .B(n12817), .Z(n12636) );
  AND U14164 ( .A(n12818), .B(n12819), .Z(n12816) );
  AND U14165 ( .A(a[49]), .B(b[9]), .Z(n12815) );
  XOR U14166 ( .A(n12821), .B(n12822), .Z(n12641) );
  AND U14167 ( .A(n12823), .B(n12824), .Z(n12821) );
  AND U14168 ( .A(a[50]), .B(b[8]), .Z(n12820) );
  XOR U14169 ( .A(n12826), .B(n12827), .Z(n12646) );
  AND U14170 ( .A(n12828), .B(n12829), .Z(n12826) );
  AND U14171 ( .A(a[51]), .B(b[7]), .Z(n12825) );
  XOR U14172 ( .A(n12831), .B(n12832), .Z(n12651) );
  AND U14173 ( .A(n12833), .B(n12834), .Z(n12831) );
  AND U14174 ( .A(a[52]), .B(b[6]), .Z(n12830) );
  XOR U14175 ( .A(n12836), .B(n12837), .Z(n12656) );
  AND U14176 ( .A(n12838), .B(n12839), .Z(n12836) );
  AND U14177 ( .A(a[53]), .B(b[5]), .Z(n12835) );
  XOR U14178 ( .A(n12841), .B(n12842), .Z(n12661) );
  AND U14179 ( .A(n12843), .B(n12844), .Z(n12841) );
  AND U14180 ( .A(a[54]), .B(b[4]), .Z(n12840) );
  XOR U14181 ( .A(n12846), .B(n12847), .Z(n12666) );
  AND U14182 ( .A(n12680), .B(n12678), .Z(n12846) );
  AND U14183 ( .A(b[2]), .B(a[55]), .Z(n12848) );
  XOR U14184 ( .A(n12843), .B(n12847), .Z(n12849) );
  XOR U14185 ( .A(n12850), .B(n12851), .Z(n12847) );
  NANDN U14186 ( .A(n12682), .B(n12681), .Z(n12851) );
  XOR U14187 ( .A(n12852), .B(n12853), .Z(n12681) );
  NAND U14188 ( .A(a[55]), .B(b[1]), .Z(n12853) );
  XOR U14189 ( .A(n12854), .B(n12855), .Z(n12682) );
  XOR U14190 ( .A(n12852), .B(n12856), .Z(n12855) );
  IV U14191 ( .A(n12850), .Z(n12852) );
  ANDN U14192 ( .B(n5277), .A(n5279), .Z(n12850) );
  NAND U14193 ( .A(a[55]), .B(b[0]), .Z(n5279) );
  XNOR U14194 ( .A(n12857), .B(n12858), .Z(n5277) );
  XOR U14195 ( .A(n12838), .B(n12842), .Z(n12859) );
  XOR U14196 ( .A(n12833), .B(n12837), .Z(n12860) );
  XOR U14197 ( .A(n12828), .B(n12832), .Z(n12861) );
  XOR U14198 ( .A(n12823), .B(n12827), .Z(n12862) );
  XOR U14199 ( .A(n12818), .B(n12822), .Z(n12863) );
  XOR U14200 ( .A(n12813), .B(n12817), .Z(n12864) );
  XOR U14201 ( .A(n12808), .B(n12812), .Z(n12865) );
  XOR U14202 ( .A(n12803), .B(n12807), .Z(n12866) );
  XOR U14203 ( .A(n12798), .B(n12802), .Z(n12867) );
  XOR U14204 ( .A(n12793), .B(n12797), .Z(n12868) );
  XOR U14205 ( .A(n12788), .B(n12792), .Z(n12869) );
  XOR U14206 ( .A(n12783), .B(n12787), .Z(n12870) );
  XOR U14207 ( .A(n12778), .B(n12782), .Z(n12871) );
  XOR U14208 ( .A(n12773), .B(n12777), .Z(n12872) );
  XOR U14209 ( .A(n12768), .B(n12772), .Z(n12873) );
  XOR U14210 ( .A(n12763), .B(n12767), .Z(n12874) );
  XOR U14211 ( .A(n12753), .B(n12762), .Z(n12875) );
  XOR U14212 ( .A(n12876), .B(n12752), .Z(n12753) );
  AND U14213 ( .A(b[20]), .B(a[37]), .Z(n12876) );
  XNOR U14214 ( .A(n12752), .B(n12758), .Z(n12877) );
  XNOR U14215 ( .A(n12757), .B(n12749), .Z(n12878) );
  XNOR U14216 ( .A(n12748), .B(n12744), .Z(n12879) );
  XNOR U14217 ( .A(n12743), .B(n12739), .Z(n12880) );
  XNOR U14218 ( .A(n12738), .B(n12734), .Z(n12881) );
  XNOR U14219 ( .A(n12733), .B(n12729), .Z(n12882) );
  XNOR U14220 ( .A(n12728), .B(n12724), .Z(n12883) );
  XOR U14221 ( .A(n12723), .B(n12720), .Z(n12884) );
  XOR U14222 ( .A(n12885), .B(n12886), .Z(n12720) );
  XOR U14223 ( .A(n12718), .B(n12887), .Z(n12886) );
  XOR U14224 ( .A(n12888), .B(n12889), .Z(n12887) );
  XOR U14225 ( .A(n12890), .B(n12891), .Z(n12889) );
  NAND U14226 ( .A(a[27]), .B(b[30]), .Z(n12891) );
  AND U14227 ( .A(a[26]), .B(b[31]), .Z(n12890) );
  XOR U14228 ( .A(n12892), .B(n12888), .Z(n12885) );
  XOR U14229 ( .A(n12893), .B(n12894), .Z(n12888) );
  ANDN U14230 ( .B(n12895), .A(n12896), .Z(n12893) );
  AND U14231 ( .A(a[28]), .B(b[29]), .Z(n12892) );
  XOR U14232 ( .A(n12897), .B(n12718), .Z(n12719) );
  XOR U14233 ( .A(n12898), .B(n12899), .Z(n12718) );
  AND U14234 ( .A(n12900), .B(n12901), .Z(n12898) );
  AND U14235 ( .A(a[29]), .B(b[28]), .Z(n12897) );
  XOR U14236 ( .A(n12902), .B(n12723), .Z(n12725) );
  XOR U14237 ( .A(n12903), .B(n12904), .Z(n12723) );
  AND U14238 ( .A(n12905), .B(n12906), .Z(n12903) );
  AND U14239 ( .A(b[27]), .B(a[30]), .Z(n12902) );
  XOR U14240 ( .A(n12907), .B(n12728), .Z(n12730) );
  XOR U14241 ( .A(n12908), .B(n12909), .Z(n12728) );
  AND U14242 ( .A(n12910), .B(n12911), .Z(n12908) );
  AND U14243 ( .A(a[31]), .B(b[26]), .Z(n12907) );
  XOR U14244 ( .A(n12912), .B(n12733), .Z(n12735) );
  XOR U14245 ( .A(n12913), .B(n12914), .Z(n12733) );
  AND U14246 ( .A(n12915), .B(n12916), .Z(n12913) );
  AND U14247 ( .A(a[32]), .B(b[25]), .Z(n12912) );
  XOR U14248 ( .A(n12917), .B(n12738), .Z(n12740) );
  XOR U14249 ( .A(n12918), .B(n12919), .Z(n12738) );
  AND U14250 ( .A(n12920), .B(n12921), .Z(n12918) );
  AND U14251 ( .A(a[33]), .B(b[24]), .Z(n12917) );
  XOR U14252 ( .A(n12922), .B(n12743), .Z(n12745) );
  XOR U14253 ( .A(n12923), .B(n12924), .Z(n12743) );
  AND U14254 ( .A(n12925), .B(n12926), .Z(n12923) );
  AND U14255 ( .A(a[34]), .B(b[23]), .Z(n12922) );
  XOR U14256 ( .A(n12927), .B(n12748), .Z(n12750) );
  XOR U14257 ( .A(n12928), .B(n12929), .Z(n12748) );
  AND U14258 ( .A(n12930), .B(n12931), .Z(n12928) );
  AND U14259 ( .A(a[35]), .B(b[22]), .Z(n12927) );
  XOR U14260 ( .A(n12932), .B(n12933), .Z(n12752) );
  AND U14261 ( .A(n12934), .B(n12935), .Z(n12932) );
  XOR U14262 ( .A(n12936), .B(n12757), .Z(n12759) );
  XOR U14263 ( .A(n12937), .B(n12938), .Z(n12757) );
  AND U14264 ( .A(n12939), .B(n12940), .Z(n12937) );
  AND U14265 ( .A(a[36]), .B(b[21]), .Z(n12936) );
  XOR U14266 ( .A(n12942), .B(n12943), .Z(n12762) );
  AND U14267 ( .A(n12944), .B(n12945), .Z(n12942) );
  AND U14268 ( .A(a[38]), .B(b[19]), .Z(n12941) );
  XOR U14269 ( .A(n12947), .B(n12948), .Z(n12767) );
  AND U14270 ( .A(n12949), .B(n12950), .Z(n12947) );
  AND U14271 ( .A(a[39]), .B(b[18]), .Z(n12946) );
  XOR U14272 ( .A(n12952), .B(n12953), .Z(n12772) );
  AND U14273 ( .A(n12954), .B(n12955), .Z(n12952) );
  AND U14274 ( .A(a[40]), .B(b[17]), .Z(n12951) );
  XOR U14275 ( .A(n12957), .B(n12958), .Z(n12777) );
  AND U14276 ( .A(n12959), .B(n12960), .Z(n12957) );
  AND U14277 ( .A(a[41]), .B(b[16]), .Z(n12956) );
  XOR U14278 ( .A(n12962), .B(n12963), .Z(n12782) );
  AND U14279 ( .A(n12964), .B(n12965), .Z(n12962) );
  AND U14280 ( .A(a[42]), .B(b[15]), .Z(n12961) );
  XOR U14281 ( .A(n12967), .B(n12968), .Z(n12787) );
  AND U14282 ( .A(n12969), .B(n12970), .Z(n12967) );
  AND U14283 ( .A(a[43]), .B(b[14]), .Z(n12966) );
  XOR U14284 ( .A(n12972), .B(n12973), .Z(n12792) );
  AND U14285 ( .A(n12974), .B(n12975), .Z(n12972) );
  AND U14286 ( .A(a[44]), .B(b[13]), .Z(n12971) );
  XOR U14287 ( .A(n12977), .B(n12978), .Z(n12797) );
  AND U14288 ( .A(n12979), .B(n12980), .Z(n12977) );
  AND U14289 ( .A(a[45]), .B(b[12]), .Z(n12976) );
  XOR U14290 ( .A(n12982), .B(n12983), .Z(n12802) );
  AND U14291 ( .A(n12984), .B(n12985), .Z(n12982) );
  AND U14292 ( .A(a[46]), .B(b[11]), .Z(n12981) );
  XOR U14293 ( .A(n12987), .B(n12988), .Z(n12807) );
  AND U14294 ( .A(n12989), .B(n12990), .Z(n12987) );
  AND U14295 ( .A(a[47]), .B(b[10]), .Z(n12986) );
  XOR U14296 ( .A(n12992), .B(n12993), .Z(n12812) );
  AND U14297 ( .A(n12994), .B(n12995), .Z(n12992) );
  AND U14298 ( .A(a[48]), .B(b[9]), .Z(n12991) );
  XOR U14299 ( .A(n12997), .B(n12998), .Z(n12817) );
  AND U14300 ( .A(n12999), .B(n13000), .Z(n12997) );
  AND U14301 ( .A(a[49]), .B(b[8]), .Z(n12996) );
  XOR U14302 ( .A(n13002), .B(n13003), .Z(n12822) );
  AND U14303 ( .A(n13004), .B(n13005), .Z(n13002) );
  AND U14304 ( .A(a[50]), .B(b[7]), .Z(n13001) );
  XOR U14305 ( .A(n13007), .B(n13008), .Z(n12827) );
  AND U14306 ( .A(n13009), .B(n13010), .Z(n13007) );
  AND U14307 ( .A(a[51]), .B(b[6]), .Z(n13006) );
  XOR U14308 ( .A(n13012), .B(n13013), .Z(n12832) );
  AND U14309 ( .A(n13014), .B(n13015), .Z(n13012) );
  AND U14310 ( .A(a[52]), .B(b[5]), .Z(n13011) );
  XOR U14311 ( .A(n13017), .B(n13018), .Z(n12837) );
  AND U14312 ( .A(n13019), .B(n13020), .Z(n13017) );
  AND U14313 ( .A(a[53]), .B(b[4]), .Z(n13016) );
  XOR U14314 ( .A(n13022), .B(n13023), .Z(n12842) );
  AND U14315 ( .A(n12856), .B(n12854), .Z(n13022) );
  AND U14316 ( .A(b[2]), .B(a[54]), .Z(n13024) );
  XOR U14317 ( .A(n13019), .B(n13023), .Z(n13025) );
  XOR U14318 ( .A(n13026), .B(n13027), .Z(n13023) );
  NANDN U14319 ( .A(n12858), .B(n12857), .Z(n13027) );
  XOR U14320 ( .A(n13028), .B(n13029), .Z(n12857) );
  NAND U14321 ( .A(a[54]), .B(b[1]), .Z(n13029) );
  XOR U14322 ( .A(n13030), .B(n13031), .Z(n12858) );
  XOR U14323 ( .A(n13028), .B(n13032), .Z(n13031) );
  IV U14324 ( .A(n13026), .Z(n13028) );
  ANDN U14325 ( .B(n5282), .A(n5284), .Z(n13026) );
  NAND U14326 ( .A(a[54]), .B(b[0]), .Z(n5284) );
  XNOR U14327 ( .A(n13033), .B(n13034), .Z(n5282) );
  XOR U14328 ( .A(n13014), .B(n13018), .Z(n13035) );
  XOR U14329 ( .A(n13009), .B(n13013), .Z(n13036) );
  XOR U14330 ( .A(n13004), .B(n13008), .Z(n13037) );
  XOR U14331 ( .A(n12999), .B(n13003), .Z(n13038) );
  XOR U14332 ( .A(n12994), .B(n12998), .Z(n13039) );
  XOR U14333 ( .A(n12989), .B(n12993), .Z(n13040) );
  XOR U14334 ( .A(n12984), .B(n12988), .Z(n13041) );
  XOR U14335 ( .A(n12979), .B(n12983), .Z(n13042) );
  XOR U14336 ( .A(n12974), .B(n12978), .Z(n13043) );
  XOR U14337 ( .A(n12969), .B(n12973), .Z(n13044) );
  XOR U14338 ( .A(n12964), .B(n12968), .Z(n13045) );
  XOR U14339 ( .A(n12959), .B(n12963), .Z(n13046) );
  XOR U14340 ( .A(n12954), .B(n12958), .Z(n13047) );
  XOR U14341 ( .A(n12949), .B(n12953), .Z(n13048) );
  XOR U14342 ( .A(n12944), .B(n12948), .Z(n13049) );
  XOR U14343 ( .A(n12934), .B(n12943), .Z(n13050) );
  XOR U14344 ( .A(n13051), .B(n12933), .Z(n12934) );
  AND U14345 ( .A(b[19]), .B(a[37]), .Z(n13051) );
  XNOR U14346 ( .A(n12933), .B(n12939), .Z(n13052) );
  XNOR U14347 ( .A(n12938), .B(n12930), .Z(n13053) );
  XNOR U14348 ( .A(n12929), .B(n12925), .Z(n13054) );
  XNOR U14349 ( .A(n12924), .B(n12920), .Z(n13055) );
  XNOR U14350 ( .A(n12919), .B(n12915), .Z(n13056) );
  XNOR U14351 ( .A(n12914), .B(n12910), .Z(n13057) );
  XNOR U14352 ( .A(n12909), .B(n12905), .Z(n13058) );
  XNOR U14353 ( .A(n12904), .B(n12900), .Z(n13059) );
  XOR U14354 ( .A(n12899), .B(n12896), .Z(n13060) );
  XOR U14355 ( .A(n13061), .B(n13062), .Z(n12896) );
  XOR U14356 ( .A(n12894), .B(n13063), .Z(n13062) );
  XOR U14357 ( .A(n13064), .B(n13065), .Z(n13063) );
  XOR U14358 ( .A(n13066), .B(n13067), .Z(n13065) );
  NAND U14359 ( .A(a[26]), .B(b[30]), .Z(n13067) );
  AND U14360 ( .A(a[25]), .B(b[31]), .Z(n13066) );
  XOR U14361 ( .A(n13068), .B(n13064), .Z(n13061) );
  XOR U14362 ( .A(n13069), .B(n13070), .Z(n13064) );
  ANDN U14363 ( .B(n13071), .A(n13072), .Z(n13069) );
  AND U14364 ( .A(a[27]), .B(b[29]), .Z(n13068) );
  XOR U14365 ( .A(n13073), .B(n12894), .Z(n12895) );
  XOR U14366 ( .A(n13074), .B(n13075), .Z(n12894) );
  AND U14367 ( .A(n13076), .B(n13077), .Z(n13074) );
  AND U14368 ( .A(b[28]), .B(a[28]), .Z(n13073) );
  XOR U14369 ( .A(n13078), .B(n12899), .Z(n12901) );
  XOR U14370 ( .A(n13079), .B(n13080), .Z(n12899) );
  AND U14371 ( .A(n13081), .B(n13082), .Z(n13079) );
  AND U14372 ( .A(a[29]), .B(b[27]), .Z(n13078) );
  XOR U14373 ( .A(n13083), .B(n12904), .Z(n12906) );
  XOR U14374 ( .A(n13084), .B(n13085), .Z(n12904) );
  AND U14375 ( .A(n13086), .B(n13087), .Z(n13084) );
  AND U14376 ( .A(b[26]), .B(a[30]), .Z(n13083) );
  XOR U14377 ( .A(n13088), .B(n12909), .Z(n12911) );
  XOR U14378 ( .A(n13089), .B(n13090), .Z(n12909) );
  AND U14379 ( .A(n13091), .B(n13092), .Z(n13089) );
  AND U14380 ( .A(a[31]), .B(b[25]), .Z(n13088) );
  XOR U14381 ( .A(n13093), .B(n12914), .Z(n12916) );
  XOR U14382 ( .A(n13094), .B(n13095), .Z(n12914) );
  AND U14383 ( .A(n13096), .B(n13097), .Z(n13094) );
  AND U14384 ( .A(a[32]), .B(b[24]), .Z(n13093) );
  XOR U14385 ( .A(n13098), .B(n12919), .Z(n12921) );
  XOR U14386 ( .A(n13099), .B(n13100), .Z(n12919) );
  AND U14387 ( .A(n13101), .B(n13102), .Z(n13099) );
  AND U14388 ( .A(a[33]), .B(b[23]), .Z(n13098) );
  XOR U14389 ( .A(n13103), .B(n12924), .Z(n12926) );
  XOR U14390 ( .A(n13104), .B(n13105), .Z(n12924) );
  AND U14391 ( .A(n13106), .B(n13107), .Z(n13104) );
  AND U14392 ( .A(a[34]), .B(b[22]), .Z(n13103) );
  XOR U14393 ( .A(n13108), .B(n12929), .Z(n12931) );
  XOR U14394 ( .A(n13109), .B(n13110), .Z(n12929) );
  AND U14395 ( .A(n13111), .B(n13112), .Z(n13109) );
  AND U14396 ( .A(a[35]), .B(b[21]), .Z(n13108) );
  XOR U14397 ( .A(n13113), .B(n13114), .Z(n12933) );
  AND U14398 ( .A(n13115), .B(n13116), .Z(n13113) );
  XOR U14399 ( .A(n13117), .B(n12938), .Z(n12940) );
  XOR U14400 ( .A(n13118), .B(n13119), .Z(n12938) );
  AND U14401 ( .A(n13120), .B(n13121), .Z(n13118) );
  AND U14402 ( .A(a[36]), .B(b[20]), .Z(n13117) );
  XOR U14403 ( .A(n13123), .B(n13124), .Z(n12943) );
  AND U14404 ( .A(n13125), .B(n13126), .Z(n13123) );
  AND U14405 ( .A(a[38]), .B(b[18]), .Z(n13122) );
  XOR U14406 ( .A(n13128), .B(n13129), .Z(n12948) );
  AND U14407 ( .A(n13130), .B(n13131), .Z(n13128) );
  AND U14408 ( .A(a[39]), .B(b[17]), .Z(n13127) );
  XOR U14409 ( .A(n13133), .B(n13134), .Z(n12953) );
  AND U14410 ( .A(n13135), .B(n13136), .Z(n13133) );
  AND U14411 ( .A(a[40]), .B(b[16]), .Z(n13132) );
  XOR U14412 ( .A(n13138), .B(n13139), .Z(n12958) );
  AND U14413 ( .A(n13140), .B(n13141), .Z(n13138) );
  AND U14414 ( .A(a[41]), .B(b[15]), .Z(n13137) );
  XOR U14415 ( .A(n13143), .B(n13144), .Z(n12963) );
  AND U14416 ( .A(n13145), .B(n13146), .Z(n13143) );
  AND U14417 ( .A(a[42]), .B(b[14]), .Z(n13142) );
  XOR U14418 ( .A(n13148), .B(n13149), .Z(n12968) );
  AND U14419 ( .A(n13150), .B(n13151), .Z(n13148) );
  AND U14420 ( .A(a[43]), .B(b[13]), .Z(n13147) );
  XOR U14421 ( .A(n13153), .B(n13154), .Z(n12973) );
  AND U14422 ( .A(n13155), .B(n13156), .Z(n13153) );
  AND U14423 ( .A(a[44]), .B(b[12]), .Z(n13152) );
  XOR U14424 ( .A(n13158), .B(n13159), .Z(n12978) );
  AND U14425 ( .A(n13160), .B(n13161), .Z(n13158) );
  AND U14426 ( .A(a[45]), .B(b[11]), .Z(n13157) );
  XOR U14427 ( .A(n13163), .B(n13164), .Z(n12983) );
  AND U14428 ( .A(n13165), .B(n13166), .Z(n13163) );
  AND U14429 ( .A(a[46]), .B(b[10]), .Z(n13162) );
  XOR U14430 ( .A(n13168), .B(n13169), .Z(n12988) );
  AND U14431 ( .A(n13170), .B(n13171), .Z(n13168) );
  AND U14432 ( .A(a[47]), .B(b[9]), .Z(n13167) );
  XOR U14433 ( .A(n13173), .B(n13174), .Z(n12993) );
  AND U14434 ( .A(n13175), .B(n13176), .Z(n13173) );
  AND U14435 ( .A(a[48]), .B(b[8]), .Z(n13172) );
  XOR U14436 ( .A(n13178), .B(n13179), .Z(n12998) );
  AND U14437 ( .A(n13180), .B(n13181), .Z(n13178) );
  AND U14438 ( .A(a[49]), .B(b[7]), .Z(n13177) );
  XOR U14439 ( .A(n13183), .B(n13184), .Z(n13003) );
  AND U14440 ( .A(n13185), .B(n13186), .Z(n13183) );
  AND U14441 ( .A(a[50]), .B(b[6]), .Z(n13182) );
  XOR U14442 ( .A(n13188), .B(n13189), .Z(n13008) );
  AND U14443 ( .A(n13190), .B(n13191), .Z(n13188) );
  AND U14444 ( .A(a[51]), .B(b[5]), .Z(n13187) );
  XOR U14445 ( .A(n13193), .B(n13194), .Z(n13013) );
  AND U14446 ( .A(n13195), .B(n13196), .Z(n13193) );
  AND U14447 ( .A(a[52]), .B(b[4]), .Z(n13192) );
  XOR U14448 ( .A(n13198), .B(n13199), .Z(n13018) );
  AND U14449 ( .A(n13032), .B(n13030), .Z(n13198) );
  AND U14450 ( .A(b[2]), .B(a[53]), .Z(n13200) );
  XOR U14451 ( .A(n13195), .B(n13199), .Z(n13201) );
  XOR U14452 ( .A(n13202), .B(n13203), .Z(n13199) );
  NANDN U14453 ( .A(n13034), .B(n13033), .Z(n13203) );
  XOR U14454 ( .A(n13204), .B(n13205), .Z(n13033) );
  NAND U14455 ( .A(a[53]), .B(b[1]), .Z(n13205) );
  XOR U14456 ( .A(n13206), .B(n13207), .Z(n13034) );
  XOR U14457 ( .A(n13204), .B(n13208), .Z(n13207) );
  IV U14458 ( .A(n13202), .Z(n13204) );
  ANDN U14459 ( .B(n5287), .A(n5289), .Z(n13202) );
  NAND U14460 ( .A(a[53]), .B(b[0]), .Z(n5289) );
  XNOR U14461 ( .A(n13209), .B(n13210), .Z(n5287) );
  XOR U14462 ( .A(n13190), .B(n13194), .Z(n13211) );
  XOR U14463 ( .A(n13185), .B(n13189), .Z(n13212) );
  XOR U14464 ( .A(n13180), .B(n13184), .Z(n13213) );
  XOR U14465 ( .A(n13175), .B(n13179), .Z(n13214) );
  XOR U14466 ( .A(n13170), .B(n13174), .Z(n13215) );
  XOR U14467 ( .A(n13165), .B(n13169), .Z(n13216) );
  XOR U14468 ( .A(n13160), .B(n13164), .Z(n13217) );
  XOR U14469 ( .A(n13155), .B(n13159), .Z(n13218) );
  XOR U14470 ( .A(n13150), .B(n13154), .Z(n13219) );
  XOR U14471 ( .A(n13145), .B(n13149), .Z(n13220) );
  XOR U14472 ( .A(n13140), .B(n13144), .Z(n13221) );
  XOR U14473 ( .A(n13135), .B(n13139), .Z(n13222) );
  XOR U14474 ( .A(n13130), .B(n13134), .Z(n13223) );
  XOR U14475 ( .A(n13125), .B(n13129), .Z(n13224) );
  XOR U14476 ( .A(n13115), .B(n13124), .Z(n13225) );
  XOR U14477 ( .A(n13226), .B(n13114), .Z(n13115) );
  AND U14478 ( .A(b[18]), .B(a[37]), .Z(n13226) );
  XNOR U14479 ( .A(n13114), .B(n13120), .Z(n13227) );
  XNOR U14480 ( .A(n13119), .B(n13111), .Z(n13228) );
  XNOR U14481 ( .A(n13110), .B(n13106), .Z(n13229) );
  XNOR U14482 ( .A(n13105), .B(n13101), .Z(n13230) );
  XNOR U14483 ( .A(n13100), .B(n13096), .Z(n13231) );
  XNOR U14484 ( .A(n13095), .B(n13091), .Z(n13232) );
  XNOR U14485 ( .A(n13090), .B(n13086), .Z(n13233) );
  XNOR U14486 ( .A(n13085), .B(n13081), .Z(n13234) );
  XNOR U14487 ( .A(n13080), .B(n13076), .Z(n13235) );
  XOR U14488 ( .A(n13075), .B(n13072), .Z(n13236) );
  XOR U14489 ( .A(n13237), .B(n13238), .Z(n13072) );
  XOR U14490 ( .A(n13070), .B(n13239), .Z(n13238) );
  XOR U14491 ( .A(n13240), .B(n13241), .Z(n13239) );
  XOR U14492 ( .A(n13242), .B(n13243), .Z(n13241) );
  NAND U14493 ( .A(a[25]), .B(b[30]), .Z(n13243) );
  AND U14494 ( .A(a[24]), .B(b[31]), .Z(n13242) );
  XOR U14495 ( .A(n13244), .B(n13240), .Z(n13237) );
  XOR U14496 ( .A(n13245), .B(n13246), .Z(n13240) );
  ANDN U14497 ( .B(n13247), .A(n13248), .Z(n13245) );
  AND U14498 ( .A(a[26]), .B(b[29]), .Z(n13244) );
  XOR U14499 ( .A(n13249), .B(n13070), .Z(n13071) );
  XOR U14500 ( .A(n13250), .B(n13251), .Z(n13070) );
  AND U14501 ( .A(n13252), .B(n13253), .Z(n13250) );
  AND U14502 ( .A(a[27]), .B(b[28]), .Z(n13249) );
  XOR U14503 ( .A(n13254), .B(n13075), .Z(n13077) );
  XOR U14504 ( .A(n13255), .B(n13256), .Z(n13075) );
  AND U14505 ( .A(n13257), .B(n13258), .Z(n13255) );
  AND U14506 ( .A(b[27]), .B(a[28]), .Z(n13254) );
  XOR U14507 ( .A(n13259), .B(n13080), .Z(n13082) );
  XOR U14508 ( .A(n13260), .B(n13261), .Z(n13080) );
  AND U14509 ( .A(n13262), .B(n13263), .Z(n13260) );
  AND U14510 ( .A(a[29]), .B(b[26]), .Z(n13259) );
  XOR U14511 ( .A(n13264), .B(n13085), .Z(n13087) );
  XOR U14512 ( .A(n13265), .B(n13266), .Z(n13085) );
  AND U14513 ( .A(n13267), .B(n13268), .Z(n13265) );
  AND U14514 ( .A(b[25]), .B(a[30]), .Z(n13264) );
  XOR U14515 ( .A(n13269), .B(n13090), .Z(n13092) );
  XOR U14516 ( .A(n13270), .B(n13271), .Z(n13090) );
  AND U14517 ( .A(n13272), .B(n13273), .Z(n13270) );
  AND U14518 ( .A(a[31]), .B(b[24]), .Z(n13269) );
  XOR U14519 ( .A(n13274), .B(n13095), .Z(n13097) );
  XOR U14520 ( .A(n13275), .B(n13276), .Z(n13095) );
  AND U14521 ( .A(n13277), .B(n13278), .Z(n13275) );
  AND U14522 ( .A(a[32]), .B(b[23]), .Z(n13274) );
  XOR U14523 ( .A(n13279), .B(n13100), .Z(n13102) );
  XOR U14524 ( .A(n13280), .B(n13281), .Z(n13100) );
  AND U14525 ( .A(n13282), .B(n13283), .Z(n13280) );
  AND U14526 ( .A(a[33]), .B(b[22]), .Z(n13279) );
  XOR U14527 ( .A(n13284), .B(n13105), .Z(n13107) );
  XOR U14528 ( .A(n13285), .B(n13286), .Z(n13105) );
  AND U14529 ( .A(n13287), .B(n13288), .Z(n13285) );
  AND U14530 ( .A(a[34]), .B(b[21]), .Z(n13284) );
  XOR U14531 ( .A(n13289), .B(n13110), .Z(n13112) );
  XOR U14532 ( .A(n13290), .B(n13291), .Z(n13110) );
  AND U14533 ( .A(n13292), .B(n13293), .Z(n13290) );
  AND U14534 ( .A(a[35]), .B(b[20]), .Z(n13289) );
  XOR U14535 ( .A(n13294), .B(n13295), .Z(n13114) );
  AND U14536 ( .A(n13296), .B(n13297), .Z(n13294) );
  XOR U14537 ( .A(n13298), .B(n13119), .Z(n13121) );
  XOR U14538 ( .A(n13299), .B(n13300), .Z(n13119) );
  AND U14539 ( .A(n13301), .B(n13302), .Z(n13299) );
  AND U14540 ( .A(a[36]), .B(b[19]), .Z(n13298) );
  XOR U14541 ( .A(n13304), .B(n13305), .Z(n13124) );
  AND U14542 ( .A(n13306), .B(n13307), .Z(n13304) );
  AND U14543 ( .A(a[38]), .B(b[17]), .Z(n13303) );
  XOR U14544 ( .A(n13309), .B(n13310), .Z(n13129) );
  AND U14545 ( .A(n13311), .B(n13312), .Z(n13309) );
  AND U14546 ( .A(a[39]), .B(b[16]), .Z(n13308) );
  XOR U14547 ( .A(n13314), .B(n13315), .Z(n13134) );
  AND U14548 ( .A(n13316), .B(n13317), .Z(n13314) );
  AND U14549 ( .A(a[40]), .B(b[15]), .Z(n13313) );
  XOR U14550 ( .A(n13319), .B(n13320), .Z(n13139) );
  AND U14551 ( .A(n13321), .B(n13322), .Z(n13319) );
  AND U14552 ( .A(a[41]), .B(b[14]), .Z(n13318) );
  XOR U14553 ( .A(n13324), .B(n13325), .Z(n13144) );
  AND U14554 ( .A(n13326), .B(n13327), .Z(n13324) );
  AND U14555 ( .A(a[42]), .B(b[13]), .Z(n13323) );
  XOR U14556 ( .A(n13329), .B(n13330), .Z(n13149) );
  AND U14557 ( .A(n13331), .B(n13332), .Z(n13329) );
  AND U14558 ( .A(a[43]), .B(b[12]), .Z(n13328) );
  XOR U14559 ( .A(n13334), .B(n13335), .Z(n13154) );
  AND U14560 ( .A(n13336), .B(n13337), .Z(n13334) );
  AND U14561 ( .A(a[44]), .B(b[11]), .Z(n13333) );
  XOR U14562 ( .A(n13339), .B(n13340), .Z(n13159) );
  AND U14563 ( .A(n13341), .B(n13342), .Z(n13339) );
  AND U14564 ( .A(a[45]), .B(b[10]), .Z(n13338) );
  XOR U14565 ( .A(n13344), .B(n13345), .Z(n13164) );
  AND U14566 ( .A(n13346), .B(n13347), .Z(n13344) );
  AND U14567 ( .A(a[46]), .B(b[9]), .Z(n13343) );
  XOR U14568 ( .A(n13349), .B(n13350), .Z(n13169) );
  AND U14569 ( .A(n13351), .B(n13352), .Z(n13349) );
  AND U14570 ( .A(a[47]), .B(b[8]), .Z(n13348) );
  XOR U14571 ( .A(n13354), .B(n13355), .Z(n13174) );
  AND U14572 ( .A(n13356), .B(n13357), .Z(n13354) );
  AND U14573 ( .A(a[48]), .B(b[7]), .Z(n13353) );
  XOR U14574 ( .A(n13359), .B(n13360), .Z(n13179) );
  AND U14575 ( .A(n13361), .B(n13362), .Z(n13359) );
  AND U14576 ( .A(a[49]), .B(b[6]), .Z(n13358) );
  XOR U14577 ( .A(n13364), .B(n13365), .Z(n13184) );
  AND U14578 ( .A(n13366), .B(n13367), .Z(n13364) );
  AND U14579 ( .A(a[50]), .B(b[5]), .Z(n13363) );
  XOR U14580 ( .A(n13369), .B(n13370), .Z(n13189) );
  AND U14581 ( .A(n13371), .B(n13372), .Z(n13369) );
  AND U14582 ( .A(a[51]), .B(b[4]), .Z(n13368) );
  XOR U14583 ( .A(n13374), .B(n13375), .Z(n13194) );
  AND U14584 ( .A(n13208), .B(n13206), .Z(n13374) );
  AND U14585 ( .A(b[2]), .B(a[52]), .Z(n13376) );
  XOR U14586 ( .A(n13371), .B(n13375), .Z(n13377) );
  XOR U14587 ( .A(n13378), .B(n13379), .Z(n13375) );
  NANDN U14588 ( .A(n13210), .B(n13209), .Z(n13379) );
  XOR U14589 ( .A(n13380), .B(n13381), .Z(n13209) );
  NAND U14590 ( .A(a[52]), .B(b[1]), .Z(n13381) );
  XOR U14591 ( .A(n13382), .B(n13383), .Z(n13210) );
  XOR U14592 ( .A(n13380), .B(n13384), .Z(n13383) );
  IV U14593 ( .A(n13378), .Z(n13380) );
  ANDN U14594 ( .B(n5292), .A(n5294), .Z(n13378) );
  NAND U14595 ( .A(a[52]), .B(b[0]), .Z(n5294) );
  XNOR U14596 ( .A(n13385), .B(n13386), .Z(n5292) );
  XOR U14597 ( .A(n13366), .B(n13370), .Z(n13387) );
  XOR U14598 ( .A(n13361), .B(n13365), .Z(n13388) );
  XOR U14599 ( .A(n13356), .B(n13360), .Z(n13389) );
  XOR U14600 ( .A(n13351), .B(n13355), .Z(n13390) );
  XOR U14601 ( .A(n13346), .B(n13350), .Z(n13391) );
  XOR U14602 ( .A(n13341), .B(n13345), .Z(n13392) );
  XOR U14603 ( .A(n13336), .B(n13340), .Z(n13393) );
  XOR U14604 ( .A(n13331), .B(n13335), .Z(n13394) );
  XOR U14605 ( .A(n13326), .B(n13330), .Z(n13395) );
  XOR U14606 ( .A(n13321), .B(n13325), .Z(n13396) );
  XOR U14607 ( .A(n13316), .B(n13320), .Z(n13397) );
  XOR U14608 ( .A(n13311), .B(n13315), .Z(n13398) );
  XOR U14609 ( .A(n13306), .B(n13310), .Z(n13399) );
  XOR U14610 ( .A(n13296), .B(n13305), .Z(n13400) );
  XOR U14611 ( .A(n13401), .B(n13295), .Z(n13296) );
  AND U14612 ( .A(b[17]), .B(a[37]), .Z(n13401) );
  XNOR U14613 ( .A(n13295), .B(n13301), .Z(n13402) );
  XNOR U14614 ( .A(n13300), .B(n13292), .Z(n13403) );
  XNOR U14615 ( .A(n13291), .B(n13287), .Z(n13404) );
  XNOR U14616 ( .A(n13286), .B(n13282), .Z(n13405) );
  XNOR U14617 ( .A(n13281), .B(n13277), .Z(n13406) );
  XNOR U14618 ( .A(n13276), .B(n13272), .Z(n13407) );
  XNOR U14619 ( .A(n13271), .B(n13267), .Z(n13408) );
  XNOR U14620 ( .A(n13266), .B(n13262), .Z(n13409) );
  XNOR U14621 ( .A(n13261), .B(n13257), .Z(n13410) );
  XNOR U14622 ( .A(n13256), .B(n13252), .Z(n13411) );
  XOR U14623 ( .A(n13251), .B(n13248), .Z(n13412) );
  XOR U14624 ( .A(n13413), .B(n13414), .Z(n13248) );
  XOR U14625 ( .A(n13246), .B(n13415), .Z(n13414) );
  XOR U14626 ( .A(n13416), .B(n13417), .Z(n13415) );
  XOR U14627 ( .A(n13418), .B(n13419), .Z(n13417) );
  NAND U14628 ( .A(a[24]), .B(b[30]), .Z(n13419) );
  AND U14629 ( .A(a[23]), .B(b[31]), .Z(n13418) );
  XOR U14630 ( .A(n13420), .B(n13416), .Z(n13413) );
  XOR U14631 ( .A(n13421), .B(n13422), .Z(n13416) );
  ANDN U14632 ( .B(n13423), .A(n13424), .Z(n13421) );
  AND U14633 ( .A(a[25]), .B(b[29]), .Z(n13420) );
  XOR U14634 ( .A(n13425), .B(n13246), .Z(n13247) );
  XOR U14635 ( .A(n13426), .B(n13427), .Z(n13246) );
  AND U14636 ( .A(n13428), .B(n13429), .Z(n13426) );
  AND U14637 ( .A(a[26]), .B(b[28]), .Z(n13425) );
  XOR U14638 ( .A(n13430), .B(n13251), .Z(n13253) );
  XOR U14639 ( .A(n13431), .B(n13432), .Z(n13251) );
  AND U14640 ( .A(n13433), .B(n13434), .Z(n13431) );
  AND U14641 ( .A(a[27]), .B(b[27]), .Z(n13430) );
  XOR U14642 ( .A(n13435), .B(n13256), .Z(n13258) );
  XOR U14643 ( .A(n13436), .B(n13437), .Z(n13256) );
  AND U14644 ( .A(n13438), .B(n13439), .Z(n13436) );
  AND U14645 ( .A(b[26]), .B(a[28]), .Z(n13435) );
  XOR U14646 ( .A(n13440), .B(n13261), .Z(n13263) );
  XOR U14647 ( .A(n13441), .B(n13442), .Z(n13261) );
  AND U14648 ( .A(n13443), .B(n13444), .Z(n13441) );
  AND U14649 ( .A(a[29]), .B(b[25]), .Z(n13440) );
  XOR U14650 ( .A(n13445), .B(n13266), .Z(n13268) );
  XOR U14651 ( .A(n13446), .B(n13447), .Z(n13266) );
  AND U14652 ( .A(n13448), .B(n13449), .Z(n13446) );
  AND U14653 ( .A(b[24]), .B(a[30]), .Z(n13445) );
  XOR U14654 ( .A(n13450), .B(n13271), .Z(n13273) );
  XOR U14655 ( .A(n13451), .B(n13452), .Z(n13271) );
  AND U14656 ( .A(n13453), .B(n13454), .Z(n13451) );
  AND U14657 ( .A(a[31]), .B(b[23]), .Z(n13450) );
  XOR U14658 ( .A(n13455), .B(n13276), .Z(n13278) );
  XOR U14659 ( .A(n13456), .B(n13457), .Z(n13276) );
  AND U14660 ( .A(n13458), .B(n13459), .Z(n13456) );
  AND U14661 ( .A(a[32]), .B(b[22]), .Z(n13455) );
  XOR U14662 ( .A(n13460), .B(n13281), .Z(n13283) );
  XOR U14663 ( .A(n13461), .B(n13462), .Z(n13281) );
  AND U14664 ( .A(n13463), .B(n13464), .Z(n13461) );
  AND U14665 ( .A(a[33]), .B(b[21]), .Z(n13460) );
  XOR U14666 ( .A(n13465), .B(n13286), .Z(n13288) );
  XOR U14667 ( .A(n13466), .B(n13467), .Z(n13286) );
  AND U14668 ( .A(n13468), .B(n13469), .Z(n13466) );
  AND U14669 ( .A(a[34]), .B(b[20]), .Z(n13465) );
  XOR U14670 ( .A(n13470), .B(n13291), .Z(n13293) );
  XOR U14671 ( .A(n13471), .B(n13472), .Z(n13291) );
  AND U14672 ( .A(n13473), .B(n13474), .Z(n13471) );
  AND U14673 ( .A(a[35]), .B(b[19]), .Z(n13470) );
  XOR U14674 ( .A(n13475), .B(n13476), .Z(n13295) );
  AND U14675 ( .A(n13477), .B(n13478), .Z(n13475) );
  XOR U14676 ( .A(n13479), .B(n13300), .Z(n13302) );
  XOR U14677 ( .A(n13480), .B(n13481), .Z(n13300) );
  AND U14678 ( .A(n13482), .B(n13483), .Z(n13480) );
  AND U14679 ( .A(a[36]), .B(b[18]), .Z(n13479) );
  XOR U14680 ( .A(n13485), .B(n13486), .Z(n13305) );
  AND U14681 ( .A(n13487), .B(n13488), .Z(n13485) );
  AND U14682 ( .A(a[38]), .B(b[16]), .Z(n13484) );
  XOR U14683 ( .A(n13490), .B(n13491), .Z(n13310) );
  AND U14684 ( .A(n13492), .B(n13493), .Z(n13490) );
  AND U14685 ( .A(a[39]), .B(b[15]), .Z(n13489) );
  XOR U14686 ( .A(n13495), .B(n13496), .Z(n13315) );
  AND U14687 ( .A(n13497), .B(n13498), .Z(n13495) );
  AND U14688 ( .A(a[40]), .B(b[14]), .Z(n13494) );
  XOR U14689 ( .A(n13500), .B(n13501), .Z(n13320) );
  AND U14690 ( .A(n13502), .B(n13503), .Z(n13500) );
  AND U14691 ( .A(a[41]), .B(b[13]), .Z(n13499) );
  XOR U14692 ( .A(n13505), .B(n13506), .Z(n13325) );
  AND U14693 ( .A(n13507), .B(n13508), .Z(n13505) );
  AND U14694 ( .A(a[42]), .B(b[12]), .Z(n13504) );
  XOR U14695 ( .A(n13510), .B(n13511), .Z(n13330) );
  AND U14696 ( .A(n13512), .B(n13513), .Z(n13510) );
  AND U14697 ( .A(a[43]), .B(b[11]), .Z(n13509) );
  XOR U14698 ( .A(n13515), .B(n13516), .Z(n13335) );
  AND U14699 ( .A(n13517), .B(n13518), .Z(n13515) );
  AND U14700 ( .A(a[44]), .B(b[10]), .Z(n13514) );
  XOR U14701 ( .A(n13520), .B(n13521), .Z(n13340) );
  AND U14702 ( .A(n13522), .B(n13523), .Z(n13520) );
  AND U14703 ( .A(a[45]), .B(b[9]), .Z(n13519) );
  XOR U14704 ( .A(n13525), .B(n13526), .Z(n13345) );
  AND U14705 ( .A(n13527), .B(n13528), .Z(n13525) );
  AND U14706 ( .A(a[46]), .B(b[8]), .Z(n13524) );
  XOR U14707 ( .A(n13530), .B(n13531), .Z(n13350) );
  AND U14708 ( .A(n13532), .B(n13533), .Z(n13530) );
  AND U14709 ( .A(a[47]), .B(b[7]), .Z(n13529) );
  XOR U14710 ( .A(n13535), .B(n13536), .Z(n13355) );
  AND U14711 ( .A(n13537), .B(n13538), .Z(n13535) );
  AND U14712 ( .A(a[48]), .B(b[6]), .Z(n13534) );
  XOR U14713 ( .A(n13540), .B(n13541), .Z(n13360) );
  AND U14714 ( .A(n13542), .B(n13543), .Z(n13540) );
  AND U14715 ( .A(a[49]), .B(b[5]), .Z(n13539) );
  XOR U14716 ( .A(n13545), .B(n13546), .Z(n13365) );
  AND U14717 ( .A(n13547), .B(n13548), .Z(n13545) );
  AND U14718 ( .A(a[50]), .B(b[4]), .Z(n13544) );
  XOR U14719 ( .A(n13550), .B(n13551), .Z(n13370) );
  AND U14720 ( .A(n13384), .B(n13382), .Z(n13550) );
  AND U14721 ( .A(b[2]), .B(a[51]), .Z(n13552) );
  XOR U14722 ( .A(n13547), .B(n13551), .Z(n13553) );
  XOR U14723 ( .A(n13554), .B(n13555), .Z(n13551) );
  NANDN U14724 ( .A(n13386), .B(n13385), .Z(n13555) );
  XOR U14725 ( .A(n13556), .B(n13557), .Z(n13385) );
  NAND U14726 ( .A(a[51]), .B(b[1]), .Z(n13557) );
  XOR U14727 ( .A(n13558), .B(n13559), .Z(n13386) );
  XOR U14728 ( .A(n13556), .B(n13560), .Z(n13559) );
  IV U14729 ( .A(n13554), .Z(n13556) );
  ANDN U14730 ( .B(n5297), .A(n5299), .Z(n13554) );
  NAND U14731 ( .A(a[51]), .B(b[0]), .Z(n5299) );
  XNOR U14732 ( .A(n13561), .B(n13562), .Z(n5297) );
  XOR U14733 ( .A(n13542), .B(n13546), .Z(n13563) );
  XOR U14734 ( .A(n13537), .B(n13541), .Z(n13564) );
  XOR U14735 ( .A(n13532), .B(n13536), .Z(n13565) );
  XOR U14736 ( .A(n13527), .B(n13531), .Z(n13566) );
  XOR U14737 ( .A(n13522), .B(n13526), .Z(n13567) );
  XOR U14738 ( .A(n13517), .B(n13521), .Z(n13568) );
  XOR U14739 ( .A(n13512), .B(n13516), .Z(n13569) );
  XOR U14740 ( .A(n13507), .B(n13511), .Z(n13570) );
  XOR U14741 ( .A(n13502), .B(n13506), .Z(n13571) );
  XOR U14742 ( .A(n13497), .B(n13501), .Z(n13572) );
  XOR U14743 ( .A(n13492), .B(n13496), .Z(n13573) );
  XOR U14744 ( .A(n13487), .B(n13491), .Z(n13574) );
  XOR U14745 ( .A(n13477), .B(n13486), .Z(n13575) );
  XOR U14746 ( .A(n13576), .B(n13476), .Z(n13477) );
  AND U14747 ( .A(b[16]), .B(a[37]), .Z(n13576) );
  XNOR U14748 ( .A(n13476), .B(n13482), .Z(n13577) );
  XNOR U14749 ( .A(n13481), .B(n13473), .Z(n13578) );
  XNOR U14750 ( .A(n13472), .B(n13468), .Z(n13579) );
  XNOR U14751 ( .A(n13467), .B(n13463), .Z(n13580) );
  XNOR U14752 ( .A(n13462), .B(n13458), .Z(n13581) );
  XNOR U14753 ( .A(n13457), .B(n13453), .Z(n13582) );
  XNOR U14754 ( .A(n13452), .B(n13448), .Z(n13583) );
  XNOR U14755 ( .A(n13447), .B(n13443), .Z(n13584) );
  XNOR U14756 ( .A(n13442), .B(n13438), .Z(n13585) );
  XNOR U14757 ( .A(n13437), .B(n13433), .Z(n13586) );
  XNOR U14758 ( .A(n13432), .B(n13428), .Z(n13587) );
  XOR U14759 ( .A(n13427), .B(n13424), .Z(n13588) );
  XOR U14760 ( .A(n13589), .B(n13590), .Z(n13424) );
  XOR U14761 ( .A(n13422), .B(n13591), .Z(n13590) );
  XOR U14762 ( .A(n13592), .B(n13593), .Z(n13591) );
  XOR U14763 ( .A(n13594), .B(n13595), .Z(n13593) );
  NAND U14764 ( .A(a[23]), .B(b[30]), .Z(n13595) );
  AND U14765 ( .A(a[22]), .B(b[31]), .Z(n13594) );
  XOR U14766 ( .A(n13596), .B(n13592), .Z(n13589) );
  XOR U14767 ( .A(n13597), .B(n13598), .Z(n13592) );
  ANDN U14768 ( .B(n13599), .A(n13600), .Z(n13597) );
  AND U14769 ( .A(a[24]), .B(b[29]), .Z(n13596) );
  XOR U14770 ( .A(n13601), .B(n13422), .Z(n13423) );
  XOR U14771 ( .A(n13602), .B(n13603), .Z(n13422) );
  AND U14772 ( .A(n13604), .B(n13605), .Z(n13602) );
  AND U14773 ( .A(a[25]), .B(b[28]), .Z(n13601) );
  XOR U14774 ( .A(n13606), .B(n13427), .Z(n13429) );
  XOR U14775 ( .A(n13607), .B(n13608), .Z(n13427) );
  AND U14776 ( .A(n13609), .B(n13610), .Z(n13607) );
  AND U14777 ( .A(a[26]), .B(b[27]), .Z(n13606) );
  XOR U14778 ( .A(n13611), .B(n13432), .Z(n13434) );
  XOR U14779 ( .A(n13612), .B(n13613), .Z(n13432) );
  AND U14780 ( .A(n13614), .B(n13615), .Z(n13612) );
  AND U14781 ( .A(a[27]), .B(b[26]), .Z(n13611) );
  XOR U14782 ( .A(n13616), .B(n13437), .Z(n13439) );
  XOR U14783 ( .A(n13617), .B(n13618), .Z(n13437) );
  AND U14784 ( .A(n13619), .B(n13620), .Z(n13617) );
  AND U14785 ( .A(b[25]), .B(a[28]), .Z(n13616) );
  XOR U14786 ( .A(n13621), .B(n13442), .Z(n13444) );
  XOR U14787 ( .A(n13622), .B(n13623), .Z(n13442) );
  AND U14788 ( .A(n13624), .B(n13625), .Z(n13622) );
  AND U14789 ( .A(a[29]), .B(b[24]), .Z(n13621) );
  XOR U14790 ( .A(n13626), .B(n13447), .Z(n13449) );
  XOR U14791 ( .A(n13627), .B(n13628), .Z(n13447) );
  AND U14792 ( .A(n13629), .B(n13630), .Z(n13627) );
  AND U14793 ( .A(b[23]), .B(a[30]), .Z(n13626) );
  XOR U14794 ( .A(n13631), .B(n13452), .Z(n13454) );
  XOR U14795 ( .A(n13632), .B(n13633), .Z(n13452) );
  AND U14796 ( .A(n13634), .B(n13635), .Z(n13632) );
  AND U14797 ( .A(a[31]), .B(b[22]), .Z(n13631) );
  XOR U14798 ( .A(n13636), .B(n13457), .Z(n13459) );
  XOR U14799 ( .A(n13637), .B(n13638), .Z(n13457) );
  AND U14800 ( .A(n13639), .B(n13640), .Z(n13637) );
  AND U14801 ( .A(a[32]), .B(b[21]), .Z(n13636) );
  XOR U14802 ( .A(n13641), .B(n13462), .Z(n13464) );
  XOR U14803 ( .A(n13642), .B(n13643), .Z(n13462) );
  AND U14804 ( .A(n13644), .B(n13645), .Z(n13642) );
  AND U14805 ( .A(a[33]), .B(b[20]), .Z(n13641) );
  XOR U14806 ( .A(n13646), .B(n13467), .Z(n13469) );
  XOR U14807 ( .A(n13647), .B(n13648), .Z(n13467) );
  AND U14808 ( .A(n13649), .B(n13650), .Z(n13647) );
  AND U14809 ( .A(a[34]), .B(b[19]), .Z(n13646) );
  XOR U14810 ( .A(n13651), .B(n13472), .Z(n13474) );
  XOR U14811 ( .A(n13652), .B(n13653), .Z(n13472) );
  AND U14812 ( .A(n13654), .B(n13655), .Z(n13652) );
  AND U14813 ( .A(a[35]), .B(b[18]), .Z(n13651) );
  XOR U14814 ( .A(n13656), .B(n13657), .Z(n13476) );
  AND U14815 ( .A(n13658), .B(n13659), .Z(n13656) );
  XOR U14816 ( .A(n13660), .B(n13481), .Z(n13483) );
  XOR U14817 ( .A(n13661), .B(n13662), .Z(n13481) );
  AND U14818 ( .A(n13663), .B(n13664), .Z(n13661) );
  AND U14819 ( .A(a[36]), .B(b[17]), .Z(n13660) );
  XOR U14820 ( .A(n13666), .B(n13667), .Z(n13486) );
  AND U14821 ( .A(n13668), .B(n13669), .Z(n13666) );
  AND U14822 ( .A(a[38]), .B(b[15]), .Z(n13665) );
  XOR U14823 ( .A(n13671), .B(n13672), .Z(n13491) );
  AND U14824 ( .A(n13673), .B(n13674), .Z(n13671) );
  AND U14825 ( .A(a[39]), .B(b[14]), .Z(n13670) );
  XOR U14826 ( .A(n13676), .B(n13677), .Z(n13496) );
  AND U14827 ( .A(n13678), .B(n13679), .Z(n13676) );
  AND U14828 ( .A(a[40]), .B(b[13]), .Z(n13675) );
  XOR U14829 ( .A(n13681), .B(n13682), .Z(n13501) );
  AND U14830 ( .A(n13683), .B(n13684), .Z(n13681) );
  AND U14831 ( .A(a[41]), .B(b[12]), .Z(n13680) );
  XOR U14832 ( .A(n13686), .B(n13687), .Z(n13506) );
  AND U14833 ( .A(n13688), .B(n13689), .Z(n13686) );
  AND U14834 ( .A(a[42]), .B(b[11]), .Z(n13685) );
  XOR U14835 ( .A(n13691), .B(n13692), .Z(n13511) );
  AND U14836 ( .A(n13693), .B(n13694), .Z(n13691) );
  AND U14837 ( .A(a[43]), .B(b[10]), .Z(n13690) );
  XOR U14838 ( .A(n13696), .B(n13697), .Z(n13516) );
  AND U14839 ( .A(n13698), .B(n13699), .Z(n13696) );
  AND U14840 ( .A(a[44]), .B(b[9]), .Z(n13695) );
  XOR U14841 ( .A(n13701), .B(n13702), .Z(n13521) );
  AND U14842 ( .A(n13703), .B(n13704), .Z(n13701) );
  AND U14843 ( .A(a[45]), .B(b[8]), .Z(n13700) );
  XOR U14844 ( .A(n13706), .B(n13707), .Z(n13526) );
  AND U14845 ( .A(n13708), .B(n13709), .Z(n13706) );
  AND U14846 ( .A(a[46]), .B(b[7]), .Z(n13705) );
  XOR U14847 ( .A(n13711), .B(n13712), .Z(n13531) );
  AND U14848 ( .A(n13713), .B(n13714), .Z(n13711) );
  AND U14849 ( .A(a[47]), .B(b[6]), .Z(n13710) );
  XOR U14850 ( .A(n13716), .B(n13717), .Z(n13536) );
  AND U14851 ( .A(n13718), .B(n13719), .Z(n13716) );
  AND U14852 ( .A(a[48]), .B(b[5]), .Z(n13715) );
  XOR U14853 ( .A(n13721), .B(n13722), .Z(n13541) );
  AND U14854 ( .A(n13723), .B(n13724), .Z(n13721) );
  AND U14855 ( .A(a[49]), .B(b[4]), .Z(n13720) );
  XOR U14856 ( .A(n13726), .B(n13727), .Z(n13546) );
  AND U14857 ( .A(n13560), .B(n13558), .Z(n13726) );
  AND U14858 ( .A(b[2]), .B(a[50]), .Z(n13728) );
  XOR U14859 ( .A(n13723), .B(n13727), .Z(n13729) );
  XOR U14860 ( .A(n13730), .B(n13731), .Z(n13727) );
  NANDN U14861 ( .A(n13562), .B(n13561), .Z(n13731) );
  XOR U14862 ( .A(n13732), .B(n13733), .Z(n13561) );
  NAND U14863 ( .A(a[50]), .B(b[1]), .Z(n13733) );
  XOR U14864 ( .A(n13734), .B(n13735), .Z(n13562) );
  XOR U14865 ( .A(n13732), .B(n13736), .Z(n13735) );
  IV U14866 ( .A(n13730), .Z(n13732) );
  ANDN U14867 ( .B(n5302), .A(n5304), .Z(n13730) );
  NAND U14868 ( .A(a[50]), .B(b[0]), .Z(n5304) );
  XNOR U14869 ( .A(n13737), .B(n13738), .Z(n5302) );
  XOR U14870 ( .A(n13718), .B(n13722), .Z(n13739) );
  XOR U14871 ( .A(n13713), .B(n13717), .Z(n13740) );
  XOR U14872 ( .A(n13708), .B(n13712), .Z(n13741) );
  XOR U14873 ( .A(n13703), .B(n13707), .Z(n13742) );
  XOR U14874 ( .A(n13698), .B(n13702), .Z(n13743) );
  XOR U14875 ( .A(n13693), .B(n13697), .Z(n13744) );
  XOR U14876 ( .A(n13688), .B(n13692), .Z(n13745) );
  XOR U14877 ( .A(n13683), .B(n13687), .Z(n13746) );
  XOR U14878 ( .A(n13678), .B(n13682), .Z(n13747) );
  XOR U14879 ( .A(n13673), .B(n13677), .Z(n13748) );
  XOR U14880 ( .A(n13668), .B(n13672), .Z(n13749) );
  XOR U14881 ( .A(n13658), .B(n13667), .Z(n13750) );
  XOR U14882 ( .A(n13751), .B(n13657), .Z(n13658) );
  AND U14883 ( .A(b[15]), .B(a[37]), .Z(n13751) );
  XNOR U14884 ( .A(n13657), .B(n13663), .Z(n13752) );
  XNOR U14885 ( .A(n13662), .B(n13654), .Z(n13753) );
  XNOR U14886 ( .A(n13653), .B(n13649), .Z(n13754) );
  XNOR U14887 ( .A(n13648), .B(n13644), .Z(n13755) );
  XNOR U14888 ( .A(n13643), .B(n13639), .Z(n13756) );
  XNOR U14889 ( .A(n13638), .B(n13634), .Z(n13757) );
  XNOR U14890 ( .A(n13633), .B(n13629), .Z(n13758) );
  XNOR U14891 ( .A(n13628), .B(n13624), .Z(n13759) );
  XNOR U14892 ( .A(n13623), .B(n13619), .Z(n13760) );
  XNOR U14893 ( .A(n13618), .B(n13614), .Z(n13761) );
  XNOR U14894 ( .A(n13613), .B(n13609), .Z(n13762) );
  XNOR U14895 ( .A(n13608), .B(n13604), .Z(n13763) );
  XOR U14896 ( .A(n13603), .B(n13600), .Z(n13764) );
  XOR U14897 ( .A(n13765), .B(n13766), .Z(n13600) );
  XOR U14898 ( .A(n13598), .B(n13767), .Z(n13766) );
  XOR U14899 ( .A(n13768), .B(n13769), .Z(n13767) );
  XOR U14900 ( .A(n13770), .B(n13771), .Z(n13769) );
  NAND U14901 ( .A(a[22]), .B(b[30]), .Z(n13771) );
  AND U14902 ( .A(a[21]), .B(b[31]), .Z(n13770) );
  XOR U14903 ( .A(n13772), .B(n13768), .Z(n13765) );
  XOR U14904 ( .A(n13773), .B(n13774), .Z(n13768) );
  ANDN U14905 ( .B(n13775), .A(n13776), .Z(n13773) );
  AND U14906 ( .A(a[23]), .B(b[29]), .Z(n13772) );
  XOR U14907 ( .A(n13777), .B(n13598), .Z(n13599) );
  XOR U14908 ( .A(n13778), .B(n13779), .Z(n13598) );
  AND U14909 ( .A(n13780), .B(n13781), .Z(n13778) );
  AND U14910 ( .A(a[24]), .B(b[28]), .Z(n13777) );
  XOR U14911 ( .A(n13782), .B(n13603), .Z(n13605) );
  XOR U14912 ( .A(n13783), .B(n13784), .Z(n13603) );
  AND U14913 ( .A(n13785), .B(n13786), .Z(n13783) );
  AND U14914 ( .A(a[25]), .B(b[27]), .Z(n13782) );
  XOR U14915 ( .A(n13787), .B(n13608), .Z(n13610) );
  XOR U14916 ( .A(n13788), .B(n13789), .Z(n13608) );
  AND U14917 ( .A(n13790), .B(n13791), .Z(n13788) );
  AND U14918 ( .A(b[26]), .B(a[26]), .Z(n13787) );
  XOR U14919 ( .A(n13792), .B(n13613), .Z(n13615) );
  XOR U14920 ( .A(n13793), .B(n13794), .Z(n13613) );
  AND U14921 ( .A(n13795), .B(n13796), .Z(n13793) );
  AND U14922 ( .A(a[27]), .B(b[25]), .Z(n13792) );
  XOR U14923 ( .A(n13797), .B(n13618), .Z(n13620) );
  XOR U14924 ( .A(n13798), .B(n13799), .Z(n13618) );
  AND U14925 ( .A(n13800), .B(n13801), .Z(n13798) );
  AND U14926 ( .A(b[24]), .B(a[28]), .Z(n13797) );
  XOR U14927 ( .A(n13802), .B(n13623), .Z(n13625) );
  XOR U14928 ( .A(n13803), .B(n13804), .Z(n13623) );
  AND U14929 ( .A(n13805), .B(n13806), .Z(n13803) );
  AND U14930 ( .A(a[29]), .B(b[23]), .Z(n13802) );
  XOR U14931 ( .A(n13807), .B(n13628), .Z(n13630) );
  XOR U14932 ( .A(n13808), .B(n13809), .Z(n13628) );
  AND U14933 ( .A(n13810), .B(n13811), .Z(n13808) );
  AND U14934 ( .A(b[22]), .B(a[30]), .Z(n13807) );
  XOR U14935 ( .A(n13812), .B(n13633), .Z(n13635) );
  XOR U14936 ( .A(n13813), .B(n13814), .Z(n13633) );
  AND U14937 ( .A(n13815), .B(n13816), .Z(n13813) );
  AND U14938 ( .A(a[31]), .B(b[21]), .Z(n13812) );
  XOR U14939 ( .A(n13817), .B(n13638), .Z(n13640) );
  XOR U14940 ( .A(n13818), .B(n13819), .Z(n13638) );
  AND U14941 ( .A(n13820), .B(n13821), .Z(n13818) );
  AND U14942 ( .A(a[32]), .B(b[20]), .Z(n13817) );
  XOR U14943 ( .A(n13822), .B(n13643), .Z(n13645) );
  XOR U14944 ( .A(n13823), .B(n13824), .Z(n13643) );
  AND U14945 ( .A(n13825), .B(n13826), .Z(n13823) );
  AND U14946 ( .A(a[33]), .B(b[19]), .Z(n13822) );
  XOR U14947 ( .A(n13827), .B(n13648), .Z(n13650) );
  XOR U14948 ( .A(n13828), .B(n13829), .Z(n13648) );
  AND U14949 ( .A(n13830), .B(n13831), .Z(n13828) );
  AND U14950 ( .A(a[34]), .B(b[18]), .Z(n13827) );
  XOR U14951 ( .A(n13832), .B(n13653), .Z(n13655) );
  XOR U14952 ( .A(n13833), .B(n13834), .Z(n13653) );
  AND U14953 ( .A(n13835), .B(n13836), .Z(n13833) );
  AND U14954 ( .A(a[35]), .B(b[17]), .Z(n13832) );
  XOR U14955 ( .A(n13837), .B(n13838), .Z(n13657) );
  AND U14956 ( .A(n13839), .B(n13840), .Z(n13837) );
  XOR U14957 ( .A(n13841), .B(n13662), .Z(n13664) );
  XOR U14958 ( .A(n13842), .B(n13843), .Z(n13662) );
  AND U14959 ( .A(n13844), .B(n13845), .Z(n13842) );
  AND U14960 ( .A(a[36]), .B(b[16]), .Z(n13841) );
  XOR U14961 ( .A(n13847), .B(n13848), .Z(n13667) );
  AND U14962 ( .A(n13849), .B(n13850), .Z(n13847) );
  AND U14963 ( .A(a[38]), .B(b[14]), .Z(n13846) );
  XOR U14964 ( .A(n13852), .B(n13853), .Z(n13672) );
  AND U14965 ( .A(n13854), .B(n13855), .Z(n13852) );
  AND U14966 ( .A(a[39]), .B(b[13]), .Z(n13851) );
  XOR U14967 ( .A(n13857), .B(n13858), .Z(n13677) );
  AND U14968 ( .A(n13859), .B(n13860), .Z(n13857) );
  AND U14969 ( .A(a[40]), .B(b[12]), .Z(n13856) );
  XOR U14970 ( .A(n13862), .B(n13863), .Z(n13682) );
  AND U14971 ( .A(n13864), .B(n13865), .Z(n13862) );
  AND U14972 ( .A(a[41]), .B(b[11]), .Z(n13861) );
  XOR U14973 ( .A(n13867), .B(n13868), .Z(n13687) );
  AND U14974 ( .A(n13869), .B(n13870), .Z(n13867) );
  AND U14975 ( .A(a[42]), .B(b[10]), .Z(n13866) );
  XOR U14976 ( .A(n13872), .B(n13873), .Z(n13692) );
  AND U14977 ( .A(n13874), .B(n13875), .Z(n13872) );
  AND U14978 ( .A(a[43]), .B(b[9]), .Z(n13871) );
  XOR U14979 ( .A(n13877), .B(n13878), .Z(n13697) );
  AND U14980 ( .A(n13879), .B(n13880), .Z(n13877) );
  AND U14981 ( .A(a[44]), .B(b[8]), .Z(n13876) );
  XOR U14982 ( .A(n13882), .B(n13883), .Z(n13702) );
  AND U14983 ( .A(n13884), .B(n13885), .Z(n13882) );
  AND U14984 ( .A(a[45]), .B(b[7]), .Z(n13881) );
  XOR U14985 ( .A(n13887), .B(n13888), .Z(n13707) );
  AND U14986 ( .A(n13889), .B(n13890), .Z(n13887) );
  AND U14987 ( .A(a[46]), .B(b[6]), .Z(n13886) );
  XOR U14988 ( .A(n13892), .B(n13893), .Z(n13712) );
  AND U14989 ( .A(n13894), .B(n13895), .Z(n13892) );
  AND U14990 ( .A(a[47]), .B(b[5]), .Z(n13891) );
  XOR U14991 ( .A(n13897), .B(n13898), .Z(n13717) );
  AND U14992 ( .A(n13899), .B(n13900), .Z(n13897) );
  AND U14993 ( .A(a[48]), .B(b[4]), .Z(n13896) );
  XOR U14994 ( .A(n13902), .B(n13903), .Z(n13722) );
  AND U14995 ( .A(n13736), .B(n13734), .Z(n13902) );
  AND U14996 ( .A(b[2]), .B(a[49]), .Z(n13904) );
  XOR U14997 ( .A(n13899), .B(n13903), .Z(n13905) );
  XOR U14998 ( .A(n13906), .B(n13907), .Z(n13903) );
  NANDN U14999 ( .A(n13738), .B(n13737), .Z(n13907) );
  XOR U15000 ( .A(n13908), .B(n13909), .Z(n13737) );
  NAND U15001 ( .A(a[49]), .B(b[1]), .Z(n13909) );
  XOR U15002 ( .A(n13910), .B(n13911), .Z(n13738) );
  XOR U15003 ( .A(n13908), .B(n13912), .Z(n13911) );
  IV U15004 ( .A(n13906), .Z(n13908) );
  ANDN U15005 ( .B(n5307), .A(n5309), .Z(n13906) );
  NAND U15006 ( .A(a[49]), .B(b[0]), .Z(n5309) );
  XNOR U15007 ( .A(n13913), .B(n13914), .Z(n5307) );
  XOR U15008 ( .A(n13894), .B(n13898), .Z(n13915) );
  XOR U15009 ( .A(n13889), .B(n13893), .Z(n13916) );
  XOR U15010 ( .A(n13884), .B(n13888), .Z(n13917) );
  XOR U15011 ( .A(n13879), .B(n13883), .Z(n13918) );
  XOR U15012 ( .A(n13874), .B(n13878), .Z(n13919) );
  XOR U15013 ( .A(n13869), .B(n13873), .Z(n13920) );
  XOR U15014 ( .A(n13864), .B(n13868), .Z(n13921) );
  XOR U15015 ( .A(n13859), .B(n13863), .Z(n13922) );
  XOR U15016 ( .A(n13854), .B(n13858), .Z(n13923) );
  XOR U15017 ( .A(n13849), .B(n13853), .Z(n13924) );
  XOR U15018 ( .A(n13839), .B(n13848), .Z(n13925) );
  XOR U15019 ( .A(n13926), .B(n13838), .Z(n13839) );
  AND U15020 ( .A(b[14]), .B(a[37]), .Z(n13926) );
  XNOR U15021 ( .A(n13838), .B(n13844), .Z(n13927) );
  XNOR U15022 ( .A(n13843), .B(n13835), .Z(n13928) );
  XNOR U15023 ( .A(n13834), .B(n13830), .Z(n13929) );
  XNOR U15024 ( .A(n13829), .B(n13825), .Z(n13930) );
  XNOR U15025 ( .A(n13824), .B(n13820), .Z(n13931) );
  XNOR U15026 ( .A(n13819), .B(n13815), .Z(n13932) );
  XNOR U15027 ( .A(n13814), .B(n13810), .Z(n13933) );
  XNOR U15028 ( .A(n13809), .B(n13805), .Z(n13934) );
  XNOR U15029 ( .A(n13804), .B(n13800), .Z(n13935) );
  XNOR U15030 ( .A(n13799), .B(n13795), .Z(n13936) );
  XNOR U15031 ( .A(n13794), .B(n13790), .Z(n13937) );
  XNOR U15032 ( .A(n13789), .B(n13785), .Z(n13938) );
  XNOR U15033 ( .A(n13784), .B(n13780), .Z(n13939) );
  XOR U15034 ( .A(n13779), .B(n13776), .Z(n13940) );
  XOR U15035 ( .A(n13941), .B(n13942), .Z(n13776) );
  XOR U15036 ( .A(n13774), .B(n13943), .Z(n13942) );
  XOR U15037 ( .A(n13944), .B(n13945), .Z(n13943) );
  XOR U15038 ( .A(n13946), .B(n13947), .Z(n13945) );
  NAND U15039 ( .A(a[21]), .B(b[30]), .Z(n13947) );
  AND U15040 ( .A(a[20]), .B(b[31]), .Z(n13946) );
  XOR U15041 ( .A(n13948), .B(n13944), .Z(n13941) );
  XOR U15042 ( .A(n13949), .B(n13950), .Z(n13944) );
  ANDN U15043 ( .B(n13951), .A(n13952), .Z(n13949) );
  AND U15044 ( .A(a[22]), .B(b[29]), .Z(n13948) );
  XOR U15045 ( .A(n13953), .B(n13774), .Z(n13775) );
  XOR U15046 ( .A(n13954), .B(n13955), .Z(n13774) );
  AND U15047 ( .A(n13956), .B(n13957), .Z(n13954) );
  AND U15048 ( .A(a[23]), .B(b[28]), .Z(n13953) );
  XOR U15049 ( .A(n13958), .B(n13779), .Z(n13781) );
  XOR U15050 ( .A(n13959), .B(n13960), .Z(n13779) );
  AND U15051 ( .A(n13961), .B(n13962), .Z(n13959) );
  AND U15052 ( .A(a[24]), .B(b[27]), .Z(n13958) );
  XOR U15053 ( .A(n13963), .B(n13784), .Z(n13786) );
  XOR U15054 ( .A(n13964), .B(n13965), .Z(n13784) );
  AND U15055 ( .A(n13966), .B(n13967), .Z(n13964) );
  AND U15056 ( .A(a[25]), .B(b[26]), .Z(n13963) );
  XOR U15057 ( .A(n13968), .B(n13789), .Z(n13791) );
  XOR U15058 ( .A(n13969), .B(n13970), .Z(n13789) );
  AND U15059 ( .A(n13971), .B(n13972), .Z(n13969) );
  AND U15060 ( .A(b[25]), .B(a[26]), .Z(n13968) );
  XOR U15061 ( .A(n13973), .B(n13794), .Z(n13796) );
  XOR U15062 ( .A(n13974), .B(n13975), .Z(n13794) );
  AND U15063 ( .A(n13976), .B(n13977), .Z(n13974) );
  AND U15064 ( .A(a[27]), .B(b[24]), .Z(n13973) );
  XOR U15065 ( .A(n13978), .B(n13799), .Z(n13801) );
  XOR U15066 ( .A(n13979), .B(n13980), .Z(n13799) );
  AND U15067 ( .A(n13981), .B(n13982), .Z(n13979) );
  AND U15068 ( .A(b[23]), .B(a[28]), .Z(n13978) );
  XOR U15069 ( .A(n13983), .B(n13804), .Z(n13806) );
  XOR U15070 ( .A(n13984), .B(n13985), .Z(n13804) );
  AND U15071 ( .A(n13986), .B(n13987), .Z(n13984) );
  AND U15072 ( .A(a[29]), .B(b[22]), .Z(n13983) );
  XOR U15073 ( .A(n13988), .B(n13809), .Z(n13811) );
  XOR U15074 ( .A(n13989), .B(n13990), .Z(n13809) );
  AND U15075 ( .A(n13991), .B(n13992), .Z(n13989) );
  AND U15076 ( .A(b[21]), .B(a[30]), .Z(n13988) );
  XOR U15077 ( .A(n13993), .B(n13814), .Z(n13816) );
  XOR U15078 ( .A(n13994), .B(n13995), .Z(n13814) );
  AND U15079 ( .A(n13996), .B(n13997), .Z(n13994) );
  AND U15080 ( .A(a[31]), .B(b[20]), .Z(n13993) );
  XOR U15081 ( .A(n13998), .B(n13819), .Z(n13821) );
  XOR U15082 ( .A(n13999), .B(n14000), .Z(n13819) );
  AND U15083 ( .A(n14001), .B(n14002), .Z(n13999) );
  AND U15084 ( .A(a[32]), .B(b[19]), .Z(n13998) );
  XOR U15085 ( .A(n14003), .B(n13824), .Z(n13826) );
  XOR U15086 ( .A(n14004), .B(n14005), .Z(n13824) );
  AND U15087 ( .A(n14006), .B(n14007), .Z(n14004) );
  AND U15088 ( .A(a[33]), .B(b[18]), .Z(n14003) );
  XOR U15089 ( .A(n14008), .B(n13829), .Z(n13831) );
  XOR U15090 ( .A(n14009), .B(n14010), .Z(n13829) );
  AND U15091 ( .A(n14011), .B(n14012), .Z(n14009) );
  AND U15092 ( .A(a[34]), .B(b[17]), .Z(n14008) );
  XOR U15093 ( .A(n14013), .B(n13834), .Z(n13836) );
  XOR U15094 ( .A(n14014), .B(n14015), .Z(n13834) );
  AND U15095 ( .A(n14016), .B(n14017), .Z(n14014) );
  AND U15096 ( .A(a[35]), .B(b[16]), .Z(n14013) );
  XOR U15097 ( .A(n14018), .B(n14019), .Z(n13838) );
  AND U15098 ( .A(n14020), .B(n14021), .Z(n14018) );
  XOR U15099 ( .A(n14022), .B(n13843), .Z(n13845) );
  XOR U15100 ( .A(n14023), .B(n14024), .Z(n13843) );
  AND U15101 ( .A(n14025), .B(n14026), .Z(n14023) );
  AND U15102 ( .A(a[36]), .B(b[15]), .Z(n14022) );
  XOR U15103 ( .A(n14028), .B(n14029), .Z(n13848) );
  AND U15104 ( .A(n14030), .B(n14031), .Z(n14028) );
  AND U15105 ( .A(a[38]), .B(b[13]), .Z(n14027) );
  XOR U15106 ( .A(n14033), .B(n14034), .Z(n13853) );
  AND U15107 ( .A(n14035), .B(n14036), .Z(n14033) );
  AND U15108 ( .A(a[39]), .B(b[12]), .Z(n14032) );
  XOR U15109 ( .A(n14038), .B(n14039), .Z(n13858) );
  AND U15110 ( .A(n14040), .B(n14041), .Z(n14038) );
  AND U15111 ( .A(a[40]), .B(b[11]), .Z(n14037) );
  XOR U15112 ( .A(n14043), .B(n14044), .Z(n13863) );
  AND U15113 ( .A(n14045), .B(n14046), .Z(n14043) );
  AND U15114 ( .A(a[41]), .B(b[10]), .Z(n14042) );
  XOR U15115 ( .A(n14048), .B(n14049), .Z(n13868) );
  AND U15116 ( .A(n14050), .B(n14051), .Z(n14048) );
  AND U15117 ( .A(a[42]), .B(b[9]), .Z(n14047) );
  XOR U15118 ( .A(n14053), .B(n14054), .Z(n13873) );
  AND U15119 ( .A(n14055), .B(n14056), .Z(n14053) );
  AND U15120 ( .A(a[43]), .B(b[8]), .Z(n14052) );
  XOR U15121 ( .A(n14058), .B(n14059), .Z(n13878) );
  AND U15122 ( .A(n14060), .B(n14061), .Z(n14058) );
  AND U15123 ( .A(a[44]), .B(b[7]), .Z(n14057) );
  XOR U15124 ( .A(n14063), .B(n14064), .Z(n13883) );
  AND U15125 ( .A(n14065), .B(n14066), .Z(n14063) );
  AND U15126 ( .A(a[45]), .B(b[6]), .Z(n14062) );
  XOR U15127 ( .A(n14068), .B(n14069), .Z(n13888) );
  AND U15128 ( .A(n14070), .B(n14071), .Z(n14068) );
  AND U15129 ( .A(a[46]), .B(b[5]), .Z(n14067) );
  XOR U15130 ( .A(n14073), .B(n14074), .Z(n13893) );
  AND U15131 ( .A(n14075), .B(n14076), .Z(n14073) );
  AND U15132 ( .A(a[47]), .B(b[4]), .Z(n14072) );
  XOR U15133 ( .A(n14078), .B(n14079), .Z(n13898) );
  AND U15134 ( .A(n13912), .B(n13910), .Z(n14078) );
  AND U15135 ( .A(b[2]), .B(a[48]), .Z(n14080) );
  XOR U15136 ( .A(n14075), .B(n14079), .Z(n14081) );
  XOR U15137 ( .A(n14082), .B(n14083), .Z(n14079) );
  NANDN U15138 ( .A(n13914), .B(n13913), .Z(n14083) );
  XOR U15139 ( .A(n14084), .B(n14085), .Z(n13913) );
  NAND U15140 ( .A(a[48]), .B(b[1]), .Z(n14085) );
  XOR U15141 ( .A(n14086), .B(n14087), .Z(n13914) );
  XOR U15142 ( .A(n14084), .B(n14088), .Z(n14087) );
  IV U15143 ( .A(n14082), .Z(n14084) );
  ANDN U15144 ( .B(n5312), .A(n5314), .Z(n14082) );
  NAND U15145 ( .A(a[48]), .B(b[0]), .Z(n5314) );
  XNOR U15146 ( .A(n14089), .B(n14090), .Z(n5312) );
  XOR U15147 ( .A(n14070), .B(n14074), .Z(n14091) );
  XOR U15148 ( .A(n14065), .B(n14069), .Z(n14092) );
  XOR U15149 ( .A(n14060), .B(n14064), .Z(n14093) );
  XOR U15150 ( .A(n14055), .B(n14059), .Z(n14094) );
  XOR U15151 ( .A(n14050), .B(n14054), .Z(n14095) );
  XOR U15152 ( .A(n14045), .B(n14049), .Z(n14096) );
  XOR U15153 ( .A(n14040), .B(n14044), .Z(n14097) );
  XOR U15154 ( .A(n14035), .B(n14039), .Z(n14098) );
  XOR U15155 ( .A(n14030), .B(n14034), .Z(n14099) );
  XOR U15156 ( .A(n14020), .B(n14029), .Z(n14100) );
  XOR U15157 ( .A(n14101), .B(n14019), .Z(n14020) );
  AND U15158 ( .A(b[13]), .B(a[37]), .Z(n14101) );
  XNOR U15159 ( .A(n14019), .B(n14025), .Z(n14102) );
  XNOR U15160 ( .A(n14024), .B(n14016), .Z(n14103) );
  XNOR U15161 ( .A(n14015), .B(n14011), .Z(n14104) );
  XNOR U15162 ( .A(n14010), .B(n14006), .Z(n14105) );
  XNOR U15163 ( .A(n14005), .B(n14001), .Z(n14106) );
  XNOR U15164 ( .A(n14000), .B(n13996), .Z(n14107) );
  XNOR U15165 ( .A(n13995), .B(n13991), .Z(n14108) );
  XNOR U15166 ( .A(n13990), .B(n13986), .Z(n14109) );
  XNOR U15167 ( .A(n13985), .B(n13981), .Z(n14110) );
  XNOR U15168 ( .A(n13980), .B(n13976), .Z(n14111) );
  XNOR U15169 ( .A(n13975), .B(n13971), .Z(n14112) );
  XNOR U15170 ( .A(n13970), .B(n13966), .Z(n14113) );
  XNOR U15171 ( .A(n13965), .B(n13961), .Z(n14114) );
  XNOR U15172 ( .A(n13960), .B(n13956), .Z(n14115) );
  XOR U15173 ( .A(n13955), .B(n13952), .Z(n14116) );
  XOR U15174 ( .A(n14117), .B(n14118), .Z(n13952) );
  XOR U15175 ( .A(n13950), .B(n14119), .Z(n14118) );
  XOR U15176 ( .A(n14120), .B(n14121), .Z(n14119) );
  XOR U15177 ( .A(n14122), .B(n14123), .Z(n14121) );
  NAND U15178 ( .A(a[20]), .B(b[30]), .Z(n14123) );
  AND U15179 ( .A(a[19]), .B(b[31]), .Z(n14122) );
  XOR U15180 ( .A(n14124), .B(n14120), .Z(n14117) );
  XOR U15181 ( .A(n14125), .B(n14126), .Z(n14120) );
  ANDN U15182 ( .B(n14127), .A(n14128), .Z(n14125) );
  AND U15183 ( .A(a[21]), .B(b[29]), .Z(n14124) );
  XOR U15184 ( .A(n14129), .B(n13950), .Z(n13951) );
  XOR U15185 ( .A(n14130), .B(n14131), .Z(n13950) );
  AND U15186 ( .A(n14132), .B(n14133), .Z(n14130) );
  AND U15187 ( .A(a[22]), .B(b[28]), .Z(n14129) );
  XOR U15188 ( .A(n14134), .B(n13955), .Z(n13957) );
  XOR U15189 ( .A(n14135), .B(n14136), .Z(n13955) );
  AND U15190 ( .A(n14137), .B(n14138), .Z(n14135) );
  AND U15191 ( .A(a[23]), .B(b[27]), .Z(n14134) );
  XOR U15192 ( .A(n14139), .B(n13960), .Z(n13962) );
  XOR U15193 ( .A(n14140), .B(n14141), .Z(n13960) );
  AND U15194 ( .A(n14142), .B(n14143), .Z(n14140) );
  AND U15195 ( .A(a[24]), .B(b[26]), .Z(n14139) );
  XOR U15196 ( .A(n14144), .B(n13965), .Z(n13967) );
  XOR U15197 ( .A(n14145), .B(n14146), .Z(n13965) );
  AND U15198 ( .A(n14147), .B(n14148), .Z(n14145) );
  AND U15199 ( .A(a[25]), .B(b[25]), .Z(n14144) );
  XOR U15200 ( .A(n14149), .B(n13970), .Z(n13972) );
  XOR U15201 ( .A(n14150), .B(n14151), .Z(n13970) );
  AND U15202 ( .A(n14152), .B(n14153), .Z(n14150) );
  AND U15203 ( .A(b[24]), .B(a[26]), .Z(n14149) );
  XOR U15204 ( .A(n14154), .B(n13975), .Z(n13977) );
  XOR U15205 ( .A(n14155), .B(n14156), .Z(n13975) );
  AND U15206 ( .A(n14157), .B(n14158), .Z(n14155) );
  AND U15207 ( .A(a[27]), .B(b[23]), .Z(n14154) );
  XOR U15208 ( .A(n14159), .B(n13980), .Z(n13982) );
  XOR U15209 ( .A(n14160), .B(n14161), .Z(n13980) );
  AND U15210 ( .A(n14162), .B(n14163), .Z(n14160) );
  AND U15211 ( .A(b[22]), .B(a[28]), .Z(n14159) );
  XOR U15212 ( .A(n14164), .B(n13985), .Z(n13987) );
  XOR U15213 ( .A(n14165), .B(n14166), .Z(n13985) );
  AND U15214 ( .A(n14167), .B(n14168), .Z(n14165) );
  AND U15215 ( .A(a[29]), .B(b[21]), .Z(n14164) );
  XOR U15216 ( .A(n14169), .B(n13990), .Z(n13992) );
  XOR U15217 ( .A(n14170), .B(n14171), .Z(n13990) );
  AND U15218 ( .A(n14172), .B(n14173), .Z(n14170) );
  AND U15219 ( .A(b[20]), .B(a[30]), .Z(n14169) );
  XOR U15220 ( .A(n14174), .B(n13995), .Z(n13997) );
  XOR U15221 ( .A(n14175), .B(n14176), .Z(n13995) );
  AND U15222 ( .A(n14177), .B(n14178), .Z(n14175) );
  AND U15223 ( .A(a[31]), .B(b[19]), .Z(n14174) );
  XOR U15224 ( .A(n14179), .B(n14000), .Z(n14002) );
  XOR U15225 ( .A(n14180), .B(n14181), .Z(n14000) );
  AND U15226 ( .A(n14182), .B(n14183), .Z(n14180) );
  AND U15227 ( .A(a[32]), .B(b[18]), .Z(n14179) );
  XOR U15228 ( .A(n14184), .B(n14005), .Z(n14007) );
  XOR U15229 ( .A(n14185), .B(n14186), .Z(n14005) );
  AND U15230 ( .A(n14187), .B(n14188), .Z(n14185) );
  AND U15231 ( .A(a[33]), .B(b[17]), .Z(n14184) );
  XOR U15232 ( .A(n14189), .B(n14010), .Z(n14012) );
  XOR U15233 ( .A(n14190), .B(n14191), .Z(n14010) );
  AND U15234 ( .A(n14192), .B(n14193), .Z(n14190) );
  AND U15235 ( .A(a[34]), .B(b[16]), .Z(n14189) );
  XOR U15236 ( .A(n14194), .B(n14015), .Z(n14017) );
  XOR U15237 ( .A(n14195), .B(n14196), .Z(n14015) );
  AND U15238 ( .A(n14197), .B(n14198), .Z(n14195) );
  AND U15239 ( .A(a[35]), .B(b[15]), .Z(n14194) );
  XOR U15240 ( .A(n14199), .B(n14200), .Z(n14019) );
  AND U15241 ( .A(n14201), .B(n14202), .Z(n14199) );
  XOR U15242 ( .A(n14203), .B(n14024), .Z(n14026) );
  XOR U15243 ( .A(n14204), .B(n14205), .Z(n14024) );
  AND U15244 ( .A(n14206), .B(n14207), .Z(n14204) );
  AND U15245 ( .A(a[36]), .B(b[14]), .Z(n14203) );
  XOR U15246 ( .A(n14209), .B(n14210), .Z(n14029) );
  AND U15247 ( .A(n14211), .B(n14212), .Z(n14209) );
  AND U15248 ( .A(a[38]), .B(b[12]), .Z(n14208) );
  XOR U15249 ( .A(n14214), .B(n14215), .Z(n14034) );
  AND U15250 ( .A(n14216), .B(n14217), .Z(n14214) );
  AND U15251 ( .A(a[39]), .B(b[11]), .Z(n14213) );
  XOR U15252 ( .A(n14219), .B(n14220), .Z(n14039) );
  AND U15253 ( .A(n14221), .B(n14222), .Z(n14219) );
  AND U15254 ( .A(a[40]), .B(b[10]), .Z(n14218) );
  XOR U15255 ( .A(n14224), .B(n14225), .Z(n14044) );
  AND U15256 ( .A(n14226), .B(n14227), .Z(n14224) );
  AND U15257 ( .A(a[41]), .B(b[9]), .Z(n14223) );
  XOR U15258 ( .A(n14229), .B(n14230), .Z(n14049) );
  AND U15259 ( .A(n14231), .B(n14232), .Z(n14229) );
  AND U15260 ( .A(a[42]), .B(b[8]), .Z(n14228) );
  XOR U15261 ( .A(n14234), .B(n14235), .Z(n14054) );
  AND U15262 ( .A(n14236), .B(n14237), .Z(n14234) );
  AND U15263 ( .A(a[43]), .B(b[7]), .Z(n14233) );
  XOR U15264 ( .A(n14239), .B(n14240), .Z(n14059) );
  AND U15265 ( .A(n14241), .B(n14242), .Z(n14239) );
  AND U15266 ( .A(a[44]), .B(b[6]), .Z(n14238) );
  XOR U15267 ( .A(n14244), .B(n14245), .Z(n14064) );
  AND U15268 ( .A(n14246), .B(n14247), .Z(n14244) );
  AND U15269 ( .A(a[45]), .B(b[5]), .Z(n14243) );
  XOR U15270 ( .A(n14249), .B(n14250), .Z(n14069) );
  AND U15271 ( .A(n14251), .B(n14252), .Z(n14249) );
  AND U15272 ( .A(a[46]), .B(b[4]), .Z(n14248) );
  XOR U15273 ( .A(n14254), .B(n14255), .Z(n14074) );
  AND U15274 ( .A(n14088), .B(n14086), .Z(n14254) );
  AND U15275 ( .A(b[2]), .B(a[47]), .Z(n14256) );
  XOR U15276 ( .A(n14251), .B(n14255), .Z(n14257) );
  XOR U15277 ( .A(n14258), .B(n14259), .Z(n14255) );
  NANDN U15278 ( .A(n14090), .B(n14089), .Z(n14259) );
  XOR U15279 ( .A(n14260), .B(n14261), .Z(n14089) );
  NAND U15280 ( .A(a[47]), .B(b[1]), .Z(n14261) );
  XOR U15281 ( .A(n14262), .B(n14263), .Z(n14090) );
  XOR U15282 ( .A(n14260), .B(n14264), .Z(n14263) );
  IV U15283 ( .A(n14258), .Z(n14260) );
  ANDN U15284 ( .B(n5317), .A(n5319), .Z(n14258) );
  NAND U15285 ( .A(a[47]), .B(b[0]), .Z(n5319) );
  XNOR U15286 ( .A(n14265), .B(n14266), .Z(n5317) );
  XOR U15287 ( .A(n14246), .B(n14250), .Z(n14267) );
  XOR U15288 ( .A(n14241), .B(n14245), .Z(n14268) );
  XOR U15289 ( .A(n14236), .B(n14240), .Z(n14269) );
  XOR U15290 ( .A(n14231), .B(n14235), .Z(n14270) );
  XOR U15291 ( .A(n14226), .B(n14230), .Z(n14271) );
  XOR U15292 ( .A(n14221), .B(n14225), .Z(n14272) );
  XOR U15293 ( .A(n14216), .B(n14220), .Z(n14273) );
  XOR U15294 ( .A(n14211), .B(n14215), .Z(n14274) );
  XOR U15295 ( .A(n14201), .B(n14210), .Z(n14275) );
  XOR U15296 ( .A(n14276), .B(n14200), .Z(n14201) );
  AND U15297 ( .A(b[12]), .B(a[37]), .Z(n14276) );
  XNOR U15298 ( .A(n14200), .B(n14206), .Z(n14277) );
  XNOR U15299 ( .A(n14205), .B(n14197), .Z(n14278) );
  XNOR U15300 ( .A(n14196), .B(n14192), .Z(n14279) );
  XNOR U15301 ( .A(n14191), .B(n14187), .Z(n14280) );
  XNOR U15302 ( .A(n14186), .B(n14182), .Z(n14281) );
  XNOR U15303 ( .A(n14181), .B(n14177), .Z(n14282) );
  XNOR U15304 ( .A(n14176), .B(n14172), .Z(n14283) );
  XNOR U15305 ( .A(n14171), .B(n14167), .Z(n14284) );
  XNOR U15306 ( .A(n14166), .B(n14162), .Z(n14285) );
  XNOR U15307 ( .A(n14161), .B(n14157), .Z(n14286) );
  XNOR U15308 ( .A(n14156), .B(n14152), .Z(n14287) );
  XNOR U15309 ( .A(n14151), .B(n14147), .Z(n14288) );
  XNOR U15310 ( .A(n14146), .B(n14142), .Z(n14289) );
  XNOR U15311 ( .A(n14141), .B(n14137), .Z(n14290) );
  XNOR U15312 ( .A(n14136), .B(n14132), .Z(n14291) );
  XOR U15313 ( .A(n14131), .B(n14128), .Z(n14292) );
  XOR U15314 ( .A(n14293), .B(n14294), .Z(n14128) );
  XOR U15315 ( .A(n14126), .B(n14295), .Z(n14294) );
  XOR U15316 ( .A(n14296), .B(n14297), .Z(n14295) );
  XOR U15317 ( .A(n14298), .B(n14299), .Z(n14297) );
  NAND U15318 ( .A(a[19]), .B(b[30]), .Z(n14299) );
  AND U15319 ( .A(a[18]), .B(b[31]), .Z(n14298) );
  XOR U15320 ( .A(n14300), .B(n14296), .Z(n14293) );
  XOR U15321 ( .A(n14301), .B(n14302), .Z(n14296) );
  ANDN U15322 ( .B(n14303), .A(n14304), .Z(n14301) );
  AND U15323 ( .A(a[20]), .B(b[29]), .Z(n14300) );
  XOR U15324 ( .A(n14305), .B(n14126), .Z(n14127) );
  XOR U15325 ( .A(n14306), .B(n14307), .Z(n14126) );
  AND U15326 ( .A(n14308), .B(n14309), .Z(n14306) );
  AND U15327 ( .A(a[21]), .B(b[28]), .Z(n14305) );
  XOR U15328 ( .A(n14310), .B(n14131), .Z(n14133) );
  XOR U15329 ( .A(n14311), .B(n14312), .Z(n14131) );
  AND U15330 ( .A(n14313), .B(n14314), .Z(n14311) );
  AND U15331 ( .A(a[22]), .B(b[27]), .Z(n14310) );
  XOR U15332 ( .A(n14315), .B(n14136), .Z(n14138) );
  XOR U15333 ( .A(n14316), .B(n14317), .Z(n14136) );
  AND U15334 ( .A(n14318), .B(n14319), .Z(n14316) );
  AND U15335 ( .A(a[23]), .B(b[26]), .Z(n14315) );
  XOR U15336 ( .A(n14320), .B(n14141), .Z(n14143) );
  XOR U15337 ( .A(n14321), .B(n14322), .Z(n14141) );
  AND U15338 ( .A(n14323), .B(n14324), .Z(n14321) );
  AND U15339 ( .A(a[24]), .B(b[25]), .Z(n14320) );
  XOR U15340 ( .A(n14325), .B(n14146), .Z(n14148) );
  XOR U15341 ( .A(n14326), .B(n14327), .Z(n14146) );
  AND U15342 ( .A(n14328), .B(n14329), .Z(n14326) );
  AND U15343 ( .A(a[25]), .B(b[24]), .Z(n14325) );
  XOR U15344 ( .A(n14330), .B(n14151), .Z(n14153) );
  XOR U15345 ( .A(n14331), .B(n14332), .Z(n14151) );
  AND U15346 ( .A(n14333), .B(n14334), .Z(n14331) );
  AND U15347 ( .A(b[23]), .B(a[26]), .Z(n14330) );
  XOR U15348 ( .A(n14335), .B(n14156), .Z(n14158) );
  XOR U15349 ( .A(n14336), .B(n14337), .Z(n14156) );
  AND U15350 ( .A(n14338), .B(n14339), .Z(n14336) );
  AND U15351 ( .A(a[27]), .B(b[22]), .Z(n14335) );
  XOR U15352 ( .A(n14340), .B(n14161), .Z(n14163) );
  XOR U15353 ( .A(n14341), .B(n14342), .Z(n14161) );
  AND U15354 ( .A(n14343), .B(n14344), .Z(n14341) );
  AND U15355 ( .A(b[21]), .B(a[28]), .Z(n14340) );
  XOR U15356 ( .A(n14345), .B(n14166), .Z(n14168) );
  XOR U15357 ( .A(n14346), .B(n14347), .Z(n14166) );
  AND U15358 ( .A(n14348), .B(n14349), .Z(n14346) );
  AND U15359 ( .A(a[29]), .B(b[20]), .Z(n14345) );
  XOR U15360 ( .A(n14350), .B(n14171), .Z(n14173) );
  XOR U15361 ( .A(n14351), .B(n14352), .Z(n14171) );
  AND U15362 ( .A(n14353), .B(n14354), .Z(n14351) );
  AND U15363 ( .A(b[19]), .B(a[30]), .Z(n14350) );
  XOR U15364 ( .A(n14355), .B(n14176), .Z(n14178) );
  XOR U15365 ( .A(n14356), .B(n14357), .Z(n14176) );
  AND U15366 ( .A(n14358), .B(n14359), .Z(n14356) );
  AND U15367 ( .A(a[31]), .B(b[18]), .Z(n14355) );
  XOR U15368 ( .A(n14360), .B(n14181), .Z(n14183) );
  XOR U15369 ( .A(n14361), .B(n14362), .Z(n14181) );
  AND U15370 ( .A(n14363), .B(n14364), .Z(n14361) );
  AND U15371 ( .A(a[32]), .B(b[17]), .Z(n14360) );
  XOR U15372 ( .A(n14365), .B(n14186), .Z(n14188) );
  XOR U15373 ( .A(n14366), .B(n14367), .Z(n14186) );
  AND U15374 ( .A(n14368), .B(n14369), .Z(n14366) );
  AND U15375 ( .A(a[33]), .B(b[16]), .Z(n14365) );
  XOR U15376 ( .A(n14370), .B(n14191), .Z(n14193) );
  XOR U15377 ( .A(n14371), .B(n14372), .Z(n14191) );
  AND U15378 ( .A(n14373), .B(n14374), .Z(n14371) );
  AND U15379 ( .A(a[34]), .B(b[15]), .Z(n14370) );
  XOR U15380 ( .A(n14375), .B(n14196), .Z(n14198) );
  XOR U15381 ( .A(n14376), .B(n14377), .Z(n14196) );
  AND U15382 ( .A(n14378), .B(n14379), .Z(n14376) );
  AND U15383 ( .A(a[35]), .B(b[14]), .Z(n14375) );
  XOR U15384 ( .A(n14380), .B(n14381), .Z(n14200) );
  AND U15385 ( .A(n14382), .B(n14383), .Z(n14380) );
  XOR U15386 ( .A(n14384), .B(n14205), .Z(n14207) );
  XOR U15387 ( .A(n14385), .B(n14386), .Z(n14205) );
  AND U15388 ( .A(n14387), .B(n14388), .Z(n14385) );
  AND U15389 ( .A(a[36]), .B(b[13]), .Z(n14384) );
  XOR U15390 ( .A(n14390), .B(n14391), .Z(n14210) );
  AND U15391 ( .A(n14392), .B(n14393), .Z(n14390) );
  AND U15392 ( .A(a[38]), .B(b[11]), .Z(n14389) );
  XOR U15393 ( .A(n14395), .B(n14396), .Z(n14215) );
  AND U15394 ( .A(n14397), .B(n14398), .Z(n14395) );
  AND U15395 ( .A(a[39]), .B(b[10]), .Z(n14394) );
  XOR U15396 ( .A(n14400), .B(n14401), .Z(n14220) );
  AND U15397 ( .A(n14402), .B(n14403), .Z(n14400) );
  AND U15398 ( .A(a[40]), .B(b[9]), .Z(n14399) );
  XOR U15399 ( .A(n14405), .B(n14406), .Z(n14225) );
  AND U15400 ( .A(n14407), .B(n14408), .Z(n14405) );
  AND U15401 ( .A(a[41]), .B(b[8]), .Z(n14404) );
  XOR U15402 ( .A(n14410), .B(n14411), .Z(n14230) );
  AND U15403 ( .A(n14412), .B(n14413), .Z(n14410) );
  AND U15404 ( .A(a[42]), .B(b[7]), .Z(n14409) );
  XOR U15405 ( .A(n14415), .B(n14416), .Z(n14235) );
  AND U15406 ( .A(n14417), .B(n14418), .Z(n14415) );
  AND U15407 ( .A(a[43]), .B(b[6]), .Z(n14414) );
  XOR U15408 ( .A(n14420), .B(n14421), .Z(n14240) );
  AND U15409 ( .A(n14422), .B(n14423), .Z(n14420) );
  AND U15410 ( .A(a[44]), .B(b[5]), .Z(n14419) );
  XOR U15411 ( .A(n14425), .B(n14426), .Z(n14245) );
  AND U15412 ( .A(n14427), .B(n14428), .Z(n14425) );
  AND U15413 ( .A(a[45]), .B(b[4]), .Z(n14424) );
  XOR U15414 ( .A(n14430), .B(n14431), .Z(n14250) );
  AND U15415 ( .A(n14264), .B(n14262), .Z(n14430) );
  AND U15416 ( .A(b[2]), .B(a[46]), .Z(n14432) );
  XOR U15417 ( .A(n14427), .B(n14431), .Z(n14433) );
  XOR U15418 ( .A(n14434), .B(n14435), .Z(n14431) );
  NANDN U15419 ( .A(n14266), .B(n14265), .Z(n14435) );
  XOR U15420 ( .A(n14436), .B(n14437), .Z(n14265) );
  NAND U15421 ( .A(a[46]), .B(b[1]), .Z(n14437) );
  XOR U15422 ( .A(n14438), .B(n14439), .Z(n14266) );
  XOR U15423 ( .A(n14436), .B(n14440), .Z(n14439) );
  IV U15424 ( .A(n14434), .Z(n14436) );
  ANDN U15425 ( .B(n5322), .A(n5324), .Z(n14434) );
  NAND U15426 ( .A(a[46]), .B(b[0]), .Z(n5324) );
  XNOR U15427 ( .A(n14441), .B(n14442), .Z(n5322) );
  XOR U15428 ( .A(n14422), .B(n14426), .Z(n14443) );
  XOR U15429 ( .A(n14417), .B(n14421), .Z(n14444) );
  XOR U15430 ( .A(n14412), .B(n14416), .Z(n14445) );
  XOR U15431 ( .A(n14407), .B(n14411), .Z(n14446) );
  XOR U15432 ( .A(n14402), .B(n14406), .Z(n14447) );
  XOR U15433 ( .A(n14397), .B(n14401), .Z(n14448) );
  XOR U15434 ( .A(n14392), .B(n14396), .Z(n14449) );
  XOR U15435 ( .A(n14382), .B(n14391), .Z(n14450) );
  XOR U15436 ( .A(n14451), .B(n14381), .Z(n14382) );
  AND U15437 ( .A(b[11]), .B(a[37]), .Z(n14451) );
  XNOR U15438 ( .A(n14381), .B(n14387), .Z(n14452) );
  XNOR U15439 ( .A(n14386), .B(n14378), .Z(n14453) );
  XNOR U15440 ( .A(n14377), .B(n14373), .Z(n14454) );
  XNOR U15441 ( .A(n14372), .B(n14368), .Z(n14455) );
  XNOR U15442 ( .A(n14367), .B(n14363), .Z(n14456) );
  XNOR U15443 ( .A(n14362), .B(n14358), .Z(n14457) );
  XNOR U15444 ( .A(n14357), .B(n14353), .Z(n14458) );
  XNOR U15445 ( .A(n14352), .B(n14348), .Z(n14459) );
  XNOR U15446 ( .A(n14347), .B(n14343), .Z(n14460) );
  XNOR U15447 ( .A(n14342), .B(n14338), .Z(n14461) );
  XNOR U15448 ( .A(n14337), .B(n14333), .Z(n14462) );
  XNOR U15449 ( .A(n14332), .B(n14328), .Z(n14463) );
  XNOR U15450 ( .A(n14327), .B(n14323), .Z(n14464) );
  XNOR U15451 ( .A(n14322), .B(n14318), .Z(n14465) );
  XNOR U15452 ( .A(n14317), .B(n14313), .Z(n14466) );
  XNOR U15453 ( .A(n14312), .B(n14308), .Z(n14467) );
  XOR U15454 ( .A(n14307), .B(n14304), .Z(n14468) );
  XOR U15455 ( .A(n14469), .B(n14470), .Z(n14304) );
  XOR U15456 ( .A(n14302), .B(n14471), .Z(n14470) );
  XOR U15457 ( .A(n14472), .B(n14473), .Z(n14471) );
  XOR U15458 ( .A(n14474), .B(n14475), .Z(n14473) );
  NAND U15459 ( .A(a[18]), .B(b[30]), .Z(n14475) );
  AND U15460 ( .A(a[17]), .B(b[31]), .Z(n14474) );
  XOR U15461 ( .A(n14476), .B(n14472), .Z(n14469) );
  XOR U15462 ( .A(n14477), .B(n14478), .Z(n14472) );
  ANDN U15463 ( .B(n14479), .A(n14480), .Z(n14477) );
  AND U15464 ( .A(a[19]), .B(b[29]), .Z(n14476) );
  XOR U15465 ( .A(n14481), .B(n14302), .Z(n14303) );
  XOR U15466 ( .A(n14482), .B(n14483), .Z(n14302) );
  AND U15467 ( .A(n14484), .B(n14485), .Z(n14482) );
  AND U15468 ( .A(a[20]), .B(b[28]), .Z(n14481) );
  XOR U15469 ( .A(n14486), .B(n14307), .Z(n14309) );
  XOR U15470 ( .A(n14487), .B(n14488), .Z(n14307) );
  AND U15471 ( .A(n14489), .B(n14490), .Z(n14487) );
  AND U15472 ( .A(a[21]), .B(b[27]), .Z(n14486) );
  XOR U15473 ( .A(n14491), .B(n14312), .Z(n14314) );
  XOR U15474 ( .A(n14492), .B(n14493), .Z(n14312) );
  AND U15475 ( .A(n14494), .B(n14495), .Z(n14492) );
  AND U15476 ( .A(a[22]), .B(b[26]), .Z(n14491) );
  XOR U15477 ( .A(n14496), .B(n14317), .Z(n14319) );
  XOR U15478 ( .A(n14497), .B(n14498), .Z(n14317) );
  AND U15479 ( .A(n14499), .B(n14500), .Z(n14497) );
  AND U15480 ( .A(a[23]), .B(b[25]), .Z(n14496) );
  XOR U15481 ( .A(n14501), .B(n14322), .Z(n14324) );
  XOR U15482 ( .A(n14502), .B(n14503), .Z(n14322) );
  AND U15483 ( .A(n14504), .B(n14505), .Z(n14502) );
  AND U15484 ( .A(b[24]), .B(a[24]), .Z(n14501) );
  XOR U15485 ( .A(n14506), .B(n14327), .Z(n14329) );
  XOR U15486 ( .A(n14507), .B(n14508), .Z(n14327) );
  AND U15487 ( .A(n14509), .B(n14510), .Z(n14507) );
  AND U15488 ( .A(a[25]), .B(b[23]), .Z(n14506) );
  XOR U15489 ( .A(n14511), .B(n14332), .Z(n14334) );
  XOR U15490 ( .A(n14512), .B(n14513), .Z(n14332) );
  AND U15491 ( .A(n14514), .B(n14515), .Z(n14512) );
  AND U15492 ( .A(b[22]), .B(a[26]), .Z(n14511) );
  XOR U15493 ( .A(n14516), .B(n14337), .Z(n14339) );
  XOR U15494 ( .A(n14517), .B(n14518), .Z(n14337) );
  AND U15495 ( .A(n14519), .B(n14520), .Z(n14517) );
  AND U15496 ( .A(a[27]), .B(b[21]), .Z(n14516) );
  XOR U15497 ( .A(n14521), .B(n14342), .Z(n14344) );
  XOR U15498 ( .A(n14522), .B(n14523), .Z(n14342) );
  AND U15499 ( .A(n14524), .B(n14525), .Z(n14522) );
  AND U15500 ( .A(b[20]), .B(a[28]), .Z(n14521) );
  XOR U15501 ( .A(n14526), .B(n14347), .Z(n14349) );
  XOR U15502 ( .A(n14527), .B(n14528), .Z(n14347) );
  AND U15503 ( .A(n14529), .B(n14530), .Z(n14527) );
  AND U15504 ( .A(a[29]), .B(b[19]), .Z(n14526) );
  XOR U15505 ( .A(n14531), .B(n14352), .Z(n14354) );
  XOR U15506 ( .A(n14532), .B(n14533), .Z(n14352) );
  AND U15507 ( .A(n14534), .B(n14535), .Z(n14532) );
  AND U15508 ( .A(b[18]), .B(a[30]), .Z(n14531) );
  XOR U15509 ( .A(n14536), .B(n14357), .Z(n14359) );
  XOR U15510 ( .A(n14537), .B(n14538), .Z(n14357) );
  AND U15511 ( .A(n14539), .B(n14540), .Z(n14537) );
  AND U15512 ( .A(a[31]), .B(b[17]), .Z(n14536) );
  XOR U15513 ( .A(n14541), .B(n14362), .Z(n14364) );
  XOR U15514 ( .A(n14542), .B(n14543), .Z(n14362) );
  AND U15515 ( .A(n14544), .B(n14545), .Z(n14542) );
  AND U15516 ( .A(a[32]), .B(b[16]), .Z(n14541) );
  XOR U15517 ( .A(n14546), .B(n14367), .Z(n14369) );
  XOR U15518 ( .A(n14547), .B(n14548), .Z(n14367) );
  AND U15519 ( .A(n14549), .B(n14550), .Z(n14547) );
  AND U15520 ( .A(a[33]), .B(b[15]), .Z(n14546) );
  XOR U15521 ( .A(n14551), .B(n14372), .Z(n14374) );
  XOR U15522 ( .A(n14552), .B(n14553), .Z(n14372) );
  AND U15523 ( .A(n14554), .B(n14555), .Z(n14552) );
  AND U15524 ( .A(a[34]), .B(b[14]), .Z(n14551) );
  XOR U15525 ( .A(n14556), .B(n14377), .Z(n14379) );
  XOR U15526 ( .A(n14557), .B(n14558), .Z(n14377) );
  AND U15527 ( .A(n14559), .B(n14560), .Z(n14557) );
  AND U15528 ( .A(a[35]), .B(b[13]), .Z(n14556) );
  XOR U15529 ( .A(n14561), .B(n14562), .Z(n14381) );
  AND U15530 ( .A(n14563), .B(n14564), .Z(n14561) );
  XOR U15531 ( .A(n14565), .B(n14386), .Z(n14388) );
  XOR U15532 ( .A(n14566), .B(n14567), .Z(n14386) );
  AND U15533 ( .A(n14568), .B(n14569), .Z(n14566) );
  AND U15534 ( .A(a[36]), .B(b[12]), .Z(n14565) );
  XOR U15535 ( .A(n14571), .B(n14572), .Z(n14391) );
  AND U15536 ( .A(n14573), .B(n14574), .Z(n14571) );
  AND U15537 ( .A(a[38]), .B(b[10]), .Z(n14570) );
  XOR U15538 ( .A(n14576), .B(n14577), .Z(n14396) );
  AND U15539 ( .A(n14578), .B(n14579), .Z(n14576) );
  AND U15540 ( .A(a[39]), .B(b[9]), .Z(n14575) );
  XOR U15541 ( .A(n14581), .B(n14582), .Z(n14401) );
  AND U15542 ( .A(n14583), .B(n14584), .Z(n14581) );
  AND U15543 ( .A(a[40]), .B(b[8]), .Z(n14580) );
  XOR U15544 ( .A(n14586), .B(n14587), .Z(n14406) );
  AND U15545 ( .A(n14588), .B(n14589), .Z(n14586) );
  AND U15546 ( .A(a[41]), .B(b[7]), .Z(n14585) );
  XOR U15547 ( .A(n14591), .B(n14592), .Z(n14411) );
  AND U15548 ( .A(n14593), .B(n14594), .Z(n14591) );
  AND U15549 ( .A(a[42]), .B(b[6]), .Z(n14590) );
  XOR U15550 ( .A(n14596), .B(n14597), .Z(n14416) );
  AND U15551 ( .A(n14598), .B(n14599), .Z(n14596) );
  AND U15552 ( .A(a[43]), .B(b[5]), .Z(n14595) );
  XOR U15553 ( .A(n14601), .B(n14602), .Z(n14421) );
  AND U15554 ( .A(n14603), .B(n14604), .Z(n14601) );
  AND U15555 ( .A(a[44]), .B(b[4]), .Z(n14600) );
  XOR U15556 ( .A(n14606), .B(n14607), .Z(n14426) );
  AND U15557 ( .A(n14440), .B(n14438), .Z(n14606) );
  AND U15558 ( .A(b[2]), .B(a[45]), .Z(n14608) );
  XOR U15559 ( .A(n14603), .B(n14607), .Z(n14609) );
  XOR U15560 ( .A(n14610), .B(n14611), .Z(n14607) );
  NANDN U15561 ( .A(n14442), .B(n14441), .Z(n14611) );
  XOR U15562 ( .A(n14612), .B(n14613), .Z(n14441) );
  NAND U15563 ( .A(a[45]), .B(b[1]), .Z(n14613) );
  XOR U15564 ( .A(n14614), .B(n14615), .Z(n14442) );
  XOR U15565 ( .A(n14612), .B(n14616), .Z(n14615) );
  IV U15566 ( .A(n14610), .Z(n14612) );
  ANDN U15567 ( .B(n5327), .A(n5329), .Z(n14610) );
  NAND U15568 ( .A(a[45]), .B(b[0]), .Z(n5329) );
  XNOR U15569 ( .A(n14617), .B(n14618), .Z(n5327) );
  XOR U15570 ( .A(n14598), .B(n14602), .Z(n14619) );
  XOR U15571 ( .A(n14593), .B(n14597), .Z(n14620) );
  XOR U15572 ( .A(n14588), .B(n14592), .Z(n14621) );
  XOR U15573 ( .A(n14583), .B(n14587), .Z(n14622) );
  XOR U15574 ( .A(n14578), .B(n14582), .Z(n14623) );
  XOR U15575 ( .A(n14573), .B(n14577), .Z(n14624) );
  XOR U15576 ( .A(n14563), .B(n14572), .Z(n14625) );
  XOR U15577 ( .A(n14626), .B(n14562), .Z(n14563) );
  AND U15578 ( .A(b[10]), .B(a[37]), .Z(n14626) );
  XNOR U15579 ( .A(n14562), .B(n14568), .Z(n14627) );
  XNOR U15580 ( .A(n14567), .B(n14559), .Z(n14628) );
  XNOR U15581 ( .A(n14558), .B(n14554), .Z(n14629) );
  XNOR U15582 ( .A(n14553), .B(n14549), .Z(n14630) );
  XNOR U15583 ( .A(n14548), .B(n14544), .Z(n14631) );
  XNOR U15584 ( .A(n14543), .B(n14539), .Z(n14632) );
  XNOR U15585 ( .A(n14538), .B(n14534), .Z(n14633) );
  XNOR U15586 ( .A(n14533), .B(n14529), .Z(n14634) );
  XNOR U15587 ( .A(n14528), .B(n14524), .Z(n14635) );
  XNOR U15588 ( .A(n14523), .B(n14519), .Z(n14636) );
  XNOR U15589 ( .A(n14518), .B(n14514), .Z(n14637) );
  XNOR U15590 ( .A(n14513), .B(n14509), .Z(n14638) );
  XNOR U15591 ( .A(n14508), .B(n14504), .Z(n14639) );
  XNOR U15592 ( .A(n14503), .B(n14499), .Z(n14640) );
  XNOR U15593 ( .A(n14498), .B(n14494), .Z(n14641) );
  XNOR U15594 ( .A(n14493), .B(n14489), .Z(n14642) );
  XNOR U15595 ( .A(n14488), .B(n14484), .Z(n14643) );
  XOR U15596 ( .A(n14483), .B(n14480), .Z(n14644) );
  XOR U15597 ( .A(n14645), .B(n14646), .Z(n14480) );
  XOR U15598 ( .A(n14478), .B(n14647), .Z(n14646) );
  XOR U15599 ( .A(n14648), .B(n14649), .Z(n14647) );
  XOR U15600 ( .A(n14650), .B(n14651), .Z(n14649) );
  NAND U15601 ( .A(a[17]), .B(b[30]), .Z(n14651) );
  AND U15602 ( .A(a[16]), .B(b[31]), .Z(n14650) );
  XOR U15603 ( .A(n14652), .B(n14648), .Z(n14645) );
  XOR U15604 ( .A(n14653), .B(n14654), .Z(n14648) );
  ANDN U15605 ( .B(n14655), .A(n14656), .Z(n14653) );
  AND U15606 ( .A(a[18]), .B(b[29]), .Z(n14652) );
  XOR U15607 ( .A(n14657), .B(n14478), .Z(n14479) );
  XOR U15608 ( .A(n14658), .B(n14659), .Z(n14478) );
  AND U15609 ( .A(n14660), .B(n14661), .Z(n14658) );
  AND U15610 ( .A(a[19]), .B(b[28]), .Z(n14657) );
  XOR U15611 ( .A(n14662), .B(n14483), .Z(n14485) );
  XOR U15612 ( .A(n14663), .B(n14664), .Z(n14483) );
  AND U15613 ( .A(n14665), .B(n14666), .Z(n14663) );
  AND U15614 ( .A(a[20]), .B(b[27]), .Z(n14662) );
  XOR U15615 ( .A(n14667), .B(n14488), .Z(n14490) );
  XOR U15616 ( .A(n14668), .B(n14669), .Z(n14488) );
  AND U15617 ( .A(n14670), .B(n14671), .Z(n14668) );
  AND U15618 ( .A(a[21]), .B(b[26]), .Z(n14667) );
  XOR U15619 ( .A(n14672), .B(n14493), .Z(n14495) );
  XOR U15620 ( .A(n14673), .B(n14674), .Z(n14493) );
  AND U15621 ( .A(n14675), .B(n14676), .Z(n14673) );
  AND U15622 ( .A(a[22]), .B(b[25]), .Z(n14672) );
  XOR U15623 ( .A(n14677), .B(n14498), .Z(n14500) );
  XOR U15624 ( .A(n14678), .B(n14679), .Z(n14498) );
  AND U15625 ( .A(n14680), .B(n14681), .Z(n14678) );
  AND U15626 ( .A(a[23]), .B(b[24]), .Z(n14677) );
  XOR U15627 ( .A(n14682), .B(n14503), .Z(n14505) );
  XOR U15628 ( .A(n14683), .B(n14684), .Z(n14503) );
  AND U15629 ( .A(n14685), .B(n14686), .Z(n14683) );
  AND U15630 ( .A(b[23]), .B(a[24]), .Z(n14682) );
  XOR U15631 ( .A(n14687), .B(n14508), .Z(n14510) );
  XOR U15632 ( .A(n14688), .B(n14689), .Z(n14508) );
  AND U15633 ( .A(n14690), .B(n14691), .Z(n14688) );
  AND U15634 ( .A(a[25]), .B(b[22]), .Z(n14687) );
  XOR U15635 ( .A(n14692), .B(n14513), .Z(n14515) );
  XOR U15636 ( .A(n14693), .B(n14694), .Z(n14513) );
  AND U15637 ( .A(n14695), .B(n14696), .Z(n14693) );
  AND U15638 ( .A(b[21]), .B(a[26]), .Z(n14692) );
  XOR U15639 ( .A(n14697), .B(n14518), .Z(n14520) );
  XOR U15640 ( .A(n14698), .B(n14699), .Z(n14518) );
  AND U15641 ( .A(n14700), .B(n14701), .Z(n14698) );
  AND U15642 ( .A(a[27]), .B(b[20]), .Z(n14697) );
  XOR U15643 ( .A(n14702), .B(n14523), .Z(n14525) );
  XOR U15644 ( .A(n14703), .B(n14704), .Z(n14523) );
  AND U15645 ( .A(n14705), .B(n14706), .Z(n14703) );
  AND U15646 ( .A(b[19]), .B(a[28]), .Z(n14702) );
  XOR U15647 ( .A(n14707), .B(n14528), .Z(n14530) );
  XOR U15648 ( .A(n14708), .B(n14709), .Z(n14528) );
  AND U15649 ( .A(n14710), .B(n14711), .Z(n14708) );
  AND U15650 ( .A(a[29]), .B(b[18]), .Z(n14707) );
  XOR U15651 ( .A(n14712), .B(n14533), .Z(n14535) );
  XOR U15652 ( .A(n14713), .B(n14714), .Z(n14533) );
  AND U15653 ( .A(n14715), .B(n14716), .Z(n14713) );
  AND U15654 ( .A(b[17]), .B(a[30]), .Z(n14712) );
  XOR U15655 ( .A(n14717), .B(n14538), .Z(n14540) );
  XOR U15656 ( .A(n14718), .B(n14719), .Z(n14538) );
  AND U15657 ( .A(n14720), .B(n14721), .Z(n14718) );
  AND U15658 ( .A(a[31]), .B(b[16]), .Z(n14717) );
  XOR U15659 ( .A(n14722), .B(n14543), .Z(n14545) );
  XOR U15660 ( .A(n14723), .B(n14724), .Z(n14543) );
  AND U15661 ( .A(n14725), .B(n14726), .Z(n14723) );
  AND U15662 ( .A(a[32]), .B(b[15]), .Z(n14722) );
  XOR U15663 ( .A(n14727), .B(n14548), .Z(n14550) );
  XOR U15664 ( .A(n14728), .B(n14729), .Z(n14548) );
  AND U15665 ( .A(n14730), .B(n14731), .Z(n14728) );
  AND U15666 ( .A(a[33]), .B(b[14]), .Z(n14727) );
  XOR U15667 ( .A(n14732), .B(n14553), .Z(n14555) );
  XOR U15668 ( .A(n14733), .B(n14734), .Z(n14553) );
  AND U15669 ( .A(n14735), .B(n14736), .Z(n14733) );
  AND U15670 ( .A(a[34]), .B(b[13]), .Z(n14732) );
  XOR U15671 ( .A(n14737), .B(n14558), .Z(n14560) );
  XOR U15672 ( .A(n14738), .B(n14739), .Z(n14558) );
  AND U15673 ( .A(n14740), .B(n14741), .Z(n14738) );
  AND U15674 ( .A(a[35]), .B(b[12]), .Z(n14737) );
  XOR U15675 ( .A(n14742), .B(n14743), .Z(n14562) );
  AND U15676 ( .A(n14744), .B(n14745), .Z(n14742) );
  XOR U15677 ( .A(n14746), .B(n14567), .Z(n14569) );
  XOR U15678 ( .A(n14747), .B(n14748), .Z(n14567) );
  AND U15679 ( .A(n14749), .B(n14750), .Z(n14747) );
  AND U15680 ( .A(a[36]), .B(b[11]), .Z(n14746) );
  XOR U15681 ( .A(n14752), .B(n14753), .Z(n14572) );
  AND U15682 ( .A(n14754), .B(n14755), .Z(n14752) );
  AND U15683 ( .A(a[38]), .B(b[9]), .Z(n14751) );
  XOR U15684 ( .A(n14757), .B(n14758), .Z(n14577) );
  AND U15685 ( .A(n14759), .B(n14760), .Z(n14757) );
  AND U15686 ( .A(a[39]), .B(b[8]), .Z(n14756) );
  XOR U15687 ( .A(n14762), .B(n14763), .Z(n14582) );
  AND U15688 ( .A(n14764), .B(n14765), .Z(n14762) );
  AND U15689 ( .A(a[40]), .B(b[7]), .Z(n14761) );
  XOR U15690 ( .A(n14767), .B(n14768), .Z(n14587) );
  AND U15691 ( .A(n14769), .B(n14770), .Z(n14767) );
  AND U15692 ( .A(a[41]), .B(b[6]), .Z(n14766) );
  XOR U15693 ( .A(n14772), .B(n14773), .Z(n14592) );
  AND U15694 ( .A(n14774), .B(n14775), .Z(n14772) );
  AND U15695 ( .A(a[42]), .B(b[5]), .Z(n14771) );
  XOR U15696 ( .A(n14777), .B(n14778), .Z(n14597) );
  AND U15697 ( .A(n14779), .B(n14780), .Z(n14777) );
  AND U15698 ( .A(a[43]), .B(b[4]), .Z(n14776) );
  XOR U15699 ( .A(n14782), .B(n14783), .Z(n14602) );
  AND U15700 ( .A(n14616), .B(n14614), .Z(n14782) );
  AND U15701 ( .A(b[2]), .B(a[44]), .Z(n14784) );
  XOR U15702 ( .A(n14779), .B(n14783), .Z(n14785) );
  XOR U15703 ( .A(n14786), .B(n14787), .Z(n14783) );
  NANDN U15704 ( .A(n14618), .B(n14617), .Z(n14787) );
  XOR U15705 ( .A(n14788), .B(n14789), .Z(n14617) );
  NAND U15706 ( .A(a[44]), .B(b[1]), .Z(n14789) );
  XOR U15707 ( .A(n14790), .B(n14791), .Z(n14618) );
  XOR U15708 ( .A(n14788), .B(n14792), .Z(n14791) );
  IV U15709 ( .A(n14786), .Z(n14788) );
  ANDN U15710 ( .B(n5332), .A(n5334), .Z(n14786) );
  NAND U15711 ( .A(a[44]), .B(b[0]), .Z(n5334) );
  XNOR U15712 ( .A(n14793), .B(n14794), .Z(n5332) );
  XOR U15713 ( .A(n14774), .B(n14778), .Z(n14795) );
  XOR U15714 ( .A(n14769), .B(n14773), .Z(n14796) );
  XOR U15715 ( .A(n14764), .B(n14768), .Z(n14797) );
  XOR U15716 ( .A(n14759), .B(n14763), .Z(n14798) );
  XOR U15717 ( .A(n14754), .B(n14758), .Z(n14799) );
  XOR U15718 ( .A(n14744), .B(n14753), .Z(n14800) );
  XOR U15719 ( .A(n14801), .B(n14743), .Z(n14744) );
  AND U15720 ( .A(b[9]), .B(a[37]), .Z(n14801) );
  XNOR U15721 ( .A(n14743), .B(n14749), .Z(n14802) );
  XNOR U15722 ( .A(n14748), .B(n14740), .Z(n14803) );
  XNOR U15723 ( .A(n14739), .B(n14735), .Z(n14804) );
  XNOR U15724 ( .A(n14734), .B(n14730), .Z(n14805) );
  XNOR U15725 ( .A(n14729), .B(n14725), .Z(n14806) );
  XNOR U15726 ( .A(n14724), .B(n14720), .Z(n14807) );
  XNOR U15727 ( .A(n14719), .B(n14715), .Z(n14808) );
  XNOR U15728 ( .A(n14714), .B(n14710), .Z(n14809) );
  XNOR U15729 ( .A(n14709), .B(n14705), .Z(n14810) );
  XNOR U15730 ( .A(n14704), .B(n14700), .Z(n14811) );
  XNOR U15731 ( .A(n14699), .B(n14695), .Z(n14812) );
  XNOR U15732 ( .A(n14694), .B(n14690), .Z(n14813) );
  XNOR U15733 ( .A(n14689), .B(n14685), .Z(n14814) );
  XNOR U15734 ( .A(n14684), .B(n14680), .Z(n14815) );
  XNOR U15735 ( .A(n14679), .B(n14675), .Z(n14816) );
  XNOR U15736 ( .A(n14674), .B(n14670), .Z(n14817) );
  XNOR U15737 ( .A(n14669), .B(n14665), .Z(n14818) );
  XNOR U15738 ( .A(n14664), .B(n14660), .Z(n14819) );
  XOR U15739 ( .A(n14659), .B(n14656), .Z(n14820) );
  XOR U15740 ( .A(n14821), .B(n14822), .Z(n14656) );
  XOR U15741 ( .A(n14654), .B(n14823), .Z(n14822) );
  XOR U15742 ( .A(n14824), .B(n14825), .Z(n14823) );
  XOR U15743 ( .A(n14826), .B(n14827), .Z(n14825) );
  NAND U15744 ( .A(a[16]), .B(b[30]), .Z(n14827) );
  AND U15745 ( .A(a[15]), .B(b[31]), .Z(n14826) );
  XOR U15746 ( .A(n14828), .B(n14824), .Z(n14821) );
  XOR U15747 ( .A(n14829), .B(n14830), .Z(n14824) );
  ANDN U15748 ( .B(n14831), .A(n14832), .Z(n14829) );
  AND U15749 ( .A(a[17]), .B(b[29]), .Z(n14828) );
  XOR U15750 ( .A(n14833), .B(n14654), .Z(n14655) );
  XOR U15751 ( .A(n14834), .B(n14835), .Z(n14654) );
  AND U15752 ( .A(n14836), .B(n14837), .Z(n14834) );
  AND U15753 ( .A(a[18]), .B(b[28]), .Z(n14833) );
  XOR U15754 ( .A(n14838), .B(n14659), .Z(n14661) );
  XOR U15755 ( .A(n14839), .B(n14840), .Z(n14659) );
  AND U15756 ( .A(n14841), .B(n14842), .Z(n14839) );
  AND U15757 ( .A(a[19]), .B(b[27]), .Z(n14838) );
  XOR U15758 ( .A(n14843), .B(n14664), .Z(n14666) );
  XOR U15759 ( .A(n14844), .B(n14845), .Z(n14664) );
  AND U15760 ( .A(n14846), .B(n14847), .Z(n14844) );
  AND U15761 ( .A(a[20]), .B(b[26]), .Z(n14843) );
  XOR U15762 ( .A(n14848), .B(n14669), .Z(n14671) );
  XOR U15763 ( .A(n14849), .B(n14850), .Z(n14669) );
  AND U15764 ( .A(n14851), .B(n14852), .Z(n14849) );
  AND U15765 ( .A(a[21]), .B(b[25]), .Z(n14848) );
  XOR U15766 ( .A(n14853), .B(n14674), .Z(n14676) );
  XOR U15767 ( .A(n14854), .B(n14855), .Z(n14674) );
  AND U15768 ( .A(n14856), .B(n14857), .Z(n14854) );
  AND U15769 ( .A(a[22]), .B(b[24]), .Z(n14853) );
  XOR U15770 ( .A(n14858), .B(n14679), .Z(n14681) );
  XOR U15771 ( .A(n14859), .B(n14860), .Z(n14679) );
  AND U15772 ( .A(n14861), .B(n14862), .Z(n14859) );
  AND U15773 ( .A(a[23]), .B(b[23]), .Z(n14858) );
  XOR U15774 ( .A(n14863), .B(n14684), .Z(n14686) );
  XOR U15775 ( .A(n14864), .B(n14865), .Z(n14684) );
  AND U15776 ( .A(n14866), .B(n14867), .Z(n14864) );
  AND U15777 ( .A(b[22]), .B(a[24]), .Z(n14863) );
  XOR U15778 ( .A(n14868), .B(n14689), .Z(n14691) );
  XOR U15779 ( .A(n14869), .B(n14870), .Z(n14689) );
  AND U15780 ( .A(n14871), .B(n14872), .Z(n14869) );
  AND U15781 ( .A(a[25]), .B(b[21]), .Z(n14868) );
  XOR U15782 ( .A(n14873), .B(n14694), .Z(n14696) );
  XOR U15783 ( .A(n14874), .B(n14875), .Z(n14694) );
  AND U15784 ( .A(n14876), .B(n14877), .Z(n14874) );
  AND U15785 ( .A(b[20]), .B(a[26]), .Z(n14873) );
  XOR U15786 ( .A(n14878), .B(n14699), .Z(n14701) );
  XOR U15787 ( .A(n14879), .B(n14880), .Z(n14699) );
  AND U15788 ( .A(n14881), .B(n14882), .Z(n14879) );
  AND U15789 ( .A(a[27]), .B(b[19]), .Z(n14878) );
  XOR U15790 ( .A(n14883), .B(n14704), .Z(n14706) );
  XOR U15791 ( .A(n14884), .B(n14885), .Z(n14704) );
  AND U15792 ( .A(n14886), .B(n14887), .Z(n14884) );
  AND U15793 ( .A(b[18]), .B(a[28]), .Z(n14883) );
  XOR U15794 ( .A(n14888), .B(n14709), .Z(n14711) );
  XOR U15795 ( .A(n14889), .B(n14890), .Z(n14709) );
  AND U15796 ( .A(n14891), .B(n14892), .Z(n14889) );
  AND U15797 ( .A(a[29]), .B(b[17]), .Z(n14888) );
  XOR U15798 ( .A(n14893), .B(n14714), .Z(n14716) );
  XOR U15799 ( .A(n14894), .B(n14895), .Z(n14714) );
  AND U15800 ( .A(n14896), .B(n14897), .Z(n14894) );
  AND U15801 ( .A(b[16]), .B(a[30]), .Z(n14893) );
  XOR U15802 ( .A(n14898), .B(n14719), .Z(n14721) );
  XOR U15803 ( .A(n14899), .B(n14900), .Z(n14719) );
  AND U15804 ( .A(n14901), .B(n14902), .Z(n14899) );
  AND U15805 ( .A(a[31]), .B(b[15]), .Z(n14898) );
  XOR U15806 ( .A(n14903), .B(n14724), .Z(n14726) );
  XOR U15807 ( .A(n14904), .B(n14905), .Z(n14724) );
  AND U15808 ( .A(n14906), .B(n14907), .Z(n14904) );
  AND U15809 ( .A(a[32]), .B(b[14]), .Z(n14903) );
  XOR U15810 ( .A(n14908), .B(n14729), .Z(n14731) );
  XOR U15811 ( .A(n14909), .B(n14910), .Z(n14729) );
  AND U15812 ( .A(n14911), .B(n14912), .Z(n14909) );
  AND U15813 ( .A(a[33]), .B(b[13]), .Z(n14908) );
  XOR U15814 ( .A(n14913), .B(n14734), .Z(n14736) );
  XOR U15815 ( .A(n14914), .B(n14915), .Z(n14734) );
  AND U15816 ( .A(n14916), .B(n14917), .Z(n14914) );
  AND U15817 ( .A(a[34]), .B(b[12]), .Z(n14913) );
  XOR U15818 ( .A(n14918), .B(n14739), .Z(n14741) );
  XOR U15819 ( .A(n14919), .B(n14920), .Z(n14739) );
  AND U15820 ( .A(n14921), .B(n14922), .Z(n14919) );
  AND U15821 ( .A(a[35]), .B(b[11]), .Z(n14918) );
  XOR U15822 ( .A(n14923), .B(n14924), .Z(n14743) );
  AND U15823 ( .A(n14925), .B(n14926), .Z(n14923) );
  XOR U15824 ( .A(n14927), .B(n14748), .Z(n14750) );
  XOR U15825 ( .A(n14928), .B(n14929), .Z(n14748) );
  AND U15826 ( .A(n14930), .B(n14931), .Z(n14928) );
  AND U15827 ( .A(a[36]), .B(b[10]), .Z(n14927) );
  XOR U15828 ( .A(n14933), .B(n14934), .Z(n14753) );
  AND U15829 ( .A(n14935), .B(n14936), .Z(n14933) );
  AND U15830 ( .A(a[38]), .B(b[8]), .Z(n14932) );
  XOR U15831 ( .A(n14938), .B(n14939), .Z(n14758) );
  AND U15832 ( .A(n14940), .B(n14941), .Z(n14938) );
  AND U15833 ( .A(a[39]), .B(b[7]), .Z(n14937) );
  XOR U15834 ( .A(n14943), .B(n14944), .Z(n14763) );
  AND U15835 ( .A(n14945), .B(n14946), .Z(n14943) );
  AND U15836 ( .A(a[40]), .B(b[6]), .Z(n14942) );
  XOR U15837 ( .A(n14948), .B(n14949), .Z(n14768) );
  AND U15838 ( .A(n14950), .B(n14951), .Z(n14948) );
  AND U15839 ( .A(a[41]), .B(b[5]), .Z(n14947) );
  XOR U15840 ( .A(n14953), .B(n14954), .Z(n14773) );
  AND U15841 ( .A(n14955), .B(n14956), .Z(n14953) );
  AND U15842 ( .A(a[42]), .B(b[4]), .Z(n14952) );
  XOR U15843 ( .A(n14958), .B(n14959), .Z(n14778) );
  AND U15844 ( .A(n14792), .B(n14790), .Z(n14958) );
  AND U15845 ( .A(b[2]), .B(a[43]), .Z(n14960) );
  XOR U15846 ( .A(n14955), .B(n14959), .Z(n14961) );
  XOR U15847 ( .A(n14962), .B(n14963), .Z(n14959) );
  NANDN U15848 ( .A(n14794), .B(n14793), .Z(n14963) );
  XOR U15849 ( .A(n14964), .B(n14965), .Z(n14793) );
  NAND U15850 ( .A(a[43]), .B(b[1]), .Z(n14965) );
  XOR U15851 ( .A(n14966), .B(n14967), .Z(n14794) );
  XOR U15852 ( .A(n14964), .B(n14968), .Z(n14967) );
  IV U15853 ( .A(n14962), .Z(n14964) );
  ANDN U15854 ( .B(n5337), .A(n5339), .Z(n14962) );
  NAND U15855 ( .A(a[43]), .B(b[0]), .Z(n5339) );
  XNOR U15856 ( .A(n14969), .B(n14970), .Z(n5337) );
  XOR U15857 ( .A(n14950), .B(n14954), .Z(n14971) );
  XOR U15858 ( .A(n14945), .B(n14949), .Z(n14972) );
  XOR U15859 ( .A(n14940), .B(n14944), .Z(n14973) );
  XOR U15860 ( .A(n14935), .B(n14939), .Z(n14974) );
  XOR U15861 ( .A(n14925), .B(n14934), .Z(n14975) );
  XOR U15862 ( .A(n14976), .B(n14924), .Z(n14925) );
  AND U15863 ( .A(b[8]), .B(a[37]), .Z(n14976) );
  XNOR U15864 ( .A(n14924), .B(n14930), .Z(n14977) );
  XNOR U15865 ( .A(n14929), .B(n14921), .Z(n14978) );
  XNOR U15866 ( .A(n14920), .B(n14916), .Z(n14979) );
  XNOR U15867 ( .A(n14915), .B(n14911), .Z(n14980) );
  XNOR U15868 ( .A(n14910), .B(n14906), .Z(n14981) );
  XNOR U15869 ( .A(n14905), .B(n14901), .Z(n14982) );
  XNOR U15870 ( .A(n14900), .B(n14896), .Z(n14983) );
  XNOR U15871 ( .A(n14895), .B(n14891), .Z(n14984) );
  XNOR U15872 ( .A(n14890), .B(n14886), .Z(n14985) );
  XNOR U15873 ( .A(n14885), .B(n14881), .Z(n14986) );
  XNOR U15874 ( .A(n14880), .B(n14876), .Z(n14987) );
  XNOR U15875 ( .A(n14875), .B(n14871), .Z(n14988) );
  XNOR U15876 ( .A(n14870), .B(n14866), .Z(n14989) );
  XNOR U15877 ( .A(n14865), .B(n14861), .Z(n14990) );
  XNOR U15878 ( .A(n14860), .B(n14856), .Z(n14991) );
  XNOR U15879 ( .A(n14855), .B(n14851), .Z(n14992) );
  XNOR U15880 ( .A(n14850), .B(n14846), .Z(n14993) );
  XNOR U15881 ( .A(n14845), .B(n14841), .Z(n14994) );
  XNOR U15882 ( .A(n14840), .B(n14836), .Z(n14995) );
  XOR U15883 ( .A(n14835), .B(n14832), .Z(n14996) );
  XOR U15884 ( .A(n14997), .B(n14998), .Z(n14832) );
  XOR U15885 ( .A(n14830), .B(n14999), .Z(n14998) );
  XOR U15886 ( .A(n15000), .B(n15001), .Z(n14999) );
  XOR U15887 ( .A(n15002), .B(n15003), .Z(n15001) );
  NAND U15888 ( .A(a[15]), .B(b[30]), .Z(n15003) );
  AND U15889 ( .A(a[14]), .B(b[31]), .Z(n15002) );
  XOR U15890 ( .A(n15004), .B(n15000), .Z(n14997) );
  XOR U15891 ( .A(n15005), .B(n15006), .Z(n15000) );
  ANDN U15892 ( .B(n15007), .A(n15008), .Z(n15005) );
  AND U15893 ( .A(a[16]), .B(b[29]), .Z(n15004) );
  XOR U15894 ( .A(n15009), .B(n14830), .Z(n14831) );
  XOR U15895 ( .A(n15010), .B(n15011), .Z(n14830) );
  AND U15896 ( .A(n15012), .B(n15013), .Z(n15010) );
  AND U15897 ( .A(a[17]), .B(b[28]), .Z(n15009) );
  XOR U15898 ( .A(n15014), .B(n14835), .Z(n14837) );
  XOR U15899 ( .A(n15015), .B(n15016), .Z(n14835) );
  AND U15900 ( .A(n15017), .B(n15018), .Z(n15015) );
  AND U15901 ( .A(a[18]), .B(b[27]), .Z(n15014) );
  XOR U15902 ( .A(n15019), .B(n14840), .Z(n14842) );
  XOR U15903 ( .A(n15020), .B(n15021), .Z(n14840) );
  AND U15904 ( .A(n15022), .B(n15023), .Z(n15020) );
  AND U15905 ( .A(a[19]), .B(b[26]), .Z(n15019) );
  XOR U15906 ( .A(n15024), .B(n14845), .Z(n14847) );
  XOR U15907 ( .A(n15025), .B(n15026), .Z(n14845) );
  AND U15908 ( .A(n15027), .B(n15028), .Z(n15025) );
  AND U15909 ( .A(a[20]), .B(b[25]), .Z(n15024) );
  XOR U15910 ( .A(n15029), .B(n14850), .Z(n14852) );
  XOR U15911 ( .A(n15030), .B(n15031), .Z(n14850) );
  AND U15912 ( .A(n15032), .B(n15033), .Z(n15030) );
  AND U15913 ( .A(a[21]), .B(b[24]), .Z(n15029) );
  XOR U15914 ( .A(n15034), .B(n14855), .Z(n14857) );
  XOR U15915 ( .A(n15035), .B(n15036), .Z(n14855) );
  AND U15916 ( .A(n15037), .B(n15038), .Z(n15035) );
  AND U15917 ( .A(a[22]), .B(b[23]), .Z(n15034) );
  XOR U15918 ( .A(n15039), .B(n14860), .Z(n14862) );
  XOR U15919 ( .A(n15040), .B(n15041), .Z(n14860) );
  AND U15920 ( .A(n15042), .B(n15043), .Z(n15040) );
  AND U15921 ( .A(a[23]), .B(b[22]), .Z(n15039) );
  XOR U15922 ( .A(n15044), .B(n14865), .Z(n14867) );
  XOR U15923 ( .A(n15045), .B(n15046), .Z(n14865) );
  AND U15924 ( .A(n15047), .B(n15048), .Z(n15045) );
  AND U15925 ( .A(b[21]), .B(a[24]), .Z(n15044) );
  XOR U15926 ( .A(n15049), .B(n14870), .Z(n14872) );
  XOR U15927 ( .A(n15050), .B(n15051), .Z(n14870) );
  AND U15928 ( .A(n15052), .B(n15053), .Z(n15050) );
  AND U15929 ( .A(a[25]), .B(b[20]), .Z(n15049) );
  XOR U15930 ( .A(n15054), .B(n14875), .Z(n14877) );
  XOR U15931 ( .A(n15055), .B(n15056), .Z(n14875) );
  AND U15932 ( .A(n15057), .B(n15058), .Z(n15055) );
  AND U15933 ( .A(b[19]), .B(a[26]), .Z(n15054) );
  XOR U15934 ( .A(n15059), .B(n14880), .Z(n14882) );
  XOR U15935 ( .A(n15060), .B(n15061), .Z(n14880) );
  AND U15936 ( .A(n15062), .B(n15063), .Z(n15060) );
  AND U15937 ( .A(a[27]), .B(b[18]), .Z(n15059) );
  XOR U15938 ( .A(n15064), .B(n14885), .Z(n14887) );
  XOR U15939 ( .A(n15065), .B(n15066), .Z(n14885) );
  AND U15940 ( .A(n15067), .B(n15068), .Z(n15065) );
  AND U15941 ( .A(b[17]), .B(a[28]), .Z(n15064) );
  XOR U15942 ( .A(n15069), .B(n14890), .Z(n14892) );
  XOR U15943 ( .A(n15070), .B(n15071), .Z(n14890) );
  AND U15944 ( .A(n15072), .B(n15073), .Z(n15070) );
  AND U15945 ( .A(a[29]), .B(b[16]), .Z(n15069) );
  XOR U15946 ( .A(n15074), .B(n14895), .Z(n14897) );
  XOR U15947 ( .A(n15075), .B(n15076), .Z(n14895) );
  AND U15948 ( .A(n15077), .B(n15078), .Z(n15075) );
  AND U15949 ( .A(b[15]), .B(a[30]), .Z(n15074) );
  XOR U15950 ( .A(n15079), .B(n14900), .Z(n14902) );
  XOR U15951 ( .A(n15080), .B(n15081), .Z(n14900) );
  AND U15952 ( .A(n15082), .B(n15083), .Z(n15080) );
  AND U15953 ( .A(a[31]), .B(b[14]), .Z(n15079) );
  XOR U15954 ( .A(n15084), .B(n14905), .Z(n14907) );
  XOR U15955 ( .A(n15085), .B(n15086), .Z(n14905) );
  AND U15956 ( .A(n15087), .B(n15088), .Z(n15085) );
  AND U15957 ( .A(a[32]), .B(b[13]), .Z(n15084) );
  XOR U15958 ( .A(n15089), .B(n14910), .Z(n14912) );
  XOR U15959 ( .A(n15090), .B(n15091), .Z(n14910) );
  AND U15960 ( .A(n15092), .B(n15093), .Z(n15090) );
  AND U15961 ( .A(a[33]), .B(b[12]), .Z(n15089) );
  XOR U15962 ( .A(n15094), .B(n14915), .Z(n14917) );
  XOR U15963 ( .A(n15095), .B(n15096), .Z(n14915) );
  AND U15964 ( .A(n15097), .B(n15098), .Z(n15095) );
  AND U15965 ( .A(a[34]), .B(b[11]), .Z(n15094) );
  XOR U15966 ( .A(n15099), .B(n14920), .Z(n14922) );
  XOR U15967 ( .A(n15100), .B(n15101), .Z(n14920) );
  AND U15968 ( .A(n15102), .B(n15103), .Z(n15100) );
  AND U15969 ( .A(a[35]), .B(b[10]), .Z(n15099) );
  XOR U15970 ( .A(n15104), .B(n15105), .Z(n14924) );
  AND U15971 ( .A(n15106), .B(n15107), .Z(n15104) );
  XOR U15972 ( .A(n15108), .B(n14929), .Z(n14931) );
  XOR U15973 ( .A(n15109), .B(n15110), .Z(n14929) );
  AND U15974 ( .A(n15111), .B(n15112), .Z(n15109) );
  AND U15975 ( .A(a[36]), .B(b[9]), .Z(n15108) );
  XOR U15976 ( .A(n15114), .B(n15115), .Z(n14934) );
  AND U15977 ( .A(n15116), .B(n15117), .Z(n15114) );
  AND U15978 ( .A(a[38]), .B(b[7]), .Z(n15113) );
  XOR U15979 ( .A(n15119), .B(n15120), .Z(n14939) );
  AND U15980 ( .A(n15121), .B(n15122), .Z(n15119) );
  AND U15981 ( .A(a[39]), .B(b[6]), .Z(n15118) );
  XOR U15982 ( .A(n15124), .B(n15125), .Z(n14944) );
  AND U15983 ( .A(n15126), .B(n15127), .Z(n15124) );
  AND U15984 ( .A(a[40]), .B(b[5]), .Z(n15123) );
  XOR U15985 ( .A(n15129), .B(n15130), .Z(n14949) );
  AND U15986 ( .A(n15131), .B(n15132), .Z(n15129) );
  AND U15987 ( .A(a[41]), .B(b[4]), .Z(n15128) );
  XOR U15988 ( .A(n15134), .B(n15135), .Z(n14954) );
  AND U15989 ( .A(n14968), .B(n14966), .Z(n15134) );
  AND U15990 ( .A(b[2]), .B(a[42]), .Z(n15136) );
  XOR U15991 ( .A(n15131), .B(n15135), .Z(n15137) );
  XOR U15992 ( .A(n15138), .B(n15139), .Z(n15135) );
  NANDN U15993 ( .A(n14970), .B(n14969), .Z(n15139) );
  XOR U15994 ( .A(n15140), .B(n15141), .Z(n14969) );
  NAND U15995 ( .A(a[42]), .B(b[1]), .Z(n15141) );
  XOR U15996 ( .A(n15142), .B(n15143), .Z(n14970) );
  XOR U15997 ( .A(n15140), .B(n15144), .Z(n15143) );
  IV U15998 ( .A(n15138), .Z(n15140) );
  ANDN U15999 ( .B(n5342), .A(n5344), .Z(n15138) );
  NAND U16000 ( .A(a[42]), .B(b[0]), .Z(n5344) );
  XNOR U16001 ( .A(n15145), .B(n15146), .Z(n5342) );
  XOR U16002 ( .A(n15126), .B(n15130), .Z(n15147) );
  XOR U16003 ( .A(n15121), .B(n15125), .Z(n15148) );
  XOR U16004 ( .A(n15116), .B(n15120), .Z(n15149) );
  XOR U16005 ( .A(n15106), .B(n15115), .Z(n15150) );
  XOR U16006 ( .A(n15151), .B(n15105), .Z(n15106) );
  AND U16007 ( .A(b[7]), .B(a[37]), .Z(n15151) );
  XNOR U16008 ( .A(n15105), .B(n15111), .Z(n15152) );
  XNOR U16009 ( .A(n15110), .B(n15102), .Z(n15153) );
  XNOR U16010 ( .A(n15101), .B(n15097), .Z(n15154) );
  XNOR U16011 ( .A(n15096), .B(n15092), .Z(n15155) );
  XNOR U16012 ( .A(n15091), .B(n15087), .Z(n15156) );
  XNOR U16013 ( .A(n15086), .B(n15082), .Z(n15157) );
  XNOR U16014 ( .A(n15081), .B(n15077), .Z(n15158) );
  XNOR U16015 ( .A(n15076), .B(n15072), .Z(n15159) );
  XNOR U16016 ( .A(n15071), .B(n15067), .Z(n15160) );
  XNOR U16017 ( .A(n15066), .B(n15062), .Z(n15161) );
  XNOR U16018 ( .A(n15061), .B(n15057), .Z(n15162) );
  XNOR U16019 ( .A(n15056), .B(n15052), .Z(n15163) );
  XNOR U16020 ( .A(n15051), .B(n15047), .Z(n15164) );
  XNOR U16021 ( .A(n15046), .B(n15042), .Z(n15165) );
  XNOR U16022 ( .A(n15041), .B(n15037), .Z(n15166) );
  XNOR U16023 ( .A(n15036), .B(n15032), .Z(n15167) );
  XNOR U16024 ( .A(n15031), .B(n15027), .Z(n15168) );
  XNOR U16025 ( .A(n15026), .B(n15022), .Z(n15169) );
  XNOR U16026 ( .A(n15021), .B(n15017), .Z(n15170) );
  XNOR U16027 ( .A(n15016), .B(n15012), .Z(n15171) );
  XOR U16028 ( .A(n15011), .B(n15008), .Z(n15172) );
  XOR U16029 ( .A(n15173), .B(n15174), .Z(n15008) );
  XOR U16030 ( .A(n15006), .B(n15175), .Z(n15174) );
  XOR U16031 ( .A(n15176), .B(n15177), .Z(n15175) );
  XOR U16032 ( .A(n15178), .B(n15179), .Z(n15177) );
  NAND U16033 ( .A(a[14]), .B(b[30]), .Z(n15179) );
  AND U16034 ( .A(a[13]), .B(b[31]), .Z(n15178) );
  XOR U16035 ( .A(n15180), .B(n15176), .Z(n15173) );
  XOR U16036 ( .A(n15181), .B(n15182), .Z(n15176) );
  ANDN U16037 ( .B(n15183), .A(n15184), .Z(n15181) );
  AND U16038 ( .A(a[15]), .B(b[29]), .Z(n15180) );
  XOR U16039 ( .A(n15185), .B(n15006), .Z(n15007) );
  XOR U16040 ( .A(n15186), .B(n15187), .Z(n15006) );
  AND U16041 ( .A(n15188), .B(n15189), .Z(n15186) );
  AND U16042 ( .A(a[16]), .B(b[28]), .Z(n15185) );
  XOR U16043 ( .A(n15190), .B(n15011), .Z(n15013) );
  XOR U16044 ( .A(n15191), .B(n15192), .Z(n15011) );
  AND U16045 ( .A(n15193), .B(n15194), .Z(n15191) );
  AND U16046 ( .A(a[17]), .B(b[27]), .Z(n15190) );
  XOR U16047 ( .A(n15195), .B(n15016), .Z(n15018) );
  XOR U16048 ( .A(n15196), .B(n15197), .Z(n15016) );
  AND U16049 ( .A(n15198), .B(n15199), .Z(n15196) );
  AND U16050 ( .A(a[18]), .B(b[26]), .Z(n15195) );
  XOR U16051 ( .A(n15200), .B(n15021), .Z(n15023) );
  XOR U16052 ( .A(n15201), .B(n15202), .Z(n15021) );
  AND U16053 ( .A(n15203), .B(n15204), .Z(n15201) );
  AND U16054 ( .A(a[19]), .B(b[25]), .Z(n15200) );
  XOR U16055 ( .A(n15205), .B(n15026), .Z(n15028) );
  XOR U16056 ( .A(n15206), .B(n15207), .Z(n15026) );
  AND U16057 ( .A(n15208), .B(n15209), .Z(n15206) );
  AND U16058 ( .A(a[20]), .B(b[24]), .Z(n15205) );
  XOR U16059 ( .A(n15210), .B(n15031), .Z(n15033) );
  XOR U16060 ( .A(n15211), .B(n15212), .Z(n15031) );
  AND U16061 ( .A(n15213), .B(n15214), .Z(n15211) );
  AND U16062 ( .A(a[21]), .B(b[23]), .Z(n15210) );
  XOR U16063 ( .A(n15215), .B(n15036), .Z(n15038) );
  XOR U16064 ( .A(n15216), .B(n15217), .Z(n15036) );
  AND U16065 ( .A(n15218), .B(n15219), .Z(n15216) );
  AND U16066 ( .A(b[22]), .B(a[22]), .Z(n15215) );
  XOR U16067 ( .A(n15220), .B(n15041), .Z(n15043) );
  XOR U16068 ( .A(n15221), .B(n15222), .Z(n15041) );
  AND U16069 ( .A(n15223), .B(n15224), .Z(n15221) );
  AND U16070 ( .A(a[23]), .B(b[21]), .Z(n15220) );
  XOR U16071 ( .A(n15225), .B(n15046), .Z(n15048) );
  XOR U16072 ( .A(n15226), .B(n15227), .Z(n15046) );
  AND U16073 ( .A(n15228), .B(n15229), .Z(n15226) );
  AND U16074 ( .A(b[20]), .B(a[24]), .Z(n15225) );
  XOR U16075 ( .A(n15230), .B(n15051), .Z(n15053) );
  XOR U16076 ( .A(n15231), .B(n15232), .Z(n15051) );
  AND U16077 ( .A(n15233), .B(n15234), .Z(n15231) );
  AND U16078 ( .A(a[25]), .B(b[19]), .Z(n15230) );
  XOR U16079 ( .A(n15235), .B(n15056), .Z(n15058) );
  XOR U16080 ( .A(n15236), .B(n15237), .Z(n15056) );
  AND U16081 ( .A(n15238), .B(n15239), .Z(n15236) );
  AND U16082 ( .A(b[18]), .B(a[26]), .Z(n15235) );
  XOR U16083 ( .A(n15240), .B(n15061), .Z(n15063) );
  XOR U16084 ( .A(n15241), .B(n15242), .Z(n15061) );
  AND U16085 ( .A(n15243), .B(n15244), .Z(n15241) );
  AND U16086 ( .A(a[27]), .B(b[17]), .Z(n15240) );
  XOR U16087 ( .A(n15245), .B(n15066), .Z(n15068) );
  XOR U16088 ( .A(n15246), .B(n15247), .Z(n15066) );
  AND U16089 ( .A(n15248), .B(n15249), .Z(n15246) );
  AND U16090 ( .A(b[16]), .B(a[28]), .Z(n15245) );
  XOR U16091 ( .A(n15250), .B(n15071), .Z(n15073) );
  XOR U16092 ( .A(n15251), .B(n15252), .Z(n15071) );
  AND U16093 ( .A(n15253), .B(n15254), .Z(n15251) );
  AND U16094 ( .A(a[29]), .B(b[15]), .Z(n15250) );
  XOR U16095 ( .A(n15255), .B(n15076), .Z(n15078) );
  XOR U16096 ( .A(n15256), .B(n15257), .Z(n15076) );
  AND U16097 ( .A(n15258), .B(n15259), .Z(n15256) );
  AND U16098 ( .A(b[14]), .B(a[30]), .Z(n15255) );
  XOR U16099 ( .A(n15260), .B(n15081), .Z(n15083) );
  XOR U16100 ( .A(n15261), .B(n15262), .Z(n15081) );
  AND U16101 ( .A(n15263), .B(n15264), .Z(n15261) );
  AND U16102 ( .A(a[31]), .B(b[13]), .Z(n15260) );
  XOR U16103 ( .A(n15265), .B(n15086), .Z(n15088) );
  XOR U16104 ( .A(n15266), .B(n15267), .Z(n15086) );
  AND U16105 ( .A(n15268), .B(n15269), .Z(n15266) );
  AND U16106 ( .A(a[32]), .B(b[12]), .Z(n15265) );
  XOR U16107 ( .A(n15270), .B(n15091), .Z(n15093) );
  XOR U16108 ( .A(n15271), .B(n15272), .Z(n15091) );
  AND U16109 ( .A(n15273), .B(n15274), .Z(n15271) );
  AND U16110 ( .A(a[33]), .B(b[11]), .Z(n15270) );
  XOR U16111 ( .A(n15275), .B(n15096), .Z(n15098) );
  XOR U16112 ( .A(n15276), .B(n15277), .Z(n15096) );
  AND U16113 ( .A(n15278), .B(n15279), .Z(n15276) );
  AND U16114 ( .A(a[34]), .B(b[10]), .Z(n15275) );
  XOR U16115 ( .A(n15280), .B(n15101), .Z(n15103) );
  XOR U16116 ( .A(n15281), .B(n15282), .Z(n15101) );
  AND U16117 ( .A(n15283), .B(n15284), .Z(n15281) );
  AND U16118 ( .A(a[35]), .B(b[9]), .Z(n15280) );
  XOR U16119 ( .A(n15285), .B(n15286), .Z(n15105) );
  AND U16120 ( .A(n15287), .B(n15288), .Z(n15285) );
  XOR U16121 ( .A(n15289), .B(n15110), .Z(n15112) );
  XOR U16122 ( .A(n15290), .B(n15291), .Z(n15110) );
  AND U16123 ( .A(n15292), .B(n15293), .Z(n15290) );
  AND U16124 ( .A(a[36]), .B(b[8]), .Z(n15289) );
  XOR U16125 ( .A(n15295), .B(n15296), .Z(n15115) );
  AND U16126 ( .A(n15297), .B(n15298), .Z(n15295) );
  AND U16127 ( .A(a[38]), .B(b[6]), .Z(n15294) );
  XOR U16128 ( .A(n15300), .B(n15301), .Z(n15120) );
  AND U16129 ( .A(n15302), .B(n15303), .Z(n15300) );
  AND U16130 ( .A(a[39]), .B(b[5]), .Z(n15299) );
  XOR U16131 ( .A(n15305), .B(n15306), .Z(n15125) );
  AND U16132 ( .A(n15307), .B(n15308), .Z(n15305) );
  AND U16133 ( .A(a[40]), .B(b[4]), .Z(n15304) );
  XOR U16134 ( .A(n15310), .B(n15311), .Z(n15130) );
  AND U16135 ( .A(n15144), .B(n15142), .Z(n15310) );
  AND U16136 ( .A(b[2]), .B(a[41]), .Z(n15312) );
  XOR U16137 ( .A(n15307), .B(n15311), .Z(n15313) );
  XOR U16138 ( .A(n15314), .B(n15315), .Z(n15311) );
  NANDN U16139 ( .A(n15146), .B(n15145), .Z(n15315) );
  XOR U16140 ( .A(n15316), .B(n15317), .Z(n15145) );
  NAND U16141 ( .A(a[41]), .B(b[1]), .Z(n15317) );
  XOR U16142 ( .A(n15318), .B(n15319), .Z(n15146) );
  XOR U16143 ( .A(n15316), .B(n15320), .Z(n15319) );
  IV U16144 ( .A(n15314), .Z(n15316) );
  ANDN U16145 ( .B(n5347), .A(n5349), .Z(n15314) );
  NAND U16146 ( .A(a[41]), .B(b[0]), .Z(n5349) );
  XNOR U16147 ( .A(n15321), .B(n15322), .Z(n5347) );
  XOR U16148 ( .A(n15302), .B(n15306), .Z(n15323) );
  XOR U16149 ( .A(n15297), .B(n15301), .Z(n15324) );
  XOR U16150 ( .A(n15287), .B(n15296), .Z(n15325) );
  XOR U16151 ( .A(n15326), .B(n15286), .Z(n15287) );
  AND U16152 ( .A(b[6]), .B(a[37]), .Z(n15326) );
  XNOR U16153 ( .A(n15286), .B(n15292), .Z(n15327) );
  XNOR U16154 ( .A(n15291), .B(n15283), .Z(n15328) );
  XNOR U16155 ( .A(n15282), .B(n15278), .Z(n15329) );
  XNOR U16156 ( .A(n15277), .B(n15273), .Z(n15330) );
  XNOR U16157 ( .A(n15272), .B(n15268), .Z(n15331) );
  XNOR U16158 ( .A(n15267), .B(n15263), .Z(n15332) );
  XNOR U16159 ( .A(n15262), .B(n15258), .Z(n15333) );
  XNOR U16160 ( .A(n15257), .B(n15253), .Z(n15334) );
  XNOR U16161 ( .A(n15252), .B(n15248), .Z(n15335) );
  XNOR U16162 ( .A(n15247), .B(n15243), .Z(n15336) );
  XNOR U16163 ( .A(n15242), .B(n15238), .Z(n15337) );
  XNOR U16164 ( .A(n15237), .B(n15233), .Z(n15338) );
  XNOR U16165 ( .A(n15232), .B(n15228), .Z(n15339) );
  XNOR U16166 ( .A(n15227), .B(n15223), .Z(n15340) );
  XNOR U16167 ( .A(n15222), .B(n15218), .Z(n15341) );
  XNOR U16168 ( .A(n15217), .B(n15213), .Z(n15342) );
  XNOR U16169 ( .A(n15212), .B(n15208), .Z(n15343) );
  XNOR U16170 ( .A(n15207), .B(n15203), .Z(n15344) );
  XNOR U16171 ( .A(n15202), .B(n15198), .Z(n15345) );
  XNOR U16172 ( .A(n15197), .B(n15193), .Z(n15346) );
  XNOR U16173 ( .A(n15192), .B(n15188), .Z(n15347) );
  XOR U16174 ( .A(n15187), .B(n15184), .Z(n15348) );
  XOR U16175 ( .A(n15349), .B(n15350), .Z(n15184) );
  XOR U16176 ( .A(n15182), .B(n15351), .Z(n15350) );
  XOR U16177 ( .A(n15352), .B(n15353), .Z(n15351) );
  XOR U16178 ( .A(n15354), .B(n15355), .Z(n15353) );
  NAND U16179 ( .A(a[13]), .B(b[30]), .Z(n15355) );
  AND U16180 ( .A(a[12]), .B(b[31]), .Z(n15354) );
  XOR U16181 ( .A(n15356), .B(n15352), .Z(n15349) );
  XOR U16182 ( .A(n15357), .B(n15358), .Z(n15352) );
  ANDN U16183 ( .B(n15359), .A(n15360), .Z(n15357) );
  AND U16184 ( .A(a[14]), .B(b[29]), .Z(n15356) );
  XOR U16185 ( .A(n15361), .B(n15182), .Z(n15183) );
  XOR U16186 ( .A(n15362), .B(n15363), .Z(n15182) );
  AND U16187 ( .A(n15364), .B(n15365), .Z(n15362) );
  AND U16188 ( .A(a[15]), .B(b[28]), .Z(n15361) );
  XOR U16189 ( .A(n15366), .B(n15187), .Z(n15189) );
  XOR U16190 ( .A(n15367), .B(n15368), .Z(n15187) );
  AND U16191 ( .A(n15369), .B(n15370), .Z(n15367) );
  AND U16192 ( .A(a[16]), .B(b[27]), .Z(n15366) );
  XOR U16193 ( .A(n15371), .B(n15192), .Z(n15194) );
  XOR U16194 ( .A(n15372), .B(n15373), .Z(n15192) );
  AND U16195 ( .A(n15374), .B(n15375), .Z(n15372) );
  AND U16196 ( .A(a[17]), .B(b[26]), .Z(n15371) );
  XOR U16197 ( .A(n15376), .B(n15197), .Z(n15199) );
  XOR U16198 ( .A(n15377), .B(n15378), .Z(n15197) );
  AND U16199 ( .A(n15379), .B(n15380), .Z(n15377) );
  AND U16200 ( .A(a[18]), .B(b[25]), .Z(n15376) );
  XOR U16201 ( .A(n15381), .B(n15202), .Z(n15204) );
  XOR U16202 ( .A(n15382), .B(n15383), .Z(n15202) );
  AND U16203 ( .A(n15384), .B(n15385), .Z(n15382) );
  AND U16204 ( .A(a[19]), .B(b[24]), .Z(n15381) );
  XOR U16205 ( .A(n15386), .B(n15207), .Z(n15209) );
  XOR U16206 ( .A(n15387), .B(n15388), .Z(n15207) );
  AND U16207 ( .A(n15389), .B(n15390), .Z(n15387) );
  AND U16208 ( .A(a[20]), .B(b[23]), .Z(n15386) );
  XOR U16209 ( .A(n15391), .B(n15212), .Z(n15214) );
  XOR U16210 ( .A(n15392), .B(n15393), .Z(n15212) );
  AND U16211 ( .A(n15394), .B(n15395), .Z(n15392) );
  AND U16212 ( .A(a[21]), .B(b[22]), .Z(n15391) );
  XOR U16213 ( .A(n15396), .B(n15217), .Z(n15219) );
  XOR U16214 ( .A(n15397), .B(n15398), .Z(n15217) );
  AND U16215 ( .A(n15399), .B(n15400), .Z(n15397) );
  AND U16216 ( .A(b[21]), .B(a[22]), .Z(n15396) );
  XOR U16217 ( .A(n15401), .B(n15222), .Z(n15224) );
  XOR U16218 ( .A(n15402), .B(n15403), .Z(n15222) );
  AND U16219 ( .A(n15404), .B(n15405), .Z(n15402) );
  AND U16220 ( .A(a[23]), .B(b[20]), .Z(n15401) );
  XOR U16221 ( .A(n15406), .B(n15227), .Z(n15229) );
  XOR U16222 ( .A(n15407), .B(n15408), .Z(n15227) );
  AND U16223 ( .A(n15409), .B(n15410), .Z(n15407) );
  AND U16224 ( .A(b[19]), .B(a[24]), .Z(n15406) );
  XOR U16225 ( .A(n15411), .B(n15232), .Z(n15234) );
  XOR U16226 ( .A(n15412), .B(n15413), .Z(n15232) );
  AND U16227 ( .A(n15414), .B(n15415), .Z(n15412) );
  AND U16228 ( .A(a[25]), .B(b[18]), .Z(n15411) );
  XOR U16229 ( .A(n15416), .B(n15237), .Z(n15239) );
  XOR U16230 ( .A(n15417), .B(n15418), .Z(n15237) );
  AND U16231 ( .A(n15419), .B(n15420), .Z(n15417) );
  AND U16232 ( .A(b[17]), .B(a[26]), .Z(n15416) );
  XOR U16233 ( .A(n15421), .B(n15242), .Z(n15244) );
  XOR U16234 ( .A(n15422), .B(n15423), .Z(n15242) );
  AND U16235 ( .A(n15424), .B(n15425), .Z(n15422) );
  AND U16236 ( .A(a[27]), .B(b[16]), .Z(n15421) );
  XOR U16237 ( .A(n15426), .B(n15247), .Z(n15249) );
  XOR U16238 ( .A(n15427), .B(n15428), .Z(n15247) );
  AND U16239 ( .A(n15429), .B(n15430), .Z(n15427) );
  AND U16240 ( .A(b[15]), .B(a[28]), .Z(n15426) );
  XOR U16241 ( .A(n15431), .B(n15252), .Z(n15254) );
  XOR U16242 ( .A(n15432), .B(n15433), .Z(n15252) );
  AND U16243 ( .A(n15434), .B(n15435), .Z(n15432) );
  AND U16244 ( .A(a[29]), .B(b[14]), .Z(n15431) );
  XOR U16245 ( .A(n15436), .B(n15257), .Z(n15259) );
  XOR U16246 ( .A(n15437), .B(n15438), .Z(n15257) );
  AND U16247 ( .A(n15439), .B(n15440), .Z(n15437) );
  AND U16248 ( .A(b[13]), .B(a[30]), .Z(n15436) );
  XOR U16249 ( .A(n15441), .B(n15262), .Z(n15264) );
  XOR U16250 ( .A(n15442), .B(n15443), .Z(n15262) );
  AND U16251 ( .A(n15444), .B(n15445), .Z(n15442) );
  AND U16252 ( .A(a[31]), .B(b[12]), .Z(n15441) );
  XOR U16253 ( .A(n15446), .B(n15267), .Z(n15269) );
  XOR U16254 ( .A(n15447), .B(n15448), .Z(n15267) );
  AND U16255 ( .A(n15449), .B(n15450), .Z(n15447) );
  AND U16256 ( .A(a[32]), .B(b[11]), .Z(n15446) );
  XOR U16257 ( .A(n15451), .B(n15272), .Z(n15274) );
  XOR U16258 ( .A(n15452), .B(n15453), .Z(n15272) );
  AND U16259 ( .A(n15454), .B(n15455), .Z(n15452) );
  AND U16260 ( .A(a[33]), .B(b[10]), .Z(n15451) );
  XOR U16261 ( .A(n15456), .B(n15277), .Z(n15279) );
  XOR U16262 ( .A(n15457), .B(n15458), .Z(n15277) );
  AND U16263 ( .A(n15459), .B(n15460), .Z(n15457) );
  AND U16264 ( .A(a[34]), .B(b[9]), .Z(n15456) );
  XOR U16265 ( .A(n15461), .B(n15282), .Z(n15284) );
  XOR U16266 ( .A(n15462), .B(n15463), .Z(n15282) );
  AND U16267 ( .A(n15464), .B(n15465), .Z(n15462) );
  AND U16268 ( .A(a[35]), .B(b[8]), .Z(n15461) );
  XOR U16269 ( .A(n15466), .B(n15467), .Z(n15286) );
  AND U16270 ( .A(n15468), .B(n15469), .Z(n15466) );
  XOR U16271 ( .A(n15470), .B(n15291), .Z(n15293) );
  XOR U16272 ( .A(n15471), .B(n15472), .Z(n15291) );
  AND U16273 ( .A(n15473), .B(n15474), .Z(n15471) );
  AND U16274 ( .A(a[36]), .B(b[7]), .Z(n15470) );
  XOR U16275 ( .A(n15476), .B(n15477), .Z(n15296) );
  AND U16276 ( .A(n15478), .B(n15479), .Z(n15476) );
  AND U16277 ( .A(a[38]), .B(b[5]), .Z(n15475) );
  XOR U16278 ( .A(n15481), .B(n15482), .Z(n15301) );
  AND U16279 ( .A(n15483), .B(n15484), .Z(n15481) );
  AND U16280 ( .A(a[39]), .B(b[4]), .Z(n15480) );
  XOR U16281 ( .A(n15486), .B(n15487), .Z(n15306) );
  AND U16282 ( .A(n15320), .B(n15318), .Z(n15486) );
  AND U16283 ( .A(b[2]), .B(a[40]), .Z(n15488) );
  XOR U16284 ( .A(n15483), .B(n15487), .Z(n15489) );
  XOR U16285 ( .A(n15490), .B(n15491), .Z(n15487) );
  NANDN U16286 ( .A(n15322), .B(n15321), .Z(n15491) );
  XOR U16287 ( .A(n15492), .B(n15493), .Z(n15321) );
  NAND U16288 ( .A(a[40]), .B(b[1]), .Z(n15493) );
  XOR U16289 ( .A(n15494), .B(n15495), .Z(n15322) );
  XOR U16290 ( .A(n15492), .B(n15496), .Z(n15495) );
  IV U16291 ( .A(n15490), .Z(n15492) );
  ANDN U16292 ( .B(n5352), .A(n5354), .Z(n15490) );
  NAND U16293 ( .A(a[40]), .B(b[0]), .Z(n5354) );
  XNOR U16294 ( .A(n15497), .B(n15498), .Z(n5352) );
  XOR U16295 ( .A(n15478), .B(n15482), .Z(n15499) );
  XOR U16296 ( .A(n15468), .B(n15477), .Z(n15500) );
  XOR U16297 ( .A(n15501), .B(n15467), .Z(n15468) );
  AND U16298 ( .A(b[5]), .B(a[37]), .Z(n15501) );
  XNOR U16299 ( .A(n15467), .B(n15473), .Z(n15502) );
  XNOR U16300 ( .A(n15472), .B(n15464), .Z(n15503) );
  XNOR U16301 ( .A(n15463), .B(n15459), .Z(n15504) );
  XNOR U16302 ( .A(n15458), .B(n15454), .Z(n15505) );
  XNOR U16303 ( .A(n15453), .B(n15449), .Z(n15506) );
  XNOR U16304 ( .A(n15448), .B(n15444), .Z(n15507) );
  XNOR U16305 ( .A(n15443), .B(n15439), .Z(n15508) );
  XNOR U16306 ( .A(n15438), .B(n15434), .Z(n15509) );
  XNOR U16307 ( .A(n15433), .B(n15429), .Z(n15510) );
  XNOR U16308 ( .A(n15428), .B(n15424), .Z(n15511) );
  XNOR U16309 ( .A(n15423), .B(n15419), .Z(n15512) );
  XNOR U16310 ( .A(n15418), .B(n15414), .Z(n15513) );
  XNOR U16311 ( .A(n15413), .B(n15409), .Z(n15514) );
  XNOR U16312 ( .A(n15408), .B(n15404), .Z(n15515) );
  XNOR U16313 ( .A(n15403), .B(n15399), .Z(n15516) );
  XNOR U16314 ( .A(n15398), .B(n15394), .Z(n15517) );
  XNOR U16315 ( .A(n15393), .B(n15389), .Z(n15518) );
  XNOR U16316 ( .A(n15388), .B(n15384), .Z(n15519) );
  XNOR U16317 ( .A(n15383), .B(n15379), .Z(n15520) );
  XNOR U16318 ( .A(n15378), .B(n15374), .Z(n15521) );
  XNOR U16319 ( .A(n15373), .B(n15369), .Z(n15522) );
  XNOR U16320 ( .A(n15368), .B(n15364), .Z(n15523) );
  XOR U16321 ( .A(n15363), .B(n15360), .Z(n15524) );
  XOR U16322 ( .A(n15525), .B(n15526), .Z(n15360) );
  XOR U16323 ( .A(n15358), .B(n15527), .Z(n15526) );
  XOR U16324 ( .A(n15528), .B(n15529), .Z(n15527) );
  XOR U16325 ( .A(n15530), .B(n15531), .Z(n15529) );
  NAND U16326 ( .A(a[12]), .B(b[30]), .Z(n15531) );
  AND U16327 ( .A(a[11]), .B(b[31]), .Z(n15530) );
  XOR U16328 ( .A(n15532), .B(n15528), .Z(n15525) );
  XOR U16329 ( .A(n15533), .B(n15534), .Z(n15528) );
  ANDN U16330 ( .B(n15535), .A(n15536), .Z(n15533) );
  AND U16331 ( .A(a[13]), .B(b[29]), .Z(n15532) );
  XOR U16332 ( .A(n15537), .B(n15358), .Z(n15359) );
  XOR U16333 ( .A(n15538), .B(n15539), .Z(n15358) );
  AND U16334 ( .A(n15540), .B(n15541), .Z(n15538) );
  AND U16335 ( .A(a[14]), .B(b[28]), .Z(n15537) );
  XOR U16336 ( .A(n15542), .B(n15363), .Z(n15365) );
  XOR U16337 ( .A(n15543), .B(n15544), .Z(n15363) );
  AND U16338 ( .A(n15545), .B(n15546), .Z(n15543) );
  AND U16339 ( .A(a[15]), .B(b[27]), .Z(n15542) );
  XOR U16340 ( .A(n15547), .B(n15368), .Z(n15370) );
  XOR U16341 ( .A(n15548), .B(n15549), .Z(n15368) );
  AND U16342 ( .A(n15550), .B(n15551), .Z(n15548) );
  AND U16343 ( .A(a[16]), .B(b[26]), .Z(n15547) );
  XOR U16344 ( .A(n15552), .B(n15373), .Z(n15375) );
  XOR U16345 ( .A(n15553), .B(n15554), .Z(n15373) );
  AND U16346 ( .A(n15555), .B(n15556), .Z(n15553) );
  AND U16347 ( .A(a[17]), .B(b[25]), .Z(n15552) );
  XOR U16348 ( .A(n15557), .B(n15378), .Z(n15380) );
  XOR U16349 ( .A(n15558), .B(n15559), .Z(n15378) );
  AND U16350 ( .A(n15560), .B(n15561), .Z(n15558) );
  AND U16351 ( .A(a[18]), .B(b[24]), .Z(n15557) );
  XOR U16352 ( .A(n15562), .B(n15383), .Z(n15385) );
  XOR U16353 ( .A(n15563), .B(n15564), .Z(n15383) );
  AND U16354 ( .A(n15565), .B(n15566), .Z(n15563) );
  AND U16355 ( .A(a[19]), .B(b[23]), .Z(n15562) );
  XOR U16356 ( .A(n15567), .B(n15388), .Z(n15390) );
  XOR U16357 ( .A(n15568), .B(n15569), .Z(n15388) );
  AND U16358 ( .A(n15570), .B(n15571), .Z(n15568) );
  AND U16359 ( .A(a[20]), .B(b[22]), .Z(n15567) );
  XOR U16360 ( .A(n15572), .B(n15393), .Z(n15395) );
  XOR U16361 ( .A(n15573), .B(n15574), .Z(n15393) );
  AND U16362 ( .A(n15575), .B(n15576), .Z(n15573) );
  AND U16363 ( .A(a[21]), .B(b[21]), .Z(n15572) );
  XOR U16364 ( .A(n15577), .B(n15398), .Z(n15400) );
  XOR U16365 ( .A(n15578), .B(n15579), .Z(n15398) );
  AND U16366 ( .A(n15580), .B(n15581), .Z(n15578) );
  AND U16367 ( .A(b[20]), .B(a[22]), .Z(n15577) );
  XOR U16368 ( .A(n15582), .B(n15403), .Z(n15405) );
  XOR U16369 ( .A(n15583), .B(n15584), .Z(n15403) );
  AND U16370 ( .A(n15585), .B(n15586), .Z(n15583) );
  AND U16371 ( .A(a[23]), .B(b[19]), .Z(n15582) );
  XOR U16372 ( .A(n15587), .B(n15408), .Z(n15410) );
  XOR U16373 ( .A(n15588), .B(n15589), .Z(n15408) );
  AND U16374 ( .A(n15590), .B(n15591), .Z(n15588) );
  AND U16375 ( .A(b[18]), .B(a[24]), .Z(n15587) );
  XOR U16376 ( .A(n15592), .B(n15413), .Z(n15415) );
  XOR U16377 ( .A(n15593), .B(n15594), .Z(n15413) );
  AND U16378 ( .A(n15595), .B(n15596), .Z(n15593) );
  AND U16379 ( .A(a[25]), .B(b[17]), .Z(n15592) );
  XOR U16380 ( .A(n15597), .B(n15418), .Z(n15420) );
  XOR U16381 ( .A(n15598), .B(n15599), .Z(n15418) );
  AND U16382 ( .A(n15600), .B(n15601), .Z(n15598) );
  AND U16383 ( .A(b[16]), .B(a[26]), .Z(n15597) );
  XOR U16384 ( .A(n15602), .B(n15423), .Z(n15425) );
  XOR U16385 ( .A(n15603), .B(n15604), .Z(n15423) );
  AND U16386 ( .A(n15605), .B(n15606), .Z(n15603) );
  AND U16387 ( .A(a[27]), .B(b[15]), .Z(n15602) );
  XOR U16388 ( .A(n15607), .B(n15428), .Z(n15430) );
  XOR U16389 ( .A(n15608), .B(n15609), .Z(n15428) );
  AND U16390 ( .A(n15610), .B(n15611), .Z(n15608) );
  AND U16391 ( .A(b[14]), .B(a[28]), .Z(n15607) );
  XOR U16392 ( .A(n15612), .B(n15433), .Z(n15435) );
  XOR U16393 ( .A(n15613), .B(n15614), .Z(n15433) );
  AND U16394 ( .A(n15615), .B(n15616), .Z(n15613) );
  AND U16395 ( .A(a[29]), .B(b[13]), .Z(n15612) );
  XOR U16396 ( .A(n15617), .B(n15438), .Z(n15440) );
  XOR U16397 ( .A(n15618), .B(n15619), .Z(n15438) );
  AND U16398 ( .A(n15620), .B(n15621), .Z(n15618) );
  AND U16399 ( .A(b[12]), .B(a[30]), .Z(n15617) );
  XOR U16400 ( .A(n15622), .B(n15443), .Z(n15445) );
  XOR U16401 ( .A(n15623), .B(n15624), .Z(n15443) );
  AND U16402 ( .A(n15625), .B(n15626), .Z(n15623) );
  AND U16403 ( .A(a[31]), .B(b[11]), .Z(n15622) );
  XOR U16404 ( .A(n15627), .B(n15448), .Z(n15450) );
  XOR U16405 ( .A(n15628), .B(n15629), .Z(n15448) );
  AND U16406 ( .A(n15630), .B(n15631), .Z(n15628) );
  AND U16407 ( .A(a[32]), .B(b[10]), .Z(n15627) );
  XOR U16408 ( .A(n15632), .B(n15453), .Z(n15455) );
  XOR U16409 ( .A(n15633), .B(n15634), .Z(n15453) );
  AND U16410 ( .A(n15635), .B(n15636), .Z(n15633) );
  AND U16411 ( .A(a[33]), .B(b[9]), .Z(n15632) );
  XOR U16412 ( .A(n15637), .B(n15458), .Z(n15460) );
  XOR U16413 ( .A(n15638), .B(n15639), .Z(n15458) );
  AND U16414 ( .A(n15640), .B(n15641), .Z(n15638) );
  AND U16415 ( .A(a[34]), .B(b[8]), .Z(n15637) );
  XOR U16416 ( .A(n15642), .B(n15463), .Z(n15465) );
  XOR U16417 ( .A(n15643), .B(n15644), .Z(n15463) );
  AND U16418 ( .A(n15645), .B(n15646), .Z(n15643) );
  AND U16419 ( .A(a[35]), .B(b[7]), .Z(n15642) );
  XOR U16420 ( .A(n15647), .B(n15648), .Z(n15467) );
  AND U16421 ( .A(n15649), .B(n15650), .Z(n15647) );
  XOR U16422 ( .A(n15651), .B(n15472), .Z(n15474) );
  XOR U16423 ( .A(n15652), .B(n15653), .Z(n15472) );
  AND U16424 ( .A(n15654), .B(n15655), .Z(n15652) );
  AND U16425 ( .A(a[36]), .B(b[6]), .Z(n15651) );
  XOR U16426 ( .A(n15657), .B(n15658), .Z(n15477) );
  AND U16427 ( .A(n15659), .B(n15660), .Z(n15657) );
  AND U16428 ( .A(a[38]), .B(b[4]), .Z(n15656) );
  XOR U16429 ( .A(n15662), .B(n15663), .Z(n15482) );
  AND U16430 ( .A(n15496), .B(n15494), .Z(n15662) );
  AND U16431 ( .A(b[2]), .B(a[39]), .Z(n15664) );
  XOR U16432 ( .A(n15659), .B(n15663), .Z(n15665) );
  XOR U16433 ( .A(n15666), .B(n15667), .Z(n15663) );
  NANDN U16434 ( .A(n15498), .B(n15497), .Z(n15667) );
  XOR U16435 ( .A(n15668), .B(n15669), .Z(n15497) );
  NAND U16436 ( .A(a[39]), .B(b[1]), .Z(n15669) );
  XOR U16437 ( .A(n15670), .B(n15671), .Z(n15498) );
  XOR U16438 ( .A(n15668), .B(n15672), .Z(n15671) );
  IV U16439 ( .A(n15666), .Z(n15668) );
  ANDN U16440 ( .B(n5357), .A(n5359), .Z(n15666) );
  NAND U16441 ( .A(a[39]), .B(b[0]), .Z(n5359) );
  XNOR U16442 ( .A(n15673), .B(n15674), .Z(n5357) );
  XOR U16443 ( .A(n15649), .B(n15658), .Z(n15675) );
  XOR U16444 ( .A(n15676), .B(n15648), .Z(n15649) );
  AND U16445 ( .A(b[4]), .B(a[37]), .Z(n15676) );
  XNOR U16446 ( .A(n15648), .B(n15654), .Z(n15677) );
  XNOR U16447 ( .A(n15653), .B(n15645), .Z(n15678) );
  XNOR U16448 ( .A(n15644), .B(n15640), .Z(n15679) );
  XNOR U16449 ( .A(n15639), .B(n15635), .Z(n15680) );
  XNOR U16450 ( .A(n15634), .B(n15630), .Z(n15681) );
  XNOR U16451 ( .A(n15629), .B(n15625), .Z(n15682) );
  XNOR U16452 ( .A(n15624), .B(n15620), .Z(n15683) );
  XNOR U16453 ( .A(n15619), .B(n15615), .Z(n15684) );
  XNOR U16454 ( .A(n15614), .B(n15610), .Z(n15685) );
  XNOR U16455 ( .A(n15609), .B(n15605), .Z(n15686) );
  XNOR U16456 ( .A(n15604), .B(n15600), .Z(n15687) );
  XNOR U16457 ( .A(n15599), .B(n15595), .Z(n15688) );
  XNOR U16458 ( .A(n15594), .B(n15590), .Z(n15689) );
  XNOR U16459 ( .A(n15589), .B(n15585), .Z(n15690) );
  XNOR U16460 ( .A(n15584), .B(n15580), .Z(n15691) );
  XNOR U16461 ( .A(n15579), .B(n15575), .Z(n15692) );
  XNOR U16462 ( .A(n15574), .B(n15570), .Z(n15693) );
  XNOR U16463 ( .A(n15569), .B(n15565), .Z(n15694) );
  XNOR U16464 ( .A(n15564), .B(n15560), .Z(n15695) );
  XNOR U16465 ( .A(n15559), .B(n15555), .Z(n15696) );
  XNOR U16466 ( .A(n15554), .B(n15550), .Z(n15697) );
  XNOR U16467 ( .A(n15549), .B(n15545), .Z(n15698) );
  XNOR U16468 ( .A(n15544), .B(n15540), .Z(n15699) );
  XOR U16469 ( .A(n15539), .B(n15536), .Z(n15700) );
  XOR U16470 ( .A(n15701), .B(n15702), .Z(n15536) );
  XOR U16471 ( .A(n15534), .B(n15703), .Z(n15702) );
  XOR U16472 ( .A(n15704), .B(n15705), .Z(n15703) );
  XOR U16473 ( .A(n15706), .B(n15707), .Z(n15705) );
  NAND U16474 ( .A(a[11]), .B(b[30]), .Z(n15707) );
  AND U16475 ( .A(a[10]), .B(b[31]), .Z(n15706) );
  XOR U16476 ( .A(n15708), .B(n15704), .Z(n15701) );
  XOR U16477 ( .A(n15709), .B(n15710), .Z(n15704) );
  ANDN U16478 ( .B(n15711), .A(n15712), .Z(n15709) );
  AND U16479 ( .A(a[12]), .B(b[29]), .Z(n15708) );
  XOR U16480 ( .A(n15713), .B(n15534), .Z(n15535) );
  XOR U16481 ( .A(n15714), .B(n15715), .Z(n15534) );
  AND U16482 ( .A(n15716), .B(n15717), .Z(n15714) );
  AND U16483 ( .A(a[13]), .B(b[28]), .Z(n15713) );
  XOR U16484 ( .A(n15718), .B(n15539), .Z(n15541) );
  XOR U16485 ( .A(n15719), .B(n15720), .Z(n15539) );
  AND U16486 ( .A(n15721), .B(n15722), .Z(n15719) );
  AND U16487 ( .A(a[14]), .B(b[27]), .Z(n15718) );
  XOR U16488 ( .A(n15723), .B(n15544), .Z(n15546) );
  XOR U16489 ( .A(n15724), .B(n15725), .Z(n15544) );
  AND U16490 ( .A(n15726), .B(n15727), .Z(n15724) );
  AND U16491 ( .A(a[15]), .B(b[26]), .Z(n15723) );
  XOR U16492 ( .A(n15728), .B(n15549), .Z(n15551) );
  XOR U16493 ( .A(n15729), .B(n15730), .Z(n15549) );
  AND U16494 ( .A(n15731), .B(n15732), .Z(n15729) );
  AND U16495 ( .A(a[16]), .B(b[25]), .Z(n15728) );
  XOR U16496 ( .A(n15733), .B(n15554), .Z(n15556) );
  XOR U16497 ( .A(n15734), .B(n15735), .Z(n15554) );
  AND U16498 ( .A(n15736), .B(n15737), .Z(n15734) );
  AND U16499 ( .A(a[17]), .B(b[24]), .Z(n15733) );
  XOR U16500 ( .A(n15738), .B(n15559), .Z(n15561) );
  XOR U16501 ( .A(n15739), .B(n15740), .Z(n15559) );
  AND U16502 ( .A(n15741), .B(n15742), .Z(n15739) );
  AND U16503 ( .A(a[18]), .B(b[23]), .Z(n15738) );
  XOR U16504 ( .A(n15743), .B(n15564), .Z(n15566) );
  XOR U16505 ( .A(n15744), .B(n15745), .Z(n15564) );
  AND U16506 ( .A(n15746), .B(n15747), .Z(n15744) );
  AND U16507 ( .A(a[19]), .B(b[22]), .Z(n15743) );
  XOR U16508 ( .A(n15748), .B(n15569), .Z(n15571) );
  XOR U16509 ( .A(n15749), .B(n15750), .Z(n15569) );
  AND U16510 ( .A(n15751), .B(n15752), .Z(n15749) );
  AND U16511 ( .A(a[20]), .B(b[21]), .Z(n15748) );
  XOR U16512 ( .A(n15753), .B(n15574), .Z(n15576) );
  XOR U16513 ( .A(n15754), .B(n15755), .Z(n15574) );
  AND U16514 ( .A(n15756), .B(n15757), .Z(n15754) );
  AND U16515 ( .A(a[21]), .B(b[20]), .Z(n15753) );
  XOR U16516 ( .A(n15758), .B(n15579), .Z(n15581) );
  XOR U16517 ( .A(n15759), .B(n15760), .Z(n15579) );
  AND U16518 ( .A(n15761), .B(n15762), .Z(n15759) );
  AND U16519 ( .A(b[19]), .B(a[22]), .Z(n15758) );
  XOR U16520 ( .A(n15763), .B(n15584), .Z(n15586) );
  XOR U16521 ( .A(n15764), .B(n15765), .Z(n15584) );
  AND U16522 ( .A(n15766), .B(n15767), .Z(n15764) );
  AND U16523 ( .A(a[23]), .B(b[18]), .Z(n15763) );
  XOR U16524 ( .A(n15768), .B(n15589), .Z(n15591) );
  XOR U16525 ( .A(n15769), .B(n15770), .Z(n15589) );
  AND U16526 ( .A(n15771), .B(n15772), .Z(n15769) );
  AND U16527 ( .A(b[17]), .B(a[24]), .Z(n15768) );
  XOR U16528 ( .A(n15773), .B(n15594), .Z(n15596) );
  XOR U16529 ( .A(n15774), .B(n15775), .Z(n15594) );
  AND U16530 ( .A(n15776), .B(n15777), .Z(n15774) );
  AND U16531 ( .A(a[25]), .B(b[16]), .Z(n15773) );
  XOR U16532 ( .A(n15778), .B(n15599), .Z(n15601) );
  XOR U16533 ( .A(n15779), .B(n15780), .Z(n15599) );
  AND U16534 ( .A(n15781), .B(n15782), .Z(n15779) );
  AND U16535 ( .A(b[15]), .B(a[26]), .Z(n15778) );
  XOR U16536 ( .A(n15783), .B(n15604), .Z(n15606) );
  XOR U16537 ( .A(n15784), .B(n15785), .Z(n15604) );
  AND U16538 ( .A(n15786), .B(n15787), .Z(n15784) );
  AND U16539 ( .A(a[27]), .B(b[14]), .Z(n15783) );
  XOR U16540 ( .A(n15788), .B(n15609), .Z(n15611) );
  XOR U16541 ( .A(n15789), .B(n15790), .Z(n15609) );
  AND U16542 ( .A(n15791), .B(n15792), .Z(n15789) );
  AND U16543 ( .A(b[13]), .B(a[28]), .Z(n15788) );
  XOR U16544 ( .A(n15793), .B(n15614), .Z(n15616) );
  XOR U16545 ( .A(n15794), .B(n15795), .Z(n15614) );
  AND U16546 ( .A(n15796), .B(n15797), .Z(n15794) );
  AND U16547 ( .A(a[29]), .B(b[12]), .Z(n15793) );
  XOR U16548 ( .A(n15798), .B(n15619), .Z(n15621) );
  XOR U16549 ( .A(n15799), .B(n15800), .Z(n15619) );
  AND U16550 ( .A(n15801), .B(n15802), .Z(n15799) );
  AND U16551 ( .A(b[11]), .B(a[30]), .Z(n15798) );
  XOR U16552 ( .A(n15803), .B(n15624), .Z(n15626) );
  XOR U16553 ( .A(n15804), .B(n15805), .Z(n15624) );
  AND U16554 ( .A(n15806), .B(n15807), .Z(n15804) );
  AND U16555 ( .A(a[31]), .B(b[10]), .Z(n15803) );
  XOR U16556 ( .A(n15808), .B(n15629), .Z(n15631) );
  XOR U16557 ( .A(n15809), .B(n15810), .Z(n15629) );
  AND U16558 ( .A(n15811), .B(n15812), .Z(n15809) );
  AND U16559 ( .A(a[32]), .B(b[9]), .Z(n15808) );
  XOR U16560 ( .A(n15813), .B(n15634), .Z(n15636) );
  XOR U16561 ( .A(n15814), .B(n15815), .Z(n15634) );
  AND U16562 ( .A(n15816), .B(n15817), .Z(n15814) );
  AND U16563 ( .A(a[33]), .B(b[8]), .Z(n15813) );
  XOR U16564 ( .A(n15818), .B(n15639), .Z(n15641) );
  XOR U16565 ( .A(n15819), .B(n15820), .Z(n15639) );
  AND U16566 ( .A(n15821), .B(n15822), .Z(n15819) );
  AND U16567 ( .A(a[34]), .B(b[7]), .Z(n15818) );
  XOR U16568 ( .A(n15823), .B(n15644), .Z(n15646) );
  XOR U16569 ( .A(n15824), .B(n15825), .Z(n15644) );
  AND U16570 ( .A(n15826), .B(n15827), .Z(n15824) );
  AND U16571 ( .A(a[35]), .B(b[6]), .Z(n15823) );
  XOR U16572 ( .A(n15828), .B(n15829), .Z(n15648) );
  AND U16573 ( .A(n15830), .B(n15831), .Z(n15828) );
  XOR U16574 ( .A(n15832), .B(n15653), .Z(n15655) );
  XOR U16575 ( .A(n15833), .B(n15834), .Z(n15653) );
  AND U16576 ( .A(n15835), .B(n15836), .Z(n15833) );
  AND U16577 ( .A(a[36]), .B(b[5]), .Z(n15832) );
  XOR U16578 ( .A(n15838), .B(n15839), .Z(n15658) );
  AND U16579 ( .A(n15672), .B(n15670), .Z(n15838) );
  AND U16580 ( .A(b[2]), .B(a[38]), .Z(n15840) );
  XOR U16581 ( .A(n15830), .B(n15839), .Z(n15841) );
  XOR U16582 ( .A(n15842), .B(n15843), .Z(n15839) );
  NANDN U16583 ( .A(n15674), .B(n15673), .Z(n15843) );
  XOR U16584 ( .A(n15844), .B(n15845), .Z(n15673) );
  NAND U16585 ( .A(a[38]), .B(b[1]), .Z(n15845) );
  XOR U16586 ( .A(n15846), .B(n15847), .Z(n15674) );
  XOR U16587 ( .A(n15844), .B(n15848), .Z(n15847) );
  IV U16588 ( .A(n15842), .Z(n15844) );
  ANDN U16589 ( .B(n5362), .A(n5364), .Z(n15842) );
  NAND U16590 ( .A(a[38]), .B(b[0]), .Z(n5364) );
  XNOR U16591 ( .A(n15849), .B(n15850), .Z(n5362) );
  XOR U16592 ( .A(n15851), .B(n15829), .Z(n15830) );
  AND U16593 ( .A(b[3]), .B(a[37]), .Z(n15851) );
  XNOR U16594 ( .A(n15829), .B(n15835), .Z(n15852) );
  XNOR U16595 ( .A(n15834), .B(n15826), .Z(n15853) );
  XNOR U16596 ( .A(n15825), .B(n15821), .Z(n15854) );
  XNOR U16597 ( .A(n15820), .B(n15816), .Z(n15855) );
  XNOR U16598 ( .A(n15815), .B(n15811), .Z(n15856) );
  XNOR U16599 ( .A(n15810), .B(n15806), .Z(n15857) );
  XNOR U16600 ( .A(n15805), .B(n15801), .Z(n15858) );
  XNOR U16601 ( .A(n15800), .B(n15796), .Z(n15859) );
  XNOR U16602 ( .A(n15795), .B(n15791), .Z(n15860) );
  XNOR U16603 ( .A(n15790), .B(n15786), .Z(n15861) );
  XNOR U16604 ( .A(n15785), .B(n15781), .Z(n15862) );
  XNOR U16605 ( .A(n15780), .B(n15776), .Z(n15863) );
  XNOR U16606 ( .A(n15775), .B(n15771), .Z(n15864) );
  XNOR U16607 ( .A(n15770), .B(n15766), .Z(n15865) );
  XNOR U16608 ( .A(n15765), .B(n15761), .Z(n15866) );
  XNOR U16609 ( .A(n15760), .B(n15756), .Z(n15867) );
  XNOR U16610 ( .A(n15755), .B(n15751), .Z(n15868) );
  XNOR U16611 ( .A(n15750), .B(n15746), .Z(n15869) );
  XNOR U16612 ( .A(n15745), .B(n15741), .Z(n15870) );
  XNOR U16613 ( .A(n15740), .B(n15736), .Z(n15871) );
  XNOR U16614 ( .A(n15735), .B(n15731), .Z(n15872) );
  XNOR U16615 ( .A(n15730), .B(n15726), .Z(n15873) );
  XNOR U16616 ( .A(n15725), .B(n15721), .Z(n15874) );
  XNOR U16617 ( .A(n15720), .B(n15716), .Z(n15875) );
  XOR U16618 ( .A(n15715), .B(n15712), .Z(n15876) );
  XOR U16619 ( .A(n15877), .B(n15878), .Z(n15712) );
  XOR U16620 ( .A(n15710), .B(n15879), .Z(n15878) );
  XOR U16621 ( .A(n15880), .B(n15881), .Z(n15879) );
  XOR U16622 ( .A(n15882), .B(n15883), .Z(n15881) );
  NAND U16623 ( .A(a[10]), .B(b[30]), .Z(n15883) );
  AND U16624 ( .A(a[9]), .B(b[31]), .Z(n15882) );
  XOR U16625 ( .A(n15884), .B(n15880), .Z(n15877) );
  XOR U16626 ( .A(n15885), .B(n15886), .Z(n15880) );
  ANDN U16627 ( .B(n15887), .A(n15888), .Z(n15885) );
  AND U16628 ( .A(a[11]), .B(b[29]), .Z(n15884) );
  XOR U16629 ( .A(n15889), .B(n15710), .Z(n15711) );
  XOR U16630 ( .A(n15890), .B(n15891), .Z(n15710) );
  AND U16631 ( .A(n15892), .B(n15893), .Z(n15890) );
  AND U16632 ( .A(a[12]), .B(b[28]), .Z(n15889) );
  XOR U16633 ( .A(n15894), .B(n15715), .Z(n15717) );
  XOR U16634 ( .A(n15895), .B(n15896), .Z(n15715) );
  AND U16635 ( .A(n15897), .B(n15898), .Z(n15895) );
  AND U16636 ( .A(a[13]), .B(b[27]), .Z(n15894) );
  XOR U16637 ( .A(n15899), .B(n15720), .Z(n15722) );
  XOR U16638 ( .A(n15900), .B(n15901), .Z(n15720) );
  AND U16639 ( .A(n15902), .B(n15903), .Z(n15900) );
  AND U16640 ( .A(a[14]), .B(b[26]), .Z(n15899) );
  XOR U16641 ( .A(n15904), .B(n15725), .Z(n15727) );
  XOR U16642 ( .A(n15905), .B(n15906), .Z(n15725) );
  AND U16643 ( .A(n15907), .B(n15908), .Z(n15905) );
  AND U16644 ( .A(a[15]), .B(b[25]), .Z(n15904) );
  XOR U16645 ( .A(n15909), .B(n15730), .Z(n15732) );
  XOR U16646 ( .A(n15910), .B(n15911), .Z(n15730) );
  AND U16647 ( .A(n15912), .B(n15913), .Z(n15910) );
  AND U16648 ( .A(a[16]), .B(b[24]), .Z(n15909) );
  XOR U16649 ( .A(n15914), .B(n15735), .Z(n15737) );
  XOR U16650 ( .A(n15915), .B(n15916), .Z(n15735) );
  AND U16651 ( .A(n15917), .B(n15918), .Z(n15915) );
  AND U16652 ( .A(a[17]), .B(b[23]), .Z(n15914) );
  XOR U16653 ( .A(n15919), .B(n15740), .Z(n15742) );
  XOR U16654 ( .A(n15920), .B(n15921), .Z(n15740) );
  AND U16655 ( .A(n15922), .B(n15923), .Z(n15920) );
  AND U16656 ( .A(a[18]), .B(b[22]), .Z(n15919) );
  XOR U16657 ( .A(n15924), .B(n15745), .Z(n15747) );
  XOR U16658 ( .A(n15925), .B(n15926), .Z(n15745) );
  AND U16659 ( .A(n15927), .B(n15928), .Z(n15925) );
  AND U16660 ( .A(a[19]), .B(b[21]), .Z(n15924) );
  XOR U16661 ( .A(n15929), .B(n15750), .Z(n15752) );
  XOR U16662 ( .A(n15930), .B(n15931), .Z(n15750) );
  AND U16663 ( .A(n15932), .B(n15933), .Z(n15930) );
  AND U16664 ( .A(b[20]), .B(a[20]), .Z(n15929) );
  XOR U16665 ( .A(n15934), .B(n15755), .Z(n15757) );
  XOR U16666 ( .A(n15935), .B(n15936), .Z(n15755) );
  AND U16667 ( .A(n15937), .B(n15938), .Z(n15935) );
  AND U16668 ( .A(a[21]), .B(b[19]), .Z(n15934) );
  XOR U16669 ( .A(n15939), .B(n15760), .Z(n15762) );
  XOR U16670 ( .A(n15940), .B(n15941), .Z(n15760) );
  AND U16671 ( .A(n15942), .B(n15943), .Z(n15940) );
  AND U16672 ( .A(b[18]), .B(a[22]), .Z(n15939) );
  XOR U16673 ( .A(n15944), .B(n15765), .Z(n15767) );
  XOR U16674 ( .A(n15945), .B(n15946), .Z(n15765) );
  AND U16675 ( .A(n15947), .B(n15948), .Z(n15945) );
  AND U16676 ( .A(a[23]), .B(b[17]), .Z(n15944) );
  XOR U16677 ( .A(n15949), .B(n15770), .Z(n15772) );
  XOR U16678 ( .A(n15950), .B(n15951), .Z(n15770) );
  AND U16679 ( .A(n15952), .B(n15953), .Z(n15950) );
  AND U16680 ( .A(b[16]), .B(a[24]), .Z(n15949) );
  XOR U16681 ( .A(n15954), .B(n15775), .Z(n15777) );
  XOR U16682 ( .A(n15955), .B(n15956), .Z(n15775) );
  AND U16683 ( .A(n15957), .B(n15958), .Z(n15955) );
  AND U16684 ( .A(a[25]), .B(b[15]), .Z(n15954) );
  XOR U16685 ( .A(n15959), .B(n15780), .Z(n15782) );
  XOR U16686 ( .A(n15960), .B(n15961), .Z(n15780) );
  AND U16687 ( .A(n15962), .B(n15963), .Z(n15960) );
  AND U16688 ( .A(b[14]), .B(a[26]), .Z(n15959) );
  XOR U16689 ( .A(n15964), .B(n15785), .Z(n15787) );
  XOR U16690 ( .A(n15965), .B(n15966), .Z(n15785) );
  AND U16691 ( .A(n15967), .B(n15968), .Z(n15965) );
  AND U16692 ( .A(a[27]), .B(b[13]), .Z(n15964) );
  XOR U16693 ( .A(n15969), .B(n15790), .Z(n15792) );
  XOR U16694 ( .A(n15970), .B(n15971), .Z(n15790) );
  AND U16695 ( .A(n15972), .B(n15973), .Z(n15970) );
  AND U16696 ( .A(b[12]), .B(a[28]), .Z(n15969) );
  XOR U16697 ( .A(n15974), .B(n15795), .Z(n15797) );
  XOR U16698 ( .A(n15975), .B(n15976), .Z(n15795) );
  AND U16699 ( .A(n15977), .B(n15978), .Z(n15975) );
  AND U16700 ( .A(a[29]), .B(b[11]), .Z(n15974) );
  XOR U16701 ( .A(n15979), .B(n15800), .Z(n15802) );
  XOR U16702 ( .A(n15980), .B(n15981), .Z(n15800) );
  AND U16703 ( .A(n15982), .B(n15983), .Z(n15980) );
  AND U16704 ( .A(b[10]), .B(a[30]), .Z(n15979) );
  XOR U16705 ( .A(n15984), .B(n15805), .Z(n15807) );
  XOR U16706 ( .A(n15985), .B(n15986), .Z(n15805) );
  AND U16707 ( .A(n15987), .B(n15988), .Z(n15985) );
  AND U16708 ( .A(a[31]), .B(b[9]), .Z(n15984) );
  XOR U16709 ( .A(n15989), .B(n15810), .Z(n15812) );
  XOR U16710 ( .A(n15990), .B(n15991), .Z(n15810) );
  AND U16711 ( .A(n15992), .B(n15993), .Z(n15990) );
  AND U16712 ( .A(a[32]), .B(b[8]), .Z(n15989) );
  XOR U16713 ( .A(n15994), .B(n15815), .Z(n15817) );
  XOR U16714 ( .A(n15995), .B(n15996), .Z(n15815) );
  AND U16715 ( .A(n15997), .B(n15998), .Z(n15995) );
  AND U16716 ( .A(a[33]), .B(b[7]), .Z(n15994) );
  XOR U16717 ( .A(n15999), .B(n15820), .Z(n15822) );
  XOR U16718 ( .A(n16000), .B(n16001), .Z(n15820) );
  AND U16719 ( .A(n16002), .B(n16003), .Z(n16000) );
  AND U16720 ( .A(a[34]), .B(b[6]), .Z(n15999) );
  XOR U16721 ( .A(n16004), .B(n15825), .Z(n15827) );
  XOR U16722 ( .A(n16005), .B(n16006), .Z(n15825) );
  AND U16723 ( .A(n16007), .B(n16008), .Z(n16005) );
  AND U16724 ( .A(a[35]), .B(b[5]), .Z(n16004) );
  XNOR U16725 ( .A(n16009), .B(n16010), .Z(n15829) );
  AND U16726 ( .A(n15848), .B(n15846), .Z(n16009) );
  XNOR U16727 ( .A(n16011), .B(n16012), .Z(n15846) );
  XOR U16728 ( .A(n16010), .B(n16013), .Z(n16012) );
  XNOR U16729 ( .A(n16014), .B(n16010), .Z(n15848) );
  XOR U16730 ( .A(n16015), .B(n16016), .Z(n16010) );
  NANDN U16731 ( .A(n15850), .B(n15849), .Z(n16016) );
  XNOR U16732 ( .A(n16017), .B(n16018), .Z(n15849) );
  XNOR U16733 ( .A(n16015), .B(n16019), .Z(n16018) );
  XOR U16734 ( .A(n16015), .B(n16020), .Z(n15850) );
  NAND U16735 ( .A(b[1]), .B(a[37]), .Z(n16020) );
  ANDN U16736 ( .B(n5367), .A(n5369), .Z(n16015) );
  NAND U16737 ( .A(a[37]), .B(b[0]), .Z(n5369) );
  XOR U16738 ( .A(n16021), .B(n16022), .Z(n5367) );
  AND U16739 ( .A(b[2]), .B(a[37]), .Z(n16014) );
  XOR U16740 ( .A(n16023), .B(n15834), .Z(n15836) );
  XOR U16741 ( .A(n16024), .B(n16025), .Z(n15834) );
  AND U16742 ( .A(n16013), .B(n16011), .Z(n16024) );
  XOR U16743 ( .A(n16026), .B(n16025), .Z(n16011) );
  AND U16744 ( .A(a[36]), .B(b[3]), .Z(n16026) );
  XNOR U16745 ( .A(n16025), .B(n16007), .Z(n16027) );
  XNOR U16746 ( .A(n16006), .B(n16002), .Z(n16028) );
  XNOR U16747 ( .A(n16001), .B(n15997), .Z(n16029) );
  XNOR U16748 ( .A(n15996), .B(n15992), .Z(n16030) );
  XNOR U16749 ( .A(n15991), .B(n15987), .Z(n16031) );
  XNOR U16750 ( .A(n15986), .B(n15982), .Z(n16032) );
  XNOR U16751 ( .A(n15981), .B(n15977), .Z(n16033) );
  XNOR U16752 ( .A(n15976), .B(n15972), .Z(n16034) );
  XNOR U16753 ( .A(n15971), .B(n15967), .Z(n16035) );
  XNOR U16754 ( .A(n15966), .B(n15962), .Z(n16036) );
  XNOR U16755 ( .A(n15961), .B(n15957), .Z(n16037) );
  XNOR U16756 ( .A(n15956), .B(n15952), .Z(n16038) );
  XNOR U16757 ( .A(n15951), .B(n15947), .Z(n16039) );
  XNOR U16758 ( .A(n15946), .B(n15942), .Z(n16040) );
  XNOR U16759 ( .A(n15941), .B(n15937), .Z(n16041) );
  XNOR U16760 ( .A(n15936), .B(n15932), .Z(n16042) );
  XNOR U16761 ( .A(n15931), .B(n15927), .Z(n16043) );
  XNOR U16762 ( .A(n15926), .B(n15922), .Z(n16044) );
  XNOR U16763 ( .A(n15921), .B(n15917), .Z(n16045) );
  XNOR U16764 ( .A(n15916), .B(n15912), .Z(n16046) );
  XNOR U16765 ( .A(n15911), .B(n15907), .Z(n16047) );
  XNOR U16766 ( .A(n15906), .B(n15902), .Z(n16048) );
  XNOR U16767 ( .A(n15901), .B(n15897), .Z(n16049) );
  XNOR U16768 ( .A(n15896), .B(n15892), .Z(n16050) );
  XOR U16769 ( .A(n15891), .B(n15888), .Z(n16051) );
  XOR U16770 ( .A(n16052), .B(n16053), .Z(n15888) );
  XOR U16771 ( .A(n15886), .B(n16054), .Z(n16053) );
  XOR U16772 ( .A(n16055), .B(n16056), .Z(n16054) );
  XOR U16773 ( .A(n16057), .B(n16058), .Z(n16056) );
  NAND U16774 ( .A(a[9]), .B(b[30]), .Z(n16058) );
  AND U16775 ( .A(a[8]), .B(b[31]), .Z(n16057) );
  XOR U16776 ( .A(n16059), .B(n16055), .Z(n16052) );
  XOR U16777 ( .A(n16060), .B(n16061), .Z(n16055) );
  ANDN U16778 ( .B(n16062), .A(n16063), .Z(n16060) );
  AND U16779 ( .A(a[10]), .B(b[29]), .Z(n16059) );
  XOR U16780 ( .A(n16064), .B(n15886), .Z(n15887) );
  XOR U16781 ( .A(n16065), .B(n16066), .Z(n15886) );
  AND U16782 ( .A(n16067), .B(n16068), .Z(n16065) );
  AND U16783 ( .A(a[11]), .B(b[28]), .Z(n16064) );
  XOR U16784 ( .A(n16069), .B(n15891), .Z(n15893) );
  XOR U16785 ( .A(n16070), .B(n16071), .Z(n15891) );
  AND U16786 ( .A(n16072), .B(n16073), .Z(n16070) );
  AND U16787 ( .A(a[12]), .B(b[27]), .Z(n16069) );
  XOR U16788 ( .A(n16074), .B(n15896), .Z(n15898) );
  XOR U16789 ( .A(n16075), .B(n16076), .Z(n15896) );
  AND U16790 ( .A(n16077), .B(n16078), .Z(n16075) );
  AND U16791 ( .A(a[13]), .B(b[26]), .Z(n16074) );
  XOR U16792 ( .A(n16079), .B(n15901), .Z(n15903) );
  XOR U16793 ( .A(n16080), .B(n16081), .Z(n15901) );
  AND U16794 ( .A(n16082), .B(n16083), .Z(n16080) );
  AND U16795 ( .A(a[14]), .B(b[25]), .Z(n16079) );
  XOR U16796 ( .A(n16084), .B(n15906), .Z(n15908) );
  XOR U16797 ( .A(n16085), .B(n16086), .Z(n15906) );
  AND U16798 ( .A(n16087), .B(n16088), .Z(n16085) );
  AND U16799 ( .A(a[15]), .B(b[24]), .Z(n16084) );
  XOR U16800 ( .A(n16089), .B(n15911), .Z(n15913) );
  XOR U16801 ( .A(n16090), .B(n16091), .Z(n15911) );
  AND U16802 ( .A(n16092), .B(n16093), .Z(n16090) );
  AND U16803 ( .A(a[16]), .B(b[23]), .Z(n16089) );
  XOR U16804 ( .A(n16094), .B(n15916), .Z(n15918) );
  XOR U16805 ( .A(n16095), .B(n16096), .Z(n15916) );
  AND U16806 ( .A(n16097), .B(n16098), .Z(n16095) );
  AND U16807 ( .A(a[17]), .B(b[22]), .Z(n16094) );
  XOR U16808 ( .A(n16099), .B(n15921), .Z(n15923) );
  XOR U16809 ( .A(n16100), .B(n16101), .Z(n15921) );
  AND U16810 ( .A(n16102), .B(n16103), .Z(n16100) );
  AND U16811 ( .A(a[18]), .B(b[21]), .Z(n16099) );
  XOR U16812 ( .A(n16104), .B(n15926), .Z(n15928) );
  XOR U16813 ( .A(n16105), .B(n16106), .Z(n15926) );
  AND U16814 ( .A(n16107), .B(n16108), .Z(n16105) );
  AND U16815 ( .A(a[19]), .B(b[20]), .Z(n16104) );
  XOR U16816 ( .A(n16109), .B(n15931), .Z(n15933) );
  XOR U16817 ( .A(n16110), .B(n16111), .Z(n15931) );
  AND U16818 ( .A(n16112), .B(n16113), .Z(n16110) );
  AND U16819 ( .A(b[19]), .B(a[20]), .Z(n16109) );
  XOR U16820 ( .A(n16114), .B(n15936), .Z(n15938) );
  XOR U16821 ( .A(n16115), .B(n16116), .Z(n15936) );
  AND U16822 ( .A(n16117), .B(n16118), .Z(n16115) );
  AND U16823 ( .A(a[21]), .B(b[18]), .Z(n16114) );
  XOR U16824 ( .A(n16119), .B(n15941), .Z(n15943) );
  XOR U16825 ( .A(n16120), .B(n16121), .Z(n15941) );
  AND U16826 ( .A(n16122), .B(n16123), .Z(n16120) );
  AND U16827 ( .A(b[17]), .B(a[22]), .Z(n16119) );
  XOR U16828 ( .A(n16124), .B(n15946), .Z(n15948) );
  XOR U16829 ( .A(n16125), .B(n16126), .Z(n15946) );
  AND U16830 ( .A(n16127), .B(n16128), .Z(n16125) );
  AND U16831 ( .A(a[23]), .B(b[16]), .Z(n16124) );
  XOR U16832 ( .A(n16129), .B(n15951), .Z(n15953) );
  XOR U16833 ( .A(n16130), .B(n16131), .Z(n15951) );
  AND U16834 ( .A(n16132), .B(n16133), .Z(n16130) );
  AND U16835 ( .A(b[15]), .B(a[24]), .Z(n16129) );
  XOR U16836 ( .A(n16134), .B(n15956), .Z(n15958) );
  XOR U16837 ( .A(n16135), .B(n16136), .Z(n15956) );
  AND U16838 ( .A(n16137), .B(n16138), .Z(n16135) );
  AND U16839 ( .A(a[25]), .B(b[14]), .Z(n16134) );
  XOR U16840 ( .A(n16139), .B(n15961), .Z(n15963) );
  XOR U16841 ( .A(n16140), .B(n16141), .Z(n15961) );
  AND U16842 ( .A(n16142), .B(n16143), .Z(n16140) );
  AND U16843 ( .A(b[13]), .B(a[26]), .Z(n16139) );
  XOR U16844 ( .A(n16144), .B(n15966), .Z(n15968) );
  XOR U16845 ( .A(n16145), .B(n16146), .Z(n15966) );
  AND U16846 ( .A(n16147), .B(n16148), .Z(n16145) );
  AND U16847 ( .A(a[27]), .B(b[12]), .Z(n16144) );
  XOR U16848 ( .A(n16149), .B(n15971), .Z(n15973) );
  XOR U16849 ( .A(n16150), .B(n16151), .Z(n15971) );
  AND U16850 ( .A(n16152), .B(n16153), .Z(n16150) );
  AND U16851 ( .A(b[11]), .B(a[28]), .Z(n16149) );
  XOR U16852 ( .A(n16154), .B(n15976), .Z(n15978) );
  XOR U16853 ( .A(n16155), .B(n16156), .Z(n15976) );
  AND U16854 ( .A(n16157), .B(n16158), .Z(n16155) );
  AND U16855 ( .A(a[29]), .B(b[10]), .Z(n16154) );
  XOR U16856 ( .A(n16159), .B(n15981), .Z(n15983) );
  XOR U16857 ( .A(n16160), .B(n16161), .Z(n15981) );
  AND U16858 ( .A(n16162), .B(n16163), .Z(n16160) );
  AND U16859 ( .A(b[9]), .B(a[30]), .Z(n16159) );
  XOR U16860 ( .A(n16164), .B(n15986), .Z(n15988) );
  XOR U16861 ( .A(n16165), .B(n16166), .Z(n15986) );
  AND U16862 ( .A(n16167), .B(n16168), .Z(n16165) );
  AND U16863 ( .A(a[31]), .B(b[8]), .Z(n16164) );
  XOR U16864 ( .A(n16169), .B(n15991), .Z(n15993) );
  XOR U16865 ( .A(n16170), .B(n16171), .Z(n15991) );
  AND U16866 ( .A(n16172), .B(n16173), .Z(n16170) );
  AND U16867 ( .A(a[32]), .B(b[7]), .Z(n16169) );
  XOR U16868 ( .A(n16174), .B(n15996), .Z(n15998) );
  XOR U16869 ( .A(n16175), .B(n16176), .Z(n15996) );
  AND U16870 ( .A(n16177), .B(n16178), .Z(n16175) );
  AND U16871 ( .A(a[33]), .B(b[6]), .Z(n16174) );
  XOR U16872 ( .A(n16179), .B(n16001), .Z(n16003) );
  XOR U16873 ( .A(n16180), .B(n16181), .Z(n16001) );
  AND U16874 ( .A(n16182), .B(n16183), .Z(n16180) );
  AND U16875 ( .A(a[34]), .B(b[5]), .Z(n16179) );
  XNOR U16876 ( .A(n16184), .B(n16185), .Z(n16025) );
  AND U16877 ( .A(n16019), .B(n16017), .Z(n16184) );
  XNOR U16878 ( .A(n16186), .B(n16187), .Z(n16017) );
  XOR U16879 ( .A(n16185), .B(n16188), .Z(n16187) );
  XNOR U16880 ( .A(n16189), .B(n16185), .Z(n16019) );
  XNOR U16881 ( .A(n16190), .B(n16191), .Z(n16185) );
  OR U16882 ( .A(n16022), .B(n16021), .Z(n16191) );
  XNOR U16883 ( .A(n16190), .B(n16192), .Z(n16021) );
  NAND U16884 ( .A(a[36]), .B(b[1]), .Z(n16192) );
  XOR U16885 ( .A(n16193), .B(n16194), .Z(n16022) );
  XOR U16886 ( .A(n16190), .B(n16195), .Z(n16194) );
  NANDN U16887 ( .A(n5374), .B(n5372), .Z(n16190) );
  XNOR U16888 ( .A(n16196), .B(n16197), .Z(n5372) );
  NAND U16889 ( .A(a[36]), .B(b[0]), .Z(n5374) );
  AND U16890 ( .A(b[2]), .B(a[36]), .Z(n16189) );
  XOR U16891 ( .A(n16198), .B(n16006), .Z(n16008) );
  XNOR U16892 ( .A(n16199), .B(n16200), .Z(n16006) );
  AND U16893 ( .A(n16188), .B(n16186), .Z(n16199) );
  XNOR U16894 ( .A(n16201), .B(n16200), .Z(n16186) );
  AND U16895 ( .A(a[35]), .B(b[3]), .Z(n16201) );
  XOR U16896 ( .A(n16200), .B(n16182), .Z(n16202) );
  XNOR U16897 ( .A(n16181), .B(n16177), .Z(n16203) );
  XNOR U16898 ( .A(n16176), .B(n16172), .Z(n16204) );
  XNOR U16899 ( .A(n16171), .B(n16167), .Z(n16205) );
  XNOR U16900 ( .A(n16166), .B(n16162), .Z(n16206) );
  XNOR U16901 ( .A(n16161), .B(n16157), .Z(n16207) );
  XNOR U16902 ( .A(n16156), .B(n16152), .Z(n16208) );
  XNOR U16903 ( .A(n16151), .B(n16147), .Z(n16209) );
  XNOR U16904 ( .A(n16146), .B(n16142), .Z(n16210) );
  XNOR U16905 ( .A(n16141), .B(n16137), .Z(n16211) );
  XNOR U16906 ( .A(n16136), .B(n16132), .Z(n16212) );
  XNOR U16907 ( .A(n16131), .B(n16127), .Z(n16213) );
  XNOR U16908 ( .A(n16126), .B(n16122), .Z(n16214) );
  XNOR U16909 ( .A(n16121), .B(n16117), .Z(n16215) );
  XNOR U16910 ( .A(n16116), .B(n16112), .Z(n16216) );
  XNOR U16911 ( .A(n16111), .B(n16107), .Z(n16217) );
  XNOR U16912 ( .A(n16106), .B(n16102), .Z(n16218) );
  XNOR U16913 ( .A(n16101), .B(n16097), .Z(n16219) );
  XNOR U16914 ( .A(n16096), .B(n16092), .Z(n16220) );
  XNOR U16915 ( .A(n16091), .B(n16087), .Z(n16221) );
  XNOR U16916 ( .A(n16086), .B(n16082), .Z(n16222) );
  XNOR U16917 ( .A(n16081), .B(n16077), .Z(n16223) );
  XNOR U16918 ( .A(n16076), .B(n16072), .Z(n16224) );
  XNOR U16919 ( .A(n16071), .B(n16067), .Z(n16225) );
  XOR U16920 ( .A(n16066), .B(n16063), .Z(n16226) );
  XOR U16921 ( .A(n16227), .B(n16228), .Z(n16063) );
  XOR U16922 ( .A(n16061), .B(n16229), .Z(n16228) );
  XNOR U16923 ( .A(n16230), .B(n16231), .Z(n16229) );
  XOR U16924 ( .A(n16232), .B(n16233), .Z(n16231) );
  NAND U16925 ( .A(a[8]), .B(b[30]), .Z(n16233) );
  AND U16926 ( .A(a[7]), .B(b[31]), .Z(n16232) );
  XNOR U16927 ( .A(n16234), .B(n16230), .Z(n16227) );
  XNOR U16928 ( .A(n16235), .B(n16236), .Z(n16230) );
  ANDN U16929 ( .B(n16237), .A(n16238), .Z(n16235) );
  AND U16930 ( .A(a[9]), .B(b[29]), .Z(n16234) );
  XOR U16931 ( .A(n16239), .B(n16061), .Z(n16062) );
  XOR U16932 ( .A(n16240), .B(n16241), .Z(n16061) );
  AND U16933 ( .A(n16242), .B(n16243), .Z(n16240) );
  AND U16934 ( .A(a[10]), .B(b[28]), .Z(n16239) );
  XOR U16935 ( .A(n16244), .B(n16066), .Z(n16068) );
  XOR U16936 ( .A(n16245), .B(n16246), .Z(n16066) );
  AND U16937 ( .A(n16247), .B(n16248), .Z(n16245) );
  AND U16938 ( .A(a[11]), .B(b[27]), .Z(n16244) );
  XOR U16939 ( .A(n16249), .B(n16071), .Z(n16073) );
  XOR U16940 ( .A(n16250), .B(n16251), .Z(n16071) );
  AND U16941 ( .A(n16252), .B(n16253), .Z(n16250) );
  AND U16942 ( .A(a[12]), .B(b[26]), .Z(n16249) );
  XOR U16943 ( .A(n16254), .B(n16076), .Z(n16078) );
  XOR U16944 ( .A(n16255), .B(n16256), .Z(n16076) );
  AND U16945 ( .A(n16257), .B(n16258), .Z(n16255) );
  AND U16946 ( .A(a[13]), .B(b[25]), .Z(n16254) );
  XOR U16947 ( .A(n16259), .B(n16081), .Z(n16083) );
  XOR U16948 ( .A(n16260), .B(n16261), .Z(n16081) );
  AND U16949 ( .A(n16262), .B(n16263), .Z(n16260) );
  AND U16950 ( .A(a[14]), .B(b[24]), .Z(n16259) );
  XOR U16951 ( .A(n16264), .B(n16086), .Z(n16088) );
  XOR U16952 ( .A(n16265), .B(n16266), .Z(n16086) );
  AND U16953 ( .A(n16267), .B(n16268), .Z(n16265) );
  AND U16954 ( .A(a[15]), .B(b[23]), .Z(n16264) );
  XOR U16955 ( .A(n16269), .B(n16091), .Z(n16093) );
  XOR U16956 ( .A(n16270), .B(n16271), .Z(n16091) );
  AND U16957 ( .A(n16272), .B(n16273), .Z(n16270) );
  AND U16958 ( .A(a[16]), .B(b[22]), .Z(n16269) );
  XOR U16959 ( .A(n16274), .B(n16096), .Z(n16098) );
  XOR U16960 ( .A(n16275), .B(n16276), .Z(n16096) );
  AND U16961 ( .A(n16277), .B(n16278), .Z(n16275) );
  AND U16962 ( .A(a[17]), .B(b[21]), .Z(n16274) );
  XOR U16963 ( .A(n16279), .B(n16101), .Z(n16103) );
  XOR U16964 ( .A(n16280), .B(n16281), .Z(n16101) );
  AND U16965 ( .A(n16282), .B(n16283), .Z(n16280) );
  AND U16966 ( .A(a[18]), .B(b[20]), .Z(n16279) );
  XOR U16967 ( .A(n16284), .B(n16106), .Z(n16108) );
  XOR U16968 ( .A(n16285), .B(n16286), .Z(n16106) );
  AND U16969 ( .A(n16287), .B(n16288), .Z(n16285) );
  AND U16970 ( .A(a[19]), .B(b[19]), .Z(n16284) );
  XOR U16971 ( .A(n16289), .B(n16111), .Z(n16113) );
  XOR U16972 ( .A(n16290), .B(n16291), .Z(n16111) );
  AND U16973 ( .A(n16292), .B(n16293), .Z(n16290) );
  AND U16974 ( .A(b[18]), .B(a[20]), .Z(n16289) );
  XOR U16975 ( .A(n16294), .B(n16116), .Z(n16118) );
  XOR U16976 ( .A(n16295), .B(n16296), .Z(n16116) );
  AND U16977 ( .A(n16297), .B(n16298), .Z(n16295) );
  AND U16978 ( .A(a[21]), .B(b[17]), .Z(n16294) );
  XOR U16979 ( .A(n16299), .B(n16121), .Z(n16123) );
  XOR U16980 ( .A(n16300), .B(n16301), .Z(n16121) );
  AND U16981 ( .A(n16302), .B(n16303), .Z(n16300) );
  AND U16982 ( .A(b[16]), .B(a[22]), .Z(n16299) );
  XOR U16983 ( .A(n16304), .B(n16126), .Z(n16128) );
  XOR U16984 ( .A(n16305), .B(n16306), .Z(n16126) );
  AND U16985 ( .A(n16307), .B(n16308), .Z(n16305) );
  AND U16986 ( .A(a[23]), .B(b[15]), .Z(n16304) );
  XOR U16987 ( .A(n16309), .B(n16131), .Z(n16133) );
  XOR U16988 ( .A(n16310), .B(n16311), .Z(n16131) );
  AND U16989 ( .A(n16312), .B(n16313), .Z(n16310) );
  AND U16990 ( .A(b[14]), .B(a[24]), .Z(n16309) );
  XOR U16991 ( .A(n16314), .B(n16136), .Z(n16138) );
  XOR U16992 ( .A(n16315), .B(n16316), .Z(n16136) );
  AND U16993 ( .A(n16317), .B(n16318), .Z(n16315) );
  AND U16994 ( .A(a[25]), .B(b[13]), .Z(n16314) );
  XOR U16995 ( .A(n16319), .B(n16141), .Z(n16143) );
  XOR U16996 ( .A(n16320), .B(n16321), .Z(n16141) );
  AND U16997 ( .A(n16322), .B(n16323), .Z(n16320) );
  AND U16998 ( .A(b[12]), .B(a[26]), .Z(n16319) );
  XOR U16999 ( .A(n16324), .B(n16146), .Z(n16148) );
  XOR U17000 ( .A(n16325), .B(n16326), .Z(n16146) );
  AND U17001 ( .A(n16327), .B(n16328), .Z(n16325) );
  AND U17002 ( .A(a[27]), .B(b[11]), .Z(n16324) );
  XOR U17003 ( .A(n16329), .B(n16151), .Z(n16153) );
  XOR U17004 ( .A(n16330), .B(n16331), .Z(n16151) );
  AND U17005 ( .A(n16332), .B(n16333), .Z(n16330) );
  AND U17006 ( .A(b[10]), .B(a[28]), .Z(n16329) );
  XOR U17007 ( .A(n16334), .B(n16156), .Z(n16158) );
  XOR U17008 ( .A(n16335), .B(n16336), .Z(n16156) );
  AND U17009 ( .A(n16337), .B(n16338), .Z(n16335) );
  AND U17010 ( .A(a[29]), .B(b[9]), .Z(n16334) );
  XOR U17011 ( .A(n16339), .B(n16161), .Z(n16163) );
  XOR U17012 ( .A(n16340), .B(n16341), .Z(n16161) );
  AND U17013 ( .A(n16342), .B(n16343), .Z(n16340) );
  AND U17014 ( .A(b[8]), .B(a[30]), .Z(n16339) );
  XOR U17015 ( .A(n16344), .B(n16166), .Z(n16168) );
  XOR U17016 ( .A(n16345), .B(n16346), .Z(n16166) );
  AND U17017 ( .A(n16347), .B(n16348), .Z(n16345) );
  AND U17018 ( .A(a[31]), .B(b[7]), .Z(n16344) );
  XOR U17019 ( .A(n16349), .B(n16171), .Z(n16173) );
  XOR U17020 ( .A(n16350), .B(n16351), .Z(n16171) );
  AND U17021 ( .A(n16352), .B(n16353), .Z(n16350) );
  AND U17022 ( .A(a[32]), .B(b[6]), .Z(n16349) );
  XOR U17023 ( .A(n16354), .B(n16176), .Z(n16178) );
  XOR U17024 ( .A(n16355), .B(n16356), .Z(n16176) );
  AND U17025 ( .A(n16357), .B(n16358), .Z(n16355) );
  AND U17026 ( .A(a[33]), .B(b[5]), .Z(n16354) );
  XOR U17027 ( .A(n16359), .B(n16360), .Z(n16200) );
  AND U17028 ( .A(n16195), .B(n16193), .Z(n16359) );
  AND U17029 ( .A(b[2]), .B(a[35]), .Z(n16361) );
  XNOR U17030 ( .A(n16362), .B(n16363), .Z(n16195) );
  XOR U17031 ( .A(n16364), .B(n16360), .Z(n16363) );
  XOR U17032 ( .A(n16365), .B(n16366), .Z(n16360) );
  NANDN U17033 ( .A(n16196), .B(n16197), .Z(n16366) );
  XNOR U17034 ( .A(n16367), .B(n16368), .Z(n16197) );
  XNOR U17035 ( .A(n16365), .B(n16369), .Z(n16368) );
  NAND U17036 ( .A(a[35]), .B(b[1]), .Z(n16370) );
  ANDN U17037 ( .B(n5377), .A(n5379), .Z(n16365) );
  NAND U17038 ( .A(a[35]), .B(b[0]), .Z(n5379) );
  XNOR U17039 ( .A(n16371), .B(n16372), .Z(n5377) );
  XOR U17040 ( .A(n16373), .B(n16181), .Z(n16183) );
  XOR U17041 ( .A(n16374), .B(n16375), .Z(n16181) );
  AND U17042 ( .A(n16362), .B(n16364), .Z(n16374) );
  XOR U17043 ( .A(n16357), .B(n16377), .Z(n16376) );
  XOR U17044 ( .A(n16352), .B(n16379), .Z(n16378) );
  XOR U17045 ( .A(n16347), .B(n16381), .Z(n16380) );
  XOR U17046 ( .A(n16342), .B(n16383), .Z(n16382) );
  XOR U17047 ( .A(n16337), .B(n16385), .Z(n16384) );
  XOR U17048 ( .A(n16332), .B(n16387), .Z(n16386) );
  XOR U17049 ( .A(n16327), .B(n16389), .Z(n16388) );
  XOR U17050 ( .A(n16322), .B(n16391), .Z(n16390) );
  XOR U17051 ( .A(n16317), .B(n16393), .Z(n16392) );
  XOR U17052 ( .A(n16312), .B(n16395), .Z(n16394) );
  XOR U17053 ( .A(n16307), .B(n16397), .Z(n16396) );
  XOR U17054 ( .A(n16302), .B(n16399), .Z(n16398) );
  XOR U17055 ( .A(n16297), .B(n16401), .Z(n16400) );
  XOR U17056 ( .A(n16292), .B(n16403), .Z(n16402) );
  XOR U17057 ( .A(n16287), .B(n16405), .Z(n16404) );
  XOR U17058 ( .A(n16282), .B(n16407), .Z(n16406) );
  XOR U17059 ( .A(n16277), .B(n16409), .Z(n16408) );
  XOR U17060 ( .A(n16272), .B(n16411), .Z(n16410) );
  XOR U17061 ( .A(n16267), .B(n16413), .Z(n16412) );
  XOR U17062 ( .A(n16262), .B(n16415), .Z(n16414) );
  XOR U17063 ( .A(n16257), .B(n16417), .Z(n16416) );
  XOR U17064 ( .A(n16252), .B(n16419), .Z(n16418) );
  XOR U17065 ( .A(n16247), .B(n16421), .Z(n16420) );
  XOR U17066 ( .A(n16242), .B(n16423), .Z(n16422) );
  XNOR U17067 ( .A(n16238), .B(n16425), .Z(n16424) );
  XOR U17068 ( .A(n16426), .B(n16427), .Z(n16238) );
  XOR U17069 ( .A(n16428), .B(n16429), .Z(n16427) );
  XNOR U17070 ( .A(n16430), .B(n16431), .Z(n16428) );
  XOR U17071 ( .A(n16432), .B(n16433), .Z(n16431) );
  AND U17072 ( .A(a[6]), .B(b[31]), .Z(n16433) );
  AND U17073 ( .A(a[7]), .B(b[30]), .Z(n16432) );
  XNOR U17074 ( .A(n16434), .B(n16430), .Z(n16426) );
  XNOR U17075 ( .A(n16435), .B(n16436), .Z(n16430) );
  ANDN U17076 ( .B(n16437), .A(n16438), .Z(n16435) );
  AND U17077 ( .A(a[8]), .B(b[29]), .Z(n16434) );
  XOR U17078 ( .A(n16439), .B(n16236), .Z(n16237) );
  IV U17079 ( .A(n16429), .Z(n16236) );
  XOR U17080 ( .A(n16440), .B(n16441), .Z(n16429) );
  AND U17081 ( .A(n16442), .B(n16443), .Z(n16440) );
  AND U17082 ( .A(a[9]), .B(b[28]), .Z(n16439) );
  XOR U17083 ( .A(n16444), .B(n16241), .Z(n16243) );
  IV U17084 ( .A(n16425), .Z(n16241) );
  XOR U17085 ( .A(n16445), .B(n16446), .Z(n16425) );
  AND U17086 ( .A(n16447), .B(n16448), .Z(n16445) );
  AND U17087 ( .A(a[10]), .B(b[27]), .Z(n16444) );
  XOR U17088 ( .A(n16449), .B(n16246), .Z(n16248) );
  IV U17089 ( .A(n16423), .Z(n16246) );
  XOR U17090 ( .A(n16450), .B(n16451), .Z(n16423) );
  AND U17091 ( .A(n16452), .B(n16453), .Z(n16450) );
  AND U17092 ( .A(a[11]), .B(b[26]), .Z(n16449) );
  XOR U17093 ( .A(n16454), .B(n16251), .Z(n16253) );
  IV U17094 ( .A(n16421), .Z(n16251) );
  XOR U17095 ( .A(n16455), .B(n16456), .Z(n16421) );
  AND U17096 ( .A(n16457), .B(n16458), .Z(n16455) );
  AND U17097 ( .A(a[12]), .B(b[25]), .Z(n16454) );
  XOR U17098 ( .A(n16459), .B(n16256), .Z(n16258) );
  IV U17099 ( .A(n16419), .Z(n16256) );
  XOR U17100 ( .A(n16460), .B(n16461), .Z(n16419) );
  AND U17101 ( .A(n16462), .B(n16463), .Z(n16460) );
  AND U17102 ( .A(a[13]), .B(b[24]), .Z(n16459) );
  XOR U17103 ( .A(n16464), .B(n16261), .Z(n16263) );
  IV U17104 ( .A(n16417), .Z(n16261) );
  XOR U17105 ( .A(n16465), .B(n16466), .Z(n16417) );
  AND U17106 ( .A(n16467), .B(n16468), .Z(n16465) );
  AND U17107 ( .A(a[14]), .B(b[23]), .Z(n16464) );
  XOR U17108 ( .A(n16469), .B(n16266), .Z(n16268) );
  IV U17109 ( .A(n16415), .Z(n16266) );
  XOR U17110 ( .A(n16470), .B(n16471), .Z(n16415) );
  AND U17111 ( .A(n16472), .B(n16473), .Z(n16470) );
  AND U17112 ( .A(a[15]), .B(b[22]), .Z(n16469) );
  XOR U17113 ( .A(n16474), .B(n16271), .Z(n16273) );
  IV U17114 ( .A(n16413), .Z(n16271) );
  XOR U17115 ( .A(n16475), .B(n16476), .Z(n16413) );
  AND U17116 ( .A(n16477), .B(n16478), .Z(n16475) );
  AND U17117 ( .A(a[16]), .B(b[21]), .Z(n16474) );
  XOR U17118 ( .A(n16479), .B(n16276), .Z(n16278) );
  IV U17119 ( .A(n16411), .Z(n16276) );
  XOR U17120 ( .A(n16480), .B(n16481), .Z(n16411) );
  AND U17121 ( .A(n16482), .B(n16483), .Z(n16480) );
  AND U17122 ( .A(a[17]), .B(b[20]), .Z(n16479) );
  XOR U17123 ( .A(n16484), .B(n16281), .Z(n16283) );
  IV U17124 ( .A(n16409), .Z(n16281) );
  XOR U17125 ( .A(n16485), .B(n16486), .Z(n16409) );
  AND U17126 ( .A(n16487), .B(n16488), .Z(n16485) );
  AND U17127 ( .A(a[18]), .B(b[19]), .Z(n16484) );
  XOR U17128 ( .A(n16489), .B(n16286), .Z(n16288) );
  IV U17129 ( .A(n16407), .Z(n16286) );
  XOR U17130 ( .A(n16490), .B(n16491), .Z(n16407) );
  AND U17131 ( .A(n16492), .B(n16493), .Z(n16490) );
  AND U17132 ( .A(a[19]), .B(b[18]), .Z(n16489) );
  XOR U17133 ( .A(n16494), .B(n16291), .Z(n16293) );
  IV U17134 ( .A(n16405), .Z(n16291) );
  XOR U17135 ( .A(n16495), .B(n16496), .Z(n16405) );
  AND U17136 ( .A(n16497), .B(n16498), .Z(n16495) );
  AND U17137 ( .A(b[17]), .B(a[20]), .Z(n16494) );
  XOR U17138 ( .A(n16499), .B(n16296), .Z(n16298) );
  IV U17139 ( .A(n16403), .Z(n16296) );
  XOR U17140 ( .A(n16500), .B(n16501), .Z(n16403) );
  AND U17141 ( .A(n16502), .B(n16503), .Z(n16500) );
  AND U17142 ( .A(a[21]), .B(b[16]), .Z(n16499) );
  XOR U17143 ( .A(n16504), .B(n16301), .Z(n16303) );
  IV U17144 ( .A(n16401), .Z(n16301) );
  XOR U17145 ( .A(n16505), .B(n16506), .Z(n16401) );
  AND U17146 ( .A(n16507), .B(n16508), .Z(n16505) );
  AND U17147 ( .A(b[15]), .B(a[22]), .Z(n16504) );
  XOR U17148 ( .A(n16509), .B(n16306), .Z(n16308) );
  IV U17149 ( .A(n16399), .Z(n16306) );
  XOR U17150 ( .A(n16510), .B(n16511), .Z(n16399) );
  AND U17151 ( .A(n16512), .B(n16513), .Z(n16510) );
  AND U17152 ( .A(a[23]), .B(b[14]), .Z(n16509) );
  XOR U17153 ( .A(n16514), .B(n16311), .Z(n16313) );
  IV U17154 ( .A(n16397), .Z(n16311) );
  XOR U17155 ( .A(n16515), .B(n16516), .Z(n16397) );
  AND U17156 ( .A(n16517), .B(n16518), .Z(n16515) );
  AND U17157 ( .A(b[13]), .B(a[24]), .Z(n16514) );
  XOR U17158 ( .A(n16519), .B(n16316), .Z(n16318) );
  IV U17159 ( .A(n16395), .Z(n16316) );
  XOR U17160 ( .A(n16520), .B(n16521), .Z(n16395) );
  AND U17161 ( .A(n16522), .B(n16523), .Z(n16520) );
  AND U17162 ( .A(a[25]), .B(b[12]), .Z(n16519) );
  XOR U17163 ( .A(n16524), .B(n16321), .Z(n16323) );
  IV U17164 ( .A(n16393), .Z(n16321) );
  XOR U17165 ( .A(n16525), .B(n16526), .Z(n16393) );
  AND U17166 ( .A(n16527), .B(n16528), .Z(n16525) );
  AND U17167 ( .A(b[11]), .B(a[26]), .Z(n16524) );
  XOR U17168 ( .A(n16529), .B(n16326), .Z(n16328) );
  IV U17169 ( .A(n16391), .Z(n16326) );
  XOR U17170 ( .A(n16530), .B(n16531), .Z(n16391) );
  AND U17171 ( .A(n16532), .B(n16533), .Z(n16530) );
  AND U17172 ( .A(a[27]), .B(b[10]), .Z(n16529) );
  XOR U17173 ( .A(n16534), .B(n16331), .Z(n16333) );
  IV U17174 ( .A(n16389), .Z(n16331) );
  XOR U17175 ( .A(n16535), .B(n16536), .Z(n16389) );
  AND U17176 ( .A(n16537), .B(n16538), .Z(n16535) );
  AND U17177 ( .A(b[9]), .B(a[28]), .Z(n16534) );
  XOR U17178 ( .A(n16539), .B(n16336), .Z(n16338) );
  IV U17179 ( .A(n16387), .Z(n16336) );
  XOR U17180 ( .A(n16540), .B(n16541), .Z(n16387) );
  AND U17181 ( .A(n16542), .B(n16543), .Z(n16540) );
  AND U17182 ( .A(a[29]), .B(b[8]), .Z(n16539) );
  XOR U17183 ( .A(n16544), .B(n16341), .Z(n16343) );
  IV U17184 ( .A(n16385), .Z(n16341) );
  XOR U17185 ( .A(n16545), .B(n16546), .Z(n16385) );
  AND U17186 ( .A(n16547), .B(n16548), .Z(n16545) );
  AND U17187 ( .A(b[7]), .B(a[30]), .Z(n16544) );
  XOR U17188 ( .A(n16549), .B(n16346), .Z(n16348) );
  IV U17189 ( .A(n16383), .Z(n16346) );
  XOR U17190 ( .A(n16550), .B(n16551), .Z(n16383) );
  AND U17191 ( .A(n16552), .B(n16553), .Z(n16550) );
  AND U17192 ( .A(a[31]), .B(b[6]), .Z(n16549) );
  XOR U17193 ( .A(n16554), .B(n16351), .Z(n16353) );
  IV U17194 ( .A(n16381), .Z(n16351) );
  XOR U17195 ( .A(n16555), .B(n16556), .Z(n16381) );
  AND U17196 ( .A(n16557), .B(n16558), .Z(n16555) );
  AND U17197 ( .A(a[32]), .B(b[5]), .Z(n16554) );
  XOR U17198 ( .A(n16559), .B(n16356), .Z(n16358) );
  IV U17199 ( .A(n16379), .Z(n16356) );
  XOR U17200 ( .A(n16560), .B(n16561), .Z(n16379) );
  AND U17201 ( .A(n16562), .B(n16563), .Z(n16560) );
  AND U17202 ( .A(a[33]), .B(b[4]), .Z(n16559) );
  XOR U17203 ( .A(n16564), .B(n16375), .Z(n16362) );
  IV U17204 ( .A(n16377), .Z(n16375) );
  XOR U17205 ( .A(n16565), .B(n16566), .Z(n16377) );
  AND U17206 ( .A(n16369), .B(n16367), .Z(n16565) );
  AND U17207 ( .A(b[2]), .B(a[34]), .Z(n16567) );
  XOR U17208 ( .A(n16562), .B(n16566), .Z(n16568) );
  XOR U17209 ( .A(n16569), .B(n16570), .Z(n16566) );
  NANDN U17210 ( .A(n16372), .B(n16371), .Z(n16570) );
  XOR U17211 ( .A(n16571), .B(n16572), .Z(n16371) );
  NAND U17212 ( .A(a[34]), .B(b[1]), .Z(n16572) );
  XOR U17213 ( .A(n16573), .B(n16574), .Z(n16372) );
  XOR U17214 ( .A(n16571), .B(n16575), .Z(n16574) );
  IV U17215 ( .A(n16569), .Z(n16571) );
  ANDN U17216 ( .B(n5382), .A(n5384), .Z(n16569) );
  NAND U17217 ( .A(a[34]), .B(b[0]), .Z(n5384) );
  XNOR U17218 ( .A(n16576), .B(n16577), .Z(n5382) );
  XOR U17219 ( .A(n16557), .B(n16561), .Z(n16578) );
  XOR U17220 ( .A(n16552), .B(n16556), .Z(n16579) );
  XOR U17221 ( .A(n16547), .B(n16551), .Z(n16580) );
  XOR U17222 ( .A(n16542), .B(n16546), .Z(n16581) );
  XOR U17223 ( .A(n16537), .B(n16541), .Z(n16582) );
  XOR U17224 ( .A(n16532), .B(n16536), .Z(n16583) );
  XOR U17225 ( .A(n16527), .B(n16531), .Z(n16584) );
  XOR U17226 ( .A(n16522), .B(n16526), .Z(n16585) );
  XOR U17227 ( .A(n16517), .B(n16521), .Z(n16586) );
  XOR U17228 ( .A(n16512), .B(n16516), .Z(n16587) );
  XOR U17229 ( .A(n16507), .B(n16511), .Z(n16588) );
  XOR U17230 ( .A(n16502), .B(n16506), .Z(n16589) );
  XOR U17231 ( .A(n16497), .B(n16501), .Z(n16590) );
  XOR U17232 ( .A(n16492), .B(n16496), .Z(n16591) );
  XOR U17233 ( .A(n16487), .B(n16491), .Z(n16592) );
  XOR U17234 ( .A(n16482), .B(n16486), .Z(n16593) );
  XOR U17235 ( .A(n16477), .B(n16481), .Z(n16594) );
  XOR U17236 ( .A(n16472), .B(n16476), .Z(n16595) );
  XOR U17237 ( .A(n16467), .B(n16471), .Z(n16596) );
  XOR U17238 ( .A(n16462), .B(n16466), .Z(n16597) );
  XOR U17239 ( .A(n16457), .B(n16461), .Z(n16598) );
  XOR U17240 ( .A(n16452), .B(n16456), .Z(n16599) );
  XOR U17241 ( .A(n16447), .B(n16451), .Z(n16600) );
  XOR U17242 ( .A(n16442), .B(n16446), .Z(n16601) );
  XNOR U17243 ( .A(n16438), .B(n16441), .Z(n16602) );
  XOR U17244 ( .A(n16603), .B(n16604), .Z(n16438) );
  XOR U17245 ( .A(n16605), .B(n16606), .Z(n16604) );
  XNOR U17246 ( .A(n16607), .B(n16608), .Z(n16605) );
  XOR U17247 ( .A(n16609), .B(n16610), .Z(n16608) );
  AND U17248 ( .A(a[6]), .B(b[30]), .Z(n16610) );
  AND U17249 ( .A(a[5]), .B(b[31]), .Z(n16609) );
  XNOR U17250 ( .A(n16611), .B(n16607), .Z(n16603) );
  XNOR U17251 ( .A(n16612), .B(n16613), .Z(n16607) );
  ANDN U17252 ( .B(n16614), .A(n16615), .Z(n16612) );
  AND U17253 ( .A(a[7]), .B(b[29]), .Z(n16611) );
  XOR U17254 ( .A(n16616), .B(n16436), .Z(n16437) );
  IV U17255 ( .A(n16606), .Z(n16436) );
  XOR U17256 ( .A(n16617), .B(n16618), .Z(n16606) );
  AND U17257 ( .A(n16619), .B(n16620), .Z(n16617) );
  AND U17258 ( .A(a[8]), .B(b[28]), .Z(n16616) );
  XOR U17259 ( .A(n16622), .B(n16623), .Z(n16441) );
  AND U17260 ( .A(n16624), .B(n16625), .Z(n16622) );
  AND U17261 ( .A(a[9]), .B(b[27]), .Z(n16621) );
  XOR U17262 ( .A(n16627), .B(n16628), .Z(n16446) );
  AND U17263 ( .A(n16629), .B(n16630), .Z(n16627) );
  AND U17264 ( .A(a[10]), .B(b[26]), .Z(n16626) );
  XOR U17265 ( .A(n16632), .B(n16633), .Z(n16451) );
  AND U17266 ( .A(n16634), .B(n16635), .Z(n16632) );
  AND U17267 ( .A(a[11]), .B(b[25]), .Z(n16631) );
  XOR U17268 ( .A(n16637), .B(n16638), .Z(n16456) );
  AND U17269 ( .A(n16639), .B(n16640), .Z(n16637) );
  AND U17270 ( .A(a[12]), .B(b[24]), .Z(n16636) );
  XOR U17271 ( .A(n16642), .B(n16643), .Z(n16461) );
  AND U17272 ( .A(n16644), .B(n16645), .Z(n16642) );
  AND U17273 ( .A(a[13]), .B(b[23]), .Z(n16641) );
  XOR U17274 ( .A(n16647), .B(n16648), .Z(n16466) );
  AND U17275 ( .A(n16649), .B(n16650), .Z(n16647) );
  AND U17276 ( .A(a[14]), .B(b[22]), .Z(n16646) );
  XOR U17277 ( .A(n16652), .B(n16653), .Z(n16471) );
  AND U17278 ( .A(n16654), .B(n16655), .Z(n16652) );
  AND U17279 ( .A(a[15]), .B(b[21]), .Z(n16651) );
  XOR U17280 ( .A(n16657), .B(n16658), .Z(n16476) );
  AND U17281 ( .A(n16659), .B(n16660), .Z(n16657) );
  AND U17282 ( .A(a[16]), .B(b[20]), .Z(n16656) );
  XOR U17283 ( .A(n16662), .B(n16663), .Z(n16481) );
  AND U17284 ( .A(n16664), .B(n16665), .Z(n16662) );
  AND U17285 ( .A(a[17]), .B(b[19]), .Z(n16661) );
  XOR U17286 ( .A(n16667), .B(n16668), .Z(n16486) );
  AND U17287 ( .A(n16669), .B(n16670), .Z(n16667) );
  AND U17288 ( .A(b[18]), .B(a[18]), .Z(n16666) );
  XOR U17289 ( .A(n16672), .B(n16673), .Z(n16491) );
  AND U17290 ( .A(n16674), .B(n16675), .Z(n16672) );
  AND U17291 ( .A(a[19]), .B(b[17]), .Z(n16671) );
  XOR U17292 ( .A(n16677), .B(n16678), .Z(n16496) );
  AND U17293 ( .A(n16679), .B(n16680), .Z(n16677) );
  AND U17294 ( .A(b[16]), .B(a[20]), .Z(n16676) );
  XOR U17295 ( .A(n16682), .B(n16683), .Z(n16501) );
  AND U17296 ( .A(n16684), .B(n16685), .Z(n16682) );
  AND U17297 ( .A(a[21]), .B(b[15]), .Z(n16681) );
  XOR U17298 ( .A(n16687), .B(n16688), .Z(n16506) );
  AND U17299 ( .A(n16689), .B(n16690), .Z(n16687) );
  AND U17300 ( .A(b[14]), .B(a[22]), .Z(n16686) );
  XOR U17301 ( .A(n16692), .B(n16693), .Z(n16511) );
  AND U17302 ( .A(n16694), .B(n16695), .Z(n16692) );
  AND U17303 ( .A(a[23]), .B(b[13]), .Z(n16691) );
  XOR U17304 ( .A(n16697), .B(n16698), .Z(n16516) );
  AND U17305 ( .A(n16699), .B(n16700), .Z(n16697) );
  AND U17306 ( .A(b[12]), .B(a[24]), .Z(n16696) );
  XOR U17307 ( .A(n16702), .B(n16703), .Z(n16521) );
  AND U17308 ( .A(n16704), .B(n16705), .Z(n16702) );
  AND U17309 ( .A(a[25]), .B(b[11]), .Z(n16701) );
  XOR U17310 ( .A(n16707), .B(n16708), .Z(n16526) );
  AND U17311 ( .A(n16709), .B(n16710), .Z(n16707) );
  AND U17312 ( .A(b[10]), .B(a[26]), .Z(n16706) );
  XOR U17313 ( .A(n16712), .B(n16713), .Z(n16531) );
  AND U17314 ( .A(n16714), .B(n16715), .Z(n16712) );
  AND U17315 ( .A(a[27]), .B(b[9]), .Z(n16711) );
  XOR U17316 ( .A(n16717), .B(n16718), .Z(n16536) );
  AND U17317 ( .A(n16719), .B(n16720), .Z(n16717) );
  AND U17318 ( .A(b[8]), .B(a[28]), .Z(n16716) );
  XOR U17319 ( .A(n16722), .B(n16723), .Z(n16541) );
  AND U17320 ( .A(n16724), .B(n16725), .Z(n16722) );
  AND U17321 ( .A(a[29]), .B(b[7]), .Z(n16721) );
  XOR U17322 ( .A(n16727), .B(n16728), .Z(n16546) );
  AND U17323 ( .A(n16729), .B(n16730), .Z(n16727) );
  AND U17324 ( .A(b[6]), .B(a[30]), .Z(n16726) );
  XOR U17325 ( .A(n16732), .B(n16733), .Z(n16551) );
  AND U17326 ( .A(n16734), .B(n16735), .Z(n16732) );
  AND U17327 ( .A(a[31]), .B(b[5]), .Z(n16731) );
  XOR U17328 ( .A(n16737), .B(n16738), .Z(n16556) );
  AND U17329 ( .A(n16739), .B(n16740), .Z(n16737) );
  AND U17330 ( .A(a[32]), .B(b[4]), .Z(n16736) );
  XOR U17331 ( .A(n16742), .B(n16743), .Z(n16561) );
  AND U17332 ( .A(n16575), .B(n16573), .Z(n16742) );
  AND U17333 ( .A(b[2]), .B(a[33]), .Z(n16744) );
  XOR U17334 ( .A(n16739), .B(n16743), .Z(n16745) );
  XOR U17335 ( .A(n16746), .B(n16747), .Z(n16743) );
  NANDN U17336 ( .A(n16577), .B(n16576), .Z(n16747) );
  XOR U17337 ( .A(n16748), .B(n16749), .Z(n16576) );
  NAND U17338 ( .A(a[33]), .B(b[1]), .Z(n16749) );
  XOR U17339 ( .A(n16750), .B(n16751), .Z(n16577) );
  XOR U17340 ( .A(n16748), .B(n16752), .Z(n16751) );
  IV U17341 ( .A(n16746), .Z(n16748) );
  ANDN U17342 ( .B(n5387), .A(n5389), .Z(n16746) );
  NAND U17343 ( .A(a[33]), .B(b[0]), .Z(n5389) );
  XNOR U17344 ( .A(n16753), .B(n16754), .Z(n5387) );
  XOR U17345 ( .A(n16734), .B(n16738), .Z(n16755) );
  XOR U17346 ( .A(n16729), .B(n16733), .Z(n16756) );
  XOR U17347 ( .A(n16724), .B(n16728), .Z(n16757) );
  XOR U17348 ( .A(n16719), .B(n16723), .Z(n16758) );
  XOR U17349 ( .A(n16714), .B(n16718), .Z(n16759) );
  XOR U17350 ( .A(n16709), .B(n16713), .Z(n16760) );
  XOR U17351 ( .A(n16704), .B(n16708), .Z(n16761) );
  XOR U17352 ( .A(n16699), .B(n16703), .Z(n16762) );
  XOR U17353 ( .A(n16694), .B(n16698), .Z(n16763) );
  XOR U17354 ( .A(n16689), .B(n16693), .Z(n16764) );
  XOR U17355 ( .A(n16684), .B(n16688), .Z(n16765) );
  XOR U17356 ( .A(n16679), .B(n16683), .Z(n16766) );
  XOR U17357 ( .A(n16674), .B(n16678), .Z(n16767) );
  XOR U17358 ( .A(n16669), .B(n16673), .Z(n16768) );
  XOR U17359 ( .A(n16664), .B(n16668), .Z(n16769) );
  XOR U17360 ( .A(n16659), .B(n16663), .Z(n16770) );
  XOR U17361 ( .A(n16654), .B(n16658), .Z(n16771) );
  XOR U17362 ( .A(n16649), .B(n16653), .Z(n16772) );
  XOR U17363 ( .A(n16644), .B(n16648), .Z(n16773) );
  XOR U17364 ( .A(n16639), .B(n16643), .Z(n16774) );
  XOR U17365 ( .A(n16634), .B(n16638), .Z(n16775) );
  XOR U17366 ( .A(n16629), .B(n16633), .Z(n16776) );
  XOR U17367 ( .A(n16624), .B(n16628), .Z(n16777) );
  XOR U17368 ( .A(n16619), .B(n16623), .Z(n16778) );
  XNOR U17369 ( .A(n16615), .B(n16618), .Z(n16779) );
  XOR U17370 ( .A(n16780), .B(n16781), .Z(n16615) );
  XOR U17371 ( .A(n16782), .B(n16783), .Z(n16781) );
  XOR U17372 ( .A(n16784), .B(n16785), .Z(n16782) );
  AND U17373 ( .A(a[6]), .B(b[29]), .Z(n16784) );
  XOR U17374 ( .A(n16785), .B(n16786), .Z(n16780) );
  XOR U17375 ( .A(n16787), .B(n16788), .Z(n16786) );
  AND U17376 ( .A(a[5]), .B(b[30]), .Z(n16788) );
  AND U17377 ( .A(a[4]), .B(b[31]), .Z(n16787) );
  XOR U17378 ( .A(n16789), .B(n16790), .Z(n16785) );
  ANDN U17379 ( .B(n16791), .A(n16792), .Z(n16789) );
  XOR U17380 ( .A(n16793), .B(n16613), .Z(n16614) );
  IV U17381 ( .A(n16783), .Z(n16613) );
  XOR U17382 ( .A(n16794), .B(n16795), .Z(n16783) );
  ANDN U17383 ( .B(n16796), .A(n16797), .Z(n16794) );
  AND U17384 ( .A(a[7]), .B(b[28]), .Z(n16793) );
  XOR U17385 ( .A(n16799), .B(n16800), .Z(n16618) );
  AND U17386 ( .A(n16801), .B(n16802), .Z(n16799) );
  AND U17387 ( .A(a[8]), .B(b[27]), .Z(n16798) );
  XOR U17388 ( .A(n16804), .B(n16805), .Z(n16623) );
  AND U17389 ( .A(n16806), .B(n16807), .Z(n16804) );
  AND U17390 ( .A(a[9]), .B(b[26]), .Z(n16803) );
  XOR U17391 ( .A(n16809), .B(n16810), .Z(n16628) );
  AND U17392 ( .A(n16811), .B(n16812), .Z(n16809) );
  AND U17393 ( .A(a[10]), .B(b[25]), .Z(n16808) );
  XOR U17394 ( .A(n16814), .B(n16815), .Z(n16633) );
  AND U17395 ( .A(n16816), .B(n16817), .Z(n16814) );
  AND U17396 ( .A(a[11]), .B(b[24]), .Z(n16813) );
  XOR U17397 ( .A(n16819), .B(n16820), .Z(n16638) );
  AND U17398 ( .A(n16821), .B(n16822), .Z(n16819) );
  AND U17399 ( .A(a[12]), .B(b[23]), .Z(n16818) );
  XOR U17400 ( .A(n16824), .B(n16825), .Z(n16643) );
  AND U17401 ( .A(n16826), .B(n16827), .Z(n16824) );
  AND U17402 ( .A(a[13]), .B(b[22]), .Z(n16823) );
  XOR U17403 ( .A(n16829), .B(n16830), .Z(n16648) );
  AND U17404 ( .A(n16831), .B(n16832), .Z(n16829) );
  AND U17405 ( .A(a[14]), .B(b[21]), .Z(n16828) );
  XOR U17406 ( .A(n16834), .B(n16835), .Z(n16653) );
  AND U17407 ( .A(n16836), .B(n16837), .Z(n16834) );
  AND U17408 ( .A(a[15]), .B(b[20]), .Z(n16833) );
  XOR U17409 ( .A(n16839), .B(n16840), .Z(n16658) );
  AND U17410 ( .A(n16841), .B(n16842), .Z(n16839) );
  AND U17411 ( .A(a[16]), .B(b[19]), .Z(n16838) );
  XOR U17412 ( .A(n16844), .B(n16845), .Z(n16663) );
  AND U17413 ( .A(n16846), .B(n16847), .Z(n16844) );
  AND U17414 ( .A(a[17]), .B(b[18]), .Z(n16843) );
  XOR U17415 ( .A(n16849), .B(n16850), .Z(n16668) );
  AND U17416 ( .A(n16851), .B(n16852), .Z(n16849) );
  AND U17417 ( .A(b[17]), .B(a[18]), .Z(n16848) );
  XOR U17418 ( .A(n16854), .B(n16855), .Z(n16673) );
  AND U17419 ( .A(n16856), .B(n16857), .Z(n16854) );
  AND U17420 ( .A(a[19]), .B(b[16]), .Z(n16853) );
  XOR U17421 ( .A(n16859), .B(n16860), .Z(n16678) );
  AND U17422 ( .A(n16861), .B(n16862), .Z(n16859) );
  AND U17423 ( .A(b[15]), .B(a[20]), .Z(n16858) );
  XOR U17424 ( .A(n16864), .B(n16865), .Z(n16683) );
  AND U17425 ( .A(n16866), .B(n16867), .Z(n16864) );
  AND U17426 ( .A(a[21]), .B(b[14]), .Z(n16863) );
  XOR U17427 ( .A(n16869), .B(n16870), .Z(n16688) );
  AND U17428 ( .A(n16871), .B(n16872), .Z(n16869) );
  AND U17429 ( .A(b[13]), .B(a[22]), .Z(n16868) );
  XOR U17430 ( .A(n16874), .B(n16875), .Z(n16693) );
  AND U17431 ( .A(n16876), .B(n16877), .Z(n16874) );
  AND U17432 ( .A(a[23]), .B(b[12]), .Z(n16873) );
  XOR U17433 ( .A(n16879), .B(n16880), .Z(n16698) );
  AND U17434 ( .A(n16881), .B(n16882), .Z(n16879) );
  AND U17435 ( .A(b[11]), .B(a[24]), .Z(n16878) );
  XOR U17436 ( .A(n16884), .B(n16885), .Z(n16703) );
  AND U17437 ( .A(n16886), .B(n16887), .Z(n16884) );
  AND U17438 ( .A(a[25]), .B(b[10]), .Z(n16883) );
  XOR U17439 ( .A(n16889), .B(n16890), .Z(n16708) );
  AND U17440 ( .A(n16891), .B(n16892), .Z(n16889) );
  AND U17441 ( .A(b[9]), .B(a[26]), .Z(n16888) );
  XOR U17442 ( .A(n16894), .B(n16895), .Z(n16713) );
  AND U17443 ( .A(n16896), .B(n16897), .Z(n16894) );
  AND U17444 ( .A(a[27]), .B(b[8]), .Z(n16893) );
  XOR U17445 ( .A(n16899), .B(n16900), .Z(n16718) );
  AND U17446 ( .A(n16901), .B(n16902), .Z(n16899) );
  AND U17447 ( .A(b[7]), .B(a[28]), .Z(n16898) );
  XOR U17448 ( .A(n16904), .B(n16905), .Z(n16723) );
  AND U17449 ( .A(n16906), .B(n16907), .Z(n16904) );
  AND U17450 ( .A(a[29]), .B(b[6]), .Z(n16903) );
  XOR U17451 ( .A(n16909), .B(n16910), .Z(n16728) );
  AND U17452 ( .A(n16911), .B(n16912), .Z(n16909) );
  AND U17453 ( .A(b[5]), .B(a[30]), .Z(n16908) );
  XOR U17454 ( .A(n16914), .B(n16915), .Z(n16733) );
  AND U17455 ( .A(n16916), .B(n16917), .Z(n16914) );
  AND U17456 ( .A(a[31]), .B(b[4]), .Z(n16913) );
  XOR U17457 ( .A(n16919), .B(n16920), .Z(n16738) );
  AND U17458 ( .A(n16752), .B(n16750), .Z(n16919) );
  AND U17459 ( .A(b[2]), .B(a[32]), .Z(n16921) );
  XOR U17460 ( .A(n16916), .B(n16920), .Z(n16922) );
  XOR U17461 ( .A(n16923), .B(n16924), .Z(n16920) );
  NANDN U17462 ( .A(n16754), .B(n16753), .Z(n16924) );
  XOR U17463 ( .A(n16925), .B(n16926), .Z(n16753) );
  NAND U17464 ( .A(a[32]), .B(b[1]), .Z(n16926) );
  XOR U17465 ( .A(n16927), .B(n16928), .Z(n16754) );
  XOR U17466 ( .A(n16925), .B(n16929), .Z(n16928) );
  IV U17467 ( .A(n16923), .Z(n16925) );
  ANDN U17468 ( .B(n5392), .A(n5394), .Z(n16923) );
  NAND U17469 ( .A(a[32]), .B(b[0]), .Z(n5394) );
  XNOR U17470 ( .A(n16930), .B(n16931), .Z(n5392) );
  XOR U17471 ( .A(n16911), .B(n16915), .Z(n16932) );
  XOR U17472 ( .A(n16906), .B(n16910), .Z(n16933) );
  XOR U17473 ( .A(n16901), .B(n16905), .Z(n16934) );
  XOR U17474 ( .A(n16896), .B(n16900), .Z(n16935) );
  XOR U17475 ( .A(n16891), .B(n16895), .Z(n16936) );
  XOR U17476 ( .A(n16886), .B(n16890), .Z(n16937) );
  XOR U17477 ( .A(n16881), .B(n16885), .Z(n16938) );
  XOR U17478 ( .A(n16876), .B(n16880), .Z(n16939) );
  XOR U17479 ( .A(n16871), .B(n16875), .Z(n16940) );
  XOR U17480 ( .A(n16866), .B(n16870), .Z(n16941) );
  XOR U17481 ( .A(n16861), .B(n16865), .Z(n16942) );
  XOR U17482 ( .A(n16856), .B(n16860), .Z(n16943) );
  XOR U17483 ( .A(n16851), .B(n16855), .Z(n16944) );
  XOR U17484 ( .A(n16846), .B(n16850), .Z(n16945) );
  XOR U17485 ( .A(n16841), .B(n16845), .Z(n16946) );
  XOR U17486 ( .A(n16836), .B(n16840), .Z(n16947) );
  XOR U17487 ( .A(n16831), .B(n16835), .Z(n16948) );
  XOR U17488 ( .A(n16826), .B(n16830), .Z(n16949) );
  XOR U17489 ( .A(n16821), .B(n16825), .Z(n16950) );
  XOR U17490 ( .A(n16816), .B(n16820), .Z(n16951) );
  XOR U17491 ( .A(n16811), .B(n16815), .Z(n16952) );
  XOR U17492 ( .A(n16806), .B(n16810), .Z(n16953) );
  XOR U17493 ( .A(n16801), .B(n16805), .Z(n16954) );
  XNOR U17494 ( .A(n16797), .B(n16800), .Z(n16955) );
  XNOR U17495 ( .A(n16792), .B(n16956), .Z(n16797) );
  XOR U17496 ( .A(n16791), .B(n16795), .Z(n16956) );
  XOR U17497 ( .A(n16957), .B(n16790), .Z(n16791) );
  AND U17498 ( .A(a[6]), .B(b[28]), .Z(n16957) );
  XOR U17499 ( .A(n16958), .B(n16959), .Z(n16792) );
  XOR U17500 ( .A(n16790), .B(n16960), .Z(n16959) );
  XOR U17501 ( .A(n16961), .B(n16962), .Z(n16960) );
  XOR U17502 ( .A(n16963), .B(n16964), .Z(n16962) );
  NAND U17503 ( .A(a[4]), .B(b[30]), .Z(n16964) );
  AND U17504 ( .A(a[3]), .B(b[31]), .Z(n16963) );
  XOR U17505 ( .A(n16965), .B(n16966), .Z(n16790) );
  AND U17506 ( .A(n16967), .B(n16968), .Z(n16965) );
  XOR U17507 ( .A(n16969), .B(n16961), .Z(n16958) );
  XOR U17508 ( .A(n16970), .B(n16971), .Z(n16961) );
  ANDN U17509 ( .B(n16972), .A(n16973), .Z(n16970) );
  AND U17510 ( .A(a[5]), .B(b[29]), .Z(n16969) );
  XOR U17511 ( .A(n16975), .B(n16976), .Z(n16795) );
  AND U17512 ( .A(n16977), .B(n16978), .Z(n16975) );
  AND U17513 ( .A(a[7]), .B(b[27]), .Z(n16974) );
  XOR U17514 ( .A(n16980), .B(n16981), .Z(n16800) );
  AND U17515 ( .A(n16982), .B(n16983), .Z(n16980) );
  AND U17516 ( .A(a[8]), .B(b[26]), .Z(n16979) );
  XOR U17517 ( .A(n16985), .B(n16986), .Z(n16805) );
  AND U17518 ( .A(n16987), .B(n16988), .Z(n16985) );
  AND U17519 ( .A(a[9]), .B(b[25]), .Z(n16984) );
  XOR U17520 ( .A(n16990), .B(n16991), .Z(n16810) );
  AND U17521 ( .A(n16992), .B(n16993), .Z(n16990) );
  AND U17522 ( .A(a[10]), .B(b[24]), .Z(n16989) );
  XOR U17523 ( .A(n16995), .B(n16996), .Z(n16815) );
  AND U17524 ( .A(n16997), .B(n16998), .Z(n16995) );
  AND U17525 ( .A(a[11]), .B(b[23]), .Z(n16994) );
  XOR U17526 ( .A(n17000), .B(n17001), .Z(n16820) );
  AND U17527 ( .A(n17002), .B(n17003), .Z(n17000) );
  AND U17528 ( .A(a[12]), .B(b[22]), .Z(n16999) );
  XOR U17529 ( .A(n17005), .B(n17006), .Z(n16825) );
  AND U17530 ( .A(n17007), .B(n17008), .Z(n17005) );
  AND U17531 ( .A(a[13]), .B(b[21]), .Z(n17004) );
  XOR U17532 ( .A(n17010), .B(n17011), .Z(n16830) );
  AND U17533 ( .A(n17012), .B(n17013), .Z(n17010) );
  AND U17534 ( .A(a[14]), .B(b[20]), .Z(n17009) );
  XOR U17535 ( .A(n17015), .B(n17016), .Z(n16835) );
  AND U17536 ( .A(n17017), .B(n17018), .Z(n17015) );
  AND U17537 ( .A(a[15]), .B(b[19]), .Z(n17014) );
  XOR U17538 ( .A(n17020), .B(n17021), .Z(n16840) );
  AND U17539 ( .A(n17022), .B(n17023), .Z(n17020) );
  AND U17540 ( .A(a[16]), .B(b[18]), .Z(n17019) );
  XOR U17541 ( .A(n17025), .B(n17026), .Z(n16845) );
  AND U17542 ( .A(n17027), .B(n17028), .Z(n17025) );
  AND U17543 ( .A(a[17]), .B(b[17]), .Z(n17024) );
  XOR U17544 ( .A(n17030), .B(n17031), .Z(n16850) );
  AND U17545 ( .A(n17032), .B(n17033), .Z(n17030) );
  AND U17546 ( .A(b[16]), .B(a[18]), .Z(n17029) );
  XOR U17547 ( .A(n17035), .B(n17036), .Z(n16855) );
  AND U17548 ( .A(n17037), .B(n17038), .Z(n17035) );
  AND U17549 ( .A(a[19]), .B(b[15]), .Z(n17034) );
  XOR U17550 ( .A(n17040), .B(n17041), .Z(n16860) );
  AND U17551 ( .A(n17042), .B(n17043), .Z(n17040) );
  AND U17552 ( .A(b[14]), .B(a[20]), .Z(n17039) );
  XOR U17553 ( .A(n17045), .B(n17046), .Z(n16865) );
  AND U17554 ( .A(n17047), .B(n17048), .Z(n17045) );
  AND U17555 ( .A(a[21]), .B(b[13]), .Z(n17044) );
  XOR U17556 ( .A(n17050), .B(n17051), .Z(n16870) );
  AND U17557 ( .A(n17052), .B(n17053), .Z(n17050) );
  AND U17558 ( .A(b[12]), .B(a[22]), .Z(n17049) );
  XOR U17559 ( .A(n17055), .B(n17056), .Z(n16875) );
  AND U17560 ( .A(n17057), .B(n17058), .Z(n17055) );
  AND U17561 ( .A(a[23]), .B(b[11]), .Z(n17054) );
  XOR U17562 ( .A(n17060), .B(n17061), .Z(n16880) );
  AND U17563 ( .A(n17062), .B(n17063), .Z(n17060) );
  AND U17564 ( .A(b[10]), .B(a[24]), .Z(n17059) );
  XOR U17565 ( .A(n17065), .B(n17066), .Z(n16885) );
  AND U17566 ( .A(n17067), .B(n17068), .Z(n17065) );
  AND U17567 ( .A(a[25]), .B(b[9]), .Z(n17064) );
  XOR U17568 ( .A(n17070), .B(n17071), .Z(n16890) );
  AND U17569 ( .A(n17072), .B(n17073), .Z(n17070) );
  AND U17570 ( .A(b[8]), .B(a[26]), .Z(n17069) );
  XOR U17571 ( .A(n17075), .B(n17076), .Z(n16895) );
  AND U17572 ( .A(n17077), .B(n17078), .Z(n17075) );
  AND U17573 ( .A(a[27]), .B(b[7]), .Z(n17074) );
  XOR U17574 ( .A(n17080), .B(n17081), .Z(n16900) );
  AND U17575 ( .A(n17082), .B(n17083), .Z(n17080) );
  AND U17576 ( .A(b[6]), .B(a[28]), .Z(n17079) );
  XOR U17577 ( .A(n17085), .B(n17086), .Z(n16905) );
  AND U17578 ( .A(n17087), .B(n17088), .Z(n17085) );
  AND U17579 ( .A(a[29]), .B(b[5]), .Z(n17084) );
  XOR U17580 ( .A(n17090), .B(n17091), .Z(n16910) );
  AND U17581 ( .A(n17092), .B(n17093), .Z(n17090) );
  AND U17582 ( .A(b[4]), .B(a[30]), .Z(n17089) );
  XOR U17583 ( .A(n17095), .B(n17096), .Z(n16915) );
  AND U17584 ( .A(n16929), .B(n16927), .Z(n17095) );
  AND U17585 ( .A(b[2]), .B(a[31]), .Z(n17097) );
  XOR U17586 ( .A(n17092), .B(n17096), .Z(n17098) );
  XOR U17587 ( .A(n17099), .B(n17100), .Z(n17096) );
  NANDN U17588 ( .A(n16931), .B(n16930), .Z(n17100) );
  XOR U17589 ( .A(n17101), .B(n17102), .Z(n16930) );
  NAND U17590 ( .A(a[31]), .B(b[1]), .Z(n17102) );
  XOR U17591 ( .A(n17103), .B(n17104), .Z(n16931) );
  XOR U17592 ( .A(n17101), .B(n17105), .Z(n17104) );
  IV U17593 ( .A(n17099), .Z(n17101) );
  ANDN U17594 ( .B(n17106), .A(n17107), .Z(n17099) );
  XOR U17595 ( .A(n17087), .B(n17091), .Z(n17108) );
  XOR U17596 ( .A(n17082), .B(n17086), .Z(n17109) );
  XOR U17597 ( .A(n17077), .B(n17081), .Z(n17110) );
  XOR U17598 ( .A(n17072), .B(n17076), .Z(n17111) );
  XOR U17599 ( .A(n17067), .B(n17071), .Z(n17112) );
  XOR U17600 ( .A(n17062), .B(n17066), .Z(n17113) );
  XOR U17601 ( .A(n17057), .B(n17061), .Z(n17114) );
  XOR U17602 ( .A(n17052), .B(n17056), .Z(n17115) );
  XOR U17603 ( .A(n17047), .B(n17051), .Z(n17116) );
  XOR U17604 ( .A(n17042), .B(n17046), .Z(n17117) );
  XOR U17605 ( .A(n17037), .B(n17041), .Z(n17118) );
  XOR U17606 ( .A(n17032), .B(n17036), .Z(n17119) );
  XOR U17607 ( .A(n17027), .B(n17031), .Z(n17120) );
  XOR U17608 ( .A(n17022), .B(n17026), .Z(n17121) );
  XOR U17609 ( .A(n17017), .B(n17021), .Z(n17122) );
  XOR U17610 ( .A(n17012), .B(n17016), .Z(n17123) );
  XOR U17611 ( .A(n17007), .B(n17011), .Z(n17124) );
  XOR U17612 ( .A(n17002), .B(n17006), .Z(n17125) );
  XOR U17613 ( .A(n16997), .B(n17001), .Z(n17126) );
  XOR U17614 ( .A(n16992), .B(n16996), .Z(n17127) );
  XOR U17615 ( .A(n16987), .B(n16991), .Z(n17128) );
  XOR U17616 ( .A(n16982), .B(n16986), .Z(n17129) );
  XOR U17617 ( .A(n16977), .B(n16981), .Z(n17130) );
  XOR U17618 ( .A(n16967), .B(n16976), .Z(n17131) );
  XOR U17619 ( .A(n17132), .B(n16966), .Z(n16967) );
  AND U17620 ( .A(a[6]), .B(b[27]), .Z(n17132) );
  XOR U17621 ( .A(n16966), .B(n16973), .Z(n17133) );
  XOR U17622 ( .A(n17134), .B(n17135), .Z(n16973) );
  XOR U17623 ( .A(n16971), .B(n17136), .Z(n17135) );
  XOR U17624 ( .A(n17137), .B(n17138), .Z(n17136) );
  XOR U17625 ( .A(n17139), .B(n17140), .Z(n17138) );
  NAND U17626 ( .A(a[3]), .B(b[30]), .Z(n17140) );
  AND U17627 ( .A(a[2]), .B(b[31]), .Z(n17139) );
  XOR U17628 ( .A(n17141), .B(n17137), .Z(n17134) );
  XOR U17629 ( .A(n17142), .B(n17143), .Z(n17137) );
  ANDN U17630 ( .B(n17144), .A(n17145), .Z(n17142) );
  AND U17631 ( .A(a[4]), .B(b[29]), .Z(n17141) );
  XOR U17632 ( .A(n17146), .B(n17147), .Z(n16966) );
  AND U17633 ( .A(n17148), .B(n17149), .Z(n17146) );
  XOR U17634 ( .A(n17150), .B(n16971), .Z(n16972) );
  XOR U17635 ( .A(n17151), .B(n17152), .Z(n16971) );
  AND U17636 ( .A(n17153), .B(n17154), .Z(n17151) );
  AND U17637 ( .A(a[5]), .B(b[28]), .Z(n17150) );
  XNOR U17638 ( .A(n17156), .B(n17157), .Z(n16976) );
  AND U17639 ( .A(n17158), .B(n17159), .Z(n17156) );
  AND U17640 ( .A(a[7]), .B(b[26]), .Z(n17155) );
  XNOR U17641 ( .A(n17161), .B(n17162), .Z(n16981) );
  AND U17642 ( .A(n17163), .B(n17164), .Z(n17161) );
  AND U17643 ( .A(a[8]), .B(b[25]), .Z(n17160) );
  XNOR U17644 ( .A(n17166), .B(n17167), .Z(n16986) );
  AND U17645 ( .A(n17168), .B(n17169), .Z(n17166) );
  AND U17646 ( .A(a[9]), .B(b[24]), .Z(n17165) );
  XNOR U17647 ( .A(n17171), .B(n17172), .Z(n16991) );
  AND U17648 ( .A(n17173), .B(n17174), .Z(n17171) );
  AND U17649 ( .A(a[10]), .B(b[23]), .Z(n17170) );
  XNOR U17650 ( .A(n17176), .B(n17177), .Z(n16996) );
  AND U17651 ( .A(n17178), .B(n17179), .Z(n17176) );
  AND U17652 ( .A(a[11]), .B(b[22]), .Z(n17175) );
  XNOR U17653 ( .A(n17181), .B(n17182), .Z(n17001) );
  AND U17654 ( .A(n17183), .B(n17184), .Z(n17181) );
  AND U17655 ( .A(a[12]), .B(b[21]), .Z(n17180) );
  XNOR U17656 ( .A(n17186), .B(n17187), .Z(n17006) );
  AND U17657 ( .A(n17188), .B(n17189), .Z(n17186) );
  AND U17658 ( .A(a[13]), .B(b[20]), .Z(n17185) );
  XNOR U17659 ( .A(n17191), .B(n17192), .Z(n17011) );
  AND U17660 ( .A(n17193), .B(n17194), .Z(n17191) );
  AND U17661 ( .A(a[14]), .B(b[19]), .Z(n17190) );
  XNOR U17662 ( .A(n17196), .B(n17197), .Z(n17016) );
  AND U17663 ( .A(n17198), .B(n17199), .Z(n17196) );
  AND U17664 ( .A(a[15]), .B(b[18]), .Z(n17195) );
  XNOR U17665 ( .A(n17201), .B(n17202), .Z(n17021) );
  AND U17666 ( .A(n17203), .B(n17204), .Z(n17201) );
  AND U17667 ( .A(a[16]), .B(b[17]), .Z(n17200) );
  XNOR U17668 ( .A(n17206), .B(n17207), .Z(n17026) );
  AND U17669 ( .A(n17208), .B(n17209), .Z(n17206) );
  AND U17670 ( .A(a[17]), .B(b[16]), .Z(n17205) );
  XNOR U17671 ( .A(n17211), .B(n17212), .Z(n17031) );
  AND U17672 ( .A(n17213), .B(n17214), .Z(n17211) );
  AND U17673 ( .A(b[15]), .B(a[18]), .Z(n17210) );
  XNOR U17674 ( .A(n17216), .B(n17217), .Z(n17036) );
  AND U17675 ( .A(n17218), .B(n17219), .Z(n17216) );
  AND U17676 ( .A(a[19]), .B(b[14]), .Z(n17215) );
  XNOR U17677 ( .A(n17221), .B(n17222), .Z(n17041) );
  AND U17678 ( .A(n17223), .B(n17224), .Z(n17221) );
  AND U17679 ( .A(b[13]), .B(a[20]), .Z(n17220) );
  XNOR U17680 ( .A(n17226), .B(n17227), .Z(n17046) );
  AND U17681 ( .A(n17228), .B(n17229), .Z(n17226) );
  AND U17682 ( .A(a[21]), .B(b[12]), .Z(n17225) );
  XNOR U17683 ( .A(n17231), .B(n17232), .Z(n17051) );
  AND U17684 ( .A(n17233), .B(n17234), .Z(n17231) );
  AND U17685 ( .A(b[11]), .B(a[22]), .Z(n17230) );
  XNOR U17686 ( .A(n17236), .B(n17237), .Z(n17056) );
  AND U17687 ( .A(n17238), .B(n17239), .Z(n17236) );
  AND U17688 ( .A(a[23]), .B(b[10]), .Z(n17235) );
  XNOR U17689 ( .A(n17241), .B(n17242), .Z(n17061) );
  AND U17690 ( .A(n17243), .B(n17244), .Z(n17241) );
  AND U17691 ( .A(b[9]), .B(a[24]), .Z(n17240) );
  XNOR U17692 ( .A(n17246), .B(n17247), .Z(n17066) );
  AND U17693 ( .A(n17248), .B(n17249), .Z(n17246) );
  AND U17694 ( .A(a[25]), .B(b[8]), .Z(n17245) );
  XNOR U17695 ( .A(n17251), .B(n17252), .Z(n17071) );
  AND U17696 ( .A(n17253), .B(n17254), .Z(n17251) );
  AND U17697 ( .A(b[7]), .B(a[26]), .Z(n17250) );
  XNOR U17698 ( .A(n17256), .B(n17257), .Z(n17076) );
  AND U17699 ( .A(n17258), .B(n17259), .Z(n17256) );
  AND U17700 ( .A(a[27]), .B(b[6]), .Z(n17255) );
  XNOR U17701 ( .A(n17261), .B(n17262), .Z(n17081) );
  AND U17702 ( .A(n17263), .B(n17264), .Z(n17261) );
  AND U17703 ( .A(b[5]), .B(a[28]), .Z(n17260) );
  XNOR U17704 ( .A(n17266), .B(n17267), .Z(n17086) );
  AND U17705 ( .A(n17268), .B(n17269), .Z(n17266) );
  AND U17706 ( .A(a[29]), .B(b[4]), .Z(n17265) );
  XOR U17707 ( .A(n17271), .B(n17272), .Z(n17091) );
  AND U17708 ( .A(n17105), .B(n17103), .Z(n17271) );
  AND U17709 ( .A(b[2]), .B(a[30]), .Z(n17273) );
  XOR U17710 ( .A(n17268), .B(n17272), .Z(n17274) );
  XOR U17711 ( .A(n17275), .B(n17276), .Z(n17272) );
  NANDN U17712 ( .A(n17277), .B(n17278), .Z(n17276) );
  XNOR U17713 ( .A(n17263), .B(n17267), .Z(n17279) );
  XNOR U17714 ( .A(n17258), .B(n17262), .Z(n17280) );
  XNOR U17715 ( .A(n17253), .B(n17257), .Z(n17281) );
  XNOR U17716 ( .A(n17248), .B(n17252), .Z(n17282) );
  XNOR U17717 ( .A(n17243), .B(n17247), .Z(n17283) );
  XNOR U17718 ( .A(n17238), .B(n17242), .Z(n17284) );
  XNOR U17719 ( .A(n17233), .B(n17237), .Z(n17285) );
  XNOR U17720 ( .A(n17228), .B(n17232), .Z(n17286) );
  XNOR U17721 ( .A(n17223), .B(n17227), .Z(n17287) );
  XNOR U17722 ( .A(n17218), .B(n17222), .Z(n17288) );
  XNOR U17723 ( .A(n17213), .B(n17217), .Z(n17289) );
  XNOR U17724 ( .A(n17208), .B(n17212), .Z(n17290) );
  XNOR U17725 ( .A(n17203), .B(n17207), .Z(n17291) );
  XNOR U17726 ( .A(n17198), .B(n17202), .Z(n17292) );
  XNOR U17727 ( .A(n17193), .B(n17197), .Z(n17293) );
  XNOR U17728 ( .A(n17188), .B(n17192), .Z(n17294) );
  XNOR U17729 ( .A(n17183), .B(n17187), .Z(n17295) );
  XNOR U17730 ( .A(n17178), .B(n17182), .Z(n17296) );
  XNOR U17731 ( .A(n17173), .B(n17177), .Z(n17297) );
  XNOR U17732 ( .A(n17168), .B(n17172), .Z(n17298) );
  XNOR U17733 ( .A(n17163), .B(n17167), .Z(n17299) );
  XNOR U17734 ( .A(n17158), .B(n17162), .Z(n17300) );
  XNOR U17735 ( .A(n17148), .B(n17157), .Z(n17301) );
  XOR U17736 ( .A(n17302), .B(n17147), .Z(n17148) );
  AND U17737 ( .A(a[6]), .B(b[26]), .Z(n17302) );
  XNOR U17738 ( .A(n17147), .B(n17153), .Z(n17303) );
  XOR U17739 ( .A(n17152), .B(n17145), .Z(n17304) );
  XOR U17740 ( .A(n17305), .B(n17306), .Z(n17145) );
  XOR U17741 ( .A(n17143), .B(n17307), .Z(n17306) );
  XOR U17742 ( .A(n17308), .B(n17309), .Z(n17307) );
  XOR U17743 ( .A(n17310), .B(n17311), .Z(n17309) );
  NAND U17744 ( .A(a[2]), .B(b[30]), .Z(n17311) );
  AND U17745 ( .A(a[1]), .B(b[31]), .Z(n17310) );
  XOR U17746 ( .A(n17312), .B(n17308), .Z(n17305) );
  XOR U17747 ( .A(n17313), .B(n17314), .Z(n17308) );
  ANDN U17748 ( .B(n17315), .A(n17316), .Z(n17313) );
  AND U17749 ( .A(a[3]), .B(b[29]), .Z(n17312) );
  XOR U17750 ( .A(n17317), .B(n17143), .Z(n17144) );
  XOR U17751 ( .A(n17318), .B(n17319), .Z(n17143) );
  AND U17752 ( .A(n17320), .B(n17321), .Z(n17318) );
  AND U17753 ( .A(a[4]), .B(b[28]), .Z(n17317) );
  XOR U17754 ( .A(n17322), .B(n17323), .Z(n17147) );
  AND U17755 ( .A(n17324), .B(n17325), .Z(n17322) );
  XOR U17756 ( .A(n17326), .B(n17152), .Z(n17154) );
  XOR U17757 ( .A(n17327), .B(n17328), .Z(n17152) );
  AND U17758 ( .A(n17329), .B(n17330), .Z(n17327) );
  AND U17759 ( .A(a[5]), .B(b[27]), .Z(n17326) );
  XOR U17760 ( .A(n17331), .B(n17157), .Z(n17159) );
  XOR U17761 ( .A(n17332), .B(n17333), .Z(n17157) );
  AND U17762 ( .A(n17334), .B(n17335), .Z(n17332) );
  AND U17763 ( .A(a[7]), .B(b[25]), .Z(n17331) );
  XOR U17764 ( .A(n17336), .B(n17162), .Z(n17164) );
  XOR U17765 ( .A(n17337), .B(n17338), .Z(n17162) );
  AND U17766 ( .A(n17339), .B(n17340), .Z(n17337) );
  AND U17767 ( .A(a[8]), .B(b[24]), .Z(n17336) );
  XOR U17768 ( .A(n17341), .B(n17167), .Z(n17169) );
  XOR U17769 ( .A(n17342), .B(n17343), .Z(n17167) );
  AND U17770 ( .A(n17344), .B(n17345), .Z(n17342) );
  AND U17771 ( .A(a[9]), .B(b[23]), .Z(n17341) );
  XOR U17772 ( .A(n17346), .B(n17172), .Z(n17174) );
  XOR U17773 ( .A(n17347), .B(n17348), .Z(n17172) );
  AND U17774 ( .A(n17349), .B(n17350), .Z(n17347) );
  AND U17775 ( .A(a[10]), .B(b[22]), .Z(n17346) );
  XOR U17776 ( .A(n17351), .B(n17177), .Z(n17179) );
  XOR U17777 ( .A(n17352), .B(n17353), .Z(n17177) );
  AND U17778 ( .A(n17354), .B(n17355), .Z(n17352) );
  AND U17779 ( .A(a[11]), .B(b[21]), .Z(n17351) );
  XOR U17780 ( .A(n17356), .B(n17182), .Z(n17184) );
  XOR U17781 ( .A(n17357), .B(n17358), .Z(n17182) );
  AND U17782 ( .A(n17359), .B(n17360), .Z(n17357) );
  AND U17783 ( .A(a[12]), .B(b[20]), .Z(n17356) );
  XOR U17784 ( .A(n17361), .B(n17187), .Z(n17189) );
  XOR U17785 ( .A(n17362), .B(n17363), .Z(n17187) );
  AND U17786 ( .A(n17364), .B(n17365), .Z(n17362) );
  AND U17787 ( .A(a[13]), .B(b[19]), .Z(n17361) );
  XOR U17788 ( .A(n17366), .B(n17192), .Z(n17194) );
  XOR U17789 ( .A(n17367), .B(n17368), .Z(n17192) );
  AND U17790 ( .A(n17369), .B(n17370), .Z(n17367) );
  AND U17791 ( .A(a[14]), .B(b[18]), .Z(n17366) );
  XOR U17792 ( .A(n17371), .B(n17197), .Z(n17199) );
  XOR U17793 ( .A(n17372), .B(n17373), .Z(n17197) );
  AND U17794 ( .A(n17374), .B(n17375), .Z(n17372) );
  AND U17795 ( .A(a[15]), .B(b[17]), .Z(n17371) );
  XOR U17796 ( .A(n17376), .B(n17202), .Z(n17204) );
  XOR U17797 ( .A(n17377), .B(n17378), .Z(n17202) );
  AND U17798 ( .A(n17379), .B(n17380), .Z(n17377) );
  AND U17799 ( .A(b[16]), .B(a[16]), .Z(n17376) );
  XOR U17800 ( .A(n17381), .B(n17207), .Z(n17209) );
  XOR U17801 ( .A(n17382), .B(n17383), .Z(n17207) );
  AND U17802 ( .A(n17384), .B(n17385), .Z(n17382) );
  AND U17803 ( .A(a[17]), .B(b[15]), .Z(n17381) );
  XOR U17804 ( .A(n17386), .B(n17212), .Z(n17214) );
  XOR U17805 ( .A(n17387), .B(n17388), .Z(n17212) );
  AND U17806 ( .A(n17389), .B(n17390), .Z(n17387) );
  AND U17807 ( .A(b[14]), .B(a[18]), .Z(n17386) );
  XOR U17808 ( .A(n17391), .B(n17217), .Z(n17219) );
  XOR U17809 ( .A(n17392), .B(n17393), .Z(n17217) );
  AND U17810 ( .A(n17394), .B(n17395), .Z(n17392) );
  AND U17811 ( .A(a[19]), .B(b[13]), .Z(n17391) );
  XOR U17812 ( .A(n17396), .B(n17222), .Z(n17224) );
  XOR U17813 ( .A(n17397), .B(n17398), .Z(n17222) );
  AND U17814 ( .A(n17399), .B(n17400), .Z(n17397) );
  AND U17815 ( .A(b[12]), .B(a[20]), .Z(n17396) );
  XOR U17816 ( .A(n17401), .B(n17227), .Z(n17229) );
  XOR U17817 ( .A(n17402), .B(n17403), .Z(n17227) );
  AND U17818 ( .A(n17404), .B(n17405), .Z(n17402) );
  AND U17819 ( .A(a[21]), .B(b[11]), .Z(n17401) );
  XOR U17820 ( .A(n17406), .B(n17232), .Z(n17234) );
  XOR U17821 ( .A(n17407), .B(n17408), .Z(n17232) );
  AND U17822 ( .A(n17409), .B(n17410), .Z(n17407) );
  AND U17823 ( .A(b[10]), .B(a[22]), .Z(n17406) );
  XOR U17824 ( .A(n17411), .B(n17237), .Z(n17239) );
  XOR U17825 ( .A(n17412), .B(n17413), .Z(n17237) );
  AND U17826 ( .A(n17414), .B(n17415), .Z(n17412) );
  AND U17827 ( .A(a[23]), .B(b[9]), .Z(n17411) );
  XOR U17828 ( .A(n17416), .B(n17242), .Z(n17244) );
  XOR U17829 ( .A(n17417), .B(n17418), .Z(n17242) );
  AND U17830 ( .A(n17419), .B(n17420), .Z(n17417) );
  AND U17831 ( .A(b[8]), .B(a[24]), .Z(n17416) );
  XOR U17832 ( .A(n17421), .B(n17247), .Z(n17249) );
  XOR U17833 ( .A(n17422), .B(n17423), .Z(n17247) );
  AND U17834 ( .A(n17424), .B(n17425), .Z(n17422) );
  AND U17835 ( .A(a[25]), .B(b[7]), .Z(n17421) );
  XOR U17836 ( .A(n17426), .B(n17252), .Z(n17254) );
  XOR U17837 ( .A(n17427), .B(n17428), .Z(n17252) );
  AND U17838 ( .A(n17429), .B(n17430), .Z(n17427) );
  AND U17839 ( .A(b[6]), .B(a[26]), .Z(n17426) );
  XOR U17840 ( .A(n17431), .B(n17257), .Z(n17259) );
  XOR U17841 ( .A(n17432), .B(n17433), .Z(n17257) );
  AND U17842 ( .A(n17434), .B(n17435), .Z(n17432) );
  AND U17843 ( .A(a[27]), .B(b[5]), .Z(n17431) );
  XOR U17844 ( .A(n17436), .B(n17262), .Z(n17264) );
  XOR U17845 ( .A(n17437), .B(n17438), .Z(n17262) );
  AND U17846 ( .A(n17439), .B(n17440), .Z(n17437) );
  AND U17847 ( .A(b[4]), .B(a[28]), .Z(n17436) );
  XOR U17848 ( .A(n17441), .B(n17267), .Z(n17269) );
  XNOR U17849 ( .A(n17442), .B(n17443), .Z(n17267) );
  AND U17850 ( .A(n17444), .B(n17445), .Z(n17442) );
  AND U17851 ( .A(a[29]), .B(b[3]), .Z(n17441) );
  AND U17852 ( .A(b[3]), .B(a[30]), .Z(n17270) );
  AND U17853 ( .A(a[31]), .B(b[3]), .Z(n17094) );
  AND U17854 ( .A(a[32]), .B(b[3]), .Z(n16918) );
  AND U17855 ( .A(a[33]), .B(b[3]), .Z(n16741) );
  AND U17856 ( .A(a[34]), .B(b[3]), .Z(n16564) );
  AND U17857 ( .A(a[34]), .B(b[4]), .Z(n16373) );
  AND U17858 ( .A(a[35]), .B(b[4]), .Z(n16198) );
  AND U17859 ( .A(a[36]), .B(b[4]), .Z(n16023) );
  AND U17860 ( .A(a[38]), .B(b[3]), .Z(n15837) );
  AND U17861 ( .A(a[39]), .B(b[3]), .Z(n15661) );
  AND U17862 ( .A(a[40]), .B(b[3]), .Z(n15485) );
  AND U17863 ( .A(a[41]), .B(b[3]), .Z(n15309) );
  AND U17864 ( .A(a[42]), .B(b[3]), .Z(n15133) );
  AND U17865 ( .A(a[43]), .B(b[3]), .Z(n14957) );
  AND U17866 ( .A(a[44]), .B(b[3]), .Z(n14781) );
  AND U17867 ( .A(a[45]), .B(b[3]), .Z(n14605) );
  AND U17868 ( .A(a[46]), .B(b[3]), .Z(n14429) );
  AND U17869 ( .A(a[47]), .B(b[3]), .Z(n14253) );
  AND U17870 ( .A(a[48]), .B(b[3]), .Z(n14077) );
  AND U17871 ( .A(a[49]), .B(b[3]), .Z(n13901) );
  AND U17872 ( .A(a[50]), .B(b[3]), .Z(n13725) );
  AND U17873 ( .A(a[51]), .B(b[3]), .Z(n13549) );
  AND U17874 ( .A(a[52]), .B(b[3]), .Z(n13373) );
  AND U17875 ( .A(a[53]), .B(b[3]), .Z(n13197) );
  AND U17876 ( .A(a[54]), .B(b[3]), .Z(n13021) );
  AND U17877 ( .A(a[55]), .B(b[3]), .Z(n12845) );
  AND U17878 ( .A(a[56]), .B(b[3]), .Z(n12669) );
  AND U17879 ( .A(a[57]), .B(b[3]), .Z(n12493) );
  AND U17880 ( .A(a[58]), .B(b[3]), .Z(n12317) );
  AND U17881 ( .A(a[59]), .B(b[3]), .Z(n12141) );
  AND U17882 ( .A(a[60]), .B(b[3]), .Z(n11965) );
  AND U17883 ( .A(a[61]), .B(b[3]), .Z(n11789) );
  AND U17884 ( .A(a[62]), .B(b[3]), .Z(n11613) );
  AND U17885 ( .A(a[63]), .B(b[3]), .Z(n11437) );
  AND U17886 ( .A(a[64]), .B(b[3]), .Z(n11260) );
  AND U17887 ( .A(a[65]), .B(b[3]), .Z(n11083) );
  AND U17888 ( .A(a[66]), .B(b[3]), .Z(n10882) );
  NAND U17889 ( .A(a[97]), .B(b[0]), .Z(n5071) );
  NAND U17890 ( .A(a[98]), .B(b[0]), .Z(n5068) );
  XOR U17891 ( .A(n17446), .B(n17447), .Z(c[99]) );
  XOR U17892 ( .A(n17448), .B(n17449), .Z(c[98]) );
  XOR U17893 ( .A(n17450), .B(n17451), .Z(c[97]) );
  XNOR U17894 ( .A(sreg[128]), .B(n17452), .Z(c[96]) );
  XOR U17895 ( .A(n5398), .B(n5397), .Z(c[127]) );
  XOR U17896 ( .A(sreg[159]), .B(n5396), .Z(n5397) );
  XOR U17897 ( .A(n17106), .B(n17453), .Z(n5398) );
  XNOR U17898 ( .A(n17107), .B(n5396), .Z(n17453) );
  XOR U17899 ( .A(n17454), .B(n17455), .Z(n5396) );
  NOR U17900 ( .A(n17456), .B(n17457), .Z(n17454) );
  NAND U17901 ( .A(a[31]), .B(b[0]), .Z(n17107) );
  XNOR U17902 ( .A(n17278), .B(n17277), .Z(n17106) );
  XOR U17903 ( .A(n17275), .B(n17458), .Z(n17277) );
  NAND U17904 ( .A(b[1]), .B(a[30]), .Z(n17458) );
  XNOR U17905 ( .A(n17445), .B(n17459), .Z(n17278) );
  XNOR U17906 ( .A(n17275), .B(n17444), .Z(n17459) );
  XNOR U17907 ( .A(n17460), .B(n17443), .Z(n17444) );
  AND U17908 ( .A(b[2]), .B(a[29]), .Z(n17460) );
  ANDN U17909 ( .B(n17461), .A(n17462), .Z(n17275) );
  XOR U17910 ( .A(n17443), .B(n17439), .Z(n17463) );
  XNOR U17911 ( .A(n17438), .B(n17434), .Z(n17464) );
  XNOR U17912 ( .A(n17433), .B(n17429), .Z(n17465) );
  XNOR U17913 ( .A(n17428), .B(n17424), .Z(n17466) );
  XNOR U17914 ( .A(n17423), .B(n17419), .Z(n17467) );
  XNOR U17915 ( .A(n17418), .B(n17414), .Z(n17468) );
  XNOR U17916 ( .A(n17413), .B(n17409), .Z(n17469) );
  XNOR U17917 ( .A(n17408), .B(n17404), .Z(n17470) );
  XNOR U17918 ( .A(n17403), .B(n17399), .Z(n17471) );
  XNOR U17919 ( .A(n17398), .B(n17394), .Z(n17472) );
  XNOR U17920 ( .A(n17393), .B(n17389), .Z(n17473) );
  XNOR U17921 ( .A(n17388), .B(n17384), .Z(n17474) );
  XNOR U17922 ( .A(n17383), .B(n17379), .Z(n17475) );
  XNOR U17923 ( .A(n17378), .B(n17374), .Z(n17476) );
  XNOR U17924 ( .A(n17373), .B(n17369), .Z(n17477) );
  XNOR U17925 ( .A(n17368), .B(n17364), .Z(n17478) );
  XNOR U17926 ( .A(n17363), .B(n17359), .Z(n17479) );
  XNOR U17927 ( .A(n17358), .B(n17354), .Z(n17480) );
  XNOR U17928 ( .A(n17353), .B(n17349), .Z(n17481) );
  XNOR U17929 ( .A(n17348), .B(n17344), .Z(n17482) );
  XNOR U17930 ( .A(n17343), .B(n17339), .Z(n17483) );
  XNOR U17931 ( .A(n17338), .B(n17334), .Z(n17484) );
  XNOR U17932 ( .A(n17333), .B(n17324), .Z(n17485) );
  XNOR U17933 ( .A(n17323), .B(n17329), .Z(n17486) );
  XNOR U17934 ( .A(n17328), .B(n17320), .Z(n17487) );
  XOR U17935 ( .A(n17319), .B(n17316), .Z(n17488) );
  XOR U17936 ( .A(n17489), .B(n17490), .Z(n17316) );
  XOR U17937 ( .A(n17314), .B(n17491), .Z(n17490) );
  XOR U17938 ( .A(n17492), .B(n17493), .Z(n17491) );
  XOR U17939 ( .A(n17494), .B(n17495), .Z(n17493) );
  NAND U17940 ( .A(a[1]), .B(b[30]), .Z(n17495) );
  AND U17941 ( .A(a[0]), .B(b[31]), .Z(n17494) );
  XOR U17942 ( .A(n17496), .B(n17492), .Z(n17489) );
  XOR U17943 ( .A(n17497), .B(n17498), .Z(n17492) );
  ANDN U17944 ( .B(n17499), .A(n17500), .Z(n17497) );
  AND U17945 ( .A(a[2]), .B(b[29]), .Z(n17496) );
  XOR U17946 ( .A(n17501), .B(n17314), .Z(n17315) );
  XOR U17947 ( .A(n17502), .B(n17503), .Z(n17314) );
  AND U17948 ( .A(n17504), .B(n17505), .Z(n17502) );
  AND U17949 ( .A(a[3]), .B(b[28]), .Z(n17501) );
  XOR U17950 ( .A(n17506), .B(n17319), .Z(n17321) );
  XOR U17951 ( .A(n17507), .B(n17508), .Z(n17319) );
  AND U17952 ( .A(n17509), .B(n17510), .Z(n17507) );
  AND U17953 ( .A(a[4]), .B(b[27]), .Z(n17506) );
  XOR U17954 ( .A(n17511), .B(n17328), .Z(n17330) );
  XOR U17955 ( .A(n17512), .B(n17513), .Z(n17328) );
  AND U17956 ( .A(n17514), .B(n17515), .Z(n17512) );
  AND U17957 ( .A(a[5]), .B(b[26]), .Z(n17511) );
  XOR U17958 ( .A(n17516), .B(n17323), .Z(n17325) );
  XOR U17959 ( .A(n17517), .B(n17518), .Z(n17323) );
  AND U17960 ( .A(n17519), .B(n17520), .Z(n17517) );
  AND U17961 ( .A(a[6]), .B(b[25]), .Z(n17516) );
  XOR U17962 ( .A(n17521), .B(n17333), .Z(n17335) );
  XOR U17963 ( .A(n17522), .B(n17523), .Z(n17333) );
  AND U17964 ( .A(n17524), .B(n17525), .Z(n17522) );
  AND U17965 ( .A(a[7]), .B(b[24]), .Z(n17521) );
  XOR U17966 ( .A(n17526), .B(n17338), .Z(n17340) );
  XOR U17967 ( .A(n17527), .B(n17528), .Z(n17338) );
  AND U17968 ( .A(n17529), .B(n17530), .Z(n17527) );
  AND U17969 ( .A(a[8]), .B(b[23]), .Z(n17526) );
  XOR U17970 ( .A(n17531), .B(n17343), .Z(n17345) );
  XOR U17971 ( .A(n17532), .B(n17533), .Z(n17343) );
  AND U17972 ( .A(n17534), .B(n17535), .Z(n17532) );
  AND U17973 ( .A(a[9]), .B(b[22]), .Z(n17531) );
  XOR U17974 ( .A(n17536), .B(n17348), .Z(n17350) );
  XOR U17975 ( .A(n17537), .B(n17538), .Z(n17348) );
  AND U17976 ( .A(n17539), .B(n17540), .Z(n17537) );
  AND U17977 ( .A(a[10]), .B(b[21]), .Z(n17536) );
  XOR U17978 ( .A(n17541), .B(n17353), .Z(n17355) );
  XOR U17979 ( .A(n17542), .B(n17543), .Z(n17353) );
  AND U17980 ( .A(n17544), .B(n17545), .Z(n17542) );
  AND U17981 ( .A(a[11]), .B(b[20]), .Z(n17541) );
  XOR U17982 ( .A(n17546), .B(n17358), .Z(n17360) );
  XOR U17983 ( .A(n17547), .B(n17548), .Z(n17358) );
  AND U17984 ( .A(n17549), .B(n17550), .Z(n17547) );
  AND U17985 ( .A(a[12]), .B(b[19]), .Z(n17546) );
  XOR U17986 ( .A(n17551), .B(n17363), .Z(n17365) );
  XOR U17987 ( .A(n17552), .B(n17553), .Z(n17363) );
  AND U17988 ( .A(n17554), .B(n17555), .Z(n17552) );
  AND U17989 ( .A(a[13]), .B(b[18]), .Z(n17551) );
  XOR U17990 ( .A(n17556), .B(n17368), .Z(n17370) );
  XOR U17991 ( .A(n17557), .B(n17558), .Z(n17368) );
  AND U17992 ( .A(n17559), .B(n17560), .Z(n17557) );
  AND U17993 ( .A(a[14]), .B(b[17]), .Z(n17556) );
  XOR U17994 ( .A(n17561), .B(n17373), .Z(n17375) );
  XOR U17995 ( .A(n17562), .B(n17563), .Z(n17373) );
  AND U17996 ( .A(n17564), .B(n17565), .Z(n17562) );
  AND U17997 ( .A(a[15]), .B(b[16]), .Z(n17561) );
  XOR U17998 ( .A(n17566), .B(n17378), .Z(n17380) );
  XOR U17999 ( .A(n17567), .B(n17568), .Z(n17378) );
  AND U18000 ( .A(n17569), .B(n17570), .Z(n17567) );
  AND U18001 ( .A(b[15]), .B(a[16]), .Z(n17566) );
  XOR U18002 ( .A(n17571), .B(n17383), .Z(n17385) );
  XOR U18003 ( .A(n17572), .B(n17573), .Z(n17383) );
  AND U18004 ( .A(n17574), .B(n17575), .Z(n17572) );
  AND U18005 ( .A(a[17]), .B(b[14]), .Z(n17571) );
  XOR U18006 ( .A(n17576), .B(n17388), .Z(n17390) );
  XOR U18007 ( .A(n17577), .B(n17578), .Z(n17388) );
  AND U18008 ( .A(n17579), .B(n17580), .Z(n17577) );
  AND U18009 ( .A(b[13]), .B(a[18]), .Z(n17576) );
  XOR U18010 ( .A(n17581), .B(n17393), .Z(n17395) );
  XOR U18011 ( .A(n17582), .B(n17583), .Z(n17393) );
  AND U18012 ( .A(n17584), .B(n17585), .Z(n17582) );
  AND U18013 ( .A(a[19]), .B(b[12]), .Z(n17581) );
  XOR U18014 ( .A(n17586), .B(n17398), .Z(n17400) );
  XOR U18015 ( .A(n17587), .B(n17588), .Z(n17398) );
  AND U18016 ( .A(n17589), .B(n17590), .Z(n17587) );
  AND U18017 ( .A(b[11]), .B(a[20]), .Z(n17586) );
  XOR U18018 ( .A(n17591), .B(n17403), .Z(n17405) );
  XOR U18019 ( .A(n17592), .B(n17593), .Z(n17403) );
  AND U18020 ( .A(n17594), .B(n17595), .Z(n17592) );
  AND U18021 ( .A(a[21]), .B(b[10]), .Z(n17591) );
  XOR U18022 ( .A(n17596), .B(n17408), .Z(n17410) );
  XOR U18023 ( .A(n17597), .B(n17598), .Z(n17408) );
  AND U18024 ( .A(n17599), .B(n17600), .Z(n17597) );
  AND U18025 ( .A(b[9]), .B(a[22]), .Z(n17596) );
  XOR U18026 ( .A(n17601), .B(n17413), .Z(n17415) );
  XOR U18027 ( .A(n17602), .B(n17603), .Z(n17413) );
  AND U18028 ( .A(n17604), .B(n17605), .Z(n17602) );
  AND U18029 ( .A(a[23]), .B(b[8]), .Z(n17601) );
  XOR U18030 ( .A(n17606), .B(n17418), .Z(n17420) );
  XOR U18031 ( .A(n17607), .B(n17608), .Z(n17418) );
  AND U18032 ( .A(n17609), .B(n17610), .Z(n17607) );
  AND U18033 ( .A(b[7]), .B(a[24]), .Z(n17606) );
  XOR U18034 ( .A(n17611), .B(n17423), .Z(n17425) );
  XOR U18035 ( .A(n17612), .B(n17613), .Z(n17423) );
  AND U18036 ( .A(n17614), .B(n17615), .Z(n17612) );
  AND U18037 ( .A(a[25]), .B(b[6]), .Z(n17611) );
  XOR U18038 ( .A(n17616), .B(n17428), .Z(n17430) );
  XOR U18039 ( .A(n17617), .B(n17618), .Z(n17428) );
  AND U18040 ( .A(n17619), .B(n17620), .Z(n17617) );
  AND U18041 ( .A(b[5]), .B(a[26]), .Z(n17616) );
  XOR U18042 ( .A(n17621), .B(n17433), .Z(n17435) );
  XOR U18043 ( .A(n17622), .B(n17623), .Z(n17433) );
  AND U18044 ( .A(n17624), .B(n17625), .Z(n17622) );
  AND U18045 ( .A(a[27]), .B(b[4]), .Z(n17621) );
  XNOR U18046 ( .A(n17626), .B(n17627), .Z(n17443) );
  NANDN U18047 ( .A(n17628), .B(n17629), .Z(n17627) );
  XOR U18048 ( .A(n17630), .B(n17438), .Z(n17440) );
  XNOR U18049 ( .A(n17631), .B(n17632), .Z(n17438) );
  AND U18050 ( .A(n17633), .B(n17634), .Z(n17631) );
  AND U18051 ( .A(b[3]), .B(a[28]), .Z(n17630) );
  XOR U18052 ( .A(n17457), .B(n17456), .Z(c[126]) );
  XOR U18053 ( .A(sreg[158]), .B(n17455), .Z(n17456) );
  XOR U18054 ( .A(n17461), .B(n17635), .Z(n17457) );
  XNOR U18055 ( .A(n17462), .B(n17455), .Z(n17635) );
  XOR U18056 ( .A(n17636), .B(n17637), .Z(n17455) );
  NOR U18057 ( .A(n17638), .B(n17639), .Z(n17636) );
  NAND U18058 ( .A(a[30]), .B(b[0]), .Z(n17462) );
  XNOR U18059 ( .A(n17628), .B(n17629), .Z(n17461) );
  XOR U18060 ( .A(n17626), .B(n17640), .Z(n17629) );
  NAND U18061 ( .A(a[29]), .B(b[1]), .Z(n17640) );
  XOR U18062 ( .A(n17634), .B(n17641), .Z(n17628) );
  XOR U18063 ( .A(n17626), .B(n17633), .Z(n17641) );
  XNOR U18064 ( .A(n17642), .B(n17632), .Z(n17633) );
  AND U18065 ( .A(b[2]), .B(a[28]), .Z(n17642) );
  NANDN U18066 ( .A(n17643), .B(n17644), .Z(n17626) );
  XOR U18067 ( .A(n17632), .B(n17624), .Z(n17645) );
  XNOR U18068 ( .A(n17623), .B(n17619), .Z(n17646) );
  XNOR U18069 ( .A(n17618), .B(n17614), .Z(n17647) );
  XNOR U18070 ( .A(n17613), .B(n17609), .Z(n17648) );
  XNOR U18071 ( .A(n17608), .B(n17604), .Z(n17649) );
  XNOR U18072 ( .A(n17603), .B(n17599), .Z(n17650) );
  XNOR U18073 ( .A(n17598), .B(n17594), .Z(n17651) );
  XNOR U18074 ( .A(n17593), .B(n17589), .Z(n17652) );
  XNOR U18075 ( .A(n17588), .B(n17584), .Z(n17653) );
  XNOR U18076 ( .A(n17583), .B(n17579), .Z(n17654) );
  XNOR U18077 ( .A(n17578), .B(n17574), .Z(n17655) );
  XNOR U18078 ( .A(n17573), .B(n17569), .Z(n17656) );
  XNOR U18079 ( .A(n17568), .B(n17564), .Z(n17657) );
  XNOR U18080 ( .A(n17563), .B(n17559), .Z(n17658) );
  XNOR U18081 ( .A(n17558), .B(n17554), .Z(n17659) );
  XNOR U18082 ( .A(n17553), .B(n17549), .Z(n17660) );
  XNOR U18083 ( .A(n17548), .B(n17544), .Z(n17661) );
  XNOR U18084 ( .A(n17543), .B(n17539), .Z(n17662) );
  XNOR U18085 ( .A(n17538), .B(n17534), .Z(n17663) );
  XNOR U18086 ( .A(n17533), .B(n17529), .Z(n17664) );
  XNOR U18087 ( .A(n17528), .B(n17524), .Z(n17665) );
  XNOR U18088 ( .A(n17523), .B(n17519), .Z(n17666) );
  XNOR U18089 ( .A(n17518), .B(n17514), .Z(n17667) );
  XNOR U18090 ( .A(n17513), .B(n17509), .Z(n17668) );
  XNOR U18091 ( .A(n17508), .B(n17504), .Z(n17669) );
  XOR U18092 ( .A(n17503), .B(n17500), .Z(n17670) );
  XOR U18093 ( .A(n17671), .B(n17672), .Z(n17500) );
  XOR U18094 ( .A(n17498), .B(n17673), .Z(n17672) );
  XOR U18095 ( .A(n17674), .B(n17675), .Z(n17673) );
  AND U18096 ( .A(a[0]), .B(b[30]), .Z(n17674) );
  XNOR U18097 ( .A(n17676), .B(n17675), .Z(n17671) );
  XNOR U18098 ( .A(n17677), .B(n17678), .Z(n17675) );
  AND U18099 ( .A(n17679), .B(n17680), .Z(n17677) );
  AND U18100 ( .A(a[1]), .B(b[29]), .Z(n17676) );
  XOR U18101 ( .A(n17681), .B(n17498), .Z(n17499) );
  XOR U18102 ( .A(n17682), .B(n17683), .Z(n17498) );
  AND U18103 ( .A(n17684), .B(n17685), .Z(n17682) );
  AND U18104 ( .A(a[2]), .B(b[28]), .Z(n17681) );
  XOR U18105 ( .A(n17686), .B(n17503), .Z(n17505) );
  XOR U18106 ( .A(n17687), .B(n17688), .Z(n17503) );
  AND U18107 ( .A(n17689), .B(n17690), .Z(n17687) );
  AND U18108 ( .A(a[3]), .B(b[27]), .Z(n17686) );
  XOR U18109 ( .A(n17691), .B(n17508), .Z(n17510) );
  XOR U18110 ( .A(n17692), .B(n17693), .Z(n17508) );
  AND U18111 ( .A(n17694), .B(n17695), .Z(n17692) );
  AND U18112 ( .A(a[4]), .B(b[26]), .Z(n17691) );
  XOR U18113 ( .A(n17696), .B(n17513), .Z(n17515) );
  XOR U18114 ( .A(n17697), .B(n17698), .Z(n17513) );
  AND U18115 ( .A(n17699), .B(n17700), .Z(n17697) );
  AND U18116 ( .A(a[5]), .B(b[25]), .Z(n17696) );
  XOR U18117 ( .A(n17701), .B(n17518), .Z(n17520) );
  XOR U18118 ( .A(n17702), .B(n17703), .Z(n17518) );
  AND U18119 ( .A(n17704), .B(n17705), .Z(n17702) );
  AND U18120 ( .A(a[6]), .B(b[24]), .Z(n17701) );
  XOR U18121 ( .A(n17706), .B(n17523), .Z(n17525) );
  XOR U18122 ( .A(n17707), .B(n17708), .Z(n17523) );
  AND U18123 ( .A(n17709), .B(n17710), .Z(n17707) );
  AND U18124 ( .A(a[7]), .B(b[23]), .Z(n17706) );
  XOR U18125 ( .A(n17711), .B(n17528), .Z(n17530) );
  XOR U18126 ( .A(n17712), .B(n17713), .Z(n17528) );
  AND U18127 ( .A(n17714), .B(n17715), .Z(n17712) );
  AND U18128 ( .A(a[8]), .B(b[22]), .Z(n17711) );
  XOR U18129 ( .A(n17716), .B(n17533), .Z(n17535) );
  XOR U18130 ( .A(n17717), .B(n17718), .Z(n17533) );
  AND U18131 ( .A(n17719), .B(n17720), .Z(n17717) );
  AND U18132 ( .A(a[9]), .B(b[21]), .Z(n17716) );
  XOR U18133 ( .A(n17721), .B(n17538), .Z(n17540) );
  XOR U18134 ( .A(n17722), .B(n17723), .Z(n17538) );
  AND U18135 ( .A(n17724), .B(n17725), .Z(n17722) );
  AND U18136 ( .A(a[10]), .B(b[20]), .Z(n17721) );
  XOR U18137 ( .A(n17726), .B(n17543), .Z(n17545) );
  XOR U18138 ( .A(n17727), .B(n17728), .Z(n17543) );
  AND U18139 ( .A(n17729), .B(n17730), .Z(n17727) );
  AND U18140 ( .A(a[11]), .B(b[19]), .Z(n17726) );
  XOR U18141 ( .A(n17731), .B(n17548), .Z(n17550) );
  XOR U18142 ( .A(n17732), .B(n17733), .Z(n17548) );
  AND U18143 ( .A(n17734), .B(n17735), .Z(n17732) );
  AND U18144 ( .A(a[12]), .B(b[18]), .Z(n17731) );
  XOR U18145 ( .A(n17736), .B(n17553), .Z(n17555) );
  XOR U18146 ( .A(n17737), .B(n17738), .Z(n17553) );
  AND U18147 ( .A(n17739), .B(n17740), .Z(n17737) );
  AND U18148 ( .A(a[13]), .B(b[17]), .Z(n17736) );
  XOR U18149 ( .A(n17741), .B(n17558), .Z(n17560) );
  XOR U18150 ( .A(n17742), .B(n17743), .Z(n17558) );
  AND U18151 ( .A(n17744), .B(n17745), .Z(n17742) );
  AND U18152 ( .A(a[14]), .B(b[16]), .Z(n17741) );
  XOR U18153 ( .A(n17746), .B(n17563), .Z(n17565) );
  XOR U18154 ( .A(n17747), .B(n17748), .Z(n17563) );
  AND U18155 ( .A(n17749), .B(n17750), .Z(n17747) );
  AND U18156 ( .A(a[15]), .B(b[15]), .Z(n17746) );
  XOR U18157 ( .A(n17751), .B(n17568), .Z(n17570) );
  XOR U18158 ( .A(n17752), .B(n17753), .Z(n17568) );
  AND U18159 ( .A(n17754), .B(n17755), .Z(n17752) );
  AND U18160 ( .A(b[14]), .B(a[16]), .Z(n17751) );
  XOR U18161 ( .A(n17756), .B(n17573), .Z(n17575) );
  XOR U18162 ( .A(n17757), .B(n17758), .Z(n17573) );
  AND U18163 ( .A(n17759), .B(n17760), .Z(n17757) );
  AND U18164 ( .A(a[17]), .B(b[13]), .Z(n17756) );
  XOR U18165 ( .A(n17761), .B(n17578), .Z(n17580) );
  XOR U18166 ( .A(n17762), .B(n17763), .Z(n17578) );
  AND U18167 ( .A(n17764), .B(n17765), .Z(n17762) );
  AND U18168 ( .A(b[12]), .B(a[18]), .Z(n17761) );
  XOR U18169 ( .A(n17766), .B(n17583), .Z(n17585) );
  XOR U18170 ( .A(n17767), .B(n17768), .Z(n17583) );
  AND U18171 ( .A(n17769), .B(n17770), .Z(n17767) );
  AND U18172 ( .A(a[19]), .B(b[11]), .Z(n17766) );
  XOR U18173 ( .A(n17771), .B(n17588), .Z(n17590) );
  XOR U18174 ( .A(n17772), .B(n17773), .Z(n17588) );
  AND U18175 ( .A(n17774), .B(n17775), .Z(n17772) );
  AND U18176 ( .A(b[10]), .B(a[20]), .Z(n17771) );
  XOR U18177 ( .A(n17776), .B(n17593), .Z(n17595) );
  XOR U18178 ( .A(n17777), .B(n17778), .Z(n17593) );
  AND U18179 ( .A(n17779), .B(n17780), .Z(n17777) );
  AND U18180 ( .A(a[21]), .B(b[9]), .Z(n17776) );
  XOR U18181 ( .A(n17781), .B(n17598), .Z(n17600) );
  XOR U18182 ( .A(n17782), .B(n17783), .Z(n17598) );
  AND U18183 ( .A(n17784), .B(n17785), .Z(n17782) );
  AND U18184 ( .A(b[8]), .B(a[22]), .Z(n17781) );
  XOR U18185 ( .A(n17786), .B(n17603), .Z(n17605) );
  XOR U18186 ( .A(n17787), .B(n17788), .Z(n17603) );
  AND U18187 ( .A(n17789), .B(n17790), .Z(n17787) );
  AND U18188 ( .A(a[23]), .B(b[7]), .Z(n17786) );
  XOR U18189 ( .A(n17791), .B(n17608), .Z(n17610) );
  XOR U18190 ( .A(n17792), .B(n17793), .Z(n17608) );
  AND U18191 ( .A(n17794), .B(n17795), .Z(n17792) );
  AND U18192 ( .A(b[6]), .B(a[24]), .Z(n17791) );
  XOR U18193 ( .A(n17796), .B(n17613), .Z(n17615) );
  XOR U18194 ( .A(n17797), .B(n17798), .Z(n17613) );
  AND U18195 ( .A(n17799), .B(n17800), .Z(n17797) );
  AND U18196 ( .A(a[25]), .B(b[5]), .Z(n17796) );
  XOR U18197 ( .A(n17801), .B(n17618), .Z(n17620) );
  XOR U18198 ( .A(n17802), .B(n17803), .Z(n17618) );
  AND U18199 ( .A(n17804), .B(n17805), .Z(n17802) );
  AND U18200 ( .A(b[4]), .B(a[26]), .Z(n17801) );
  XNOR U18201 ( .A(n17806), .B(n17807), .Z(n17632) );
  NANDN U18202 ( .A(n17808), .B(n17809), .Z(n17807) );
  XOR U18203 ( .A(n17810), .B(n17623), .Z(n17625) );
  XNOR U18204 ( .A(n17811), .B(n17812), .Z(n17623) );
  AND U18205 ( .A(n17813), .B(n17814), .Z(n17811) );
  AND U18206 ( .A(a[27]), .B(b[3]), .Z(n17810) );
  XOR U18207 ( .A(n17639), .B(n17638), .Z(c[125]) );
  XOR U18208 ( .A(sreg[157]), .B(n17637), .Z(n17638) );
  XOR U18209 ( .A(n17644), .B(n17815), .Z(n17639) );
  XNOR U18210 ( .A(n17643), .B(n17637), .Z(n17815) );
  XOR U18211 ( .A(n17816), .B(n17817), .Z(n17637) );
  NOR U18212 ( .A(n17818), .B(n17819), .Z(n17816) );
  NAND U18213 ( .A(a[29]), .B(b[0]), .Z(n17643) );
  XNOR U18214 ( .A(n17808), .B(n17809), .Z(n17644) );
  XOR U18215 ( .A(n17806), .B(n17820), .Z(n17809) );
  NAND U18216 ( .A(b[1]), .B(a[28]), .Z(n17820) );
  XOR U18217 ( .A(n17814), .B(n17821), .Z(n17808) );
  XOR U18218 ( .A(n17806), .B(n17813), .Z(n17821) );
  XNOR U18219 ( .A(n17822), .B(n17812), .Z(n17813) );
  AND U18220 ( .A(b[2]), .B(a[27]), .Z(n17822) );
  NANDN U18221 ( .A(n17823), .B(n17824), .Z(n17806) );
  XOR U18222 ( .A(n17812), .B(n17804), .Z(n17825) );
  XNOR U18223 ( .A(n17803), .B(n17799), .Z(n17826) );
  XNOR U18224 ( .A(n17798), .B(n17794), .Z(n17827) );
  XNOR U18225 ( .A(n17793), .B(n17789), .Z(n17828) );
  XNOR U18226 ( .A(n17788), .B(n17784), .Z(n17829) );
  XNOR U18227 ( .A(n17783), .B(n17779), .Z(n17830) );
  XNOR U18228 ( .A(n17778), .B(n17774), .Z(n17831) );
  XNOR U18229 ( .A(n17773), .B(n17769), .Z(n17832) );
  XNOR U18230 ( .A(n17768), .B(n17764), .Z(n17833) );
  XNOR U18231 ( .A(n17763), .B(n17759), .Z(n17834) );
  XNOR U18232 ( .A(n17758), .B(n17754), .Z(n17835) );
  XNOR U18233 ( .A(n17753), .B(n17749), .Z(n17836) );
  XNOR U18234 ( .A(n17748), .B(n17744), .Z(n17837) );
  XNOR U18235 ( .A(n17743), .B(n17739), .Z(n17838) );
  XNOR U18236 ( .A(n17738), .B(n17734), .Z(n17839) );
  XNOR U18237 ( .A(n17733), .B(n17729), .Z(n17840) );
  XNOR U18238 ( .A(n17728), .B(n17724), .Z(n17841) );
  XNOR U18239 ( .A(n17723), .B(n17719), .Z(n17842) );
  XNOR U18240 ( .A(n17718), .B(n17714), .Z(n17843) );
  XNOR U18241 ( .A(n17713), .B(n17709), .Z(n17844) );
  XNOR U18242 ( .A(n17708), .B(n17704), .Z(n17845) );
  XNOR U18243 ( .A(n17703), .B(n17699), .Z(n17846) );
  XNOR U18244 ( .A(n17698), .B(n17694), .Z(n17847) );
  XNOR U18245 ( .A(n17693), .B(n17689), .Z(n17848) );
  XNOR U18246 ( .A(n17688), .B(n17684), .Z(n17849) );
  XNOR U18247 ( .A(n17683), .B(n17679), .Z(n17850) );
  XOR U18248 ( .A(n17851), .B(n17678), .Z(n17679) );
  AND U18249 ( .A(a[0]), .B(b[29]), .Z(n17851) );
  XOR U18250 ( .A(n17852), .B(n17678), .Z(n17680) );
  XNOR U18251 ( .A(n17853), .B(n17854), .Z(n17678) );
  AND U18252 ( .A(n17855), .B(n17856), .Z(n17853) );
  AND U18253 ( .A(a[1]), .B(b[28]), .Z(n17852) );
  XOR U18254 ( .A(n17857), .B(n17683), .Z(n17685) );
  XOR U18255 ( .A(n17858), .B(n17859), .Z(n17683) );
  AND U18256 ( .A(n17860), .B(n17861), .Z(n17858) );
  AND U18257 ( .A(a[2]), .B(b[27]), .Z(n17857) );
  XOR U18258 ( .A(n17862), .B(n17688), .Z(n17690) );
  XOR U18259 ( .A(n17863), .B(n17864), .Z(n17688) );
  AND U18260 ( .A(n17865), .B(n17866), .Z(n17863) );
  AND U18261 ( .A(a[3]), .B(b[26]), .Z(n17862) );
  XOR U18262 ( .A(n17867), .B(n17693), .Z(n17695) );
  XOR U18263 ( .A(n17868), .B(n17869), .Z(n17693) );
  AND U18264 ( .A(n17870), .B(n17871), .Z(n17868) );
  AND U18265 ( .A(a[4]), .B(b[25]), .Z(n17867) );
  XOR U18266 ( .A(n17872), .B(n17698), .Z(n17700) );
  XOR U18267 ( .A(n17873), .B(n17874), .Z(n17698) );
  AND U18268 ( .A(n17875), .B(n17876), .Z(n17873) );
  AND U18269 ( .A(a[5]), .B(b[24]), .Z(n17872) );
  XOR U18270 ( .A(n17877), .B(n17703), .Z(n17705) );
  XOR U18271 ( .A(n17878), .B(n17879), .Z(n17703) );
  AND U18272 ( .A(n17880), .B(n17881), .Z(n17878) );
  AND U18273 ( .A(a[6]), .B(b[23]), .Z(n17877) );
  XOR U18274 ( .A(n17882), .B(n17708), .Z(n17710) );
  XOR U18275 ( .A(n17883), .B(n17884), .Z(n17708) );
  AND U18276 ( .A(n17885), .B(n17886), .Z(n17883) );
  AND U18277 ( .A(a[7]), .B(b[22]), .Z(n17882) );
  XOR U18278 ( .A(n17887), .B(n17713), .Z(n17715) );
  XOR U18279 ( .A(n17888), .B(n17889), .Z(n17713) );
  AND U18280 ( .A(n17890), .B(n17891), .Z(n17888) );
  AND U18281 ( .A(a[8]), .B(b[21]), .Z(n17887) );
  XOR U18282 ( .A(n17892), .B(n17718), .Z(n17720) );
  XOR U18283 ( .A(n17893), .B(n17894), .Z(n17718) );
  AND U18284 ( .A(n17895), .B(n17896), .Z(n17893) );
  AND U18285 ( .A(a[9]), .B(b[20]), .Z(n17892) );
  XOR U18286 ( .A(n17897), .B(n17723), .Z(n17725) );
  XOR U18287 ( .A(n17898), .B(n17899), .Z(n17723) );
  AND U18288 ( .A(n17900), .B(n17901), .Z(n17898) );
  AND U18289 ( .A(a[10]), .B(b[19]), .Z(n17897) );
  XOR U18290 ( .A(n17902), .B(n17728), .Z(n17730) );
  XOR U18291 ( .A(n17903), .B(n17904), .Z(n17728) );
  AND U18292 ( .A(n17905), .B(n17906), .Z(n17903) );
  AND U18293 ( .A(a[11]), .B(b[18]), .Z(n17902) );
  XOR U18294 ( .A(n17907), .B(n17733), .Z(n17735) );
  XOR U18295 ( .A(n17908), .B(n17909), .Z(n17733) );
  AND U18296 ( .A(n17910), .B(n17911), .Z(n17908) );
  AND U18297 ( .A(a[12]), .B(b[17]), .Z(n17907) );
  XOR U18298 ( .A(n17912), .B(n17738), .Z(n17740) );
  XOR U18299 ( .A(n17913), .B(n17914), .Z(n17738) );
  AND U18300 ( .A(n17915), .B(n17916), .Z(n17913) );
  AND U18301 ( .A(a[13]), .B(b[16]), .Z(n17912) );
  XOR U18302 ( .A(n17917), .B(n17743), .Z(n17745) );
  XOR U18303 ( .A(n17918), .B(n17919), .Z(n17743) );
  AND U18304 ( .A(n17920), .B(n17921), .Z(n17918) );
  AND U18305 ( .A(a[14]), .B(b[15]), .Z(n17917) );
  XOR U18306 ( .A(n17922), .B(n17748), .Z(n17750) );
  XOR U18307 ( .A(n17923), .B(n17924), .Z(n17748) );
  AND U18308 ( .A(n17925), .B(n17926), .Z(n17923) );
  AND U18309 ( .A(a[15]), .B(b[14]), .Z(n17922) );
  XOR U18310 ( .A(n17927), .B(n17753), .Z(n17755) );
  XOR U18311 ( .A(n17928), .B(n17929), .Z(n17753) );
  AND U18312 ( .A(n17930), .B(n17931), .Z(n17928) );
  AND U18313 ( .A(b[13]), .B(a[16]), .Z(n17927) );
  XOR U18314 ( .A(n17932), .B(n17758), .Z(n17760) );
  XOR U18315 ( .A(n17933), .B(n17934), .Z(n17758) );
  AND U18316 ( .A(n17935), .B(n17936), .Z(n17933) );
  AND U18317 ( .A(a[17]), .B(b[12]), .Z(n17932) );
  XOR U18318 ( .A(n17937), .B(n17763), .Z(n17765) );
  XOR U18319 ( .A(n17938), .B(n17939), .Z(n17763) );
  AND U18320 ( .A(n17940), .B(n17941), .Z(n17938) );
  AND U18321 ( .A(b[11]), .B(a[18]), .Z(n17937) );
  XOR U18322 ( .A(n17942), .B(n17768), .Z(n17770) );
  XOR U18323 ( .A(n17943), .B(n17944), .Z(n17768) );
  AND U18324 ( .A(n17945), .B(n17946), .Z(n17943) );
  AND U18325 ( .A(a[19]), .B(b[10]), .Z(n17942) );
  XOR U18326 ( .A(n17947), .B(n17773), .Z(n17775) );
  XOR U18327 ( .A(n17948), .B(n17949), .Z(n17773) );
  AND U18328 ( .A(n17950), .B(n17951), .Z(n17948) );
  AND U18329 ( .A(b[9]), .B(a[20]), .Z(n17947) );
  XOR U18330 ( .A(n17952), .B(n17778), .Z(n17780) );
  XOR U18331 ( .A(n17953), .B(n17954), .Z(n17778) );
  AND U18332 ( .A(n17955), .B(n17956), .Z(n17953) );
  AND U18333 ( .A(a[21]), .B(b[8]), .Z(n17952) );
  XOR U18334 ( .A(n17957), .B(n17783), .Z(n17785) );
  XOR U18335 ( .A(n17958), .B(n17959), .Z(n17783) );
  AND U18336 ( .A(n17960), .B(n17961), .Z(n17958) );
  AND U18337 ( .A(b[7]), .B(a[22]), .Z(n17957) );
  XOR U18338 ( .A(n17962), .B(n17788), .Z(n17790) );
  XOR U18339 ( .A(n17963), .B(n17964), .Z(n17788) );
  AND U18340 ( .A(n17965), .B(n17966), .Z(n17963) );
  AND U18341 ( .A(a[23]), .B(b[6]), .Z(n17962) );
  XOR U18342 ( .A(n17967), .B(n17793), .Z(n17795) );
  XOR U18343 ( .A(n17968), .B(n17969), .Z(n17793) );
  AND U18344 ( .A(n17970), .B(n17971), .Z(n17968) );
  AND U18345 ( .A(b[5]), .B(a[24]), .Z(n17967) );
  XOR U18346 ( .A(n17972), .B(n17798), .Z(n17800) );
  XOR U18347 ( .A(n17973), .B(n17974), .Z(n17798) );
  AND U18348 ( .A(n17975), .B(n17976), .Z(n17973) );
  AND U18349 ( .A(a[25]), .B(b[4]), .Z(n17972) );
  XNOR U18350 ( .A(n17977), .B(n17978), .Z(n17812) );
  NANDN U18351 ( .A(n17979), .B(n17980), .Z(n17978) );
  XOR U18352 ( .A(n17981), .B(n17803), .Z(n17805) );
  XNOR U18353 ( .A(n17982), .B(n17983), .Z(n17803) );
  AND U18354 ( .A(n17984), .B(n17985), .Z(n17982) );
  AND U18355 ( .A(b[3]), .B(a[26]), .Z(n17981) );
  XOR U18356 ( .A(n17819), .B(n17818), .Z(c[124]) );
  XOR U18357 ( .A(sreg[156]), .B(n17817), .Z(n17818) );
  XOR U18358 ( .A(n17824), .B(n17986), .Z(n17819) );
  XNOR U18359 ( .A(n17823), .B(n17817), .Z(n17986) );
  XOR U18360 ( .A(n17987), .B(n17988), .Z(n17817) );
  NOR U18361 ( .A(n17989), .B(n17990), .Z(n17987) );
  NAND U18362 ( .A(a[28]), .B(b[0]), .Z(n17823) );
  XNOR U18363 ( .A(n17979), .B(n17980), .Z(n17824) );
  XOR U18364 ( .A(n17977), .B(n17991), .Z(n17980) );
  NAND U18365 ( .A(a[27]), .B(b[1]), .Z(n17991) );
  XOR U18366 ( .A(n17985), .B(n17992), .Z(n17979) );
  XOR U18367 ( .A(n17977), .B(n17984), .Z(n17992) );
  XNOR U18368 ( .A(n17993), .B(n17983), .Z(n17984) );
  AND U18369 ( .A(b[2]), .B(a[26]), .Z(n17993) );
  NANDN U18370 ( .A(n17994), .B(n17995), .Z(n17977) );
  XOR U18371 ( .A(n17983), .B(n17975), .Z(n17996) );
  XNOR U18372 ( .A(n17974), .B(n17970), .Z(n17997) );
  XNOR U18373 ( .A(n17969), .B(n17965), .Z(n17998) );
  XNOR U18374 ( .A(n17964), .B(n17960), .Z(n17999) );
  XNOR U18375 ( .A(n17959), .B(n17955), .Z(n18000) );
  XNOR U18376 ( .A(n17954), .B(n17950), .Z(n18001) );
  XNOR U18377 ( .A(n17949), .B(n17945), .Z(n18002) );
  XNOR U18378 ( .A(n17944), .B(n17940), .Z(n18003) );
  XNOR U18379 ( .A(n17939), .B(n17935), .Z(n18004) );
  XNOR U18380 ( .A(n17934), .B(n17930), .Z(n18005) );
  XNOR U18381 ( .A(n17929), .B(n17925), .Z(n18006) );
  XNOR U18382 ( .A(n17924), .B(n17920), .Z(n18007) );
  XNOR U18383 ( .A(n17919), .B(n17915), .Z(n18008) );
  XNOR U18384 ( .A(n17914), .B(n17910), .Z(n18009) );
  XNOR U18385 ( .A(n17909), .B(n17905), .Z(n18010) );
  XNOR U18386 ( .A(n17904), .B(n17900), .Z(n18011) );
  XNOR U18387 ( .A(n17899), .B(n17895), .Z(n18012) );
  XNOR U18388 ( .A(n17894), .B(n17890), .Z(n18013) );
  XNOR U18389 ( .A(n17889), .B(n17885), .Z(n18014) );
  XNOR U18390 ( .A(n17884), .B(n17880), .Z(n18015) );
  XNOR U18391 ( .A(n17879), .B(n17875), .Z(n18016) );
  XNOR U18392 ( .A(n17874), .B(n17870), .Z(n18017) );
  XNOR U18393 ( .A(n17869), .B(n17865), .Z(n18018) );
  XNOR U18394 ( .A(n17864), .B(n17860), .Z(n18019) );
  XNOR U18395 ( .A(n17859), .B(n17855), .Z(n18020) );
  XNOR U18396 ( .A(n18021), .B(n17854), .Z(n17855) );
  AND U18397 ( .A(a[0]), .B(b[28]), .Z(n18021) );
  XNOR U18398 ( .A(n18022), .B(n17854), .Z(n17856) );
  XNOR U18399 ( .A(n18023), .B(n18024), .Z(n17854) );
  AND U18400 ( .A(n18025), .B(n18026), .Z(n18023) );
  AND U18401 ( .A(a[1]), .B(b[27]), .Z(n18022) );
  XOR U18402 ( .A(n18027), .B(n17859), .Z(n17861) );
  XOR U18403 ( .A(n18028), .B(n18029), .Z(n17859) );
  AND U18404 ( .A(n18030), .B(n18031), .Z(n18028) );
  AND U18405 ( .A(a[2]), .B(b[26]), .Z(n18027) );
  XOR U18406 ( .A(n18032), .B(n17864), .Z(n17866) );
  XOR U18407 ( .A(n18033), .B(n18034), .Z(n17864) );
  AND U18408 ( .A(n18035), .B(n18036), .Z(n18033) );
  AND U18409 ( .A(a[3]), .B(b[25]), .Z(n18032) );
  XOR U18410 ( .A(n18037), .B(n17869), .Z(n17871) );
  XOR U18411 ( .A(n18038), .B(n18039), .Z(n17869) );
  AND U18412 ( .A(n18040), .B(n18041), .Z(n18038) );
  AND U18413 ( .A(a[4]), .B(b[24]), .Z(n18037) );
  XOR U18414 ( .A(n18042), .B(n17874), .Z(n17876) );
  XOR U18415 ( .A(n18043), .B(n18044), .Z(n17874) );
  AND U18416 ( .A(n18045), .B(n18046), .Z(n18043) );
  AND U18417 ( .A(a[5]), .B(b[23]), .Z(n18042) );
  XOR U18418 ( .A(n18047), .B(n17879), .Z(n17881) );
  XOR U18419 ( .A(n18048), .B(n18049), .Z(n17879) );
  AND U18420 ( .A(n18050), .B(n18051), .Z(n18048) );
  AND U18421 ( .A(a[6]), .B(b[22]), .Z(n18047) );
  XOR U18422 ( .A(n18052), .B(n17884), .Z(n17886) );
  XOR U18423 ( .A(n18053), .B(n18054), .Z(n17884) );
  AND U18424 ( .A(n18055), .B(n18056), .Z(n18053) );
  AND U18425 ( .A(a[7]), .B(b[21]), .Z(n18052) );
  XOR U18426 ( .A(n18057), .B(n17889), .Z(n17891) );
  XOR U18427 ( .A(n18058), .B(n18059), .Z(n17889) );
  AND U18428 ( .A(n18060), .B(n18061), .Z(n18058) );
  AND U18429 ( .A(a[8]), .B(b[20]), .Z(n18057) );
  XOR U18430 ( .A(n18062), .B(n17894), .Z(n17896) );
  XOR U18431 ( .A(n18063), .B(n18064), .Z(n17894) );
  AND U18432 ( .A(n18065), .B(n18066), .Z(n18063) );
  AND U18433 ( .A(a[9]), .B(b[19]), .Z(n18062) );
  XOR U18434 ( .A(n18067), .B(n17899), .Z(n17901) );
  XOR U18435 ( .A(n18068), .B(n18069), .Z(n17899) );
  AND U18436 ( .A(n18070), .B(n18071), .Z(n18068) );
  AND U18437 ( .A(a[10]), .B(b[18]), .Z(n18067) );
  XOR U18438 ( .A(n18072), .B(n17904), .Z(n17906) );
  XOR U18439 ( .A(n18073), .B(n18074), .Z(n17904) );
  AND U18440 ( .A(n18075), .B(n18076), .Z(n18073) );
  AND U18441 ( .A(a[11]), .B(b[17]), .Z(n18072) );
  XOR U18442 ( .A(n18077), .B(n17909), .Z(n17911) );
  XOR U18443 ( .A(n18078), .B(n18079), .Z(n17909) );
  AND U18444 ( .A(n18080), .B(n18081), .Z(n18078) );
  AND U18445 ( .A(a[12]), .B(b[16]), .Z(n18077) );
  XOR U18446 ( .A(n18082), .B(n17914), .Z(n17916) );
  XOR U18447 ( .A(n18083), .B(n18084), .Z(n17914) );
  AND U18448 ( .A(n18085), .B(n18086), .Z(n18083) );
  AND U18449 ( .A(a[13]), .B(b[15]), .Z(n18082) );
  XOR U18450 ( .A(n18087), .B(n17919), .Z(n17921) );
  XOR U18451 ( .A(n18088), .B(n18089), .Z(n17919) );
  AND U18452 ( .A(n18090), .B(n18091), .Z(n18088) );
  AND U18453 ( .A(b[14]), .B(a[14]), .Z(n18087) );
  XOR U18454 ( .A(n18092), .B(n17924), .Z(n17926) );
  XOR U18455 ( .A(n18093), .B(n18094), .Z(n17924) );
  AND U18456 ( .A(n18095), .B(n18096), .Z(n18093) );
  AND U18457 ( .A(a[15]), .B(b[13]), .Z(n18092) );
  XOR U18458 ( .A(n18097), .B(n17929), .Z(n17931) );
  XOR U18459 ( .A(n18098), .B(n18099), .Z(n17929) );
  AND U18460 ( .A(n18100), .B(n18101), .Z(n18098) );
  AND U18461 ( .A(b[12]), .B(a[16]), .Z(n18097) );
  XOR U18462 ( .A(n18102), .B(n17934), .Z(n17936) );
  XOR U18463 ( .A(n18103), .B(n18104), .Z(n17934) );
  AND U18464 ( .A(n18105), .B(n18106), .Z(n18103) );
  AND U18465 ( .A(a[17]), .B(b[11]), .Z(n18102) );
  XOR U18466 ( .A(n18107), .B(n17939), .Z(n17941) );
  XOR U18467 ( .A(n18108), .B(n18109), .Z(n17939) );
  AND U18468 ( .A(n18110), .B(n18111), .Z(n18108) );
  AND U18469 ( .A(b[10]), .B(a[18]), .Z(n18107) );
  XOR U18470 ( .A(n18112), .B(n17944), .Z(n17946) );
  XOR U18471 ( .A(n18113), .B(n18114), .Z(n17944) );
  AND U18472 ( .A(n18115), .B(n18116), .Z(n18113) );
  AND U18473 ( .A(a[19]), .B(b[9]), .Z(n18112) );
  XOR U18474 ( .A(n18117), .B(n17949), .Z(n17951) );
  XOR U18475 ( .A(n18118), .B(n18119), .Z(n17949) );
  AND U18476 ( .A(n18120), .B(n18121), .Z(n18118) );
  AND U18477 ( .A(b[8]), .B(a[20]), .Z(n18117) );
  XOR U18478 ( .A(n18122), .B(n17954), .Z(n17956) );
  XOR U18479 ( .A(n18123), .B(n18124), .Z(n17954) );
  AND U18480 ( .A(n18125), .B(n18126), .Z(n18123) );
  AND U18481 ( .A(a[21]), .B(b[7]), .Z(n18122) );
  XOR U18482 ( .A(n18127), .B(n17959), .Z(n17961) );
  XOR U18483 ( .A(n18128), .B(n18129), .Z(n17959) );
  AND U18484 ( .A(n18130), .B(n18131), .Z(n18128) );
  AND U18485 ( .A(b[6]), .B(a[22]), .Z(n18127) );
  XOR U18486 ( .A(n18132), .B(n17964), .Z(n17966) );
  XOR U18487 ( .A(n18133), .B(n18134), .Z(n17964) );
  AND U18488 ( .A(n18135), .B(n18136), .Z(n18133) );
  AND U18489 ( .A(a[23]), .B(b[5]), .Z(n18132) );
  XOR U18490 ( .A(n18137), .B(n17969), .Z(n17971) );
  XOR U18491 ( .A(n18138), .B(n18139), .Z(n17969) );
  AND U18492 ( .A(n18140), .B(n18141), .Z(n18138) );
  AND U18493 ( .A(b[4]), .B(a[24]), .Z(n18137) );
  XNOR U18494 ( .A(n18142), .B(n18143), .Z(n17983) );
  NANDN U18495 ( .A(n18144), .B(n18145), .Z(n18143) );
  XOR U18496 ( .A(n18146), .B(n17974), .Z(n17976) );
  XNOR U18497 ( .A(n18147), .B(n18148), .Z(n17974) );
  AND U18498 ( .A(n18149), .B(n18150), .Z(n18147) );
  AND U18499 ( .A(a[25]), .B(b[3]), .Z(n18146) );
  XOR U18500 ( .A(n17990), .B(n17989), .Z(c[123]) );
  XOR U18501 ( .A(sreg[155]), .B(n17988), .Z(n17989) );
  XOR U18502 ( .A(n17995), .B(n18151), .Z(n17990) );
  XNOR U18503 ( .A(n17994), .B(n17988), .Z(n18151) );
  XOR U18504 ( .A(n18152), .B(n18153), .Z(n17988) );
  NOR U18505 ( .A(n18154), .B(n18155), .Z(n18152) );
  NAND U18506 ( .A(a[27]), .B(b[0]), .Z(n17994) );
  XNOR U18507 ( .A(n18144), .B(n18145), .Z(n17995) );
  XOR U18508 ( .A(n18142), .B(n18156), .Z(n18145) );
  NAND U18509 ( .A(b[1]), .B(a[26]), .Z(n18156) );
  XOR U18510 ( .A(n18150), .B(n18157), .Z(n18144) );
  XOR U18511 ( .A(n18142), .B(n18149), .Z(n18157) );
  XNOR U18512 ( .A(n18158), .B(n18148), .Z(n18149) );
  AND U18513 ( .A(b[2]), .B(a[25]), .Z(n18158) );
  NANDN U18514 ( .A(n18159), .B(n18160), .Z(n18142) );
  XOR U18515 ( .A(n18148), .B(n18140), .Z(n18161) );
  XNOR U18516 ( .A(n18139), .B(n18135), .Z(n18162) );
  XNOR U18517 ( .A(n18134), .B(n18130), .Z(n18163) );
  XNOR U18518 ( .A(n18129), .B(n18125), .Z(n18164) );
  XNOR U18519 ( .A(n18124), .B(n18120), .Z(n18165) );
  XNOR U18520 ( .A(n18119), .B(n18115), .Z(n18166) );
  XNOR U18521 ( .A(n18114), .B(n18110), .Z(n18167) );
  XNOR U18522 ( .A(n18109), .B(n18105), .Z(n18168) );
  XNOR U18523 ( .A(n18104), .B(n18100), .Z(n18169) );
  XNOR U18524 ( .A(n18099), .B(n18095), .Z(n18170) );
  XNOR U18525 ( .A(n18094), .B(n18090), .Z(n18171) );
  XNOR U18526 ( .A(n18089), .B(n18085), .Z(n18172) );
  XNOR U18527 ( .A(n18084), .B(n18080), .Z(n18173) );
  XNOR U18528 ( .A(n18079), .B(n18075), .Z(n18174) );
  XNOR U18529 ( .A(n18074), .B(n18070), .Z(n18175) );
  XNOR U18530 ( .A(n18069), .B(n18065), .Z(n18176) );
  XNOR U18531 ( .A(n18064), .B(n18060), .Z(n18177) );
  XNOR U18532 ( .A(n18059), .B(n18055), .Z(n18178) );
  XNOR U18533 ( .A(n18054), .B(n18050), .Z(n18179) );
  XNOR U18534 ( .A(n18049), .B(n18045), .Z(n18180) );
  XNOR U18535 ( .A(n18044), .B(n18040), .Z(n18181) );
  XNOR U18536 ( .A(n18039), .B(n18035), .Z(n18182) );
  XNOR U18537 ( .A(n18034), .B(n18030), .Z(n18183) );
  XNOR U18538 ( .A(n18029), .B(n18025), .Z(n18184) );
  XOR U18539 ( .A(n18185), .B(n18024), .Z(n18025) );
  AND U18540 ( .A(a[0]), .B(b[27]), .Z(n18185) );
  XOR U18541 ( .A(n18186), .B(n18024), .Z(n18026) );
  XNOR U18542 ( .A(n18187), .B(n18188), .Z(n18024) );
  AND U18543 ( .A(n18189), .B(n18190), .Z(n18187) );
  AND U18544 ( .A(a[1]), .B(b[26]), .Z(n18186) );
  XOR U18545 ( .A(n18191), .B(n18029), .Z(n18031) );
  XOR U18546 ( .A(n18192), .B(n18193), .Z(n18029) );
  AND U18547 ( .A(n18194), .B(n18195), .Z(n18192) );
  AND U18548 ( .A(a[2]), .B(b[25]), .Z(n18191) );
  XOR U18549 ( .A(n18196), .B(n18034), .Z(n18036) );
  XOR U18550 ( .A(n18197), .B(n18198), .Z(n18034) );
  AND U18551 ( .A(n18199), .B(n18200), .Z(n18197) );
  AND U18552 ( .A(a[3]), .B(b[24]), .Z(n18196) );
  XOR U18553 ( .A(n18201), .B(n18039), .Z(n18041) );
  XOR U18554 ( .A(n18202), .B(n18203), .Z(n18039) );
  AND U18555 ( .A(n18204), .B(n18205), .Z(n18202) );
  AND U18556 ( .A(a[4]), .B(b[23]), .Z(n18201) );
  XOR U18557 ( .A(n18206), .B(n18044), .Z(n18046) );
  XOR U18558 ( .A(n18207), .B(n18208), .Z(n18044) );
  AND U18559 ( .A(n18209), .B(n18210), .Z(n18207) );
  AND U18560 ( .A(a[5]), .B(b[22]), .Z(n18206) );
  XOR U18561 ( .A(n18211), .B(n18049), .Z(n18051) );
  XOR U18562 ( .A(n18212), .B(n18213), .Z(n18049) );
  AND U18563 ( .A(n18214), .B(n18215), .Z(n18212) );
  AND U18564 ( .A(a[6]), .B(b[21]), .Z(n18211) );
  XOR U18565 ( .A(n18216), .B(n18054), .Z(n18056) );
  XOR U18566 ( .A(n18217), .B(n18218), .Z(n18054) );
  AND U18567 ( .A(n18219), .B(n18220), .Z(n18217) );
  AND U18568 ( .A(a[7]), .B(b[20]), .Z(n18216) );
  XOR U18569 ( .A(n18221), .B(n18059), .Z(n18061) );
  XOR U18570 ( .A(n18222), .B(n18223), .Z(n18059) );
  AND U18571 ( .A(n18224), .B(n18225), .Z(n18222) );
  AND U18572 ( .A(a[8]), .B(b[19]), .Z(n18221) );
  XOR U18573 ( .A(n18226), .B(n18064), .Z(n18066) );
  XOR U18574 ( .A(n18227), .B(n18228), .Z(n18064) );
  AND U18575 ( .A(n18229), .B(n18230), .Z(n18227) );
  AND U18576 ( .A(a[9]), .B(b[18]), .Z(n18226) );
  XOR U18577 ( .A(n18231), .B(n18069), .Z(n18071) );
  XOR U18578 ( .A(n18232), .B(n18233), .Z(n18069) );
  AND U18579 ( .A(n18234), .B(n18235), .Z(n18232) );
  AND U18580 ( .A(a[10]), .B(b[17]), .Z(n18231) );
  XOR U18581 ( .A(n18236), .B(n18074), .Z(n18076) );
  XOR U18582 ( .A(n18237), .B(n18238), .Z(n18074) );
  AND U18583 ( .A(n18239), .B(n18240), .Z(n18237) );
  AND U18584 ( .A(a[11]), .B(b[16]), .Z(n18236) );
  XOR U18585 ( .A(n18241), .B(n18079), .Z(n18081) );
  XOR U18586 ( .A(n18242), .B(n18243), .Z(n18079) );
  AND U18587 ( .A(n18244), .B(n18245), .Z(n18242) );
  AND U18588 ( .A(a[12]), .B(b[15]), .Z(n18241) );
  XOR U18589 ( .A(n18246), .B(n18084), .Z(n18086) );
  XOR U18590 ( .A(n18247), .B(n18248), .Z(n18084) );
  AND U18591 ( .A(n18249), .B(n18250), .Z(n18247) );
  AND U18592 ( .A(a[13]), .B(b[14]), .Z(n18246) );
  XOR U18593 ( .A(n18251), .B(n18089), .Z(n18091) );
  XOR U18594 ( .A(n18252), .B(n18253), .Z(n18089) );
  AND U18595 ( .A(n18254), .B(n18255), .Z(n18252) );
  AND U18596 ( .A(b[13]), .B(a[14]), .Z(n18251) );
  XOR U18597 ( .A(n18256), .B(n18094), .Z(n18096) );
  XOR U18598 ( .A(n18257), .B(n18258), .Z(n18094) );
  AND U18599 ( .A(n18259), .B(n18260), .Z(n18257) );
  AND U18600 ( .A(a[15]), .B(b[12]), .Z(n18256) );
  XOR U18601 ( .A(n18261), .B(n18099), .Z(n18101) );
  XOR U18602 ( .A(n18262), .B(n18263), .Z(n18099) );
  AND U18603 ( .A(n18264), .B(n18265), .Z(n18262) );
  AND U18604 ( .A(b[11]), .B(a[16]), .Z(n18261) );
  XOR U18605 ( .A(n18266), .B(n18104), .Z(n18106) );
  XOR U18606 ( .A(n18267), .B(n18268), .Z(n18104) );
  AND U18607 ( .A(n18269), .B(n18270), .Z(n18267) );
  AND U18608 ( .A(a[17]), .B(b[10]), .Z(n18266) );
  XOR U18609 ( .A(n18271), .B(n18109), .Z(n18111) );
  XOR U18610 ( .A(n18272), .B(n18273), .Z(n18109) );
  AND U18611 ( .A(n18274), .B(n18275), .Z(n18272) );
  AND U18612 ( .A(b[9]), .B(a[18]), .Z(n18271) );
  XOR U18613 ( .A(n18276), .B(n18114), .Z(n18116) );
  XOR U18614 ( .A(n18277), .B(n18278), .Z(n18114) );
  AND U18615 ( .A(n18279), .B(n18280), .Z(n18277) );
  AND U18616 ( .A(a[19]), .B(b[8]), .Z(n18276) );
  XOR U18617 ( .A(n18281), .B(n18119), .Z(n18121) );
  XOR U18618 ( .A(n18282), .B(n18283), .Z(n18119) );
  AND U18619 ( .A(n18284), .B(n18285), .Z(n18282) );
  AND U18620 ( .A(b[7]), .B(a[20]), .Z(n18281) );
  XOR U18621 ( .A(n18286), .B(n18124), .Z(n18126) );
  XOR U18622 ( .A(n18287), .B(n18288), .Z(n18124) );
  AND U18623 ( .A(n18289), .B(n18290), .Z(n18287) );
  AND U18624 ( .A(a[21]), .B(b[6]), .Z(n18286) );
  XOR U18625 ( .A(n18291), .B(n18129), .Z(n18131) );
  XOR U18626 ( .A(n18292), .B(n18293), .Z(n18129) );
  AND U18627 ( .A(n18294), .B(n18295), .Z(n18292) );
  AND U18628 ( .A(b[5]), .B(a[22]), .Z(n18291) );
  XOR U18629 ( .A(n18296), .B(n18134), .Z(n18136) );
  XOR U18630 ( .A(n18297), .B(n18298), .Z(n18134) );
  AND U18631 ( .A(n18299), .B(n18300), .Z(n18297) );
  AND U18632 ( .A(a[23]), .B(b[4]), .Z(n18296) );
  XNOR U18633 ( .A(n18301), .B(n18302), .Z(n18148) );
  NANDN U18634 ( .A(n18303), .B(n18304), .Z(n18302) );
  XOR U18635 ( .A(n18305), .B(n18139), .Z(n18141) );
  XNOR U18636 ( .A(n18306), .B(n18307), .Z(n18139) );
  AND U18637 ( .A(n18308), .B(n18309), .Z(n18306) );
  AND U18638 ( .A(b[3]), .B(a[24]), .Z(n18305) );
  XOR U18639 ( .A(n18155), .B(n18154), .Z(c[122]) );
  XOR U18640 ( .A(sreg[154]), .B(n18153), .Z(n18154) );
  XOR U18641 ( .A(n18160), .B(n18310), .Z(n18155) );
  XNOR U18642 ( .A(n18159), .B(n18153), .Z(n18310) );
  XOR U18643 ( .A(n18311), .B(n18312), .Z(n18153) );
  NOR U18644 ( .A(n18313), .B(n18314), .Z(n18311) );
  NAND U18645 ( .A(a[26]), .B(b[0]), .Z(n18159) );
  XNOR U18646 ( .A(n18303), .B(n18304), .Z(n18160) );
  XOR U18647 ( .A(n18301), .B(n18315), .Z(n18304) );
  NAND U18648 ( .A(a[25]), .B(b[1]), .Z(n18315) );
  XOR U18649 ( .A(n18309), .B(n18316), .Z(n18303) );
  XOR U18650 ( .A(n18301), .B(n18308), .Z(n18316) );
  XNOR U18651 ( .A(n18317), .B(n18307), .Z(n18308) );
  AND U18652 ( .A(b[2]), .B(a[24]), .Z(n18317) );
  NANDN U18653 ( .A(n18318), .B(n18319), .Z(n18301) );
  XOR U18654 ( .A(n18307), .B(n18299), .Z(n18320) );
  XNOR U18655 ( .A(n18298), .B(n18294), .Z(n18321) );
  XNOR U18656 ( .A(n18293), .B(n18289), .Z(n18322) );
  XNOR U18657 ( .A(n18288), .B(n18284), .Z(n18323) );
  XNOR U18658 ( .A(n18283), .B(n18279), .Z(n18324) );
  XNOR U18659 ( .A(n18278), .B(n18274), .Z(n18325) );
  XNOR U18660 ( .A(n18273), .B(n18269), .Z(n18326) );
  XNOR U18661 ( .A(n18268), .B(n18264), .Z(n18327) );
  XNOR U18662 ( .A(n18263), .B(n18259), .Z(n18328) );
  XNOR U18663 ( .A(n18258), .B(n18254), .Z(n18329) );
  XNOR U18664 ( .A(n18253), .B(n18249), .Z(n18330) );
  XNOR U18665 ( .A(n18248), .B(n18244), .Z(n18331) );
  XNOR U18666 ( .A(n18243), .B(n18239), .Z(n18332) );
  XNOR U18667 ( .A(n18238), .B(n18234), .Z(n18333) );
  XNOR U18668 ( .A(n18233), .B(n18229), .Z(n18334) );
  XNOR U18669 ( .A(n18228), .B(n18224), .Z(n18335) );
  XNOR U18670 ( .A(n18223), .B(n18219), .Z(n18336) );
  XNOR U18671 ( .A(n18218), .B(n18214), .Z(n18337) );
  XNOR U18672 ( .A(n18213), .B(n18209), .Z(n18338) );
  XNOR U18673 ( .A(n18208), .B(n18204), .Z(n18339) );
  XNOR U18674 ( .A(n18203), .B(n18199), .Z(n18340) );
  XNOR U18675 ( .A(n18198), .B(n18194), .Z(n18341) );
  XNOR U18676 ( .A(n18193), .B(n18189), .Z(n18342) );
  XNOR U18677 ( .A(n18343), .B(n18188), .Z(n18189) );
  AND U18678 ( .A(a[0]), .B(b[26]), .Z(n18343) );
  XNOR U18679 ( .A(n18344), .B(n18188), .Z(n18190) );
  XNOR U18680 ( .A(n18345), .B(n18346), .Z(n18188) );
  AND U18681 ( .A(n18347), .B(n18348), .Z(n18345) );
  AND U18682 ( .A(a[1]), .B(b[25]), .Z(n18344) );
  XOR U18683 ( .A(n18349), .B(n18193), .Z(n18195) );
  XOR U18684 ( .A(n18350), .B(n18351), .Z(n18193) );
  AND U18685 ( .A(n18352), .B(n18353), .Z(n18350) );
  AND U18686 ( .A(a[2]), .B(b[24]), .Z(n18349) );
  XOR U18687 ( .A(n18354), .B(n18198), .Z(n18200) );
  XOR U18688 ( .A(n18355), .B(n18356), .Z(n18198) );
  AND U18689 ( .A(n18357), .B(n18358), .Z(n18355) );
  AND U18690 ( .A(a[3]), .B(b[23]), .Z(n18354) );
  XOR U18691 ( .A(n18359), .B(n18203), .Z(n18205) );
  XOR U18692 ( .A(n18360), .B(n18361), .Z(n18203) );
  AND U18693 ( .A(n18362), .B(n18363), .Z(n18360) );
  AND U18694 ( .A(a[4]), .B(b[22]), .Z(n18359) );
  XOR U18695 ( .A(n18364), .B(n18208), .Z(n18210) );
  XOR U18696 ( .A(n18365), .B(n18366), .Z(n18208) );
  AND U18697 ( .A(n18367), .B(n18368), .Z(n18365) );
  AND U18698 ( .A(a[5]), .B(b[21]), .Z(n18364) );
  XOR U18699 ( .A(n18369), .B(n18213), .Z(n18215) );
  XOR U18700 ( .A(n18370), .B(n18371), .Z(n18213) );
  AND U18701 ( .A(n18372), .B(n18373), .Z(n18370) );
  AND U18702 ( .A(a[6]), .B(b[20]), .Z(n18369) );
  XOR U18703 ( .A(n18374), .B(n18218), .Z(n18220) );
  XOR U18704 ( .A(n18375), .B(n18376), .Z(n18218) );
  AND U18705 ( .A(n18377), .B(n18378), .Z(n18375) );
  AND U18706 ( .A(a[7]), .B(b[19]), .Z(n18374) );
  XOR U18707 ( .A(n18379), .B(n18223), .Z(n18225) );
  XOR U18708 ( .A(n18380), .B(n18381), .Z(n18223) );
  AND U18709 ( .A(n18382), .B(n18383), .Z(n18380) );
  AND U18710 ( .A(a[8]), .B(b[18]), .Z(n18379) );
  XOR U18711 ( .A(n18384), .B(n18228), .Z(n18230) );
  XOR U18712 ( .A(n18385), .B(n18386), .Z(n18228) );
  AND U18713 ( .A(n18387), .B(n18388), .Z(n18385) );
  AND U18714 ( .A(a[9]), .B(b[17]), .Z(n18384) );
  XOR U18715 ( .A(n18389), .B(n18233), .Z(n18235) );
  XOR U18716 ( .A(n18390), .B(n18391), .Z(n18233) );
  AND U18717 ( .A(n18392), .B(n18393), .Z(n18390) );
  AND U18718 ( .A(a[10]), .B(b[16]), .Z(n18389) );
  XOR U18719 ( .A(n18394), .B(n18238), .Z(n18240) );
  XOR U18720 ( .A(n18395), .B(n18396), .Z(n18238) );
  AND U18721 ( .A(n18397), .B(n18398), .Z(n18395) );
  AND U18722 ( .A(a[11]), .B(b[15]), .Z(n18394) );
  XOR U18723 ( .A(n18399), .B(n18243), .Z(n18245) );
  XOR U18724 ( .A(n18400), .B(n18401), .Z(n18243) );
  AND U18725 ( .A(n18402), .B(n18403), .Z(n18400) );
  AND U18726 ( .A(a[12]), .B(b[14]), .Z(n18399) );
  XOR U18727 ( .A(n18404), .B(n18248), .Z(n18250) );
  XOR U18728 ( .A(n18405), .B(n18406), .Z(n18248) );
  AND U18729 ( .A(n18407), .B(n18408), .Z(n18405) );
  AND U18730 ( .A(a[13]), .B(b[13]), .Z(n18404) );
  XOR U18731 ( .A(n18409), .B(n18253), .Z(n18255) );
  XOR U18732 ( .A(n18410), .B(n18411), .Z(n18253) );
  AND U18733 ( .A(n18412), .B(n18413), .Z(n18410) );
  AND U18734 ( .A(b[12]), .B(a[14]), .Z(n18409) );
  XOR U18735 ( .A(n18414), .B(n18258), .Z(n18260) );
  XOR U18736 ( .A(n18415), .B(n18416), .Z(n18258) );
  AND U18737 ( .A(n18417), .B(n18418), .Z(n18415) );
  AND U18738 ( .A(a[15]), .B(b[11]), .Z(n18414) );
  XOR U18739 ( .A(n18419), .B(n18263), .Z(n18265) );
  XOR U18740 ( .A(n18420), .B(n18421), .Z(n18263) );
  AND U18741 ( .A(n18422), .B(n18423), .Z(n18420) );
  AND U18742 ( .A(b[10]), .B(a[16]), .Z(n18419) );
  XOR U18743 ( .A(n18424), .B(n18268), .Z(n18270) );
  XOR U18744 ( .A(n18425), .B(n18426), .Z(n18268) );
  AND U18745 ( .A(n18427), .B(n18428), .Z(n18425) );
  AND U18746 ( .A(a[17]), .B(b[9]), .Z(n18424) );
  XOR U18747 ( .A(n18429), .B(n18273), .Z(n18275) );
  XOR U18748 ( .A(n18430), .B(n18431), .Z(n18273) );
  AND U18749 ( .A(n18432), .B(n18433), .Z(n18430) );
  AND U18750 ( .A(b[8]), .B(a[18]), .Z(n18429) );
  XOR U18751 ( .A(n18434), .B(n18278), .Z(n18280) );
  XOR U18752 ( .A(n18435), .B(n18436), .Z(n18278) );
  AND U18753 ( .A(n18437), .B(n18438), .Z(n18435) );
  AND U18754 ( .A(a[19]), .B(b[7]), .Z(n18434) );
  XOR U18755 ( .A(n18439), .B(n18283), .Z(n18285) );
  XOR U18756 ( .A(n18440), .B(n18441), .Z(n18283) );
  AND U18757 ( .A(n18442), .B(n18443), .Z(n18440) );
  AND U18758 ( .A(b[6]), .B(a[20]), .Z(n18439) );
  XOR U18759 ( .A(n18444), .B(n18288), .Z(n18290) );
  XOR U18760 ( .A(n18445), .B(n18446), .Z(n18288) );
  AND U18761 ( .A(n18447), .B(n18448), .Z(n18445) );
  AND U18762 ( .A(a[21]), .B(b[5]), .Z(n18444) );
  XOR U18763 ( .A(n18449), .B(n18293), .Z(n18295) );
  XOR U18764 ( .A(n18450), .B(n18451), .Z(n18293) );
  AND U18765 ( .A(n18452), .B(n18453), .Z(n18450) );
  AND U18766 ( .A(b[4]), .B(a[22]), .Z(n18449) );
  XNOR U18767 ( .A(n18454), .B(n18455), .Z(n18307) );
  NANDN U18768 ( .A(n18456), .B(n18457), .Z(n18455) );
  XOR U18769 ( .A(n18458), .B(n18298), .Z(n18300) );
  XNOR U18770 ( .A(n18459), .B(n18460), .Z(n18298) );
  AND U18771 ( .A(n18461), .B(n18462), .Z(n18459) );
  AND U18772 ( .A(a[23]), .B(b[3]), .Z(n18458) );
  XOR U18773 ( .A(n18314), .B(n18313), .Z(c[121]) );
  XOR U18774 ( .A(sreg[153]), .B(n18312), .Z(n18313) );
  XOR U18775 ( .A(n18319), .B(n18463), .Z(n18314) );
  XNOR U18776 ( .A(n18318), .B(n18312), .Z(n18463) );
  XOR U18777 ( .A(n18464), .B(n18465), .Z(n18312) );
  NOR U18778 ( .A(n18466), .B(n18467), .Z(n18464) );
  NAND U18779 ( .A(a[25]), .B(b[0]), .Z(n18318) );
  XNOR U18780 ( .A(n18456), .B(n18457), .Z(n18319) );
  XOR U18781 ( .A(n18454), .B(n18468), .Z(n18457) );
  NAND U18782 ( .A(b[1]), .B(a[24]), .Z(n18468) );
  XOR U18783 ( .A(n18462), .B(n18469), .Z(n18456) );
  XOR U18784 ( .A(n18454), .B(n18461), .Z(n18469) );
  XNOR U18785 ( .A(n18470), .B(n18460), .Z(n18461) );
  AND U18786 ( .A(b[2]), .B(a[23]), .Z(n18470) );
  NANDN U18787 ( .A(n18471), .B(n18472), .Z(n18454) );
  XOR U18788 ( .A(n18460), .B(n18452), .Z(n18473) );
  XNOR U18789 ( .A(n18451), .B(n18447), .Z(n18474) );
  XNOR U18790 ( .A(n18446), .B(n18442), .Z(n18475) );
  XNOR U18791 ( .A(n18441), .B(n18437), .Z(n18476) );
  XNOR U18792 ( .A(n18436), .B(n18432), .Z(n18477) );
  XNOR U18793 ( .A(n18431), .B(n18427), .Z(n18478) );
  XNOR U18794 ( .A(n18426), .B(n18422), .Z(n18479) );
  XNOR U18795 ( .A(n18421), .B(n18417), .Z(n18480) );
  XNOR U18796 ( .A(n18416), .B(n18412), .Z(n18481) );
  XNOR U18797 ( .A(n18411), .B(n18407), .Z(n18482) );
  XNOR U18798 ( .A(n18406), .B(n18402), .Z(n18483) );
  XNOR U18799 ( .A(n18401), .B(n18397), .Z(n18484) );
  XNOR U18800 ( .A(n18396), .B(n18392), .Z(n18485) );
  XNOR U18801 ( .A(n18391), .B(n18387), .Z(n18486) );
  XNOR U18802 ( .A(n18386), .B(n18382), .Z(n18487) );
  XNOR U18803 ( .A(n18381), .B(n18377), .Z(n18488) );
  XNOR U18804 ( .A(n18376), .B(n18372), .Z(n18489) );
  XNOR U18805 ( .A(n18371), .B(n18367), .Z(n18490) );
  XNOR U18806 ( .A(n18366), .B(n18362), .Z(n18491) );
  XNOR U18807 ( .A(n18361), .B(n18357), .Z(n18492) );
  XNOR U18808 ( .A(n18356), .B(n18352), .Z(n18493) );
  XNOR U18809 ( .A(n18351), .B(n18347), .Z(n18494) );
  XOR U18810 ( .A(n18495), .B(n18346), .Z(n18347) );
  AND U18811 ( .A(a[0]), .B(b[25]), .Z(n18495) );
  XOR U18812 ( .A(n18496), .B(n18346), .Z(n18348) );
  XNOR U18813 ( .A(n18497), .B(n18498), .Z(n18346) );
  AND U18814 ( .A(n18499), .B(n18500), .Z(n18497) );
  AND U18815 ( .A(a[1]), .B(b[24]), .Z(n18496) );
  XOR U18816 ( .A(n18501), .B(n18351), .Z(n18353) );
  XOR U18817 ( .A(n18502), .B(n18503), .Z(n18351) );
  AND U18818 ( .A(n18504), .B(n18505), .Z(n18502) );
  AND U18819 ( .A(a[2]), .B(b[23]), .Z(n18501) );
  XOR U18820 ( .A(n18506), .B(n18356), .Z(n18358) );
  XOR U18821 ( .A(n18507), .B(n18508), .Z(n18356) );
  AND U18822 ( .A(n18509), .B(n18510), .Z(n18507) );
  AND U18823 ( .A(a[3]), .B(b[22]), .Z(n18506) );
  XOR U18824 ( .A(n18511), .B(n18361), .Z(n18363) );
  XOR U18825 ( .A(n18512), .B(n18513), .Z(n18361) );
  AND U18826 ( .A(n18514), .B(n18515), .Z(n18512) );
  AND U18827 ( .A(a[4]), .B(b[21]), .Z(n18511) );
  XOR U18828 ( .A(n18516), .B(n18366), .Z(n18368) );
  XOR U18829 ( .A(n18517), .B(n18518), .Z(n18366) );
  AND U18830 ( .A(n18519), .B(n18520), .Z(n18517) );
  AND U18831 ( .A(a[5]), .B(b[20]), .Z(n18516) );
  XOR U18832 ( .A(n18521), .B(n18371), .Z(n18373) );
  XOR U18833 ( .A(n18522), .B(n18523), .Z(n18371) );
  AND U18834 ( .A(n18524), .B(n18525), .Z(n18522) );
  AND U18835 ( .A(a[6]), .B(b[19]), .Z(n18521) );
  XOR U18836 ( .A(n18526), .B(n18376), .Z(n18378) );
  XOR U18837 ( .A(n18527), .B(n18528), .Z(n18376) );
  AND U18838 ( .A(n18529), .B(n18530), .Z(n18527) );
  AND U18839 ( .A(a[7]), .B(b[18]), .Z(n18526) );
  XOR U18840 ( .A(n18531), .B(n18381), .Z(n18383) );
  XOR U18841 ( .A(n18532), .B(n18533), .Z(n18381) );
  AND U18842 ( .A(n18534), .B(n18535), .Z(n18532) );
  AND U18843 ( .A(a[8]), .B(b[17]), .Z(n18531) );
  XOR U18844 ( .A(n18536), .B(n18386), .Z(n18388) );
  XOR U18845 ( .A(n18537), .B(n18538), .Z(n18386) );
  AND U18846 ( .A(n18539), .B(n18540), .Z(n18537) );
  AND U18847 ( .A(a[9]), .B(b[16]), .Z(n18536) );
  XOR U18848 ( .A(n18541), .B(n18391), .Z(n18393) );
  XOR U18849 ( .A(n18542), .B(n18543), .Z(n18391) );
  AND U18850 ( .A(n18544), .B(n18545), .Z(n18542) );
  AND U18851 ( .A(a[10]), .B(b[15]), .Z(n18541) );
  XOR U18852 ( .A(n18546), .B(n18396), .Z(n18398) );
  XOR U18853 ( .A(n18547), .B(n18548), .Z(n18396) );
  AND U18854 ( .A(n18549), .B(n18550), .Z(n18547) );
  AND U18855 ( .A(a[11]), .B(b[14]), .Z(n18546) );
  XOR U18856 ( .A(n18551), .B(n18401), .Z(n18403) );
  XOR U18857 ( .A(n18552), .B(n18553), .Z(n18401) );
  AND U18858 ( .A(n18554), .B(n18555), .Z(n18552) );
  AND U18859 ( .A(a[12]), .B(b[13]), .Z(n18551) );
  XOR U18860 ( .A(n18556), .B(n18406), .Z(n18408) );
  XOR U18861 ( .A(n18557), .B(n18558), .Z(n18406) );
  AND U18862 ( .A(n18559), .B(n18560), .Z(n18557) );
  AND U18863 ( .A(a[13]), .B(b[12]), .Z(n18556) );
  XOR U18864 ( .A(n18561), .B(n18411), .Z(n18413) );
  XOR U18865 ( .A(n18562), .B(n18563), .Z(n18411) );
  AND U18866 ( .A(n18564), .B(n18565), .Z(n18562) );
  AND U18867 ( .A(b[11]), .B(a[14]), .Z(n18561) );
  XOR U18868 ( .A(n18566), .B(n18416), .Z(n18418) );
  XOR U18869 ( .A(n18567), .B(n18568), .Z(n18416) );
  AND U18870 ( .A(n18569), .B(n18570), .Z(n18567) );
  AND U18871 ( .A(a[15]), .B(b[10]), .Z(n18566) );
  XOR U18872 ( .A(n18571), .B(n18421), .Z(n18423) );
  XOR U18873 ( .A(n18572), .B(n18573), .Z(n18421) );
  AND U18874 ( .A(n18574), .B(n18575), .Z(n18572) );
  AND U18875 ( .A(b[9]), .B(a[16]), .Z(n18571) );
  XOR U18876 ( .A(n18576), .B(n18426), .Z(n18428) );
  XOR U18877 ( .A(n18577), .B(n18578), .Z(n18426) );
  AND U18878 ( .A(n18579), .B(n18580), .Z(n18577) );
  AND U18879 ( .A(a[17]), .B(b[8]), .Z(n18576) );
  XOR U18880 ( .A(n18581), .B(n18431), .Z(n18433) );
  XOR U18881 ( .A(n18582), .B(n18583), .Z(n18431) );
  AND U18882 ( .A(n18584), .B(n18585), .Z(n18582) );
  AND U18883 ( .A(b[7]), .B(a[18]), .Z(n18581) );
  XOR U18884 ( .A(n18586), .B(n18436), .Z(n18438) );
  XOR U18885 ( .A(n18587), .B(n18588), .Z(n18436) );
  AND U18886 ( .A(n18589), .B(n18590), .Z(n18587) );
  AND U18887 ( .A(a[19]), .B(b[6]), .Z(n18586) );
  XOR U18888 ( .A(n18591), .B(n18441), .Z(n18443) );
  XOR U18889 ( .A(n18592), .B(n18593), .Z(n18441) );
  AND U18890 ( .A(n18594), .B(n18595), .Z(n18592) );
  AND U18891 ( .A(b[5]), .B(a[20]), .Z(n18591) );
  XOR U18892 ( .A(n18596), .B(n18446), .Z(n18448) );
  XOR U18893 ( .A(n18597), .B(n18598), .Z(n18446) );
  AND U18894 ( .A(n18599), .B(n18600), .Z(n18597) );
  AND U18895 ( .A(a[21]), .B(b[4]), .Z(n18596) );
  XNOR U18896 ( .A(n18601), .B(n18602), .Z(n18460) );
  NANDN U18897 ( .A(n18603), .B(n18604), .Z(n18602) );
  XOR U18898 ( .A(n18605), .B(n18451), .Z(n18453) );
  XNOR U18899 ( .A(n18606), .B(n18607), .Z(n18451) );
  AND U18900 ( .A(n18608), .B(n18609), .Z(n18606) );
  AND U18901 ( .A(b[3]), .B(a[22]), .Z(n18605) );
  XOR U18902 ( .A(n18467), .B(n18466), .Z(c[120]) );
  XOR U18903 ( .A(sreg[152]), .B(n18465), .Z(n18466) );
  XOR U18904 ( .A(n18472), .B(n18610), .Z(n18467) );
  XNOR U18905 ( .A(n18471), .B(n18465), .Z(n18610) );
  XOR U18906 ( .A(n18611), .B(n18612), .Z(n18465) );
  NOR U18907 ( .A(n18613), .B(n18614), .Z(n18611) );
  NAND U18908 ( .A(a[24]), .B(b[0]), .Z(n18471) );
  XNOR U18909 ( .A(n18603), .B(n18604), .Z(n18472) );
  XOR U18910 ( .A(n18601), .B(n18615), .Z(n18604) );
  NAND U18911 ( .A(a[23]), .B(b[1]), .Z(n18615) );
  XOR U18912 ( .A(n18609), .B(n18616), .Z(n18603) );
  XOR U18913 ( .A(n18601), .B(n18608), .Z(n18616) );
  XNOR U18914 ( .A(n18617), .B(n18607), .Z(n18608) );
  AND U18915 ( .A(b[2]), .B(a[22]), .Z(n18617) );
  NANDN U18916 ( .A(n18618), .B(n18619), .Z(n18601) );
  XOR U18917 ( .A(n18607), .B(n18599), .Z(n18620) );
  XNOR U18918 ( .A(n18598), .B(n18594), .Z(n18621) );
  XNOR U18919 ( .A(n18593), .B(n18589), .Z(n18622) );
  XNOR U18920 ( .A(n18588), .B(n18584), .Z(n18623) );
  XNOR U18921 ( .A(n18583), .B(n18579), .Z(n18624) );
  XNOR U18922 ( .A(n18578), .B(n18574), .Z(n18625) );
  XNOR U18923 ( .A(n18573), .B(n18569), .Z(n18626) );
  XNOR U18924 ( .A(n18568), .B(n18564), .Z(n18627) );
  XNOR U18925 ( .A(n18563), .B(n18559), .Z(n18628) );
  XNOR U18926 ( .A(n18558), .B(n18554), .Z(n18629) );
  XNOR U18927 ( .A(n18553), .B(n18549), .Z(n18630) );
  XNOR U18928 ( .A(n18548), .B(n18544), .Z(n18631) );
  XNOR U18929 ( .A(n18543), .B(n18539), .Z(n18632) );
  XNOR U18930 ( .A(n18538), .B(n18534), .Z(n18633) );
  XNOR U18931 ( .A(n18533), .B(n18529), .Z(n18634) );
  XNOR U18932 ( .A(n18528), .B(n18524), .Z(n18635) );
  XNOR U18933 ( .A(n18523), .B(n18519), .Z(n18636) );
  XNOR U18934 ( .A(n18518), .B(n18514), .Z(n18637) );
  XNOR U18935 ( .A(n18513), .B(n18509), .Z(n18638) );
  XNOR U18936 ( .A(n18508), .B(n18504), .Z(n18639) );
  XNOR U18937 ( .A(n18503), .B(n18499), .Z(n18640) );
  XNOR U18938 ( .A(n18641), .B(n18498), .Z(n18499) );
  AND U18939 ( .A(a[0]), .B(b[24]), .Z(n18641) );
  XNOR U18940 ( .A(n18642), .B(n18498), .Z(n18500) );
  XNOR U18941 ( .A(n18643), .B(n18644), .Z(n18498) );
  AND U18942 ( .A(n18645), .B(n18646), .Z(n18643) );
  AND U18943 ( .A(a[1]), .B(b[23]), .Z(n18642) );
  XOR U18944 ( .A(n18647), .B(n18503), .Z(n18505) );
  XOR U18945 ( .A(n18648), .B(n18649), .Z(n18503) );
  AND U18946 ( .A(n18650), .B(n18651), .Z(n18648) );
  AND U18947 ( .A(a[2]), .B(b[22]), .Z(n18647) );
  XOR U18948 ( .A(n18652), .B(n18508), .Z(n18510) );
  XOR U18949 ( .A(n18653), .B(n18654), .Z(n18508) );
  AND U18950 ( .A(n18655), .B(n18656), .Z(n18653) );
  AND U18951 ( .A(a[3]), .B(b[21]), .Z(n18652) );
  XOR U18952 ( .A(n18657), .B(n18513), .Z(n18515) );
  XOR U18953 ( .A(n18658), .B(n18659), .Z(n18513) );
  AND U18954 ( .A(n18660), .B(n18661), .Z(n18658) );
  AND U18955 ( .A(a[4]), .B(b[20]), .Z(n18657) );
  XOR U18956 ( .A(n18662), .B(n18518), .Z(n18520) );
  XOR U18957 ( .A(n18663), .B(n18664), .Z(n18518) );
  AND U18958 ( .A(n18665), .B(n18666), .Z(n18663) );
  AND U18959 ( .A(a[5]), .B(b[19]), .Z(n18662) );
  XOR U18960 ( .A(n18667), .B(n18523), .Z(n18525) );
  XOR U18961 ( .A(n18668), .B(n18669), .Z(n18523) );
  AND U18962 ( .A(n18670), .B(n18671), .Z(n18668) );
  AND U18963 ( .A(a[6]), .B(b[18]), .Z(n18667) );
  XOR U18964 ( .A(n18672), .B(n18528), .Z(n18530) );
  XOR U18965 ( .A(n18673), .B(n18674), .Z(n18528) );
  AND U18966 ( .A(n18675), .B(n18676), .Z(n18673) );
  AND U18967 ( .A(a[7]), .B(b[17]), .Z(n18672) );
  XOR U18968 ( .A(n18677), .B(n18533), .Z(n18535) );
  XOR U18969 ( .A(n18678), .B(n18679), .Z(n18533) );
  AND U18970 ( .A(n18680), .B(n18681), .Z(n18678) );
  AND U18971 ( .A(a[8]), .B(b[16]), .Z(n18677) );
  XOR U18972 ( .A(n18682), .B(n18538), .Z(n18540) );
  XOR U18973 ( .A(n18683), .B(n18684), .Z(n18538) );
  AND U18974 ( .A(n18685), .B(n18686), .Z(n18683) );
  AND U18975 ( .A(a[9]), .B(b[15]), .Z(n18682) );
  XOR U18976 ( .A(n18687), .B(n18543), .Z(n18545) );
  XOR U18977 ( .A(n18688), .B(n18689), .Z(n18543) );
  AND U18978 ( .A(n18690), .B(n18691), .Z(n18688) );
  AND U18979 ( .A(a[10]), .B(b[14]), .Z(n18687) );
  XOR U18980 ( .A(n18692), .B(n18548), .Z(n18550) );
  XOR U18981 ( .A(n18693), .B(n18694), .Z(n18548) );
  AND U18982 ( .A(n18695), .B(n18696), .Z(n18693) );
  AND U18983 ( .A(a[11]), .B(b[13]), .Z(n18692) );
  XOR U18984 ( .A(n18697), .B(n18553), .Z(n18555) );
  XOR U18985 ( .A(n18698), .B(n18699), .Z(n18553) );
  AND U18986 ( .A(n18700), .B(n18701), .Z(n18698) );
  AND U18987 ( .A(b[12]), .B(a[12]), .Z(n18697) );
  XOR U18988 ( .A(n18702), .B(n18558), .Z(n18560) );
  XOR U18989 ( .A(n18703), .B(n18704), .Z(n18558) );
  AND U18990 ( .A(n18705), .B(n18706), .Z(n18703) );
  AND U18991 ( .A(a[13]), .B(b[11]), .Z(n18702) );
  XOR U18992 ( .A(n18707), .B(n18563), .Z(n18565) );
  XOR U18993 ( .A(n18708), .B(n18709), .Z(n18563) );
  AND U18994 ( .A(n18710), .B(n18711), .Z(n18708) );
  AND U18995 ( .A(b[10]), .B(a[14]), .Z(n18707) );
  XOR U18996 ( .A(n18712), .B(n18568), .Z(n18570) );
  XOR U18997 ( .A(n18713), .B(n18714), .Z(n18568) );
  AND U18998 ( .A(n18715), .B(n18716), .Z(n18713) );
  AND U18999 ( .A(a[15]), .B(b[9]), .Z(n18712) );
  XOR U19000 ( .A(n18717), .B(n18573), .Z(n18575) );
  XOR U19001 ( .A(n18718), .B(n18719), .Z(n18573) );
  AND U19002 ( .A(n18720), .B(n18721), .Z(n18718) );
  AND U19003 ( .A(b[8]), .B(a[16]), .Z(n18717) );
  XOR U19004 ( .A(n18722), .B(n18578), .Z(n18580) );
  XOR U19005 ( .A(n18723), .B(n18724), .Z(n18578) );
  AND U19006 ( .A(n18725), .B(n18726), .Z(n18723) );
  AND U19007 ( .A(a[17]), .B(b[7]), .Z(n18722) );
  XOR U19008 ( .A(n18727), .B(n18583), .Z(n18585) );
  XOR U19009 ( .A(n18728), .B(n18729), .Z(n18583) );
  AND U19010 ( .A(n18730), .B(n18731), .Z(n18728) );
  AND U19011 ( .A(b[6]), .B(a[18]), .Z(n18727) );
  XOR U19012 ( .A(n18732), .B(n18588), .Z(n18590) );
  XOR U19013 ( .A(n18733), .B(n18734), .Z(n18588) );
  AND U19014 ( .A(n18735), .B(n18736), .Z(n18733) );
  AND U19015 ( .A(a[19]), .B(b[5]), .Z(n18732) );
  XOR U19016 ( .A(n18737), .B(n18593), .Z(n18595) );
  XOR U19017 ( .A(n18738), .B(n18739), .Z(n18593) );
  AND U19018 ( .A(n18740), .B(n18741), .Z(n18738) );
  AND U19019 ( .A(b[4]), .B(a[20]), .Z(n18737) );
  XNOR U19020 ( .A(n18742), .B(n18743), .Z(n18607) );
  NANDN U19021 ( .A(n18744), .B(n18745), .Z(n18743) );
  XOR U19022 ( .A(n18746), .B(n18598), .Z(n18600) );
  XNOR U19023 ( .A(n18747), .B(n18748), .Z(n18598) );
  AND U19024 ( .A(n18749), .B(n18750), .Z(n18747) );
  AND U19025 ( .A(a[21]), .B(b[3]), .Z(n18746) );
  XOR U19026 ( .A(n18614), .B(n18613), .Z(c[119]) );
  XOR U19027 ( .A(sreg[151]), .B(n18612), .Z(n18613) );
  XOR U19028 ( .A(n18619), .B(n18751), .Z(n18614) );
  XNOR U19029 ( .A(n18618), .B(n18612), .Z(n18751) );
  XOR U19030 ( .A(n18752), .B(n18753), .Z(n18612) );
  NOR U19031 ( .A(n18754), .B(n18755), .Z(n18752) );
  NAND U19032 ( .A(a[23]), .B(b[0]), .Z(n18618) );
  XNOR U19033 ( .A(n18744), .B(n18745), .Z(n18619) );
  XOR U19034 ( .A(n18742), .B(n18756), .Z(n18745) );
  NAND U19035 ( .A(b[1]), .B(a[22]), .Z(n18756) );
  XOR U19036 ( .A(n18750), .B(n18757), .Z(n18744) );
  XOR U19037 ( .A(n18742), .B(n18749), .Z(n18757) );
  XNOR U19038 ( .A(n18758), .B(n18748), .Z(n18749) );
  AND U19039 ( .A(b[2]), .B(a[21]), .Z(n18758) );
  NANDN U19040 ( .A(n18759), .B(n18760), .Z(n18742) );
  XOR U19041 ( .A(n18748), .B(n18740), .Z(n18761) );
  XNOR U19042 ( .A(n18739), .B(n18735), .Z(n18762) );
  XNOR U19043 ( .A(n18734), .B(n18730), .Z(n18763) );
  XNOR U19044 ( .A(n18729), .B(n18725), .Z(n18764) );
  XNOR U19045 ( .A(n18724), .B(n18720), .Z(n18765) );
  XNOR U19046 ( .A(n18719), .B(n18715), .Z(n18766) );
  XNOR U19047 ( .A(n18714), .B(n18710), .Z(n18767) );
  XNOR U19048 ( .A(n18709), .B(n18705), .Z(n18768) );
  XNOR U19049 ( .A(n18704), .B(n18700), .Z(n18769) );
  XNOR U19050 ( .A(n18699), .B(n18695), .Z(n18770) );
  XNOR U19051 ( .A(n18694), .B(n18690), .Z(n18771) );
  XNOR U19052 ( .A(n18689), .B(n18685), .Z(n18772) );
  XNOR U19053 ( .A(n18684), .B(n18680), .Z(n18773) );
  XNOR U19054 ( .A(n18679), .B(n18675), .Z(n18774) );
  XNOR U19055 ( .A(n18674), .B(n18670), .Z(n18775) );
  XNOR U19056 ( .A(n18669), .B(n18665), .Z(n18776) );
  XNOR U19057 ( .A(n18664), .B(n18660), .Z(n18777) );
  XNOR U19058 ( .A(n18659), .B(n18655), .Z(n18778) );
  XNOR U19059 ( .A(n18654), .B(n18650), .Z(n18779) );
  XNOR U19060 ( .A(n18649), .B(n18645), .Z(n18780) );
  XOR U19061 ( .A(n18781), .B(n18644), .Z(n18645) );
  AND U19062 ( .A(a[0]), .B(b[23]), .Z(n18781) );
  XOR U19063 ( .A(n18782), .B(n18644), .Z(n18646) );
  XNOR U19064 ( .A(n18783), .B(n18784), .Z(n18644) );
  AND U19065 ( .A(n18785), .B(n18786), .Z(n18783) );
  AND U19066 ( .A(a[1]), .B(b[22]), .Z(n18782) );
  XOR U19067 ( .A(n18787), .B(n18649), .Z(n18651) );
  XOR U19068 ( .A(n18788), .B(n18789), .Z(n18649) );
  AND U19069 ( .A(n18790), .B(n18791), .Z(n18788) );
  AND U19070 ( .A(a[2]), .B(b[21]), .Z(n18787) );
  XOR U19071 ( .A(n18792), .B(n18654), .Z(n18656) );
  XOR U19072 ( .A(n18793), .B(n18794), .Z(n18654) );
  AND U19073 ( .A(n18795), .B(n18796), .Z(n18793) );
  AND U19074 ( .A(a[3]), .B(b[20]), .Z(n18792) );
  XOR U19075 ( .A(n18797), .B(n18659), .Z(n18661) );
  XOR U19076 ( .A(n18798), .B(n18799), .Z(n18659) );
  AND U19077 ( .A(n18800), .B(n18801), .Z(n18798) );
  AND U19078 ( .A(a[4]), .B(b[19]), .Z(n18797) );
  XOR U19079 ( .A(n18802), .B(n18664), .Z(n18666) );
  XOR U19080 ( .A(n18803), .B(n18804), .Z(n18664) );
  AND U19081 ( .A(n18805), .B(n18806), .Z(n18803) );
  AND U19082 ( .A(a[5]), .B(b[18]), .Z(n18802) );
  XOR U19083 ( .A(n18807), .B(n18669), .Z(n18671) );
  XOR U19084 ( .A(n18808), .B(n18809), .Z(n18669) );
  AND U19085 ( .A(n18810), .B(n18811), .Z(n18808) );
  AND U19086 ( .A(a[6]), .B(b[17]), .Z(n18807) );
  XOR U19087 ( .A(n18812), .B(n18674), .Z(n18676) );
  XOR U19088 ( .A(n18813), .B(n18814), .Z(n18674) );
  AND U19089 ( .A(n18815), .B(n18816), .Z(n18813) );
  AND U19090 ( .A(a[7]), .B(b[16]), .Z(n18812) );
  XOR U19091 ( .A(n18817), .B(n18679), .Z(n18681) );
  XOR U19092 ( .A(n18818), .B(n18819), .Z(n18679) );
  AND U19093 ( .A(n18820), .B(n18821), .Z(n18818) );
  AND U19094 ( .A(a[8]), .B(b[15]), .Z(n18817) );
  XOR U19095 ( .A(n18822), .B(n18684), .Z(n18686) );
  XOR U19096 ( .A(n18823), .B(n18824), .Z(n18684) );
  AND U19097 ( .A(n18825), .B(n18826), .Z(n18823) );
  AND U19098 ( .A(a[9]), .B(b[14]), .Z(n18822) );
  XOR U19099 ( .A(n18827), .B(n18689), .Z(n18691) );
  XOR U19100 ( .A(n18828), .B(n18829), .Z(n18689) );
  AND U19101 ( .A(n18830), .B(n18831), .Z(n18828) );
  AND U19102 ( .A(a[10]), .B(b[13]), .Z(n18827) );
  XOR U19103 ( .A(n18832), .B(n18694), .Z(n18696) );
  XOR U19104 ( .A(n18833), .B(n18834), .Z(n18694) );
  AND U19105 ( .A(n18835), .B(n18836), .Z(n18833) );
  AND U19106 ( .A(a[11]), .B(b[12]), .Z(n18832) );
  XOR U19107 ( .A(n18837), .B(n18699), .Z(n18701) );
  XOR U19108 ( .A(n18838), .B(n18839), .Z(n18699) );
  AND U19109 ( .A(n18840), .B(n18841), .Z(n18838) );
  AND U19110 ( .A(b[11]), .B(a[12]), .Z(n18837) );
  XOR U19111 ( .A(n18842), .B(n18704), .Z(n18706) );
  XOR U19112 ( .A(n18843), .B(n18844), .Z(n18704) );
  AND U19113 ( .A(n18845), .B(n18846), .Z(n18843) );
  AND U19114 ( .A(a[13]), .B(b[10]), .Z(n18842) );
  XOR U19115 ( .A(n18847), .B(n18709), .Z(n18711) );
  XOR U19116 ( .A(n18848), .B(n18849), .Z(n18709) );
  AND U19117 ( .A(n18850), .B(n18851), .Z(n18848) );
  AND U19118 ( .A(b[9]), .B(a[14]), .Z(n18847) );
  XOR U19119 ( .A(n18852), .B(n18714), .Z(n18716) );
  XOR U19120 ( .A(n18853), .B(n18854), .Z(n18714) );
  AND U19121 ( .A(n18855), .B(n18856), .Z(n18853) );
  AND U19122 ( .A(a[15]), .B(b[8]), .Z(n18852) );
  XOR U19123 ( .A(n18857), .B(n18719), .Z(n18721) );
  XOR U19124 ( .A(n18858), .B(n18859), .Z(n18719) );
  AND U19125 ( .A(n18860), .B(n18861), .Z(n18858) );
  AND U19126 ( .A(b[7]), .B(a[16]), .Z(n18857) );
  XOR U19127 ( .A(n18862), .B(n18724), .Z(n18726) );
  XOR U19128 ( .A(n18863), .B(n18864), .Z(n18724) );
  AND U19129 ( .A(n18865), .B(n18866), .Z(n18863) );
  AND U19130 ( .A(a[17]), .B(b[6]), .Z(n18862) );
  XOR U19131 ( .A(n18867), .B(n18729), .Z(n18731) );
  XOR U19132 ( .A(n18868), .B(n18869), .Z(n18729) );
  AND U19133 ( .A(n18870), .B(n18871), .Z(n18868) );
  AND U19134 ( .A(b[5]), .B(a[18]), .Z(n18867) );
  XOR U19135 ( .A(n18872), .B(n18734), .Z(n18736) );
  XOR U19136 ( .A(n18873), .B(n18874), .Z(n18734) );
  AND U19137 ( .A(n18875), .B(n18876), .Z(n18873) );
  AND U19138 ( .A(a[19]), .B(b[4]), .Z(n18872) );
  XNOR U19139 ( .A(n18877), .B(n18878), .Z(n18748) );
  NANDN U19140 ( .A(n18879), .B(n18880), .Z(n18878) );
  XOR U19141 ( .A(n18881), .B(n18739), .Z(n18741) );
  XNOR U19142 ( .A(n18882), .B(n18883), .Z(n18739) );
  AND U19143 ( .A(n18884), .B(n18885), .Z(n18882) );
  AND U19144 ( .A(b[3]), .B(a[20]), .Z(n18881) );
  XOR U19145 ( .A(n18755), .B(n18754), .Z(c[118]) );
  XOR U19146 ( .A(sreg[150]), .B(n18753), .Z(n18754) );
  XOR U19147 ( .A(n18760), .B(n18886), .Z(n18755) );
  XNOR U19148 ( .A(n18759), .B(n18753), .Z(n18886) );
  XOR U19149 ( .A(n18887), .B(n18888), .Z(n18753) );
  NOR U19150 ( .A(n18889), .B(n18890), .Z(n18887) );
  NAND U19151 ( .A(a[22]), .B(b[0]), .Z(n18759) );
  XNOR U19152 ( .A(n18879), .B(n18880), .Z(n18760) );
  XOR U19153 ( .A(n18877), .B(n18891), .Z(n18880) );
  NAND U19154 ( .A(a[21]), .B(b[1]), .Z(n18891) );
  XOR U19155 ( .A(n18885), .B(n18892), .Z(n18879) );
  XOR U19156 ( .A(n18877), .B(n18884), .Z(n18892) );
  XNOR U19157 ( .A(n18893), .B(n18883), .Z(n18884) );
  AND U19158 ( .A(b[2]), .B(a[20]), .Z(n18893) );
  NANDN U19159 ( .A(n18894), .B(n18895), .Z(n18877) );
  XOR U19160 ( .A(n18883), .B(n18875), .Z(n18896) );
  XNOR U19161 ( .A(n18874), .B(n18870), .Z(n18897) );
  XNOR U19162 ( .A(n18869), .B(n18865), .Z(n18898) );
  XNOR U19163 ( .A(n18864), .B(n18860), .Z(n18899) );
  XNOR U19164 ( .A(n18859), .B(n18855), .Z(n18900) );
  XNOR U19165 ( .A(n18854), .B(n18850), .Z(n18901) );
  XNOR U19166 ( .A(n18849), .B(n18845), .Z(n18902) );
  XNOR U19167 ( .A(n18844), .B(n18840), .Z(n18903) );
  XNOR U19168 ( .A(n18839), .B(n18835), .Z(n18904) );
  XNOR U19169 ( .A(n18834), .B(n18830), .Z(n18905) );
  XNOR U19170 ( .A(n18829), .B(n18825), .Z(n18906) );
  XNOR U19171 ( .A(n18824), .B(n18820), .Z(n18907) );
  XNOR U19172 ( .A(n18819), .B(n18815), .Z(n18908) );
  XNOR U19173 ( .A(n18814), .B(n18810), .Z(n18909) );
  XNOR U19174 ( .A(n18809), .B(n18805), .Z(n18910) );
  XNOR U19175 ( .A(n18804), .B(n18800), .Z(n18911) );
  XNOR U19176 ( .A(n18799), .B(n18795), .Z(n18912) );
  XNOR U19177 ( .A(n18794), .B(n18790), .Z(n18913) );
  XNOR U19178 ( .A(n18789), .B(n18785), .Z(n18914) );
  XNOR U19179 ( .A(n18915), .B(n18784), .Z(n18785) );
  AND U19180 ( .A(a[0]), .B(b[22]), .Z(n18915) );
  XNOR U19181 ( .A(n18916), .B(n18784), .Z(n18786) );
  XNOR U19182 ( .A(n18917), .B(n18918), .Z(n18784) );
  AND U19183 ( .A(n18919), .B(n18920), .Z(n18917) );
  AND U19184 ( .A(a[1]), .B(b[21]), .Z(n18916) );
  XOR U19185 ( .A(n18921), .B(n18789), .Z(n18791) );
  XOR U19186 ( .A(n18922), .B(n18923), .Z(n18789) );
  AND U19187 ( .A(n18924), .B(n18925), .Z(n18922) );
  AND U19188 ( .A(a[2]), .B(b[20]), .Z(n18921) );
  XOR U19189 ( .A(n18926), .B(n18794), .Z(n18796) );
  XOR U19190 ( .A(n18927), .B(n18928), .Z(n18794) );
  AND U19191 ( .A(n18929), .B(n18930), .Z(n18927) );
  AND U19192 ( .A(a[3]), .B(b[19]), .Z(n18926) );
  XOR U19193 ( .A(n18931), .B(n18799), .Z(n18801) );
  XOR U19194 ( .A(n18932), .B(n18933), .Z(n18799) );
  AND U19195 ( .A(n18934), .B(n18935), .Z(n18932) );
  AND U19196 ( .A(a[4]), .B(b[18]), .Z(n18931) );
  XOR U19197 ( .A(n18936), .B(n18804), .Z(n18806) );
  XOR U19198 ( .A(n18937), .B(n18938), .Z(n18804) );
  AND U19199 ( .A(n18939), .B(n18940), .Z(n18937) );
  AND U19200 ( .A(a[5]), .B(b[17]), .Z(n18936) );
  XOR U19201 ( .A(n18941), .B(n18809), .Z(n18811) );
  XOR U19202 ( .A(n18942), .B(n18943), .Z(n18809) );
  AND U19203 ( .A(n18944), .B(n18945), .Z(n18942) );
  AND U19204 ( .A(a[6]), .B(b[16]), .Z(n18941) );
  XOR U19205 ( .A(n18946), .B(n18814), .Z(n18816) );
  XOR U19206 ( .A(n18947), .B(n18948), .Z(n18814) );
  AND U19207 ( .A(n18949), .B(n18950), .Z(n18947) );
  AND U19208 ( .A(a[7]), .B(b[15]), .Z(n18946) );
  XOR U19209 ( .A(n18951), .B(n18819), .Z(n18821) );
  XOR U19210 ( .A(n18952), .B(n18953), .Z(n18819) );
  AND U19211 ( .A(n18954), .B(n18955), .Z(n18952) );
  AND U19212 ( .A(a[8]), .B(b[14]), .Z(n18951) );
  XOR U19213 ( .A(n18956), .B(n18824), .Z(n18826) );
  XOR U19214 ( .A(n18957), .B(n18958), .Z(n18824) );
  AND U19215 ( .A(n18959), .B(n18960), .Z(n18957) );
  AND U19216 ( .A(a[9]), .B(b[13]), .Z(n18956) );
  XOR U19217 ( .A(n18961), .B(n18829), .Z(n18831) );
  XOR U19218 ( .A(n18962), .B(n18963), .Z(n18829) );
  AND U19219 ( .A(n18964), .B(n18965), .Z(n18962) );
  AND U19220 ( .A(a[10]), .B(b[12]), .Z(n18961) );
  XOR U19221 ( .A(n18966), .B(n18834), .Z(n18836) );
  XOR U19222 ( .A(n18967), .B(n18968), .Z(n18834) );
  AND U19223 ( .A(n18969), .B(n18970), .Z(n18967) );
  AND U19224 ( .A(a[11]), .B(b[11]), .Z(n18966) );
  XOR U19225 ( .A(n18971), .B(n18839), .Z(n18841) );
  XOR U19226 ( .A(n18972), .B(n18973), .Z(n18839) );
  AND U19227 ( .A(n18974), .B(n18975), .Z(n18972) );
  AND U19228 ( .A(b[10]), .B(a[12]), .Z(n18971) );
  XOR U19229 ( .A(n18976), .B(n18844), .Z(n18846) );
  XOR U19230 ( .A(n18977), .B(n18978), .Z(n18844) );
  AND U19231 ( .A(n18979), .B(n18980), .Z(n18977) );
  AND U19232 ( .A(a[13]), .B(b[9]), .Z(n18976) );
  XOR U19233 ( .A(n18981), .B(n18849), .Z(n18851) );
  XOR U19234 ( .A(n18982), .B(n18983), .Z(n18849) );
  AND U19235 ( .A(n18984), .B(n18985), .Z(n18982) );
  AND U19236 ( .A(b[8]), .B(a[14]), .Z(n18981) );
  XOR U19237 ( .A(n18986), .B(n18854), .Z(n18856) );
  XOR U19238 ( .A(n18987), .B(n18988), .Z(n18854) );
  AND U19239 ( .A(n18989), .B(n18990), .Z(n18987) );
  AND U19240 ( .A(a[15]), .B(b[7]), .Z(n18986) );
  XOR U19241 ( .A(n18991), .B(n18859), .Z(n18861) );
  XOR U19242 ( .A(n18992), .B(n18993), .Z(n18859) );
  AND U19243 ( .A(n18994), .B(n18995), .Z(n18992) );
  AND U19244 ( .A(b[6]), .B(a[16]), .Z(n18991) );
  XOR U19245 ( .A(n18996), .B(n18864), .Z(n18866) );
  XOR U19246 ( .A(n18997), .B(n18998), .Z(n18864) );
  AND U19247 ( .A(n18999), .B(n19000), .Z(n18997) );
  AND U19248 ( .A(a[17]), .B(b[5]), .Z(n18996) );
  XOR U19249 ( .A(n19001), .B(n18869), .Z(n18871) );
  XOR U19250 ( .A(n19002), .B(n19003), .Z(n18869) );
  AND U19251 ( .A(n19004), .B(n19005), .Z(n19002) );
  AND U19252 ( .A(b[4]), .B(a[18]), .Z(n19001) );
  XNOR U19253 ( .A(n19006), .B(n19007), .Z(n18883) );
  NANDN U19254 ( .A(n19008), .B(n19009), .Z(n19007) );
  XOR U19255 ( .A(n19010), .B(n18874), .Z(n18876) );
  XNOR U19256 ( .A(n19011), .B(n19012), .Z(n18874) );
  AND U19257 ( .A(n19013), .B(n19014), .Z(n19011) );
  AND U19258 ( .A(a[19]), .B(b[3]), .Z(n19010) );
  XOR U19259 ( .A(n18890), .B(n18889), .Z(c[117]) );
  XOR U19260 ( .A(sreg[149]), .B(n18888), .Z(n18889) );
  XOR U19261 ( .A(n18895), .B(n19015), .Z(n18890) );
  XNOR U19262 ( .A(n18894), .B(n18888), .Z(n19015) );
  XOR U19263 ( .A(n19016), .B(n19017), .Z(n18888) );
  NOR U19264 ( .A(n19018), .B(n19019), .Z(n19016) );
  NAND U19265 ( .A(a[21]), .B(b[0]), .Z(n18894) );
  XNOR U19266 ( .A(n19008), .B(n19009), .Z(n18895) );
  XOR U19267 ( .A(n19006), .B(n19020), .Z(n19009) );
  NAND U19268 ( .A(b[1]), .B(a[20]), .Z(n19020) );
  XOR U19269 ( .A(n19014), .B(n19021), .Z(n19008) );
  XOR U19270 ( .A(n19006), .B(n19013), .Z(n19021) );
  XNOR U19271 ( .A(n19022), .B(n19012), .Z(n19013) );
  AND U19272 ( .A(b[2]), .B(a[19]), .Z(n19022) );
  NANDN U19273 ( .A(n19023), .B(n19024), .Z(n19006) );
  XOR U19274 ( .A(n19012), .B(n19004), .Z(n19025) );
  XNOR U19275 ( .A(n19003), .B(n18999), .Z(n19026) );
  XNOR U19276 ( .A(n18998), .B(n18994), .Z(n19027) );
  XNOR U19277 ( .A(n18993), .B(n18989), .Z(n19028) );
  XNOR U19278 ( .A(n18988), .B(n18984), .Z(n19029) );
  XNOR U19279 ( .A(n18983), .B(n18979), .Z(n19030) );
  XNOR U19280 ( .A(n18978), .B(n18974), .Z(n19031) );
  XNOR U19281 ( .A(n18973), .B(n18969), .Z(n19032) );
  XNOR U19282 ( .A(n18968), .B(n18964), .Z(n19033) );
  XNOR U19283 ( .A(n18963), .B(n18959), .Z(n19034) );
  XNOR U19284 ( .A(n18958), .B(n18954), .Z(n19035) );
  XNOR U19285 ( .A(n18953), .B(n18949), .Z(n19036) );
  XNOR U19286 ( .A(n18948), .B(n18944), .Z(n19037) );
  XNOR U19287 ( .A(n18943), .B(n18939), .Z(n19038) );
  XNOR U19288 ( .A(n18938), .B(n18934), .Z(n19039) );
  XNOR U19289 ( .A(n18933), .B(n18929), .Z(n19040) );
  XNOR U19290 ( .A(n18928), .B(n18924), .Z(n19041) );
  XNOR U19291 ( .A(n18923), .B(n18919), .Z(n19042) );
  XOR U19292 ( .A(n19043), .B(n18918), .Z(n18919) );
  AND U19293 ( .A(a[0]), .B(b[21]), .Z(n19043) );
  XOR U19294 ( .A(n19044), .B(n18918), .Z(n18920) );
  XNOR U19295 ( .A(n19045), .B(n19046), .Z(n18918) );
  AND U19296 ( .A(n19047), .B(n19048), .Z(n19045) );
  AND U19297 ( .A(a[1]), .B(b[20]), .Z(n19044) );
  XOR U19298 ( .A(n19049), .B(n18923), .Z(n18925) );
  XOR U19299 ( .A(n19050), .B(n19051), .Z(n18923) );
  AND U19300 ( .A(n19052), .B(n19053), .Z(n19050) );
  AND U19301 ( .A(a[2]), .B(b[19]), .Z(n19049) );
  XOR U19302 ( .A(n19054), .B(n18928), .Z(n18930) );
  XOR U19303 ( .A(n19055), .B(n19056), .Z(n18928) );
  AND U19304 ( .A(n19057), .B(n19058), .Z(n19055) );
  AND U19305 ( .A(a[3]), .B(b[18]), .Z(n19054) );
  XOR U19306 ( .A(n19059), .B(n18933), .Z(n18935) );
  XOR U19307 ( .A(n19060), .B(n19061), .Z(n18933) );
  AND U19308 ( .A(n19062), .B(n19063), .Z(n19060) );
  AND U19309 ( .A(a[4]), .B(b[17]), .Z(n19059) );
  XOR U19310 ( .A(n19064), .B(n18938), .Z(n18940) );
  XOR U19311 ( .A(n19065), .B(n19066), .Z(n18938) );
  AND U19312 ( .A(n19067), .B(n19068), .Z(n19065) );
  AND U19313 ( .A(a[5]), .B(b[16]), .Z(n19064) );
  XOR U19314 ( .A(n19069), .B(n18943), .Z(n18945) );
  XOR U19315 ( .A(n19070), .B(n19071), .Z(n18943) );
  AND U19316 ( .A(n19072), .B(n19073), .Z(n19070) );
  AND U19317 ( .A(a[6]), .B(b[15]), .Z(n19069) );
  XOR U19318 ( .A(n19074), .B(n18948), .Z(n18950) );
  XOR U19319 ( .A(n19075), .B(n19076), .Z(n18948) );
  AND U19320 ( .A(n19077), .B(n19078), .Z(n19075) );
  AND U19321 ( .A(a[7]), .B(b[14]), .Z(n19074) );
  XOR U19322 ( .A(n19079), .B(n18953), .Z(n18955) );
  XOR U19323 ( .A(n19080), .B(n19081), .Z(n18953) );
  AND U19324 ( .A(n19082), .B(n19083), .Z(n19080) );
  AND U19325 ( .A(a[8]), .B(b[13]), .Z(n19079) );
  XOR U19326 ( .A(n19084), .B(n18958), .Z(n18960) );
  XOR U19327 ( .A(n19085), .B(n19086), .Z(n18958) );
  AND U19328 ( .A(n19087), .B(n19088), .Z(n19085) );
  AND U19329 ( .A(a[9]), .B(b[12]), .Z(n19084) );
  XOR U19330 ( .A(n19089), .B(n18963), .Z(n18965) );
  XOR U19331 ( .A(n19090), .B(n19091), .Z(n18963) );
  AND U19332 ( .A(n19092), .B(n19093), .Z(n19090) );
  AND U19333 ( .A(a[10]), .B(b[11]), .Z(n19089) );
  XOR U19334 ( .A(n19094), .B(n18968), .Z(n18970) );
  XOR U19335 ( .A(n19095), .B(n19096), .Z(n18968) );
  AND U19336 ( .A(n19097), .B(n19098), .Z(n19095) );
  AND U19337 ( .A(a[11]), .B(b[10]), .Z(n19094) );
  XOR U19338 ( .A(n19099), .B(n18973), .Z(n18975) );
  XOR U19339 ( .A(n19100), .B(n19101), .Z(n18973) );
  AND U19340 ( .A(n19102), .B(n19103), .Z(n19100) );
  AND U19341 ( .A(b[9]), .B(a[12]), .Z(n19099) );
  XOR U19342 ( .A(n19104), .B(n18978), .Z(n18980) );
  XOR U19343 ( .A(n19105), .B(n19106), .Z(n18978) );
  AND U19344 ( .A(n19107), .B(n19108), .Z(n19105) );
  AND U19345 ( .A(a[13]), .B(b[8]), .Z(n19104) );
  XOR U19346 ( .A(n19109), .B(n18983), .Z(n18985) );
  XOR U19347 ( .A(n19110), .B(n19111), .Z(n18983) );
  AND U19348 ( .A(n19112), .B(n19113), .Z(n19110) );
  AND U19349 ( .A(b[7]), .B(a[14]), .Z(n19109) );
  XOR U19350 ( .A(n19114), .B(n18988), .Z(n18990) );
  XOR U19351 ( .A(n19115), .B(n19116), .Z(n18988) );
  AND U19352 ( .A(n19117), .B(n19118), .Z(n19115) );
  AND U19353 ( .A(a[15]), .B(b[6]), .Z(n19114) );
  XOR U19354 ( .A(n19119), .B(n18993), .Z(n18995) );
  XOR U19355 ( .A(n19120), .B(n19121), .Z(n18993) );
  AND U19356 ( .A(n19122), .B(n19123), .Z(n19120) );
  AND U19357 ( .A(b[5]), .B(a[16]), .Z(n19119) );
  XOR U19358 ( .A(n19124), .B(n18998), .Z(n19000) );
  XOR U19359 ( .A(n19125), .B(n19126), .Z(n18998) );
  AND U19360 ( .A(n19127), .B(n19128), .Z(n19125) );
  AND U19361 ( .A(a[17]), .B(b[4]), .Z(n19124) );
  XNOR U19362 ( .A(n19129), .B(n19130), .Z(n19012) );
  NANDN U19363 ( .A(n19131), .B(n19132), .Z(n19130) );
  XOR U19364 ( .A(n19133), .B(n19003), .Z(n19005) );
  XNOR U19365 ( .A(n19134), .B(n19135), .Z(n19003) );
  AND U19366 ( .A(n19136), .B(n19137), .Z(n19134) );
  AND U19367 ( .A(b[3]), .B(a[18]), .Z(n19133) );
  XOR U19368 ( .A(n19019), .B(n19018), .Z(c[116]) );
  XOR U19369 ( .A(sreg[148]), .B(n19017), .Z(n19018) );
  XOR U19370 ( .A(n19024), .B(n19138), .Z(n19019) );
  XNOR U19371 ( .A(n19023), .B(n19017), .Z(n19138) );
  XOR U19372 ( .A(n19139), .B(n19140), .Z(n19017) );
  NOR U19373 ( .A(n19141), .B(n19142), .Z(n19139) );
  NAND U19374 ( .A(a[20]), .B(b[0]), .Z(n19023) );
  XNOR U19375 ( .A(n19131), .B(n19132), .Z(n19024) );
  XOR U19376 ( .A(n19129), .B(n19143), .Z(n19132) );
  NAND U19377 ( .A(a[19]), .B(b[1]), .Z(n19143) );
  XOR U19378 ( .A(n19137), .B(n19144), .Z(n19131) );
  XOR U19379 ( .A(n19129), .B(n19136), .Z(n19144) );
  XNOR U19380 ( .A(n19145), .B(n19135), .Z(n19136) );
  AND U19381 ( .A(b[2]), .B(a[18]), .Z(n19145) );
  NANDN U19382 ( .A(n19146), .B(n19147), .Z(n19129) );
  XOR U19383 ( .A(n19135), .B(n19127), .Z(n19148) );
  XNOR U19384 ( .A(n19126), .B(n19122), .Z(n19149) );
  XNOR U19385 ( .A(n19121), .B(n19117), .Z(n19150) );
  XNOR U19386 ( .A(n19116), .B(n19112), .Z(n19151) );
  XNOR U19387 ( .A(n19111), .B(n19107), .Z(n19152) );
  XNOR U19388 ( .A(n19106), .B(n19102), .Z(n19153) );
  XNOR U19389 ( .A(n19101), .B(n19097), .Z(n19154) );
  XNOR U19390 ( .A(n19096), .B(n19092), .Z(n19155) );
  XNOR U19391 ( .A(n19091), .B(n19087), .Z(n19156) );
  XNOR U19392 ( .A(n19086), .B(n19082), .Z(n19157) );
  XNOR U19393 ( .A(n19081), .B(n19077), .Z(n19158) );
  XNOR U19394 ( .A(n19076), .B(n19072), .Z(n19159) );
  XNOR U19395 ( .A(n19071), .B(n19067), .Z(n19160) );
  XNOR U19396 ( .A(n19066), .B(n19062), .Z(n19161) );
  XNOR U19397 ( .A(n19061), .B(n19057), .Z(n19162) );
  XNOR U19398 ( .A(n19056), .B(n19052), .Z(n19163) );
  XNOR U19399 ( .A(n19051), .B(n19047), .Z(n19164) );
  XNOR U19400 ( .A(n19165), .B(n19046), .Z(n19047) );
  AND U19401 ( .A(a[0]), .B(b[20]), .Z(n19165) );
  XNOR U19402 ( .A(n19166), .B(n19046), .Z(n19048) );
  XNOR U19403 ( .A(n19167), .B(n19168), .Z(n19046) );
  AND U19404 ( .A(n19169), .B(n19170), .Z(n19167) );
  AND U19405 ( .A(a[1]), .B(b[19]), .Z(n19166) );
  XOR U19406 ( .A(n19171), .B(n19051), .Z(n19053) );
  XOR U19407 ( .A(n19172), .B(n19173), .Z(n19051) );
  AND U19408 ( .A(n19174), .B(n19175), .Z(n19172) );
  AND U19409 ( .A(a[2]), .B(b[18]), .Z(n19171) );
  XOR U19410 ( .A(n19176), .B(n19056), .Z(n19058) );
  XOR U19411 ( .A(n19177), .B(n19178), .Z(n19056) );
  AND U19412 ( .A(n19179), .B(n19180), .Z(n19177) );
  AND U19413 ( .A(a[3]), .B(b[17]), .Z(n19176) );
  XOR U19414 ( .A(n19181), .B(n19061), .Z(n19063) );
  XOR U19415 ( .A(n19182), .B(n19183), .Z(n19061) );
  AND U19416 ( .A(n19184), .B(n19185), .Z(n19182) );
  AND U19417 ( .A(a[4]), .B(b[16]), .Z(n19181) );
  XOR U19418 ( .A(n19186), .B(n19066), .Z(n19068) );
  XOR U19419 ( .A(n19187), .B(n19188), .Z(n19066) );
  AND U19420 ( .A(n19189), .B(n19190), .Z(n19187) );
  AND U19421 ( .A(a[5]), .B(b[15]), .Z(n19186) );
  XOR U19422 ( .A(n19191), .B(n19071), .Z(n19073) );
  XOR U19423 ( .A(n19192), .B(n19193), .Z(n19071) );
  AND U19424 ( .A(n19194), .B(n19195), .Z(n19192) );
  AND U19425 ( .A(a[6]), .B(b[14]), .Z(n19191) );
  XOR U19426 ( .A(n19196), .B(n19076), .Z(n19078) );
  XOR U19427 ( .A(n19197), .B(n19198), .Z(n19076) );
  AND U19428 ( .A(n19199), .B(n19200), .Z(n19197) );
  AND U19429 ( .A(a[7]), .B(b[13]), .Z(n19196) );
  XOR U19430 ( .A(n19201), .B(n19081), .Z(n19083) );
  XOR U19431 ( .A(n19202), .B(n19203), .Z(n19081) );
  AND U19432 ( .A(n19204), .B(n19205), .Z(n19202) );
  AND U19433 ( .A(a[8]), .B(b[12]), .Z(n19201) );
  XOR U19434 ( .A(n19206), .B(n19086), .Z(n19088) );
  XOR U19435 ( .A(n19207), .B(n19208), .Z(n19086) );
  AND U19436 ( .A(n19209), .B(n19210), .Z(n19207) );
  AND U19437 ( .A(a[9]), .B(b[11]), .Z(n19206) );
  XOR U19438 ( .A(n19211), .B(n19091), .Z(n19093) );
  XOR U19439 ( .A(n19212), .B(n19213), .Z(n19091) );
  AND U19440 ( .A(n19214), .B(n19215), .Z(n19212) );
  AND U19441 ( .A(b[10]), .B(a[10]), .Z(n19211) );
  XOR U19442 ( .A(n19216), .B(n19096), .Z(n19098) );
  XOR U19443 ( .A(n19217), .B(n19218), .Z(n19096) );
  AND U19444 ( .A(n19219), .B(n19220), .Z(n19217) );
  AND U19445 ( .A(a[11]), .B(b[9]), .Z(n19216) );
  XOR U19446 ( .A(n19221), .B(n19101), .Z(n19103) );
  XOR U19447 ( .A(n19222), .B(n19223), .Z(n19101) );
  AND U19448 ( .A(n19224), .B(n19225), .Z(n19222) );
  AND U19449 ( .A(b[8]), .B(a[12]), .Z(n19221) );
  XOR U19450 ( .A(n19226), .B(n19106), .Z(n19108) );
  XOR U19451 ( .A(n19227), .B(n19228), .Z(n19106) );
  AND U19452 ( .A(n19229), .B(n19230), .Z(n19227) );
  AND U19453 ( .A(a[13]), .B(b[7]), .Z(n19226) );
  XOR U19454 ( .A(n19231), .B(n19111), .Z(n19113) );
  XOR U19455 ( .A(n19232), .B(n19233), .Z(n19111) );
  AND U19456 ( .A(n19234), .B(n19235), .Z(n19232) );
  AND U19457 ( .A(b[6]), .B(a[14]), .Z(n19231) );
  XOR U19458 ( .A(n19236), .B(n19116), .Z(n19118) );
  XOR U19459 ( .A(n19237), .B(n19238), .Z(n19116) );
  AND U19460 ( .A(n19239), .B(n19240), .Z(n19237) );
  AND U19461 ( .A(a[15]), .B(b[5]), .Z(n19236) );
  XOR U19462 ( .A(n19241), .B(n19121), .Z(n19123) );
  XOR U19463 ( .A(n19242), .B(n19243), .Z(n19121) );
  AND U19464 ( .A(n19244), .B(n19245), .Z(n19242) );
  AND U19465 ( .A(b[4]), .B(a[16]), .Z(n19241) );
  XNOR U19466 ( .A(n19246), .B(n19247), .Z(n19135) );
  NANDN U19467 ( .A(n19248), .B(n19249), .Z(n19247) );
  XOR U19468 ( .A(n19250), .B(n19126), .Z(n19128) );
  XNOR U19469 ( .A(n19251), .B(n19252), .Z(n19126) );
  AND U19470 ( .A(n19253), .B(n19254), .Z(n19251) );
  AND U19471 ( .A(a[17]), .B(b[3]), .Z(n19250) );
  XOR U19472 ( .A(n19142), .B(n19141), .Z(c[115]) );
  XOR U19473 ( .A(sreg[147]), .B(n19140), .Z(n19141) );
  XOR U19474 ( .A(n19147), .B(n19255), .Z(n19142) );
  XNOR U19475 ( .A(n19146), .B(n19140), .Z(n19255) );
  XOR U19476 ( .A(n19256), .B(n19257), .Z(n19140) );
  NOR U19477 ( .A(n19258), .B(n19259), .Z(n19256) );
  NAND U19478 ( .A(a[19]), .B(b[0]), .Z(n19146) );
  XNOR U19479 ( .A(n19248), .B(n19249), .Z(n19147) );
  XOR U19480 ( .A(n19246), .B(n19260), .Z(n19249) );
  NAND U19481 ( .A(b[1]), .B(a[18]), .Z(n19260) );
  XOR U19482 ( .A(n19254), .B(n19261), .Z(n19248) );
  XOR U19483 ( .A(n19246), .B(n19253), .Z(n19261) );
  XNOR U19484 ( .A(n19262), .B(n19252), .Z(n19253) );
  AND U19485 ( .A(b[2]), .B(a[17]), .Z(n19262) );
  NANDN U19486 ( .A(n19263), .B(n19264), .Z(n19246) );
  XOR U19487 ( .A(n19252), .B(n19244), .Z(n19265) );
  XNOR U19488 ( .A(n19243), .B(n19239), .Z(n19266) );
  XNOR U19489 ( .A(n19238), .B(n19234), .Z(n19267) );
  XNOR U19490 ( .A(n19233), .B(n19229), .Z(n19268) );
  XNOR U19491 ( .A(n19228), .B(n19224), .Z(n19269) );
  XNOR U19492 ( .A(n19223), .B(n19219), .Z(n19270) );
  XNOR U19493 ( .A(n19218), .B(n19214), .Z(n19271) );
  XNOR U19494 ( .A(n19213), .B(n19209), .Z(n19272) );
  XNOR U19495 ( .A(n19208), .B(n19204), .Z(n19273) );
  XNOR U19496 ( .A(n19203), .B(n19199), .Z(n19274) );
  XNOR U19497 ( .A(n19198), .B(n19194), .Z(n19275) );
  XNOR U19498 ( .A(n19193), .B(n19189), .Z(n19276) );
  XNOR U19499 ( .A(n19188), .B(n19184), .Z(n19277) );
  XNOR U19500 ( .A(n19183), .B(n19179), .Z(n19278) );
  XNOR U19501 ( .A(n19178), .B(n19174), .Z(n19279) );
  XNOR U19502 ( .A(n19173), .B(n19169), .Z(n19280) );
  XOR U19503 ( .A(n19281), .B(n19168), .Z(n19169) );
  AND U19504 ( .A(a[0]), .B(b[19]), .Z(n19281) );
  XOR U19505 ( .A(n19282), .B(n19168), .Z(n19170) );
  XNOR U19506 ( .A(n19283), .B(n19284), .Z(n19168) );
  AND U19507 ( .A(n19285), .B(n19286), .Z(n19283) );
  AND U19508 ( .A(a[1]), .B(b[18]), .Z(n19282) );
  XOR U19509 ( .A(n19287), .B(n19173), .Z(n19175) );
  XOR U19510 ( .A(n19288), .B(n19289), .Z(n19173) );
  AND U19511 ( .A(n19290), .B(n19291), .Z(n19288) );
  AND U19512 ( .A(a[2]), .B(b[17]), .Z(n19287) );
  XOR U19513 ( .A(n19292), .B(n19178), .Z(n19180) );
  XOR U19514 ( .A(n19293), .B(n19294), .Z(n19178) );
  AND U19515 ( .A(n19295), .B(n19296), .Z(n19293) );
  AND U19516 ( .A(a[3]), .B(b[16]), .Z(n19292) );
  XOR U19517 ( .A(n19297), .B(n19183), .Z(n19185) );
  XOR U19518 ( .A(n19298), .B(n19299), .Z(n19183) );
  AND U19519 ( .A(n19300), .B(n19301), .Z(n19298) );
  AND U19520 ( .A(a[4]), .B(b[15]), .Z(n19297) );
  XOR U19521 ( .A(n19302), .B(n19188), .Z(n19190) );
  XOR U19522 ( .A(n19303), .B(n19304), .Z(n19188) );
  AND U19523 ( .A(n19305), .B(n19306), .Z(n19303) );
  AND U19524 ( .A(a[5]), .B(b[14]), .Z(n19302) );
  XOR U19525 ( .A(n19307), .B(n19193), .Z(n19195) );
  XOR U19526 ( .A(n19308), .B(n19309), .Z(n19193) );
  AND U19527 ( .A(n19310), .B(n19311), .Z(n19308) );
  AND U19528 ( .A(a[6]), .B(b[13]), .Z(n19307) );
  XOR U19529 ( .A(n19312), .B(n19198), .Z(n19200) );
  XOR U19530 ( .A(n19313), .B(n19314), .Z(n19198) );
  AND U19531 ( .A(n19315), .B(n19316), .Z(n19313) );
  AND U19532 ( .A(a[7]), .B(b[12]), .Z(n19312) );
  XOR U19533 ( .A(n19317), .B(n19203), .Z(n19205) );
  XOR U19534 ( .A(n19318), .B(n19319), .Z(n19203) );
  AND U19535 ( .A(n19320), .B(n19321), .Z(n19318) );
  AND U19536 ( .A(a[8]), .B(b[11]), .Z(n19317) );
  XOR U19537 ( .A(n19322), .B(n19208), .Z(n19210) );
  XOR U19538 ( .A(n19323), .B(n19324), .Z(n19208) );
  AND U19539 ( .A(n19325), .B(n19326), .Z(n19323) );
  AND U19540 ( .A(a[9]), .B(b[10]), .Z(n19322) );
  XOR U19541 ( .A(n19327), .B(n19213), .Z(n19215) );
  XOR U19542 ( .A(n19328), .B(n19329), .Z(n19213) );
  AND U19543 ( .A(n19330), .B(n19331), .Z(n19328) );
  AND U19544 ( .A(b[9]), .B(a[10]), .Z(n19327) );
  XOR U19545 ( .A(n19332), .B(n19218), .Z(n19220) );
  XOR U19546 ( .A(n19333), .B(n19334), .Z(n19218) );
  AND U19547 ( .A(n19335), .B(n19336), .Z(n19333) );
  AND U19548 ( .A(a[11]), .B(b[8]), .Z(n19332) );
  XOR U19549 ( .A(n19337), .B(n19223), .Z(n19225) );
  XOR U19550 ( .A(n19338), .B(n19339), .Z(n19223) );
  AND U19551 ( .A(n19340), .B(n19341), .Z(n19338) );
  AND U19552 ( .A(b[7]), .B(a[12]), .Z(n19337) );
  XOR U19553 ( .A(n19342), .B(n19228), .Z(n19230) );
  XOR U19554 ( .A(n19343), .B(n19344), .Z(n19228) );
  AND U19555 ( .A(n19345), .B(n19346), .Z(n19343) );
  AND U19556 ( .A(a[13]), .B(b[6]), .Z(n19342) );
  XOR U19557 ( .A(n19347), .B(n19233), .Z(n19235) );
  XOR U19558 ( .A(n19348), .B(n19349), .Z(n19233) );
  AND U19559 ( .A(n19350), .B(n19351), .Z(n19348) );
  AND U19560 ( .A(b[5]), .B(a[14]), .Z(n19347) );
  XOR U19561 ( .A(n19352), .B(n19238), .Z(n19240) );
  XOR U19562 ( .A(n19353), .B(n19354), .Z(n19238) );
  AND U19563 ( .A(n19355), .B(n19356), .Z(n19353) );
  AND U19564 ( .A(a[15]), .B(b[4]), .Z(n19352) );
  XNOR U19565 ( .A(n19357), .B(n19358), .Z(n19252) );
  NANDN U19566 ( .A(n19359), .B(n19360), .Z(n19358) );
  XOR U19567 ( .A(n19361), .B(n19243), .Z(n19245) );
  XNOR U19568 ( .A(n19362), .B(n19363), .Z(n19243) );
  AND U19569 ( .A(n19364), .B(n19365), .Z(n19362) );
  AND U19570 ( .A(b[3]), .B(a[16]), .Z(n19361) );
  XOR U19571 ( .A(n19259), .B(n19258), .Z(c[114]) );
  XOR U19572 ( .A(sreg[146]), .B(n19257), .Z(n19258) );
  XOR U19573 ( .A(n19264), .B(n19366), .Z(n19259) );
  XNOR U19574 ( .A(n19263), .B(n19257), .Z(n19366) );
  XOR U19575 ( .A(n19367), .B(n19368), .Z(n19257) );
  NOR U19576 ( .A(n19369), .B(n19370), .Z(n19367) );
  NAND U19577 ( .A(a[18]), .B(b[0]), .Z(n19263) );
  XNOR U19578 ( .A(n19359), .B(n19360), .Z(n19264) );
  XOR U19579 ( .A(n19357), .B(n19371), .Z(n19360) );
  NAND U19580 ( .A(a[17]), .B(b[1]), .Z(n19371) );
  XOR U19581 ( .A(n19365), .B(n19372), .Z(n19359) );
  XOR U19582 ( .A(n19357), .B(n19364), .Z(n19372) );
  XNOR U19583 ( .A(n19373), .B(n19363), .Z(n19364) );
  AND U19584 ( .A(b[2]), .B(a[16]), .Z(n19373) );
  NANDN U19585 ( .A(n19374), .B(n19375), .Z(n19357) );
  XOR U19586 ( .A(n19363), .B(n19355), .Z(n19376) );
  XNOR U19587 ( .A(n19354), .B(n19350), .Z(n19377) );
  XNOR U19588 ( .A(n19349), .B(n19345), .Z(n19378) );
  XNOR U19589 ( .A(n19344), .B(n19340), .Z(n19379) );
  XNOR U19590 ( .A(n19339), .B(n19335), .Z(n19380) );
  XNOR U19591 ( .A(n19334), .B(n19330), .Z(n19381) );
  XNOR U19592 ( .A(n19329), .B(n19325), .Z(n19382) );
  XNOR U19593 ( .A(n19324), .B(n19320), .Z(n19383) );
  XNOR U19594 ( .A(n19319), .B(n19315), .Z(n19384) );
  XNOR U19595 ( .A(n19314), .B(n19310), .Z(n19385) );
  XNOR U19596 ( .A(n19309), .B(n19305), .Z(n19386) );
  XNOR U19597 ( .A(n19304), .B(n19300), .Z(n19387) );
  XNOR U19598 ( .A(n19299), .B(n19295), .Z(n19388) );
  XNOR U19599 ( .A(n19294), .B(n19290), .Z(n19389) );
  XNOR U19600 ( .A(n19289), .B(n19285), .Z(n19390) );
  XNOR U19601 ( .A(n19391), .B(n19284), .Z(n19285) );
  AND U19602 ( .A(a[0]), .B(b[18]), .Z(n19391) );
  XNOR U19603 ( .A(n19392), .B(n19284), .Z(n19286) );
  XNOR U19604 ( .A(n19393), .B(n19394), .Z(n19284) );
  AND U19605 ( .A(n19395), .B(n19396), .Z(n19393) );
  AND U19606 ( .A(a[1]), .B(b[17]), .Z(n19392) );
  XOR U19607 ( .A(n19397), .B(n19289), .Z(n19291) );
  XOR U19608 ( .A(n19398), .B(n19399), .Z(n19289) );
  AND U19609 ( .A(n19400), .B(n19401), .Z(n19398) );
  AND U19610 ( .A(a[2]), .B(b[16]), .Z(n19397) );
  XOR U19611 ( .A(n19402), .B(n19294), .Z(n19296) );
  XOR U19612 ( .A(n19403), .B(n19404), .Z(n19294) );
  AND U19613 ( .A(n19405), .B(n19406), .Z(n19403) );
  AND U19614 ( .A(a[3]), .B(b[15]), .Z(n19402) );
  XOR U19615 ( .A(n19407), .B(n19299), .Z(n19301) );
  XOR U19616 ( .A(n19408), .B(n19409), .Z(n19299) );
  AND U19617 ( .A(n19410), .B(n19411), .Z(n19408) );
  AND U19618 ( .A(a[4]), .B(b[14]), .Z(n19407) );
  XOR U19619 ( .A(n19412), .B(n19304), .Z(n19306) );
  XOR U19620 ( .A(n19413), .B(n19414), .Z(n19304) );
  AND U19621 ( .A(n19415), .B(n19416), .Z(n19413) );
  AND U19622 ( .A(a[5]), .B(b[13]), .Z(n19412) );
  XOR U19623 ( .A(n19417), .B(n19309), .Z(n19311) );
  XOR U19624 ( .A(n19418), .B(n19419), .Z(n19309) );
  AND U19625 ( .A(n19420), .B(n19421), .Z(n19418) );
  AND U19626 ( .A(a[6]), .B(b[12]), .Z(n19417) );
  XOR U19627 ( .A(n19422), .B(n19314), .Z(n19316) );
  XOR U19628 ( .A(n19423), .B(n19424), .Z(n19314) );
  AND U19629 ( .A(n19425), .B(n19426), .Z(n19423) );
  AND U19630 ( .A(a[7]), .B(b[11]), .Z(n19422) );
  XOR U19631 ( .A(n19427), .B(n19319), .Z(n19321) );
  XOR U19632 ( .A(n19428), .B(n19429), .Z(n19319) );
  AND U19633 ( .A(n19430), .B(n19431), .Z(n19428) );
  AND U19634 ( .A(a[8]), .B(b[10]), .Z(n19427) );
  XOR U19635 ( .A(n19432), .B(n19324), .Z(n19326) );
  XOR U19636 ( .A(n19433), .B(n19434), .Z(n19324) );
  AND U19637 ( .A(n19435), .B(n19436), .Z(n19433) );
  AND U19638 ( .A(a[9]), .B(b[9]), .Z(n19432) );
  XOR U19639 ( .A(n19437), .B(n19329), .Z(n19331) );
  XOR U19640 ( .A(n19438), .B(n19439), .Z(n19329) );
  AND U19641 ( .A(n19440), .B(n19441), .Z(n19438) );
  AND U19642 ( .A(b[8]), .B(a[10]), .Z(n19437) );
  XOR U19643 ( .A(n19442), .B(n19334), .Z(n19336) );
  XOR U19644 ( .A(n19443), .B(n19444), .Z(n19334) );
  AND U19645 ( .A(n19445), .B(n19446), .Z(n19443) );
  AND U19646 ( .A(a[11]), .B(b[7]), .Z(n19442) );
  XOR U19647 ( .A(n19447), .B(n19339), .Z(n19341) );
  XOR U19648 ( .A(n19448), .B(n19449), .Z(n19339) );
  AND U19649 ( .A(n19450), .B(n19451), .Z(n19448) );
  AND U19650 ( .A(b[6]), .B(a[12]), .Z(n19447) );
  XOR U19651 ( .A(n19452), .B(n19344), .Z(n19346) );
  XOR U19652 ( .A(n19453), .B(n19454), .Z(n19344) );
  AND U19653 ( .A(n19455), .B(n19456), .Z(n19453) );
  AND U19654 ( .A(a[13]), .B(b[5]), .Z(n19452) );
  XOR U19655 ( .A(n19457), .B(n19349), .Z(n19351) );
  XOR U19656 ( .A(n19458), .B(n19459), .Z(n19349) );
  AND U19657 ( .A(n19460), .B(n19461), .Z(n19458) );
  AND U19658 ( .A(b[4]), .B(a[14]), .Z(n19457) );
  XNOR U19659 ( .A(n19462), .B(n19463), .Z(n19363) );
  NANDN U19660 ( .A(n19464), .B(n19465), .Z(n19463) );
  XOR U19661 ( .A(n19466), .B(n19354), .Z(n19356) );
  XNOR U19662 ( .A(n19467), .B(n19468), .Z(n19354) );
  AND U19663 ( .A(n19469), .B(n19470), .Z(n19467) );
  AND U19664 ( .A(a[15]), .B(b[3]), .Z(n19466) );
  XOR U19665 ( .A(n19370), .B(n19369), .Z(c[113]) );
  XOR U19666 ( .A(sreg[145]), .B(n19368), .Z(n19369) );
  XOR U19667 ( .A(n19375), .B(n19471), .Z(n19370) );
  XNOR U19668 ( .A(n19374), .B(n19368), .Z(n19471) );
  XOR U19669 ( .A(n19472), .B(n19473), .Z(n19368) );
  NOR U19670 ( .A(n19474), .B(n19475), .Z(n19472) );
  NAND U19671 ( .A(a[17]), .B(b[0]), .Z(n19374) );
  XNOR U19672 ( .A(n19464), .B(n19465), .Z(n19375) );
  XOR U19673 ( .A(n19462), .B(n19476), .Z(n19465) );
  NAND U19674 ( .A(b[1]), .B(a[16]), .Z(n19476) );
  XOR U19675 ( .A(n19470), .B(n19477), .Z(n19464) );
  XOR U19676 ( .A(n19462), .B(n19469), .Z(n19477) );
  XNOR U19677 ( .A(n19478), .B(n19468), .Z(n19469) );
  AND U19678 ( .A(b[2]), .B(a[15]), .Z(n19478) );
  NANDN U19679 ( .A(n19479), .B(n19480), .Z(n19462) );
  XOR U19680 ( .A(n19468), .B(n19460), .Z(n19481) );
  XNOR U19681 ( .A(n19459), .B(n19455), .Z(n19482) );
  XNOR U19682 ( .A(n19454), .B(n19450), .Z(n19483) );
  XNOR U19683 ( .A(n19449), .B(n19445), .Z(n19484) );
  XNOR U19684 ( .A(n19444), .B(n19440), .Z(n19485) );
  XNOR U19685 ( .A(n19439), .B(n19435), .Z(n19486) );
  XNOR U19686 ( .A(n19434), .B(n19430), .Z(n19487) );
  XNOR U19687 ( .A(n19429), .B(n19425), .Z(n19488) );
  XNOR U19688 ( .A(n19424), .B(n19420), .Z(n19489) );
  XNOR U19689 ( .A(n19419), .B(n19415), .Z(n19490) );
  XNOR U19690 ( .A(n19414), .B(n19410), .Z(n19491) );
  XNOR U19691 ( .A(n19409), .B(n19405), .Z(n19492) );
  XNOR U19692 ( .A(n19404), .B(n19400), .Z(n19493) );
  XNOR U19693 ( .A(n19399), .B(n19395), .Z(n19494) );
  XOR U19694 ( .A(n19495), .B(n19394), .Z(n19395) );
  AND U19695 ( .A(a[0]), .B(b[17]), .Z(n19495) );
  XOR U19696 ( .A(n19496), .B(n19394), .Z(n19396) );
  XNOR U19697 ( .A(n19497), .B(n19498), .Z(n19394) );
  AND U19698 ( .A(n19499), .B(n19500), .Z(n19497) );
  AND U19699 ( .A(a[1]), .B(b[16]), .Z(n19496) );
  XOR U19700 ( .A(n19501), .B(n19399), .Z(n19401) );
  XOR U19701 ( .A(n19502), .B(n19503), .Z(n19399) );
  AND U19702 ( .A(n19504), .B(n19505), .Z(n19502) );
  AND U19703 ( .A(a[2]), .B(b[15]), .Z(n19501) );
  XOR U19704 ( .A(n19506), .B(n19404), .Z(n19406) );
  XOR U19705 ( .A(n19507), .B(n19508), .Z(n19404) );
  AND U19706 ( .A(n19509), .B(n19510), .Z(n19507) );
  AND U19707 ( .A(a[3]), .B(b[14]), .Z(n19506) );
  XOR U19708 ( .A(n19511), .B(n19409), .Z(n19411) );
  XOR U19709 ( .A(n19512), .B(n19513), .Z(n19409) );
  AND U19710 ( .A(n19514), .B(n19515), .Z(n19512) );
  AND U19711 ( .A(a[4]), .B(b[13]), .Z(n19511) );
  XOR U19712 ( .A(n19516), .B(n19414), .Z(n19416) );
  XOR U19713 ( .A(n19517), .B(n19518), .Z(n19414) );
  AND U19714 ( .A(n19519), .B(n19520), .Z(n19517) );
  AND U19715 ( .A(a[5]), .B(b[12]), .Z(n19516) );
  XOR U19716 ( .A(n19521), .B(n19419), .Z(n19421) );
  XOR U19717 ( .A(n19522), .B(n19523), .Z(n19419) );
  AND U19718 ( .A(n19524), .B(n19525), .Z(n19522) );
  AND U19719 ( .A(a[6]), .B(b[11]), .Z(n19521) );
  XOR U19720 ( .A(n19526), .B(n19424), .Z(n19426) );
  XOR U19721 ( .A(n19527), .B(n19528), .Z(n19424) );
  AND U19722 ( .A(n19529), .B(n19530), .Z(n19527) );
  AND U19723 ( .A(a[7]), .B(b[10]), .Z(n19526) );
  XOR U19724 ( .A(n19531), .B(n19429), .Z(n19431) );
  XOR U19725 ( .A(n19532), .B(n19533), .Z(n19429) );
  AND U19726 ( .A(n19534), .B(n19535), .Z(n19532) );
  AND U19727 ( .A(a[8]), .B(b[9]), .Z(n19531) );
  XOR U19728 ( .A(n19536), .B(n19434), .Z(n19436) );
  XOR U19729 ( .A(n19537), .B(n19538), .Z(n19434) );
  AND U19730 ( .A(n19539), .B(n19540), .Z(n19537) );
  AND U19731 ( .A(a[9]), .B(b[8]), .Z(n19536) );
  XOR U19732 ( .A(n19541), .B(n19439), .Z(n19441) );
  XOR U19733 ( .A(n19542), .B(n19543), .Z(n19439) );
  AND U19734 ( .A(n19544), .B(n19545), .Z(n19542) );
  AND U19735 ( .A(b[7]), .B(a[10]), .Z(n19541) );
  XOR U19736 ( .A(n19546), .B(n19444), .Z(n19446) );
  XOR U19737 ( .A(n19547), .B(n19548), .Z(n19444) );
  AND U19738 ( .A(n19549), .B(n19550), .Z(n19547) );
  AND U19739 ( .A(a[11]), .B(b[6]), .Z(n19546) );
  XOR U19740 ( .A(n19551), .B(n19449), .Z(n19451) );
  XOR U19741 ( .A(n19552), .B(n19553), .Z(n19449) );
  AND U19742 ( .A(n19554), .B(n19555), .Z(n19552) );
  AND U19743 ( .A(b[5]), .B(a[12]), .Z(n19551) );
  XOR U19744 ( .A(n19556), .B(n19454), .Z(n19456) );
  XOR U19745 ( .A(n19557), .B(n19558), .Z(n19454) );
  AND U19746 ( .A(n19559), .B(n19560), .Z(n19557) );
  AND U19747 ( .A(a[13]), .B(b[4]), .Z(n19556) );
  XNOR U19748 ( .A(n19561), .B(n19562), .Z(n19468) );
  NANDN U19749 ( .A(n19563), .B(n19564), .Z(n19562) );
  XOR U19750 ( .A(n19565), .B(n19459), .Z(n19461) );
  XNOR U19751 ( .A(n19566), .B(n19567), .Z(n19459) );
  AND U19752 ( .A(n19568), .B(n19569), .Z(n19566) );
  AND U19753 ( .A(b[3]), .B(a[14]), .Z(n19565) );
  XOR U19754 ( .A(n19475), .B(n19474), .Z(c[112]) );
  XOR U19755 ( .A(sreg[144]), .B(n19473), .Z(n19474) );
  XOR U19756 ( .A(n19480), .B(n19570), .Z(n19475) );
  XNOR U19757 ( .A(n19479), .B(n19473), .Z(n19570) );
  XOR U19758 ( .A(n19571), .B(n19572), .Z(n19473) );
  NOR U19759 ( .A(n19573), .B(n19574), .Z(n19571) );
  NAND U19760 ( .A(a[16]), .B(b[0]), .Z(n19479) );
  XNOR U19761 ( .A(n19563), .B(n19564), .Z(n19480) );
  XOR U19762 ( .A(n19561), .B(n19575), .Z(n19564) );
  NAND U19763 ( .A(a[15]), .B(b[1]), .Z(n19575) );
  XOR U19764 ( .A(n19569), .B(n19576), .Z(n19563) );
  XOR U19765 ( .A(n19561), .B(n19568), .Z(n19576) );
  XNOR U19766 ( .A(n19577), .B(n19567), .Z(n19568) );
  AND U19767 ( .A(b[2]), .B(a[14]), .Z(n19577) );
  NANDN U19768 ( .A(n19578), .B(n19579), .Z(n19561) );
  XOR U19769 ( .A(n19567), .B(n19559), .Z(n19580) );
  XNOR U19770 ( .A(n19558), .B(n19554), .Z(n19581) );
  XNOR U19771 ( .A(n19553), .B(n19549), .Z(n19582) );
  XNOR U19772 ( .A(n19548), .B(n19544), .Z(n19583) );
  XNOR U19773 ( .A(n19543), .B(n19539), .Z(n19584) );
  XNOR U19774 ( .A(n19538), .B(n19534), .Z(n19585) );
  XNOR U19775 ( .A(n19533), .B(n19529), .Z(n19586) );
  XNOR U19776 ( .A(n19528), .B(n19524), .Z(n19587) );
  XNOR U19777 ( .A(n19523), .B(n19519), .Z(n19588) );
  XNOR U19778 ( .A(n19518), .B(n19514), .Z(n19589) );
  XNOR U19779 ( .A(n19513), .B(n19509), .Z(n19590) );
  XNOR U19780 ( .A(n19508), .B(n19504), .Z(n19591) );
  XNOR U19781 ( .A(n19503), .B(n19499), .Z(n19592) );
  XNOR U19782 ( .A(n19593), .B(n19498), .Z(n19499) );
  AND U19783 ( .A(a[0]), .B(b[16]), .Z(n19593) );
  XNOR U19784 ( .A(n19594), .B(n19498), .Z(n19500) );
  XNOR U19785 ( .A(n19595), .B(n19596), .Z(n19498) );
  AND U19786 ( .A(n19597), .B(n19598), .Z(n19595) );
  AND U19787 ( .A(a[1]), .B(b[15]), .Z(n19594) );
  XOR U19788 ( .A(n19599), .B(n19503), .Z(n19505) );
  XOR U19789 ( .A(n19600), .B(n19601), .Z(n19503) );
  AND U19790 ( .A(n19602), .B(n19603), .Z(n19600) );
  AND U19791 ( .A(a[2]), .B(b[14]), .Z(n19599) );
  XOR U19792 ( .A(n19604), .B(n19508), .Z(n19510) );
  XOR U19793 ( .A(n19605), .B(n19606), .Z(n19508) );
  AND U19794 ( .A(n19607), .B(n19608), .Z(n19605) );
  AND U19795 ( .A(a[3]), .B(b[13]), .Z(n19604) );
  XOR U19796 ( .A(n19609), .B(n19513), .Z(n19515) );
  XOR U19797 ( .A(n19610), .B(n19611), .Z(n19513) );
  AND U19798 ( .A(n19612), .B(n19613), .Z(n19610) );
  AND U19799 ( .A(a[4]), .B(b[12]), .Z(n19609) );
  XOR U19800 ( .A(n19614), .B(n19518), .Z(n19520) );
  XOR U19801 ( .A(n19615), .B(n19616), .Z(n19518) );
  AND U19802 ( .A(n19617), .B(n19618), .Z(n19615) );
  AND U19803 ( .A(a[5]), .B(b[11]), .Z(n19614) );
  XOR U19804 ( .A(n19619), .B(n19523), .Z(n19525) );
  XOR U19805 ( .A(n19620), .B(n19621), .Z(n19523) );
  AND U19806 ( .A(n19622), .B(n19623), .Z(n19620) );
  AND U19807 ( .A(a[6]), .B(b[10]), .Z(n19619) );
  XOR U19808 ( .A(n19624), .B(n19528), .Z(n19530) );
  XOR U19809 ( .A(n19625), .B(n19626), .Z(n19528) );
  AND U19810 ( .A(n19627), .B(n19628), .Z(n19625) );
  AND U19811 ( .A(a[7]), .B(b[9]), .Z(n19624) );
  XOR U19812 ( .A(n19629), .B(n19533), .Z(n19535) );
  XOR U19813 ( .A(n19630), .B(n19631), .Z(n19533) );
  AND U19814 ( .A(n19632), .B(n19633), .Z(n19630) );
  AND U19815 ( .A(b[8]), .B(a[8]), .Z(n19629) );
  XOR U19816 ( .A(n19634), .B(n19538), .Z(n19540) );
  XOR U19817 ( .A(n19635), .B(n19636), .Z(n19538) );
  AND U19818 ( .A(n19637), .B(n19638), .Z(n19635) );
  AND U19819 ( .A(a[9]), .B(b[7]), .Z(n19634) );
  XOR U19820 ( .A(n19639), .B(n19543), .Z(n19545) );
  XOR U19821 ( .A(n19640), .B(n19641), .Z(n19543) );
  AND U19822 ( .A(n19642), .B(n19643), .Z(n19640) );
  AND U19823 ( .A(b[6]), .B(a[10]), .Z(n19639) );
  XOR U19824 ( .A(n19644), .B(n19548), .Z(n19550) );
  XOR U19825 ( .A(n19645), .B(n19646), .Z(n19548) );
  AND U19826 ( .A(n19647), .B(n19648), .Z(n19645) );
  AND U19827 ( .A(a[11]), .B(b[5]), .Z(n19644) );
  XOR U19828 ( .A(n19649), .B(n19553), .Z(n19555) );
  XOR U19829 ( .A(n19650), .B(n19651), .Z(n19553) );
  AND U19830 ( .A(n19652), .B(n19653), .Z(n19650) );
  AND U19831 ( .A(b[4]), .B(a[12]), .Z(n19649) );
  XNOR U19832 ( .A(n19654), .B(n19655), .Z(n19567) );
  NANDN U19833 ( .A(n19656), .B(n19657), .Z(n19655) );
  XOR U19834 ( .A(n19658), .B(n19558), .Z(n19560) );
  XNOR U19835 ( .A(n19659), .B(n19660), .Z(n19558) );
  AND U19836 ( .A(n19661), .B(n19662), .Z(n19659) );
  AND U19837 ( .A(a[13]), .B(b[3]), .Z(n19658) );
  XOR U19838 ( .A(n19574), .B(n19573), .Z(c[111]) );
  XOR U19839 ( .A(sreg[143]), .B(n19572), .Z(n19573) );
  XOR U19840 ( .A(n19579), .B(n19663), .Z(n19574) );
  XNOR U19841 ( .A(n19578), .B(n19572), .Z(n19663) );
  XOR U19842 ( .A(n19664), .B(n19665), .Z(n19572) );
  NOR U19843 ( .A(n19666), .B(n19667), .Z(n19664) );
  NAND U19844 ( .A(a[15]), .B(b[0]), .Z(n19578) );
  XNOR U19845 ( .A(n19656), .B(n19657), .Z(n19579) );
  XOR U19846 ( .A(n19654), .B(n19668), .Z(n19657) );
  NAND U19847 ( .A(b[1]), .B(a[14]), .Z(n19668) );
  XOR U19848 ( .A(n19662), .B(n19669), .Z(n19656) );
  XOR U19849 ( .A(n19654), .B(n19661), .Z(n19669) );
  XNOR U19850 ( .A(n19670), .B(n19660), .Z(n19661) );
  AND U19851 ( .A(b[2]), .B(a[13]), .Z(n19670) );
  NANDN U19852 ( .A(n19671), .B(n19672), .Z(n19654) );
  XOR U19853 ( .A(n19660), .B(n19652), .Z(n19673) );
  XNOR U19854 ( .A(n19651), .B(n19647), .Z(n19674) );
  XNOR U19855 ( .A(n19646), .B(n19642), .Z(n19675) );
  XNOR U19856 ( .A(n19641), .B(n19637), .Z(n19676) );
  XNOR U19857 ( .A(n19636), .B(n19632), .Z(n19677) );
  XNOR U19858 ( .A(n19631), .B(n19627), .Z(n19678) );
  XNOR U19859 ( .A(n19626), .B(n19622), .Z(n19679) );
  XNOR U19860 ( .A(n19621), .B(n19617), .Z(n19680) );
  XNOR U19861 ( .A(n19616), .B(n19612), .Z(n19681) );
  XNOR U19862 ( .A(n19611), .B(n19607), .Z(n19682) );
  XNOR U19863 ( .A(n19606), .B(n19602), .Z(n19683) );
  XNOR U19864 ( .A(n19601), .B(n19597), .Z(n19684) );
  XOR U19865 ( .A(n19685), .B(n19596), .Z(n19597) );
  AND U19866 ( .A(a[0]), .B(b[15]), .Z(n19685) );
  XOR U19867 ( .A(n19686), .B(n19596), .Z(n19598) );
  XNOR U19868 ( .A(n19687), .B(n19688), .Z(n19596) );
  AND U19869 ( .A(n19689), .B(n19690), .Z(n19687) );
  AND U19870 ( .A(a[1]), .B(b[14]), .Z(n19686) );
  XOR U19871 ( .A(n19691), .B(n19601), .Z(n19603) );
  XOR U19872 ( .A(n19692), .B(n19693), .Z(n19601) );
  AND U19873 ( .A(n19694), .B(n19695), .Z(n19692) );
  AND U19874 ( .A(a[2]), .B(b[13]), .Z(n19691) );
  XOR U19875 ( .A(n19696), .B(n19606), .Z(n19608) );
  XOR U19876 ( .A(n19697), .B(n19698), .Z(n19606) );
  AND U19877 ( .A(n19699), .B(n19700), .Z(n19697) );
  AND U19878 ( .A(a[3]), .B(b[12]), .Z(n19696) );
  XOR U19879 ( .A(n19701), .B(n19611), .Z(n19613) );
  XOR U19880 ( .A(n19702), .B(n19703), .Z(n19611) );
  AND U19881 ( .A(n19704), .B(n19705), .Z(n19702) );
  AND U19882 ( .A(a[4]), .B(b[11]), .Z(n19701) );
  XOR U19883 ( .A(n19706), .B(n19616), .Z(n19618) );
  XOR U19884 ( .A(n19707), .B(n19708), .Z(n19616) );
  AND U19885 ( .A(n19709), .B(n19710), .Z(n19707) );
  AND U19886 ( .A(a[5]), .B(b[10]), .Z(n19706) );
  XOR U19887 ( .A(n19711), .B(n19621), .Z(n19623) );
  XOR U19888 ( .A(n19712), .B(n19713), .Z(n19621) );
  AND U19889 ( .A(n19714), .B(n19715), .Z(n19712) );
  AND U19890 ( .A(a[6]), .B(b[9]), .Z(n19711) );
  XOR U19891 ( .A(n19716), .B(n19626), .Z(n19628) );
  XOR U19892 ( .A(n19717), .B(n19718), .Z(n19626) );
  AND U19893 ( .A(n19719), .B(n19720), .Z(n19717) );
  AND U19894 ( .A(a[7]), .B(b[8]), .Z(n19716) );
  XOR U19895 ( .A(n19721), .B(n19631), .Z(n19633) );
  XOR U19896 ( .A(n19722), .B(n19723), .Z(n19631) );
  AND U19897 ( .A(n19724), .B(n19725), .Z(n19722) );
  AND U19898 ( .A(b[7]), .B(a[8]), .Z(n19721) );
  XOR U19899 ( .A(n19726), .B(n19636), .Z(n19638) );
  XOR U19900 ( .A(n19727), .B(n19728), .Z(n19636) );
  AND U19901 ( .A(n19729), .B(n19730), .Z(n19727) );
  AND U19902 ( .A(a[9]), .B(b[6]), .Z(n19726) );
  XOR U19903 ( .A(n19731), .B(n19641), .Z(n19643) );
  XOR U19904 ( .A(n19732), .B(n19733), .Z(n19641) );
  AND U19905 ( .A(n19734), .B(n19735), .Z(n19732) );
  AND U19906 ( .A(b[5]), .B(a[10]), .Z(n19731) );
  XOR U19907 ( .A(n19736), .B(n19646), .Z(n19648) );
  XOR U19908 ( .A(n19737), .B(n19738), .Z(n19646) );
  AND U19909 ( .A(n19739), .B(n19740), .Z(n19737) );
  AND U19910 ( .A(a[11]), .B(b[4]), .Z(n19736) );
  XNOR U19911 ( .A(n19741), .B(n19742), .Z(n19660) );
  NANDN U19912 ( .A(n19743), .B(n19744), .Z(n19742) );
  XOR U19913 ( .A(n19745), .B(n19651), .Z(n19653) );
  XNOR U19914 ( .A(n19746), .B(n19747), .Z(n19651) );
  AND U19915 ( .A(n19748), .B(n19749), .Z(n19746) );
  AND U19916 ( .A(b[3]), .B(a[12]), .Z(n19745) );
  XOR U19917 ( .A(n19667), .B(n19666), .Z(c[110]) );
  XOR U19918 ( .A(sreg[142]), .B(n19665), .Z(n19666) );
  XOR U19919 ( .A(n19672), .B(n19750), .Z(n19667) );
  XNOR U19920 ( .A(n19671), .B(n19665), .Z(n19750) );
  XOR U19921 ( .A(n19751), .B(n19752), .Z(n19665) );
  NOR U19922 ( .A(n19753), .B(n19754), .Z(n19751) );
  NAND U19923 ( .A(a[14]), .B(b[0]), .Z(n19671) );
  XNOR U19924 ( .A(n19743), .B(n19744), .Z(n19672) );
  XOR U19925 ( .A(n19741), .B(n19755), .Z(n19744) );
  NAND U19926 ( .A(a[13]), .B(b[1]), .Z(n19755) );
  XOR U19927 ( .A(n19749), .B(n19756), .Z(n19743) );
  XOR U19928 ( .A(n19741), .B(n19748), .Z(n19756) );
  XNOR U19929 ( .A(n19757), .B(n19747), .Z(n19748) );
  AND U19930 ( .A(b[2]), .B(a[12]), .Z(n19757) );
  NANDN U19931 ( .A(n19758), .B(n19759), .Z(n19741) );
  XOR U19932 ( .A(n19747), .B(n19739), .Z(n19760) );
  XNOR U19933 ( .A(n19738), .B(n19734), .Z(n19761) );
  XNOR U19934 ( .A(n19733), .B(n19729), .Z(n19762) );
  XNOR U19935 ( .A(n19728), .B(n19724), .Z(n19763) );
  XNOR U19936 ( .A(n19723), .B(n19719), .Z(n19764) );
  XNOR U19937 ( .A(n19718), .B(n19714), .Z(n19765) );
  XNOR U19938 ( .A(n19713), .B(n19709), .Z(n19766) );
  XNOR U19939 ( .A(n19708), .B(n19704), .Z(n19767) );
  XNOR U19940 ( .A(n19703), .B(n19699), .Z(n19768) );
  XNOR U19941 ( .A(n19698), .B(n19694), .Z(n19769) );
  XNOR U19942 ( .A(n19693), .B(n19689), .Z(n19770) );
  XNOR U19943 ( .A(n19771), .B(n19688), .Z(n19689) );
  AND U19944 ( .A(a[0]), .B(b[14]), .Z(n19771) );
  XNOR U19945 ( .A(n19772), .B(n19688), .Z(n19690) );
  XNOR U19946 ( .A(n19773), .B(n19774), .Z(n19688) );
  AND U19947 ( .A(n19775), .B(n19776), .Z(n19773) );
  AND U19948 ( .A(a[1]), .B(b[13]), .Z(n19772) );
  XOR U19949 ( .A(n19777), .B(n19693), .Z(n19695) );
  XOR U19950 ( .A(n19778), .B(n19779), .Z(n19693) );
  AND U19951 ( .A(n19780), .B(n19781), .Z(n19778) );
  AND U19952 ( .A(a[2]), .B(b[12]), .Z(n19777) );
  XOR U19953 ( .A(n19782), .B(n19698), .Z(n19700) );
  XOR U19954 ( .A(n19783), .B(n19784), .Z(n19698) );
  AND U19955 ( .A(n19785), .B(n19786), .Z(n19783) );
  AND U19956 ( .A(a[3]), .B(b[11]), .Z(n19782) );
  XOR U19957 ( .A(n19787), .B(n19703), .Z(n19705) );
  XOR U19958 ( .A(n19788), .B(n19789), .Z(n19703) );
  AND U19959 ( .A(n19790), .B(n19791), .Z(n19788) );
  AND U19960 ( .A(a[4]), .B(b[10]), .Z(n19787) );
  XOR U19961 ( .A(n19792), .B(n19708), .Z(n19710) );
  XOR U19962 ( .A(n19793), .B(n19794), .Z(n19708) );
  AND U19963 ( .A(n19795), .B(n19796), .Z(n19793) );
  AND U19964 ( .A(a[5]), .B(b[9]), .Z(n19792) );
  XOR U19965 ( .A(n19797), .B(n19713), .Z(n19715) );
  XOR U19966 ( .A(n19798), .B(n19799), .Z(n19713) );
  AND U19967 ( .A(n19800), .B(n19801), .Z(n19798) );
  AND U19968 ( .A(a[6]), .B(b[8]), .Z(n19797) );
  XOR U19969 ( .A(n19802), .B(n19718), .Z(n19720) );
  XOR U19970 ( .A(n19803), .B(n19804), .Z(n19718) );
  AND U19971 ( .A(n19805), .B(n19806), .Z(n19803) );
  AND U19972 ( .A(a[7]), .B(b[7]), .Z(n19802) );
  XOR U19973 ( .A(n19807), .B(n19723), .Z(n19725) );
  XOR U19974 ( .A(n19808), .B(n19809), .Z(n19723) );
  AND U19975 ( .A(n19810), .B(n19811), .Z(n19808) );
  AND U19976 ( .A(b[6]), .B(a[8]), .Z(n19807) );
  XOR U19977 ( .A(n19812), .B(n19728), .Z(n19730) );
  XOR U19978 ( .A(n19813), .B(n19814), .Z(n19728) );
  AND U19979 ( .A(n19815), .B(n19816), .Z(n19813) );
  AND U19980 ( .A(a[9]), .B(b[5]), .Z(n19812) );
  XOR U19981 ( .A(n19817), .B(n19733), .Z(n19735) );
  XOR U19982 ( .A(n19818), .B(n19819), .Z(n19733) );
  AND U19983 ( .A(n19820), .B(n19821), .Z(n19818) );
  AND U19984 ( .A(b[4]), .B(a[10]), .Z(n19817) );
  XNOR U19985 ( .A(n19822), .B(n19823), .Z(n19747) );
  NANDN U19986 ( .A(n19824), .B(n19825), .Z(n19823) );
  XOR U19987 ( .A(n19826), .B(n19738), .Z(n19740) );
  XNOR U19988 ( .A(n19827), .B(n19828), .Z(n19738) );
  AND U19989 ( .A(n19829), .B(n19830), .Z(n19827) );
  AND U19990 ( .A(a[11]), .B(b[3]), .Z(n19826) );
  XOR U19991 ( .A(n19754), .B(n19753), .Z(c[109]) );
  XOR U19992 ( .A(sreg[141]), .B(n19752), .Z(n19753) );
  XOR U19993 ( .A(n19759), .B(n19831), .Z(n19754) );
  XNOR U19994 ( .A(n19758), .B(n19752), .Z(n19831) );
  XOR U19995 ( .A(n19832), .B(n19833), .Z(n19752) );
  NOR U19996 ( .A(n19834), .B(n19835), .Z(n19832) );
  NAND U19997 ( .A(a[13]), .B(b[0]), .Z(n19758) );
  XNOR U19998 ( .A(n19824), .B(n19825), .Z(n19759) );
  XOR U19999 ( .A(n19822), .B(n19836), .Z(n19825) );
  NAND U20000 ( .A(b[1]), .B(a[12]), .Z(n19836) );
  XOR U20001 ( .A(n19830), .B(n19837), .Z(n19824) );
  XOR U20002 ( .A(n19822), .B(n19829), .Z(n19837) );
  XNOR U20003 ( .A(n19838), .B(n19828), .Z(n19829) );
  AND U20004 ( .A(b[2]), .B(a[11]), .Z(n19838) );
  NANDN U20005 ( .A(n19839), .B(n19840), .Z(n19822) );
  XOR U20006 ( .A(n19828), .B(n19820), .Z(n19841) );
  XNOR U20007 ( .A(n19819), .B(n19815), .Z(n19842) );
  XNOR U20008 ( .A(n19814), .B(n19810), .Z(n19843) );
  XNOR U20009 ( .A(n19809), .B(n19805), .Z(n19844) );
  XNOR U20010 ( .A(n19804), .B(n19800), .Z(n19845) );
  XNOR U20011 ( .A(n19799), .B(n19795), .Z(n19846) );
  XNOR U20012 ( .A(n19794), .B(n19790), .Z(n19847) );
  XNOR U20013 ( .A(n19789), .B(n19785), .Z(n19848) );
  XNOR U20014 ( .A(n19784), .B(n19780), .Z(n19849) );
  XNOR U20015 ( .A(n19779), .B(n19775), .Z(n19850) );
  XOR U20016 ( .A(n19851), .B(n19774), .Z(n19775) );
  AND U20017 ( .A(a[0]), .B(b[13]), .Z(n19851) );
  XOR U20018 ( .A(n19852), .B(n19774), .Z(n19776) );
  XNOR U20019 ( .A(n19853), .B(n19854), .Z(n19774) );
  AND U20020 ( .A(n19855), .B(n19856), .Z(n19853) );
  AND U20021 ( .A(a[1]), .B(b[12]), .Z(n19852) );
  XOR U20022 ( .A(n19857), .B(n19779), .Z(n19781) );
  XOR U20023 ( .A(n19858), .B(n19859), .Z(n19779) );
  AND U20024 ( .A(n19860), .B(n19861), .Z(n19858) );
  AND U20025 ( .A(a[2]), .B(b[11]), .Z(n19857) );
  XOR U20026 ( .A(n19862), .B(n19784), .Z(n19786) );
  XOR U20027 ( .A(n19863), .B(n19864), .Z(n19784) );
  AND U20028 ( .A(n19865), .B(n19866), .Z(n19863) );
  AND U20029 ( .A(a[3]), .B(b[10]), .Z(n19862) );
  XOR U20030 ( .A(n19867), .B(n19789), .Z(n19791) );
  XOR U20031 ( .A(n19868), .B(n19869), .Z(n19789) );
  AND U20032 ( .A(n19870), .B(n19871), .Z(n19868) );
  AND U20033 ( .A(a[4]), .B(b[9]), .Z(n19867) );
  XOR U20034 ( .A(n19872), .B(n19794), .Z(n19796) );
  XOR U20035 ( .A(n19873), .B(n19874), .Z(n19794) );
  AND U20036 ( .A(n19875), .B(n19876), .Z(n19873) );
  AND U20037 ( .A(a[5]), .B(b[8]), .Z(n19872) );
  XOR U20038 ( .A(n19877), .B(n19799), .Z(n19801) );
  XOR U20039 ( .A(n19878), .B(n19879), .Z(n19799) );
  AND U20040 ( .A(n19880), .B(n19881), .Z(n19878) );
  AND U20041 ( .A(a[6]), .B(b[7]), .Z(n19877) );
  XOR U20042 ( .A(n19882), .B(n19804), .Z(n19806) );
  XOR U20043 ( .A(n19883), .B(n19884), .Z(n19804) );
  AND U20044 ( .A(n19885), .B(n19886), .Z(n19883) );
  AND U20045 ( .A(a[7]), .B(b[6]), .Z(n19882) );
  XOR U20046 ( .A(n19887), .B(n19809), .Z(n19811) );
  XOR U20047 ( .A(n19888), .B(n19889), .Z(n19809) );
  AND U20048 ( .A(n19890), .B(n19891), .Z(n19888) );
  AND U20049 ( .A(b[5]), .B(a[8]), .Z(n19887) );
  XOR U20050 ( .A(n19892), .B(n19814), .Z(n19816) );
  XOR U20051 ( .A(n19893), .B(n19894), .Z(n19814) );
  AND U20052 ( .A(n19895), .B(n19896), .Z(n19893) );
  AND U20053 ( .A(a[9]), .B(b[4]), .Z(n19892) );
  XNOR U20054 ( .A(n19897), .B(n19898), .Z(n19828) );
  NANDN U20055 ( .A(n19899), .B(n19900), .Z(n19898) );
  XOR U20056 ( .A(n19901), .B(n19819), .Z(n19821) );
  XNOR U20057 ( .A(n19902), .B(n19903), .Z(n19819) );
  AND U20058 ( .A(n19904), .B(n19905), .Z(n19902) );
  AND U20059 ( .A(b[3]), .B(a[10]), .Z(n19901) );
  XOR U20060 ( .A(n19835), .B(n19834), .Z(c[108]) );
  XOR U20061 ( .A(sreg[140]), .B(n19833), .Z(n19834) );
  XOR U20062 ( .A(n19840), .B(n19906), .Z(n19835) );
  XNOR U20063 ( .A(n19839), .B(n19833), .Z(n19906) );
  XOR U20064 ( .A(n19907), .B(n19908), .Z(n19833) );
  NOR U20065 ( .A(n19909), .B(n19910), .Z(n19907) );
  NAND U20066 ( .A(a[12]), .B(b[0]), .Z(n19839) );
  XNOR U20067 ( .A(n19899), .B(n19900), .Z(n19840) );
  XOR U20068 ( .A(n19897), .B(n19911), .Z(n19900) );
  NAND U20069 ( .A(a[11]), .B(b[1]), .Z(n19911) );
  XOR U20070 ( .A(n19905), .B(n19912), .Z(n19899) );
  XOR U20071 ( .A(n19897), .B(n19904), .Z(n19912) );
  XNOR U20072 ( .A(n19913), .B(n19903), .Z(n19904) );
  AND U20073 ( .A(b[2]), .B(a[10]), .Z(n19913) );
  NANDN U20074 ( .A(n19914), .B(n19915), .Z(n19897) );
  XOR U20075 ( .A(n19903), .B(n19895), .Z(n19916) );
  XNOR U20076 ( .A(n19894), .B(n19890), .Z(n19917) );
  XNOR U20077 ( .A(n19889), .B(n19885), .Z(n19918) );
  XNOR U20078 ( .A(n19884), .B(n19880), .Z(n19919) );
  XNOR U20079 ( .A(n19879), .B(n19875), .Z(n19920) );
  XNOR U20080 ( .A(n19874), .B(n19870), .Z(n19921) );
  XNOR U20081 ( .A(n19869), .B(n19865), .Z(n19922) );
  XNOR U20082 ( .A(n19864), .B(n19860), .Z(n19923) );
  XNOR U20083 ( .A(n19859), .B(n19855), .Z(n19924) );
  XNOR U20084 ( .A(n19925), .B(n19854), .Z(n19855) );
  AND U20085 ( .A(a[0]), .B(b[12]), .Z(n19925) );
  XNOR U20086 ( .A(n19926), .B(n19854), .Z(n19856) );
  XNOR U20087 ( .A(n19927), .B(n19928), .Z(n19854) );
  AND U20088 ( .A(n19929), .B(n19930), .Z(n19927) );
  AND U20089 ( .A(a[1]), .B(b[11]), .Z(n19926) );
  XOR U20090 ( .A(n19931), .B(n19859), .Z(n19861) );
  XOR U20091 ( .A(n19932), .B(n19933), .Z(n19859) );
  AND U20092 ( .A(n19934), .B(n19935), .Z(n19932) );
  AND U20093 ( .A(a[2]), .B(b[10]), .Z(n19931) );
  XOR U20094 ( .A(n19936), .B(n19864), .Z(n19866) );
  XOR U20095 ( .A(n19937), .B(n19938), .Z(n19864) );
  AND U20096 ( .A(n19939), .B(n19940), .Z(n19937) );
  AND U20097 ( .A(a[3]), .B(b[9]), .Z(n19936) );
  XOR U20098 ( .A(n19941), .B(n19869), .Z(n19871) );
  XOR U20099 ( .A(n19942), .B(n19943), .Z(n19869) );
  AND U20100 ( .A(n19944), .B(n19945), .Z(n19942) );
  AND U20101 ( .A(a[4]), .B(b[8]), .Z(n19941) );
  XOR U20102 ( .A(n19946), .B(n19874), .Z(n19876) );
  XOR U20103 ( .A(n19947), .B(n19948), .Z(n19874) );
  AND U20104 ( .A(n19949), .B(n19950), .Z(n19947) );
  AND U20105 ( .A(a[5]), .B(b[7]), .Z(n19946) );
  XOR U20106 ( .A(n19951), .B(n19879), .Z(n19881) );
  XOR U20107 ( .A(n19952), .B(n19953), .Z(n19879) );
  AND U20108 ( .A(n19954), .B(n19955), .Z(n19952) );
  AND U20109 ( .A(b[6]), .B(a[6]), .Z(n19951) );
  XOR U20110 ( .A(n19956), .B(n19884), .Z(n19886) );
  XOR U20111 ( .A(n19957), .B(n19958), .Z(n19884) );
  AND U20112 ( .A(n19959), .B(n19960), .Z(n19957) );
  AND U20113 ( .A(a[7]), .B(b[5]), .Z(n19956) );
  XOR U20114 ( .A(n19961), .B(n19889), .Z(n19891) );
  XOR U20115 ( .A(n19962), .B(n19963), .Z(n19889) );
  AND U20116 ( .A(n19964), .B(n19965), .Z(n19962) );
  AND U20117 ( .A(b[4]), .B(a[8]), .Z(n19961) );
  XNOR U20118 ( .A(n19966), .B(n19967), .Z(n19903) );
  NANDN U20119 ( .A(n19968), .B(n19969), .Z(n19967) );
  XOR U20120 ( .A(n19970), .B(n19894), .Z(n19896) );
  XNOR U20121 ( .A(n19971), .B(n19972), .Z(n19894) );
  AND U20122 ( .A(n19973), .B(n19974), .Z(n19971) );
  AND U20123 ( .A(a[9]), .B(b[3]), .Z(n19970) );
  XOR U20124 ( .A(n19910), .B(n19909), .Z(c[107]) );
  XOR U20125 ( .A(sreg[139]), .B(n19908), .Z(n19909) );
  XOR U20126 ( .A(n19915), .B(n19975), .Z(n19910) );
  XNOR U20127 ( .A(n19914), .B(n19908), .Z(n19975) );
  XOR U20128 ( .A(n19976), .B(n19977), .Z(n19908) );
  NOR U20129 ( .A(n19978), .B(n19979), .Z(n19976) );
  NAND U20130 ( .A(a[11]), .B(b[0]), .Z(n19914) );
  XNOR U20131 ( .A(n19968), .B(n19969), .Z(n19915) );
  XOR U20132 ( .A(n19966), .B(n19980), .Z(n19969) );
  NAND U20133 ( .A(b[1]), .B(a[10]), .Z(n19980) );
  XOR U20134 ( .A(n19974), .B(n19981), .Z(n19968) );
  XOR U20135 ( .A(n19966), .B(n19973), .Z(n19981) );
  XNOR U20136 ( .A(n19982), .B(n19972), .Z(n19973) );
  AND U20137 ( .A(b[2]), .B(a[9]), .Z(n19982) );
  NANDN U20138 ( .A(n19983), .B(n19984), .Z(n19966) );
  XOR U20139 ( .A(n19972), .B(n19964), .Z(n19985) );
  XNOR U20140 ( .A(n19963), .B(n19959), .Z(n19986) );
  XNOR U20141 ( .A(n19958), .B(n19954), .Z(n19987) );
  XNOR U20142 ( .A(n19953), .B(n19949), .Z(n19988) );
  XNOR U20143 ( .A(n19948), .B(n19944), .Z(n19989) );
  XNOR U20144 ( .A(n19943), .B(n19939), .Z(n19990) );
  XNOR U20145 ( .A(n19938), .B(n19934), .Z(n19991) );
  XNOR U20146 ( .A(n19933), .B(n19929), .Z(n19992) );
  XOR U20147 ( .A(n19993), .B(n19928), .Z(n19929) );
  AND U20148 ( .A(a[0]), .B(b[11]), .Z(n19993) );
  XOR U20149 ( .A(n19994), .B(n19928), .Z(n19930) );
  XNOR U20150 ( .A(n19995), .B(n19996), .Z(n19928) );
  AND U20151 ( .A(n19997), .B(n19998), .Z(n19995) );
  AND U20152 ( .A(a[1]), .B(b[10]), .Z(n19994) );
  XOR U20153 ( .A(n19999), .B(n19933), .Z(n19935) );
  XOR U20154 ( .A(n20000), .B(n20001), .Z(n19933) );
  AND U20155 ( .A(n20002), .B(n20003), .Z(n20000) );
  AND U20156 ( .A(a[2]), .B(b[9]), .Z(n19999) );
  XOR U20157 ( .A(n20004), .B(n19938), .Z(n19940) );
  XOR U20158 ( .A(n20005), .B(n20006), .Z(n19938) );
  AND U20159 ( .A(n20007), .B(n20008), .Z(n20005) );
  AND U20160 ( .A(a[3]), .B(b[8]), .Z(n20004) );
  XOR U20161 ( .A(n20009), .B(n19943), .Z(n19945) );
  XOR U20162 ( .A(n20010), .B(n20011), .Z(n19943) );
  AND U20163 ( .A(n20012), .B(n20013), .Z(n20010) );
  AND U20164 ( .A(a[4]), .B(b[7]), .Z(n20009) );
  XOR U20165 ( .A(n20014), .B(n19948), .Z(n19950) );
  XOR U20166 ( .A(n20015), .B(n20016), .Z(n19948) );
  AND U20167 ( .A(n20017), .B(n20018), .Z(n20015) );
  AND U20168 ( .A(a[5]), .B(b[6]), .Z(n20014) );
  XOR U20169 ( .A(n20019), .B(n19953), .Z(n19955) );
  XOR U20170 ( .A(n20020), .B(n20021), .Z(n19953) );
  AND U20171 ( .A(n20022), .B(n20023), .Z(n20020) );
  AND U20172 ( .A(b[5]), .B(a[6]), .Z(n20019) );
  XOR U20173 ( .A(n20024), .B(n19958), .Z(n19960) );
  XOR U20174 ( .A(n20025), .B(n20026), .Z(n19958) );
  AND U20175 ( .A(n20027), .B(n20028), .Z(n20025) );
  AND U20176 ( .A(a[7]), .B(b[4]), .Z(n20024) );
  XNOR U20177 ( .A(n20029), .B(n20030), .Z(n19972) );
  NANDN U20178 ( .A(n20031), .B(n20032), .Z(n20030) );
  XOR U20179 ( .A(n20033), .B(n19963), .Z(n19965) );
  XNOR U20180 ( .A(n20034), .B(n20035), .Z(n19963) );
  AND U20181 ( .A(n20036), .B(n20037), .Z(n20034) );
  AND U20182 ( .A(b[3]), .B(a[8]), .Z(n20033) );
  XOR U20183 ( .A(n19979), .B(n19978), .Z(c[106]) );
  XOR U20184 ( .A(sreg[138]), .B(n19977), .Z(n19978) );
  XOR U20185 ( .A(n19984), .B(n20038), .Z(n19979) );
  XNOR U20186 ( .A(n19983), .B(n19977), .Z(n20038) );
  XOR U20187 ( .A(n20039), .B(n20040), .Z(n19977) );
  NOR U20188 ( .A(n20041), .B(n20042), .Z(n20039) );
  NAND U20189 ( .A(a[10]), .B(b[0]), .Z(n19983) );
  XNOR U20190 ( .A(n20031), .B(n20032), .Z(n19984) );
  XOR U20191 ( .A(n20029), .B(n20043), .Z(n20032) );
  NAND U20192 ( .A(a[9]), .B(b[1]), .Z(n20043) );
  XOR U20193 ( .A(n20037), .B(n20044), .Z(n20031) );
  XOR U20194 ( .A(n20029), .B(n20036), .Z(n20044) );
  XNOR U20195 ( .A(n20045), .B(n20035), .Z(n20036) );
  AND U20196 ( .A(b[2]), .B(a[8]), .Z(n20045) );
  NANDN U20197 ( .A(n20046), .B(n20047), .Z(n20029) );
  XOR U20198 ( .A(n20035), .B(n20027), .Z(n20048) );
  XNOR U20199 ( .A(n20026), .B(n20022), .Z(n20049) );
  XNOR U20200 ( .A(n20021), .B(n20017), .Z(n20050) );
  XNOR U20201 ( .A(n20016), .B(n20012), .Z(n20051) );
  XNOR U20202 ( .A(n20011), .B(n20007), .Z(n20052) );
  XNOR U20203 ( .A(n20006), .B(n20002), .Z(n20053) );
  XNOR U20204 ( .A(n20001), .B(n19997), .Z(n20054) );
  XNOR U20205 ( .A(n20055), .B(n19996), .Z(n19997) );
  AND U20206 ( .A(a[0]), .B(b[10]), .Z(n20055) );
  XNOR U20207 ( .A(n20056), .B(n19996), .Z(n19998) );
  XNOR U20208 ( .A(n20057), .B(n20058), .Z(n19996) );
  AND U20209 ( .A(n20059), .B(n20060), .Z(n20057) );
  AND U20210 ( .A(a[1]), .B(b[9]), .Z(n20056) );
  XOR U20211 ( .A(n20061), .B(n20001), .Z(n20003) );
  XOR U20212 ( .A(n20062), .B(n20063), .Z(n20001) );
  AND U20213 ( .A(n20064), .B(n20065), .Z(n20062) );
  AND U20214 ( .A(a[2]), .B(b[8]), .Z(n20061) );
  XOR U20215 ( .A(n20066), .B(n20006), .Z(n20008) );
  XOR U20216 ( .A(n20067), .B(n20068), .Z(n20006) );
  AND U20217 ( .A(n20069), .B(n20070), .Z(n20067) );
  AND U20218 ( .A(a[3]), .B(b[7]), .Z(n20066) );
  XOR U20219 ( .A(n20071), .B(n20011), .Z(n20013) );
  XOR U20220 ( .A(n20072), .B(n20073), .Z(n20011) );
  AND U20221 ( .A(n20074), .B(n20075), .Z(n20072) );
  AND U20222 ( .A(a[4]), .B(b[6]), .Z(n20071) );
  XOR U20223 ( .A(n20076), .B(n20016), .Z(n20018) );
  XOR U20224 ( .A(n20077), .B(n20078), .Z(n20016) );
  AND U20225 ( .A(n20079), .B(n20080), .Z(n20077) );
  AND U20226 ( .A(a[5]), .B(b[5]), .Z(n20076) );
  XOR U20227 ( .A(n20081), .B(n20021), .Z(n20023) );
  XOR U20228 ( .A(n20082), .B(n20083), .Z(n20021) );
  AND U20229 ( .A(n20084), .B(n20085), .Z(n20082) );
  AND U20230 ( .A(b[4]), .B(a[6]), .Z(n20081) );
  XNOR U20231 ( .A(n20086), .B(n20087), .Z(n20035) );
  NANDN U20232 ( .A(n20088), .B(n20089), .Z(n20087) );
  XOR U20233 ( .A(n20090), .B(n20026), .Z(n20028) );
  XNOR U20234 ( .A(n20091), .B(n20092), .Z(n20026) );
  AND U20235 ( .A(n20093), .B(n20094), .Z(n20091) );
  AND U20236 ( .A(a[7]), .B(b[3]), .Z(n20090) );
  XOR U20237 ( .A(n20042), .B(n20041), .Z(c[105]) );
  XOR U20238 ( .A(sreg[137]), .B(n20040), .Z(n20041) );
  XOR U20239 ( .A(n20047), .B(n20095), .Z(n20042) );
  XNOR U20240 ( .A(n20046), .B(n20040), .Z(n20095) );
  XOR U20241 ( .A(n20096), .B(n20097), .Z(n20040) );
  NOR U20242 ( .A(n20098), .B(n20099), .Z(n20096) );
  NAND U20243 ( .A(a[9]), .B(b[0]), .Z(n20046) );
  XNOR U20244 ( .A(n20088), .B(n20089), .Z(n20047) );
  XOR U20245 ( .A(n20086), .B(n20100), .Z(n20089) );
  NAND U20246 ( .A(b[1]), .B(a[8]), .Z(n20100) );
  XOR U20247 ( .A(n20094), .B(n20101), .Z(n20088) );
  XOR U20248 ( .A(n20086), .B(n20093), .Z(n20101) );
  XNOR U20249 ( .A(n20102), .B(n20092), .Z(n20093) );
  AND U20250 ( .A(b[2]), .B(a[7]), .Z(n20102) );
  NANDN U20251 ( .A(n20103), .B(n20104), .Z(n20086) );
  XOR U20252 ( .A(n20092), .B(n20084), .Z(n20105) );
  XNOR U20253 ( .A(n20083), .B(n20079), .Z(n20106) );
  XNOR U20254 ( .A(n20078), .B(n20074), .Z(n20107) );
  XNOR U20255 ( .A(n20073), .B(n20069), .Z(n20108) );
  XNOR U20256 ( .A(n20068), .B(n20064), .Z(n20109) );
  XNOR U20257 ( .A(n20063), .B(n20059), .Z(n20110) );
  XOR U20258 ( .A(n20111), .B(n20058), .Z(n20059) );
  AND U20259 ( .A(a[0]), .B(b[9]), .Z(n20111) );
  XOR U20260 ( .A(n20112), .B(n20058), .Z(n20060) );
  XNOR U20261 ( .A(n20113), .B(n20114), .Z(n20058) );
  AND U20262 ( .A(n20115), .B(n20116), .Z(n20113) );
  AND U20263 ( .A(a[1]), .B(b[8]), .Z(n20112) );
  XOR U20264 ( .A(n20117), .B(n20063), .Z(n20065) );
  XOR U20265 ( .A(n20118), .B(n20119), .Z(n20063) );
  AND U20266 ( .A(n20120), .B(n20121), .Z(n20118) );
  AND U20267 ( .A(a[2]), .B(b[7]), .Z(n20117) );
  XOR U20268 ( .A(n20122), .B(n20068), .Z(n20070) );
  XOR U20269 ( .A(n20123), .B(n20124), .Z(n20068) );
  AND U20270 ( .A(n20125), .B(n20126), .Z(n20123) );
  AND U20271 ( .A(a[3]), .B(b[6]), .Z(n20122) );
  XOR U20272 ( .A(n20127), .B(n20073), .Z(n20075) );
  XOR U20273 ( .A(n20128), .B(n20129), .Z(n20073) );
  AND U20274 ( .A(n20130), .B(n20131), .Z(n20128) );
  AND U20275 ( .A(a[4]), .B(b[5]), .Z(n20127) );
  XOR U20276 ( .A(n20132), .B(n20078), .Z(n20080) );
  XOR U20277 ( .A(n20133), .B(n20134), .Z(n20078) );
  AND U20278 ( .A(n20135), .B(n20136), .Z(n20133) );
  AND U20279 ( .A(a[5]), .B(b[4]), .Z(n20132) );
  XNOR U20280 ( .A(n20137), .B(n20138), .Z(n20092) );
  NANDN U20281 ( .A(n20139), .B(n20140), .Z(n20138) );
  XOR U20282 ( .A(n20141), .B(n20083), .Z(n20085) );
  XNOR U20283 ( .A(n20142), .B(n20143), .Z(n20083) );
  AND U20284 ( .A(n20144), .B(n20145), .Z(n20142) );
  AND U20285 ( .A(b[3]), .B(a[6]), .Z(n20141) );
  XOR U20286 ( .A(n20099), .B(n20098), .Z(c[104]) );
  XOR U20287 ( .A(sreg[136]), .B(n20097), .Z(n20098) );
  XOR U20288 ( .A(n20104), .B(n20146), .Z(n20099) );
  XNOR U20289 ( .A(n20103), .B(n20097), .Z(n20146) );
  XOR U20290 ( .A(n20147), .B(n20148), .Z(n20097) );
  NOR U20291 ( .A(n20149), .B(n20150), .Z(n20147) );
  NAND U20292 ( .A(a[8]), .B(b[0]), .Z(n20103) );
  XNOR U20293 ( .A(n20139), .B(n20140), .Z(n20104) );
  XOR U20294 ( .A(n20137), .B(n20151), .Z(n20140) );
  NAND U20295 ( .A(a[7]), .B(b[1]), .Z(n20151) );
  XOR U20296 ( .A(n20145), .B(n20152), .Z(n20139) );
  XOR U20297 ( .A(n20137), .B(n20144), .Z(n20152) );
  XNOR U20298 ( .A(n20153), .B(n20143), .Z(n20144) );
  AND U20299 ( .A(b[2]), .B(a[6]), .Z(n20153) );
  NANDN U20300 ( .A(n20154), .B(n20155), .Z(n20137) );
  XOR U20301 ( .A(n20143), .B(n20135), .Z(n20156) );
  XNOR U20302 ( .A(n20134), .B(n20130), .Z(n20157) );
  XNOR U20303 ( .A(n20129), .B(n20125), .Z(n20158) );
  XNOR U20304 ( .A(n20124), .B(n20120), .Z(n20159) );
  XNOR U20305 ( .A(n20119), .B(n20115), .Z(n20160) );
  XNOR U20306 ( .A(n20161), .B(n20114), .Z(n20115) );
  AND U20307 ( .A(a[0]), .B(b[8]), .Z(n20161) );
  XNOR U20308 ( .A(n20162), .B(n20114), .Z(n20116) );
  XNOR U20309 ( .A(n20163), .B(n20164), .Z(n20114) );
  AND U20310 ( .A(n20165), .B(n20166), .Z(n20163) );
  AND U20311 ( .A(a[1]), .B(b[7]), .Z(n20162) );
  XOR U20312 ( .A(n20167), .B(n20119), .Z(n20121) );
  XOR U20313 ( .A(n20168), .B(n20169), .Z(n20119) );
  AND U20314 ( .A(n20170), .B(n20171), .Z(n20168) );
  AND U20315 ( .A(a[2]), .B(b[6]), .Z(n20167) );
  XOR U20316 ( .A(n20172), .B(n20124), .Z(n20126) );
  XOR U20317 ( .A(n20173), .B(n20174), .Z(n20124) );
  AND U20318 ( .A(n20175), .B(n20176), .Z(n20173) );
  AND U20319 ( .A(a[3]), .B(b[5]), .Z(n20172) );
  XOR U20320 ( .A(n20177), .B(n20129), .Z(n20131) );
  XOR U20321 ( .A(n20178), .B(n20179), .Z(n20129) );
  AND U20322 ( .A(n20180), .B(n20181), .Z(n20178) );
  AND U20323 ( .A(b[4]), .B(a[4]), .Z(n20177) );
  XNOR U20324 ( .A(n20182), .B(n20183), .Z(n20143) );
  NANDN U20325 ( .A(n20184), .B(n20185), .Z(n20183) );
  XOR U20326 ( .A(n20186), .B(n20134), .Z(n20136) );
  XNOR U20327 ( .A(n20187), .B(n20188), .Z(n20134) );
  AND U20328 ( .A(n20189), .B(n20190), .Z(n20187) );
  AND U20329 ( .A(a[5]), .B(b[3]), .Z(n20186) );
  XOR U20330 ( .A(n20150), .B(n20149), .Z(c[103]) );
  XOR U20331 ( .A(sreg[135]), .B(n20148), .Z(n20149) );
  XOR U20332 ( .A(n20155), .B(n20191), .Z(n20150) );
  XNOR U20333 ( .A(n20154), .B(n20148), .Z(n20191) );
  XOR U20334 ( .A(n20192), .B(n20193), .Z(n20148) );
  NOR U20335 ( .A(n20194), .B(n20195), .Z(n20192) );
  NAND U20336 ( .A(a[7]), .B(b[0]), .Z(n20154) );
  XNOR U20337 ( .A(n20184), .B(n20185), .Z(n20155) );
  XOR U20338 ( .A(n20182), .B(n20196), .Z(n20185) );
  NAND U20339 ( .A(b[1]), .B(a[6]), .Z(n20196) );
  XOR U20340 ( .A(n20190), .B(n20197), .Z(n20184) );
  XOR U20341 ( .A(n20182), .B(n20189), .Z(n20197) );
  XNOR U20342 ( .A(n20198), .B(n20188), .Z(n20189) );
  AND U20343 ( .A(b[2]), .B(a[5]), .Z(n20198) );
  NANDN U20344 ( .A(n20199), .B(n20200), .Z(n20182) );
  XOR U20345 ( .A(n20188), .B(n20180), .Z(n20201) );
  XNOR U20346 ( .A(n20179), .B(n20175), .Z(n20202) );
  XNOR U20347 ( .A(n20174), .B(n20170), .Z(n20203) );
  XNOR U20348 ( .A(n20169), .B(n20165), .Z(n20204) );
  XOR U20349 ( .A(n20205), .B(n20164), .Z(n20165) );
  AND U20350 ( .A(a[0]), .B(b[7]), .Z(n20205) );
  XOR U20351 ( .A(n20206), .B(n20164), .Z(n20166) );
  XNOR U20352 ( .A(n20207), .B(n20208), .Z(n20164) );
  AND U20353 ( .A(n20209), .B(n20210), .Z(n20207) );
  AND U20354 ( .A(a[1]), .B(b[6]), .Z(n20206) );
  XOR U20355 ( .A(n20211), .B(n20169), .Z(n20171) );
  XOR U20356 ( .A(n20212), .B(n20213), .Z(n20169) );
  AND U20357 ( .A(n20214), .B(n20215), .Z(n20212) );
  AND U20358 ( .A(a[2]), .B(b[5]), .Z(n20211) );
  XOR U20359 ( .A(n20216), .B(n20174), .Z(n20176) );
  XOR U20360 ( .A(n20217), .B(n20218), .Z(n20174) );
  AND U20361 ( .A(n20219), .B(n20220), .Z(n20217) );
  AND U20362 ( .A(a[3]), .B(b[4]), .Z(n20216) );
  XNOR U20363 ( .A(n20221), .B(n20222), .Z(n20188) );
  NANDN U20364 ( .A(n20223), .B(n20224), .Z(n20222) );
  XOR U20365 ( .A(n20225), .B(n20179), .Z(n20181) );
  XNOR U20366 ( .A(n20226), .B(n20227), .Z(n20179) );
  AND U20367 ( .A(n20228), .B(n20229), .Z(n20226) );
  AND U20368 ( .A(b[3]), .B(a[4]), .Z(n20225) );
  XOR U20369 ( .A(n20195), .B(n20194), .Z(c[102]) );
  XOR U20370 ( .A(sreg[134]), .B(n20193), .Z(n20194) );
  XOR U20371 ( .A(n20200), .B(n20230), .Z(n20195) );
  XNOR U20372 ( .A(n20199), .B(n20193), .Z(n20230) );
  XOR U20373 ( .A(n20231), .B(n20232), .Z(n20193) );
  NOR U20374 ( .A(n20233), .B(n20234), .Z(n20231) );
  NAND U20375 ( .A(a[6]), .B(b[0]), .Z(n20199) );
  XNOR U20376 ( .A(n20223), .B(n20224), .Z(n20200) );
  XOR U20377 ( .A(n20221), .B(n20235), .Z(n20224) );
  NAND U20378 ( .A(a[5]), .B(b[1]), .Z(n20235) );
  XOR U20379 ( .A(n20229), .B(n20236), .Z(n20223) );
  XOR U20380 ( .A(n20221), .B(n20228), .Z(n20236) );
  XNOR U20381 ( .A(n20237), .B(n20227), .Z(n20228) );
  AND U20382 ( .A(b[2]), .B(a[4]), .Z(n20237) );
  NANDN U20383 ( .A(n20238), .B(n20239), .Z(n20221) );
  XOR U20384 ( .A(n20227), .B(n20219), .Z(n20240) );
  XNOR U20385 ( .A(n20218), .B(n20214), .Z(n20241) );
  XNOR U20386 ( .A(n20213), .B(n20209), .Z(n20242) );
  XNOR U20387 ( .A(n20243), .B(n20208), .Z(n20209) );
  AND U20388 ( .A(a[0]), .B(b[6]), .Z(n20243) );
  XNOR U20389 ( .A(n20244), .B(n20208), .Z(n20210) );
  XNOR U20390 ( .A(n20245), .B(n20246), .Z(n20208) );
  AND U20391 ( .A(n20247), .B(n20248), .Z(n20245) );
  AND U20392 ( .A(a[1]), .B(b[5]), .Z(n20244) );
  XOR U20393 ( .A(n20249), .B(n20213), .Z(n20215) );
  XOR U20394 ( .A(n20250), .B(n20251), .Z(n20213) );
  AND U20395 ( .A(n20252), .B(n20253), .Z(n20250) );
  AND U20396 ( .A(a[2]), .B(b[4]), .Z(n20249) );
  XNOR U20397 ( .A(n20254), .B(n20255), .Z(n20227) );
  NANDN U20398 ( .A(n20256), .B(n20257), .Z(n20255) );
  XOR U20399 ( .A(n20258), .B(n20218), .Z(n20220) );
  XNOR U20400 ( .A(n20259), .B(n20260), .Z(n20218) );
  AND U20401 ( .A(n20261), .B(n20262), .Z(n20259) );
  AND U20402 ( .A(a[3]), .B(b[3]), .Z(n20258) );
  XOR U20403 ( .A(n20234), .B(n20233), .Z(c[101]) );
  XOR U20404 ( .A(sreg[133]), .B(n20232), .Z(n20233) );
  XOR U20405 ( .A(n20239), .B(n20263), .Z(n20234) );
  XNOR U20406 ( .A(n20238), .B(n20232), .Z(n20263) );
  XOR U20407 ( .A(n20264), .B(n20265), .Z(n20232) );
  NOR U20408 ( .A(n20266), .B(n20267), .Z(n20264) );
  NAND U20409 ( .A(a[5]), .B(b[0]), .Z(n20238) );
  XNOR U20410 ( .A(n20256), .B(n20257), .Z(n20239) );
  XOR U20411 ( .A(n20254), .B(n20268), .Z(n20257) );
  NAND U20412 ( .A(b[1]), .B(a[4]), .Z(n20268) );
  XOR U20413 ( .A(n20262), .B(n20269), .Z(n20256) );
  XOR U20414 ( .A(n20254), .B(n20261), .Z(n20269) );
  XNOR U20415 ( .A(n20270), .B(n20260), .Z(n20261) );
  AND U20416 ( .A(b[2]), .B(a[3]), .Z(n20270) );
  NANDN U20417 ( .A(n20271), .B(n20272), .Z(n20254) );
  XOR U20418 ( .A(n20260), .B(n20252), .Z(n20273) );
  XNOR U20419 ( .A(n20251), .B(n20247), .Z(n20274) );
  XOR U20420 ( .A(n20275), .B(n20246), .Z(n20247) );
  AND U20421 ( .A(a[0]), .B(b[5]), .Z(n20275) );
  XOR U20422 ( .A(n20276), .B(n20246), .Z(n20248) );
  XNOR U20423 ( .A(n20277), .B(n20278), .Z(n20246) );
  AND U20424 ( .A(n20279), .B(n20280), .Z(n20277) );
  AND U20425 ( .A(a[1]), .B(b[4]), .Z(n20276) );
  XNOR U20426 ( .A(n20281), .B(n20282), .Z(n20260) );
  NANDN U20427 ( .A(n20283), .B(n20284), .Z(n20282) );
  XOR U20428 ( .A(n20285), .B(n20251), .Z(n20253) );
  XNOR U20429 ( .A(n20286), .B(n20287), .Z(n20251) );
  AND U20430 ( .A(n20288), .B(n20289), .Z(n20286) );
  AND U20431 ( .A(a[2]), .B(b[3]), .Z(n20285) );
  XOR U20432 ( .A(n20267), .B(n20266), .Z(c[100]) );
  XOR U20433 ( .A(sreg[132]), .B(n20265), .Z(n20266) );
  XOR U20434 ( .A(n20272), .B(n20290), .Z(n20267) );
  XNOR U20435 ( .A(n20271), .B(n20265), .Z(n20290) );
  XOR U20436 ( .A(n20291), .B(n20292), .Z(n20265) );
  NOR U20437 ( .A(n17447), .B(n17446), .Z(n20291) );
  XOR U20438 ( .A(n20293), .B(n20294), .Z(n17446) );
  XNOR U20439 ( .A(n20295), .B(n20292), .Z(n20294) );
  XOR U20440 ( .A(sreg[131]), .B(n20292), .Z(n17447) );
  XOR U20441 ( .A(n20296), .B(n20297), .Z(n20292) );
  NOR U20442 ( .A(n17449), .B(n17448), .Z(n20296) );
  XOR U20443 ( .A(n20298), .B(n20299), .Z(n17448) );
  XOR U20444 ( .A(sreg[130]), .B(n20297), .Z(n17449) );
  XOR U20445 ( .A(n20301), .B(n20302), .Z(n20297) );
  NAND U20446 ( .A(n17450), .B(n17451), .Z(n20302) );
  XOR U20447 ( .A(sreg[129]), .B(n20301), .Z(n17451) );
  XNOR U20448 ( .A(n20301), .B(n20303), .Z(n17450) );
  XNOR U20449 ( .A(n20304), .B(n20305), .Z(n20303) );
  ANDN U20450 ( .B(sreg[128]), .A(n17452), .Z(n20301) );
  NAND U20451 ( .A(a[0]), .B(b[0]), .Z(n17452) );
  NAND U20452 ( .A(a[4]), .B(b[0]), .Z(n20271) );
  XNOR U20453 ( .A(n20283), .B(n20284), .Z(n20272) );
  XOR U20454 ( .A(n20281), .B(n20306), .Z(n20284) );
  NAND U20455 ( .A(a[3]), .B(b[1]), .Z(n20306) );
  XOR U20456 ( .A(n20289), .B(n20307), .Z(n20283) );
  XOR U20457 ( .A(n20281), .B(n20288), .Z(n20307) );
  XNOR U20458 ( .A(n20308), .B(n20287), .Z(n20288) );
  AND U20459 ( .A(b[2]), .B(a[2]), .Z(n20308) );
  NANDN U20460 ( .A(n20295), .B(n20293), .Z(n20281) );
  XNOR U20461 ( .A(n20309), .B(n20310), .Z(n20293) );
  NAND U20462 ( .A(a[3]), .B(b[0]), .Z(n20295) );
  XOR U20463 ( .A(n20287), .B(n20279), .Z(n20311) );
  XNOR U20464 ( .A(n20312), .B(n20278), .Z(n20279) );
  AND U20465 ( .A(a[0]), .B(b[4]), .Z(n20312) );
  XNOR U20466 ( .A(n20313), .B(n20314), .Z(n20287) );
  NANDN U20467 ( .A(n20309), .B(n20310), .Z(n20314) );
  XOR U20468 ( .A(n20313), .B(n20315), .Z(n20310) );
  NAND U20469 ( .A(b[1]), .B(a[2]), .Z(n20315) );
  XOR U20470 ( .A(n20316), .B(n20317), .Z(n20309) );
  XOR U20471 ( .A(n20313), .B(n20318), .Z(n20317) );
  NANDN U20472 ( .A(n20300), .B(n20298), .Z(n20313) );
  XNOR U20473 ( .A(n20319), .B(n20320), .Z(n20298) );
  NAND U20474 ( .A(a[2]), .B(b[0]), .Z(n20300) );
  XNOR U20475 ( .A(n20321), .B(n20278), .Z(n20280) );
  XNOR U20476 ( .A(n20322), .B(n20323), .Z(n20278) );
  AND U20477 ( .A(n20318), .B(n20316), .Z(n20322) );
  XOR U20478 ( .A(n20324), .B(n20323), .Z(n20316) );
  AND U20479 ( .A(a[0]), .B(b[3]), .Z(n20324) );
  XOR U20480 ( .A(n20325), .B(n20323), .Z(n20318) );
  XOR U20481 ( .A(n20326), .B(n20327), .Z(n20323) );
  NANDN U20482 ( .A(n20319), .B(n20320), .Z(n20327) );
  XOR U20483 ( .A(n20326), .B(n20328), .Z(n20320) );
  NAND U20484 ( .A(a[1]), .B(b[1]), .Z(n20328) );
  XNOR U20485 ( .A(n20326), .B(n20329), .Z(n20319) );
  NAND U20486 ( .A(b[2]), .B(a[0]), .Z(n20329) );
  OR U20487 ( .A(n20304), .B(n20305), .Z(n20326) );
  NAND U20488 ( .A(a[0]), .B(b[1]), .Z(n20305) );
  NAND U20489 ( .A(a[1]), .B(b[0]), .Z(n20304) );
  AND U20490 ( .A(b[2]), .B(a[1]), .Z(n20325) );
  AND U20491 ( .A(a[1]), .B(b[3]), .Z(n20321) );
endmodule

