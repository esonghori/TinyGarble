
module sum_N128_CC1 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506;

  XNOR U2 ( .A(a[3]), .B(n499), .Z(n67) );
  XNOR U3 ( .A(a[6]), .B(n490), .Z(n34) );
  XNOR U4 ( .A(a[9]), .B(n481), .Z(n1) );
  XNOR U5 ( .A(a[12]), .B(n472), .Z(n97) );
  XNOR U6 ( .A(a[15]), .B(n463), .Z(n94) );
  XNOR U7 ( .A(a[18]), .B(n454), .Z(n91) );
  XNOR U8 ( .A(a[21]), .B(n445), .Z(n87) );
  XNOR U9 ( .A(a[24]), .B(n436), .Z(n84) );
  XNOR U10 ( .A(a[27]), .B(n427), .Z(n81) );
  XNOR U11 ( .A(a[30]), .B(n418), .Z(n77) );
  XNOR U12 ( .A(a[33]), .B(n409), .Z(n74) );
  XNOR U13 ( .A(a[36]), .B(n400), .Z(n71) );
  XNOR U14 ( .A(a[39]), .B(n391), .Z(n68) );
  XNOR U15 ( .A(a[42]), .B(n382), .Z(n64) );
  XNOR U16 ( .A(a[45]), .B(n373), .Z(n61) );
  XNOR U17 ( .A(a[48]), .B(n364), .Z(n58) );
  XNOR U18 ( .A(a[51]), .B(n355), .Z(n54) );
  XNOR U19 ( .A(a[54]), .B(n346), .Z(n51) );
  XNOR U20 ( .A(a[57]), .B(n337), .Z(n48) );
  XNOR U21 ( .A(a[60]), .B(n328), .Z(n44) );
  XNOR U22 ( .A(a[63]), .B(n319), .Z(n41) );
  XNOR U23 ( .A(a[66]), .B(n310), .Z(n38) );
  XNOR U24 ( .A(a[69]), .B(n301), .Z(n35) );
  XNOR U25 ( .A(a[72]), .B(n292), .Z(n31) );
  XNOR U26 ( .A(a[75]), .B(n283), .Z(n28) );
  XNOR U27 ( .A(a[78]), .B(n274), .Z(n25) );
  XNOR U28 ( .A(a[81]), .B(n265), .Z(n21) );
  XNOR U29 ( .A(a[84]), .B(n256), .Z(n18) );
  XNOR U30 ( .A(a[87]), .B(n247), .Z(n15) );
  XNOR U31 ( .A(a[90]), .B(n238), .Z(n11) );
  XNOR U32 ( .A(a[93]), .B(n229), .Z(n8) );
  XNOR U33 ( .A(a[96]), .B(n220), .Z(n5) );
  XNOR U34 ( .A(a[99]), .B(n211), .Z(n2) );
  XNOR U35 ( .A(a[102]), .B(n199), .Z(n201) );
  XNOR U36 ( .A(a[105]), .B(n187), .Z(n189) );
  XNOR U37 ( .A(a[108]), .B(n175), .Z(n177) );
  XNOR U38 ( .A(a[111]), .B(n162), .Z(n164) );
  XNOR U39 ( .A(a[114]), .B(n150), .Z(n152) );
  XNOR U40 ( .A(a[117]), .B(n138), .Z(n140) );
  XNOR U41 ( .A(a[120]), .B(n125), .Z(n127) );
  XNOR U42 ( .A(a[123]), .B(n113), .Z(n115) );
  XNOR U43 ( .A(a[4]), .B(n496), .Z(n56) );
  XNOR U44 ( .A(a[7]), .B(n487), .Z(n23) );
  XNOR U45 ( .A(a[10]), .B(n478), .Z(n173) );
  XNOR U46 ( .A(a[13]), .B(n469), .Z(n96) );
  XNOR U47 ( .A(a[16]), .B(n460), .Z(n93) );
  XNOR U48 ( .A(a[19]), .B(n451), .Z(n90) );
  XNOR U49 ( .A(a[22]), .B(n442), .Z(n86) );
  XNOR U50 ( .A(a[25]), .B(n433), .Z(n83) );
  XNOR U51 ( .A(a[28]), .B(n424), .Z(n80) );
  XNOR U52 ( .A(a[31]), .B(n415), .Z(n76) );
  XNOR U53 ( .A(a[34]), .B(n406), .Z(n73) );
  XNOR U54 ( .A(a[37]), .B(n397), .Z(n70) );
  XNOR U55 ( .A(a[40]), .B(n388), .Z(n66) );
  XNOR U56 ( .A(a[43]), .B(n379), .Z(n63) );
  XNOR U57 ( .A(a[46]), .B(n370), .Z(n60) );
  XNOR U58 ( .A(a[49]), .B(n361), .Z(n57) );
  XNOR U59 ( .A(a[52]), .B(n352), .Z(n53) );
  XNOR U60 ( .A(a[55]), .B(n343), .Z(n50) );
  XNOR U61 ( .A(a[58]), .B(n334), .Z(n47) );
  XNOR U62 ( .A(a[61]), .B(n325), .Z(n43) );
  XNOR U63 ( .A(a[64]), .B(n316), .Z(n40) );
  XNOR U64 ( .A(a[67]), .B(n307), .Z(n37) );
  XNOR U65 ( .A(a[70]), .B(n298), .Z(n33) );
  XNOR U66 ( .A(a[73]), .B(n289), .Z(n30) );
  XNOR U67 ( .A(a[76]), .B(n280), .Z(n27) );
  XNOR U68 ( .A(a[79]), .B(n271), .Z(n24) );
  XNOR U69 ( .A(a[82]), .B(n262), .Z(n20) );
  XNOR U70 ( .A(a[85]), .B(n253), .Z(n17) );
  XNOR U71 ( .A(a[88]), .B(n244), .Z(n14) );
  XNOR U72 ( .A(a[91]), .B(n235), .Z(n10) );
  XNOR U73 ( .A(a[94]), .B(n226), .Z(n7) );
  XNOR U74 ( .A(a[97]), .B(n217), .Z(n4) );
  XNOR U75 ( .A(a[100]), .B(n207), .Z(n209) );
  XNOR U76 ( .A(a[103]), .B(n195), .Z(n197) );
  XNOR U77 ( .A(a[106]), .B(n183), .Z(n185) );
  XNOR U78 ( .A(a[109]), .B(n170), .Z(n172) );
  XNOR U79 ( .A(a[112]), .B(n158), .Z(n160) );
  XNOR U80 ( .A(a[115]), .B(n146), .Z(n148) );
  XNOR U81 ( .A(a[118]), .B(n134), .Z(n136) );
  XNOR U82 ( .A(a[121]), .B(n121), .Z(n123) );
  XNOR U83 ( .A(a[124]), .B(n109), .Z(n111) );
  XNOR U84 ( .A(a[2]), .B(n502), .Z(n78) );
  XNOR U85 ( .A(a[5]), .B(n493), .Z(n45) );
  XNOR U86 ( .A(a[8]), .B(n484), .Z(n12) );
  XNOR U87 ( .A(a[11]), .B(n475), .Z(n132) );
  XNOR U88 ( .A(a[14]), .B(n466), .Z(n95) );
  XNOR U89 ( .A(a[17]), .B(n457), .Z(n92) );
  XNOR U90 ( .A(a[20]), .B(n448), .Z(n88) );
  XNOR U91 ( .A(a[23]), .B(n439), .Z(n85) );
  XNOR U92 ( .A(a[26]), .B(n430), .Z(n82) );
  XNOR U93 ( .A(a[29]), .B(n421), .Z(n79) );
  XNOR U94 ( .A(a[32]), .B(n412), .Z(n75) );
  XNOR U95 ( .A(a[35]), .B(n403), .Z(n72) );
  XNOR U96 ( .A(a[38]), .B(n394), .Z(n69) );
  XNOR U97 ( .A(a[41]), .B(n385), .Z(n65) );
  XNOR U98 ( .A(a[44]), .B(n376), .Z(n62) );
  XNOR U99 ( .A(a[47]), .B(n367), .Z(n59) );
  XNOR U100 ( .A(a[50]), .B(n358), .Z(n55) );
  XNOR U101 ( .A(a[53]), .B(n349), .Z(n52) );
  XNOR U102 ( .A(a[56]), .B(n340), .Z(n49) );
  XNOR U103 ( .A(a[59]), .B(n331), .Z(n46) );
  XNOR U104 ( .A(a[62]), .B(n322), .Z(n42) );
  XNOR U105 ( .A(a[65]), .B(n313), .Z(n39) );
  XNOR U106 ( .A(a[68]), .B(n304), .Z(n36) );
  XNOR U107 ( .A(a[71]), .B(n295), .Z(n32) );
  XNOR U108 ( .A(a[74]), .B(n286), .Z(n29) );
  XNOR U109 ( .A(a[77]), .B(n277), .Z(n26) );
  XNOR U110 ( .A(a[80]), .B(n268), .Z(n22) );
  XNOR U111 ( .A(a[83]), .B(n259), .Z(n19) );
  XNOR U112 ( .A(a[86]), .B(n250), .Z(n16) );
  XNOR U113 ( .A(a[89]), .B(n241), .Z(n13) );
  XNOR U114 ( .A(a[92]), .B(n232), .Z(n9) );
  XNOR U115 ( .A(a[95]), .B(n223), .Z(n6) );
  XNOR U116 ( .A(a[98]), .B(n214), .Z(n3) );
  XNOR U117 ( .A(a[101]), .B(n203), .Z(n205) );
  XNOR U118 ( .A(a[104]), .B(n191), .Z(n193) );
  XNOR U119 ( .A(a[107]), .B(n179), .Z(n181) );
  XNOR U120 ( .A(a[110]), .B(n166), .Z(n168) );
  XNOR U121 ( .A(a[113]), .B(n154), .Z(n156) );
  XNOR U122 ( .A(a[116]), .B(n142), .Z(n144) );
  XNOR U123 ( .A(a[119]), .B(n129), .Z(n131) );
  XNOR U124 ( .A(a[122]), .B(n117), .Z(n119) );
  XNOR U125 ( .A(a[125]), .B(n105), .Z(n107) );
  XNOR U126 ( .A(b[9]), .B(n1), .Z(c[9]) );
  XNOR U127 ( .A(b[99]), .B(n2), .Z(c[99]) );
  XNOR U128 ( .A(b[98]), .B(n3), .Z(c[98]) );
  XNOR U129 ( .A(b[97]), .B(n4), .Z(c[97]) );
  XNOR U130 ( .A(b[96]), .B(n5), .Z(c[96]) );
  XNOR U131 ( .A(b[95]), .B(n6), .Z(c[95]) );
  XNOR U132 ( .A(b[94]), .B(n7), .Z(c[94]) );
  XNOR U133 ( .A(b[93]), .B(n8), .Z(c[93]) );
  XNOR U134 ( .A(b[92]), .B(n9), .Z(c[92]) );
  XNOR U135 ( .A(b[91]), .B(n10), .Z(c[91]) );
  XNOR U136 ( .A(b[90]), .B(n11), .Z(c[90]) );
  XNOR U137 ( .A(b[8]), .B(n12), .Z(c[8]) );
  XNOR U138 ( .A(b[89]), .B(n13), .Z(c[89]) );
  XNOR U139 ( .A(b[88]), .B(n14), .Z(c[88]) );
  XNOR U140 ( .A(b[87]), .B(n15), .Z(c[87]) );
  XNOR U141 ( .A(b[86]), .B(n16), .Z(c[86]) );
  XNOR U142 ( .A(b[85]), .B(n17), .Z(c[85]) );
  XNOR U143 ( .A(b[84]), .B(n18), .Z(c[84]) );
  XNOR U144 ( .A(b[83]), .B(n19), .Z(c[83]) );
  XNOR U145 ( .A(b[82]), .B(n20), .Z(c[82]) );
  XNOR U146 ( .A(b[81]), .B(n21), .Z(c[81]) );
  XNOR U147 ( .A(b[80]), .B(n22), .Z(c[80]) );
  XNOR U148 ( .A(b[7]), .B(n23), .Z(c[7]) );
  XNOR U149 ( .A(b[79]), .B(n24), .Z(c[79]) );
  XNOR U150 ( .A(b[78]), .B(n25), .Z(c[78]) );
  XNOR U151 ( .A(b[77]), .B(n26), .Z(c[77]) );
  XNOR U152 ( .A(b[76]), .B(n27), .Z(c[76]) );
  XNOR U153 ( .A(b[75]), .B(n28), .Z(c[75]) );
  XNOR U154 ( .A(b[74]), .B(n29), .Z(c[74]) );
  XNOR U155 ( .A(b[73]), .B(n30), .Z(c[73]) );
  XNOR U156 ( .A(b[72]), .B(n31), .Z(c[72]) );
  XNOR U157 ( .A(b[71]), .B(n32), .Z(c[71]) );
  XNOR U158 ( .A(b[70]), .B(n33), .Z(c[70]) );
  XNOR U159 ( .A(b[6]), .B(n34), .Z(c[6]) );
  XNOR U160 ( .A(b[69]), .B(n35), .Z(c[69]) );
  XNOR U161 ( .A(b[68]), .B(n36), .Z(c[68]) );
  XNOR U162 ( .A(b[67]), .B(n37), .Z(c[67]) );
  XNOR U163 ( .A(b[66]), .B(n38), .Z(c[66]) );
  XNOR U164 ( .A(b[65]), .B(n39), .Z(c[65]) );
  XNOR U165 ( .A(b[64]), .B(n40), .Z(c[64]) );
  XNOR U166 ( .A(b[63]), .B(n41), .Z(c[63]) );
  XNOR U167 ( .A(b[62]), .B(n42), .Z(c[62]) );
  XNOR U168 ( .A(b[61]), .B(n43), .Z(c[61]) );
  XNOR U169 ( .A(b[60]), .B(n44), .Z(c[60]) );
  XNOR U170 ( .A(b[5]), .B(n45), .Z(c[5]) );
  XNOR U171 ( .A(b[59]), .B(n46), .Z(c[59]) );
  XNOR U172 ( .A(b[58]), .B(n47), .Z(c[58]) );
  XNOR U173 ( .A(b[57]), .B(n48), .Z(c[57]) );
  XNOR U174 ( .A(b[56]), .B(n49), .Z(c[56]) );
  XNOR U175 ( .A(b[55]), .B(n50), .Z(c[55]) );
  XNOR U176 ( .A(b[54]), .B(n51), .Z(c[54]) );
  XNOR U177 ( .A(b[53]), .B(n52), .Z(c[53]) );
  XNOR U178 ( .A(b[52]), .B(n53), .Z(c[52]) );
  XNOR U179 ( .A(b[51]), .B(n54), .Z(c[51]) );
  XNOR U180 ( .A(b[50]), .B(n55), .Z(c[50]) );
  XNOR U181 ( .A(b[4]), .B(n56), .Z(c[4]) );
  XNOR U182 ( .A(b[49]), .B(n57), .Z(c[49]) );
  XNOR U183 ( .A(b[48]), .B(n58), .Z(c[48]) );
  XNOR U184 ( .A(b[47]), .B(n59), .Z(c[47]) );
  XNOR U185 ( .A(b[46]), .B(n60), .Z(c[46]) );
  XNOR U186 ( .A(b[45]), .B(n61), .Z(c[45]) );
  XNOR U187 ( .A(b[44]), .B(n62), .Z(c[44]) );
  XNOR U188 ( .A(b[43]), .B(n63), .Z(c[43]) );
  XNOR U189 ( .A(b[42]), .B(n64), .Z(c[42]) );
  XNOR U190 ( .A(b[41]), .B(n65), .Z(c[41]) );
  XNOR U191 ( .A(b[40]), .B(n66), .Z(c[40]) );
  XNOR U192 ( .A(b[3]), .B(n67), .Z(c[3]) );
  XNOR U193 ( .A(b[39]), .B(n68), .Z(c[39]) );
  XNOR U194 ( .A(b[38]), .B(n69), .Z(c[38]) );
  XNOR U195 ( .A(b[37]), .B(n70), .Z(c[37]) );
  XNOR U196 ( .A(b[36]), .B(n71), .Z(c[36]) );
  XNOR U197 ( .A(b[35]), .B(n72), .Z(c[35]) );
  XNOR U198 ( .A(b[34]), .B(n73), .Z(c[34]) );
  XNOR U199 ( .A(b[33]), .B(n74), .Z(c[33]) );
  XNOR U200 ( .A(b[32]), .B(n75), .Z(c[32]) );
  XNOR U201 ( .A(b[31]), .B(n76), .Z(c[31]) );
  XNOR U202 ( .A(b[30]), .B(n77), .Z(c[30]) );
  XNOR U203 ( .A(b[2]), .B(n78), .Z(c[2]) );
  XNOR U204 ( .A(b[29]), .B(n79), .Z(c[29]) );
  XNOR U205 ( .A(b[28]), .B(n80), .Z(c[28]) );
  XNOR U206 ( .A(b[27]), .B(n81), .Z(c[27]) );
  XNOR U207 ( .A(b[26]), .B(n82), .Z(c[26]) );
  XNOR U208 ( .A(b[25]), .B(n83), .Z(c[25]) );
  XNOR U209 ( .A(b[24]), .B(n84), .Z(c[24]) );
  XNOR U210 ( .A(b[23]), .B(n85), .Z(c[23]) );
  XNOR U211 ( .A(b[22]), .B(n86), .Z(c[22]) );
  XNOR U212 ( .A(b[21]), .B(n87), .Z(c[21]) );
  XNOR U213 ( .A(b[20]), .B(n88), .Z(c[20]) );
  XNOR U214 ( .A(b[1]), .B(n89), .Z(c[1]) );
  XNOR U215 ( .A(b[19]), .B(n90), .Z(c[19]) );
  XNOR U216 ( .A(b[18]), .B(n91), .Z(c[18]) );
  XNOR U217 ( .A(b[17]), .B(n92), .Z(c[17]) );
  XNOR U218 ( .A(b[16]), .B(n93), .Z(c[16]) );
  XNOR U219 ( .A(b[15]), .B(n94), .Z(c[15]) );
  XNOR U220 ( .A(b[14]), .B(n95), .Z(c[14]) );
  XNOR U221 ( .A(b[13]), .B(n96), .Z(c[13]) );
  XNOR U222 ( .A(b[12]), .B(n97), .Z(c[12]) );
  XOR U223 ( .A(n98), .B(n99), .Z(c[127]) );
  XOR U224 ( .A(n100), .B(n101), .Z(n99) );
  ANDN U225 ( .B(n102), .A(n103), .Z(n100) );
  XOR U226 ( .A(b[126]), .B(n101), .Z(n102) );
  XOR U227 ( .A(b[127]), .B(a[127]), .Z(n98) );
  XNOR U228 ( .A(b[126]), .B(n103), .Z(c[126]) );
  XNOR U229 ( .A(a[126]), .B(n101), .Z(n103) );
  XOR U230 ( .A(n104), .B(n105), .Z(n101) );
  ANDN U231 ( .B(n106), .A(n107), .Z(n104) );
  XOR U232 ( .A(b[125]), .B(n105), .Z(n106) );
  XNOR U233 ( .A(b[125]), .B(n107), .Z(c[125]) );
  XOR U234 ( .A(n108), .B(n109), .Z(n105) );
  ANDN U235 ( .B(n110), .A(n111), .Z(n108) );
  XOR U236 ( .A(b[124]), .B(n109), .Z(n110) );
  XNOR U237 ( .A(b[124]), .B(n111), .Z(c[124]) );
  XOR U238 ( .A(n112), .B(n113), .Z(n109) );
  ANDN U239 ( .B(n114), .A(n115), .Z(n112) );
  XOR U240 ( .A(b[123]), .B(n113), .Z(n114) );
  XNOR U241 ( .A(b[123]), .B(n115), .Z(c[123]) );
  XOR U242 ( .A(n116), .B(n117), .Z(n113) );
  ANDN U243 ( .B(n118), .A(n119), .Z(n116) );
  XOR U244 ( .A(b[122]), .B(n117), .Z(n118) );
  XNOR U245 ( .A(b[122]), .B(n119), .Z(c[122]) );
  XOR U246 ( .A(n120), .B(n121), .Z(n117) );
  ANDN U247 ( .B(n122), .A(n123), .Z(n120) );
  XOR U248 ( .A(b[121]), .B(n121), .Z(n122) );
  XNOR U249 ( .A(b[121]), .B(n123), .Z(c[121]) );
  XOR U250 ( .A(n124), .B(n125), .Z(n121) );
  ANDN U251 ( .B(n126), .A(n127), .Z(n124) );
  XOR U252 ( .A(b[120]), .B(n125), .Z(n126) );
  XNOR U253 ( .A(b[120]), .B(n127), .Z(c[120]) );
  XOR U254 ( .A(n128), .B(n129), .Z(n125) );
  ANDN U255 ( .B(n130), .A(n131), .Z(n128) );
  XOR U256 ( .A(b[119]), .B(n129), .Z(n130) );
  XNOR U257 ( .A(b[11]), .B(n132), .Z(c[11]) );
  XNOR U258 ( .A(b[119]), .B(n131), .Z(c[119]) );
  XOR U259 ( .A(n133), .B(n134), .Z(n129) );
  ANDN U260 ( .B(n135), .A(n136), .Z(n133) );
  XOR U261 ( .A(b[118]), .B(n134), .Z(n135) );
  XNOR U262 ( .A(b[118]), .B(n136), .Z(c[118]) );
  XOR U263 ( .A(n137), .B(n138), .Z(n134) );
  ANDN U264 ( .B(n139), .A(n140), .Z(n137) );
  XOR U265 ( .A(b[117]), .B(n138), .Z(n139) );
  XNOR U266 ( .A(b[117]), .B(n140), .Z(c[117]) );
  XOR U267 ( .A(n141), .B(n142), .Z(n138) );
  ANDN U268 ( .B(n143), .A(n144), .Z(n141) );
  XOR U269 ( .A(b[116]), .B(n142), .Z(n143) );
  XNOR U270 ( .A(b[116]), .B(n144), .Z(c[116]) );
  XOR U271 ( .A(n145), .B(n146), .Z(n142) );
  ANDN U272 ( .B(n147), .A(n148), .Z(n145) );
  XOR U273 ( .A(b[115]), .B(n146), .Z(n147) );
  XNOR U274 ( .A(b[115]), .B(n148), .Z(c[115]) );
  XOR U275 ( .A(n149), .B(n150), .Z(n146) );
  ANDN U276 ( .B(n151), .A(n152), .Z(n149) );
  XOR U277 ( .A(b[114]), .B(n150), .Z(n151) );
  XNOR U278 ( .A(b[114]), .B(n152), .Z(c[114]) );
  XOR U279 ( .A(n153), .B(n154), .Z(n150) );
  ANDN U280 ( .B(n155), .A(n156), .Z(n153) );
  XOR U281 ( .A(b[113]), .B(n154), .Z(n155) );
  XNOR U282 ( .A(b[113]), .B(n156), .Z(c[113]) );
  XOR U283 ( .A(n157), .B(n158), .Z(n154) );
  ANDN U284 ( .B(n159), .A(n160), .Z(n157) );
  XOR U285 ( .A(b[112]), .B(n158), .Z(n159) );
  XNOR U286 ( .A(b[112]), .B(n160), .Z(c[112]) );
  XOR U287 ( .A(n161), .B(n162), .Z(n158) );
  ANDN U288 ( .B(n163), .A(n164), .Z(n161) );
  XOR U289 ( .A(b[111]), .B(n162), .Z(n163) );
  XNOR U290 ( .A(b[111]), .B(n164), .Z(c[111]) );
  XOR U291 ( .A(n165), .B(n166), .Z(n162) );
  ANDN U292 ( .B(n167), .A(n168), .Z(n165) );
  XOR U293 ( .A(b[110]), .B(n166), .Z(n167) );
  XNOR U294 ( .A(b[110]), .B(n168), .Z(c[110]) );
  XOR U295 ( .A(n169), .B(n170), .Z(n166) );
  ANDN U296 ( .B(n171), .A(n172), .Z(n169) );
  XOR U297 ( .A(b[109]), .B(n170), .Z(n171) );
  XNOR U298 ( .A(b[10]), .B(n173), .Z(c[10]) );
  XNOR U299 ( .A(b[109]), .B(n172), .Z(c[109]) );
  XOR U300 ( .A(n174), .B(n175), .Z(n170) );
  ANDN U301 ( .B(n176), .A(n177), .Z(n174) );
  XOR U302 ( .A(b[108]), .B(n175), .Z(n176) );
  XNOR U303 ( .A(b[108]), .B(n177), .Z(c[108]) );
  XOR U304 ( .A(n178), .B(n179), .Z(n175) );
  ANDN U305 ( .B(n180), .A(n181), .Z(n178) );
  XOR U306 ( .A(b[107]), .B(n179), .Z(n180) );
  XNOR U307 ( .A(b[107]), .B(n181), .Z(c[107]) );
  XOR U308 ( .A(n182), .B(n183), .Z(n179) );
  ANDN U309 ( .B(n184), .A(n185), .Z(n182) );
  XOR U310 ( .A(b[106]), .B(n183), .Z(n184) );
  XNOR U311 ( .A(b[106]), .B(n185), .Z(c[106]) );
  XOR U312 ( .A(n186), .B(n187), .Z(n183) );
  ANDN U313 ( .B(n188), .A(n189), .Z(n186) );
  XOR U314 ( .A(b[105]), .B(n187), .Z(n188) );
  XNOR U315 ( .A(b[105]), .B(n189), .Z(c[105]) );
  XOR U316 ( .A(n190), .B(n191), .Z(n187) );
  ANDN U317 ( .B(n192), .A(n193), .Z(n190) );
  XOR U318 ( .A(b[104]), .B(n191), .Z(n192) );
  XNOR U319 ( .A(b[104]), .B(n193), .Z(c[104]) );
  XOR U320 ( .A(n194), .B(n195), .Z(n191) );
  ANDN U321 ( .B(n196), .A(n197), .Z(n194) );
  XOR U322 ( .A(b[103]), .B(n195), .Z(n196) );
  XNOR U323 ( .A(b[103]), .B(n197), .Z(c[103]) );
  XOR U324 ( .A(n198), .B(n199), .Z(n195) );
  ANDN U325 ( .B(n200), .A(n201), .Z(n198) );
  XOR U326 ( .A(b[102]), .B(n199), .Z(n200) );
  XNOR U327 ( .A(b[102]), .B(n201), .Z(c[102]) );
  XOR U328 ( .A(n202), .B(n203), .Z(n199) );
  ANDN U329 ( .B(n204), .A(n205), .Z(n202) );
  XOR U330 ( .A(b[101]), .B(n203), .Z(n204) );
  XNOR U331 ( .A(b[101]), .B(n205), .Z(c[101]) );
  XOR U332 ( .A(n206), .B(n207), .Z(n203) );
  ANDN U333 ( .B(n208), .A(n209), .Z(n206) );
  XOR U334 ( .A(b[100]), .B(n207), .Z(n208) );
  XNOR U335 ( .A(b[100]), .B(n209), .Z(c[100]) );
  XOR U336 ( .A(n210), .B(n211), .Z(n207) );
  ANDN U337 ( .B(n212), .A(n2), .Z(n210) );
  XOR U338 ( .A(b[99]), .B(n211), .Z(n212) );
  XOR U339 ( .A(n213), .B(n214), .Z(n211) );
  ANDN U340 ( .B(n215), .A(n3), .Z(n213) );
  XOR U341 ( .A(b[98]), .B(n214), .Z(n215) );
  XOR U342 ( .A(n216), .B(n217), .Z(n214) );
  ANDN U343 ( .B(n218), .A(n4), .Z(n216) );
  XOR U344 ( .A(b[97]), .B(n217), .Z(n218) );
  XOR U345 ( .A(n219), .B(n220), .Z(n217) );
  ANDN U346 ( .B(n221), .A(n5), .Z(n219) );
  XOR U347 ( .A(b[96]), .B(n220), .Z(n221) );
  XOR U348 ( .A(n222), .B(n223), .Z(n220) );
  ANDN U349 ( .B(n224), .A(n6), .Z(n222) );
  XOR U350 ( .A(b[95]), .B(n223), .Z(n224) );
  XOR U351 ( .A(n225), .B(n226), .Z(n223) );
  ANDN U352 ( .B(n227), .A(n7), .Z(n225) );
  XOR U353 ( .A(b[94]), .B(n226), .Z(n227) );
  XOR U354 ( .A(n228), .B(n229), .Z(n226) );
  ANDN U355 ( .B(n230), .A(n8), .Z(n228) );
  XOR U356 ( .A(b[93]), .B(n229), .Z(n230) );
  XOR U357 ( .A(n231), .B(n232), .Z(n229) );
  ANDN U358 ( .B(n233), .A(n9), .Z(n231) );
  XOR U359 ( .A(b[92]), .B(n232), .Z(n233) );
  XOR U360 ( .A(n234), .B(n235), .Z(n232) );
  ANDN U361 ( .B(n236), .A(n10), .Z(n234) );
  XOR U362 ( .A(b[91]), .B(n235), .Z(n236) );
  XOR U363 ( .A(n237), .B(n238), .Z(n235) );
  ANDN U364 ( .B(n239), .A(n11), .Z(n237) );
  XOR U365 ( .A(b[90]), .B(n238), .Z(n239) );
  XOR U366 ( .A(n240), .B(n241), .Z(n238) );
  ANDN U367 ( .B(n242), .A(n13), .Z(n240) );
  XOR U368 ( .A(b[89]), .B(n241), .Z(n242) );
  XOR U369 ( .A(n243), .B(n244), .Z(n241) );
  ANDN U370 ( .B(n245), .A(n14), .Z(n243) );
  XOR U371 ( .A(b[88]), .B(n244), .Z(n245) );
  XOR U372 ( .A(n246), .B(n247), .Z(n244) );
  ANDN U373 ( .B(n248), .A(n15), .Z(n246) );
  XOR U374 ( .A(b[87]), .B(n247), .Z(n248) );
  XOR U375 ( .A(n249), .B(n250), .Z(n247) );
  ANDN U376 ( .B(n251), .A(n16), .Z(n249) );
  XOR U377 ( .A(b[86]), .B(n250), .Z(n251) );
  XOR U378 ( .A(n252), .B(n253), .Z(n250) );
  ANDN U379 ( .B(n254), .A(n17), .Z(n252) );
  XOR U380 ( .A(b[85]), .B(n253), .Z(n254) );
  XOR U381 ( .A(n255), .B(n256), .Z(n253) );
  ANDN U382 ( .B(n257), .A(n18), .Z(n255) );
  XOR U383 ( .A(b[84]), .B(n256), .Z(n257) );
  XOR U384 ( .A(n258), .B(n259), .Z(n256) );
  ANDN U385 ( .B(n260), .A(n19), .Z(n258) );
  XOR U386 ( .A(b[83]), .B(n259), .Z(n260) );
  XOR U387 ( .A(n261), .B(n262), .Z(n259) );
  ANDN U388 ( .B(n263), .A(n20), .Z(n261) );
  XOR U389 ( .A(b[82]), .B(n262), .Z(n263) );
  XOR U390 ( .A(n264), .B(n265), .Z(n262) );
  ANDN U391 ( .B(n266), .A(n21), .Z(n264) );
  XOR U392 ( .A(b[81]), .B(n265), .Z(n266) );
  XOR U393 ( .A(n267), .B(n268), .Z(n265) );
  ANDN U394 ( .B(n269), .A(n22), .Z(n267) );
  XOR U395 ( .A(b[80]), .B(n268), .Z(n269) );
  XOR U396 ( .A(n270), .B(n271), .Z(n268) );
  ANDN U397 ( .B(n272), .A(n24), .Z(n270) );
  XOR U398 ( .A(b[79]), .B(n271), .Z(n272) );
  XOR U399 ( .A(n273), .B(n274), .Z(n271) );
  ANDN U400 ( .B(n275), .A(n25), .Z(n273) );
  XOR U401 ( .A(b[78]), .B(n274), .Z(n275) );
  XOR U402 ( .A(n276), .B(n277), .Z(n274) );
  ANDN U403 ( .B(n278), .A(n26), .Z(n276) );
  XOR U404 ( .A(b[77]), .B(n277), .Z(n278) );
  XOR U405 ( .A(n279), .B(n280), .Z(n277) );
  ANDN U406 ( .B(n281), .A(n27), .Z(n279) );
  XOR U407 ( .A(b[76]), .B(n280), .Z(n281) );
  XOR U408 ( .A(n282), .B(n283), .Z(n280) );
  ANDN U409 ( .B(n284), .A(n28), .Z(n282) );
  XOR U410 ( .A(b[75]), .B(n283), .Z(n284) );
  XOR U411 ( .A(n285), .B(n286), .Z(n283) );
  ANDN U412 ( .B(n287), .A(n29), .Z(n285) );
  XOR U413 ( .A(b[74]), .B(n286), .Z(n287) );
  XOR U414 ( .A(n288), .B(n289), .Z(n286) );
  ANDN U415 ( .B(n290), .A(n30), .Z(n288) );
  XOR U416 ( .A(b[73]), .B(n289), .Z(n290) );
  XOR U417 ( .A(n291), .B(n292), .Z(n289) );
  ANDN U418 ( .B(n293), .A(n31), .Z(n291) );
  XOR U419 ( .A(b[72]), .B(n292), .Z(n293) );
  XOR U420 ( .A(n294), .B(n295), .Z(n292) );
  ANDN U421 ( .B(n296), .A(n32), .Z(n294) );
  XOR U422 ( .A(b[71]), .B(n295), .Z(n296) );
  XOR U423 ( .A(n297), .B(n298), .Z(n295) );
  ANDN U424 ( .B(n299), .A(n33), .Z(n297) );
  XOR U425 ( .A(b[70]), .B(n298), .Z(n299) );
  XOR U426 ( .A(n300), .B(n301), .Z(n298) );
  ANDN U427 ( .B(n302), .A(n35), .Z(n300) );
  XOR U428 ( .A(b[69]), .B(n301), .Z(n302) );
  XOR U429 ( .A(n303), .B(n304), .Z(n301) );
  ANDN U430 ( .B(n305), .A(n36), .Z(n303) );
  XOR U431 ( .A(b[68]), .B(n304), .Z(n305) );
  XOR U432 ( .A(n306), .B(n307), .Z(n304) );
  ANDN U433 ( .B(n308), .A(n37), .Z(n306) );
  XOR U434 ( .A(b[67]), .B(n307), .Z(n308) );
  XOR U435 ( .A(n309), .B(n310), .Z(n307) );
  ANDN U436 ( .B(n311), .A(n38), .Z(n309) );
  XOR U437 ( .A(b[66]), .B(n310), .Z(n311) );
  XOR U438 ( .A(n312), .B(n313), .Z(n310) );
  ANDN U439 ( .B(n314), .A(n39), .Z(n312) );
  XOR U440 ( .A(b[65]), .B(n313), .Z(n314) );
  XOR U441 ( .A(n315), .B(n316), .Z(n313) );
  ANDN U442 ( .B(n317), .A(n40), .Z(n315) );
  XOR U443 ( .A(b[64]), .B(n316), .Z(n317) );
  XOR U444 ( .A(n318), .B(n319), .Z(n316) );
  ANDN U445 ( .B(n320), .A(n41), .Z(n318) );
  XOR U446 ( .A(b[63]), .B(n319), .Z(n320) );
  XOR U447 ( .A(n321), .B(n322), .Z(n319) );
  ANDN U448 ( .B(n323), .A(n42), .Z(n321) );
  XOR U449 ( .A(b[62]), .B(n322), .Z(n323) );
  XOR U450 ( .A(n324), .B(n325), .Z(n322) );
  ANDN U451 ( .B(n326), .A(n43), .Z(n324) );
  XOR U452 ( .A(b[61]), .B(n325), .Z(n326) );
  XOR U453 ( .A(n327), .B(n328), .Z(n325) );
  ANDN U454 ( .B(n329), .A(n44), .Z(n327) );
  XOR U455 ( .A(b[60]), .B(n328), .Z(n329) );
  XOR U456 ( .A(n330), .B(n331), .Z(n328) );
  ANDN U457 ( .B(n332), .A(n46), .Z(n330) );
  XOR U458 ( .A(b[59]), .B(n331), .Z(n332) );
  XOR U459 ( .A(n333), .B(n334), .Z(n331) );
  ANDN U460 ( .B(n335), .A(n47), .Z(n333) );
  XOR U461 ( .A(b[58]), .B(n334), .Z(n335) );
  XOR U462 ( .A(n336), .B(n337), .Z(n334) );
  ANDN U463 ( .B(n338), .A(n48), .Z(n336) );
  XOR U464 ( .A(b[57]), .B(n337), .Z(n338) );
  XOR U465 ( .A(n339), .B(n340), .Z(n337) );
  ANDN U466 ( .B(n341), .A(n49), .Z(n339) );
  XOR U467 ( .A(b[56]), .B(n340), .Z(n341) );
  XOR U468 ( .A(n342), .B(n343), .Z(n340) );
  ANDN U469 ( .B(n344), .A(n50), .Z(n342) );
  XOR U470 ( .A(b[55]), .B(n343), .Z(n344) );
  XOR U471 ( .A(n345), .B(n346), .Z(n343) );
  ANDN U472 ( .B(n347), .A(n51), .Z(n345) );
  XOR U473 ( .A(b[54]), .B(n346), .Z(n347) );
  XOR U474 ( .A(n348), .B(n349), .Z(n346) );
  ANDN U475 ( .B(n350), .A(n52), .Z(n348) );
  XOR U476 ( .A(b[53]), .B(n349), .Z(n350) );
  XOR U477 ( .A(n351), .B(n352), .Z(n349) );
  ANDN U478 ( .B(n353), .A(n53), .Z(n351) );
  XOR U479 ( .A(b[52]), .B(n352), .Z(n353) );
  XOR U480 ( .A(n354), .B(n355), .Z(n352) );
  ANDN U481 ( .B(n356), .A(n54), .Z(n354) );
  XOR U482 ( .A(b[51]), .B(n355), .Z(n356) );
  XOR U483 ( .A(n357), .B(n358), .Z(n355) );
  ANDN U484 ( .B(n359), .A(n55), .Z(n357) );
  XOR U485 ( .A(b[50]), .B(n358), .Z(n359) );
  XOR U486 ( .A(n360), .B(n361), .Z(n358) );
  ANDN U487 ( .B(n362), .A(n57), .Z(n360) );
  XOR U488 ( .A(b[49]), .B(n361), .Z(n362) );
  XOR U489 ( .A(n363), .B(n364), .Z(n361) );
  ANDN U490 ( .B(n365), .A(n58), .Z(n363) );
  XOR U491 ( .A(b[48]), .B(n364), .Z(n365) );
  XOR U492 ( .A(n366), .B(n367), .Z(n364) );
  ANDN U493 ( .B(n368), .A(n59), .Z(n366) );
  XOR U494 ( .A(b[47]), .B(n367), .Z(n368) );
  XOR U495 ( .A(n369), .B(n370), .Z(n367) );
  ANDN U496 ( .B(n371), .A(n60), .Z(n369) );
  XOR U497 ( .A(b[46]), .B(n370), .Z(n371) );
  XOR U498 ( .A(n372), .B(n373), .Z(n370) );
  ANDN U499 ( .B(n374), .A(n61), .Z(n372) );
  XOR U500 ( .A(b[45]), .B(n373), .Z(n374) );
  XOR U501 ( .A(n375), .B(n376), .Z(n373) );
  ANDN U502 ( .B(n377), .A(n62), .Z(n375) );
  XOR U503 ( .A(b[44]), .B(n376), .Z(n377) );
  XOR U504 ( .A(n378), .B(n379), .Z(n376) );
  ANDN U505 ( .B(n380), .A(n63), .Z(n378) );
  XOR U506 ( .A(b[43]), .B(n379), .Z(n380) );
  XOR U507 ( .A(n381), .B(n382), .Z(n379) );
  ANDN U508 ( .B(n383), .A(n64), .Z(n381) );
  XOR U509 ( .A(b[42]), .B(n382), .Z(n383) );
  XOR U510 ( .A(n384), .B(n385), .Z(n382) );
  ANDN U511 ( .B(n386), .A(n65), .Z(n384) );
  XOR U512 ( .A(b[41]), .B(n385), .Z(n386) );
  XOR U513 ( .A(n387), .B(n388), .Z(n385) );
  ANDN U514 ( .B(n389), .A(n66), .Z(n387) );
  XOR U515 ( .A(b[40]), .B(n388), .Z(n389) );
  XOR U516 ( .A(n390), .B(n391), .Z(n388) );
  ANDN U517 ( .B(n392), .A(n68), .Z(n390) );
  XOR U518 ( .A(b[39]), .B(n391), .Z(n392) );
  XOR U519 ( .A(n393), .B(n394), .Z(n391) );
  ANDN U520 ( .B(n395), .A(n69), .Z(n393) );
  XOR U521 ( .A(b[38]), .B(n394), .Z(n395) );
  XOR U522 ( .A(n396), .B(n397), .Z(n394) );
  ANDN U523 ( .B(n398), .A(n70), .Z(n396) );
  XOR U524 ( .A(b[37]), .B(n397), .Z(n398) );
  XOR U525 ( .A(n399), .B(n400), .Z(n397) );
  ANDN U526 ( .B(n401), .A(n71), .Z(n399) );
  XOR U527 ( .A(b[36]), .B(n400), .Z(n401) );
  XOR U528 ( .A(n402), .B(n403), .Z(n400) );
  ANDN U529 ( .B(n404), .A(n72), .Z(n402) );
  XOR U530 ( .A(b[35]), .B(n403), .Z(n404) );
  XOR U531 ( .A(n405), .B(n406), .Z(n403) );
  ANDN U532 ( .B(n407), .A(n73), .Z(n405) );
  XOR U533 ( .A(b[34]), .B(n406), .Z(n407) );
  XOR U534 ( .A(n408), .B(n409), .Z(n406) );
  ANDN U535 ( .B(n410), .A(n74), .Z(n408) );
  XOR U536 ( .A(b[33]), .B(n409), .Z(n410) );
  XOR U537 ( .A(n411), .B(n412), .Z(n409) );
  ANDN U538 ( .B(n413), .A(n75), .Z(n411) );
  XOR U539 ( .A(b[32]), .B(n412), .Z(n413) );
  XOR U540 ( .A(n414), .B(n415), .Z(n412) );
  ANDN U541 ( .B(n416), .A(n76), .Z(n414) );
  XOR U542 ( .A(b[31]), .B(n415), .Z(n416) );
  XOR U543 ( .A(n417), .B(n418), .Z(n415) );
  ANDN U544 ( .B(n419), .A(n77), .Z(n417) );
  XOR U545 ( .A(b[30]), .B(n418), .Z(n419) );
  XOR U546 ( .A(n420), .B(n421), .Z(n418) );
  ANDN U547 ( .B(n422), .A(n79), .Z(n420) );
  XOR U548 ( .A(b[29]), .B(n421), .Z(n422) );
  XOR U549 ( .A(n423), .B(n424), .Z(n421) );
  ANDN U550 ( .B(n425), .A(n80), .Z(n423) );
  XOR U551 ( .A(b[28]), .B(n424), .Z(n425) );
  XOR U552 ( .A(n426), .B(n427), .Z(n424) );
  ANDN U553 ( .B(n428), .A(n81), .Z(n426) );
  XOR U554 ( .A(b[27]), .B(n427), .Z(n428) );
  XOR U555 ( .A(n429), .B(n430), .Z(n427) );
  ANDN U556 ( .B(n431), .A(n82), .Z(n429) );
  XOR U557 ( .A(b[26]), .B(n430), .Z(n431) );
  XOR U558 ( .A(n432), .B(n433), .Z(n430) );
  ANDN U559 ( .B(n434), .A(n83), .Z(n432) );
  XOR U560 ( .A(b[25]), .B(n433), .Z(n434) );
  XOR U561 ( .A(n435), .B(n436), .Z(n433) );
  ANDN U562 ( .B(n437), .A(n84), .Z(n435) );
  XOR U563 ( .A(b[24]), .B(n436), .Z(n437) );
  XOR U564 ( .A(n438), .B(n439), .Z(n436) );
  ANDN U565 ( .B(n440), .A(n85), .Z(n438) );
  XOR U566 ( .A(b[23]), .B(n439), .Z(n440) );
  XOR U567 ( .A(n441), .B(n442), .Z(n439) );
  ANDN U568 ( .B(n443), .A(n86), .Z(n441) );
  XOR U569 ( .A(b[22]), .B(n442), .Z(n443) );
  XOR U570 ( .A(n444), .B(n445), .Z(n442) );
  ANDN U571 ( .B(n446), .A(n87), .Z(n444) );
  XOR U572 ( .A(b[21]), .B(n445), .Z(n446) );
  XOR U573 ( .A(n447), .B(n448), .Z(n445) );
  ANDN U574 ( .B(n449), .A(n88), .Z(n447) );
  XOR U575 ( .A(b[20]), .B(n448), .Z(n449) );
  XOR U576 ( .A(n450), .B(n451), .Z(n448) );
  ANDN U577 ( .B(n452), .A(n90), .Z(n450) );
  XOR U578 ( .A(b[19]), .B(n451), .Z(n452) );
  XOR U579 ( .A(n453), .B(n454), .Z(n451) );
  ANDN U580 ( .B(n455), .A(n91), .Z(n453) );
  XOR U581 ( .A(b[18]), .B(n454), .Z(n455) );
  XOR U582 ( .A(n456), .B(n457), .Z(n454) );
  ANDN U583 ( .B(n458), .A(n92), .Z(n456) );
  XOR U584 ( .A(b[17]), .B(n457), .Z(n458) );
  XOR U585 ( .A(n459), .B(n460), .Z(n457) );
  ANDN U586 ( .B(n461), .A(n93), .Z(n459) );
  XOR U587 ( .A(b[16]), .B(n460), .Z(n461) );
  XOR U588 ( .A(n462), .B(n463), .Z(n460) );
  ANDN U589 ( .B(n464), .A(n94), .Z(n462) );
  XOR U590 ( .A(b[15]), .B(n463), .Z(n464) );
  XOR U591 ( .A(n465), .B(n466), .Z(n463) );
  ANDN U592 ( .B(n467), .A(n95), .Z(n465) );
  XOR U593 ( .A(b[14]), .B(n466), .Z(n467) );
  XOR U594 ( .A(n468), .B(n469), .Z(n466) );
  ANDN U595 ( .B(n470), .A(n96), .Z(n468) );
  XOR U596 ( .A(b[13]), .B(n469), .Z(n470) );
  XOR U597 ( .A(n471), .B(n472), .Z(n469) );
  ANDN U598 ( .B(n473), .A(n97), .Z(n471) );
  XOR U599 ( .A(b[12]), .B(n472), .Z(n473) );
  XOR U600 ( .A(n474), .B(n475), .Z(n472) );
  ANDN U601 ( .B(n476), .A(n132), .Z(n474) );
  XOR U602 ( .A(b[11]), .B(n475), .Z(n476) );
  XOR U603 ( .A(n477), .B(n478), .Z(n475) );
  ANDN U604 ( .B(n479), .A(n173), .Z(n477) );
  XOR U605 ( .A(b[10]), .B(n478), .Z(n479) );
  XOR U606 ( .A(n480), .B(n481), .Z(n478) );
  ANDN U607 ( .B(n482), .A(n1), .Z(n480) );
  XOR U608 ( .A(b[9]), .B(n481), .Z(n482) );
  XOR U609 ( .A(n483), .B(n484), .Z(n481) );
  ANDN U610 ( .B(n485), .A(n12), .Z(n483) );
  XOR U611 ( .A(b[8]), .B(n484), .Z(n485) );
  XOR U612 ( .A(n486), .B(n487), .Z(n484) );
  ANDN U613 ( .B(n488), .A(n23), .Z(n486) );
  XOR U614 ( .A(b[7]), .B(n487), .Z(n488) );
  XOR U615 ( .A(n489), .B(n490), .Z(n487) );
  ANDN U616 ( .B(n491), .A(n34), .Z(n489) );
  XOR U617 ( .A(b[6]), .B(n490), .Z(n491) );
  XOR U618 ( .A(n492), .B(n493), .Z(n490) );
  ANDN U619 ( .B(n494), .A(n45), .Z(n492) );
  XOR U620 ( .A(b[5]), .B(n493), .Z(n494) );
  XOR U621 ( .A(n495), .B(n496), .Z(n493) );
  ANDN U622 ( .B(n497), .A(n56), .Z(n495) );
  XOR U623 ( .A(b[4]), .B(n496), .Z(n497) );
  XOR U624 ( .A(n498), .B(n499), .Z(n496) );
  ANDN U625 ( .B(n500), .A(n67), .Z(n498) );
  XOR U626 ( .A(b[3]), .B(n499), .Z(n500) );
  XOR U627 ( .A(n501), .B(n502), .Z(n499) );
  ANDN U628 ( .B(n503), .A(n78), .Z(n501) );
  XOR U629 ( .A(b[2]), .B(n502), .Z(n503) );
  XNOR U630 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U631 ( .A(n89), .B(n506), .Z(n505) );
  XOR U632 ( .A(b[1]), .B(n504), .Z(n506) );
  XNOR U633 ( .A(a[1]), .B(n504), .Z(n89) );
  AND U634 ( .A(b[0]), .B(a[0]), .Z(n504) );
  XOR U635 ( .A(b[0]), .B(a[0]), .Z(c[0]) );
endmodule

