
module stackMachine_N32 ( clk, rst, x, opcode, o );
  input [31:0] x;
  input [2:0] opcode;
  output [31:0] o;
  input clk, rst;
  wire   \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \stack[0][31] , \stack[0][30] , \stack[0][29] , \stack[0][28] ,
         \stack[0][27] , \stack[0][26] , \stack[0][25] , \stack[0][24] ,
         \stack[0][23] , \stack[0][22] , \stack[0][21] , \stack[0][20] ,
         \stack[0][19] , \stack[0][18] , \stack[0][17] , \stack[0][16] ,
         \stack[0][15] , \stack[0][14] , \stack[0][13] , \stack[0][12] ,
         \stack[0][11] , \stack[0][10] , \stack[0][9] , \stack[0][8] ,
         \stack[0][7] , \stack[0][6] , \stack[0][5] , \stack[0][4] ,
         \stack[0][3] , \stack[0][2] , \stack[0][1] , \stack[0][0] , n1989,
         n1996, n2003, n2012, n2021, n2030, n2039, n2048, n2057, n2066, n2075,
         n2084, n2093, n2102, n2111, n2120, n2129, n2138, n2147, n2156, n2165,
         n2174, n2183, n2192, n2201, n2210, n2219, n2228, n2237, n2246, n2255,
         n2264, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026;

  DFF \stack_reg[0][0]  ( .D(n2499), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][0] ) );
  DFF \stack_reg[1][0]  ( .D(n2467), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][0] ) );
  DFF \stack_reg[0][31]  ( .D(n2468), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][31] ) );
  DFF \stack_reg[1][31]  ( .D(n2436), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][31] ) );
  DFF \stack_reg[0][1]  ( .D(n2498), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][1] ) );
  DFF \stack_reg[1][1]  ( .D(n2466), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][1] ) );
  DFF \stack_reg[2][1]  ( .D(n2434), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][1] ) );
  DFF \stack_reg[3][1]  ( .D(n2402), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][1] ) );
  DFF \stack_reg[4][1]  ( .D(n2370), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][1] ) );
  DFF \stack_reg[5][1]  ( .D(n2338), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][1] ) );
  DFF \stack_reg[6][1]  ( .D(n2306), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][1] ) );
  DFF \stack_reg[7][1]  ( .D(n2264), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][1] ) );
  DFF \stack_reg[0][2]  ( .D(n2497), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][2] ) );
  DFF \stack_reg[1][2]  ( .D(n2465), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][2] ) );
  DFF \stack_reg[2][2]  ( .D(n2433), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][2] ) );
  DFF \stack_reg[3][2]  ( .D(n2401), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][2] ) );
  DFF \stack_reg[4][2]  ( .D(n2369), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][2] ) );
  DFF \stack_reg[5][2]  ( .D(n2337), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][2] ) );
  DFF \stack_reg[6][2]  ( .D(n2305), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][2] ) );
  DFF \stack_reg[7][2]  ( .D(n2255), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][2] ) );
  DFF \stack_reg[0][3]  ( .D(n2496), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][3] ) );
  DFF \stack_reg[1][3]  ( .D(n2464), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][3] ) );
  DFF \stack_reg[2][3]  ( .D(n2432), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][3] ) );
  DFF \stack_reg[3][3]  ( .D(n2400), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][3] ) );
  DFF \stack_reg[4][3]  ( .D(n2368), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][3] ) );
  DFF \stack_reg[5][3]  ( .D(n2336), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][3] ) );
  DFF \stack_reg[6][3]  ( .D(n2304), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][3] ) );
  DFF \stack_reg[7][3]  ( .D(n2246), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][3] ) );
  DFF \stack_reg[0][4]  ( .D(n2495), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][4] ) );
  DFF \stack_reg[1][4]  ( .D(n2463), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][4] ) );
  DFF \stack_reg[2][4]  ( .D(n2431), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][4] ) );
  DFF \stack_reg[3][4]  ( .D(n2399), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][4] ) );
  DFF \stack_reg[4][4]  ( .D(n2367), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][4] ) );
  DFF \stack_reg[5][4]  ( .D(n2335), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][4] ) );
  DFF \stack_reg[6][4]  ( .D(n2303), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][4] ) );
  DFF \stack_reg[7][4]  ( .D(n2237), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][4] ) );
  DFF \stack_reg[0][5]  ( .D(n2494), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][5] ) );
  DFF \stack_reg[1][5]  ( .D(n2462), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][5] ) );
  DFF \stack_reg[2][5]  ( .D(n2430), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][5] ) );
  DFF \stack_reg[3][5]  ( .D(n2398), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][5] ) );
  DFF \stack_reg[4][5]  ( .D(n2366), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][5] ) );
  DFF \stack_reg[5][5]  ( .D(n2334), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][5] ) );
  DFF \stack_reg[6][5]  ( .D(n2302), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][5] ) );
  DFF \stack_reg[7][5]  ( .D(n2228), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][5] ) );
  DFF \stack_reg[0][6]  ( .D(n2493), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][6] ) );
  DFF \stack_reg[1][6]  ( .D(n2461), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][6] ) );
  DFF \stack_reg[2][6]  ( .D(n2429), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][6] ) );
  DFF \stack_reg[3][6]  ( .D(n2397), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][6] ) );
  DFF \stack_reg[4][6]  ( .D(n2365), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][6] ) );
  DFF \stack_reg[5][6]  ( .D(n2333), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][6] ) );
  DFF \stack_reg[6][6]  ( .D(n2301), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][6] ) );
  DFF \stack_reg[7][6]  ( .D(n2219), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][6] ) );
  DFF \stack_reg[0][7]  ( .D(n2492), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][7] ) );
  DFF \stack_reg[1][7]  ( .D(n2460), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][7] ) );
  DFF \stack_reg[2][7]  ( .D(n2428), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][7] ) );
  DFF \stack_reg[3][7]  ( .D(n2396), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][7] ) );
  DFF \stack_reg[4][7]  ( .D(n2364), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][7] ) );
  DFF \stack_reg[5][7]  ( .D(n2332), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][7] ) );
  DFF \stack_reg[6][7]  ( .D(n2300), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][7] ) );
  DFF \stack_reg[7][7]  ( .D(n2210), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][7] ) );
  DFF \stack_reg[0][8]  ( .D(n2491), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][8] ) );
  DFF \stack_reg[1][8]  ( .D(n2459), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][8] ) );
  DFF \stack_reg[2][8]  ( .D(n2427), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][8] ) );
  DFF \stack_reg[3][8]  ( .D(n2395), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][8] ) );
  DFF \stack_reg[4][8]  ( .D(n2363), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][8] ) );
  DFF \stack_reg[5][8]  ( .D(n2331), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][8] ) );
  DFF \stack_reg[6][8]  ( .D(n2299), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][8] ) );
  DFF \stack_reg[7][8]  ( .D(n2201), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][8] ) );
  DFF \stack_reg[0][9]  ( .D(n2490), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][9] ) );
  DFF \stack_reg[1][9]  ( .D(n2458), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][9] ) );
  DFF \stack_reg[2][9]  ( .D(n2426), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][9] ) );
  DFF \stack_reg[3][9]  ( .D(n2394), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][9] ) );
  DFF \stack_reg[4][9]  ( .D(n2362), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][9] ) );
  DFF \stack_reg[5][9]  ( .D(n2330), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][9] ) );
  DFF \stack_reg[6][9]  ( .D(n2298), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][9] ) );
  DFF \stack_reg[7][9]  ( .D(n2192), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][9] ) );
  DFF \stack_reg[0][10]  ( .D(n2489), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][10] ) );
  DFF \stack_reg[1][10]  ( .D(n2457), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][10] ) );
  DFF \stack_reg[2][10]  ( .D(n2425), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][10] ) );
  DFF \stack_reg[3][10]  ( .D(n2393), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][10] ) );
  DFF \stack_reg[4][10]  ( .D(n2361), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][10] ) );
  DFF \stack_reg[5][10]  ( .D(n2329), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][10] ) );
  DFF \stack_reg[6][10]  ( .D(n2297), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][10] ) );
  DFF \stack_reg[7][10]  ( .D(n2183), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][10] ) );
  DFF \stack_reg[0][11]  ( .D(n2488), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][11] ) );
  DFF \stack_reg[1][11]  ( .D(n2456), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][11] ) );
  DFF \stack_reg[2][11]  ( .D(n2424), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][11] ) );
  DFF \stack_reg[3][11]  ( .D(n2392), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][11] ) );
  DFF \stack_reg[4][11]  ( .D(n2360), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][11] ) );
  DFF \stack_reg[5][11]  ( .D(n2328), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][11] ) );
  DFF \stack_reg[6][11]  ( .D(n2296), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][11] ) );
  DFF \stack_reg[7][11]  ( .D(n2174), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][11] ) );
  DFF \stack_reg[0][12]  ( .D(n2487), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][12] ) );
  DFF \stack_reg[1][12]  ( .D(n2455), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][12] ) );
  DFF \stack_reg[2][12]  ( .D(n2423), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][12] ) );
  DFF \stack_reg[3][12]  ( .D(n2391), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][12] ) );
  DFF \stack_reg[4][12]  ( .D(n2359), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][12] ) );
  DFF \stack_reg[5][12]  ( .D(n2327), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][12] ) );
  DFF \stack_reg[6][12]  ( .D(n2295), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][12] ) );
  DFF \stack_reg[7][12]  ( .D(n2165), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][12] ) );
  DFF \stack_reg[0][13]  ( .D(n2486), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][13] ) );
  DFF \stack_reg[1][13]  ( .D(n2454), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][13] ) );
  DFF \stack_reg[2][13]  ( .D(n2422), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][13] ) );
  DFF \stack_reg[3][13]  ( .D(n2390), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][13] ) );
  DFF \stack_reg[4][13]  ( .D(n2358), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][13] ) );
  DFF \stack_reg[5][13]  ( .D(n2326), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][13] ) );
  DFF \stack_reg[6][13]  ( .D(n2294), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][13] ) );
  DFF \stack_reg[7][13]  ( .D(n2156), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][13] ) );
  DFF \stack_reg[0][14]  ( .D(n2485), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][14] ) );
  DFF \stack_reg[1][14]  ( .D(n2453), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][14] ) );
  DFF \stack_reg[2][14]  ( .D(n2421), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][14] ) );
  DFF \stack_reg[3][14]  ( .D(n2389), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][14] ) );
  DFF \stack_reg[4][14]  ( .D(n2357), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][14] ) );
  DFF \stack_reg[5][14]  ( .D(n2325), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][14] ) );
  DFF \stack_reg[6][14]  ( .D(n2293), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][14] ) );
  DFF \stack_reg[7][14]  ( .D(n2147), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][14] ) );
  DFF \stack_reg[0][15]  ( .D(n2484), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][15] ) );
  DFF \stack_reg[1][15]  ( .D(n2452), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][15] ) );
  DFF \stack_reg[2][15]  ( .D(n2420), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][15] ) );
  DFF \stack_reg[3][15]  ( .D(n2388), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][15] ) );
  DFF \stack_reg[4][15]  ( .D(n2356), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][15] ) );
  DFF \stack_reg[5][15]  ( .D(n2324), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][15] ) );
  DFF \stack_reg[6][15]  ( .D(n2292), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][15] ) );
  DFF \stack_reg[7][15]  ( .D(n2138), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][15] ) );
  DFF \stack_reg[0][16]  ( .D(n2483), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][16] ) );
  DFF \stack_reg[1][16]  ( .D(n2451), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][16] ) );
  DFF \stack_reg[2][16]  ( .D(n2419), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][16] ) );
  DFF \stack_reg[3][16]  ( .D(n2387), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][16] ) );
  DFF \stack_reg[4][16]  ( .D(n2355), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][16] ) );
  DFF \stack_reg[5][16]  ( .D(n2323), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][16] ) );
  DFF \stack_reg[6][16]  ( .D(n2291), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][16] ) );
  DFF \stack_reg[7][16]  ( .D(n2129), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][16] ) );
  DFF \stack_reg[0][17]  ( .D(n2482), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][17] ) );
  DFF \stack_reg[1][17]  ( .D(n2450), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][17] ) );
  DFF \stack_reg[2][17]  ( .D(n2418), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][17] ) );
  DFF \stack_reg[3][17]  ( .D(n2386), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][17] ) );
  DFF \stack_reg[4][17]  ( .D(n2354), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][17] ) );
  DFF \stack_reg[5][17]  ( .D(n2322), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][17] ) );
  DFF \stack_reg[6][17]  ( .D(n2290), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][17] ) );
  DFF \stack_reg[7][17]  ( .D(n2120), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][17] ) );
  DFF \stack_reg[0][18]  ( .D(n2481), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][18] ) );
  DFF \stack_reg[1][18]  ( .D(n2449), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][18] ) );
  DFF \stack_reg[2][18]  ( .D(n2417), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][18] ) );
  DFF \stack_reg[3][18]  ( .D(n2385), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][18] ) );
  DFF \stack_reg[4][18]  ( .D(n2353), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][18] ) );
  DFF \stack_reg[5][18]  ( .D(n2321), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][18] ) );
  DFF \stack_reg[6][18]  ( .D(n2289), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][18] ) );
  DFF \stack_reg[7][18]  ( .D(n2111), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][18] ) );
  DFF \stack_reg[0][19]  ( .D(n2480), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][19] ) );
  DFF \stack_reg[1][19]  ( .D(n2448), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][19] ) );
  DFF \stack_reg[2][19]  ( .D(n2416), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][19] ) );
  DFF \stack_reg[3][19]  ( .D(n2384), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][19] ) );
  DFF \stack_reg[4][19]  ( .D(n2352), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][19] ) );
  DFF \stack_reg[5][19]  ( .D(n2320), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][19] ) );
  DFF \stack_reg[6][19]  ( .D(n2288), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][19] ) );
  DFF \stack_reg[7][19]  ( .D(n2102), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][19] ) );
  DFF \stack_reg[0][20]  ( .D(n2479), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][20] ) );
  DFF \stack_reg[1][20]  ( .D(n2447), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][20] ) );
  DFF \stack_reg[2][20]  ( .D(n2415), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][20] ) );
  DFF \stack_reg[3][20]  ( .D(n2383), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][20] ) );
  DFF \stack_reg[4][20]  ( .D(n2351), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][20] ) );
  DFF \stack_reg[5][20]  ( .D(n2319), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][20] ) );
  DFF \stack_reg[6][20]  ( .D(n2287), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][20] ) );
  DFF \stack_reg[7][20]  ( .D(n2093), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][20] ) );
  DFF \stack_reg[0][21]  ( .D(n2478), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][21] ) );
  DFF \stack_reg[1][21]  ( .D(n2446), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][21] ) );
  DFF \stack_reg[2][21]  ( .D(n2414), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][21] ) );
  DFF \stack_reg[3][21]  ( .D(n2382), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][21] ) );
  DFF \stack_reg[4][21]  ( .D(n2350), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][21] ) );
  DFF \stack_reg[5][21]  ( .D(n2318), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][21] ) );
  DFF \stack_reg[6][21]  ( .D(n2286), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][21] ) );
  DFF \stack_reg[7][21]  ( .D(n2084), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][21] ) );
  DFF \stack_reg[0][22]  ( .D(n2477), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][22] ) );
  DFF \stack_reg[1][22]  ( .D(n2445), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][22] ) );
  DFF \stack_reg[2][22]  ( .D(n2413), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][22] ) );
  DFF \stack_reg[3][22]  ( .D(n2381), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][22] ) );
  DFF \stack_reg[4][22]  ( .D(n2349), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][22] ) );
  DFF \stack_reg[5][22]  ( .D(n2317), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][22] ) );
  DFF \stack_reg[6][22]  ( .D(n2285), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][22] ) );
  DFF \stack_reg[7][22]  ( .D(n2075), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][22] ) );
  DFF \stack_reg[0][23]  ( .D(n2476), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][23] ) );
  DFF \stack_reg[1][23]  ( .D(n2444), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][23] ) );
  DFF \stack_reg[2][23]  ( .D(n2412), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][23] ) );
  DFF \stack_reg[3][23]  ( .D(n2380), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][23] ) );
  DFF \stack_reg[4][23]  ( .D(n2348), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][23] ) );
  DFF \stack_reg[5][23]  ( .D(n2316), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][23] ) );
  DFF \stack_reg[6][23]  ( .D(n2284), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][23] ) );
  DFF \stack_reg[7][23]  ( .D(n2066), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][23] ) );
  DFF \stack_reg[0][24]  ( .D(n2475), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][24] ) );
  DFF \stack_reg[1][24]  ( .D(n2443), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][24] ) );
  DFF \stack_reg[2][24]  ( .D(n2411), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][24] ) );
  DFF \stack_reg[3][24]  ( .D(n2379), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][24] ) );
  DFF \stack_reg[4][24]  ( .D(n2347), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][24] ) );
  DFF \stack_reg[5][24]  ( .D(n2315), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][24] ) );
  DFF \stack_reg[6][24]  ( .D(n2283), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][24] ) );
  DFF \stack_reg[7][24]  ( .D(n2057), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][24] ) );
  DFF \stack_reg[0][25]  ( .D(n2474), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][25] ) );
  DFF \stack_reg[1][25]  ( .D(n2442), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][25] ) );
  DFF \stack_reg[2][25]  ( .D(n2410), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][25] ) );
  DFF \stack_reg[3][25]  ( .D(n2378), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][25] ) );
  DFF \stack_reg[4][25]  ( .D(n2346), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][25] ) );
  DFF \stack_reg[5][25]  ( .D(n2314), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][25] ) );
  DFF \stack_reg[6][25]  ( .D(n2282), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][25] ) );
  DFF \stack_reg[7][25]  ( .D(n2048), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][25] ) );
  DFF \stack_reg[0][26]  ( .D(n2473), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][26] ) );
  DFF \stack_reg[1][26]  ( .D(n2441), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][26] ) );
  DFF \stack_reg[2][26]  ( .D(n2409), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][26] ) );
  DFF \stack_reg[3][26]  ( .D(n2377), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][26] ) );
  DFF \stack_reg[4][26]  ( .D(n2345), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][26] ) );
  DFF \stack_reg[5][26]  ( .D(n2313), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][26] ) );
  DFF \stack_reg[6][26]  ( .D(n2281), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][26] ) );
  DFF \stack_reg[7][26]  ( .D(n2039), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][26] ) );
  DFF \stack_reg[0][27]  ( .D(n2472), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][27] ) );
  DFF \stack_reg[1][27]  ( .D(n2440), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][27] ) );
  DFF \stack_reg[2][27]  ( .D(n2408), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][27] ) );
  DFF \stack_reg[3][27]  ( .D(n2376), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][27] ) );
  DFF \stack_reg[4][27]  ( .D(n2344), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][27] ) );
  DFF \stack_reg[5][27]  ( .D(n2312), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][27] ) );
  DFF \stack_reg[6][27]  ( .D(n2280), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][27] ) );
  DFF \stack_reg[7][27]  ( .D(n2030), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][27] ) );
  DFF \stack_reg[0][28]  ( .D(n2471), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][28] ) );
  DFF \stack_reg[1][28]  ( .D(n2439), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][28] ) );
  DFF \stack_reg[2][28]  ( .D(n2407), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][28] ) );
  DFF \stack_reg[3][28]  ( .D(n2375), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][28] ) );
  DFF \stack_reg[4][28]  ( .D(n2343), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][28] ) );
  DFF \stack_reg[5][28]  ( .D(n2311), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][28] ) );
  DFF \stack_reg[6][28]  ( .D(n2279), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][28] ) );
  DFF \stack_reg[7][28]  ( .D(n2021), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][28] ) );
  DFF \stack_reg[0][29]  ( .D(n2470), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][29] ) );
  DFF \stack_reg[1][29]  ( .D(n2438), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][29] ) );
  DFF \stack_reg[2][29]  ( .D(n2406), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][29] ) );
  DFF \stack_reg[3][29]  ( .D(n2374), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][29] ) );
  DFF \stack_reg[4][29]  ( .D(n2342), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][29] ) );
  DFF \stack_reg[5][29]  ( .D(n2310), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][29] ) );
  DFF \stack_reg[6][29]  ( .D(n2278), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][29] ) );
  DFF \stack_reg[7][29]  ( .D(n2012), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][29] ) );
  DFF \stack_reg[0][30]  ( .D(n2469), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][30] ) );
  DFF \stack_reg[1][30]  ( .D(n2437), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][30] ) );
  DFF \stack_reg[2][30]  ( .D(n2405), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][30] ) );
  DFF \stack_reg[3][30]  ( .D(n2373), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][30] ) );
  DFF \stack_reg[4][30]  ( .D(n2341), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][30] ) );
  DFF \stack_reg[5][30]  ( .D(n2309), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][30] ) );
  DFF \stack_reg[6][30]  ( .D(n2277), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][30] ) );
  DFF \stack_reg[7][30]  ( .D(n2003), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][30] ) );
  DFF \stack_reg[2][31]  ( .D(n2404), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][31] ) );
  DFF \stack_reg[3][31]  ( .D(n2372), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][31] ) );
  DFF \stack_reg[4][31]  ( .D(n2340), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][31] ) );
  DFF \stack_reg[5][31]  ( .D(n2308), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][31] ) );
  DFF \stack_reg[6][31]  ( .D(n2276), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][31] ) );
  DFF \stack_reg[7][31]  ( .D(n1996), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][31] ) );
  DFF \stack_reg[2][0]  ( .D(n2435), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][0] ) );
  DFF \stack_reg[3][0]  ( .D(n2403), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][0] ) );
  DFF \stack_reg[4][0]  ( .D(n2371), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][0] ) );
  DFF \stack_reg[5][0]  ( .D(n2339), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][0] ) );
  DFF \stack_reg[6][0]  ( .D(n2307), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][0] ) );
  DFF \stack_reg[7][0]  ( .D(n1989), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][0] ) );
  OR U2528 ( .A(n3366), .B(n3365), .Z(n3368) );
  OR U2529 ( .A(n4003), .B(n4005), .Z(n4203) );
  OR U2530 ( .A(n3458), .B(n3457), .Z(n3460) );
  OR U2531 ( .A(n3492), .B(n3491), .Z(n3494) );
  NANDN U2532 ( .A(n3636), .B(n3635), .Z(n3638) );
  AND U2533 ( .A(\stack[1][0] ), .B(\stack[0][30] ), .Z(n3323) );
  NANDN U2534 ( .A(n2831), .B(n2833), .Z(n6772) );
  XNOR U2535 ( .A(\stack[1][31] ), .B(\stack[0][31] ), .Z(n3349) );
  OR U2536 ( .A(n3472), .B(n3471), .Z(n3474) );
  OR U2537 ( .A(n3434), .B(n3433), .Z(n3436) );
  OR U2538 ( .A(n3422), .B(n3421), .Z(n3424) );
  OR U2539 ( .A(n3518), .B(n3517), .Z(n3520) );
  OR U2540 ( .A(n3408), .B(n3407), .Z(n3410) );
  OR U2541 ( .A(n3544), .B(n3543), .Z(n3546) );
  OR U2542 ( .A(n4763), .B(n4765), .Z(n4933) );
  OR U2543 ( .A(n3394), .B(n3393), .Z(n3396) );
  OR U2544 ( .A(n3570), .B(n3569), .Z(n3572) );
  OR U2545 ( .A(n3380), .B(n3379), .Z(n3382) );
  OR U2546 ( .A(n4398), .B(n4400), .Z(n4583) );
  OR U2547 ( .A(n3596), .B(n3595), .Z(n3598) );
  OR U2548 ( .A(n3622), .B(n3621), .Z(n3624) );
  NANDN U2549 ( .A(n2819), .B(n2821), .Z(n3714) );
  NANDN U2550 ( .A(n2619), .B(n2621), .Z(n6807) );
  OR U2551 ( .A(\stack[0][30] ), .B(\stack[1][30] ), .Z(n3328) );
  OR U2552 ( .A(\stack[0][29] ), .B(\stack[1][29] ), .Z(n3305) );
  OR U2553 ( .A(\stack[0][28] ), .B(\stack[1][28] ), .Z(n3282) );
  NANDN U2554 ( .A(\stack[0][2] ), .B(n2660), .Z(n2659) );
  OR U2555 ( .A(\stack[0][31] ), .B(\stack[1][31] ), .Z(n6668) );
  NANDN U2556 ( .A(n2500), .B(n2501), .Z(o[9]) );
  NANDN U2557 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2558 ( .A(n2504), .B(n2505), .Z(o[8]) );
  NANDN U2559 ( .A(n2506), .B(n2503), .Z(n2505) );
  NANDN U2560 ( .A(n2507), .B(n2508), .Z(o[7]) );
  NANDN U2561 ( .A(n2509), .B(n2503), .Z(n2508) );
  NANDN U2562 ( .A(n2510), .B(n2511), .Z(o[6]) );
  NANDN U2563 ( .A(n2512), .B(n2503), .Z(n2511) );
  NANDN U2564 ( .A(n2513), .B(n2514), .Z(o[5]) );
  NANDN U2565 ( .A(n2515), .B(n2503), .Z(n2514) );
  NANDN U2566 ( .A(n2516), .B(n2517), .Z(o[4]) );
  NANDN U2567 ( .A(n2518), .B(n2503), .Z(n2517) );
  NANDN U2568 ( .A(n2519), .B(n2520), .Z(o[3]) );
  NANDN U2569 ( .A(n2521), .B(n2503), .Z(n2520) );
  NANDN U2570 ( .A(n2522), .B(n2523), .Z(o[31]) );
  NANDN U2571 ( .A(n2524), .B(n2503), .Z(n2523) );
  NANDN U2572 ( .A(n2525), .B(n2526), .Z(o[30]) );
  NANDN U2573 ( .A(n2527), .B(n2503), .Z(n2526) );
  NANDN U2574 ( .A(n2528), .B(n2529), .Z(o[2]) );
  NANDN U2575 ( .A(n2530), .B(n2503), .Z(n2529) );
  NANDN U2576 ( .A(n2531), .B(n2532), .Z(o[29]) );
  NANDN U2577 ( .A(n2533), .B(n2503), .Z(n2532) );
  NANDN U2578 ( .A(n2534), .B(n2535), .Z(o[28]) );
  NANDN U2579 ( .A(n2536), .B(n2503), .Z(n2535) );
  NANDN U2580 ( .A(n2537), .B(n2538), .Z(o[27]) );
  NANDN U2581 ( .A(n2539), .B(n2503), .Z(n2538) );
  NANDN U2582 ( .A(n2540), .B(n2541), .Z(o[26]) );
  NANDN U2583 ( .A(n2542), .B(n2503), .Z(n2541) );
  NANDN U2584 ( .A(n2543), .B(n2544), .Z(o[25]) );
  NANDN U2585 ( .A(n2545), .B(n2503), .Z(n2544) );
  NANDN U2586 ( .A(n2546), .B(n2547), .Z(o[24]) );
  NANDN U2587 ( .A(n2548), .B(n2503), .Z(n2547) );
  NANDN U2588 ( .A(n2549), .B(n2550), .Z(o[23]) );
  NANDN U2589 ( .A(n2551), .B(n2503), .Z(n2550) );
  NANDN U2590 ( .A(n2552), .B(n2553), .Z(o[22]) );
  NANDN U2591 ( .A(n2554), .B(n2503), .Z(n2553) );
  NANDN U2592 ( .A(n2555), .B(n2556), .Z(o[21]) );
  NANDN U2593 ( .A(n2557), .B(n2503), .Z(n2556) );
  NANDN U2594 ( .A(n2558), .B(n2559), .Z(o[20]) );
  NANDN U2595 ( .A(n2560), .B(n2503), .Z(n2559) );
  NANDN U2596 ( .A(n2561), .B(n2562), .Z(o[1]) );
  NANDN U2597 ( .A(n2563), .B(n2503), .Z(n2562) );
  NANDN U2598 ( .A(n2564), .B(n2565), .Z(o[19]) );
  NANDN U2599 ( .A(n2566), .B(n2503), .Z(n2565) );
  NANDN U2600 ( .A(n2567), .B(n2568), .Z(o[18]) );
  NANDN U2601 ( .A(n2569), .B(n2503), .Z(n2568) );
  NANDN U2602 ( .A(n2570), .B(n2571), .Z(o[17]) );
  NANDN U2603 ( .A(n2572), .B(n2503), .Z(n2571) );
  NANDN U2604 ( .A(n2573), .B(n2574), .Z(o[16]) );
  NANDN U2605 ( .A(n2575), .B(n2503), .Z(n2574) );
  NANDN U2606 ( .A(n2576), .B(n2577), .Z(o[15]) );
  NANDN U2607 ( .A(n2578), .B(n2503), .Z(n2577) );
  NANDN U2608 ( .A(n2579), .B(n2580), .Z(o[14]) );
  NANDN U2609 ( .A(n2581), .B(n2503), .Z(n2580) );
  NANDN U2610 ( .A(n2582), .B(n2583), .Z(o[13]) );
  NANDN U2611 ( .A(n2584), .B(n2503), .Z(n2583) );
  NANDN U2612 ( .A(n2585), .B(n2586), .Z(o[12]) );
  NANDN U2613 ( .A(n2587), .B(n2503), .Z(n2586) );
  NANDN U2614 ( .A(n2588), .B(n2589), .Z(o[11]) );
  NANDN U2615 ( .A(n2590), .B(n2503), .Z(n2589) );
  NANDN U2616 ( .A(n2591), .B(n2592), .Z(o[10]) );
  NANDN U2617 ( .A(n2593), .B(n2503), .Z(n2592) );
  NANDN U2618 ( .A(n2594), .B(n2595), .Z(o[0]) );
  NANDN U2619 ( .A(n2596), .B(n2503), .Z(n2595) );
  NAND U2620 ( .A(n2597), .B(n2598), .Z(n2499) );
  NANDN U2621 ( .A(n2599), .B(\stack[0][0] ), .Z(n2598) );
  ANDN U2622 ( .B(n2600), .A(n2594), .Z(n2597) );
  ANDN U2623 ( .B(x[0]), .A(n2503), .Z(n2594) );
  NANDN U2624 ( .A(n2596), .B(n2601), .Z(n2600) );
  AND U2625 ( .A(n2602), .B(n2603), .Z(n2596) );
  AND U2626 ( .A(n2604), .B(n2605), .Z(n2603) );
  NAND U2627 ( .A(n2606), .B(n2607), .Z(n2605) );
  AND U2628 ( .A(\stack[0][0] ), .B(\stack[1][0] ), .Z(n2606) );
  AND U2629 ( .A(n2608), .B(n2609), .Z(n2604) );
  NAND U2630 ( .A(\stack[1][0] ), .B(n2610), .Z(n2609) );
  ANDN U2631 ( .B(\stack[0][0] ), .A(n2611), .Z(n2610) );
  NAND U2632 ( .A(n2612), .B(n2613), .Z(n2608) );
  NAND U2633 ( .A(n2614), .B(n2615), .Z(n2612) );
  AND U2634 ( .A(n2616), .B(n2617), .Z(n2602) );
  NAND U2635 ( .A(\stack[0][0] ), .B(n2618), .Z(n2617) );
  XOR U2636 ( .A(n2619), .B(n2620), .Z(n2616) );
  XNOR U2637 ( .A(n2621), .B(n2622), .Z(n2620) );
  NAND U2638 ( .A(n2623), .B(n2624), .Z(n2498) );
  NANDN U2639 ( .A(n2599), .B(\stack[0][1] ), .Z(n2624) );
  ANDN U2640 ( .B(n2625), .A(n2561), .Z(n2623) );
  ANDN U2641 ( .B(x[1]), .A(n2503), .Z(n2561) );
  NANDN U2642 ( .A(n2563), .B(n2601), .Z(n2625) );
  AND U2643 ( .A(n2626), .B(n2627), .Z(n2563) );
  AND U2644 ( .A(n2628), .B(n2629), .Z(n2627) );
  NAND U2645 ( .A(n2630), .B(n2607), .Z(n2629) );
  XOR U2646 ( .A(n2631), .B(n2632), .Z(n2630) );
  AND U2647 ( .A(n2633), .B(n2634), .Z(n2628) );
  NAND U2648 ( .A(\stack[1][1] ), .B(n2635), .Z(n2634) );
  ANDN U2649 ( .B(\stack[0][1] ), .A(n2611), .Z(n2635) );
  NAND U2650 ( .A(n2636), .B(n2613), .Z(n2633) );
  NANDN U2651 ( .A(\stack[0][1] ), .B(n2637), .Z(n2636) );
  AND U2652 ( .A(n2638), .B(n2639), .Z(n2626) );
  NAND U2653 ( .A(\stack[0][1] ), .B(n2618), .Z(n2639) );
  XNOR U2654 ( .A(n2640), .B(n2641), .Z(n2638) );
  XNOR U2655 ( .A(n2642), .B(n2643), .Z(n2641) );
  NAND U2656 ( .A(n2644), .B(n2645), .Z(n2497) );
  NANDN U2657 ( .A(n2599), .B(\stack[0][2] ), .Z(n2645) );
  ANDN U2658 ( .B(n2646), .A(n2528), .Z(n2644) );
  ANDN U2659 ( .B(x[2]), .A(n2503), .Z(n2528) );
  NANDN U2660 ( .A(n2530), .B(n2601), .Z(n2646) );
  AND U2661 ( .A(n2647), .B(n2648), .Z(n2530) );
  AND U2662 ( .A(n2649), .B(n2650), .Z(n2648) );
  NAND U2663 ( .A(n2651), .B(n2607), .Z(n2650) );
  XNOR U2664 ( .A(n2652), .B(n2653), .Z(n2651) );
  XNOR U2665 ( .A(n2654), .B(n2655), .Z(n2653) );
  AND U2666 ( .A(n2656), .B(n2657), .Z(n2649) );
  NAND U2667 ( .A(\stack[1][2] ), .B(n2658), .Z(n2657) );
  ANDN U2668 ( .B(\stack[0][2] ), .A(n2611), .Z(n2658) );
  NAND U2669 ( .A(n2659), .B(n2613), .Z(n2656) );
  AND U2670 ( .A(n2661), .B(n2662), .Z(n2647) );
  NAND U2671 ( .A(\stack[0][2] ), .B(n2618), .Z(n2662) );
  XNOR U2672 ( .A(n2663), .B(n2664), .Z(n2661) );
  XNOR U2673 ( .A(n2665), .B(n2666), .Z(n2664) );
  NAND U2674 ( .A(n2667), .B(n2668), .Z(n2496) );
  NANDN U2675 ( .A(n2599), .B(\stack[0][3] ), .Z(n2668) );
  ANDN U2676 ( .B(n2669), .A(n2519), .Z(n2667) );
  ANDN U2677 ( .B(x[3]), .A(n2503), .Z(n2519) );
  NANDN U2678 ( .A(n2521), .B(n2601), .Z(n2669) );
  AND U2679 ( .A(n2670), .B(n2671), .Z(n2521) );
  AND U2680 ( .A(n2672), .B(n2673), .Z(n2671) );
  NAND U2681 ( .A(n2674), .B(n2607), .Z(n2673) );
  XNOR U2682 ( .A(n2675), .B(n2676), .Z(n2674) );
  XNOR U2683 ( .A(n2677), .B(n2678), .Z(n2676) );
  AND U2684 ( .A(n2679), .B(n2680), .Z(n2672) );
  NAND U2685 ( .A(\stack[1][3] ), .B(n2681), .Z(n2680) );
  ANDN U2686 ( .B(\stack[0][3] ), .A(n2611), .Z(n2681) );
  NAND U2687 ( .A(n2682), .B(n2613), .Z(n2679) );
  NAND U2688 ( .A(n2683), .B(n2684), .Z(n2682) );
  AND U2689 ( .A(n2685), .B(n2686), .Z(n2670) );
  NAND U2690 ( .A(\stack[0][3] ), .B(n2618), .Z(n2686) );
  XNOR U2691 ( .A(n2687), .B(n2688), .Z(n2685) );
  XNOR U2692 ( .A(n2689), .B(n2690), .Z(n2688) );
  NAND U2693 ( .A(n2691), .B(n2692), .Z(n2495) );
  NANDN U2694 ( .A(n2599), .B(\stack[0][4] ), .Z(n2692) );
  ANDN U2695 ( .B(n2693), .A(n2516), .Z(n2691) );
  ANDN U2696 ( .B(x[4]), .A(n2503), .Z(n2516) );
  NANDN U2697 ( .A(n2518), .B(n2601), .Z(n2693) );
  AND U2698 ( .A(n2694), .B(n2695), .Z(n2518) );
  AND U2699 ( .A(n2696), .B(n2697), .Z(n2695) );
  NAND U2700 ( .A(n2698), .B(n2607), .Z(n2697) );
  XOR U2701 ( .A(n2699), .B(n2700), .Z(n2698) );
  XNOR U2702 ( .A(n2701), .B(n2702), .Z(n2700) );
  AND U2703 ( .A(n2703), .B(n2704), .Z(n2696) );
  NAND U2704 ( .A(\stack[1][4] ), .B(n2705), .Z(n2704) );
  ANDN U2705 ( .B(\stack[0][4] ), .A(n2611), .Z(n2705) );
  NAND U2706 ( .A(n2706), .B(n2613), .Z(n2703) );
  NAND U2707 ( .A(n2707), .B(n2708), .Z(n2706) );
  AND U2708 ( .A(n2709), .B(n2710), .Z(n2694) );
  NAND U2709 ( .A(\stack[0][4] ), .B(n2618), .Z(n2710) );
  XNOR U2710 ( .A(n2711), .B(n2712), .Z(n2709) );
  XNOR U2711 ( .A(n2713), .B(n2714), .Z(n2712) );
  NAND U2712 ( .A(n2715), .B(n2716), .Z(n2494) );
  NANDN U2713 ( .A(n2599), .B(\stack[0][5] ), .Z(n2716) );
  ANDN U2714 ( .B(n2717), .A(n2513), .Z(n2715) );
  ANDN U2715 ( .B(x[5]), .A(n2503), .Z(n2513) );
  NANDN U2716 ( .A(n2515), .B(n2601), .Z(n2717) );
  AND U2717 ( .A(n2718), .B(n2719), .Z(n2515) );
  AND U2718 ( .A(n2720), .B(n2721), .Z(n2719) );
  NAND U2719 ( .A(n2722), .B(n2607), .Z(n2721) );
  XNOR U2720 ( .A(n2723), .B(n2724), .Z(n2722) );
  XOR U2721 ( .A(n2725), .B(n2726), .Z(n2724) );
  AND U2722 ( .A(n2727), .B(n2728), .Z(n2720) );
  NAND U2723 ( .A(\stack[0][5] ), .B(n2729), .Z(n2728) );
  ANDN U2724 ( .B(\stack[1][5] ), .A(n2611), .Z(n2729) );
  NAND U2725 ( .A(n2730), .B(n2613), .Z(n2727) );
  NAND U2726 ( .A(n2731), .B(n2732), .Z(n2730) );
  AND U2727 ( .A(n2733), .B(n2734), .Z(n2718) );
  NAND U2728 ( .A(\stack[0][5] ), .B(n2618), .Z(n2734) );
  XNOR U2729 ( .A(n2735), .B(n2736), .Z(n2733) );
  XNOR U2730 ( .A(n2737), .B(n2738), .Z(n2736) );
  NAND U2731 ( .A(n2739), .B(n2740), .Z(n2493) );
  NANDN U2732 ( .A(n2599), .B(\stack[0][6] ), .Z(n2740) );
  ANDN U2733 ( .B(n2741), .A(n2510), .Z(n2739) );
  ANDN U2734 ( .B(x[6]), .A(n2503), .Z(n2510) );
  NANDN U2735 ( .A(n2512), .B(n2601), .Z(n2741) );
  AND U2736 ( .A(n2742), .B(n2743), .Z(n2512) );
  AND U2737 ( .A(n2744), .B(n2745), .Z(n2743) );
  NAND U2738 ( .A(n2746), .B(n2607), .Z(n2745) );
  XOR U2739 ( .A(n2747), .B(n2748), .Z(n2746) );
  XNOR U2740 ( .A(n2749), .B(n2750), .Z(n2748) );
  AND U2741 ( .A(n2751), .B(n2752), .Z(n2744) );
  NAND U2742 ( .A(\stack[0][6] ), .B(n2753), .Z(n2752) );
  ANDN U2743 ( .B(\stack[1][6] ), .A(n2611), .Z(n2753) );
  NAND U2744 ( .A(n2754), .B(n2613), .Z(n2751) );
  NAND U2745 ( .A(n2755), .B(n2756), .Z(n2754) );
  AND U2746 ( .A(n2757), .B(n2758), .Z(n2742) );
  NAND U2747 ( .A(\stack[0][6] ), .B(n2618), .Z(n2758) );
  XNOR U2748 ( .A(n2759), .B(n2760), .Z(n2757) );
  XNOR U2749 ( .A(n2761), .B(n2762), .Z(n2760) );
  NAND U2750 ( .A(n2763), .B(n2764), .Z(n2492) );
  NANDN U2751 ( .A(n2599), .B(\stack[0][7] ), .Z(n2764) );
  ANDN U2752 ( .B(n2765), .A(n2507), .Z(n2763) );
  ANDN U2753 ( .B(x[7]), .A(n2503), .Z(n2507) );
  NANDN U2754 ( .A(n2509), .B(n2601), .Z(n2765) );
  AND U2755 ( .A(n2766), .B(n2767), .Z(n2509) );
  AND U2756 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2757 ( .A(n2770), .B(n2607), .Z(n2769) );
  XNOR U2758 ( .A(n2771), .B(n2772), .Z(n2770) );
  XOR U2759 ( .A(n2773), .B(n2774), .Z(n2772) );
  AND U2760 ( .A(n2775), .B(n2776), .Z(n2768) );
  NAND U2761 ( .A(\stack[0][7] ), .B(n2777), .Z(n2776) );
  ANDN U2762 ( .B(\stack[1][7] ), .A(n2611), .Z(n2777) );
  NAND U2763 ( .A(n2778), .B(n2613), .Z(n2775) );
  NAND U2764 ( .A(n2779), .B(n2780), .Z(n2778) );
  AND U2765 ( .A(n2781), .B(n2782), .Z(n2766) );
  NAND U2766 ( .A(\stack[0][7] ), .B(n2618), .Z(n2782) );
  XNOR U2767 ( .A(n2783), .B(n2784), .Z(n2781) );
  XNOR U2768 ( .A(n2785), .B(n2786), .Z(n2784) );
  NAND U2769 ( .A(n2787), .B(n2788), .Z(n2491) );
  NANDN U2770 ( .A(n2599), .B(\stack[0][8] ), .Z(n2788) );
  ANDN U2771 ( .B(n2789), .A(n2504), .Z(n2787) );
  ANDN U2772 ( .B(x[8]), .A(n2503), .Z(n2504) );
  NANDN U2773 ( .A(n2506), .B(n2601), .Z(n2789) );
  AND U2774 ( .A(n2790), .B(n2791), .Z(n2506) );
  AND U2775 ( .A(n2792), .B(n2793), .Z(n2791) );
  NAND U2776 ( .A(n2794), .B(n2607), .Z(n2793) );
  XOR U2777 ( .A(n2795), .B(n2796), .Z(n2794) );
  XNOR U2778 ( .A(n2797), .B(n2798), .Z(n2796) );
  AND U2779 ( .A(n2799), .B(n2800), .Z(n2792) );
  NAND U2780 ( .A(\stack[0][8] ), .B(n2801), .Z(n2800) );
  ANDN U2781 ( .B(\stack[1][8] ), .A(n2611), .Z(n2801) );
  NAND U2782 ( .A(n2802), .B(n2613), .Z(n2799) );
  NAND U2783 ( .A(n2803), .B(n2804), .Z(n2802) );
  AND U2784 ( .A(n2805), .B(n2806), .Z(n2790) );
  NAND U2785 ( .A(\stack[0][8] ), .B(n2618), .Z(n2806) );
  XNOR U2786 ( .A(n2807), .B(n2808), .Z(n2805) );
  XNOR U2787 ( .A(n2809), .B(n2810), .Z(n2808) );
  NAND U2788 ( .A(n2811), .B(n2812), .Z(n2490) );
  NANDN U2789 ( .A(n2599), .B(\stack[0][9] ), .Z(n2812) );
  ANDN U2790 ( .B(n2813), .A(n2500), .Z(n2811) );
  ANDN U2791 ( .B(x[9]), .A(n2503), .Z(n2500) );
  NANDN U2792 ( .A(n2502), .B(n2601), .Z(n2813) );
  AND U2793 ( .A(n2814), .B(n2815), .Z(n2502) );
  AND U2794 ( .A(n2816), .B(n2817), .Z(n2815) );
  NAND U2795 ( .A(n2818), .B(n2607), .Z(n2817) );
  XOR U2796 ( .A(n2819), .B(n2820), .Z(n2818) );
  XNOR U2797 ( .A(n2821), .B(n2822), .Z(n2820) );
  AND U2798 ( .A(n2823), .B(n2824), .Z(n2816) );
  NAND U2799 ( .A(\stack[1][9] ), .B(n2825), .Z(n2824) );
  ANDN U2800 ( .B(\stack[0][9] ), .A(n2611), .Z(n2825) );
  NAND U2801 ( .A(n2826), .B(n2613), .Z(n2823) );
  NAND U2802 ( .A(n2827), .B(n2828), .Z(n2826) );
  AND U2803 ( .A(n2829), .B(n2830), .Z(n2814) );
  NAND U2804 ( .A(\stack[0][9] ), .B(n2618), .Z(n2830) );
  XOR U2805 ( .A(n2831), .B(n2832), .Z(n2829) );
  XNOR U2806 ( .A(n2833), .B(n2834), .Z(n2832) );
  NAND U2807 ( .A(n2835), .B(n2836), .Z(n2489) );
  NANDN U2808 ( .A(n2599), .B(\stack[0][10] ), .Z(n2836) );
  ANDN U2809 ( .B(n2837), .A(n2591), .Z(n2835) );
  ANDN U2810 ( .B(x[10]), .A(n2503), .Z(n2591) );
  NANDN U2811 ( .A(n2593), .B(n2601), .Z(n2837) );
  AND U2812 ( .A(n2838), .B(n2839), .Z(n2593) );
  AND U2813 ( .A(n2840), .B(n2841), .Z(n2839) );
  NAND U2814 ( .A(n2842), .B(n2607), .Z(n2841) );
  XOR U2815 ( .A(n2843), .B(n2844), .Z(n2842) );
  XNOR U2816 ( .A(n2845), .B(n2846), .Z(n2844) );
  AND U2817 ( .A(n2847), .B(n2848), .Z(n2840) );
  NAND U2818 ( .A(\stack[1][10] ), .B(n2849), .Z(n2848) );
  ANDN U2819 ( .B(\stack[0][10] ), .A(n2611), .Z(n2849) );
  NAND U2820 ( .A(n2850), .B(n2613), .Z(n2847) );
  NAND U2821 ( .A(n2851), .B(n2852), .Z(n2850) );
  AND U2822 ( .A(n2853), .B(n2854), .Z(n2838) );
  NAND U2823 ( .A(\stack[0][10] ), .B(n2618), .Z(n2854) );
  XNOR U2824 ( .A(n2855), .B(n2856), .Z(n2853) );
  XNOR U2825 ( .A(n2857), .B(n2858), .Z(n2856) );
  NAND U2826 ( .A(n2859), .B(n2860), .Z(n2488) );
  NANDN U2827 ( .A(n2599), .B(\stack[0][11] ), .Z(n2860) );
  ANDN U2828 ( .B(n2861), .A(n2588), .Z(n2859) );
  ANDN U2829 ( .B(x[11]), .A(n2503), .Z(n2588) );
  NANDN U2830 ( .A(n2590), .B(n2601), .Z(n2861) );
  AND U2831 ( .A(n2862), .B(n2863), .Z(n2590) );
  AND U2832 ( .A(n2864), .B(n2865), .Z(n2863) );
  NAND U2833 ( .A(n2866), .B(n2607), .Z(n2865) );
  XNOR U2834 ( .A(n2867), .B(n2868), .Z(n2866) );
  XOR U2835 ( .A(n2869), .B(n2870), .Z(n2868) );
  AND U2836 ( .A(n2871), .B(n2872), .Z(n2864) );
  NAND U2837 ( .A(\stack[1][11] ), .B(n2873), .Z(n2872) );
  ANDN U2838 ( .B(\stack[0][11] ), .A(n2611), .Z(n2873) );
  NAND U2839 ( .A(n2874), .B(n2613), .Z(n2871) );
  NAND U2840 ( .A(n2875), .B(n2876), .Z(n2874) );
  AND U2841 ( .A(n2877), .B(n2878), .Z(n2862) );
  NAND U2842 ( .A(\stack[0][11] ), .B(n2618), .Z(n2878) );
  XNOR U2843 ( .A(n2879), .B(n2880), .Z(n2877) );
  XNOR U2844 ( .A(n2881), .B(n2882), .Z(n2880) );
  NAND U2845 ( .A(n2883), .B(n2884), .Z(n2487) );
  NANDN U2846 ( .A(n2599), .B(\stack[0][12] ), .Z(n2884) );
  ANDN U2847 ( .B(n2885), .A(n2585), .Z(n2883) );
  ANDN U2848 ( .B(x[12]), .A(n2503), .Z(n2585) );
  NANDN U2849 ( .A(n2587), .B(n2601), .Z(n2885) );
  AND U2850 ( .A(n2886), .B(n2887), .Z(n2587) );
  AND U2851 ( .A(n2888), .B(n2889), .Z(n2887) );
  NAND U2852 ( .A(n2890), .B(n2607), .Z(n2889) );
  XOR U2853 ( .A(n2891), .B(n2892), .Z(n2890) );
  XNOR U2854 ( .A(n2893), .B(n2894), .Z(n2892) );
  AND U2855 ( .A(n2895), .B(n2896), .Z(n2888) );
  NAND U2856 ( .A(\stack[1][12] ), .B(n2897), .Z(n2896) );
  ANDN U2857 ( .B(\stack[0][12] ), .A(n2611), .Z(n2897) );
  NAND U2858 ( .A(n2898), .B(n2613), .Z(n2895) );
  NAND U2859 ( .A(n2899), .B(n2900), .Z(n2898) );
  AND U2860 ( .A(n2901), .B(n2902), .Z(n2886) );
  NAND U2861 ( .A(\stack[0][12] ), .B(n2618), .Z(n2902) );
  XNOR U2862 ( .A(n2903), .B(n2904), .Z(n2901) );
  XNOR U2863 ( .A(n2905), .B(n2906), .Z(n2904) );
  NAND U2864 ( .A(n2907), .B(n2908), .Z(n2486) );
  NANDN U2865 ( .A(n2599), .B(\stack[0][13] ), .Z(n2908) );
  ANDN U2866 ( .B(n2909), .A(n2582), .Z(n2907) );
  ANDN U2867 ( .B(x[13]), .A(n2503), .Z(n2582) );
  NANDN U2868 ( .A(n2584), .B(n2601), .Z(n2909) );
  AND U2869 ( .A(n2910), .B(n2911), .Z(n2584) );
  AND U2870 ( .A(n2912), .B(n2913), .Z(n2911) );
  NAND U2871 ( .A(n2914), .B(n2607), .Z(n2913) );
  XOR U2872 ( .A(n2915), .B(n2916), .Z(n2914) );
  XNOR U2873 ( .A(n2917), .B(n2918), .Z(n2916) );
  AND U2874 ( .A(n2919), .B(n2920), .Z(n2912) );
  NAND U2875 ( .A(\stack[1][13] ), .B(n2921), .Z(n2920) );
  ANDN U2876 ( .B(\stack[0][13] ), .A(n2611), .Z(n2921) );
  NAND U2877 ( .A(n2922), .B(n2613), .Z(n2919) );
  NAND U2878 ( .A(n2923), .B(n2924), .Z(n2922) );
  AND U2879 ( .A(n2925), .B(n2926), .Z(n2910) );
  NAND U2880 ( .A(\stack[0][13] ), .B(n2618), .Z(n2926) );
  XNOR U2881 ( .A(n2927), .B(n2928), .Z(n2925) );
  XNOR U2882 ( .A(n2929), .B(n2930), .Z(n2928) );
  NAND U2883 ( .A(n2931), .B(n2932), .Z(n2485) );
  NANDN U2884 ( .A(n2599), .B(\stack[0][14] ), .Z(n2932) );
  ANDN U2885 ( .B(n2933), .A(n2579), .Z(n2931) );
  ANDN U2886 ( .B(x[14]), .A(n2503), .Z(n2579) );
  NANDN U2887 ( .A(n2581), .B(n2601), .Z(n2933) );
  AND U2888 ( .A(n2934), .B(n2935), .Z(n2581) );
  AND U2889 ( .A(n2936), .B(n2937), .Z(n2935) );
  NAND U2890 ( .A(n2938), .B(n2607), .Z(n2937) );
  XOR U2891 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR U2892 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2893 ( .A(n2943), .B(n2944), .Z(n2936) );
  NAND U2894 ( .A(\stack[1][14] ), .B(n2945), .Z(n2944) );
  ANDN U2895 ( .B(\stack[0][14] ), .A(n2611), .Z(n2945) );
  NAND U2896 ( .A(n2946), .B(n2613), .Z(n2943) );
  NAND U2897 ( .A(n2947), .B(n2948), .Z(n2946) );
  AND U2898 ( .A(n2949), .B(n2950), .Z(n2934) );
  NAND U2899 ( .A(\stack[0][14] ), .B(n2618), .Z(n2950) );
  XNOR U2900 ( .A(n2951), .B(n2952), .Z(n2949) );
  XNOR U2901 ( .A(n2953), .B(n2954), .Z(n2952) );
  NAND U2902 ( .A(n2955), .B(n2956), .Z(n2484) );
  NANDN U2903 ( .A(n2599), .B(\stack[0][15] ), .Z(n2956) );
  ANDN U2904 ( .B(n2957), .A(n2576), .Z(n2955) );
  ANDN U2905 ( .B(x[15]), .A(n2503), .Z(n2576) );
  NANDN U2906 ( .A(n2578), .B(n2601), .Z(n2957) );
  AND U2907 ( .A(n2958), .B(n2959), .Z(n2578) );
  AND U2908 ( .A(n2960), .B(n2961), .Z(n2959) );
  NAND U2909 ( .A(n2962), .B(n2607), .Z(n2961) );
  XOR U2910 ( .A(n2963), .B(n2964), .Z(n2962) );
  XNOR U2911 ( .A(n2965), .B(n2966), .Z(n2964) );
  AND U2912 ( .A(n2967), .B(n2968), .Z(n2960) );
  NAND U2913 ( .A(\stack[1][15] ), .B(n2969), .Z(n2968) );
  ANDN U2914 ( .B(\stack[0][15] ), .A(n2611), .Z(n2969) );
  NAND U2915 ( .A(n2970), .B(n2613), .Z(n2967) );
  NAND U2916 ( .A(n2971), .B(n2972), .Z(n2970) );
  AND U2917 ( .A(n2973), .B(n2974), .Z(n2958) );
  NAND U2918 ( .A(\stack[0][15] ), .B(n2618), .Z(n2974) );
  XNOR U2919 ( .A(n2975), .B(n2976), .Z(n2973) );
  XNOR U2920 ( .A(n2977), .B(n2978), .Z(n2976) );
  NAND U2921 ( .A(n2979), .B(n2980), .Z(n2483) );
  NANDN U2922 ( .A(n2599), .B(\stack[0][16] ), .Z(n2980) );
  ANDN U2923 ( .B(n2981), .A(n2573), .Z(n2979) );
  ANDN U2924 ( .B(x[16]), .A(n2503), .Z(n2573) );
  NANDN U2925 ( .A(n2575), .B(n2601), .Z(n2981) );
  AND U2926 ( .A(n2982), .B(n2983), .Z(n2575) );
  AND U2927 ( .A(n2984), .B(n2985), .Z(n2983) );
  NAND U2928 ( .A(n2986), .B(n2607), .Z(n2985) );
  XOR U2929 ( .A(n2987), .B(n2988), .Z(n2986) );
  XOR U2930 ( .A(n2989), .B(n2990), .Z(n2988) );
  AND U2931 ( .A(n2991), .B(n2992), .Z(n2984) );
  NAND U2932 ( .A(\stack[0][16] ), .B(n2993), .Z(n2992) );
  ANDN U2933 ( .B(\stack[1][16] ), .A(n2611), .Z(n2993) );
  NAND U2934 ( .A(n2994), .B(n2613), .Z(n2991) );
  NAND U2935 ( .A(n2995), .B(n2996), .Z(n2994) );
  AND U2936 ( .A(n2997), .B(n2998), .Z(n2982) );
  NAND U2937 ( .A(\stack[0][16] ), .B(n2618), .Z(n2998) );
  XNOR U2938 ( .A(n2999), .B(n3000), .Z(n2997) );
  XNOR U2939 ( .A(n3001), .B(n3002), .Z(n3000) );
  NAND U2940 ( .A(n3003), .B(n3004), .Z(n2482) );
  NANDN U2941 ( .A(n2599), .B(\stack[0][17] ), .Z(n3004) );
  ANDN U2942 ( .B(n3005), .A(n2570), .Z(n3003) );
  ANDN U2943 ( .B(x[17]), .A(n2503), .Z(n2570) );
  NANDN U2944 ( .A(n2572), .B(n2601), .Z(n3005) );
  AND U2945 ( .A(n3006), .B(n3007), .Z(n2572) );
  AND U2946 ( .A(n3008), .B(n3009), .Z(n3007) );
  NAND U2947 ( .A(n3010), .B(n2607), .Z(n3009) );
  XOR U2948 ( .A(n3011), .B(n3012), .Z(n3010) );
  XNOR U2949 ( .A(n3013), .B(n3014), .Z(n3012) );
  AND U2950 ( .A(n3015), .B(n3016), .Z(n3008) );
  NAND U2951 ( .A(\stack[0][17] ), .B(n3017), .Z(n3016) );
  ANDN U2952 ( .B(\stack[1][17] ), .A(n2611), .Z(n3017) );
  NAND U2953 ( .A(n3018), .B(n2613), .Z(n3015) );
  NAND U2954 ( .A(n3019), .B(n3020), .Z(n3018) );
  AND U2955 ( .A(n3021), .B(n3022), .Z(n3006) );
  NAND U2956 ( .A(\stack[0][17] ), .B(n2618), .Z(n3022) );
  XNOR U2957 ( .A(n3023), .B(n3024), .Z(n3021) );
  XNOR U2958 ( .A(n3025), .B(n3026), .Z(n3024) );
  NAND U2959 ( .A(n3027), .B(n3028), .Z(n2481) );
  NANDN U2960 ( .A(n2599), .B(\stack[0][18] ), .Z(n3028) );
  ANDN U2961 ( .B(n3029), .A(n2567), .Z(n3027) );
  ANDN U2962 ( .B(x[18]), .A(n2503), .Z(n2567) );
  NANDN U2963 ( .A(n2569), .B(n2601), .Z(n3029) );
  AND U2964 ( .A(n3030), .B(n3031), .Z(n2569) );
  AND U2965 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U2966 ( .A(n3034), .B(n2607), .Z(n3033) );
  XOR U2967 ( .A(n3035), .B(n3036), .Z(n3034) );
  XOR U2968 ( .A(n3037), .B(n3038), .Z(n3036) );
  AND U2969 ( .A(n3039), .B(n3040), .Z(n3032) );
  NAND U2970 ( .A(\stack[0][18] ), .B(n3041), .Z(n3040) );
  ANDN U2971 ( .B(\stack[1][18] ), .A(n2611), .Z(n3041) );
  NAND U2972 ( .A(n3042), .B(n2613), .Z(n3039) );
  NAND U2973 ( .A(n3043), .B(n3044), .Z(n3042) );
  AND U2974 ( .A(n3045), .B(n3046), .Z(n3030) );
  NAND U2975 ( .A(\stack[0][18] ), .B(n2618), .Z(n3046) );
  XNOR U2976 ( .A(n3047), .B(n3048), .Z(n3045) );
  XNOR U2977 ( .A(n3049), .B(n3050), .Z(n3048) );
  NAND U2978 ( .A(n3051), .B(n3052), .Z(n2480) );
  NANDN U2979 ( .A(n2599), .B(\stack[0][19] ), .Z(n3052) );
  ANDN U2980 ( .B(n3053), .A(n2564), .Z(n3051) );
  ANDN U2981 ( .B(x[19]), .A(n2503), .Z(n2564) );
  NANDN U2982 ( .A(n2566), .B(n2601), .Z(n3053) );
  AND U2983 ( .A(n3054), .B(n3055), .Z(n2566) );
  AND U2984 ( .A(n3056), .B(n3057), .Z(n3055) );
  NAND U2985 ( .A(n3058), .B(n2607), .Z(n3057) );
  XOR U2986 ( .A(n3059), .B(n3060), .Z(n3058) );
  XNOR U2987 ( .A(n3061), .B(n3062), .Z(n3060) );
  AND U2988 ( .A(n3063), .B(n3064), .Z(n3056) );
  NAND U2989 ( .A(\stack[0][19] ), .B(n3065), .Z(n3064) );
  ANDN U2990 ( .B(\stack[1][19] ), .A(n2611), .Z(n3065) );
  NAND U2991 ( .A(n3066), .B(n2613), .Z(n3063) );
  NAND U2992 ( .A(n3067), .B(n3068), .Z(n3066) );
  AND U2993 ( .A(n3069), .B(n3070), .Z(n3054) );
  NAND U2994 ( .A(\stack[0][19] ), .B(n2618), .Z(n3070) );
  XNOR U2995 ( .A(n3071), .B(n3072), .Z(n3069) );
  XNOR U2996 ( .A(n3073), .B(n3074), .Z(n3072) );
  NAND U2997 ( .A(n3075), .B(n3076), .Z(n2479) );
  NANDN U2998 ( .A(n2599), .B(\stack[0][20] ), .Z(n3076) );
  ANDN U2999 ( .B(n3077), .A(n2558), .Z(n3075) );
  ANDN U3000 ( .B(x[20]), .A(n2503), .Z(n2558) );
  NANDN U3001 ( .A(n2560), .B(n2601), .Z(n3077) );
  AND U3002 ( .A(n3078), .B(n3079), .Z(n2560) );
  AND U3003 ( .A(n3080), .B(n3081), .Z(n3079) );
  NAND U3004 ( .A(n3082), .B(n2607), .Z(n3081) );
  XOR U3005 ( .A(n3083), .B(n3084), .Z(n3082) );
  XOR U3006 ( .A(n3085), .B(n3086), .Z(n3084) );
  AND U3007 ( .A(n3087), .B(n3088), .Z(n3080) );
  NAND U3008 ( .A(\stack[0][20] ), .B(n3089), .Z(n3088) );
  ANDN U3009 ( .B(\stack[1][20] ), .A(n2611), .Z(n3089) );
  NAND U3010 ( .A(n3090), .B(n2613), .Z(n3087) );
  NAND U3011 ( .A(n3091), .B(n3092), .Z(n3090) );
  AND U3012 ( .A(n3093), .B(n3094), .Z(n3078) );
  NAND U3013 ( .A(\stack[0][20] ), .B(n2618), .Z(n3094) );
  XNOR U3014 ( .A(n3095), .B(n3096), .Z(n3093) );
  XNOR U3015 ( .A(n3097), .B(n3098), .Z(n3096) );
  NAND U3016 ( .A(n3099), .B(n3100), .Z(n2478) );
  NANDN U3017 ( .A(n2599), .B(\stack[0][21] ), .Z(n3100) );
  ANDN U3018 ( .B(n3101), .A(n2555), .Z(n3099) );
  ANDN U3019 ( .B(x[21]), .A(n2503), .Z(n2555) );
  NANDN U3020 ( .A(n2557), .B(n2601), .Z(n3101) );
  AND U3021 ( .A(n3102), .B(n3103), .Z(n2557) );
  AND U3022 ( .A(n3104), .B(n3105), .Z(n3103) );
  NAND U3023 ( .A(n3106), .B(n2607), .Z(n3105) );
  XOR U3024 ( .A(n3107), .B(n3108), .Z(n3106) );
  XNOR U3025 ( .A(n3109), .B(n3110), .Z(n3108) );
  AND U3026 ( .A(n3111), .B(n3112), .Z(n3104) );
  NAND U3027 ( .A(\stack[0][21] ), .B(n3113), .Z(n3112) );
  ANDN U3028 ( .B(\stack[1][21] ), .A(n2611), .Z(n3113) );
  NAND U3029 ( .A(n3114), .B(n2613), .Z(n3111) );
  NAND U3030 ( .A(n3115), .B(n3116), .Z(n3114) );
  AND U3031 ( .A(n3117), .B(n3118), .Z(n3102) );
  NAND U3032 ( .A(\stack[0][21] ), .B(n2618), .Z(n3118) );
  XNOR U3033 ( .A(n3119), .B(n3120), .Z(n3117) );
  XNOR U3034 ( .A(n3121), .B(n3122), .Z(n3120) );
  NAND U3035 ( .A(n3123), .B(n3124), .Z(n2477) );
  NANDN U3036 ( .A(n2599), .B(\stack[0][22] ), .Z(n3124) );
  ANDN U3037 ( .B(n3125), .A(n2552), .Z(n3123) );
  ANDN U3038 ( .B(x[22]), .A(n2503), .Z(n2552) );
  NANDN U3039 ( .A(n2554), .B(n2601), .Z(n3125) );
  AND U3040 ( .A(n3126), .B(n3127), .Z(n2554) );
  AND U3041 ( .A(n3128), .B(n3129), .Z(n3127) );
  NAND U3042 ( .A(n3130), .B(n2607), .Z(n3129) );
  XOR U3043 ( .A(n3131), .B(n3132), .Z(n3130) );
  XOR U3044 ( .A(n3133), .B(n3134), .Z(n3132) );
  AND U3045 ( .A(n3135), .B(n3136), .Z(n3128) );
  NAND U3046 ( .A(\stack[0][22] ), .B(n3137), .Z(n3136) );
  ANDN U3047 ( .B(\stack[1][22] ), .A(n2611), .Z(n3137) );
  NAND U3048 ( .A(n3138), .B(n2613), .Z(n3135) );
  NAND U3049 ( .A(n3139), .B(n3140), .Z(n3138) );
  AND U3050 ( .A(n3141), .B(n3142), .Z(n3126) );
  NAND U3051 ( .A(\stack[0][22] ), .B(n2618), .Z(n3142) );
  XNOR U3052 ( .A(n3143), .B(n3144), .Z(n3141) );
  XNOR U3053 ( .A(n3145), .B(n3146), .Z(n3144) );
  NAND U3054 ( .A(n3147), .B(n3148), .Z(n2476) );
  NANDN U3055 ( .A(n2599), .B(\stack[0][23] ), .Z(n3148) );
  ANDN U3056 ( .B(n3149), .A(n2549), .Z(n3147) );
  ANDN U3057 ( .B(x[23]), .A(n2503), .Z(n2549) );
  NANDN U3058 ( .A(n2551), .B(n2601), .Z(n3149) );
  AND U3059 ( .A(n3150), .B(n3151), .Z(n2551) );
  AND U3060 ( .A(n3152), .B(n3153), .Z(n3151) );
  NAND U3061 ( .A(n3154), .B(n2607), .Z(n3153) );
  XOR U3062 ( .A(n3155), .B(n3156), .Z(n3154) );
  XNOR U3063 ( .A(n3157), .B(n3158), .Z(n3156) );
  AND U3064 ( .A(n3159), .B(n3160), .Z(n3152) );
  NAND U3065 ( .A(\stack[0][23] ), .B(n3161), .Z(n3160) );
  ANDN U3066 ( .B(\stack[1][23] ), .A(n2611), .Z(n3161) );
  NAND U3067 ( .A(n3162), .B(n2613), .Z(n3159) );
  NAND U3068 ( .A(n3163), .B(n3164), .Z(n3162) );
  AND U3069 ( .A(n3165), .B(n3166), .Z(n3150) );
  NAND U3070 ( .A(\stack[0][23] ), .B(n2618), .Z(n3166) );
  XNOR U3071 ( .A(n3167), .B(n3168), .Z(n3165) );
  XNOR U3072 ( .A(n3169), .B(n3170), .Z(n3168) );
  NAND U3073 ( .A(n3171), .B(n3172), .Z(n2475) );
  NANDN U3074 ( .A(n2599), .B(\stack[0][24] ), .Z(n3172) );
  ANDN U3075 ( .B(n3173), .A(n2546), .Z(n3171) );
  ANDN U3076 ( .B(x[24]), .A(n2503), .Z(n2546) );
  NANDN U3077 ( .A(n2548), .B(n2601), .Z(n3173) );
  AND U3078 ( .A(n3174), .B(n3175), .Z(n2548) );
  AND U3079 ( .A(n3176), .B(n3177), .Z(n3175) );
  NAND U3080 ( .A(n3178), .B(n2607), .Z(n3177) );
  XOR U3081 ( .A(n3179), .B(n3180), .Z(n3178) );
  XOR U3082 ( .A(n3181), .B(n3182), .Z(n3180) );
  AND U3083 ( .A(n3183), .B(n3184), .Z(n3176) );
  NAND U3084 ( .A(\stack[0][24] ), .B(n3185), .Z(n3184) );
  ANDN U3085 ( .B(\stack[1][24] ), .A(n2611), .Z(n3185) );
  NAND U3086 ( .A(n3186), .B(n2613), .Z(n3183) );
  NAND U3087 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3088 ( .A(n3189), .B(n3190), .Z(n3174) );
  NAND U3089 ( .A(\stack[0][24] ), .B(n2618), .Z(n3190) );
  XNOR U3090 ( .A(n3191), .B(n3192), .Z(n3189) );
  XNOR U3091 ( .A(n3193), .B(n3194), .Z(n3192) );
  NAND U3092 ( .A(n3195), .B(n3196), .Z(n2474) );
  NANDN U3093 ( .A(n2599), .B(\stack[0][25] ), .Z(n3196) );
  ANDN U3094 ( .B(n3197), .A(n2543), .Z(n3195) );
  ANDN U3095 ( .B(x[25]), .A(n2503), .Z(n2543) );
  NANDN U3096 ( .A(n2545), .B(n2601), .Z(n3197) );
  AND U3097 ( .A(n3198), .B(n3199), .Z(n2545) );
  AND U3098 ( .A(n3200), .B(n3201), .Z(n3199) );
  NAND U3099 ( .A(n3202), .B(n2607), .Z(n3201) );
  XOR U3100 ( .A(n3203), .B(n3204), .Z(n3202) );
  XNOR U3101 ( .A(n3205), .B(n3206), .Z(n3204) );
  AND U3102 ( .A(n3207), .B(n3208), .Z(n3200) );
  NAND U3103 ( .A(\stack[0][25] ), .B(n3209), .Z(n3208) );
  ANDN U3104 ( .B(\stack[1][25] ), .A(n2611), .Z(n3209) );
  NAND U3105 ( .A(n3210), .B(n2613), .Z(n3207) );
  NAND U3106 ( .A(n3211), .B(n3212), .Z(n3210) );
  AND U3107 ( .A(n3213), .B(n3214), .Z(n3198) );
  NAND U3108 ( .A(\stack[0][25] ), .B(n2618), .Z(n3214) );
  XNOR U3109 ( .A(n3215), .B(n3216), .Z(n3213) );
  XNOR U3110 ( .A(n3217), .B(n3218), .Z(n3216) );
  NAND U3111 ( .A(n3219), .B(n3220), .Z(n2473) );
  NANDN U3112 ( .A(n2599), .B(\stack[0][26] ), .Z(n3220) );
  ANDN U3113 ( .B(n3221), .A(n2540), .Z(n3219) );
  ANDN U3114 ( .B(x[26]), .A(n2503), .Z(n2540) );
  NANDN U3115 ( .A(n2542), .B(n2601), .Z(n3221) );
  AND U3116 ( .A(n3222), .B(n3223), .Z(n2542) );
  AND U3117 ( .A(n3224), .B(n3225), .Z(n3223) );
  NAND U3118 ( .A(n3226), .B(n2607), .Z(n3225) );
  XOR U3119 ( .A(n3227), .B(n3228), .Z(n3226) );
  XOR U3120 ( .A(n3229), .B(n3230), .Z(n3228) );
  AND U3121 ( .A(n3231), .B(n3232), .Z(n3224) );
  NAND U3122 ( .A(\stack[0][26] ), .B(n3233), .Z(n3232) );
  ANDN U3123 ( .B(\stack[1][26] ), .A(n2611), .Z(n3233) );
  NAND U3124 ( .A(n3234), .B(n2613), .Z(n3231) );
  NAND U3125 ( .A(n3235), .B(n3236), .Z(n3234) );
  AND U3126 ( .A(n3237), .B(n3238), .Z(n3222) );
  NAND U3127 ( .A(\stack[0][26] ), .B(n2618), .Z(n3238) );
  XNOR U3128 ( .A(n3239), .B(n3240), .Z(n3237) );
  XNOR U3129 ( .A(n3241), .B(n3242), .Z(n3240) );
  NAND U3130 ( .A(n3243), .B(n3244), .Z(n2472) );
  NANDN U3131 ( .A(n2599), .B(\stack[0][27] ), .Z(n3244) );
  ANDN U3132 ( .B(n3245), .A(n2537), .Z(n3243) );
  ANDN U3133 ( .B(x[27]), .A(n2503), .Z(n2537) );
  NANDN U3134 ( .A(n2539), .B(n2601), .Z(n3245) );
  AND U3135 ( .A(n3246), .B(n3247), .Z(n2539) );
  AND U3136 ( .A(n3248), .B(n3249), .Z(n3247) );
  NAND U3137 ( .A(n3250), .B(n2607), .Z(n3249) );
  XOR U3138 ( .A(n3251), .B(n3252), .Z(n3250) );
  XNOR U3139 ( .A(n3253), .B(n3254), .Z(n3252) );
  AND U3140 ( .A(n3255), .B(n3256), .Z(n3248) );
  NAND U3141 ( .A(\stack[0][27] ), .B(n3257), .Z(n3256) );
  ANDN U3142 ( .B(\stack[1][27] ), .A(n2611), .Z(n3257) );
  NAND U3143 ( .A(n3258), .B(n2613), .Z(n3255) );
  NAND U3144 ( .A(n3259), .B(n3260), .Z(n3258) );
  AND U3145 ( .A(n3261), .B(n3262), .Z(n3246) );
  NAND U3146 ( .A(\stack[0][27] ), .B(n2618), .Z(n3262) );
  XNOR U3147 ( .A(n3263), .B(n3264), .Z(n3261) );
  XNOR U3148 ( .A(n3265), .B(n3266), .Z(n3264) );
  NAND U3149 ( .A(n3267), .B(n3268), .Z(n2471) );
  NANDN U3150 ( .A(n2599), .B(\stack[0][28] ), .Z(n3268) );
  ANDN U3151 ( .B(n3269), .A(n2534), .Z(n3267) );
  ANDN U3152 ( .B(x[28]), .A(n2503), .Z(n2534) );
  NANDN U3153 ( .A(n2536), .B(n2601), .Z(n3269) );
  AND U3154 ( .A(n3270), .B(n3271), .Z(n2536) );
  AND U3155 ( .A(n3272), .B(n3273), .Z(n3271) );
  NAND U3156 ( .A(n3274), .B(n2607), .Z(n3273) );
  XOR U3157 ( .A(n3275), .B(n3276), .Z(n3274) );
  XOR U3158 ( .A(n3277), .B(n3278), .Z(n3276) );
  AND U3159 ( .A(n3279), .B(n3280), .Z(n3272) );
  NAND U3160 ( .A(\stack[1][28] ), .B(n3281), .Z(n3280) );
  ANDN U3161 ( .B(\stack[0][28] ), .A(n2611), .Z(n3281) );
  NAND U3162 ( .A(n3282), .B(n2613), .Z(n3279) );
  AND U3163 ( .A(n3284), .B(n3285), .Z(n3270) );
  NAND U3164 ( .A(\stack[0][28] ), .B(n2618), .Z(n3285) );
  XNOR U3165 ( .A(n3286), .B(n3287), .Z(n3284) );
  XNOR U3166 ( .A(n3288), .B(n3289), .Z(n3287) );
  NAND U3167 ( .A(n3290), .B(n3291), .Z(n2470) );
  NANDN U3168 ( .A(n2599), .B(\stack[0][29] ), .Z(n3291) );
  ANDN U3169 ( .B(n3292), .A(n2531), .Z(n3290) );
  ANDN U3170 ( .B(x[29]), .A(n2503), .Z(n2531) );
  NANDN U3171 ( .A(n2533), .B(n2601), .Z(n3292) );
  AND U3172 ( .A(n3293), .B(n3294), .Z(n2533) );
  AND U3173 ( .A(n3295), .B(n3296), .Z(n3294) );
  NAND U3174 ( .A(n3297), .B(n2607), .Z(n3296) );
  XOR U3175 ( .A(n3298), .B(n3299), .Z(n3297) );
  XNOR U3176 ( .A(n3300), .B(n3301), .Z(n3299) );
  AND U3177 ( .A(n3302), .B(n3303), .Z(n3295) );
  NAND U3178 ( .A(\stack[0][29] ), .B(n3304), .Z(n3303) );
  ANDN U3179 ( .B(\stack[1][29] ), .A(n2611), .Z(n3304) );
  NAND U3180 ( .A(n3305), .B(n2613), .Z(n3302) );
  AND U3181 ( .A(n3307), .B(n3308), .Z(n3293) );
  NAND U3182 ( .A(\stack[0][29] ), .B(n2618), .Z(n3308) );
  XNOR U3183 ( .A(n3309), .B(n3310), .Z(n3307) );
  XNOR U3184 ( .A(n3311), .B(n3312), .Z(n3310) );
  NAND U3185 ( .A(n3313), .B(n3314), .Z(n2469) );
  NANDN U3186 ( .A(n2599), .B(\stack[0][30] ), .Z(n3314) );
  ANDN U3187 ( .B(n3315), .A(n2525), .Z(n3313) );
  ANDN U3188 ( .B(x[30]), .A(n2503), .Z(n2525) );
  NANDN U3189 ( .A(n2527), .B(n2601), .Z(n3315) );
  AND U3190 ( .A(n3316), .B(n3317), .Z(n2527) );
  AND U3191 ( .A(n3318), .B(n3319), .Z(n3317) );
  NAND U3192 ( .A(n3320), .B(n2607), .Z(n3319) );
  XOR U3193 ( .A(n3321), .B(n3322), .Z(n3320) );
  XNOR U3194 ( .A(n3323), .B(n3324), .Z(n3322) );
  AND U3195 ( .A(n3325), .B(n3326), .Z(n3318) );
  NAND U3196 ( .A(\stack[0][30] ), .B(n3327), .Z(n3326) );
  ANDN U3197 ( .B(\stack[1][30] ), .A(n2611), .Z(n3327) );
  NAND U3198 ( .A(n3328), .B(n2613), .Z(n3325) );
  AND U3199 ( .A(n3329), .B(n3330), .Z(n3316) );
  NAND U3200 ( .A(\stack[0][30] ), .B(n2618), .Z(n3330) );
  XOR U3201 ( .A(n3331), .B(n3332), .Z(n3329) );
  XOR U3202 ( .A(n3333), .B(n3334), .Z(n3332) );
  NAND U3203 ( .A(n3335), .B(n3336), .Z(n2468) );
  NANDN U3204 ( .A(n2599), .B(\stack[0][31] ), .Z(n3336) );
  NANDN U3205 ( .A(n3337), .B(n3338), .Z(n2599) );
  ANDN U3206 ( .B(n2503), .A(n3339), .Z(n3338) );
  ANDN U3207 ( .B(n3340), .A(n2522), .Z(n3335) );
  ANDN U3208 ( .B(x[31]), .A(n2503), .Z(n2522) );
  NANDN U3209 ( .A(n2524), .B(n2601), .Z(n3340) );
  OR U3210 ( .A(n3339), .B(n3337), .Z(n2601) );
  AND U3211 ( .A(n3341), .B(n3342), .Z(n2524) );
  AND U3212 ( .A(n3343), .B(n3344), .Z(n3342) );
  NAND U3213 ( .A(n3345), .B(n2607), .Z(n3344) );
  AND U3214 ( .A(n3346), .B(n3347), .Z(n3345) );
  NANDN U3215 ( .A(n3348), .B(n3349), .Z(n3347) );
  NAND U3216 ( .A(n3350), .B(n3348), .Z(n3346) );
  XOR U3217 ( .A(n3351), .B(n3352), .Z(n3348) );
  XOR U3218 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U3219 ( .A(n3355), .B(n3356), .Z(n3354) );
  XOR U3220 ( .A(n3357), .B(n3358), .Z(n3356) );
  XOR U3221 ( .A(n3359), .B(n3360), .Z(n3358) );
  XOR U3222 ( .A(n3361), .B(n3362), .Z(n3360) );
  NAND U3223 ( .A(n3363), .B(n3364), .Z(n3362) );
  NAND U3224 ( .A(n3365), .B(n3366), .Z(n3364) );
  NANDN U3225 ( .A(n3367), .B(n3368), .Z(n3363) );
  AND U3226 ( .A(\stack[1][1] ), .B(\stack[0][30] ), .Z(n3361) );
  XOR U3227 ( .A(n3369), .B(n3370), .Z(n3359) );
  XOR U3228 ( .A(n3371), .B(n3372), .Z(n3370) );
  XOR U3229 ( .A(n3373), .B(n3374), .Z(n3372) );
  XOR U3230 ( .A(n3375), .B(n3376), .Z(n3374) );
  AND U3231 ( .A(n3377), .B(n3378), .Z(n3376) );
  NAND U3232 ( .A(n3379), .B(n3380), .Z(n3378) );
  NANDN U3233 ( .A(n3381), .B(n3382), .Z(n3377) );
  AND U3234 ( .A(\stack[1][3] ), .B(\stack[0][28] ), .Z(n3375) );
  XOR U3235 ( .A(n3383), .B(n3384), .Z(n3373) );
  XOR U3236 ( .A(n3385), .B(n3386), .Z(n3384) );
  XOR U3237 ( .A(n3387), .B(n3388), .Z(n3386) );
  XOR U3238 ( .A(n3389), .B(n3390), .Z(n3388) );
  AND U3239 ( .A(n3391), .B(n3392), .Z(n3390) );
  NAND U3240 ( .A(n3393), .B(n3394), .Z(n3392) );
  NANDN U3241 ( .A(n3395), .B(n3396), .Z(n3391) );
  AND U3242 ( .A(\stack[1][7] ), .B(\stack[0][24] ), .Z(n3389) );
  XOR U3243 ( .A(n3397), .B(n3398), .Z(n3387) );
  XOR U3244 ( .A(n3399), .B(n3400), .Z(n3398) );
  XOR U3245 ( .A(n3401), .B(n3402), .Z(n3400) );
  XOR U3246 ( .A(n3403), .B(n3404), .Z(n3402) );
  AND U3247 ( .A(n3405), .B(n3406), .Z(n3404) );
  NAND U3248 ( .A(n3407), .B(n3408), .Z(n3406) );
  NANDN U3249 ( .A(n3409), .B(n3410), .Z(n3405) );
  AND U3250 ( .A(\stack[1][11] ), .B(\stack[0][20] ), .Z(n3403) );
  XOR U3251 ( .A(n3411), .B(n3412), .Z(n3401) );
  XOR U3252 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U3253 ( .A(n3415), .B(n3416), .Z(n3414) );
  XOR U3254 ( .A(n3417), .B(n3418), .Z(n3416) );
  AND U3255 ( .A(n3419), .B(n3420), .Z(n3418) );
  NAND U3256 ( .A(n3421), .B(n3422), .Z(n3420) );
  NANDN U3257 ( .A(n3423), .B(n3424), .Z(n3419) );
  AND U3258 ( .A(\stack[1][15] ), .B(\stack[0][16] ), .Z(n3417) );
  XOR U3259 ( .A(n3425), .B(n3426), .Z(n3415) );
  XOR U3260 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR U3261 ( .A(n3429), .B(n3430), .Z(n3428) );
  AND U3262 ( .A(n3431), .B(n3432), .Z(n3430) );
  NAND U3263 ( .A(n3433), .B(n3434), .Z(n3432) );
  NANDN U3264 ( .A(n3435), .B(n3436), .Z(n3431) );
  AND U3265 ( .A(\stack[1][19] ), .B(\stack[0][12] ), .Z(n3429) );
  XOR U3266 ( .A(n3437), .B(n3438), .Z(n3427) );
  XOR U3267 ( .A(n3439), .B(n3440), .Z(n3438) );
  XOR U3268 ( .A(n3441), .B(n3442), .Z(n3440) );
  XOR U3269 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U3270 ( .A(n3445), .B(n3446), .Z(n3444) );
  AND U3271 ( .A(\stack[0][2] ), .B(\stack[1][29] ), .Z(n3446) );
  ANDN U3272 ( .B(n3447), .A(n3448), .Z(n3445) );
  AND U3273 ( .A(\stack[0][0] ), .B(\stack[1][30] ), .Z(n3447) );
  XOR U3274 ( .A(n3449), .B(n3450), .Z(n3443) );
  AND U3275 ( .A(n2614), .B(\stack[1][31] ), .Z(n3450) );
  IV U3276 ( .A(\stack[0][0] ), .Z(n2614) );
  AND U3277 ( .A(\stack[0][1] ), .B(\stack[1][30] ), .Z(n3449) );
  XOR U3278 ( .A(n3451), .B(n3452), .Z(n3441) );
  XOR U3279 ( .A(n3453), .B(n3454), .Z(n3452) );
  AND U3280 ( .A(n3455), .B(n3456), .Z(n3454) );
  NAND U3281 ( .A(n3457), .B(n3458), .Z(n3456) );
  NANDN U3282 ( .A(n3459), .B(n3460), .Z(n3455) );
  AND U3283 ( .A(\stack[0][4] ), .B(\stack[1][27] ), .Z(n3453) );
  XOR U3284 ( .A(n3461), .B(n3462), .Z(n3451) );
  AND U3285 ( .A(n3463), .B(n3464), .Z(n3462) );
  NAND U3286 ( .A(n3465), .B(n3466), .Z(n3464) );
  NANDN U3287 ( .A(n3467), .B(n3468), .Z(n3463) );
  OR U3288 ( .A(n3465), .B(n3466), .Z(n3468) );
  AND U3289 ( .A(\stack[0][3] ), .B(\stack[1][28] ), .Z(n3461) );
  AND U3290 ( .A(n3469), .B(n3470), .Z(n3439) );
  NAND U3291 ( .A(n3471), .B(n3472), .Z(n3470) );
  NANDN U3292 ( .A(n3473), .B(n3474), .Z(n3469) );
  XOR U3293 ( .A(n3475), .B(n3476), .Z(n3437) );
  XOR U3294 ( .A(n3477), .B(n3478), .Z(n3476) );
  AND U3295 ( .A(n3479), .B(n3480), .Z(n3478) );
  NANDN U3296 ( .A(n3481), .B(n3482), .Z(n3480) );
  NANDN U3297 ( .A(n3483), .B(n3484), .Z(n3479) );
  NANDN U3298 ( .A(n3482), .B(n3481), .Z(n3484) );
  AND U3299 ( .A(\stack[0][7] ), .B(\stack[1][24] ), .Z(n3477) );
  AND U3300 ( .A(\stack[0][8] ), .B(\stack[1][23] ), .Z(n3475) );
  XOR U3301 ( .A(n3485), .B(n3486), .Z(n3425) );
  XOR U3302 ( .A(n3487), .B(n3488), .Z(n3486) );
  AND U3303 ( .A(n3489), .B(n3490), .Z(n3488) );
  NAND U3304 ( .A(n3491), .B(n3492), .Z(n3490) );
  NANDN U3305 ( .A(n3493), .B(n3494), .Z(n3489) );
  AND U3306 ( .A(\stack[0][6] ), .B(\stack[1][25] ), .Z(n3487) );
  XOR U3307 ( .A(n3495), .B(n3496), .Z(n3485) );
  AND U3308 ( .A(n3497), .B(n3498), .Z(n3496) );
  NANDN U3309 ( .A(n3499), .B(n3500), .Z(n3498) );
  NANDN U3310 ( .A(n3501), .B(n3502), .Z(n3497) );
  NANDN U3311 ( .A(n3500), .B(n3499), .Z(n3502) );
  AND U3312 ( .A(\stack[0][5] ), .B(\stack[1][26] ), .Z(n3495) );
  XOR U3313 ( .A(n3503), .B(n3504), .Z(n3413) );
  AND U3314 ( .A(n3505), .B(n3506), .Z(n3504) );
  NANDN U3315 ( .A(n3507), .B(n3508), .Z(n3506) );
  NANDN U3316 ( .A(n3509), .B(n3510), .Z(n3505) );
  NANDN U3317 ( .A(n3508), .B(n3507), .Z(n3510) );
  AND U3318 ( .A(\stack[1][20] ), .B(\stack[0][11] ), .Z(n3503) );
  XOR U3319 ( .A(n3511), .B(n3512), .Z(n3411) );
  XOR U3320 ( .A(n3513), .B(n3514), .Z(n3512) );
  AND U3321 ( .A(n3515), .B(n3516), .Z(n3514) );
  NAND U3322 ( .A(n3517), .B(n3518), .Z(n3516) );
  NANDN U3323 ( .A(n3519), .B(n3520), .Z(n3515) );
  AND U3324 ( .A(\stack[1][21] ), .B(\stack[0][10] ), .Z(n3513) );
  XOR U3325 ( .A(n3521), .B(n3522), .Z(n3511) );
  AND U3326 ( .A(n3523), .B(n3524), .Z(n3522) );
  NANDN U3327 ( .A(n3525), .B(n3526), .Z(n3524) );
  NANDN U3328 ( .A(n3527), .B(n3528), .Z(n3523) );
  NANDN U3329 ( .A(n3526), .B(n3525), .Z(n3528) );
  AND U3330 ( .A(\stack[0][9] ), .B(\stack[1][22] ), .Z(n3521) );
  XOR U3331 ( .A(n3529), .B(n3530), .Z(n3399) );
  AND U3332 ( .A(n3531), .B(n3532), .Z(n3530) );
  NANDN U3333 ( .A(n3533), .B(n3534), .Z(n3532) );
  NANDN U3334 ( .A(n3535), .B(n3536), .Z(n3531) );
  NANDN U3335 ( .A(n3534), .B(n3533), .Z(n3536) );
  AND U3336 ( .A(\stack[1][16] ), .B(\stack[0][15] ), .Z(n3529) );
  XOR U3337 ( .A(n3537), .B(n3538), .Z(n3397) );
  XOR U3338 ( .A(n3539), .B(n3540), .Z(n3538) );
  AND U3339 ( .A(n3541), .B(n3542), .Z(n3540) );
  NAND U3340 ( .A(n3543), .B(n3544), .Z(n3542) );
  NANDN U3341 ( .A(n3545), .B(n3546), .Z(n3541) );
  AND U3342 ( .A(\stack[1][17] ), .B(\stack[0][14] ), .Z(n3539) );
  XOR U3343 ( .A(n3547), .B(n3548), .Z(n3537) );
  AND U3344 ( .A(n3549), .B(n3550), .Z(n3548) );
  NANDN U3345 ( .A(n3551), .B(n3552), .Z(n3550) );
  NANDN U3346 ( .A(n3553), .B(n3554), .Z(n3549) );
  NANDN U3347 ( .A(n3552), .B(n3551), .Z(n3554) );
  AND U3348 ( .A(\stack[1][18] ), .B(\stack[0][13] ), .Z(n3547) );
  XOR U3349 ( .A(n3555), .B(n3556), .Z(n3385) );
  AND U3350 ( .A(n3557), .B(n3558), .Z(n3556) );
  NANDN U3351 ( .A(n3559), .B(n3560), .Z(n3558) );
  NANDN U3352 ( .A(n3561), .B(n3562), .Z(n3557) );
  NANDN U3353 ( .A(n3560), .B(n3559), .Z(n3562) );
  AND U3354 ( .A(\stack[1][12] ), .B(\stack[0][19] ), .Z(n3555) );
  XOR U3355 ( .A(n3563), .B(n3564), .Z(n3383) );
  XOR U3356 ( .A(n3565), .B(n3566), .Z(n3564) );
  AND U3357 ( .A(n3567), .B(n3568), .Z(n3566) );
  NAND U3358 ( .A(n3569), .B(n3570), .Z(n3568) );
  NANDN U3359 ( .A(n3571), .B(n3572), .Z(n3567) );
  AND U3360 ( .A(\stack[1][13] ), .B(\stack[0][18] ), .Z(n3565) );
  XOR U3361 ( .A(n3573), .B(n3574), .Z(n3563) );
  AND U3362 ( .A(n3575), .B(n3576), .Z(n3574) );
  NANDN U3363 ( .A(n3577), .B(n3578), .Z(n3576) );
  NANDN U3364 ( .A(n3579), .B(n3580), .Z(n3575) );
  NANDN U3365 ( .A(n3578), .B(n3577), .Z(n3580) );
  AND U3366 ( .A(\stack[1][14] ), .B(\stack[0][17] ), .Z(n3573) );
  XOR U3367 ( .A(n3581), .B(n3582), .Z(n3371) );
  AND U3368 ( .A(n3583), .B(n3584), .Z(n3582) );
  NANDN U3369 ( .A(n3585), .B(n3586), .Z(n3584) );
  NANDN U3370 ( .A(n3587), .B(n3588), .Z(n3583) );
  NANDN U3371 ( .A(n3586), .B(n3585), .Z(n3588) );
  AND U3372 ( .A(\stack[1][8] ), .B(\stack[0][23] ), .Z(n3581) );
  XOR U3373 ( .A(n3589), .B(n3590), .Z(n3369) );
  XOR U3374 ( .A(n3591), .B(n3592), .Z(n3590) );
  AND U3375 ( .A(n3593), .B(n3594), .Z(n3592) );
  NAND U3376 ( .A(n3595), .B(n3596), .Z(n3594) );
  NANDN U3377 ( .A(n3597), .B(n3598), .Z(n3593) );
  AND U3378 ( .A(\stack[1][9] ), .B(\stack[0][22] ), .Z(n3591) );
  XOR U3379 ( .A(n3599), .B(n3600), .Z(n3589) );
  AND U3380 ( .A(n3601), .B(n3602), .Z(n3600) );
  NANDN U3381 ( .A(n3603), .B(n3604), .Z(n3602) );
  NANDN U3382 ( .A(n3605), .B(n3606), .Z(n3601) );
  NANDN U3383 ( .A(n3604), .B(n3603), .Z(n3606) );
  AND U3384 ( .A(\stack[1][10] ), .B(\stack[0][21] ), .Z(n3599) );
  XOR U3385 ( .A(n3607), .B(n3608), .Z(n3357) );
  AND U3386 ( .A(n3609), .B(n3610), .Z(n3608) );
  NANDN U3387 ( .A(n3611), .B(n3612), .Z(n3610) );
  NANDN U3388 ( .A(n3613), .B(n3614), .Z(n3609) );
  NANDN U3389 ( .A(n3612), .B(n3611), .Z(n3614) );
  AND U3390 ( .A(\stack[1][4] ), .B(\stack[0][27] ), .Z(n3607) );
  XOR U3391 ( .A(n3615), .B(n3616), .Z(n3355) );
  XOR U3392 ( .A(n3617), .B(n3618), .Z(n3616) );
  AND U3393 ( .A(n3619), .B(n3620), .Z(n3618) );
  NAND U3394 ( .A(n3621), .B(n3622), .Z(n3620) );
  NANDN U3395 ( .A(n3623), .B(n3624), .Z(n3619) );
  AND U3396 ( .A(\stack[1][5] ), .B(\stack[0][26] ), .Z(n3617) );
  XOR U3397 ( .A(n3625), .B(n3626), .Z(n3615) );
  AND U3398 ( .A(n3627), .B(n3628), .Z(n3626) );
  NANDN U3399 ( .A(n3629), .B(n3630), .Z(n3628) );
  NANDN U3400 ( .A(n3631), .B(n3632), .Z(n3627) );
  NANDN U3401 ( .A(n3630), .B(n3629), .Z(n3632) );
  AND U3402 ( .A(\stack[1][6] ), .B(\stack[0][25] ), .Z(n3625) );
  AND U3403 ( .A(n3633), .B(n3634), .Z(n3353) );
  NANDN U3404 ( .A(n3635), .B(n3636), .Z(n3634) );
  NANDN U3405 ( .A(n3637), .B(n3638), .Z(n3633) );
  XOR U3406 ( .A(n3639), .B(n3640), .Z(n3351) );
  AND U3407 ( .A(\stack[1][2] ), .B(\stack[0][29] ), .Z(n3640) );
  AND U3408 ( .A(n3641), .B(n3642), .Z(n3639) );
  NAND U3409 ( .A(n3643), .B(n3324), .Z(n3642) );
  NAND U3410 ( .A(n3644), .B(n3645), .Z(n3324) );
  NANDN U3411 ( .A(n3301), .B(n3646), .Z(n3645) );
  OR U3412 ( .A(n3300), .B(n3298), .Z(n3646) );
  AND U3413 ( .A(n3647), .B(n3648), .Z(n3301) );
  NANDN U3414 ( .A(n3275), .B(n3649), .Z(n3648) );
  NAND U3415 ( .A(n3650), .B(n3278), .Z(n3647) );
  NAND U3416 ( .A(n3651), .B(n3652), .Z(n3278) );
  NANDN U3417 ( .A(n3254), .B(n3653), .Z(n3652) );
  OR U3418 ( .A(n3253), .B(n3251), .Z(n3653) );
  AND U3419 ( .A(n3654), .B(n3655), .Z(n3254) );
  NANDN U3420 ( .A(n3227), .B(n3656), .Z(n3655) );
  NAND U3421 ( .A(n3657), .B(n3230), .Z(n3654) );
  NAND U3422 ( .A(n3658), .B(n3659), .Z(n3230) );
  NANDN U3423 ( .A(n3206), .B(n3660), .Z(n3659) );
  OR U3424 ( .A(n3205), .B(n3203), .Z(n3660) );
  AND U3425 ( .A(n3661), .B(n3662), .Z(n3206) );
  NANDN U3426 ( .A(n3179), .B(n3663), .Z(n3662) );
  NAND U3427 ( .A(n3664), .B(n3182), .Z(n3661) );
  NAND U3428 ( .A(n3665), .B(n3666), .Z(n3182) );
  NANDN U3429 ( .A(n3158), .B(n3667), .Z(n3666) );
  OR U3430 ( .A(n3157), .B(n3155), .Z(n3667) );
  AND U3431 ( .A(n3668), .B(n3669), .Z(n3158) );
  NANDN U3432 ( .A(n3131), .B(n3670), .Z(n3669) );
  NAND U3433 ( .A(n3671), .B(n3134), .Z(n3668) );
  NAND U3434 ( .A(n3672), .B(n3673), .Z(n3134) );
  NANDN U3435 ( .A(n3110), .B(n3674), .Z(n3673) );
  OR U3436 ( .A(n3109), .B(n3107), .Z(n3674) );
  AND U3437 ( .A(n3675), .B(n3676), .Z(n3110) );
  NANDN U3438 ( .A(n3083), .B(n3677), .Z(n3676) );
  NAND U3439 ( .A(n3678), .B(n3086), .Z(n3675) );
  NAND U3440 ( .A(n3679), .B(n3680), .Z(n3086) );
  NANDN U3441 ( .A(n3062), .B(n3681), .Z(n3680) );
  OR U3442 ( .A(n3061), .B(n3059), .Z(n3681) );
  AND U3443 ( .A(n3682), .B(n3683), .Z(n3062) );
  NANDN U3444 ( .A(n3035), .B(n3684), .Z(n3683) );
  NAND U3445 ( .A(n3685), .B(n3038), .Z(n3682) );
  NAND U3446 ( .A(n3686), .B(n3687), .Z(n3038) );
  NANDN U3447 ( .A(n3014), .B(n3688), .Z(n3687) );
  OR U3448 ( .A(n3013), .B(n3011), .Z(n3688) );
  AND U3449 ( .A(n3689), .B(n3690), .Z(n3014) );
  NANDN U3450 ( .A(n2987), .B(n3691), .Z(n3690) );
  NAND U3451 ( .A(n3692), .B(n2990), .Z(n3689) );
  NAND U3452 ( .A(n3693), .B(n3694), .Z(n2990) );
  NANDN U3453 ( .A(n2966), .B(n3695), .Z(n3694) );
  OR U3454 ( .A(n2965), .B(n2963), .Z(n3695) );
  AND U3455 ( .A(n3696), .B(n3697), .Z(n2966) );
  NANDN U3456 ( .A(n2939), .B(n3698), .Z(n3697) );
  NAND U3457 ( .A(n3699), .B(n2942), .Z(n3696) );
  NAND U3458 ( .A(n3700), .B(n3701), .Z(n2942) );
  NANDN U3459 ( .A(n2918), .B(n3702), .Z(n3701) );
  OR U3460 ( .A(n2917), .B(n2915), .Z(n3702) );
  AND U3461 ( .A(n3703), .B(n3704), .Z(n2918) );
  OR U3462 ( .A(n2891), .B(n2893), .Z(n3704) );
  NANDN U3463 ( .A(n2894), .B(n3705), .Z(n3703) );
  NAND U3464 ( .A(n2891), .B(n2893), .Z(n3705) );
  AND U3465 ( .A(n3706), .B(n3707), .Z(n2893) );
  OR U3466 ( .A(n2867), .B(n2869), .Z(n3707) );
  NANDN U3467 ( .A(n2870), .B(n3708), .Z(n3706) );
  NAND U3468 ( .A(n2867), .B(n2869), .Z(n3708) );
  AND U3469 ( .A(n3709), .B(n3710), .Z(n2869) );
  OR U3470 ( .A(n2843), .B(n2845), .Z(n3710) );
  NANDN U3471 ( .A(n2846), .B(n3711), .Z(n3709) );
  NAND U3472 ( .A(n2843), .B(n2845), .Z(n3711) );
  AND U3473 ( .A(n3712), .B(n3713), .Z(n2845) );
  NANDN U3474 ( .A(n2821), .B(n2819), .Z(n3713) );
  NAND U3475 ( .A(n3714), .B(n2822), .Z(n3712) );
  ANDN U3476 ( .B(\stack[0][9] ), .A(n2615), .Z(n2822) );
  AND U3477 ( .A(n3715), .B(n3716), .Z(n2821) );
  OR U3478 ( .A(n2795), .B(n2797), .Z(n3716) );
  NANDN U3479 ( .A(n2798), .B(n3717), .Z(n3715) );
  NAND U3480 ( .A(n2795), .B(n2797), .Z(n3717) );
  AND U3481 ( .A(n3718), .B(n3719), .Z(n2797) );
  OR U3482 ( .A(n2771), .B(n2773), .Z(n3719) );
  NANDN U3483 ( .A(n2774), .B(n3720), .Z(n3718) );
  NAND U3484 ( .A(n2771), .B(n2773), .Z(n3720) );
  AND U3485 ( .A(n3721), .B(n3722), .Z(n2773) );
  OR U3486 ( .A(n2747), .B(n2749), .Z(n3722) );
  NANDN U3487 ( .A(n2750), .B(n3723), .Z(n3721) );
  NAND U3488 ( .A(n2747), .B(n2749), .Z(n3723) );
  AND U3489 ( .A(n3724), .B(n3725), .Z(n2749) );
  OR U3490 ( .A(n2723), .B(n2725), .Z(n3725) );
  NANDN U3491 ( .A(n2726), .B(n3726), .Z(n3724) );
  NAND U3492 ( .A(n2723), .B(n2725), .Z(n3726) );
  AND U3493 ( .A(n3727), .B(n3728), .Z(n2725) );
  OR U3494 ( .A(n2699), .B(n2701), .Z(n3728) );
  NANDN U3495 ( .A(n2702), .B(n3729), .Z(n3727) );
  NAND U3496 ( .A(n2699), .B(n2701), .Z(n3729) );
  AND U3497 ( .A(n3730), .B(n3731), .Z(n2701) );
  NANDN U3498 ( .A(n2675), .B(n2677), .Z(n3731) );
  NANDN U3499 ( .A(n2678), .B(n3732), .Z(n3730) );
  NANDN U3500 ( .A(n2677), .B(n2675), .Z(n3732) );
  XNOR U3501 ( .A(n3733), .B(n3734), .Z(n2675) );
  XNOR U3502 ( .A(n3735), .B(n3736), .Z(n3734) );
  AND U3503 ( .A(\stack[1][0] ), .B(\stack[0][3] ), .Z(n2677) );
  AND U3504 ( .A(n3737), .B(n3738), .Z(n2678) );
  NANDN U3505 ( .A(n2652), .B(n2654), .Z(n3738) );
  NANDN U3506 ( .A(n2655), .B(n3739), .Z(n3737) );
  NANDN U3507 ( .A(n2654), .B(n2652), .Z(n3739) );
  XNOR U3508 ( .A(n3740), .B(n3741), .Z(n2652) );
  NAND U3509 ( .A(\stack[0][0] ), .B(\stack[1][2] ), .Z(n3741) );
  NOR U3510 ( .A(n2631), .B(n2632), .Z(n2654) );
  NAND U3511 ( .A(\stack[1][0] ), .B(\stack[0][1] ), .Z(n2632) );
  NAND U3512 ( .A(\stack[1][1] ), .B(\stack[0][0] ), .Z(n2631) );
  NAND U3513 ( .A(\stack[1][0] ), .B(\stack[0][2] ), .Z(n2655) );
  XOR U3514 ( .A(n3742), .B(n3743), .Z(n2699) );
  XNOR U3515 ( .A(n3744), .B(n3745), .Z(n3743) );
  NAND U3516 ( .A(\stack[1][0] ), .B(\stack[0][4] ), .Z(n2702) );
  XOR U3517 ( .A(n3746), .B(n3747), .Z(n2723) );
  XOR U3518 ( .A(n3748), .B(n3749), .Z(n3747) );
  NAND U3519 ( .A(\stack[0][5] ), .B(\stack[1][0] ), .Z(n2726) );
  XOR U3520 ( .A(n3750), .B(n3751), .Z(n2747) );
  XNOR U3521 ( .A(n3752), .B(n3753), .Z(n3751) );
  NAND U3522 ( .A(\stack[1][0] ), .B(\stack[0][6] ), .Z(n2750) );
  XOR U3523 ( .A(n3754), .B(n3755), .Z(n2771) );
  XOR U3524 ( .A(n3756), .B(n3757), .Z(n3755) );
  NAND U3525 ( .A(\stack[0][7] ), .B(\stack[1][0] ), .Z(n2774) );
  XOR U3526 ( .A(n3758), .B(n3759), .Z(n2795) );
  XNOR U3527 ( .A(n3760), .B(n3761), .Z(n3759) );
  NAND U3528 ( .A(\stack[1][0] ), .B(\stack[0][8] ), .Z(n2798) );
  XOR U3529 ( .A(n3762), .B(n3763), .Z(n2819) );
  XNOR U3530 ( .A(n3764), .B(n3765), .Z(n3763) );
  XOR U3531 ( .A(n3766), .B(n3767), .Z(n2843) );
  XNOR U3532 ( .A(n3768), .B(n3769), .Z(n3767) );
  NAND U3533 ( .A(\stack[0][10] ), .B(\stack[1][0] ), .Z(n2846) );
  XOR U3534 ( .A(n3770), .B(n3771), .Z(n2867) );
  XOR U3535 ( .A(n3772), .B(n3773), .Z(n3771) );
  NAND U3536 ( .A(\stack[1][0] ), .B(\stack[0][11] ), .Z(n2870) );
  XOR U3537 ( .A(n3774), .B(n3775), .Z(n2891) );
  XNOR U3538 ( .A(n3776), .B(n3777), .Z(n3775) );
  NAND U3539 ( .A(\stack[0][12] ), .B(\stack[1][0] ), .Z(n2894) );
  NAND U3540 ( .A(n2915), .B(n2917), .Z(n3700) );
  ANDN U3541 ( .B(\stack[1][0] ), .A(n2923), .Z(n2917) );
  XNOR U3542 ( .A(n3778), .B(n3779), .Z(n2915) );
  XOR U3543 ( .A(n3780), .B(n3781), .Z(n3779) );
  NAND U3544 ( .A(n2941), .B(n2939), .Z(n3699) );
  XOR U3545 ( .A(n3782), .B(n3783), .Z(n2939) );
  XNOR U3546 ( .A(n3784), .B(n3785), .Z(n3783) );
  IV U3547 ( .A(n3698), .Z(n2941) );
  NOR U3548 ( .A(n2947), .B(n2615), .Z(n3698) );
  NAND U3549 ( .A(n2963), .B(n2965), .Z(n3693) );
  ANDN U3550 ( .B(\stack[1][0] ), .A(n2971), .Z(n2965) );
  XNOR U3551 ( .A(n3786), .B(n3787), .Z(n2963) );
  XOR U3552 ( .A(n3788), .B(n3789), .Z(n3787) );
  NAND U3553 ( .A(n2989), .B(n2987), .Z(n3692) );
  XOR U3554 ( .A(n3790), .B(n3791), .Z(n2987) );
  XNOR U3555 ( .A(n3792), .B(n3793), .Z(n3791) );
  IV U3556 ( .A(n3691), .Z(n2989) );
  NOR U3557 ( .A(n2995), .B(n2615), .Z(n3691) );
  NAND U3558 ( .A(n3011), .B(n3013), .Z(n3686) );
  ANDN U3559 ( .B(\stack[1][0] ), .A(n3019), .Z(n3013) );
  XNOR U3560 ( .A(n3794), .B(n3795), .Z(n3011) );
  XOR U3561 ( .A(n3796), .B(n3797), .Z(n3795) );
  NAND U3562 ( .A(n3037), .B(n3035), .Z(n3685) );
  XOR U3563 ( .A(n3798), .B(n3799), .Z(n3035) );
  XNOR U3564 ( .A(n3800), .B(n3801), .Z(n3799) );
  IV U3565 ( .A(n3684), .Z(n3037) );
  NOR U3566 ( .A(n3043), .B(n2615), .Z(n3684) );
  NAND U3567 ( .A(n3059), .B(n3061), .Z(n3679) );
  ANDN U3568 ( .B(\stack[1][0] ), .A(n3067), .Z(n3061) );
  XNOR U3569 ( .A(n3802), .B(n3803), .Z(n3059) );
  XOR U3570 ( .A(n3804), .B(n3805), .Z(n3803) );
  NAND U3571 ( .A(n3085), .B(n3083), .Z(n3678) );
  XOR U3572 ( .A(n3806), .B(n3807), .Z(n3083) );
  XNOR U3573 ( .A(n3808), .B(n3809), .Z(n3807) );
  IV U3574 ( .A(n3677), .Z(n3085) );
  NOR U3575 ( .A(n3091), .B(n2615), .Z(n3677) );
  NAND U3576 ( .A(n3107), .B(n3109), .Z(n3672) );
  ANDN U3577 ( .B(\stack[1][0] ), .A(n3115), .Z(n3109) );
  XNOR U3578 ( .A(n3810), .B(n3811), .Z(n3107) );
  XOR U3579 ( .A(n3812), .B(n3813), .Z(n3811) );
  NAND U3580 ( .A(n3133), .B(n3131), .Z(n3671) );
  XOR U3581 ( .A(n3814), .B(n3815), .Z(n3131) );
  XNOR U3582 ( .A(n3816), .B(n3817), .Z(n3815) );
  IV U3583 ( .A(n3670), .Z(n3133) );
  NOR U3584 ( .A(n3139), .B(n2615), .Z(n3670) );
  NAND U3585 ( .A(n3155), .B(n3157), .Z(n3665) );
  ANDN U3586 ( .B(\stack[1][0] ), .A(n3163), .Z(n3157) );
  XNOR U3587 ( .A(n3818), .B(n3819), .Z(n3155) );
  XOR U3588 ( .A(n3820), .B(n3821), .Z(n3819) );
  NAND U3589 ( .A(n3181), .B(n3179), .Z(n3664) );
  XOR U3590 ( .A(n3822), .B(n3823), .Z(n3179) );
  XNOR U3591 ( .A(n3824), .B(n3825), .Z(n3823) );
  IV U3592 ( .A(n3663), .Z(n3181) );
  NOR U3593 ( .A(n3187), .B(n2615), .Z(n3663) );
  NAND U3594 ( .A(n3203), .B(n3205), .Z(n3658) );
  ANDN U3595 ( .B(\stack[1][0] ), .A(n3211), .Z(n3205) );
  XNOR U3596 ( .A(n3826), .B(n3827), .Z(n3203) );
  XOR U3597 ( .A(n3828), .B(n3829), .Z(n3827) );
  NAND U3598 ( .A(n3229), .B(n3227), .Z(n3657) );
  XOR U3599 ( .A(n3830), .B(n3831), .Z(n3227) );
  XNOR U3600 ( .A(n3832), .B(n3833), .Z(n3831) );
  IV U3601 ( .A(n3656), .Z(n3229) );
  NOR U3602 ( .A(n3235), .B(n2615), .Z(n3656) );
  NAND U3603 ( .A(n3251), .B(n3253), .Z(n3651) );
  ANDN U3604 ( .B(\stack[1][0] ), .A(n3259), .Z(n3253) );
  XNOR U3605 ( .A(n3834), .B(n3835), .Z(n3251) );
  XOR U3606 ( .A(n3836), .B(n3837), .Z(n3835) );
  NAND U3607 ( .A(n3277), .B(n3275), .Z(n3650) );
  XOR U3608 ( .A(n3838), .B(n3839), .Z(n3275) );
  XNOR U3609 ( .A(n3840), .B(n3841), .Z(n3839) );
  IV U3610 ( .A(n3649), .Z(n3277) );
  NOR U3611 ( .A(n3283), .B(n2615), .Z(n3649) );
  NAND U3612 ( .A(n3298), .B(n3300), .Z(n3644) );
  ANDN U3613 ( .B(\stack[1][0] ), .A(n3306), .Z(n3300) );
  XNOR U3614 ( .A(n3842), .B(n3843), .Z(n3298) );
  XOR U3615 ( .A(n3844), .B(n3845), .Z(n3843) );
  NANDN U3616 ( .A(n3323), .B(n3321), .Z(n3643) );
  AND U3617 ( .A(n3846), .B(n3847), .Z(n3641) );
  NAND U3618 ( .A(\stack[0][31] ), .B(n2615), .Z(n3847) );
  IV U3619 ( .A(\stack[1][0] ), .Z(n2615) );
  NANDN U3620 ( .A(n3321), .B(n3323), .Z(n3846) );
  XNOR U3621 ( .A(n3366), .B(n3848), .Z(n3321) );
  XNOR U3622 ( .A(n3365), .B(n3367), .Z(n3848) );
  AND U3623 ( .A(n3849), .B(n3850), .Z(n3367) );
  NANDN U3624 ( .A(n3842), .B(n3851), .Z(n3850) );
  NANDN U3625 ( .A(n3845), .B(n3852), .Z(n3849) );
  NAND U3626 ( .A(n3844), .B(n3842), .Z(n3852) );
  XOR U3627 ( .A(n3853), .B(n3854), .Z(n3842) );
  XNOR U3628 ( .A(n3855), .B(n3856), .Z(n3854) );
  IV U3629 ( .A(n3851), .Z(n3844) );
  NOR U3630 ( .A(n3283), .B(n2637), .Z(n3851) );
  AND U3631 ( .A(n3857), .B(n3858), .Z(n3845) );
  NANDN U3632 ( .A(n3838), .B(n3840), .Z(n3858) );
  NANDN U3633 ( .A(n3841), .B(n3859), .Z(n3857) );
  NANDN U3634 ( .A(n3840), .B(n3838), .Z(n3859) );
  XOR U3635 ( .A(n3860), .B(n3861), .Z(n3838) );
  XOR U3636 ( .A(n3862), .B(n3863), .Z(n3861) );
  AND U3637 ( .A(\stack[0][27] ), .B(\stack[1][1] ), .Z(n3840) );
  AND U3638 ( .A(n3864), .B(n3865), .Z(n3841) );
  NANDN U3639 ( .A(n3834), .B(n3866), .Z(n3865) );
  NANDN U3640 ( .A(n3837), .B(n3867), .Z(n3864) );
  NAND U3641 ( .A(n3836), .B(n3834), .Z(n3867) );
  XOR U3642 ( .A(n3868), .B(n3869), .Z(n3834) );
  XNOR U3643 ( .A(n3870), .B(n3871), .Z(n3869) );
  IV U3644 ( .A(n3866), .Z(n3836) );
  NOR U3645 ( .A(n3235), .B(n2637), .Z(n3866) );
  AND U3646 ( .A(n3872), .B(n3873), .Z(n3837) );
  NANDN U3647 ( .A(n3830), .B(n3832), .Z(n3873) );
  NANDN U3648 ( .A(n3833), .B(n3874), .Z(n3872) );
  NANDN U3649 ( .A(n3832), .B(n3830), .Z(n3874) );
  XOR U3650 ( .A(n3875), .B(n3876), .Z(n3830) );
  XOR U3651 ( .A(n3877), .B(n3878), .Z(n3876) );
  AND U3652 ( .A(\stack[0][25] ), .B(\stack[1][1] ), .Z(n3832) );
  AND U3653 ( .A(n3879), .B(n3880), .Z(n3833) );
  NANDN U3654 ( .A(n3826), .B(n3881), .Z(n3880) );
  NANDN U3655 ( .A(n3829), .B(n3882), .Z(n3879) );
  NAND U3656 ( .A(n3828), .B(n3826), .Z(n3882) );
  XOR U3657 ( .A(n3883), .B(n3884), .Z(n3826) );
  XNOR U3658 ( .A(n3885), .B(n3886), .Z(n3884) );
  IV U3659 ( .A(n3881), .Z(n3828) );
  NOR U3660 ( .A(n3187), .B(n2637), .Z(n3881) );
  AND U3661 ( .A(n3887), .B(n3888), .Z(n3829) );
  NANDN U3662 ( .A(n3822), .B(n3824), .Z(n3888) );
  NANDN U3663 ( .A(n3825), .B(n3889), .Z(n3887) );
  NANDN U3664 ( .A(n3824), .B(n3822), .Z(n3889) );
  XOR U3665 ( .A(n3890), .B(n3891), .Z(n3822) );
  XOR U3666 ( .A(n3892), .B(n3893), .Z(n3891) );
  AND U3667 ( .A(\stack[0][23] ), .B(\stack[1][1] ), .Z(n3824) );
  AND U3668 ( .A(n3894), .B(n3895), .Z(n3825) );
  NANDN U3669 ( .A(n3818), .B(n3896), .Z(n3895) );
  NANDN U3670 ( .A(n3821), .B(n3897), .Z(n3894) );
  NAND U3671 ( .A(n3820), .B(n3818), .Z(n3897) );
  XOR U3672 ( .A(n3898), .B(n3899), .Z(n3818) );
  XNOR U3673 ( .A(n3900), .B(n3901), .Z(n3899) );
  IV U3674 ( .A(n3896), .Z(n3820) );
  NOR U3675 ( .A(n3139), .B(n2637), .Z(n3896) );
  AND U3676 ( .A(n3902), .B(n3903), .Z(n3821) );
  NANDN U3677 ( .A(n3814), .B(n3816), .Z(n3903) );
  NANDN U3678 ( .A(n3817), .B(n3904), .Z(n3902) );
  NANDN U3679 ( .A(n3816), .B(n3814), .Z(n3904) );
  XOR U3680 ( .A(n3905), .B(n3906), .Z(n3814) );
  XOR U3681 ( .A(n3907), .B(n3908), .Z(n3906) );
  AND U3682 ( .A(\stack[0][21] ), .B(\stack[1][1] ), .Z(n3816) );
  AND U3683 ( .A(n3909), .B(n3910), .Z(n3817) );
  NANDN U3684 ( .A(n3810), .B(n3911), .Z(n3910) );
  NANDN U3685 ( .A(n3813), .B(n3912), .Z(n3909) );
  NAND U3686 ( .A(n3812), .B(n3810), .Z(n3912) );
  XOR U3687 ( .A(n3913), .B(n3914), .Z(n3810) );
  XNOR U3688 ( .A(n3915), .B(n3916), .Z(n3914) );
  IV U3689 ( .A(n3911), .Z(n3812) );
  NOR U3690 ( .A(n3091), .B(n2637), .Z(n3911) );
  AND U3691 ( .A(n3917), .B(n3918), .Z(n3813) );
  NANDN U3692 ( .A(n3806), .B(n3808), .Z(n3918) );
  NANDN U3693 ( .A(n3809), .B(n3919), .Z(n3917) );
  NANDN U3694 ( .A(n3808), .B(n3806), .Z(n3919) );
  XOR U3695 ( .A(n3920), .B(n3921), .Z(n3806) );
  XOR U3696 ( .A(n3922), .B(n3923), .Z(n3921) );
  AND U3697 ( .A(\stack[0][19] ), .B(\stack[1][1] ), .Z(n3808) );
  AND U3698 ( .A(n3924), .B(n3925), .Z(n3809) );
  NANDN U3699 ( .A(n3802), .B(n3926), .Z(n3925) );
  NANDN U3700 ( .A(n3805), .B(n3927), .Z(n3924) );
  NAND U3701 ( .A(n3804), .B(n3802), .Z(n3927) );
  XOR U3702 ( .A(n3928), .B(n3929), .Z(n3802) );
  XNOR U3703 ( .A(n3930), .B(n3931), .Z(n3929) );
  IV U3704 ( .A(n3926), .Z(n3804) );
  NOR U3705 ( .A(n3043), .B(n2637), .Z(n3926) );
  AND U3706 ( .A(n3932), .B(n3933), .Z(n3805) );
  NANDN U3707 ( .A(n3798), .B(n3800), .Z(n3933) );
  NANDN U3708 ( .A(n3801), .B(n3934), .Z(n3932) );
  NANDN U3709 ( .A(n3800), .B(n3798), .Z(n3934) );
  XOR U3710 ( .A(n3935), .B(n3936), .Z(n3798) );
  XOR U3711 ( .A(n3937), .B(n3938), .Z(n3936) );
  AND U3712 ( .A(\stack[0][17] ), .B(\stack[1][1] ), .Z(n3800) );
  AND U3713 ( .A(n3939), .B(n3940), .Z(n3801) );
  NANDN U3714 ( .A(n3794), .B(n3941), .Z(n3940) );
  NANDN U3715 ( .A(n3797), .B(n3942), .Z(n3939) );
  NAND U3716 ( .A(n3796), .B(n3794), .Z(n3942) );
  XOR U3717 ( .A(n3943), .B(n3944), .Z(n3794) );
  XNOR U3718 ( .A(n3945), .B(n3946), .Z(n3944) );
  IV U3719 ( .A(n3941), .Z(n3796) );
  NOR U3720 ( .A(n2995), .B(n2637), .Z(n3941) );
  AND U3721 ( .A(n3947), .B(n3948), .Z(n3797) );
  NANDN U3722 ( .A(n3790), .B(n3792), .Z(n3948) );
  NANDN U3723 ( .A(n3793), .B(n3949), .Z(n3947) );
  NANDN U3724 ( .A(n3792), .B(n3790), .Z(n3949) );
  XOR U3725 ( .A(n3950), .B(n3951), .Z(n3790) );
  XOR U3726 ( .A(n3952), .B(n3953), .Z(n3951) );
  AND U3727 ( .A(\stack[0][15] ), .B(\stack[1][1] ), .Z(n3792) );
  AND U3728 ( .A(n3954), .B(n3955), .Z(n3793) );
  NANDN U3729 ( .A(n3786), .B(n3956), .Z(n3955) );
  NANDN U3730 ( .A(n3789), .B(n3957), .Z(n3954) );
  NAND U3731 ( .A(n3788), .B(n3786), .Z(n3957) );
  XOR U3732 ( .A(n3958), .B(n3959), .Z(n3786) );
  XNOR U3733 ( .A(n3960), .B(n3961), .Z(n3959) );
  IV U3734 ( .A(n3956), .Z(n3788) );
  NOR U3735 ( .A(n2947), .B(n2637), .Z(n3956) );
  AND U3736 ( .A(n3962), .B(n3963), .Z(n3789) );
  NANDN U3737 ( .A(n3782), .B(n3784), .Z(n3963) );
  NANDN U3738 ( .A(n3785), .B(n3964), .Z(n3962) );
  NANDN U3739 ( .A(n3784), .B(n3782), .Z(n3964) );
  XOR U3740 ( .A(n3965), .B(n3966), .Z(n3782) );
  XOR U3741 ( .A(n3967), .B(n3968), .Z(n3966) );
  AND U3742 ( .A(\stack[0][13] ), .B(\stack[1][1] ), .Z(n3784) );
  AND U3743 ( .A(n3969), .B(n3970), .Z(n3785) );
  NANDN U3744 ( .A(n3778), .B(n3971), .Z(n3970) );
  NANDN U3745 ( .A(n3781), .B(n3972), .Z(n3969) );
  NAND U3746 ( .A(n3780), .B(n3778), .Z(n3972) );
  XOR U3747 ( .A(n3973), .B(n3974), .Z(n3778) );
  XNOR U3748 ( .A(n3975), .B(n3976), .Z(n3974) );
  IV U3749 ( .A(n3971), .Z(n3780) );
  NOR U3750 ( .A(n2899), .B(n2637), .Z(n3971) );
  AND U3751 ( .A(n3977), .B(n3978), .Z(n3781) );
  NANDN U3752 ( .A(n3774), .B(n3776), .Z(n3978) );
  NANDN U3753 ( .A(n3777), .B(n3979), .Z(n3977) );
  NANDN U3754 ( .A(n3776), .B(n3774), .Z(n3979) );
  XOR U3755 ( .A(n3980), .B(n3981), .Z(n3774) );
  XOR U3756 ( .A(n3982), .B(n3983), .Z(n3981) );
  AND U3757 ( .A(\stack[0][11] ), .B(\stack[1][1] ), .Z(n3776) );
  AND U3758 ( .A(n3984), .B(n3985), .Z(n3777) );
  NANDN U3759 ( .A(n3770), .B(n3986), .Z(n3985) );
  NANDN U3760 ( .A(n3773), .B(n3987), .Z(n3984) );
  NAND U3761 ( .A(n3772), .B(n3770), .Z(n3987) );
  XOR U3762 ( .A(n3988), .B(n3989), .Z(n3770) );
  XNOR U3763 ( .A(n3990), .B(n3991), .Z(n3989) );
  IV U3764 ( .A(n3986), .Z(n3772) );
  NOR U3765 ( .A(n2851), .B(n2637), .Z(n3986) );
  AND U3766 ( .A(n3992), .B(n3993), .Z(n3773) );
  NANDN U3767 ( .A(n3766), .B(n3768), .Z(n3993) );
  NANDN U3768 ( .A(n3769), .B(n3994), .Z(n3992) );
  NANDN U3769 ( .A(n3768), .B(n3766), .Z(n3994) );
  XOR U3770 ( .A(n3995), .B(n3996), .Z(n3766) );
  XOR U3771 ( .A(n3997), .B(n3998), .Z(n3996) );
  AND U3772 ( .A(\stack[1][1] ), .B(\stack[0][9] ), .Z(n3768) );
  AND U3773 ( .A(n3999), .B(n4000), .Z(n3769) );
  NAND U3774 ( .A(n3762), .B(n3764), .Z(n4000) );
  IV U3775 ( .A(n4001), .Z(n3762) );
  NANDN U3776 ( .A(n3765), .B(n4002), .Z(n3999) );
  NANDN U3777 ( .A(n3764), .B(n4001), .Z(n4002) );
  XNOR U3778 ( .A(n4003), .B(n4004), .Z(n4001) );
  XNOR U3779 ( .A(n4005), .B(n4006), .Z(n4004) );
  ANDN U3780 ( .B(\stack[0][8] ), .A(n2637), .Z(n3764) );
  AND U3781 ( .A(n4007), .B(n4008), .Z(n3765) );
  NANDN U3782 ( .A(n3758), .B(n3760), .Z(n4008) );
  NANDN U3783 ( .A(n3761), .B(n4009), .Z(n4007) );
  NANDN U3784 ( .A(n3760), .B(n3758), .Z(n4009) );
  XOR U3785 ( .A(n4010), .B(n4011), .Z(n3758) );
  XOR U3786 ( .A(n4012), .B(n4013), .Z(n4011) );
  AND U3787 ( .A(\stack[1][1] ), .B(\stack[0][7] ), .Z(n3760) );
  AND U3788 ( .A(n4014), .B(n4015), .Z(n3761) );
  NANDN U3789 ( .A(n3754), .B(n4016), .Z(n4015) );
  NANDN U3790 ( .A(n3757), .B(n4017), .Z(n4014) );
  NAND U3791 ( .A(n3756), .B(n3754), .Z(n4017) );
  XOR U3792 ( .A(n4018), .B(n4019), .Z(n3754) );
  XNOR U3793 ( .A(n4020), .B(n4021), .Z(n4019) );
  IV U3794 ( .A(n4016), .Z(n3756) );
  NOR U3795 ( .A(n2637), .B(n2755), .Z(n4016) );
  AND U3796 ( .A(n4022), .B(n4023), .Z(n3757) );
  NANDN U3797 ( .A(n3750), .B(n3752), .Z(n4023) );
  NANDN U3798 ( .A(n3753), .B(n4024), .Z(n4022) );
  NANDN U3799 ( .A(n3752), .B(n3750), .Z(n4024) );
  XOR U3800 ( .A(n4025), .B(n4026), .Z(n3750) );
  XOR U3801 ( .A(n4027), .B(n4028), .Z(n4026) );
  AND U3802 ( .A(\stack[1][1] ), .B(\stack[0][5] ), .Z(n3752) );
  AND U3803 ( .A(n4029), .B(n4030), .Z(n3753) );
  NANDN U3804 ( .A(n3746), .B(n4031), .Z(n4030) );
  NANDN U3805 ( .A(n3749), .B(n4032), .Z(n4029) );
  NAND U3806 ( .A(n3748), .B(n3746), .Z(n4032) );
  XOR U3807 ( .A(n4033), .B(n4034), .Z(n3746) );
  XNOR U3808 ( .A(n4035), .B(n4036), .Z(n4034) );
  IV U3809 ( .A(n4031), .Z(n3748) );
  NOR U3810 ( .A(n2637), .B(n2707), .Z(n4031) );
  AND U3811 ( .A(n4037), .B(n4038), .Z(n3749) );
  NANDN U3812 ( .A(n3742), .B(n3744), .Z(n4038) );
  NANDN U3813 ( .A(n3745), .B(n4039), .Z(n4037) );
  NANDN U3814 ( .A(n3744), .B(n3742), .Z(n4039) );
  XNOR U3815 ( .A(n4040), .B(n4041), .Z(n3742) );
  XNOR U3816 ( .A(n4042), .B(n4043), .Z(n4041) );
  AND U3817 ( .A(\stack[1][1] ), .B(\stack[0][3] ), .Z(n3744) );
  AND U3818 ( .A(n4044), .B(n4045), .Z(n3745) );
  NANDN U3819 ( .A(n3733), .B(n3735), .Z(n4045) );
  NAND U3820 ( .A(n4046), .B(n3736), .Z(n4044) );
  ANDN U3821 ( .B(n4047), .A(n3740), .Z(n3736) );
  NAND U3822 ( .A(\stack[1][1] ), .B(\stack[0][1] ), .Z(n3740) );
  AND U3823 ( .A(\stack[0][0] ), .B(\stack[1][2] ), .Z(n4047) );
  NANDN U3824 ( .A(n3735), .B(n3733), .Z(n4046) );
  XNOR U3825 ( .A(n4048), .B(n4049), .Z(n3733) );
  NAND U3826 ( .A(\stack[0][0] ), .B(\stack[1][3] ), .Z(n4049) );
  AND U3827 ( .A(\stack[1][1] ), .B(\stack[0][2] ), .Z(n3735) );
  NOR U3828 ( .A(n3306), .B(n2637), .Z(n3365) );
  IV U3829 ( .A(\stack[1][1] ), .Z(n2637) );
  IV U3830 ( .A(\stack[0][29] ), .Z(n3306) );
  XNOR U3831 ( .A(n3635), .B(n4050), .Z(n3366) );
  XNOR U3832 ( .A(n3636), .B(n3637), .Z(n4050) );
  AND U3833 ( .A(n4051), .B(n4052), .Z(n3637) );
  NANDN U3834 ( .A(n3853), .B(n3855), .Z(n4052) );
  NANDN U3835 ( .A(n3856), .B(n4053), .Z(n4051) );
  NANDN U3836 ( .A(n3855), .B(n3853), .Z(n4053) );
  XOR U3837 ( .A(n4054), .B(n4055), .Z(n3853) );
  XOR U3838 ( .A(n4056), .B(n4057), .Z(n4055) );
  AND U3839 ( .A(\stack[0][27] ), .B(\stack[1][2] ), .Z(n3855) );
  AND U3840 ( .A(n4058), .B(n4059), .Z(n3856) );
  NANDN U3841 ( .A(n3860), .B(n4060), .Z(n4059) );
  NANDN U3842 ( .A(n3863), .B(n4061), .Z(n4058) );
  NAND U3843 ( .A(n3862), .B(n3860), .Z(n4061) );
  XOR U3844 ( .A(n4062), .B(n4063), .Z(n3860) );
  XNOR U3845 ( .A(n4064), .B(n4065), .Z(n4063) );
  IV U3846 ( .A(n4060), .Z(n3862) );
  NOR U3847 ( .A(n3235), .B(n2660), .Z(n4060) );
  AND U3848 ( .A(n4066), .B(n4067), .Z(n3863) );
  NANDN U3849 ( .A(n3868), .B(n3870), .Z(n4067) );
  NANDN U3850 ( .A(n3871), .B(n4068), .Z(n4066) );
  NANDN U3851 ( .A(n3870), .B(n3868), .Z(n4068) );
  XOR U3852 ( .A(n4069), .B(n4070), .Z(n3868) );
  XOR U3853 ( .A(n4071), .B(n4072), .Z(n4070) );
  AND U3854 ( .A(\stack[0][25] ), .B(\stack[1][2] ), .Z(n3870) );
  AND U3855 ( .A(n4073), .B(n4074), .Z(n3871) );
  NANDN U3856 ( .A(n3875), .B(n4075), .Z(n4074) );
  NANDN U3857 ( .A(n3878), .B(n4076), .Z(n4073) );
  NAND U3858 ( .A(n3877), .B(n3875), .Z(n4076) );
  XOR U3859 ( .A(n4077), .B(n4078), .Z(n3875) );
  XNOR U3860 ( .A(n4079), .B(n4080), .Z(n4078) );
  IV U3861 ( .A(n4075), .Z(n3877) );
  NOR U3862 ( .A(n3187), .B(n2660), .Z(n4075) );
  AND U3863 ( .A(n4081), .B(n4082), .Z(n3878) );
  NANDN U3864 ( .A(n3883), .B(n3885), .Z(n4082) );
  NANDN U3865 ( .A(n3886), .B(n4083), .Z(n4081) );
  NANDN U3866 ( .A(n3885), .B(n3883), .Z(n4083) );
  XOR U3867 ( .A(n4084), .B(n4085), .Z(n3883) );
  XOR U3868 ( .A(n4086), .B(n4087), .Z(n4085) );
  AND U3869 ( .A(\stack[0][23] ), .B(\stack[1][2] ), .Z(n3885) );
  AND U3870 ( .A(n4088), .B(n4089), .Z(n3886) );
  NANDN U3871 ( .A(n3890), .B(n4090), .Z(n4089) );
  NANDN U3872 ( .A(n3893), .B(n4091), .Z(n4088) );
  NAND U3873 ( .A(n3892), .B(n3890), .Z(n4091) );
  XOR U3874 ( .A(n4092), .B(n4093), .Z(n3890) );
  XNOR U3875 ( .A(n4094), .B(n4095), .Z(n4093) );
  IV U3876 ( .A(n4090), .Z(n3892) );
  NOR U3877 ( .A(n3139), .B(n2660), .Z(n4090) );
  AND U3878 ( .A(n4096), .B(n4097), .Z(n3893) );
  NANDN U3879 ( .A(n3898), .B(n3900), .Z(n4097) );
  NANDN U3880 ( .A(n3901), .B(n4098), .Z(n4096) );
  NANDN U3881 ( .A(n3900), .B(n3898), .Z(n4098) );
  XOR U3882 ( .A(n4099), .B(n4100), .Z(n3898) );
  XOR U3883 ( .A(n4101), .B(n4102), .Z(n4100) );
  AND U3884 ( .A(\stack[0][21] ), .B(\stack[1][2] ), .Z(n3900) );
  AND U3885 ( .A(n4103), .B(n4104), .Z(n3901) );
  NANDN U3886 ( .A(n3905), .B(n4105), .Z(n4104) );
  NANDN U3887 ( .A(n3908), .B(n4106), .Z(n4103) );
  NAND U3888 ( .A(n3907), .B(n3905), .Z(n4106) );
  XOR U3889 ( .A(n4107), .B(n4108), .Z(n3905) );
  XNOR U3890 ( .A(n4109), .B(n4110), .Z(n4108) );
  IV U3891 ( .A(n4105), .Z(n3907) );
  NOR U3892 ( .A(n3091), .B(n2660), .Z(n4105) );
  AND U3893 ( .A(n4111), .B(n4112), .Z(n3908) );
  NANDN U3894 ( .A(n3913), .B(n3915), .Z(n4112) );
  NANDN U3895 ( .A(n3916), .B(n4113), .Z(n4111) );
  NANDN U3896 ( .A(n3915), .B(n3913), .Z(n4113) );
  XOR U3897 ( .A(n4114), .B(n4115), .Z(n3913) );
  XOR U3898 ( .A(n4116), .B(n4117), .Z(n4115) );
  AND U3899 ( .A(\stack[0][19] ), .B(\stack[1][2] ), .Z(n3915) );
  AND U3900 ( .A(n4118), .B(n4119), .Z(n3916) );
  NANDN U3901 ( .A(n3920), .B(n4120), .Z(n4119) );
  NANDN U3902 ( .A(n3923), .B(n4121), .Z(n4118) );
  NAND U3903 ( .A(n3922), .B(n3920), .Z(n4121) );
  XOR U3904 ( .A(n4122), .B(n4123), .Z(n3920) );
  XNOR U3905 ( .A(n4124), .B(n4125), .Z(n4123) );
  IV U3906 ( .A(n4120), .Z(n3922) );
  NOR U3907 ( .A(n3043), .B(n2660), .Z(n4120) );
  AND U3908 ( .A(n4126), .B(n4127), .Z(n3923) );
  NANDN U3909 ( .A(n3928), .B(n3930), .Z(n4127) );
  NANDN U3910 ( .A(n3931), .B(n4128), .Z(n4126) );
  NANDN U3911 ( .A(n3930), .B(n3928), .Z(n4128) );
  XOR U3912 ( .A(n4129), .B(n4130), .Z(n3928) );
  XOR U3913 ( .A(n4131), .B(n4132), .Z(n4130) );
  AND U3914 ( .A(\stack[0][17] ), .B(\stack[1][2] ), .Z(n3930) );
  AND U3915 ( .A(n4133), .B(n4134), .Z(n3931) );
  NANDN U3916 ( .A(n3935), .B(n4135), .Z(n4134) );
  NANDN U3917 ( .A(n3938), .B(n4136), .Z(n4133) );
  NAND U3918 ( .A(n3937), .B(n3935), .Z(n4136) );
  XOR U3919 ( .A(n4137), .B(n4138), .Z(n3935) );
  XNOR U3920 ( .A(n4139), .B(n4140), .Z(n4138) );
  IV U3921 ( .A(n4135), .Z(n3937) );
  NOR U3922 ( .A(n2995), .B(n2660), .Z(n4135) );
  AND U3923 ( .A(n4141), .B(n4142), .Z(n3938) );
  NANDN U3924 ( .A(n3943), .B(n3945), .Z(n4142) );
  NANDN U3925 ( .A(n3946), .B(n4143), .Z(n4141) );
  NANDN U3926 ( .A(n3945), .B(n3943), .Z(n4143) );
  XOR U3927 ( .A(n4144), .B(n4145), .Z(n3943) );
  XOR U3928 ( .A(n4146), .B(n4147), .Z(n4145) );
  AND U3929 ( .A(\stack[0][15] ), .B(\stack[1][2] ), .Z(n3945) );
  AND U3930 ( .A(n4148), .B(n4149), .Z(n3946) );
  NANDN U3931 ( .A(n3950), .B(n4150), .Z(n4149) );
  NANDN U3932 ( .A(n3953), .B(n4151), .Z(n4148) );
  NAND U3933 ( .A(n3952), .B(n3950), .Z(n4151) );
  XOR U3934 ( .A(n4152), .B(n4153), .Z(n3950) );
  XNOR U3935 ( .A(n4154), .B(n4155), .Z(n4153) );
  IV U3936 ( .A(n4150), .Z(n3952) );
  NOR U3937 ( .A(n2947), .B(n2660), .Z(n4150) );
  AND U3938 ( .A(n4156), .B(n4157), .Z(n3953) );
  NANDN U3939 ( .A(n3958), .B(n3960), .Z(n4157) );
  NANDN U3940 ( .A(n3961), .B(n4158), .Z(n4156) );
  NANDN U3941 ( .A(n3960), .B(n3958), .Z(n4158) );
  XOR U3942 ( .A(n4159), .B(n4160), .Z(n3958) );
  XOR U3943 ( .A(n4161), .B(n4162), .Z(n4160) );
  AND U3944 ( .A(\stack[0][13] ), .B(\stack[1][2] ), .Z(n3960) );
  AND U3945 ( .A(n4163), .B(n4164), .Z(n3961) );
  NANDN U3946 ( .A(n3965), .B(n4165), .Z(n4164) );
  NANDN U3947 ( .A(n3968), .B(n4166), .Z(n4163) );
  NAND U3948 ( .A(n3967), .B(n3965), .Z(n4166) );
  XOR U3949 ( .A(n4167), .B(n4168), .Z(n3965) );
  XNOR U3950 ( .A(n4169), .B(n4170), .Z(n4168) );
  IV U3951 ( .A(n4165), .Z(n3967) );
  NOR U3952 ( .A(n2899), .B(n2660), .Z(n4165) );
  AND U3953 ( .A(n4171), .B(n4172), .Z(n3968) );
  NANDN U3954 ( .A(n3973), .B(n3975), .Z(n4172) );
  NANDN U3955 ( .A(n3976), .B(n4173), .Z(n4171) );
  NANDN U3956 ( .A(n3975), .B(n3973), .Z(n4173) );
  XOR U3957 ( .A(n4174), .B(n4175), .Z(n3973) );
  XOR U3958 ( .A(n4176), .B(n4177), .Z(n4175) );
  AND U3959 ( .A(\stack[0][11] ), .B(\stack[1][2] ), .Z(n3975) );
  AND U3960 ( .A(n4178), .B(n4179), .Z(n3976) );
  NANDN U3961 ( .A(n3980), .B(n4180), .Z(n4179) );
  NANDN U3962 ( .A(n3983), .B(n4181), .Z(n4178) );
  NAND U3963 ( .A(n3982), .B(n3980), .Z(n4181) );
  XOR U3964 ( .A(n4182), .B(n4183), .Z(n3980) );
  XNOR U3965 ( .A(n4184), .B(n4185), .Z(n4183) );
  IV U3966 ( .A(n4180), .Z(n3982) );
  NOR U3967 ( .A(n2851), .B(n2660), .Z(n4180) );
  AND U3968 ( .A(n4186), .B(n4187), .Z(n3983) );
  NANDN U3969 ( .A(n3988), .B(n3990), .Z(n4187) );
  NANDN U3970 ( .A(n3991), .B(n4188), .Z(n4186) );
  NANDN U3971 ( .A(n3990), .B(n3988), .Z(n4188) );
  XOR U3972 ( .A(n4189), .B(n4190), .Z(n3988) );
  XOR U3973 ( .A(n4191), .B(n4192), .Z(n4190) );
  AND U3974 ( .A(\stack[1][2] ), .B(\stack[0][9] ), .Z(n3990) );
  AND U3975 ( .A(n4193), .B(n4194), .Z(n3991) );
  NANDN U3976 ( .A(n3995), .B(n4195), .Z(n4194) );
  NANDN U3977 ( .A(n3998), .B(n4196), .Z(n4193) );
  NAND U3978 ( .A(n3997), .B(n3995), .Z(n4196) );
  XOR U3979 ( .A(n4197), .B(n4198), .Z(n3995) );
  XNOR U3980 ( .A(n4199), .B(n4200), .Z(n4198) );
  IV U3981 ( .A(n4195), .Z(n3997) );
  NOR U3982 ( .A(n2803), .B(n2660), .Z(n4195) );
  AND U3983 ( .A(n4201), .B(n4202), .Z(n3998) );
  NAND U3984 ( .A(n4005), .B(n4003), .Z(n4202) );
  NANDN U3985 ( .A(n4006), .B(n4203), .Z(n4201) );
  NOR U3986 ( .A(n2660), .B(n2779), .Z(n4005) );
  XNOR U3987 ( .A(n4204), .B(n4205), .Z(n4003) );
  XNOR U3988 ( .A(n4206), .B(n4207), .Z(n4205) );
  AND U3989 ( .A(n4208), .B(n4209), .Z(n4006) );
  NANDN U3990 ( .A(n4010), .B(n4210), .Z(n4209) );
  NANDN U3991 ( .A(n4013), .B(n4211), .Z(n4208) );
  NAND U3992 ( .A(n4012), .B(n4010), .Z(n4211) );
  XOR U3993 ( .A(n4212), .B(n4213), .Z(n4010) );
  XNOR U3994 ( .A(n4214), .B(n4215), .Z(n4213) );
  IV U3995 ( .A(n4210), .Z(n4012) );
  NOR U3996 ( .A(n2660), .B(n2755), .Z(n4210) );
  AND U3997 ( .A(n4216), .B(n4217), .Z(n4013) );
  NANDN U3998 ( .A(n4018), .B(n4020), .Z(n4217) );
  NANDN U3999 ( .A(n4021), .B(n4218), .Z(n4216) );
  NANDN U4000 ( .A(n4020), .B(n4018), .Z(n4218) );
  XOR U4001 ( .A(n4219), .B(n4220), .Z(n4018) );
  XOR U4002 ( .A(n4221), .B(n4222), .Z(n4220) );
  AND U4003 ( .A(\stack[1][2] ), .B(\stack[0][5] ), .Z(n4020) );
  AND U4004 ( .A(n4223), .B(n4224), .Z(n4021) );
  NANDN U4005 ( .A(n4025), .B(n4225), .Z(n4224) );
  NANDN U4006 ( .A(n4028), .B(n4226), .Z(n4223) );
  NAND U4007 ( .A(n4027), .B(n4025), .Z(n4226) );
  XOR U4008 ( .A(n4227), .B(n4228), .Z(n4025) );
  XNOR U4009 ( .A(n4229), .B(n4230), .Z(n4228) );
  IV U4010 ( .A(n4225), .Z(n4027) );
  NOR U4011 ( .A(n2660), .B(n2707), .Z(n4225) );
  AND U4012 ( .A(n4231), .B(n4232), .Z(n4028) );
  NANDN U4013 ( .A(n4033), .B(n4035), .Z(n4232) );
  NANDN U4014 ( .A(n4036), .B(n4233), .Z(n4231) );
  NANDN U4015 ( .A(n4035), .B(n4033), .Z(n4233) );
  XNOR U4016 ( .A(n4234), .B(n4235), .Z(n4033) );
  XNOR U4017 ( .A(n4236), .B(n4237), .Z(n4235) );
  AND U4018 ( .A(\stack[1][2] ), .B(\stack[0][3] ), .Z(n4035) );
  AND U4019 ( .A(n4238), .B(n4239), .Z(n4036) );
  NANDN U4020 ( .A(n4040), .B(n4042), .Z(n4239) );
  NAND U4021 ( .A(n4240), .B(n4043), .Z(n4238) );
  ANDN U4022 ( .B(n4241), .A(n4048), .Z(n4043) );
  NAND U4023 ( .A(\stack[1][2] ), .B(\stack[0][1] ), .Z(n4048) );
  AND U4024 ( .A(\stack[0][0] ), .B(\stack[1][3] ), .Z(n4241) );
  NANDN U4025 ( .A(n4042), .B(n4040), .Z(n4240) );
  XNOR U4026 ( .A(n4242), .B(n4243), .Z(n4040) );
  NAND U4027 ( .A(\stack[0][0] ), .B(\stack[1][4] ), .Z(n4243) );
  AND U4028 ( .A(\stack[1][2] ), .B(\stack[0][2] ), .Z(n4042) );
  NOR U4029 ( .A(n3283), .B(n2660), .Z(n3636) );
  IV U4030 ( .A(\stack[1][2] ), .Z(n2660) );
  IV U4031 ( .A(\stack[0][28] ), .Z(n3283) );
  XNOR U4032 ( .A(n3380), .B(n4244), .Z(n3635) );
  XNOR U4033 ( .A(n3379), .B(n3381), .Z(n4244) );
  AND U4034 ( .A(n4245), .B(n4246), .Z(n3381) );
  NANDN U4035 ( .A(n4054), .B(n4247), .Z(n4246) );
  NANDN U4036 ( .A(n4057), .B(n4248), .Z(n4245) );
  NAND U4037 ( .A(n4056), .B(n4054), .Z(n4248) );
  XOR U4038 ( .A(n4249), .B(n4250), .Z(n4054) );
  XNOR U4039 ( .A(n4251), .B(n4252), .Z(n4250) );
  IV U4040 ( .A(n4247), .Z(n4056) );
  NOR U4041 ( .A(n3235), .B(n2684), .Z(n4247) );
  AND U4042 ( .A(n4253), .B(n4254), .Z(n4057) );
  NANDN U4043 ( .A(n4062), .B(n4064), .Z(n4254) );
  NANDN U4044 ( .A(n4065), .B(n4255), .Z(n4253) );
  NANDN U4045 ( .A(n4064), .B(n4062), .Z(n4255) );
  XOR U4046 ( .A(n4256), .B(n4257), .Z(n4062) );
  XOR U4047 ( .A(n4258), .B(n4259), .Z(n4257) );
  AND U4048 ( .A(\stack[0][25] ), .B(\stack[1][3] ), .Z(n4064) );
  AND U4049 ( .A(n4260), .B(n4261), .Z(n4065) );
  NANDN U4050 ( .A(n4069), .B(n4262), .Z(n4261) );
  NANDN U4051 ( .A(n4072), .B(n4263), .Z(n4260) );
  NAND U4052 ( .A(n4071), .B(n4069), .Z(n4263) );
  XOR U4053 ( .A(n4264), .B(n4265), .Z(n4069) );
  XNOR U4054 ( .A(n4266), .B(n4267), .Z(n4265) );
  IV U4055 ( .A(n4262), .Z(n4071) );
  NOR U4056 ( .A(n3187), .B(n2684), .Z(n4262) );
  AND U4057 ( .A(n4268), .B(n4269), .Z(n4072) );
  NANDN U4058 ( .A(n4077), .B(n4079), .Z(n4269) );
  NANDN U4059 ( .A(n4080), .B(n4270), .Z(n4268) );
  NANDN U4060 ( .A(n4079), .B(n4077), .Z(n4270) );
  XOR U4061 ( .A(n4271), .B(n4272), .Z(n4077) );
  XOR U4062 ( .A(n4273), .B(n4274), .Z(n4272) );
  AND U4063 ( .A(\stack[0][23] ), .B(\stack[1][3] ), .Z(n4079) );
  AND U4064 ( .A(n4275), .B(n4276), .Z(n4080) );
  NANDN U4065 ( .A(n4084), .B(n4277), .Z(n4276) );
  NANDN U4066 ( .A(n4087), .B(n4278), .Z(n4275) );
  NAND U4067 ( .A(n4086), .B(n4084), .Z(n4278) );
  XOR U4068 ( .A(n4279), .B(n4280), .Z(n4084) );
  XNOR U4069 ( .A(n4281), .B(n4282), .Z(n4280) );
  IV U4070 ( .A(n4277), .Z(n4086) );
  NOR U4071 ( .A(n3139), .B(n2684), .Z(n4277) );
  AND U4072 ( .A(n4283), .B(n4284), .Z(n4087) );
  NANDN U4073 ( .A(n4092), .B(n4094), .Z(n4284) );
  NANDN U4074 ( .A(n4095), .B(n4285), .Z(n4283) );
  NANDN U4075 ( .A(n4094), .B(n4092), .Z(n4285) );
  XOR U4076 ( .A(n4286), .B(n4287), .Z(n4092) );
  XOR U4077 ( .A(n4288), .B(n4289), .Z(n4287) );
  AND U4078 ( .A(\stack[0][21] ), .B(\stack[1][3] ), .Z(n4094) );
  AND U4079 ( .A(n4290), .B(n4291), .Z(n4095) );
  NANDN U4080 ( .A(n4099), .B(n4292), .Z(n4291) );
  NANDN U4081 ( .A(n4102), .B(n4293), .Z(n4290) );
  NAND U4082 ( .A(n4101), .B(n4099), .Z(n4293) );
  XOR U4083 ( .A(n4294), .B(n4295), .Z(n4099) );
  XNOR U4084 ( .A(n4296), .B(n4297), .Z(n4295) );
  IV U4085 ( .A(n4292), .Z(n4101) );
  NOR U4086 ( .A(n3091), .B(n2684), .Z(n4292) );
  AND U4087 ( .A(n4298), .B(n4299), .Z(n4102) );
  NANDN U4088 ( .A(n4107), .B(n4109), .Z(n4299) );
  NANDN U4089 ( .A(n4110), .B(n4300), .Z(n4298) );
  NANDN U4090 ( .A(n4109), .B(n4107), .Z(n4300) );
  XOR U4091 ( .A(n4301), .B(n4302), .Z(n4107) );
  XOR U4092 ( .A(n4303), .B(n4304), .Z(n4302) );
  AND U4093 ( .A(\stack[0][19] ), .B(\stack[1][3] ), .Z(n4109) );
  AND U4094 ( .A(n4305), .B(n4306), .Z(n4110) );
  NANDN U4095 ( .A(n4114), .B(n4307), .Z(n4306) );
  NANDN U4096 ( .A(n4117), .B(n4308), .Z(n4305) );
  NAND U4097 ( .A(n4116), .B(n4114), .Z(n4308) );
  XOR U4098 ( .A(n4309), .B(n4310), .Z(n4114) );
  XNOR U4099 ( .A(n4311), .B(n4312), .Z(n4310) );
  IV U4100 ( .A(n4307), .Z(n4116) );
  NOR U4101 ( .A(n3043), .B(n2684), .Z(n4307) );
  AND U4102 ( .A(n4313), .B(n4314), .Z(n4117) );
  NANDN U4103 ( .A(n4122), .B(n4124), .Z(n4314) );
  NANDN U4104 ( .A(n4125), .B(n4315), .Z(n4313) );
  NANDN U4105 ( .A(n4124), .B(n4122), .Z(n4315) );
  XOR U4106 ( .A(n4316), .B(n4317), .Z(n4122) );
  XOR U4107 ( .A(n4318), .B(n4319), .Z(n4317) );
  AND U4108 ( .A(\stack[0][17] ), .B(\stack[1][3] ), .Z(n4124) );
  AND U4109 ( .A(n4320), .B(n4321), .Z(n4125) );
  NANDN U4110 ( .A(n4129), .B(n4322), .Z(n4321) );
  NANDN U4111 ( .A(n4132), .B(n4323), .Z(n4320) );
  NAND U4112 ( .A(n4131), .B(n4129), .Z(n4323) );
  XOR U4113 ( .A(n4324), .B(n4325), .Z(n4129) );
  XNOR U4114 ( .A(n4326), .B(n4327), .Z(n4325) );
  IV U4115 ( .A(n4322), .Z(n4131) );
  NOR U4116 ( .A(n2995), .B(n2684), .Z(n4322) );
  AND U4117 ( .A(n4328), .B(n4329), .Z(n4132) );
  NANDN U4118 ( .A(n4137), .B(n4139), .Z(n4329) );
  NANDN U4119 ( .A(n4140), .B(n4330), .Z(n4328) );
  NANDN U4120 ( .A(n4139), .B(n4137), .Z(n4330) );
  XOR U4121 ( .A(n4331), .B(n4332), .Z(n4137) );
  XOR U4122 ( .A(n4333), .B(n4334), .Z(n4332) );
  AND U4123 ( .A(\stack[0][15] ), .B(\stack[1][3] ), .Z(n4139) );
  AND U4124 ( .A(n4335), .B(n4336), .Z(n4140) );
  NANDN U4125 ( .A(n4144), .B(n4337), .Z(n4336) );
  NANDN U4126 ( .A(n4147), .B(n4338), .Z(n4335) );
  NAND U4127 ( .A(n4146), .B(n4144), .Z(n4338) );
  XOR U4128 ( .A(n4339), .B(n4340), .Z(n4144) );
  XNOR U4129 ( .A(n4341), .B(n4342), .Z(n4340) );
  IV U4130 ( .A(n4337), .Z(n4146) );
  NOR U4131 ( .A(n2947), .B(n2684), .Z(n4337) );
  AND U4132 ( .A(n4343), .B(n4344), .Z(n4147) );
  NANDN U4133 ( .A(n4152), .B(n4154), .Z(n4344) );
  NANDN U4134 ( .A(n4155), .B(n4345), .Z(n4343) );
  NANDN U4135 ( .A(n4154), .B(n4152), .Z(n4345) );
  XOR U4136 ( .A(n4346), .B(n4347), .Z(n4152) );
  XOR U4137 ( .A(n4348), .B(n4349), .Z(n4347) );
  AND U4138 ( .A(\stack[0][13] ), .B(\stack[1][3] ), .Z(n4154) );
  AND U4139 ( .A(n4350), .B(n4351), .Z(n4155) );
  NANDN U4140 ( .A(n4159), .B(n4352), .Z(n4351) );
  NANDN U4141 ( .A(n4162), .B(n4353), .Z(n4350) );
  NAND U4142 ( .A(n4161), .B(n4159), .Z(n4353) );
  XOR U4143 ( .A(n4354), .B(n4355), .Z(n4159) );
  XNOR U4144 ( .A(n4356), .B(n4357), .Z(n4355) );
  IV U4145 ( .A(n4352), .Z(n4161) );
  NOR U4146 ( .A(n2899), .B(n2684), .Z(n4352) );
  AND U4147 ( .A(n4358), .B(n4359), .Z(n4162) );
  NANDN U4148 ( .A(n4167), .B(n4169), .Z(n4359) );
  NANDN U4149 ( .A(n4170), .B(n4360), .Z(n4358) );
  NANDN U4150 ( .A(n4169), .B(n4167), .Z(n4360) );
  XOR U4151 ( .A(n4361), .B(n4362), .Z(n4167) );
  XOR U4152 ( .A(n4363), .B(n4364), .Z(n4362) );
  AND U4153 ( .A(\stack[0][11] ), .B(\stack[1][3] ), .Z(n4169) );
  AND U4154 ( .A(n4365), .B(n4366), .Z(n4170) );
  NANDN U4155 ( .A(n4174), .B(n4367), .Z(n4366) );
  NANDN U4156 ( .A(n4177), .B(n4368), .Z(n4365) );
  NAND U4157 ( .A(n4176), .B(n4174), .Z(n4368) );
  XOR U4158 ( .A(n4369), .B(n4370), .Z(n4174) );
  XNOR U4159 ( .A(n4371), .B(n4372), .Z(n4370) );
  IV U4160 ( .A(n4367), .Z(n4176) );
  NOR U4161 ( .A(n2851), .B(n2684), .Z(n4367) );
  AND U4162 ( .A(n4373), .B(n4374), .Z(n4177) );
  NANDN U4163 ( .A(n4182), .B(n4184), .Z(n4374) );
  NANDN U4164 ( .A(n4185), .B(n4375), .Z(n4373) );
  NANDN U4165 ( .A(n4184), .B(n4182), .Z(n4375) );
  XOR U4166 ( .A(n4376), .B(n4377), .Z(n4182) );
  XOR U4167 ( .A(n4378), .B(n4379), .Z(n4377) );
  AND U4168 ( .A(\stack[1][3] ), .B(\stack[0][9] ), .Z(n4184) );
  AND U4169 ( .A(n4380), .B(n4381), .Z(n4185) );
  NANDN U4170 ( .A(n4189), .B(n4382), .Z(n4381) );
  NANDN U4171 ( .A(n4192), .B(n4383), .Z(n4380) );
  NAND U4172 ( .A(n4191), .B(n4189), .Z(n4383) );
  XOR U4173 ( .A(n4384), .B(n4385), .Z(n4189) );
  XNOR U4174 ( .A(n4386), .B(n4387), .Z(n4385) );
  IV U4175 ( .A(n4382), .Z(n4191) );
  NOR U4176 ( .A(n2803), .B(n2684), .Z(n4382) );
  AND U4177 ( .A(n4388), .B(n4389), .Z(n4192) );
  NANDN U4178 ( .A(n4197), .B(n4199), .Z(n4389) );
  NANDN U4179 ( .A(n4200), .B(n4390), .Z(n4388) );
  NANDN U4180 ( .A(n4199), .B(n4197), .Z(n4390) );
  XOR U4181 ( .A(n4391), .B(n4392), .Z(n4197) );
  XOR U4182 ( .A(n4393), .B(n4394), .Z(n4392) );
  AND U4183 ( .A(\stack[0][7] ), .B(\stack[1][3] ), .Z(n4199) );
  AND U4184 ( .A(n4395), .B(n4396), .Z(n4200) );
  NANDN U4185 ( .A(n4204), .B(n4206), .Z(n4396) );
  NANDN U4186 ( .A(n4207), .B(n4397), .Z(n4395) );
  NANDN U4187 ( .A(n4206), .B(n4204), .Z(n4397) );
  XNOR U4188 ( .A(n4398), .B(n4399), .Z(n4204) );
  XNOR U4189 ( .A(n4400), .B(n4401), .Z(n4399) );
  ANDN U4190 ( .B(\stack[0][6] ), .A(n2684), .Z(n4206) );
  AND U4191 ( .A(n4402), .B(n4403), .Z(n4207) );
  NANDN U4192 ( .A(n4212), .B(n4214), .Z(n4403) );
  NANDN U4193 ( .A(n4215), .B(n4404), .Z(n4402) );
  NANDN U4194 ( .A(n4214), .B(n4212), .Z(n4404) );
  XOR U4195 ( .A(n4405), .B(n4406), .Z(n4212) );
  XOR U4196 ( .A(n4407), .B(n4408), .Z(n4406) );
  AND U4197 ( .A(\stack[1][3] ), .B(\stack[0][5] ), .Z(n4214) );
  AND U4198 ( .A(n4409), .B(n4410), .Z(n4215) );
  NANDN U4199 ( .A(n4219), .B(n4411), .Z(n4410) );
  NANDN U4200 ( .A(n4222), .B(n4412), .Z(n4409) );
  NAND U4201 ( .A(n4221), .B(n4219), .Z(n4412) );
  XOR U4202 ( .A(n4413), .B(n4414), .Z(n4219) );
  XNOR U4203 ( .A(n4415), .B(n4416), .Z(n4414) );
  IV U4204 ( .A(n4411), .Z(n4221) );
  NOR U4205 ( .A(n2684), .B(n2707), .Z(n4411) );
  AND U4206 ( .A(n4417), .B(n4418), .Z(n4222) );
  NANDN U4207 ( .A(n4227), .B(n4229), .Z(n4418) );
  NANDN U4208 ( .A(n4230), .B(n4419), .Z(n4417) );
  NANDN U4209 ( .A(n4229), .B(n4227), .Z(n4419) );
  XNOR U4210 ( .A(n4420), .B(n4421), .Z(n4227) );
  XNOR U4211 ( .A(n4422), .B(n4423), .Z(n4421) );
  AND U4212 ( .A(\stack[1][3] ), .B(\stack[0][3] ), .Z(n4229) );
  AND U4213 ( .A(n4424), .B(n4425), .Z(n4230) );
  NANDN U4214 ( .A(n4234), .B(n4236), .Z(n4425) );
  NAND U4215 ( .A(n4426), .B(n4237), .Z(n4424) );
  ANDN U4216 ( .B(n4427), .A(n4242), .Z(n4237) );
  NAND U4217 ( .A(\stack[1][3] ), .B(\stack[0][1] ), .Z(n4242) );
  AND U4218 ( .A(\stack[0][0] ), .B(\stack[1][4] ), .Z(n4427) );
  NANDN U4219 ( .A(n4236), .B(n4234), .Z(n4426) );
  XNOR U4220 ( .A(n4428), .B(n4429), .Z(n4234) );
  NAND U4221 ( .A(\stack[0][0] ), .B(\stack[1][5] ), .Z(n4429) );
  AND U4222 ( .A(\stack[1][3] ), .B(\stack[0][2] ), .Z(n4236) );
  NOR U4223 ( .A(n3259), .B(n2684), .Z(n3379) );
  IV U4224 ( .A(\stack[1][3] ), .Z(n2684) );
  IV U4225 ( .A(\stack[0][27] ), .Z(n3259) );
  XNOR U4226 ( .A(n3611), .B(n4430), .Z(n3380) );
  XNOR U4227 ( .A(n3612), .B(n3613), .Z(n4430) );
  AND U4228 ( .A(n4431), .B(n4432), .Z(n3613) );
  NANDN U4229 ( .A(n4249), .B(n4251), .Z(n4432) );
  NANDN U4230 ( .A(n4252), .B(n4433), .Z(n4431) );
  NANDN U4231 ( .A(n4251), .B(n4249), .Z(n4433) );
  XOR U4232 ( .A(n4434), .B(n4435), .Z(n4249) );
  XOR U4233 ( .A(n4436), .B(n4437), .Z(n4435) );
  AND U4234 ( .A(\stack[0][25] ), .B(\stack[1][4] ), .Z(n4251) );
  AND U4235 ( .A(n4438), .B(n4439), .Z(n4252) );
  NANDN U4236 ( .A(n4256), .B(n4440), .Z(n4439) );
  NANDN U4237 ( .A(n4259), .B(n4441), .Z(n4438) );
  NAND U4238 ( .A(n4258), .B(n4256), .Z(n4441) );
  XOR U4239 ( .A(n4442), .B(n4443), .Z(n4256) );
  XNOR U4240 ( .A(n4444), .B(n4445), .Z(n4443) );
  IV U4241 ( .A(n4440), .Z(n4258) );
  NOR U4242 ( .A(n3187), .B(n2708), .Z(n4440) );
  AND U4243 ( .A(n4446), .B(n4447), .Z(n4259) );
  NANDN U4244 ( .A(n4264), .B(n4266), .Z(n4447) );
  NANDN U4245 ( .A(n4267), .B(n4448), .Z(n4446) );
  NANDN U4246 ( .A(n4266), .B(n4264), .Z(n4448) );
  XOR U4247 ( .A(n4449), .B(n4450), .Z(n4264) );
  XOR U4248 ( .A(n4451), .B(n4452), .Z(n4450) );
  AND U4249 ( .A(\stack[0][23] ), .B(\stack[1][4] ), .Z(n4266) );
  AND U4250 ( .A(n4453), .B(n4454), .Z(n4267) );
  NANDN U4251 ( .A(n4271), .B(n4455), .Z(n4454) );
  NANDN U4252 ( .A(n4274), .B(n4456), .Z(n4453) );
  NAND U4253 ( .A(n4273), .B(n4271), .Z(n4456) );
  XOR U4254 ( .A(n4457), .B(n4458), .Z(n4271) );
  XNOR U4255 ( .A(n4459), .B(n4460), .Z(n4458) );
  IV U4256 ( .A(n4455), .Z(n4273) );
  NOR U4257 ( .A(n3139), .B(n2708), .Z(n4455) );
  AND U4258 ( .A(n4461), .B(n4462), .Z(n4274) );
  NANDN U4259 ( .A(n4279), .B(n4281), .Z(n4462) );
  NANDN U4260 ( .A(n4282), .B(n4463), .Z(n4461) );
  NANDN U4261 ( .A(n4281), .B(n4279), .Z(n4463) );
  XOR U4262 ( .A(n4464), .B(n4465), .Z(n4279) );
  XOR U4263 ( .A(n4466), .B(n4467), .Z(n4465) );
  AND U4264 ( .A(\stack[0][21] ), .B(\stack[1][4] ), .Z(n4281) );
  AND U4265 ( .A(n4468), .B(n4469), .Z(n4282) );
  NANDN U4266 ( .A(n4286), .B(n4470), .Z(n4469) );
  NANDN U4267 ( .A(n4289), .B(n4471), .Z(n4468) );
  NAND U4268 ( .A(n4288), .B(n4286), .Z(n4471) );
  XOR U4269 ( .A(n4472), .B(n4473), .Z(n4286) );
  XNOR U4270 ( .A(n4474), .B(n4475), .Z(n4473) );
  IV U4271 ( .A(n4470), .Z(n4288) );
  NOR U4272 ( .A(n3091), .B(n2708), .Z(n4470) );
  AND U4273 ( .A(n4476), .B(n4477), .Z(n4289) );
  NANDN U4274 ( .A(n4294), .B(n4296), .Z(n4477) );
  NANDN U4275 ( .A(n4297), .B(n4478), .Z(n4476) );
  NANDN U4276 ( .A(n4296), .B(n4294), .Z(n4478) );
  XOR U4277 ( .A(n4479), .B(n4480), .Z(n4294) );
  XOR U4278 ( .A(n4481), .B(n4482), .Z(n4480) );
  AND U4279 ( .A(\stack[0][19] ), .B(\stack[1][4] ), .Z(n4296) );
  AND U4280 ( .A(n4483), .B(n4484), .Z(n4297) );
  NANDN U4281 ( .A(n4301), .B(n4485), .Z(n4484) );
  NANDN U4282 ( .A(n4304), .B(n4486), .Z(n4483) );
  NAND U4283 ( .A(n4303), .B(n4301), .Z(n4486) );
  XOR U4284 ( .A(n4487), .B(n4488), .Z(n4301) );
  XNOR U4285 ( .A(n4489), .B(n4490), .Z(n4488) );
  IV U4286 ( .A(n4485), .Z(n4303) );
  NOR U4287 ( .A(n3043), .B(n2708), .Z(n4485) );
  AND U4288 ( .A(n4491), .B(n4492), .Z(n4304) );
  NANDN U4289 ( .A(n4309), .B(n4311), .Z(n4492) );
  NANDN U4290 ( .A(n4312), .B(n4493), .Z(n4491) );
  NANDN U4291 ( .A(n4311), .B(n4309), .Z(n4493) );
  XOR U4292 ( .A(n4494), .B(n4495), .Z(n4309) );
  XOR U4293 ( .A(n4496), .B(n4497), .Z(n4495) );
  AND U4294 ( .A(\stack[0][17] ), .B(\stack[1][4] ), .Z(n4311) );
  AND U4295 ( .A(n4498), .B(n4499), .Z(n4312) );
  NANDN U4296 ( .A(n4316), .B(n4500), .Z(n4499) );
  NANDN U4297 ( .A(n4319), .B(n4501), .Z(n4498) );
  NAND U4298 ( .A(n4318), .B(n4316), .Z(n4501) );
  XOR U4299 ( .A(n4502), .B(n4503), .Z(n4316) );
  XNOR U4300 ( .A(n4504), .B(n4505), .Z(n4503) );
  IV U4301 ( .A(n4500), .Z(n4318) );
  NOR U4302 ( .A(n2995), .B(n2708), .Z(n4500) );
  AND U4303 ( .A(n4506), .B(n4507), .Z(n4319) );
  NANDN U4304 ( .A(n4324), .B(n4326), .Z(n4507) );
  NANDN U4305 ( .A(n4327), .B(n4508), .Z(n4506) );
  NANDN U4306 ( .A(n4326), .B(n4324), .Z(n4508) );
  XOR U4307 ( .A(n4509), .B(n4510), .Z(n4324) );
  XOR U4308 ( .A(n4511), .B(n4512), .Z(n4510) );
  AND U4309 ( .A(\stack[0][15] ), .B(\stack[1][4] ), .Z(n4326) );
  AND U4310 ( .A(n4513), .B(n4514), .Z(n4327) );
  NANDN U4311 ( .A(n4331), .B(n4515), .Z(n4514) );
  NANDN U4312 ( .A(n4334), .B(n4516), .Z(n4513) );
  NAND U4313 ( .A(n4333), .B(n4331), .Z(n4516) );
  XOR U4314 ( .A(n4517), .B(n4518), .Z(n4331) );
  XNOR U4315 ( .A(n4519), .B(n4520), .Z(n4518) );
  IV U4316 ( .A(n4515), .Z(n4333) );
  NOR U4317 ( .A(n2947), .B(n2708), .Z(n4515) );
  AND U4318 ( .A(n4521), .B(n4522), .Z(n4334) );
  NANDN U4319 ( .A(n4339), .B(n4341), .Z(n4522) );
  NANDN U4320 ( .A(n4342), .B(n4523), .Z(n4521) );
  NANDN U4321 ( .A(n4341), .B(n4339), .Z(n4523) );
  XOR U4322 ( .A(n4524), .B(n4525), .Z(n4339) );
  XOR U4323 ( .A(n4526), .B(n4527), .Z(n4525) );
  AND U4324 ( .A(\stack[0][13] ), .B(\stack[1][4] ), .Z(n4341) );
  AND U4325 ( .A(n4528), .B(n4529), .Z(n4342) );
  NANDN U4326 ( .A(n4346), .B(n4530), .Z(n4529) );
  NANDN U4327 ( .A(n4349), .B(n4531), .Z(n4528) );
  NAND U4328 ( .A(n4348), .B(n4346), .Z(n4531) );
  XOR U4329 ( .A(n4532), .B(n4533), .Z(n4346) );
  XNOR U4330 ( .A(n4534), .B(n4535), .Z(n4533) );
  IV U4331 ( .A(n4530), .Z(n4348) );
  NOR U4332 ( .A(n2899), .B(n2708), .Z(n4530) );
  AND U4333 ( .A(n4536), .B(n4537), .Z(n4349) );
  NANDN U4334 ( .A(n4354), .B(n4356), .Z(n4537) );
  NANDN U4335 ( .A(n4357), .B(n4538), .Z(n4536) );
  NANDN U4336 ( .A(n4356), .B(n4354), .Z(n4538) );
  XOR U4337 ( .A(n4539), .B(n4540), .Z(n4354) );
  XOR U4338 ( .A(n4541), .B(n4542), .Z(n4540) );
  AND U4339 ( .A(\stack[0][11] ), .B(\stack[1][4] ), .Z(n4356) );
  AND U4340 ( .A(n4543), .B(n4544), .Z(n4357) );
  NANDN U4341 ( .A(n4361), .B(n4545), .Z(n4544) );
  NANDN U4342 ( .A(n4364), .B(n4546), .Z(n4543) );
  NAND U4343 ( .A(n4363), .B(n4361), .Z(n4546) );
  XOR U4344 ( .A(n4547), .B(n4548), .Z(n4361) );
  XNOR U4345 ( .A(n4549), .B(n4550), .Z(n4548) );
  IV U4346 ( .A(n4545), .Z(n4363) );
  NOR U4347 ( .A(n2851), .B(n2708), .Z(n4545) );
  AND U4348 ( .A(n4551), .B(n4552), .Z(n4364) );
  NANDN U4349 ( .A(n4369), .B(n4371), .Z(n4552) );
  NANDN U4350 ( .A(n4372), .B(n4553), .Z(n4551) );
  NANDN U4351 ( .A(n4371), .B(n4369), .Z(n4553) );
  XOR U4352 ( .A(n4554), .B(n4555), .Z(n4369) );
  XOR U4353 ( .A(n4556), .B(n4557), .Z(n4555) );
  AND U4354 ( .A(\stack[1][4] ), .B(\stack[0][9] ), .Z(n4371) );
  AND U4355 ( .A(n4558), .B(n4559), .Z(n4372) );
  NANDN U4356 ( .A(n4376), .B(n4560), .Z(n4559) );
  NANDN U4357 ( .A(n4379), .B(n4561), .Z(n4558) );
  NAND U4358 ( .A(n4378), .B(n4376), .Z(n4561) );
  XOR U4359 ( .A(n4562), .B(n4563), .Z(n4376) );
  XNOR U4360 ( .A(n4564), .B(n4565), .Z(n4563) );
  IV U4361 ( .A(n4560), .Z(n4378) );
  NOR U4362 ( .A(n2803), .B(n2708), .Z(n4560) );
  AND U4363 ( .A(n4566), .B(n4567), .Z(n4379) );
  NANDN U4364 ( .A(n4384), .B(n4386), .Z(n4567) );
  NANDN U4365 ( .A(n4387), .B(n4568), .Z(n4566) );
  NANDN U4366 ( .A(n4386), .B(n4384), .Z(n4568) );
  XOR U4367 ( .A(n4569), .B(n4570), .Z(n4384) );
  XOR U4368 ( .A(n4571), .B(n4572), .Z(n4570) );
  AND U4369 ( .A(\stack[0][7] ), .B(\stack[1][4] ), .Z(n4386) );
  AND U4370 ( .A(n4573), .B(n4574), .Z(n4387) );
  NANDN U4371 ( .A(n4391), .B(n4575), .Z(n4574) );
  NANDN U4372 ( .A(n4394), .B(n4576), .Z(n4573) );
  NAND U4373 ( .A(n4393), .B(n4391), .Z(n4576) );
  XOR U4374 ( .A(n4577), .B(n4578), .Z(n4391) );
  XNOR U4375 ( .A(n4579), .B(n4580), .Z(n4578) );
  IV U4376 ( .A(n4575), .Z(n4393) );
  NOR U4377 ( .A(n2755), .B(n2708), .Z(n4575) );
  AND U4378 ( .A(n4581), .B(n4582), .Z(n4394) );
  NAND U4379 ( .A(n4400), .B(n4398), .Z(n4582) );
  NANDN U4380 ( .A(n4401), .B(n4583), .Z(n4581) );
  NOR U4381 ( .A(n2708), .B(n2731), .Z(n4400) );
  XNOR U4382 ( .A(n4584), .B(n4585), .Z(n4398) );
  XNOR U4383 ( .A(n4586), .B(n4587), .Z(n4585) );
  AND U4384 ( .A(n4588), .B(n4589), .Z(n4401) );
  NANDN U4385 ( .A(n4405), .B(n4590), .Z(n4589) );
  NANDN U4386 ( .A(n4408), .B(n4591), .Z(n4588) );
  NAND U4387 ( .A(n4407), .B(n4405), .Z(n4591) );
  XOR U4388 ( .A(n4592), .B(n4593), .Z(n4405) );
  XNOR U4389 ( .A(n4594), .B(n4595), .Z(n4593) );
  IV U4390 ( .A(n4590), .Z(n4407) );
  NOR U4391 ( .A(n2708), .B(n2707), .Z(n4590) );
  IV U4392 ( .A(\stack[1][4] ), .Z(n2708) );
  AND U4393 ( .A(n4596), .B(n4597), .Z(n4408) );
  NANDN U4394 ( .A(n4413), .B(n4415), .Z(n4597) );
  NANDN U4395 ( .A(n4416), .B(n4598), .Z(n4596) );
  NANDN U4396 ( .A(n4415), .B(n4413), .Z(n4598) );
  XNOR U4397 ( .A(n4599), .B(n4600), .Z(n4413) );
  XNOR U4398 ( .A(n4601), .B(n4602), .Z(n4600) );
  AND U4399 ( .A(\stack[1][4] ), .B(\stack[0][3] ), .Z(n4415) );
  AND U4400 ( .A(n4603), .B(n4604), .Z(n4416) );
  NANDN U4401 ( .A(n4420), .B(n4422), .Z(n4604) );
  NAND U4402 ( .A(n4605), .B(n4423), .Z(n4603) );
  ANDN U4403 ( .B(n4606), .A(n4428), .Z(n4423) );
  NAND U4404 ( .A(\stack[1][4] ), .B(\stack[0][1] ), .Z(n4428) );
  AND U4405 ( .A(\stack[0][0] ), .B(\stack[1][5] ), .Z(n4606) );
  NANDN U4406 ( .A(n4422), .B(n4420), .Z(n4605) );
  XNOR U4407 ( .A(n4607), .B(n4608), .Z(n4420) );
  NAND U4408 ( .A(\stack[0][0] ), .B(\stack[1][6] ), .Z(n4608) );
  AND U4409 ( .A(\stack[1][4] ), .B(\stack[0][2] ), .Z(n4422) );
  ANDN U4410 ( .B(\stack[1][4] ), .A(n3235), .Z(n3612) );
  IV U4411 ( .A(\stack[0][26] ), .Z(n3235) );
  XNOR U4412 ( .A(n3622), .B(n4609), .Z(n3611) );
  XNOR U4413 ( .A(n3621), .B(n3623), .Z(n4609) );
  AND U4414 ( .A(n4610), .B(n4611), .Z(n3623) );
  NANDN U4415 ( .A(n4434), .B(n4612), .Z(n4611) );
  NANDN U4416 ( .A(n4437), .B(n4613), .Z(n4610) );
  NAND U4417 ( .A(n4436), .B(n4434), .Z(n4613) );
  XOR U4418 ( .A(n4614), .B(n4615), .Z(n4434) );
  XNOR U4419 ( .A(n4616), .B(n4617), .Z(n4615) );
  IV U4420 ( .A(n4612), .Z(n4436) );
  NOR U4421 ( .A(n3187), .B(n2732), .Z(n4612) );
  AND U4422 ( .A(n4618), .B(n4619), .Z(n4437) );
  NANDN U4423 ( .A(n4442), .B(n4444), .Z(n4619) );
  NANDN U4424 ( .A(n4445), .B(n4620), .Z(n4618) );
  NANDN U4425 ( .A(n4444), .B(n4442), .Z(n4620) );
  XOR U4426 ( .A(n4621), .B(n4622), .Z(n4442) );
  XOR U4427 ( .A(n4623), .B(n4624), .Z(n4622) );
  AND U4428 ( .A(\stack[0][23] ), .B(\stack[1][5] ), .Z(n4444) );
  AND U4429 ( .A(n4625), .B(n4626), .Z(n4445) );
  NANDN U4430 ( .A(n4449), .B(n4627), .Z(n4626) );
  NANDN U4431 ( .A(n4452), .B(n4628), .Z(n4625) );
  NAND U4432 ( .A(n4451), .B(n4449), .Z(n4628) );
  XOR U4433 ( .A(n4629), .B(n4630), .Z(n4449) );
  XNOR U4434 ( .A(n4631), .B(n4632), .Z(n4630) );
  IV U4435 ( .A(n4627), .Z(n4451) );
  NOR U4436 ( .A(n3139), .B(n2732), .Z(n4627) );
  AND U4437 ( .A(n4633), .B(n4634), .Z(n4452) );
  NANDN U4438 ( .A(n4457), .B(n4459), .Z(n4634) );
  NANDN U4439 ( .A(n4460), .B(n4635), .Z(n4633) );
  NANDN U4440 ( .A(n4459), .B(n4457), .Z(n4635) );
  XOR U4441 ( .A(n4636), .B(n4637), .Z(n4457) );
  XOR U4442 ( .A(n4638), .B(n4639), .Z(n4637) );
  AND U4443 ( .A(\stack[0][21] ), .B(\stack[1][5] ), .Z(n4459) );
  AND U4444 ( .A(n4640), .B(n4641), .Z(n4460) );
  NANDN U4445 ( .A(n4464), .B(n4642), .Z(n4641) );
  NANDN U4446 ( .A(n4467), .B(n4643), .Z(n4640) );
  NAND U4447 ( .A(n4466), .B(n4464), .Z(n4643) );
  XOR U4448 ( .A(n4644), .B(n4645), .Z(n4464) );
  XNOR U4449 ( .A(n4646), .B(n4647), .Z(n4645) );
  IV U4450 ( .A(n4642), .Z(n4466) );
  NOR U4451 ( .A(n3091), .B(n2732), .Z(n4642) );
  AND U4452 ( .A(n4648), .B(n4649), .Z(n4467) );
  NANDN U4453 ( .A(n4472), .B(n4474), .Z(n4649) );
  NANDN U4454 ( .A(n4475), .B(n4650), .Z(n4648) );
  NANDN U4455 ( .A(n4474), .B(n4472), .Z(n4650) );
  XOR U4456 ( .A(n4651), .B(n4652), .Z(n4472) );
  XOR U4457 ( .A(n4653), .B(n4654), .Z(n4652) );
  AND U4458 ( .A(\stack[0][19] ), .B(\stack[1][5] ), .Z(n4474) );
  AND U4459 ( .A(n4655), .B(n4656), .Z(n4475) );
  NANDN U4460 ( .A(n4479), .B(n4657), .Z(n4656) );
  NANDN U4461 ( .A(n4482), .B(n4658), .Z(n4655) );
  NAND U4462 ( .A(n4481), .B(n4479), .Z(n4658) );
  XOR U4463 ( .A(n4659), .B(n4660), .Z(n4479) );
  XNOR U4464 ( .A(n4661), .B(n4662), .Z(n4660) );
  IV U4465 ( .A(n4657), .Z(n4481) );
  NOR U4466 ( .A(n3043), .B(n2732), .Z(n4657) );
  AND U4467 ( .A(n4663), .B(n4664), .Z(n4482) );
  NANDN U4468 ( .A(n4487), .B(n4489), .Z(n4664) );
  NANDN U4469 ( .A(n4490), .B(n4665), .Z(n4663) );
  NANDN U4470 ( .A(n4489), .B(n4487), .Z(n4665) );
  XOR U4471 ( .A(n4666), .B(n4667), .Z(n4487) );
  XOR U4472 ( .A(n4668), .B(n4669), .Z(n4667) );
  AND U4473 ( .A(\stack[0][17] ), .B(\stack[1][5] ), .Z(n4489) );
  AND U4474 ( .A(n4670), .B(n4671), .Z(n4490) );
  NANDN U4475 ( .A(n4494), .B(n4672), .Z(n4671) );
  NANDN U4476 ( .A(n4497), .B(n4673), .Z(n4670) );
  NAND U4477 ( .A(n4496), .B(n4494), .Z(n4673) );
  XOR U4478 ( .A(n4674), .B(n4675), .Z(n4494) );
  XNOR U4479 ( .A(n4676), .B(n4677), .Z(n4675) );
  IV U4480 ( .A(n4672), .Z(n4496) );
  NOR U4481 ( .A(n2995), .B(n2732), .Z(n4672) );
  AND U4482 ( .A(n4678), .B(n4679), .Z(n4497) );
  NANDN U4483 ( .A(n4502), .B(n4504), .Z(n4679) );
  NANDN U4484 ( .A(n4505), .B(n4680), .Z(n4678) );
  NANDN U4485 ( .A(n4504), .B(n4502), .Z(n4680) );
  XOR U4486 ( .A(n4681), .B(n4682), .Z(n4502) );
  XOR U4487 ( .A(n4683), .B(n4684), .Z(n4682) );
  AND U4488 ( .A(\stack[0][15] ), .B(\stack[1][5] ), .Z(n4504) );
  AND U4489 ( .A(n4685), .B(n4686), .Z(n4505) );
  NANDN U4490 ( .A(n4509), .B(n4687), .Z(n4686) );
  NANDN U4491 ( .A(n4512), .B(n4688), .Z(n4685) );
  NAND U4492 ( .A(n4511), .B(n4509), .Z(n4688) );
  XOR U4493 ( .A(n4689), .B(n4690), .Z(n4509) );
  XNOR U4494 ( .A(n4691), .B(n4692), .Z(n4690) );
  IV U4495 ( .A(n4687), .Z(n4511) );
  NOR U4496 ( .A(n2947), .B(n2732), .Z(n4687) );
  AND U4497 ( .A(n4693), .B(n4694), .Z(n4512) );
  NANDN U4498 ( .A(n4517), .B(n4519), .Z(n4694) );
  NANDN U4499 ( .A(n4520), .B(n4695), .Z(n4693) );
  NANDN U4500 ( .A(n4519), .B(n4517), .Z(n4695) );
  XOR U4501 ( .A(n4696), .B(n4697), .Z(n4517) );
  XOR U4502 ( .A(n4698), .B(n4699), .Z(n4697) );
  AND U4503 ( .A(\stack[0][13] ), .B(\stack[1][5] ), .Z(n4519) );
  AND U4504 ( .A(n4700), .B(n4701), .Z(n4520) );
  NANDN U4505 ( .A(n4524), .B(n4702), .Z(n4701) );
  NANDN U4506 ( .A(n4527), .B(n4703), .Z(n4700) );
  NAND U4507 ( .A(n4526), .B(n4524), .Z(n4703) );
  XOR U4508 ( .A(n4704), .B(n4705), .Z(n4524) );
  XNOR U4509 ( .A(n4706), .B(n4707), .Z(n4705) );
  IV U4510 ( .A(n4702), .Z(n4526) );
  NOR U4511 ( .A(n2899), .B(n2732), .Z(n4702) );
  AND U4512 ( .A(n4708), .B(n4709), .Z(n4527) );
  NANDN U4513 ( .A(n4532), .B(n4534), .Z(n4709) );
  NANDN U4514 ( .A(n4535), .B(n4710), .Z(n4708) );
  NANDN U4515 ( .A(n4534), .B(n4532), .Z(n4710) );
  XOR U4516 ( .A(n4711), .B(n4712), .Z(n4532) );
  XOR U4517 ( .A(n4713), .B(n4714), .Z(n4712) );
  AND U4518 ( .A(\stack[0][11] ), .B(\stack[1][5] ), .Z(n4534) );
  AND U4519 ( .A(n4715), .B(n4716), .Z(n4535) );
  NANDN U4520 ( .A(n4539), .B(n4717), .Z(n4716) );
  NANDN U4521 ( .A(n4542), .B(n4718), .Z(n4715) );
  NAND U4522 ( .A(n4541), .B(n4539), .Z(n4718) );
  XOR U4523 ( .A(n4719), .B(n4720), .Z(n4539) );
  XNOR U4524 ( .A(n4721), .B(n4722), .Z(n4720) );
  IV U4525 ( .A(n4717), .Z(n4541) );
  NOR U4526 ( .A(n2851), .B(n2732), .Z(n4717) );
  AND U4527 ( .A(n4723), .B(n4724), .Z(n4542) );
  NANDN U4528 ( .A(n4547), .B(n4549), .Z(n4724) );
  NANDN U4529 ( .A(n4550), .B(n4725), .Z(n4723) );
  NANDN U4530 ( .A(n4549), .B(n4547), .Z(n4725) );
  XOR U4531 ( .A(n4726), .B(n4727), .Z(n4547) );
  XOR U4532 ( .A(n4728), .B(n4729), .Z(n4727) );
  AND U4533 ( .A(\stack[1][5] ), .B(\stack[0][9] ), .Z(n4549) );
  AND U4534 ( .A(n4730), .B(n4731), .Z(n4550) );
  NANDN U4535 ( .A(n4554), .B(n4732), .Z(n4731) );
  NANDN U4536 ( .A(n4557), .B(n4733), .Z(n4730) );
  NAND U4537 ( .A(n4556), .B(n4554), .Z(n4733) );
  XOR U4538 ( .A(n4734), .B(n4735), .Z(n4554) );
  XNOR U4539 ( .A(n4736), .B(n4737), .Z(n4735) );
  IV U4540 ( .A(n4732), .Z(n4556) );
  NOR U4541 ( .A(n2803), .B(n2732), .Z(n4732) );
  AND U4542 ( .A(n4738), .B(n4739), .Z(n4557) );
  NANDN U4543 ( .A(n4562), .B(n4564), .Z(n4739) );
  NANDN U4544 ( .A(n4565), .B(n4740), .Z(n4738) );
  NANDN U4545 ( .A(n4564), .B(n4562), .Z(n4740) );
  XOR U4546 ( .A(n4741), .B(n4742), .Z(n4562) );
  XOR U4547 ( .A(n4743), .B(n4744), .Z(n4742) );
  AND U4548 ( .A(\stack[0][7] ), .B(\stack[1][5] ), .Z(n4564) );
  AND U4549 ( .A(n4745), .B(n4746), .Z(n4565) );
  NANDN U4550 ( .A(n4569), .B(n4747), .Z(n4746) );
  NANDN U4551 ( .A(n4572), .B(n4748), .Z(n4745) );
  NAND U4552 ( .A(n4571), .B(n4569), .Z(n4748) );
  XOR U4553 ( .A(n4749), .B(n4750), .Z(n4569) );
  XNOR U4554 ( .A(n4751), .B(n4752), .Z(n4750) );
  IV U4555 ( .A(n4747), .Z(n4571) );
  NOR U4556 ( .A(n2755), .B(n2732), .Z(n4747) );
  AND U4557 ( .A(n4753), .B(n4754), .Z(n4572) );
  NANDN U4558 ( .A(n4577), .B(n4579), .Z(n4754) );
  NANDN U4559 ( .A(n4580), .B(n4755), .Z(n4753) );
  NANDN U4560 ( .A(n4579), .B(n4577), .Z(n4755) );
  XOR U4561 ( .A(n4756), .B(n4757), .Z(n4577) );
  XOR U4562 ( .A(n4758), .B(n4759), .Z(n4757) );
  AND U4563 ( .A(\stack[0][5] ), .B(\stack[1][5] ), .Z(n4579) );
  AND U4564 ( .A(n4760), .B(n4761), .Z(n4580) );
  NANDN U4565 ( .A(n4584), .B(n4586), .Z(n4761) );
  NANDN U4566 ( .A(n4587), .B(n4762), .Z(n4760) );
  NANDN U4567 ( .A(n4586), .B(n4584), .Z(n4762) );
  XNOR U4568 ( .A(n4763), .B(n4764), .Z(n4584) );
  XNOR U4569 ( .A(n4765), .B(n4766), .Z(n4764) );
  ANDN U4570 ( .B(\stack[0][4] ), .A(n2732), .Z(n4586) );
  AND U4571 ( .A(n4767), .B(n4768), .Z(n4587) );
  NANDN U4572 ( .A(n4592), .B(n4594), .Z(n4768) );
  NANDN U4573 ( .A(n4595), .B(n4769), .Z(n4767) );
  NANDN U4574 ( .A(n4594), .B(n4592), .Z(n4769) );
  XNOR U4575 ( .A(n4770), .B(n4771), .Z(n4592) );
  XNOR U4576 ( .A(n4772), .B(n4773), .Z(n4771) );
  AND U4577 ( .A(\stack[1][5] ), .B(\stack[0][3] ), .Z(n4594) );
  AND U4578 ( .A(n4774), .B(n4775), .Z(n4595) );
  NANDN U4579 ( .A(n4599), .B(n4601), .Z(n4775) );
  NAND U4580 ( .A(n4776), .B(n4602), .Z(n4774) );
  ANDN U4581 ( .B(n4777), .A(n4607), .Z(n4602) );
  NAND U4582 ( .A(\stack[1][5] ), .B(\stack[0][1] ), .Z(n4607) );
  AND U4583 ( .A(\stack[0][0] ), .B(\stack[1][6] ), .Z(n4777) );
  NANDN U4584 ( .A(n4601), .B(n4599), .Z(n4776) );
  XNOR U4585 ( .A(n4778), .B(n4779), .Z(n4599) );
  NAND U4586 ( .A(\stack[0][0] ), .B(\stack[1][7] ), .Z(n4779) );
  AND U4587 ( .A(\stack[1][5] ), .B(\stack[0][2] ), .Z(n4601) );
  NOR U4588 ( .A(n3211), .B(n2732), .Z(n3621) );
  IV U4589 ( .A(\stack[1][5] ), .Z(n2732) );
  IV U4590 ( .A(\stack[0][25] ), .Z(n3211) );
  XNOR U4591 ( .A(n3629), .B(n4780), .Z(n3622) );
  XNOR U4592 ( .A(n3630), .B(n3631), .Z(n4780) );
  AND U4593 ( .A(n4781), .B(n4782), .Z(n3631) );
  NANDN U4594 ( .A(n4614), .B(n4616), .Z(n4782) );
  NANDN U4595 ( .A(n4617), .B(n4783), .Z(n4781) );
  NANDN U4596 ( .A(n4616), .B(n4614), .Z(n4783) );
  XOR U4597 ( .A(n4784), .B(n4785), .Z(n4614) );
  XOR U4598 ( .A(n4786), .B(n4787), .Z(n4785) );
  AND U4599 ( .A(\stack[0][23] ), .B(\stack[1][6] ), .Z(n4616) );
  AND U4600 ( .A(n4788), .B(n4789), .Z(n4617) );
  NANDN U4601 ( .A(n4621), .B(n4790), .Z(n4789) );
  NANDN U4602 ( .A(n4624), .B(n4791), .Z(n4788) );
  NAND U4603 ( .A(n4623), .B(n4621), .Z(n4791) );
  XOR U4604 ( .A(n4792), .B(n4793), .Z(n4621) );
  XNOR U4605 ( .A(n4794), .B(n4795), .Z(n4793) );
  IV U4606 ( .A(n4790), .Z(n4623) );
  NOR U4607 ( .A(n3139), .B(n2756), .Z(n4790) );
  AND U4608 ( .A(n4796), .B(n4797), .Z(n4624) );
  NANDN U4609 ( .A(n4629), .B(n4631), .Z(n4797) );
  NANDN U4610 ( .A(n4632), .B(n4798), .Z(n4796) );
  NANDN U4611 ( .A(n4631), .B(n4629), .Z(n4798) );
  XOR U4612 ( .A(n4799), .B(n4800), .Z(n4629) );
  XOR U4613 ( .A(n4801), .B(n4802), .Z(n4800) );
  AND U4614 ( .A(\stack[0][21] ), .B(\stack[1][6] ), .Z(n4631) );
  AND U4615 ( .A(n4803), .B(n4804), .Z(n4632) );
  NANDN U4616 ( .A(n4636), .B(n4805), .Z(n4804) );
  NANDN U4617 ( .A(n4639), .B(n4806), .Z(n4803) );
  NAND U4618 ( .A(n4638), .B(n4636), .Z(n4806) );
  XOR U4619 ( .A(n4807), .B(n4808), .Z(n4636) );
  XNOR U4620 ( .A(n4809), .B(n4810), .Z(n4808) );
  IV U4621 ( .A(n4805), .Z(n4638) );
  NOR U4622 ( .A(n3091), .B(n2756), .Z(n4805) );
  AND U4623 ( .A(n4811), .B(n4812), .Z(n4639) );
  NANDN U4624 ( .A(n4644), .B(n4646), .Z(n4812) );
  NANDN U4625 ( .A(n4647), .B(n4813), .Z(n4811) );
  NANDN U4626 ( .A(n4646), .B(n4644), .Z(n4813) );
  XOR U4627 ( .A(n4814), .B(n4815), .Z(n4644) );
  XOR U4628 ( .A(n4816), .B(n4817), .Z(n4815) );
  AND U4629 ( .A(\stack[0][19] ), .B(\stack[1][6] ), .Z(n4646) );
  AND U4630 ( .A(n4818), .B(n4819), .Z(n4647) );
  NANDN U4631 ( .A(n4651), .B(n4820), .Z(n4819) );
  NANDN U4632 ( .A(n4654), .B(n4821), .Z(n4818) );
  NAND U4633 ( .A(n4653), .B(n4651), .Z(n4821) );
  XOR U4634 ( .A(n4822), .B(n4823), .Z(n4651) );
  XNOR U4635 ( .A(n4824), .B(n4825), .Z(n4823) );
  IV U4636 ( .A(n4820), .Z(n4653) );
  NOR U4637 ( .A(n3043), .B(n2756), .Z(n4820) );
  AND U4638 ( .A(n4826), .B(n4827), .Z(n4654) );
  NANDN U4639 ( .A(n4659), .B(n4661), .Z(n4827) );
  NANDN U4640 ( .A(n4662), .B(n4828), .Z(n4826) );
  NANDN U4641 ( .A(n4661), .B(n4659), .Z(n4828) );
  XOR U4642 ( .A(n4829), .B(n4830), .Z(n4659) );
  XOR U4643 ( .A(n4831), .B(n4832), .Z(n4830) );
  AND U4644 ( .A(\stack[0][17] ), .B(\stack[1][6] ), .Z(n4661) );
  AND U4645 ( .A(n4833), .B(n4834), .Z(n4662) );
  NANDN U4646 ( .A(n4666), .B(n4835), .Z(n4834) );
  NANDN U4647 ( .A(n4669), .B(n4836), .Z(n4833) );
  NAND U4648 ( .A(n4668), .B(n4666), .Z(n4836) );
  XOR U4649 ( .A(n4837), .B(n4838), .Z(n4666) );
  XNOR U4650 ( .A(n4839), .B(n4840), .Z(n4838) );
  IV U4651 ( .A(n4835), .Z(n4668) );
  NOR U4652 ( .A(n2995), .B(n2756), .Z(n4835) );
  AND U4653 ( .A(n4841), .B(n4842), .Z(n4669) );
  NANDN U4654 ( .A(n4674), .B(n4676), .Z(n4842) );
  NANDN U4655 ( .A(n4677), .B(n4843), .Z(n4841) );
  NANDN U4656 ( .A(n4676), .B(n4674), .Z(n4843) );
  XOR U4657 ( .A(n4844), .B(n4845), .Z(n4674) );
  XOR U4658 ( .A(n4846), .B(n4847), .Z(n4845) );
  AND U4659 ( .A(\stack[0][15] ), .B(\stack[1][6] ), .Z(n4676) );
  AND U4660 ( .A(n4848), .B(n4849), .Z(n4677) );
  NANDN U4661 ( .A(n4681), .B(n4850), .Z(n4849) );
  NANDN U4662 ( .A(n4684), .B(n4851), .Z(n4848) );
  NAND U4663 ( .A(n4683), .B(n4681), .Z(n4851) );
  XOR U4664 ( .A(n4852), .B(n4853), .Z(n4681) );
  XNOR U4665 ( .A(n4854), .B(n4855), .Z(n4853) );
  IV U4666 ( .A(n4850), .Z(n4683) );
  NOR U4667 ( .A(n2947), .B(n2756), .Z(n4850) );
  AND U4668 ( .A(n4856), .B(n4857), .Z(n4684) );
  NANDN U4669 ( .A(n4689), .B(n4691), .Z(n4857) );
  NANDN U4670 ( .A(n4692), .B(n4858), .Z(n4856) );
  NANDN U4671 ( .A(n4691), .B(n4689), .Z(n4858) );
  XOR U4672 ( .A(n4859), .B(n4860), .Z(n4689) );
  XOR U4673 ( .A(n4861), .B(n4862), .Z(n4860) );
  AND U4674 ( .A(\stack[0][13] ), .B(\stack[1][6] ), .Z(n4691) );
  AND U4675 ( .A(n4863), .B(n4864), .Z(n4692) );
  NANDN U4676 ( .A(n4696), .B(n4865), .Z(n4864) );
  NANDN U4677 ( .A(n4699), .B(n4866), .Z(n4863) );
  NAND U4678 ( .A(n4698), .B(n4696), .Z(n4866) );
  XOR U4679 ( .A(n4867), .B(n4868), .Z(n4696) );
  XNOR U4680 ( .A(n4869), .B(n4870), .Z(n4868) );
  IV U4681 ( .A(n4865), .Z(n4698) );
  NOR U4682 ( .A(n2899), .B(n2756), .Z(n4865) );
  AND U4683 ( .A(n4871), .B(n4872), .Z(n4699) );
  NANDN U4684 ( .A(n4704), .B(n4706), .Z(n4872) );
  NANDN U4685 ( .A(n4707), .B(n4873), .Z(n4871) );
  NANDN U4686 ( .A(n4706), .B(n4704), .Z(n4873) );
  XOR U4687 ( .A(n4874), .B(n4875), .Z(n4704) );
  XOR U4688 ( .A(n4876), .B(n4877), .Z(n4875) );
  AND U4689 ( .A(\stack[0][11] ), .B(\stack[1][6] ), .Z(n4706) );
  AND U4690 ( .A(n4878), .B(n4879), .Z(n4707) );
  NANDN U4691 ( .A(n4711), .B(n4880), .Z(n4879) );
  NANDN U4692 ( .A(n4714), .B(n4881), .Z(n4878) );
  NAND U4693 ( .A(n4713), .B(n4711), .Z(n4881) );
  XOR U4694 ( .A(n4882), .B(n4883), .Z(n4711) );
  XNOR U4695 ( .A(n4884), .B(n4885), .Z(n4883) );
  IV U4696 ( .A(n4880), .Z(n4713) );
  NOR U4697 ( .A(n2851), .B(n2756), .Z(n4880) );
  AND U4698 ( .A(n4886), .B(n4887), .Z(n4714) );
  NANDN U4699 ( .A(n4719), .B(n4721), .Z(n4887) );
  NANDN U4700 ( .A(n4722), .B(n4888), .Z(n4886) );
  NANDN U4701 ( .A(n4721), .B(n4719), .Z(n4888) );
  XOR U4702 ( .A(n4889), .B(n4890), .Z(n4719) );
  XOR U4703 ( .A(n4891), .B(n4892), .Z(n4890) );
  AND U4704 ( .A(\stack[1][6] ), .B(\stack[0][9] ), .Z(n4721) );
  AND U4705 ( .A(n4893), .B(n4894), .Z(n4722) );
  NANDN U4706 ( .A(n4726), .B(n4895), .Z(n4894) );
  NANDN U4707 ( .A(n4729), .B(n4896), .Z(n4893) );
  NAND U4708 ( .A(n4728), .B(n4726), .Z(n4896) );
  XOR U4709 ( .A(n4897), .B(n4898), .Z(n4726) );
  XNOR U4710 ( .A(n4899), .B(n4900), .Z(n4898) );
  IV U4711 ( .A(n4895), .Z(n4728) );
  NOR U4712 ( .A(n2803), .B(n2756), .Z(n4895) );
  AND U4713 ( .A(n4901), .B(n4902), .Z(n4729) );
  NANDN U4714 ( .A(n4734), .B(n4736), .Z(n4902) );
  NANDN U4715 ( .A(n4737), .B(n4903), .Z(n4901) );
  NANDN U4716 ( .A(n4736), .B(n4734), .Z(n4903) );
  XOR U4717 ( .A(n4904), .B(n4905), .Z(n4734) );
  XOR U4718 ( .A(n4906), .B(n4907), .Z(n4905) );
  AND U4719 ( .A(\stack[0][7] ), .B(\stack[1][6] ), .Z(n4736) );
  AND U4720 ( .A(n4908), .B(n4909), .Z(n4737) );
  NANDN U4721 ( .A(n4741), .B(n4910), .Z(n4909) );
  NANDN U4722 ( .A(n4744), .B(n4911), .Z(n4908) );
  NAND U4723 ( .A(n4743), .B(n4741), .Z(n4911) );
  XOR U4724 ( .A(n4912), .B(n4913), .Z(n4741) );
  XNOR U4725 ( .A(n4914), .B(n4915), .Z(n4913) );
  IV U4726 ( .A(n4910), .Z(n4743) );
  NOR U4727 ( .A(n2755), .B(n2756), .Z(n4910) );
  AND U4728 ( .A(n4916), .B(n4917), .Z(n4744) );
  NANDN U4729 ( .A(n4749), .B(n4751), .Z(n4917) );
  NANDN U4730 ( .A(n4752), .B(n4918), .Z(n4916) );
  NANDN U4731 ( .A(n4751), .B(n4749), .Z(n4918) );
  XOR U4732 ( .A(n4919), .B(n4920), .Z(n4749) );
  XOR U4733 ( .A(n4921), .B(n4922), .Z(n4920) );
  AND U4734 ( .A(\stack[0][5] ), .B(\stack[1][6] ), .Z(n4751) );
  AND U4735 ( .A(n4923), .B(n4924), .Z(n4752) );
  NANDN U4736 ( .A(n4756), .B(n4925), .Z(n4924) );
  NANDN U4737 ( .A(n4759), .B(n4926), .Z(n4923) );
  NAND U4738 ( .A(n4758), .B(n4756), .Z(n4926) );
  XOR U4739 ( .A(n4927), .B(n4928), .Z(n4756) );
  XNOR U4740 ( .A(n4929), .B(n4930), .Z(n4928) );
  IV U4741 ( .A(n4925), .Z(n4758) );
  NOR U4742 ( .A(n2707), .B(n2756), .Z(n4925) );
  AND U4743 ( .A(n4931), .B(n4932), .Z(n4759) );
  NAND U4744 ( .A(n4765), .B(n4763), .Z(n4932) );
  NANDN U4745 ( .A(n4766), .B(n4933), .Z(n4931) );
  NOR U4746 ( .A(n2756), .B(n2683), .Z(n4765) );
  IV U4747 ( .A(\stack[1][6] ), .Z(n2756) );
  XNOR U4748 ( .A(n4934), .B(n4935), .Z(n4763) );
  XOR U4749 ( .A(n4936), .B(n4937), .Z(n4935) );
  AND U4750 ( .A(n4938), .B(n4939), .Z(n4766) );
  NANDN U4751 ( .A(n4770), .B(n4772), .Z(n4939) );
  NAND U4752 ( .A(n4940), .B(n4773), .Z(n4938) );
  ANDN U4753 ( .B(n4941), .A(n4778), .Z(n4773) );
  NAND U4754 ( .A(\stack[1][6] ), .B(\stack[0][1] ), .Z(n4778) );
  AND U4755 ( .A(\stack[0][0] ), .B(\stack[1][7] ), .Z(n4941) );
  NANDN U4756 ( .A(n4772), .B(n4770), .Z(n4940) );
  XNOR U4757 ( .A(n4942), .B(n4943), .Z(n4770) );
  NAND U4758 ( .A(\stack[1][8] ), .B(\stack[0][0] ), .Z(n4943) );
  AND U4759 ( .A(\stack[1][6] ), .B(\stack[0][2] ), .Z(n4772) );
  ANDN U4760 ( .B(\stack[1][6] ), .A(n3187), .Z(n3630) );
  IV U4761 ( .A(\stack[0][24] ), .Z(n3187) );
  XNOR U4762 ( .A(n3394), .B(n4944), .Z(n3629) );
  XNOR U4763 ( .A(n3393), .B(n3395), .Z(n4944) );
  AND U4764 ( .A(n4945), .B(n4946), .Z(n3395) );
  NANDN U4765 ( .A(n4784), .B(n4947), .Z(n4946) );
  NANDN U4766 ( .A(n4787), .B(n4948), .Z(n4945) );
  NAND U4767 ( .A(n4786), .B(n4784), .Z(n4948) );
  XOR U4768 ( .A(n4949), .B(n4950), .Z(n4784) );
  XNOR U4769 ( .A(n4951), .B(n4952), .Z(n4950) );
  IV U4770 ( .A(n4947), .Z(n4786) );
  NOR U4771 ( .A(n3139), .B(n2780), .Z(n4947) );
  AND U4772 ( .A(n4953), .B(n4954), .Z(n4787) );
  NANDN U4773 ( .A(n4792), .B(n4794), .Z(n4954) );
  NANDN U4774 ( .A(n4795), .B(n4955), .Z(n4953) );
  NANDN U4775 ( .A(n4794), .B(n4792), .Z(n4955) );
  XOR U4776 ( .A(n4956), .B(n4957), .Z(n4792) );
  XOR U4777 ( .A(n4958), .B(n4959), .Z(n4957) );
  AND U4778 ( .A(\stack[0][21] ), .B(\stack[1][7] ), .Z(n4794) );
  AND U4779 ( .A(n4960), .B(n4961), .Z(n4795) );
  NANDN U4780 ( .A(n4799), .B(n4962), .Z(n4961) );
  NANDN U4781 ( .A(n4802), .B(n4963), .Z(n4960) );
  NAND U4782 ( .A(n4801), .B(n4799), .Z(n4963) );
  XOR U4783 ( .A(n4964), .B(n4965), .Z(n4799) );
  XNOR U4784 ( .A(n4966), .B(n4967), .Z(n4965) );
  IV U4785 ( .A(n4962), .Z(n4801) );
  NOR U4786 ( .A(n3091), .B(n2780), .Z(n4962) );
  AND U4787 ( .A(n4968), .B(n4969), .Z(n4802) );
  NANDN U4788 ( .A(n4807), .B(n4809), .Z(n4969) );
  NANDN U4789 ( .A(n4810), .B(n4970), .Z(n4968) );
  NANDN U4790 ( .A(n4809), .B(n4807), .Z(n4970) );
  XOR U4791 ( .A(n4971), .B(n4972), .Z(n4807) );
  XOR U4792 ( .A(n4973), .B(n4974), .Z(n4972) );
  AND U4793 ( .A(\stack[0][19] ), .B(\stack[1][7] ), .Z(n4809) );
  AND U4794 ( .A(n4975), .B(n4976), .Z(n4810) );
  NANDN U4795 ( .A(n4814), .B(n4977), .Z(n4976) );
  NANDN U4796 ( .A(n4817), .B(n4978), .Z(n4975) );
  NAND U4797 ( .A(n4816), .B(n4814), .Z(n4978) );
  XOR U4798 ( .A(n4979), .B(n4980), .Z(n4814) );
  XNOR U4799 ( .A(n4981), .B(n4982), .Z(n4980) );
  IV U4800 ( .A(n4977), .Z(n4816) );
  NOR U4801 ( .A(n3043), .B(n2780), .Z(n4977) );
  AND U4802 ( .A(n4983), .B(n4984), .Z(n4817) );
  NANDN U4803 ( .A(n4822), .B(n4824), .Z(n4984) );
  NANDN U4804 ( .A(n4825), .B(n4985), .Z(n4983) );
  NANDN U4805 ( .A(n4824), .B(n4822), .Z(n4985) );
  XOR U4806 ( .A(n4986), .B(n4987), .Z(n4822) );
  XOR U4807 ( .A(n4988), .B(n4989), .Z(n4987) );
  AND U4808 ( .A(\stack[0][17] ), .B(\stack[1][7] ), .Z(n4824) );
  AND U4809 ( .A(n4990), .B(n4991), .Z(n4825) );
  NANDN U4810 ( .A(n4829), .B(n4992), .Z(n4991) );
  NANDN U4811 ( .A(n4832), .B(n4993), .Z(n4990) );
  NAND U4812 ( .A(n4831), .B(n4829), .Z(n4993) );
  XOR U4813 ( .A(n4994), .B(n4995), .Z(n4829) );
  XNOR U4814 ( .A(n4996), .B(n4997), .Z(n4995) );
  IV U4815 ( .A(n4992), .Z(n4831) );
  NOR U4816 ( .A(n2995), .B(n2780), .Z(n4992) );
  AND U4817 ( .A(n4998), .B(n4999), .Z(n4832) );
  NANDN U4818 ( .A(n4837), .B(n4839), .Z(n4999) );
  NANDN U4819 ( .A(n4840), .B(n5000), .Z(n4998) );
  NANDN U4820 ( .A(n4839), .B(n4837), .Z(n5000) );
  XOR U4821 ( .A(n5001), .B(n5002), .Z(n4837) );
  XOR U4822 ( .A(n5003), .B(n5004), .Z(n5002) );
  AND U4823 ( .A(\stack[0][15] ), .B(\stack[1][7] ), .Z(n4839) );
  AND U4824 ( .A(n5005), .B(n5006), .Z(n4840) );
  NANDN U4825 ( .A(n4844), .B(n5007), .Z(n5006) );
  NANDN U4826 ( .A(n4847), .B(n5008), .Z(n5005) );
  NAND U4827 ( .A(n4846), .B(n4844), .Z(n5008) );
  XOR U4828 ( .A(n5009), .B(n5010), .Z(n4844) );
  XNOR U4829 ( .A(n5011), .B(n5012), .Z(n5010) );
  IV U4830 ( .A(n5007), .Z(n4846) );
  NOR U4831 ( .A(n2947), .B(n2780), .Z(n5007) );
  AND U4832 ( .A(n5013), .B(n5014), .Z(n4847) );
  NANDN U4833 ( .A(n4852), .B(n4854), .Z(n5014) );
  NANDN U4834 ( .A(n4855), .B(n5015), .Z(n5013) );
  NANDN U4835 ( .A(n4854), .B(n4852), .Z(n5015) );
  XOR U4836 ( .A(n5016), .B(n5017), .Z(n4852) );
  XOR U4837 ( .A(n5018), .B(n5019), .Z(n5017) );
  AND U4838 ( .A(\stack[0][13] ), .B(\stack[1][7] ), .Z(n4854) );
  AND U4839 ( .A(n5020), .B(n5021), .Z(n4855) );
  NANDN U4840 ( .A(n4859), .B(n5022), .Z(n5021) );
  NANDN U4841 ( .A(n4862), .B(n5023), .Z(n5020) );
  NAND U4842 ( .A(n4861), .B(n4859), .Z(n5023) );
  XOR U4843 ( .A(n5024), .B(n5025), .Z(n4859) );
  XNOR U4844 ( .A(n5026), .B(n5027), .Z(n5025) );
  IV U4845 ( .A(n5022), .Z(n4861) );
  NOR U4846 ( .A(n2899), .B(n2780), .Z(n5022) );
  AND U4847 ( .A(n5028), .B(n5029), .Z(n4862) );
  NANDN U4848 ( .A(n4867), .B(n4869), .Z(n5029) );
  NANDN U4849 ( .A(n4870), .B(n5030), .Z(n5028) );
  NANDN U4850 ( .A(n4869), .B(n4867), .Z(n5030) );
  XOR U4851 ( .A(n5031), .B(n5032), .Z(n4867) );
  XOR U4852 ( .A(n5033), .B(n5034), .Z(n5032) );
  AND U4853 ( .A(\stack[0][11] ), .B(\stack[1][7] ), .Z(n4869) );
  AND U4854 ( .A(n5035), .B(n5036), .Z(n4870) );
  NANDN U4855 ( .A(n4874), .B(n5037), .Z(n5036) );
  NANDN U4856 ( .A(n4877), .B(n5038), .Z(n5035) );
  NAND U4857 ( .A(n4876), .B(n4874), .Z(n5038) );
  XOR U4858 ( .A(n5039), .B(n5040), .Z(n4874) );
  XNOR U4859 ( .A(n5041), .B(n5042), .Z(n5040) );
  IV U4860 ( .A(n5037), .Z(n4876) );
  NOR U4861 ( .A(n2851), .B(n2780), .Z(n5037) );
  AND U4862 ( .A(n5043), .B(n5044), .Z(n4877) );
  NANDN U4863 ( .A(n4882), .B(n4884), .Z(n5044) );
  NANDN U4864 ( .A(n4885), .B(n5045), .Z(n5043) );
  NANDN U4865 ( .A(n4884), .B(n4882), .Z(n5045) );
  XOR U4866 ( .A(n5046), .B(n5047), .Z(n4882) );
  XOR U4867 ( .A(n5048), .B(n5049), .Z(n5047) );
  AND U4868 ( .A(\stack[1][7] ), .B(\stack[0][9] ), .Z(n4884) );
  AND U4869 ( .A(n5050), .B(n5051), .Z(n4885) );
  NANDN U4870 ( .A(n4889), .B(n5052), .Z(n5051) );
  NANDN U4871 ( .A(n4892), .B(n5053), .Z(n5050) );
  NAND U4872 ( .A(n4891), .B(n4889), .Z(n5053) );
  XOR U4873 ( .A(n5054), .B(n5055), .Z(n4889) );
  XNOR U4874 ( .A(n5056), .B(n5057), .Z(n5055) );
  IV U4875 ( .A(n5052), .Z(n4891) );
  NOR U4876 ( .A(n2803), .B(n2780), .Z(n5052) );
  AND U4877 ( .A(n5058), .B(n5059), .Z(n4892) );
  NANDN U4878 ( .A(n4897), .B(n4899), .Z(n5059) );
  NANDN U4879 ( .A(n4900), .B(n5060), .Z(n5058) );
  NANDN U4880 ( .A(n4899), .B(n4897), .Z(n5060) );
  XOR U4881 ( .A(n5061), .B(n5062), .Z(n4897) );
  XOR U4882 ( .A(n5063), .B(n5064), .Z(n5062) );
  AND U4883 ( .A(\stack[0][7] ), .B(\stack[1][7] ), .Z(n4899) );
  AND U4884 ( .A(n5065), .B(n5066), .Z(n4900) );
  NANDN U4885 ( .A(n4904), .B(n5067), .Z(n5066) );
  NANDN U4886 ( .A(n4907), .B(n5068), .Z(n5065) );
  NAND U4887 ( .A(n4906), .B(n4904), .Z(n5068) );
  XOR U4888 ( .A(n5069), .B(n5070), .Z(n4904) );
  XNOR U4889 ( .A(n5071), .B(n5072), .Z(n5070) );
  IV U4890 ( .A(n5067), .Z(n4906) );
  NOR U4891 ( .A(n2755), .B(n2780), .Z(n5067) );
  AND U4892 ( .A(n5073), .B(n5074), .Z(n4907) );
  NANDN U4893 ( .A(n4912), .B(n4914), .Z(n5074) );
  NANDN U4894 ( .A(n4915), .B(n5075), .Z(n5073) );
  NANDN U4895 ( .A(n4914), .B(n4912), .Z(n5075) );
  XOR U4896 ( .A(n5076), .B(n5077), .Z(n4912) );
  XOR U4897 ( .A(n5078), .B(n5079), .Z(n5077) );
  AND U4898 ( .A(\stack[0][5] ), .B(\stack[1][7] ), .Z(n4914) );
  AND U4899 ( .A(n5080), .B(n5081), .Z(n4915) );
  NANDN U4900 ( .A(n4919), .B(n5082), .Z(n5081) );
  NANDN U4901 ( .A(n4922), .B(n5083), .Z(n5080) );
  NAND U4902 ( .A(n4921), .B(n4919), .Z(n5083) );
  XOR U4903 ( .A(n5084), .B(n5085), .Z(n4919) );
  XNOR U4904 ( .A(n5086), .B(n5087), .Z(n5085) );
  IV U4905 ( .A(n5082), .Z(n4921) );
  NOR U4906 ( .A(n2707), .B(n2780), .Z(n5082) );
  AND U4907 ( .A(n5088), .B(n5089), .Z(n4922) );
  NANDN U4908 ( .A(n4927), .B(n4929), .Z(n5089) );
  NANDN U4909 ( .A(n4930), .B(n5090), .Z(n5088) );
  NANDN U4910 ( .A(n4929), .B(n4927), .Z(n5090) );
  XNOR U4911 ( .A(n5091), .B(n5092), .Z(n4927) );
  XOR U4912 ( .A(n5093), .B(n5094), .Z(n5092) );
  AND U4913 ( .A(\stack[0][3] ), .B(\stack[1][7] ), .Z(n4929) );
  AND U4914 ( .A(n5095), .B(n5096), .Z(n4930) );
  NAND U4915 ( .A(n4934), .B(n4937), .Z(n5096) );
  NANDN U4916 ( .A(n4936), .B(n5097), .Z(n5095) );
  OR U4917 ( .A(n4934), .B(n4937), .Z(n5097) );
  AND U4918 ( .A(\stack[0][2] ), .B(\stack[1][7] ), .Z(n4937) );
  XOR U4919 ( .A(n5098), .B(n5099), .Z(n4934) );
  NAND U4920 ( .A(\stack[1][9] ), .B(\stack[0][0] ), .Z(n5099) );
  NANDN U4921 ( .A(n4942), .B(n5100), .Z(n4936) );
  AND U4922 ( .A(\stack[1][8] ), .B(\stack[0][0] ), .Z(n5100) );
  NAND U4923 ( .A(\stack[1][7] ), .B(\stack[0][1] ), .Z(n4942) );
  NOR U4924 ( .A(n3163), .B(n2780), .Z(n3393) );
  IV U4925 ( .A(\stack[1][7] ), .Z(n2780) );
  IV U4926 ( .A(\stack[0][23] ), .Z(n3163) );
  XNOR U4927 ( .A(n3585), .B(n5101), .Z(n3394) );
  XNOR U4928 ( .A(n3586), .B(n3587), .Z(n5101) );
  AND U4929 ( .A(n5102), .B(n5103), .Z(n3587) );
  NANDN U4930 ( .A(n4949), .B(n4951), .Z(n5103) );
  NANDN U4931 ( .A(n4952), .B(n5104), .Z(n5102) );
  NANDN U4932 ( .A(n4951), .B(n4949), .Z(n5104) );
  XOR U4933 ( .A(n5105), .B(n5106), .Z(n4949) );
  XOR U4934 ( .A(n5107), .B(n5108), .Z(n5106) );
  AND U4935 ( .A(\stack[0][21] ), .B(\stack[1][8] ), .Z(n4951) );
  AND U4936 ( .A(n5109), .B(n5110), .Z(n4952) );
  NANDN U4937 ( .A(n4956), .B(n5111), .Z(n5110) );
  NANDN U4938 ( .A(n4959), .B(n5112), .Z(n5109) );
  NAND U4939 ( .A(n4958), .B(n4956), .Z(n5112) );
  XOR U4940 ( .A(n5113), .B(n5114), .Z(n4956) );
  XNOR U4941 ( .A(n5115), .B(n5116), .Z(n5114) );
  IV U4942 ( .A(n5111), .Z(n4958) );
  NOR U4943 ( .A(n3091), .B(n2804), .Z(n5111) );
  AND U4944 ( .A(n5117), .B(n5118), .Z(n4959) );
  NANDN U4945 ( .A(n4964), .B(n4966), .Z(n5118) );
  NANDN U4946 ( .A(n4967), .B(n5119), .Z(n5117) );
  NANDN U4947 ( .A(n4966), .B(n4964), .Z(n5119) );
  XOR U4948 ( .A(n5120), .B(n5121), .Z(n4964) );
  XOR U4949 ( .A(n5122), .B(n5123), .Z(n5121) );
  AND U4950 ( .A(\stack[0][19] ), .B(\stack[1][8] ), .Z(n4966) );
  AND U4951 ( .A(n5124), .B(n5125), .Z(n4967) );
  NANDN U4952 ( .A(n4971), .B(n5126), .Z(n5125) );
  NANDN U4953 ( .A(n4974), .B(n5127), .Z(n5124) );
  NAND U4954 ( .A(n4973), .B(n4971), .Z(n5127) );
  XOR U4955 ( .A(n5128), .B(n5129), .Z(n4971) );
  XNOR U4956 ( .A(n5130), .B(n5131), .Z(n5129) );
  IV U4957 ( .A(n5126), .Z(n4973) );
  NOR U4958 ( .A(n3043), .B(n2804), .Z(n5126) );
  AND U4959 ( .A(n5132), .B(n5133), .Z(n4974) );
  NANDN U4960 ( .A(n4979), .B(n4981), .Z(n5133) );
  NANDN U4961 ( .A(n4982), .B(n5134), .Z(n5132) );
  NANDN U4962 ( .A(n4981), .B(n4979), .Z(n5134) );
  XOR U4963 ( .A(n5135), .B(n5136), .Z(n4979) );
  XOR U4964 ( .A(n5137), .B(n5138), .Z(n5136) );
  AND U4965 ( .A(\stack[0][17] ), .B(\stack[1][8] ), .Z(n4981) );
  AND U4966 ( .A(n5139), .B(n5140), .Z(n4982) );
  NANDN U4967 ( .A(n4986), .B(n5141), .Z(n5140) );
  NANDN U4968 ( .A(n4989), .B(n5142), .Z(n5139) );
  NAND U4969 ( .A(n4988), .B(n4986), .Z(n5142) );
  XOR U4970 ( .A(n5143), .B(n5144), .Z(n4986) );
  XNOR U4971 ( .A(n5145), .B(n5146), .Z(n5144) );
  IV U4972 ( .A(n5141), .Z(n4988) );
  NOR U4973 ( .A(n2995), .B(n2804), .Z(n5141) );
  AND U4974 ( .A(n5147), .B(n5148), .Z(n4989) );
  NANDN U4975 ( .A(n4994), .B(n4996), .Z(n5148) );
  NANDN U4976 ( .A(n4997), .B(n5149), .Z(n5147) );
  NANDN U4977 ( .A(n4996), .B(n4994), .Z(n5149) );
  XOR U4978 ( .A(n5150), .B(n5151), .Z(n4994) );
  XOR U4979 ( .A(n5152), .B(n5153), .Z(n5151) );
  AND U4980 ( .A(\stack[0][15] ), .B(\stack[1][8] ), .Z(n4996) );
  AND U4981 ( .A(n5154), .B(n5155), .Z(n4997) );
  NANDN U4982 ( .A(n5001), .B(n5156), .Z(n5155) );
  NANDN U4983 ( .A(n5004), .B(n5157), .Z(n5154) );
  NAND U4984 ( .A(n5003), .B(n5001), .Z(n5157) );
  XOR U4985 ( .A(n5158), .B(n5159), .Z(n5001) );
  XNOR U4986 ( .A(n5160), .B(n5161), .Z(n5159) );
  IV U4987 ( .A(n5156), .Z(n5003) );
  NOR U4988 ( .A(n2947), .B(n2804), .Z(n5156) );
  AND U4989 ( .A(n5162), .B(n5163), .Z(n5004) );
  NANDN U4990 ( .A(n5009), .B(n5011), .Z(n5163) );
  NANDN U4991 ( .A(n5012), .B(n5164), .Z(n5162) );
  NANDN U4992 ( .A(n5011), .B(n5009), .Z(n5164) );
  XOR U4993 ( .A(n5165), .B(n5166), .Z(n5009) );
  XOR U4994 ( .A(n5167), .B(n5168), .Z(n5166) );
  AND U4995 ( .A(\stack[0][13] ), .B(\stack[1][8] ), .Z(n5011) );
  AND U4996 ( .A(n5169), .B(n5170), .Z(n5012) );
  NANDN U4997 ( .A(n5016), .B(n5171), .Z(n5170) );
  NANDN U4998 ( .A(n5019), .B(n5172), .Z(n5169) );
  NAND U4999 ( .A(n5018), .B(n5016), .Z(n5172) );
  XOR U5000 ( .A(n5173), .B(n5174), .Z(n5016) );
  XNOR U5001 ( .A(n5175), .B(n5176), .Z(n5174) );
  IV U5002 ( .A(n5171), .Z(n5018) );
  NOR U5003 ( .A(n2899), .B(n2804), .Z(n5171) );
  AND U5004 ( .A(n5177), .B(n5178), .Z(n5019) );
  NANDN U5005 ( .A(n5024), .B(n5026), .Z(n5178) );
  NANDN U5006 ( .A(n5027), .B(n5179), .Z(n5177) );
  NANDN U5007 ( .A(n5026), .B(n5024), .Z(n5179) );
  XOR U5008 ( .A(n5180), .B(n5181), .Z(n5024) );
  XOR U5009 ( .A(n5182), .B(n5183), .Z(n5181) );
  AND U5010 ( .A(\stack[0][11] ), .B(\stack[1][8] ), .Z(n5026) );
  AND U5011 ( .A(n5184), .B(n5185), .Z(n5027) );
  NANDN U5012 ( .A(n5031), .B(n5186), .Z(n5185) );
  NANDN U5013 ( .A(n5034), .B(n5187), .Z(n5184) );
  NAND U5014 ( .A(n5033), .B(n5031), .Z(n5187) );
  XOR U5015 ( .A(n5188), .B(n5189), .Z(n5031) );
  XNOR U5016 ( .A(n5190), .B(n5191), .Z(n5189) );
  IV U5017 ( .A(n5186), .Z(n5033) );
  NOR U5018 ( .A(n2851), .B(n2804), .Z(n5186) );
  AND U5019 ( .A(n5192), .B(n5193), .Z(n5034) );
  NANDN U5020 ( .A(n5039), .B(n5041), .Z(n5193) );
  NANDN U5021 ( .A(n5042), .B(n5194), .Z(n5192) );
  NANDN U5022 ( .A(n5041), .B(n5039), .Z(n5194) );
  XOR U5023 ( .A(n5195), .B(n5196), .Z(n5039) );
  XOR U5024 ( .A(n5197), .B(n5198), .Z(n5196) );
  AND U5025 ( .A(\stack[1][8] ), .B(\stack[0][9] ), .Z(n5041) );
  AND U5026 ( .A(n5199), .B(n5200), .Z(n5042) );
  NANDN U5027 ( .A(n5046), .B(n5201), .Z(n5200) );
  NANDN U5028 ( .A(n5049), .B(n5202), .Z(n5199) );
  NAND U5029 ( .A(n5048), .B(n5046), .Z(n5202) );
  XOR U5030 ( .A(n5203), .B(n5204), .Z(n5046) );
  XNOR U5031 ( .A(n5205), .B(n5206), .Z(n5204) );
  IV U5032 ( .A(n5201), .Z(n5048) );
  NOR U5033 ( .A(n2803), .B(n2804), .Z(n5201) );
  AND U5034 ( .A(n5207), .B(n5208), .Z(n5049) );
  NANDN U5035 ( .A(n5054), .B(n5056), .Z(n5208) );
  NANDN U5036 ( .A(n5057), .B(n5209), .Z(n5207) );
  NANDN U5037 ( .A(n5056), .B(n5054), .Z(n5209) );
  XOR U5038 ( .A(n5210), .B(n5211), .Z(n5054) );
  XOR U5039 ( .A(n5212), .B(n5213), .Z(n5211) );
  AND U5040 ( .A(\stack[0][7] ), .B(\stack[1][8] ), .Z(n5056) );
  AND U5041 ( .A(n5214), .B(n5215), .Z(n5057) );
  NANDN U5042 ( .A(n5061), .B(n5216), .Z(n5215) );
  NANDN U5043 ( .A(n5064), .B(n5217), .Z(n5214) );
  NAND U5044 ( .A(n5063), .B(n5061), .Z(n5217) );
  XOR U5045 ( .A(n5218), .B(n5219), .Z(n5061) );
  XNOR U5046 ( .A(n5220), .B(n5221), .Z(n5219) );
  IV U5047 ( .A(n5216), .Z(n5063) );
  NOR U5048 ( .A(n2755), .B(n2804), .Z(n5216) );
  AND U5049 ( .A(n5222), .B(n5223), .Z(n5064) );
  NANDN U5050 ( .A(n5069), .B(n5071), .Z(n5223) );
  NANDN U5051 ( .A(n5072), .B(n5224), .Z(n5222) );
  NANDN U5052 ( .A(n5071), .B(n5069), .Z(n5224) );
  XOR U5053 ( .A(n5225), .B(n5226), .Z(n5069) );
  XOR U5054 ( .A(n5227), .B(n5228), .Z(n5226) );
  AND U5055 ( .A(\stack[0][5] ), .B(\stack[1][8] ), .Z(n5071) );
  AND U5056 ( .A(n5229), .B(n5230), .Z(n5072) );
  NANDN U5057 ( .A(n5076), .B(n5231), .Z(n5230) );
  NANDN U5058 ( .A(n5079), .B(n5232), .Z(n5229) );
  NAND U5059 ( .A(n5078), .B(n5076), .Z(n5232) );
  XOR U5060 ( .A(n5233), .B(n5234), .Z(n5076) );
  XNOR U5061 ( .A(n5235), .B(n5236), .Z(n5234) );
  IV U5062 ( .A(n5231), .Z(n5078) );
  NOR U5063 ( .A(n2707), .B(n2804), .Z(n5231) );
  IV U5064 ( .A(\stack[1][8] ), .Z(n2804) );
  AND U5065 ( .A(n5237), .B(n5238), .Z(n5079) );
  NANDN U5066 ( .A(n5084), .B(n5086), .Z(n5238) );
  NANDN U5067 ( .A(n5087), .B(n5239), .Z(n5237) );
  NANDN U5068 ( .A(n5086), .B(n5084), .Z(n5239) );
  XNOR U5069 ( .A(n5240), .B(n5241), .Z(n5084) );
  XNOR U5070 ( .A(n5242), .B(n5243), .Z(n5241) );
  AND U5071 ( .A(\stack[0][3] ), .B(\stack[1][8] ), .Z(n5086) );
  AND U5072 ( .A(n5244), .B(n5245), .Z(n5087) );
  NANDN U5073 ( .A(n5091), .B(n5093), .Z(n5245) );
  NANDN U5074 ( .A(n5094), .B(n5246), .Z(n5244) );
  NANDN U5075 ( .A(n5093), .B(n5091), .Z(n5246) );
  XNOR U5076 ( .A(n5247), .B(n5248), .Z(n5091) );
  NAND U5077 ( .A(\stack[0][0] ), .B(\stack[1][10] ), .Z(n5248) );
  AND U5078 ( .A(\stack[0][2] ), .B(\stack[1][8] ), .Z(n5093) );
  NANDN U5079 ( .A(n5098), .B(n5249), .Z(n5094) );
  AND U5080 ( .A(\stack[1][9] ), .B(\stack[0][0] ), .Z(n5249) );
  NAND U5081 ( .A(\stack[1][8] ), .B(\stack[0][1] ), .Z(n5098) );
  ANDN U5082 ( .B(\stack[1][8] ), .A(n3139), .Z(n3586) );
  IV U5083 ( .A(\stack[0][22] ), .Z(n3139) );
  XNOR U5084 ( .A(n3596), .B(n5250), .Z(n3585) );
  XNOR U5085 ( .A(n3595), .B(n3597), .Z(n5250) );
  AND U5086 ( .A(n5251), .B(n5252), .Z(n3597) );
  NANDN U5087 ( .A(n5105), .B(n5253), .Z(n5252) );
  NANDN U5088 ( .A(n5108), .B(n5254), .Z(n5251) );
  NAND U5089 ( .A(n5107), .B(n5105), .Z(n5254) );
  XOR U5090 ( .A(n5255), .B(n5256), .Z(n5105) );
  XNOR U5091 ( .A(n5257), .B(n5258), .Z(n5256) );
  IV U5092 ( .A(n5253), .Z(n5107) );
  NOR U5093 ( .A(n3091), .B(n2828), .Z(n5253) );
  IV U5094 ( .A(\stack[0][20] ), .Z(n3091) );
  AND U5095 ( .A(n5259), .B(n5260), .Z(n5108) );
  NANDN U5096 ( .A(n5113), .B(n5115), .Z(n5260) );
  NANDN U5097 ( .A(n5116), .B(n5261), .Z(n5259) );
  NANDN U5098 ( .A(n5115), .B(n5113), .Z(n5261) );
  XOR U5099 ( .A(n5262), .B(n5263), .Z(n5113) );
  XOR U5100 ( .A(n5264), .B(n5265), .Z(n5263) );
  AND U5101 ( .A(\stack[0][19] ), .B(\stack[1][9] ), .Z(n5115) );
  AND U5102 ( .A(n5266), .B(n5267), .Z(n5116) );
  NANDN U5103 ( .A(n5120), .B(n5268), .Z(n5267) );
  NANDN U5104 ( .A(n5123), .B(n5269), .Z(n5266) );
  NAND U5105 ( .A(n5122), .B(n5120), .Z(n5269) );
  XOR U5106 ( .A(n5270), .B(n5271), .Z(n5120) );
  XNOR U5107 ( .A(n5272), .B(n5273), .Z(n5271) );
  IV U5108 ( .A(n5268), .Z(n5122) );
  NOR U5109 ( .A(n3043), .B(n2828), .Z(n5268) );
  AND U5110 ( .A(n5274), .B(n5275), .Z(n5123) );
  NANDN U5111 ( .A(n5128), .B(n5130), .Z(n5275) );
  NANDN U5112 ( .A(n5131), .B(n5276), .Z(n5274) );
  NANDN U5113 ( .A(n5130), .B(n5128), .Z(n5276) );
  XOR U5114 ( .A(n5277), .B(n5278), .Z(n5128) );
  XOR U5115 ( .A(n5279), .B(n5280), .Z(n5278) );
  AND U5116 ( .A(\stack[0][17] ), .B(\stack[1][9] ), .Z(n5130) );
  AND U5117 ( .A(n5281), .B(n5282), .Z(n5131) );
  NANDN U5118 ( .A(n5135), .B(n5283), .Z(n5282) );
  NANDN U5119 ( .A(n5138), .B(n5284), .Z(n5281) );
  NAND U5120 ( .A(n5137), .B(n5135), .Z(n5284) );
  XOR U5121 ( .A(n5285), .B(n5286), .Z(n5135) );
  XNOR U5122 ( .A(n5287), .B(n5288), .Z(n5286) );
  IV U5123 ( .A(n5283), .Z(n5137) );
  NOR U5124 ( .A(n2995), .B(n2828), .Z(n5283) );
  AND U5125 ( .A(n5289), .B(n5290), .Z(n5138) );
  NANDN U5126 ( .A(n5143), .B(n5145), .Z(n5290) );
  NANDN U5127 ( .A(n5146), .B(n5291), .Z(n5289) );
  NANDN U5128 ( .A(n5145), .B(n5143), .Z(n5291) );
  XOR U5129 ( .A(n5292), .B(n5293), .Z(n5143) );
  XOR U5130 ( .A(n5294), .B(n5295), .Z(n5293) );
  AND U5131 ( .A(\stack[0][15] ), .B(\stack[1][9] ), .Z(n5145) );
  AND U5132 ( .A(n5296), .B(n5297), .Z(n5146) );
  NANDN U5133 ( .A(n5150), .B(n5298), .Z(n5297) );
  NANDN U5134 ( .A(n5153), .B(n5299), .Z(n5296) );
  NAND U5135 ( .A(n5152), .B(n5150), .Z(n5299) );
  XOR U5136 ( .A(n5300), .B(n5301), .Z(n5150) );
  XNOR U5137 ( .A(n5302), .B(n5303), .Z(n5301) );
  IV U5138 ( .A(n5298), .Z(n5152) );
  NOR U5139 ( .A(n2947), .B(n2828), .Z(n5298) );
  AND U5140 ( .A(n5304), .B(n5305), .Z(n5153) );
  NANDN U5141 ( .A(n5158), .B(n5160), .Z(n5305) );
  NANDN U5142 ( .A(n5161), .B(n5306), .Z(n5304) );
  NANDN U5143 ( .A(n5160), .B(n5158), .Z(n5306) );
  XOR U5144 ( .A(n5307), .B(n5308), .Z(n5158) );
  XOR U5145 ( .A(n5309), .B(n5310), .Z(n5308) );
  AND U5146 ( .A(\stack[0][13] ), .B(\stack[1][9] ), .Z(n5160) );
  AND U5147 ( .A(n5311), .B(n5312), .Z(n5161) );
  NANDN U5148 ( .A(n5165), .B(n5313), .Z(n5312) );
  NANDN U5149 ( .A(n5168), .B(n5314), .Z(n5311) );
  NAND U5150 ( .A(n5167), .B(n5165), .Z(n5314) );
  XOR U5151 ( .A(n5315), .B(n5316), .Z(n5165) );
  XNOR U5152 ( .A(n5317), .B(n5318), .Z(n5316) );
  IV U5153 ( .A(n5313), .Z(n5167) );
  NOR U5154 ( .A(n2899), .B(n2828), .Z(n5313) );
  AND U5155 ( .A(n5319), .B(n5320), .Z(n5168) );
  NANDN U5156 ( .A(n5173), .B(n5175), .Z(n5320) );
  NANDN U5157 ( .A(n5176), .B(n5321), .Z(n5319) );
  NANDN U5158 ( .A(n5175), .B(n5173), .Z(n5321) );
  XOR U5159 ( .A(n5322), .B(n5323), .Z(n5173) );
  XOR U5160 ( .A(n5324), .B(n5325), .Z(n5323) );
  AND U5161 ( .A(\stack[0][11] ), .B(\stack[1][9] ), .Z(n5175) );
  AND U5162 ( .A(n5326), .B(n5327), .Z(n5176) );
  NANDN U5163 ( .A(n5180), .B(n5328), .Z(n5327) );
  NANDN U5164 ( .A(n5183), .B(n5329), .Z(n5326) );
  NAND U5165 ( .A(n5182), .B(n5180), .Z(n5329) );
  XOR U5166 ( .A(n5330), .B(n5331), .Z(n5180) );
  XNOR U5167 ( .A(n5332), .B(n5333), .Z(n5331) );
  IV U5168 ( .A(n5328), .Z(n5182) );
  NOR U5169 ( .A(n2851), .B(n2828), .Z(n5328) );
  AND U5170 ( .A(n5334), .B(n5335), .Z(n5183) );
  NANDN U5171 ( .A(n5188), .B(n5190), .Z(n5335) );
  NANDN U5172 ( .A(n5191), .B(n5336), .Z(n5334) );
  NANDN U5173 ( .A(n5190), .B(n5188), .Z(n5336) );
  XOR U5174 ( .A(n5337), .B(n5338), .Z(n5188) );
  XOR U5175 ( .A(n5339), .B(n5340), .Z(n5338) );
  AND U5176 ( .A(\stack[1][9] ), .B(\stack[0][9] ), .Z(n5190) );
  AND U5177 ( .A(n5341), .B(n5342), .Z(n5191) );
  NANDN U5178 ( .A(n5195), .B(n5343), .Z(n5342) );
  NANDN U5179 ( .A(n5198), .B(n5344), .Z(n5341) );
  NAND U5180 ( .A(n5197), .B(n5195), .Z(n5344) );
  XOR U5181 ( .A(n5345), .B(n5346), .Z(n5195) );
  XNOR U5182 ( .A(n5347), .B(n5348), .Z(n5346) );
  IV U5183 ( .A(n5343), .Z(n5197) );
  NOR U5184 ( .A(n2803), .B(n2828), .Z(n5343) );
  AND U5185 ( .A(n5349), .B(n5350), .Z(n5198) );
  NANDN U5186 ( .A(n5203), .B(n5205), .Z(n5350) );
  NANDN U5187 ( .A(n5206), .B(n5351), .Z(n5349) );
  NANDN U5188 ( .A(n5205), .B(n5203), .Z(n5351) );
  XOR U5189 ( .A(n5352), .B(n5353), .Z(n5203) );
  XOR U5190 ( .A(n5354), .B(n5355), .Z(n5353) );
  AND U5191 ( .A(\stack[0][7] ), .B(\stack[1][9] ), .Z(n5205) );
  AND U5192 ( .A(n5356), .B(n5357), .Z(n5206) );
  NANDN U5193 ( .A(n5210), .B(n5358), .Z(n5357) );
  NANDN U5194 ( .A(n5213), .B(n5359), .Z(n5356) );
  NAND U5195 ( .A(n5212), .B(n5210), .Z(n5359) );
  XOR U5196 ( .A(n5360), .B(n5361), .Z(n5210) );
  XNOR U5197 ( .A(n5362), .B(n5363), .Z(n5361) );
  IV U5198 ( .A(n5358), .Z(n5212) );
  NOR U5199 ( .A(n2755), .B(n2828), .Z(n5358) );
  AND U5200 ( .A(n5364), .B(n5365), .Z(n5213) );
  NANDN U5201 ( .A(n5218), .B(n5220), .Z(n5365) );
  NANDN U5202 ( .A(n5221), .B(n5366), .Z(n5364) );
  NANDN U5203 ( .A(n5220), .B(n5218), .Z(n5366) );
  XOR U5204 ( .A(n5367), .B(n5368), .Z(n5218) );
  XOR U5205 ( .A(n5369), .B(n5370), .Z(n5368) );
  AND U5206 ( .A(\stack[0][5] ), .B(\stack[1][9] ), .Z(n5220) );
  AND U5207 ( .A(n5371), .B(n5372), .Z(n5221) );
  NANDN U5208 ( .A(n5225), .B(n5373), .Z(n5372) );
  NANDN U5209 ( .A(n5228), .B(n5374), .Z(n5371) );
  NAND U5210 ( .A(n5227), .B(n5225), .Z(n5374) );
  XOR U5211 ( .A(n5375), .B(n5376), .Z(n5225) );
  XNOR U5212 ( .A(n5377), .B(n5378), .Z(n5376) );
  IV U5213 ( .A(n5373), .Z(n5227) );
  NOR U5214 ( .A(n2707), .B(n2828), .Z(n5373) );
  AND U5215 ( .A(n5379), .B(n5380), .Z(n5228) );
  NANDN U5216 ( .A(n5233), .B(n5235), .Z(n5380) );
  NANDN U5217 ( .A(n5236), .B(n5381), .Z(n5379) );
  NANDN U5218 ( .A(n5235), .B(n5233), .Z(n5381) );
  XNOR U5219 ( .A(n5382), .B(n5383), .Z(n5233) );
  XNOR U5220 ( .A(n5384), .B(n5385), .Z(n5383) );
  AND U5221 ( .A(\stack[0][3] ), .B(\stack[1][9] ), .Z(n5235) );
  AND U5222 ( .A(n5386), .B(n5387), .Z(n5236) );
  NANDN U5223 ( .A(n5240), .B(n5242), .Z(n5387) );
  NAND U5224 ( .A(n5388), .B(n5243), .Z(n5386) );
  ANDN U5225 ( .B(n5389), .A(n5247), .Z(n5243) );
  NAND U5226 ( .A(\stack[1][9] ), .B(\stack[0][1] ), .Z(n5247) );
  AND U5227 ( .A(\stack[0][0] ), .B(\stack[1][10] ), .Z(n5389) );
  NANDN U5228 ( .A(n5242), .B(n5240), .Z(n5388) );
  XNOR U5229 ( .A(n5390), .B(n5391), .Z(n5240) );
  NAND U5230 ( .A(\stack[0][0] ), .B(\stack[1][11] ), .Z(n5391) );
  AND U5231 ( .A(\stack[0][2] ), .B(\stack[1][9] ), .Z(n5242) );
  NOR U5232 ( .A(n3115), .B(n2828), .Z(n3595) );
  IV U5233 ( .A(\stack[1][9] ), .Z(n2828) );
  IV U5234 ( .A(\stack[0][21] ), .Z(n3115) );
  XNOR U5235 ( .A(n3603), .B(n5392), .Z(n3596) );
  XNOR U5236 ( .A(n3604), .B(n3605), .Z(n5392) );
  AND U5237 ( .A(n5393), .B(n5394), .Z(n3605) );
  NANDN U5238 ( .A(n5255), .B(n5257), .Z(n5394) );
  NANDN U5239 ( .A(n5258), .B(n5395), .Z(n5393) );
  NANDN U5240 ( .A(n5257), .B(n5255), .Z(n5395) );
  XOR U5241 ( .A(n5396), .B(n5397), .Z(n5255) );
  XOR U5242 ( .A(n5398), .B(n5399), .Z(n5397) );
  AND U5243 ( .A(\stack[1][10] ), .B(\stack[0][19] ), .Z(n5257) );
  AND U5244 ( .A(n5400), .B(n5401), .Z(n5258) );
  NANDN U5245 ( .A(n5262), .B(n5402), .Z(n5401) );
  NANDN U5246 ( .A(n5265), .B(n5403), .Z(n5400) );
  NAND U5247 ( .A(n5264), .B(n5262), .Z(n5403) );
  XOR U5248 ( .A(n5404), .B(n5405), .Z(n5262) );
  XNOR U5249 ( .A(n5406), .B(n5407), .Z(n5405) );
  IV U5250 ( .A(n5402), .Z(n5264) );
  NOR U5251 ( .A(n2852), .B(n3043), .Z(n5402) );
  AND U5252 ( .A(n5408), .B(n5409), .Z(n5265) );
  NANDN U5253 ( .A(n5270), .B(n5272), .Z(n5409) );
  NANDN U5254 ( .A(n5273), .B(n5410), .Z(n5408) );
  NANDN U5255 ( .A(n5272), .B(n5270), .Z(n5410) );
  XOR U5256 ( .A(n5411), .B(n5412), .Z(n5270) );
  XOR U5257 ( .A(n5413), .B(n5414), .Z(n5412) );
  AND U5258 ( .A(\stack[1][10] ), .B(\stack[0][17] ), .Z(n5272) );
  AND U5259 ( .A(n5415), .B(n5416), .Z(n5273) );
  NANDN U5260 ( .A(n5277), .B(n5417), .Z(n5416) );
  NANDN U5261 ( .A(n5280), .B(n5418), .Z(n5415) );
  NAND U5262 ( .A(n5279), .B(n5277), .Z(n5418) );
  XOR U5263 ( .A(n5419), .B(n5420), .Z(n5277) );
  XNOR U5264 ( .A(n5421), .B(n5422), .Z(n5420) );
  IV U5265 ( .A(n5417), .Z(n5279) );
  NOR U5266 ( .A(n2852), .B(n2995), .Z(n5417) );
  AND U5267 ( .A(n5423), .B(n5424), .Z(n5280) );
  NANDN U5268 ( .A(n5285), .B(n5287), .Z(n5424) );
  NANDN U5269 ( .A(n5288), .B(n5425), .Z(n5423) );
  NANDN U5270 ( .A(n5287), .B(n5285), .Z(n5425) );
  XOR U5271 ( .A(n5426), .B(n5427), .Z(n5285) );
  XOR U5272 ( .A(n5428), .B(n5429), .Z(n5427) );
  AND U5273 ( .A(\stack[1][10] ), .B(\stack[0][15] ), .Z(n5287) );
  AND U5274 ( .A(n5430), .B(n5431), .Z(n5288) );
  NANDN U5275 ( .A(n5292), .B(n5432), .Z(n5431) );
  NANDN U5276 ( .A(n5295), .B(n5433), .Z(n5430) );
  NAND U5277 ( .A(n5294), .B(n5292), .Z(n5433) );
  XOR U5278 ( .A(n5434), .B(n5435), .Z(n5292) );
  XNOR U5279 ( .A(n5436), .B(n5437), .Z(n5435) );
  IV U5280 ( .A(n5432), .Z(n5294) );
  NOR U5281 ( .A(n2852), .B(n2947), .Z(n5432) );
  AND U5282 ( .A(n5438), .B(n5439), .Z(n5295) );
  NANDN U5283 ( .A(n5300), .B(n5302), .Z(n5439) );
  NANDN U5284 ( .A(n5303), .B(n5440), .Z(n5438) );
  NANDN U5285 ( .A(n5302), .B(n5300), .Z(n5440) );
  XOR U5286 ( .A(n5441), .B(n5442), .Z(n5300) );
  XOR U5287 ( .A(n5443), .B(n5444), .Z(n5442) );
  AND U5288 ( .A(\stack[1][10] ), .B(\stack[0][13] ), .Z(n5302) );
  AND U5289 ( .A(n5445), .B(n5446), .Z(n5303) );
  NANDN U5290 ( .A(n5307), .B(n5447), .Z(n5446) );
  NANDN U5291 ( .A(n5310), .B(n5448), .Z(n5445) );
  NAND U5292 ( .A(n5309), .B(n5307), .Z(n5448) );
  XOR U5293 ( .A(n5449), .B(n5450), .Z(n5307) );
  XNOR U5294 ( .A(n5451), .B(n5452), .Z(n5450) );
  IV U5295 ( .A(n5447), .Z(n5309) );
  NOR U5296 ( .A(n2852), .B(n2899), .Z(n5447) );
  AND U5297 ( .A(n5453), .B(n5454), .Z(n5310) );
  NANDN U5298 ( .A(n5315), .B(n5317), .Z(n5454) );
  NANDN U5299 ( .A(n5318), .B(n5455), .Z(n5453) );
  NANDN U5300 ( .A(n5317), .B(n5315), .Z(n5455) );
  XOR U5301 ( .A(n5456), .B(n5457), .Z(n5315) );
  XOR U5302 ( .A(n5458), .B(n5459), .Z(n5457) );
  AND U5303 ( .A(\stack[1][10] ), .B(\stack[0][11] ), .Z(n5317) );
  AND U5304 ( .A(n5460), .B(n5461), .Z(n5318) );
  NANDN U5305 ( .A(n5322), .B(n5462), .Z(n5461) );
  NANDN U5306 ( .A(n5325), .B(n5463), .Z(n5460) );
  NAND U5307 ( .A(n5324), .B(n5322), .Z(n5463) );
  XOR U5308 ( .A(n5464), .B(n5465), .Z(n5322) );
  XNOR U5309 ( .A(n5466), .B(n5467), .Z(n5465) );
  IV U5310 ( .A(n5462), .Z(n5324) );
  NOR U5311 ( .A(n2852), .B(n2851), .Z(n5462) );
  AND U5312 ( .A(n5468), .B(n5469), .Z(n5325) );
  NANDN U5313 ( .A(n5330), .B(n5332), .Z(n5469) );
  NANDN U5314 ( .A(n5333), .B(n5470), .Z(n5468) );
  NANDN U5315 ( .A(n5332), .B(n5330), .Z(n5470) );
  XOR U5316 ( .A(n5471), .B(n5472), .Z(n5330) );
  XOR U5317 ( .A(n5473), .B(n5474), .Z(n5472) );
  AND U5318 ( .A(\stack[1][10] ), .B(\stack[0][9] ), .Z(n5332) );
  AND U5319 ( .A(n5475), .B(n5476), .Z(n5333) );
  NANDN U5320 ( .A(n5337), .B(n5477), .Z(n5476) );
  NANDN U5321 ( .A(n5340), .B(n5478), .Z(n5475) );
  NAND U5322 ( .A(n5339), .B(n5337), .Z(n5478) );
  XOR U5323 ( .A(n5479), .B(n5480), .Z(n5337) );
  XNOR U5324 ( .A(n5481), .B(n5482), .Z(n5480) );
  IV U5325 ( .A(n5477), .Z(n5339) );
  NOR U5326 ( .A(n2852), .B(n2803), .Z(n5477) );
  AND U5327 ( .A(n5483), .B(n5484), .Z(n5340) );
  NANDN U5328 ( .A(n5345), .B(n5347), .Z(n5484) );
  NANDN U5329 ( .A(n5348), .B(n5485), .Z(n5483) );
  NANDN U5330 ( .A(n5347), .B(n5345), .Z(n5485) );
  XOR U5331 ( .A(n5486), .B(n5487), .Z(n5345) );
  XOR U5332 ( .A(n5488), .B(n5489), .Z(n5487) );
  AND U5333 ( .A(\stack[1][10] ), .B(\stack[0][7] ), .Z(n5347) );
  AND U5334 ( .A(n5490), .B(n5491), .Z(n5348) );
  NANDN U5335 ( .A(n5352), .B(n5492), .Z(n5491) );
  NANDN U5336 ( .A(n5355), .B(n5493), .Z(n5490) );
  NAND U5337 ( .A(n5354), .B(n5352), .Z(n5493) );
  XOR U5338 ( .A(n5494), .B(n5495), .Z(n5352) );
  XNOR U5339 ( .A(n5496), .B(n5497), .Z(n5495) );
  IV U5340 ( .A(n5492), .Z(n5354) );
  NOR U5341 ( .A(n2852), .B(n2755), .Z(n5492) );
  AND U5342 ( .A(n5498), .B(n5499), .Z(n5355) );
  NANDN U5343 ( .A(n5360), .B(n5362), .Z(n5499) );
  NANDN U5344 ( .A(n5363), .B(n5500), .Z(n5498) );
  NANDN U5345 ( .A(n5362), .B(n5360), .Z(n5500) );
  XOR U5346 ( .A(n5501), .B(n5502), .Z(n5360) );
  XOR U5347 ( .A(n5503), .B(n5504), .Z(n5502) );
  AND U5348 ( .A(\stack[1][10] ), .B(\stack[0][5] ), .Z(n5362) );
  AND U5349 ( .A(n5505), .B(n5506), .Z(n5363) );
  NANDN U5350 ( .A(n5367), .B(n5507), .Z(n5506) );
  NANDN U5351 ( .A(n5370), .B(n5508), .Z(n5505) );
  NAND U5352 ( .A(n5369), .B(n5367), .Z(n5508) );
  XOR U5353 ( .A(n5509), .B(n5510), .Z(n5367) );
  XNOR U5354 ( .A(n5511), .B(n5512), .Z(n5510) );
  IV U5355 ( .A(n5507), .Z(n5369) );
  NOR U5356 ( .A(n2852), .B(n2707), .Z(n5507) );
  AND U5357 ( .A(n5513), .B(n5514), .Z(n5370) );
  NANDN U5358 ( .A(n5375), .B(n5377), .Z(n5514) );
  NANDN U5359 ( .A(n5378), .B(n5515), .Z(n5513) );
  NANDN U5360 ( .A(n5377), .B(n5375), .Z(n5515) );
  XNOR U5361 ( .A(n5516), .B(n5517), .Z(n5375) );
  XNOR U5362 ( .A(n5518), .B(n5519), .Z(n5517) );
  AND U5363 ( .A(\stack[1][10] ), .B(\stack[0][3] ), .Z(n5377) );
  AND U5364 ( .A(n5520), .B(n5521), .Z(n5378) );
  NANDN U5365 ( .A(n5382), .B(n5384), .Z(n5521) );
  NAND U5366 ( .A(n5522), .B(n5385), .Z(n5520) );
  ANDN U5367 ( .B(n5523), .A(n5390), .Z(n5385) );
  NAND U5368 ( .A(\stack[1][10] ), .B(\stack[0][1] ), .Z(n5390) );
  AND U5369 ( .A(\stack[0][0] ), .B(\stack[1][11] ), .Z(n5523) );
  NANDN U5370 ( .A(n5384), .B(n5382), .Z(n5522) );
  XNOR U5371 ( .A(n5524), .B(n5525), .Z(n5382) );
  NAND U5372 ( .A(\stack[0][0] ), .B(\stack[1][12] ), .Z(n5525) );
  AND U5373 ( .A(\stack[1][10] ), .B(\stack[0][2] ), .Z(n5384) );
  ANDN U5374 ( .B(\stack[0][20] ), .A(n2852), .Z(n3604) );
  IV U5375 ( .A(\stack[1][10] ), .Z(n2852) );
  XNOR U5376 ( .A(n3408), .B(n5526), .Z(n3603) );
  XNOR U5377 ( .A(n3407), .B(n3409), .Z(n5526) );
  AND U5378 ( .A(n5527), .B(n5528), .Z(n3409) );
  NANDN U5379 ( .A(n5396), .B(n5529), .Z(n5528) );
  NANDN U5380 ( .A(n5399), .B(n5530), .Z(n5527) );
  NAND U5381 ( .A(n5398), .B(n5396), .Z(n5530) );
  XOR U5382 ( .A(n5531), .B(n5532), .Z(n5396) );
  XNOR U5383 ( .A(n5533), .B(n5534), .Z(n5532) );
  IV U5384 ( .A(n5529), .Z(n5398) );
  NOR U5385 ( .A(n2876), .B(n3043), .Z(n5529) );
  IV U5386 ( .A(\stack[0][18] ), .Z(n3043) );
  AND U5387 ( .A(n5535), .B(n5536), .Z(n5399) );
  NANDN U5388 ( .A(n5404), .B(n5406), .Z(n5536) );
  NANDN U5389 ( .A(n5407), .B(n5537), .Z(n5535) );
  NANDN U5390 ( .A(n5406), .B(n5404), .Z(n5537) );
  XOR U5391 ( .A(n5538), .B(n5539), .Z(n5404) );
  XOR U5392 ( .A(n5540), .B(n5541), .Z(n5539) );
  AND U5393 ( .A(\stack[1][11] ), .B(\stack[0][17] ), .Z(n5406) );
  AND U5394 ( .A(n5542), .B(n5543), .Z(n5407) );
  NANDN U5395 ( .A(n5411), .B(n5544), .Z(n5543) );
  NANDN U5396 ( .A(n5414), .B(n5545), .Z(n5542) );
  NAND U5397 ( .A(n5413), .B(n5411), .Z(n5545) );
  XOR U5398 ( .A(n5546), .B(n5547), .Z(n5411) );
  XNOR U5399 ( .A(n5548), .B(n5549), .Z(n5547) );
  IV U5400 ( .A(n5544), .Z(n5413) );
  NOR U5401 ( .A(n2876), .B(n2995), .Z(n5544) );
  AND U5402 ( .A(n5550), .B(n5551), .Z(n5414) );
  NANDN U5403 ( .A(n5419), .B(n5421), .Z(n5551) );
  NANDN U5404 ( .A(n5422), .B(n5552), .Z(n5550) );
  NANDN U5405 ( .A(n5421), .B(n5419), .Z(n5552) );
  XOR U5406 ( .A(n5553), .B(n5554), .Z(n5419) );
  XOR U5407 ( .A(n5555), .B(n5556), .Z(n5554) );
  AND U5408 ( .A(\stack[1][11] ), .B(\stack[0][15] ), .Z(n5421) );
  AND U5409 ( .A(n5557), .B(n5558), .Z(n5422) );
  NANDN U5410 ( .A(n5426), .B(n5559), .Z(n5558) );
  NANDN U5411 ( .A(n5429), .B(n5560), .Z(n5557) );
  NAND U5412 ( .A(n5428), .B(n5426), .Z(n5560) );
  XOR U5413 ( .A(n5561), .B(n5562), .Z(n5426) );
  XNOR U5414 ( .A(n5563), .B(n5564), .Z(n5562) );
  IV U5415 ( .A(n5559), .Z(n5428) );
  NOR U5416 ( .A(n2876), .B(n2947), .Z(n5559) );
  AND U5417 ( .A(n5565), .B(n5566), .Z(n5429) );
  NANDN U5418 ( .A(n5434), .B(n5436), .Z(n5566) );
  NANDN U5419 ( .A(n5437), .B(n5567), .Z(n5565) );
  NANDN U5420 ( .A(n5436), .B(n5434), .Z(n5567) );
  XOR U5421 ( .A(n5568), .B(n5569), .Z(n5434) );
  XOR U5422 ( .A(n5570), .B(n5571), .Z(n5569) );
  AND U5423 ( .A(\stack[1][11] ), .B(\stack[0][13] ), .Z(n5436) );
  AND U5424 ( .A(n5572), .B(n5573), .Z(n5437) );
  NANDN U5425 ( .A(n5441), .B(n5574), .Z(n5573) );
  NANDN U5426 ( .A(n5444), .B(n5575), .Z(n5572) );
  NAND U5427 ( .A(n5443), .B(n5441), .Z(n5575) );
  XOR U5428 ( .A(n5576), .B(n5577), .Z(n5441) );
  XNOR U5429 ( .A(n5578), .B(n5579), .Z(n5577) );
  IV U5430 ( .A(n5574), .Z(n5443) );
  NOR U5431 ( .A(n2876), .B(n2899), .Z(n5574) );
  AND U5432 ( .A(n5580), .B(n5581), .Z(n5444) );
  NANDN U5433 ( .A(n5449), .B(n5451), .Z(n5581) );
  NANDN U5434 ( .A(n5452), .B(n5582), .Z(n5580) );
  NANDN U5435 ( .A(n5451), .B(n5449), .Z(n5582) );
  XOR U5436 ( .A(n5583), .B(n5584), .Z(n5449) );
  XOR U5437 ( .A(n5585), .B(n5586), .Z(n5584) );
  AND U5438 ( .A(\stack[1][11] ), .B(\stack[0][11] ), .Z(n5451) );
  AND U5439 ( .A(n5587), .B(n5588), .Z(n5452) );
  NANDN U5440 ( .A(n5456), .B(n5589), .Z(n5588) );
  NANDN U5441 ( .A(n5459), .B(n5590), .Z(n5587) );
  NAND U5442 ( .A(n5458), .B(n5456), .Z(n5590) );
  XOR U5443 ( .A(n5591), .B(n5592), .Z(n5456) );
  XNOR U5444 ( .A(n5593), .B(n5594), .Z(n5592) );
  IV U5445 ( .A(n5589), .Z(n5458) );
  NOR U5446 ( .A(n2876), .B(n2851), .Z(n5589) );
  AND U5447 ( .A(n5595), .B(n5596), .Z(n5459) );
  NANDN U5448 ( .A(n5464), .B(n5466), .Z(n5596) );
  NANDN U5449 ( .A(n5467), .B(n5597), .Z(n5595) );
  NANDN U5450 ( .A(n5466), .B(n5464), .Z(n5597) );
  XOR U5451 ( .A(n5598), .B(n5599), .Z(n5464) );
  XOR U5452 ( .A(n5600), .B(n5601), .Z(n5599) );
  AND U5453 ( .A(\stack[1][11] ), .B(\stack[0][9] ), .Z(n5466) );
  AND U5454 ( .A(n5602), .B(n5603), .Z(n5467) );
  NANDN U5455 ( .A(n5471), .B(n5604), .Z(n5603) );
  NANDN U5456 ( .A(n5474), .B(n5605), .Z(n5602) );
  NAND U5457 ( .A(n5473), .B(n5471), .Z(n5605) );
  XOR U5458 ( .A(n5606), .B(n5607), .Z(n5471) );
  XNOR U5459 ( .A(n5608), .B(n5609), .Z(n5607) );
  IV U5460 ( .A(n5604), .Z(n5473) );
  NOR U5461 ( .A(n2876), .B(n2803), .Z(n5604) );
  AND U5462 ( .A(n5610), .B(n5611), .Z(n5474) );
  NANDN U5463 ( .A(n5479), .B(n5481), .Z(n5611) );
  NANDN U5464 ( .A(n5482), .B(n5612), .Z(n5610) );
  NANDN U5465 ( .A(n5481), .B(n5479), .Z(n5612) );
  XOR U5466 ( .A(n5613), .B(n5614), .Z(n5479) );
  XOR U5467 ( .A(n5615), .B(n5616), .Z(n5614) );
  AND U5468 ( .A(\stack[1][11] ), .B(\stack[0][7] ), .Z(n5481) );
  AND U5469 ( .A(n5617), .B(n5618), .Z(n5482) );
  NANDN U5470 ( .A(n5486), .B(n5619), .Z(n5618) );
  NANDN U5471 ( .A(n5489), .B(n5620), .Z(n5617) );
  NAND U5472 ( .A(n5488), .B(n5486), .Z(n5620) );
  XOR U5473 ( .A(n5621), .B(n5622), .Z(n5486) );
  XNOR U5474 ( .A(n5623), .B(n5624), .Z(n5622) );
  IV U5475 ( .A(n5619), .Z(n5488) );
  NOR U5476 ( .A(n2876), .B(n2755), .Z(n5619) );
  AND U5477 ( .A(n5625), .B(n5626), .Z(n5489) );
  NANDN U5478 ( .A(n5494), .B(n5496), .Z(n5626) );
  NANDN U5479 ( .A(n5497), .B(n5627), .Z(n5625) );
  NANDN U5480 ( .A(n5496), .B(n5494), .Z(n5627) );
  XOR U5481 ( .A(n5628), .B(n5629), .Z(n5494) );
  XOR U5482 ( .A(n5630), .B(n5631), .Z(n5629) );
  AND U5483 ( .A(\stack[1][11] ), .B(\stack[0][5] ), .Z(n5496) );
  AND U5484 ( .A(n5632), .B(n5633), .Z(n5497) );
  NANDN U5485 ( .A(n5501), .B(n5634), .Z(n5633) );
  NANDN U5486 ( .A(n5504), .B(n5635), .Z(n5632) );
  NAND U5487 ( .A(n5503), .B(n5501), .Z(n5635) );
  XOR U5488 ( .A(n5636), .B(n5637), .Z(n5501) );
  XNOR U5489 ( .A(n5638), .B(n5639), .Z(n5637) );
  IV U5490 ( .A(n5634), .Z(n5503) );
  NOR U5491 ( .A(n2876), .B(n2707), .Z(n5634) );
  AND U5492 ( .A(n5640), .B(n5641), .Z(n5504) );
  NANDN U5493 ( .A(n5509), .B(n5511), .Z(n5641) );
  NANDN U5494 ( .A(n5512), .B(n5642), .Z(n5640) );
  NANDN U5495 ( .A(n5511), .B(n5509), .Z(n5642) );
  XNOR U5496 ( .A(n5643), .B(n5644), .Z(n5509) );
  XNOR U5497 ( .A(n5645), .B(n5646), .Z(n5644) );
  AND U5498 ( .A(\stack[1][11] ), .B(\stack[0][3] ), .Z(n5511) );
  AND U5499 ( .A(n5647), .B(n5648), .Z(n5512) );
  NANDN U5500 ( .A(n5516), .B(n5518), .Z(n5648) );
  NAND U5501 ( .A(n5649), .B(n5519), .Z(n5647) );
  ANDN U5502 ( .B(n5650), .A(n5524), .Z(n5519) );
  NAND U5503 ( .A(\stack[1][11] ), .B(\stack[0][1] ), .Z(n5524) );
  AND U5504 ( .A(\stack[0][0] ), .B(\stack[1][12] ), .Z(n5650) );
  NANDN U5505 ( .A(n5518), .B(n5516), .Z(n5649) );
  XNOR U5506 ( .A(n5651), .B(n5652), .Z(n5516) );
  NAND U5507 ( .A(\stack[0][0] ), .B(\stack[1][13] ), .Z(n5652) );
  AND U5508 ( .A(\stack[1][11] ), .B(\stack[0][2] ), .Z(n5518) );
  NOR U5509 ( .A(n2876), .B(n3067), .Z(n3407) );
  IV U5510 ( .A(\stack[0][19] ), .Z(n3067) );
  IV U5511 ( .A(\stack[1][11] ), .Z(n2876) );
  XNOR U5512 ( .A(n3559), .B(n5653), .Z(n3408) );
  XNOR U5513 ( .A(n3560), .B(n3561), .Z(n5653) );
  AND U5514 ( .A(n5654), .B(n5655), .Z(n3561) );
  NANDN U5515 ( .A(n5531), .B(n5533), .Z(n5655) );
  NANDN U5516 ( .A(n5534), .B(n5656), .Z(n5654) );
  NANDN U5517 ( .A(n5533), .B(n5531), .Z(n5656) );
  XOR U5518 ( .A(n5657), .B(n5658), .Z(n5531) );
  XOR U5519 ( .A(n5659), .B(n5660), .Z(n5658) );
  AND U5520 ( .A(\stack[1][12] ), .B(\stack[0][17] ), .Z(n5533) );
  AND U5521 ( .A(n5661), .B(n5662), .Z(n5534) );
  NANDN U5522 ( .A(n5538), .B(n5663), .Z(n5662) );
  NANDN U5523 ( .A(n5541), .B(n5664), .Z(n5661) );
  NAND U5524 ( .A(n5540), .B(n5538), .Z(n5664) );
  XOR U5525 ( .A(n5665), .B(n5666), .Z(n5538) );
  XNOR U5526 ( .A(n5667), .B(n5668), .Z(n5666) );
  IV U5527 ( .A(n5663), .Z(n5540) );
  NOR U5528 ( .A(n2900), .B(n2995), .Z(n5663) );
  AND U5529 ( .A(n5669), .B(n5670), .Z(n5541) );
  NANDN U5530 ( .A(n5546), .B(n5548), .Z(n5670) );
  NANDN U5531 ( .A(n5549), .B(n5671), .Z(n5669) );
  NANDN U5532 ( .A(n5548), .B(n5546), .Z(n5671) );
  XOR U5533 ( .A(n5672), .B(n5673), .Z(n5546) );
  XOR U5534 ( .A(n5674), .B(n5675), .Z(n5673) );
  AND U5535 ( .A(\stack[1][12] ), .B(\stack[0][15] ), .Z(n5548) );
  AND U5536 ( .A(n5676), .B(n5677), .Z(n5549) );
  NANDN U5537 ( .A(n5553), .B(n5678), .Z(n5677) );
  NANDN U5538 ( .A(n5556), .B(n5679), .Z(n5676) );
  NAND U5539 ( .A(n5555), .B(n5553), .Z(n5679) );
  XOR U5540 ( .A(n5680), .B(n5681), .Z(n5553) );
  XNOR U5541 ( .A(n5682), .B(n5683), .Z(n5681) );
  IV U5542 ( .A(n5678), .Z(n5555) );
  NOR U5543 ( .A(n2900), .B(n2947), .Z(n5678) );
  AND U5544 ( .A(n5684), .B(n5685), .Z(n5556) );
  NANDN U5545 ( .A(n5561), .B(n5563), .Z(n5685) );
  NANDN U5546 ( .A(n5564), .B(n5686), .Z(n5684) );
  NANDN U5547 ( .A(n5563), .B(n5561), .Z(n5686) );
  XOR U5548 ( .A(n5687), .B(n5688), .Z(n5561) );
  XOR U5549 ( .A(n5689), .B(n5690), .Z(n5688) );
  AND U5550 ( .A(\stack[1][12] ), .B(\stack[0][13] ), .Z(n5563) );
  AND U5551 ( .A(n5691), .B(n5692), .Z(n5564) );
  NANDN U5552 ( .A(n5568), .B(n5693), .Z(n5692) );
  NANDN U5553 ( .A(n5571), .B(n5694), .Z(n5691) );
  NAND U5554 ( .A(n5570), .B(n5568), .Z(n5694) );
  XOR U5555 ( .A(n5695), .B(n5696), .Z(n5568) );
  XNOR U5556 ( .A(n5697), .B(n5698), .Z(n5696) );
  IV U5557 ( .A(n5693), .Z(n5570) );
  NOR U5558 ( .A(n2900), .B(n2899), .Z(n5693) );
  AND U5559 ( .A(n5699), .B(n5700), .Z(n5571) );
  NANDN U5560 ( .A(n5576), .B(n5578), .Z(n5700) );
  NANDN U5561 ( .A(n5579), .B(n5701), .Z(n5699) );
  NANDN U5562 ( .A(n5578), .B(n5576), .Z(n5701) );
  XOR U5563 ( .A(n5702), .B(n5703), .Z(n5576) );
  XOR U5564 ( .A(n5704), .B(n5705), .Z(n5703) );
  AND U5565 ( .A(\stack[1][12] ), .B(\stack[0][11] ), .Z(n5578) );
  AND U5566 ( .A(n5706), .B(n5707), .Z(n5579) );
  NANDN U5567 ( .A(n5583), .B(n5708), .Z(n5707) );
  NANDN U5568 ( .A(n5586), .B(n5709), .Z(n5706) );
  NAND U5569 ( .A(n5585), .B(n5583), .Z(n5709) );
  XOR U5570 ( .A(n5710), .B(n5711), .Z(n5583) );
  XNOR U5571 ( .A(n5712), .B(n5713), .Z(n5711) );
  IV U5572 ( .A(n5708), .Z(n5585) );
  NOR U5573 ( .A(n2900), .B(n2851), .Z(n5708) );
  AND U5574 ( .A(n5714), .B(n5715), .Z(n5586) );
  NANDN U5575 ( .A(n5591), .B(n5593), .Z(n5715) );
  NANDN U5576 ( .A(n5594), .B(n5716), .Z(n5714) );
  NANDN U5577 ( .A(n5593), .B(n5591), .Z(n5716) );
  XOR U5578 ( .A(n5717), .B(n5718), .Z(n5591) );
  XOR U5579 ( .A(n5719), .B(n5720), .Z(n5718) );
  AND U5580 ( .A(\stack[1][12] ), .B(\stack[0][9] ), .Z(n5593) );
  AND U5581 ( .A(n5721), .B(n5722), .Z(n5594) );
  NANDN U5582 ( .A(n5598), .B(n5723), .Z(n5722) );
  NANDN U5583 ( .A(n5601), .B(n5724), .Z(n5721) );
  NAND U5584 ( .A(n5600), .B(n5598), .Z(n5724) );
  XOR U5585 ( .A(n5725), .B(n5726), .Z(n5598) );
  XNOR U5586 ( .A(n5727), .B(n5728), .Z(n5726) );
  IV U5587 ( .A(n5723), .Z(n5600) );
  NOR U5588 ( .A(n2900), .B(n2803), .Z(n5723) );
  AND U5589 ( .A(n5729), .B(n5730), .Z(n5601) );
  NANDN U5590 ( .A(n5606), .B(n5608), .Z(n5730) );
  NANDN U5591 ( .A(n5609), .B(n5731), .Z(n5729) );
  NANDN U5592 ( .A(n5608), .B(n5606), .Z(n5731) );
  XOR U5593 ( .A(n5732), .B(n5733), .Z(n5606) );
  XOR U5594 ( .A(n5734), .B(n5735), .Z(n5733) );
  AND U5595 ( .A(\stack[1][12] ), .B(\stack[0][7] ), .Z(n5608) );
  AND U5596 ( .A(n5736), .B(n5737), .Z(n5609) );
  NANDN U5597 ( .A(n5613), .B(n5738), .Z(n5737) );
  NANDN U5598 ( .A(n5616), .B(n5739), .Z(n5736) );
  NAND U5599 ( .A(n5615), .B(n5613), .Z(n5739) );
  XOR U5600 ( .A(n5740), .B(n5741), .Z(n5613) );
  XNOR U5601 ( .A(n5742), .B(n5743), .Z(n5741) );
  IV U5602 ( .A(n5738), .Z(n5615) );
  NOR U5603 ( .A(n2900), .B(n2755), .Z(n5738) );
  AND U5604 ( .A(n5744), .B(n5745), .Z(n5616) );
  NANDN U5605 ( .A(n5621), .B(n5623), .Z(n5745) );
  NANDN U5606 ( .A(n5624), .B(n5746), .Z(n5744) );
  NANDN U5607 ( .A(n5623), .B(n5621), .Z(n5746) );
  XOR U5608 ( .A(n5747), .B(n5748), .Z(n5621) );
  XOR U5609 ( .A(n5749), .B(n5750), .Z(n5748) );
  AND U5610 ( .A(\stack[1][12] ), .B(\stack[0][5] ), .Z(n5623) );
  AND U5611 ( .A(n5751), .B(n5752), .Z(n5624) );
  NANDN U5612 ( .A(n5628), .B(n5753), .Z(n5752) );
  NANDN U5613 ( .A(n5631), .B(n5754), .Z(n5751) );
  NAND U5614 ( .A(n5630), .B(n5628), .Z(n5754) );
  XOR U5615 ( .A(n5755), .B(n5756), .Z(n5628) );
  XNOR U5616 ( .A(n5757), .B(n5758), .Z(n5756) );
  IV U5617 ( .A(n5753), .Z(n5630) );
  NOR U5618 ( .A(n2900), .B(n2707), .Z(n5753) );
  AND U5619 ( .A(n5759), .B(n5760), .Z(n5631) );
  NANDN U5620 ( .A(n5636), .B(n5638), .Z(n5760) );
  NANDN U5621 ( .A(n5639), .B(n5761), .Z(n5759) );
  NANDN U5622 ( .A(n5638), .B(n5636), .Z(n5761) );
  XNOR U5623 ( .A(n5762), .B(n5763), .Z(n5636) );
  XNOR U5624 ( .A(n5764), .B(n5765), .Z(n5763) );
  AND U5625 ( .A(\stack[1][12] ), .B(\stack[0][3] ), .Z(n5638) );
  AND U5626 ( .A(n5766), .B(n5767), .Z(n5639) );
  NANDN U5627 ( .A(n5643), .B(n5645), .Z(n5767) );
  NAND U5628 ( .A(n5768), .B(n5646), .Z(n5766) );
  ANDN U5629 ( .B(n5769), .A(n5651), .Z(n5646) );
  NAND U5630 ( .A(\stack[1][12] ), .B(\stack[0][1] ), .Z(n5651) );
  AND U5631 ( .A(\stack[0][0] ), .B(\stack[1][13] ), .Z(n5769) );
  NANDN U5632 ( .A(n5645), .B(n5643), .Z(n5768) );
  XNOR U5633 ( .A(n5770), .B(n5771), .Z(n5643) );
  NAND U5634 ( .A(\stack[0][0] ), .B(\stack[1][14] ), .Z(n5771) );
  AND U5635 ( .A(\stack[1][12] ), .B(\stack[0][2] ), .Z(n5645) );
  ANDN U5636 ( .B(\stack[0][18] ), .A(n2900), .Z(n3560) );
  IV U5637 ( .A(\stack[1][12] ), .Z(n2900) );
  XNOR U5638 ( .A(n3570), .B(n5772), .Z(n3559) );
  XNOR U5639 ( .A(n3569), .B(n3571), .Z(n5772) );
  AND U5640 ( .A(n5773), .B(n5774), .Z(n3571) );
  NANDN U5641 ( .A(n5657), .B(n5775), .Z(n5774) );
  NANDN U5642 ( .A(n5660), .B(n5776), .Z(n5773) );
  NAND U5643 ( .A(n5659), .B(n5657), .Z(n5776) );
  XOR U5644 ( .A(n5777), .B(n5778), .Z(n5657) );
  XNOR U5645 ( .A(n5779), .B(n5780), .Z(n5778) );
  IV U5646 ( .A(n5775), .Z(n5659) );
  NOR U5647 ( .A(n2924), .B(n2995), .Z(n5775) );
  IV U5648 ( .A(\stack[0][16] ), .Z(n2995) );
  AND U5649 ( .A(n5781), .B(n5782), .Z(n5660) );
  NANDN U5650 ( .A(n5665), .B(n5667), .Z(n5782) );
  NANDN U5651 ( .A(n5668), .B(n5783), .Z(n5781) );
  NANDN U5652 ( .A(n5667), .B(n5665), .Z(n5783) );
  XOR U5653 ( .A(n5784), .B(n5785), .Z(n5665) );
  XOR U5654 ( .A(n5786), .B(n5787), .Z(n5785) );
  AND U5655 ( .A(\stack[1][13] ), .B(\stack[0][15] ), .Z(n5667) );
  AND U5656 ( .A(n5788), .B(n5789), .Z(n5668) );
  NANDN U5657 ( .A(n5672), .B(n5790), .Z(n5789) );
  NANDN U5658 ( .A(n5675), .B(n5791), .Z(n5788) );
  NAND U5659 ( .A(n5674), .B(n5672), .Z(n5791) );
  XOR U5660 ( .A(n5792), .B(n5793), .Z(n5672) );
  XNOR U5661 ( .A(n5794), .B(n5795), .Z(n5793) );
  IV U5662 ( .A(n5790), .Z(n5674) );
  NOR U5663 ( .A(n2924), .B(n2947), .Z(n5790) );
  AND U5664 ( .A(n5796), .B(n5797), .Z(n5675) );
  NANDN U5665 ( .A(n5680), .B(n5682), .Z(n5797) );
  NANDN U5666 ( .A(n5683), .B(n5798), .Z(n5796) );
  NANDN U5667 ( .A(n5682), .B(n5680), .Z(n5798) );
  XOR U5668 ( .A(n5799), .B(n5800), .Z(n5680) );
  XOR U5669 ( .A(n5801), .B(n5802), .Z(n5800) );
  AND U5670 ( .A(\stack[1][13] ), .B(\stack[0][13] ), .Z(n5682) );
  AND U5671 ( .A(n5803), .B(n5804), .Z(n5683) );
  NANDN U5672 ( .A(n5687), .B(n5805), .Z(n5804) );
  NANDN U5673 ( .A(n5690), .B(n5806), .Z(n5803) );
  NAND U5674 ( .A(n5689), .B(n5687), .Z(n5806) );
  XOR U5675 ( .A(n5807), .B(n5808), .Z(n5687) );
  XNOR U5676 ( .A(n5809), .B(n5810), .Z(n5808) );
  IV U5677 ( .A(n5805), .Z(n5689) );
  NOR U5678 ( .A(n2924), .B(n2899), .Z(n5805) );
  AND U5679 ( .A(n5811), .B(n5812), .Z(n5690) );
  NANDN U5680 ( .A(n5695), .B(n5697), .Z(n5812) );
  NANDN U5681 ( .A(n5698), .B(n5813), .Z(n5811) );
  NANDN U5682 ( .A(n5697), .B(n5695), .Z(n5813) );
  XOR U5683 ( .A(n5814), .B(n5815), .Z(n5695) );
  XOR U5684 ( .A(n5816), .B(n5817), .Z(n5815) );
  AND U5685 ( .A(\stack[1][13] ), .B(\stack[0][11] ), .Z(n5697) );
  AND U5686 ( .A(n5818), .B(n5819), .Z(n5698) );
  NANDN U5687 ( .A(n5702), .B(n5820), .Z(n5819) );
  NANDN U5688 ( .A(n5705), .B(n5821), .Z(n5818) );
  NAND U5689 ( .A(n5704), .B(n5702), .Z(n5821) );
  XOR U5690 ( .A(n5822), .B(n5823), .Z(n5702) );
  XNOR U5691 ( .A(n5824), .B(n5825), .Z(n5823) );
  IV U5692 ( .A(n5820), .Z(n5704) );
  NOR U5693 ( .A(n2924), .B(n2851), .Z(n5820) );
  AND U5694 ( .A(n5826), .B(n5827), .Z(n5705) );
  NANDN U5695 ( .A(n5710), .B(n5712), .Z(n5827) );
  NANDN U5696 ( .A(n5713), .B(n5828), .Z(n5826) );
  NANDN U5697 ( .A(n5712), .B(n5710), .Z(n5828) );
  XOR U5698 ( .A(n5829), .B(n5830), .Z(n5710) );
  XOR U5699 ( .A(n5831), .B(n5832), .Z(n5830) );
  AND U5700 ( .A(\stack[1][13] ), .B(\stack[0][9] ), .Z(n5712) );
  AND U5701 ( .A(n5833), .B(n5834), .Z(n5713) );
  NANDN U5702 ( .A(n5717), .B(n5835), .Z(n5834) );
  NANDN U5703 ( .A(n5720), .B(n5836), .Z(n5833) );
  NAND U5704 ( .A(n5719), .B(n5717), .Z(n5836) );
  XOR U5705 ( .A(n5837), .B(n5838), .Z(n5717) );
  XNOR U5706 ( .A(n5839), .B(n5840), .Z(n5838) );
  IV U5707 ( .A(n5835), .Z(n5719) );
  NOR U5708 ( .A(n2924), .B(n2803), .Z(n5835) );
  AND U5709 ( .A(n5841), .B(n5842), .Z(n5720) );
  NANDN U5710 ( .A(n5725), .B(n5727), .Z(n5842) );
  NANDN U5711 ( .A(n5728), .B(n5843), .Z(n5841) );
  NANDN U5712 ( .A(n5727), .B(n5725), .Z(n5843) );
  XOR U5713 ( .A(n5844), .B(n5845), .Z(n5725) );
  XOR U5714 ( .A(n5846), .B(n5847), .Z(n5845) );
  AND U5715 ( .A(\stack[1][13] ), .B(\stack[0][7] ), .Z(n5727) );
  AND U5716 ( .A(n5848), .B(n5849), .Z(n5728) );
  NANDN U5717 ( .A(n5732), .B(n5850), .Z(n5849) );
  NANDN U5718 ( .A(n5735), .B(n5851), .Z(n5848) );
  NAND U5719 ( .A(n5734), .B(n5732), .Z(n5851) );
  XOR U5720 ( .A(n5852), .B(n5853), .Z(n5732) );
  XNOR U5721 ( .A(n5854), .B(n5855), .Z(n5853) );
  IV U5722 ( .A(n5850), .Z(n5734) );
  NOR U5723 ( .A(n2924), .B(n2755), .Z(n5850) );
  AND U5724 ( .A(n5856), .B(n5857), .Z(n5735) );
  NANDN U5725 ( .A(n5740), .B(n5742), .Z(n5857) );
  NANDN U5726 ( .A(n5743), .B(n5858), .Z(n5856) );
  NANDN U5727 ( .A(n5742), .B(n5740), .Z(n5858) );
  XOR U5728 ( .A(n5859), .B(n5860), .Z(n5740) );
  XOR U5729 ( .A(n5861), .B(n5862), .Z(n5860) );
  AND U5730 ( .A(\stack[1][13] ), .B(\stack[0][5] ), .Z(n5742) );
  AND U5731 ( .A(n5863), .B(n5864), .Z(n5743) );
  NANDN U5732 ( .A(n5747), .B(n5865), .Z(n5864) );
  NANDN U5733 ( .A(n5750), .B(n5866), .Z(n5863) );
  NAND U5734 ( .A(n5749), .B(n5747), .Z(n5866) );
  XOR U5735 ( .A(n5867), .B(n5868), .Z(n5747) );
  XNOR U5736 ( .A(n5869), .B(n5870), .Z(n5868) );
  IV U5737 ( .A(n5865), .Z(n5749) );
  NOR U5738 ( .A(n2924), .B(n2707), .Z(n5865) );
  AND U5739 ( .A(n5871), .B(n5872), .Z(n5750) );
  NANDN U5740 ( .A(n5755), .B(n5757), .Z(n5872) );
  NANDN U5741 ( .A(n5758), .B(n5873), .Z(n5871) );
  NANDN U5742 ( .A(n5757), .B(n5755), .Z(n5873) );
  XNOR U5743 ( .A(n5874), .B(n5875), .Z(n5755) );
  XNOR U5744 ( .A(n5876), .B(n5877), .Z(n5875) );
  AND U5745 ( .A(\stack[1][13] ), .B(\stack[0][3] ), .Z(n5757) );
  AND U5746 ( .A(n5878), .B(n5879), .Z(n5758) );
  NANDN U5747 ( .A(n5762), .B(n5764), .Z(n5879) );
  NAND U5748 ( .A(n5880), .B(n5765), .Z(n5878) );
  ANDN U5749 ( .B(n5881), .A(n5770), .Z(n5765) );
  NAND U5750 ( .A(\stack[1][13] ), .B(\stack[0][1] ), .Z(n5770) );
  AND U5751 ( .A(\stack[0][0] ), .B(\stack[1][14] ), .Z(n5881) );
  NANDN U5752 ( .A(n5764), .B(n5762), .Z(n5880) );
  XNOR U5753 ( .A(n5882), .B(n5883), .Z(n5762) );
  NAND U5754 ( .A(\stack[0][0] ), .B(\stack[1][15] ), .Z(n5883) );
  AND U5755 ( .A(\stack[1][13] ), .B(\stack[0][2] ), .Z(n5764) );
  NOR U5756 ( .A(n2924), .B(n3019), .Z(n3569) );
  IV U5757 ( .A(\stack[0][17] ), .Z(n3019) );
  IV U5758 ( .A(\stack[1][13] ), .Z(n2924) );
  XNOR U5759 ( .A(n3577), .B(n5884), .Z(n3570) );
  XNOR U5760 ( .A(n3578), .B(n3579), .Z(n5884) );
  AND U5761 ( .A(n5885), .B(n5886), .Z(n3579) );
  NANDN U5762 ( .A(n5777), .B(n5779), .Z(n5886) );
  NANDN U5763 ( .A(n5780), .B(n5887), .Z(n5885) );
  NANDN U5764 ( .A(n5779), .B(n5777), .Z(n5887) );
  XOR U5765 ( .A(n5888), .B(n5889), .Z(n5777) );
  XOR U5766 ( .A(n5890), .B(n5891), .Z(n5889) );
  AND U5767 ( .A(\stack[1][14] ), .B(\stack[0][15] ), .Z(n5779) );
  AND U5768 ( .A(n5892), .B(n5893), .Z(n5780) );
  NANDN U5769 ( .A(n5784), .B(n5894), .Z(n5893) );
  NANDN U5770 ( .A(n5787), .B(n5895), .Z(n5892) );
  NAND U5771 ( .A(n5786), .B(n5784), .Z(n5895) );
  XOR U5772 ( .A(n5896), .B(n5897), .Z(n5784) );
  XNOR U5773 ( .A(n5898), .B(n5899), .Z(n5897) );
  IV U5774 ( .A(n5894), .Z(n5786) );
  NOR U5775 ( .A(n2948), .B(n2947), .Z(n5894) );
  AND U5776 ( .A(n5900), .B(n5901), .Z(n5787) );
  NANDN U5777 ( .A(n5792), .B(n5794), .Z(n5901) );
  NANDN U5778 ( .A(n5795), .B(n5902), .Z(n5900) );
  NANDN U5779 ( .A(n5794), .B(n5792), .Z(n5902) );
  XOR U5780 ( .A(n5903), .B(n5904), .Z(n5792) );
  XOR U5781 ( .A(n5905), .B(n5906), .Z(n5904) );
  AND U5782 ( .A(\stack[1][14] ), .B(\stack[0][13] ), .Z(n5794) );
  AND U5783 ( .A(n5907), .B(n5908), .Z(n5795) );
  NANDN U5784 ( .A(n5799), .B(n5909), .Z(n5908) );
  NANDN U5785 ( .A(n5802), .B(n5910), .Z(n5907) );
  NAND U5786 ( .A(n5801), .B(n5799), .Z(n5910) );
  XOR U5787 ( .A(n5911), .B(n5912), .Z(n5799) );
  XNOR U5788 ( .A(n5913), .B(n5914), .Z(n5912) );
  IV U5789 ( .A(n5909), .Z(n5801) );
  NOR U5790 ( .A(n2948), .B(n2899), .Z(n5909) );
  AND U5791 ( .A(n5915), .B(n5916), .Z(n5802) );
  NANDN U5792 ( .A(n5807), .B(n5809), .Z(n5916) );
  NANDN U5793 ( .A(n5810), .B(n5917), .Z(n5915) );
  NANDN U5794 ( .A(n5809), .B(n5807), .Z(n5917) );
  XOR U5795 ( .A(n5918), .B(n5919), .Z(n5807) );
  XOR U5796 ( .A(n5920), .B(n5921), .Z(n5919) );
  AND U5797 ( .A(\stack[1][14] ), .B(\stack[0][11] ), .Z(n5809) );
  AND U5798 ( .A(n5922), .B(n5923), .Z(n5810) );
  NANDN U5799 ( .A(n5814), .B(n5924), .Z(n5923) );
  NANDN U5800 ( .A(n5817), .B(n5925), .Z(n5922) );
  NAND U5801 ( .A(n5816), .B(n5814), .Z(n5925) );
  XOR U5802 ( .A(n5926), .B(n5927), .Z(n5814) );
  XNOR U5803 ( .A(n5928), .B(n5929), .Z(n5927) );
  IV U5804 ( .A(n5924), .Z(n5816) );
  NOR U5805 ( .A(n2948), .B(n2851), .Z(n5924) );
  AND U5806 ( .A(n5930), .B(n5931), .Z(n5817) );
  NANDN U5807 ( .A(n5822), .B(n5824), .Z(n5931) );
  NANDN U5808 ( .A(n5825), .B(n5932), .Z(n5930) );
  NANDN U5809 ( .A(n5824), .B(n5822), .Z(n5932) );
  XOR U5810 ( .A(n5933), .B(n5934), .Z(n5822) );
  XOR U5811 ( .A(n5935), .B(n5936), .Z(n5934) );
  AND U5812 ( .A(\stack[1][14] ), .B(\stack[0][9] ), .Z(n5824) );
  AND U5813 ( .A(n5937), .B(n5938), .Z(n5825) );
  NANDN U5814 ( .A(n5829), .B(n5939), .Z(n5938) );
  NANDN U5815 ( .A(n5832), .B(n5940), .Z(n5937) );
  NAND U5816 ( .A(n5831), .B(n5829), .Z(n5940) );
  XOR U5817 ( .A(n5941), .B(n5942), .Z(n5829) );
  XNOR U5818 ( .A(n5943), .B(n5944), .Z(n5942) );
  IV U5819 ( .A(n5939), .Z(n5831) );
  NOR U5820 ( .A(n2948), .B(n2803), .Z(n5939) );
  AND U5821 ( .A(n5945), .B(n5946), .Z(n5832) );
  NANDN U5822 ( .A(n5837), .B(n5839), .Z(n5946) );
  NANDN U5823 ( .A(n5840), .B(n5947), .Z(n5945) );
  NANDN U5824 ( .A(n5839), .B(n5837), .Z(n5947) );
  XOR U5825 ( .A(n5948), .B(n5949), .Z(n5837) );
  XOR U5826 ( .A(n5950), .B(n5951), .Z(n5949) );
  AND U5827 ( .A(\stack[1][14] ), .B(\stack[0][7] ), .Z(n5839) );
  AND U5828 ( .A(n5952), .B(n5953), .Z(n5840) );
  NANDN U5829 ( .A(n5844), .B(n5954), .Z(n5953) );
  NANDN U5830 ( .A(n5847), .B(n5955), .Z(n5952) );
  NAND U5831 ( .A(n5846), .B(n5844), .Z(n5955) );
  XOR U5832 ( .A(n5956), .B(n5957), .Z(n5844) );
  XNOR U5833 ( .A(n5958), .B(n5959), .Z(n5957) );
  IV U5834 ( .A(n5954), .Z(n5846) );
  NOR U5835 ( .A(n2948), .B(n2755), .Z(n5954) );
  AND U5836 ( .A(n5960), .B(n5961), .Z(n5847) );
  NANDN U5837 ( .A(n5852), .B(n5854), .Z(n5961) );
  NANDN U5838 ( .A(n5855), .B(n5962), .Z(n5960) );
  NANDN U5839 ( .A(n5854), .B(n5852), .Z(n5962) );
  XOR U5840 ( .A(n5963), .B(n5964), .Z(n5852) );
  XOR U5841 ( .A(n5965), .B(n5966), .Z(n5964) );
  AND U5842 ( .A(\stack[1][14] ), .B(\stack[0][5] ), .Z(n5854) );
  AND U5843 ( .A(n5967), .B(n5968), .Z(n5855) );
  NANDN U5844 ( .A(n5859), .B(n5969), .Z(n5968) );
  NANDN U5845 ( .A(n5862), .B(n5970), .Z(n5967) );
  NAND U5846 ( .A(n5861), .B(n5859), .Z(n5970) );
  XOR U5847 ( .A(n5971), .B(n5972), .Z(n5859) );
  XNOR U5848 ( .A(n5973), .B(n5974), .Z(n5972) );
  IV U5849 ( .A(n5969), .Z(n5861) );
  NOR U5850 ( .A(n2948), .B(n2707), .Z(n5969) );
  AND U5851 ( .A(n5975), .B(n5976), .Z(n5862) );
  NANDN U5852 ( .A(n5867), .B(n5869), .Z(n5976) );
  NANDN U5853 ( .A(n5870), .B(n5977), .Z(n5975) );
  NANDN U5854 ( .A(n5869), .B(n5867), .Z(n5977) );
  XNOR U5855 ( .A(n5978), .B(n5979), .Z(n5867) );
  XNOR U5856 ( .A(n5980), .B(n5981), .Z(n5979) );
  AND U5857 ( .A(\stack[1][14] ), .B(\stack[0][3] ), .Z(n5869) );
  AND U5858 ( .A(n5982), .B(n5983), .Z(n5870) );
  NANDN U5859 ( .A(n5874), .B(n5876), .Z(n5983) );
  NAND U5860 ( .A(n5984), .B(n5877), .Z(n5982) );
  ANDN U5861 ( .B(n5985), .A(n5882), .Z(n5877) );
  NAND U5862 ( .A(\stack[1][14] ), .B(\stack[0][1] ), .Z(n5882) );
  AND U5863 ( .A(\stack[0][0] ), .B(\stack[1][15] ), .Z(n5985) );
  NANDN U5864 ( .A(n5876), .B(n5874), .Z(n5984) );
  XNOR U5865 ( .A(n5986), .B(n5987), .Z(n5874) );
  NAND U5866 ( .A(\stack[0][0] ), .B(\stack[1][16] ), .Z(n5987) );
  AND U5867 ( .A(\stack[1][14] ), .B(\stack[0][2] ), .Z(n5876) );
  ANDN U5868 ( .B(\stack[0][16] ), .A(n2948), .Z(n3578) );
  IV U5869 ( .A(\stack[1][14] ), .Z(n2948) );
  XNOR U5870 ( .A(n3422), .B(n5988), .Z(n3577) );
  XNOR U5871 ( .A(n3421), .B(n3423), .Z(n5988) );
  AND U5872 ( .A(n5989), .B(n5990), .Z(n3423) );
  NANDN U5873 ( .A(n5888), .B(n5991), .Z(n5990) );
  NANDN U5874 ( .A(n5891), .B(n5992), .Z(n5989) );
  NAND U5875 ( .A(n5890), .B(n5888), .Z(n5992) );
  XOR U5876 ( .A(n5993), .B(n5994), .Z(n5888) );
  XNOR U5877 ( .A(n5995), .B(n5996), .Z(n5994) );
  IV U5878 ( .A(n5991), .Z(n5890) );
  NOR U5879 ( .A(n2972), .B(n2947), .Z(n5991) );
  IV U5880 ( .A(\stack[0][14] ), .Z(n2947) );
  AND U5881 ( .A(n5997), .B(n5998), .Z(n5891) );
  NANDN U5882 ( .A(n5896), .B(n5898), .Z(n5998) );
  NANDN U5883 ( .A(n5899), .B(n5999), .Z(n5997) );
  NANDN U5884 ( .A(n5898), .B(n5896), .Z(n5999) );
  XOR U5885 ( .A(n6000), .B(n6001), .Z(n5896) );
  XOR U5886 ( .A(n6002), .B(n6003), .Z(n6001) );
  AND U5887 ( .A(\stack[1][15] ), .B(\stack[0][13] ), .Z(n5898) );
  AND U5888 ( .A(n6004), .B(n6005), .Z(n5899) );
  NANDN U5889 ( .A(n5903), .B(n6006), .Z(n6005) );
  NANDN U5890 ( .A(n5906), .B(n6007), .Z(n6004) );
  NAND U5891 ( .A(n5905), .B(n5903), .Z(n6007) );
  XOR U5892 ( .A(n6008), .B(n6009), .Z(n5903) );
  XNOR U5893 ( .A(n6010), .B(n6011), .Z(n6009) );
  IV U5894 ( .A(n6006), .Z(n5905) );
  NOR U5895 ( .A(n2972), .B(n2899), .Z(n6006) );
  AND U5896 ( .A(n6012), .B(n6013), .Z(n5906) );
  NANDN U5897 ( .A(n5911), .B(n5913), .Z(n6013) );
  NANDN U5898 ( .A(n5914), .B(n6014), .Z(n6012) );
  NANDN U5899 ( .A(n5913), .B(n5911), .Z(n6014) );
  XOR U5900 ( .A(n6015), .B(n6016), .Z(n5911) );
  XOR U5901 ( .A(n6017), .B(n6018), .Z(n6016) );
  AND U5902 ( .A(\stack[1][15] ), .B(\stack[0][11] ), .Z(n5913) );
  AND U5903 ( .A(n6019), .B(n6020), .Z(n5914) );
  NANDN U5904 ( .A(n5918), .B(n6021), .Z(n6020) );
  NANDN U5905 ( .A(n5921), .B(n6022), .Z(n6019) );
  NAND U5906 ( .A(n5920), .B(n5918), .Z(n6022) );
  XOR U5907 ( .A(n6023), .B(n6024), .Z(n5918) );
  XNOR U5908 ( .A(n6025), .B(n6026), .Z(n6024) );
  IV U5909 ( .A(n6021), .Z(n5920) );
  NOR U5910 ( .A(n2972), .B(n2851), .Z(n6021) );
  AND U5911 ( .A(n6027), .B(n6028), .Z(n5921) );
  NANDN U5912 ( .A(n5926), .B(n5928), .Z(n6028) );
  NANDN U5913 ( .A(n5929), .B(n6029), .Z(n6027) );
  NANDN U5914 ( .A(n5928), .B(n5926), .Z(n6029) );
  XOR U5915 ( .A(n6030), .B(n6031), .Z(n5926) );
  XOR U5916 ( .A(n6032), .B(n6033), .Z(n6031) );
  AND U5917 ( .A(\stack[1][15] ), .B(\stack[0][9] ), .Z(n5928) );
  AND U5918 ( .A(n6034), .B(n6035), .Z(n5929) );
  NANDN U5919 ( .A(n5933), .B(n6036), .Z(n6035) );
  NANDN U5920 ( .A(n5936), .B(n6037), .Z(n6034) );
  NAND U5921 ( .A(n5935), .B(n5933), .Z(n6037) );
  XOR U5922 ( .A(n6038), .B(n6039), .Z(n5933) );
  XNOR U5923 ( .A(n6040), .B(n6041), .Z(n6039) );
  IV U5924 ( .A(n6036), .Z(n5935) );
  NOR U5925 ( .A(n2972), .B(n2803), .Z(n6036) );
  AND U5926 ( .A(n6042), .B(n6043), .Z(n5936) );
  NANDN U5927 ( .A(n5941), .B(n5943), .Z(n6043) );
  NANDN U5928 ( .A(n5944), .B(n6044), .Z(n6042) );
  NANDN U5929 ( .A(n5943), .B(n5941), .Z(n6044) );
  XOR U5930 ( .A(n6045), .B(n6046), .Z(n5941) );
  XOR U5931 ( .A(n6047), .B(n6048), .Z(n6046) );
  AND U5932 ( .A(\stack[1][15] ), .B(\stack[0][7] ), .Z(n5943) );
  AND U5933 ( .A(n6049), .B(n6050), .Z(n5944) );
  NANDN U5934 ( .A(n5948), .B(n6051), .Z(n6050) );
  NANDN U5935 ( .A(n5951), .B(n6052), .Z(n6049) );
  NAND U5936 ( .A(n5950), .B(n5948), .Z(n6052) );
  XOR U5937 ( .A(n6053), .B(n6054), .Z(n5948) );
  XNOR U5938 ( .A(n6055), .B(n6056), .Z(n6054) );
  IV U5939 ( .A(n6051), .Z(n5950) );
  NOR U5940 ( .A(n2972), .B(n2755), .Z(n6051) );
  AND U5941 ( .A(n6057), .B(n6058), .Z(n5951) );
  NANDN U5942 ( .A(n5956), .B(n5958), .Z(n6058) );
  NANDN U5943 ( .A(n5959), .B(n6059), .Z(n6057) );
  NANDN U5944 ( .A(n5958), .B(n5956), .Z(n6059) );
  XOR U5945 ( .A(n6060), .B(n6061), .Z(n5956) );
  XOR U5946 ( .A(n6062), .B(n6063), .Z(n6061) );
  AND U5947 ( .A(\stack[1][15] ), .B(\stack[0][5] ), .Z(n5958) );
  AND U5948 ( .A(n6064), .B(n6065), .Z(n5959) );
  NANDN U5949 ( .A(n5963), .B(n6066), .Z(n6065) );
  NANDN U5950 ( .A(n5966), .B(n6067), .Z(n6064) );
  NAND U5951 ( .A(n5965), .B(n5963), .Z(n6067) );
  XOR U5952 ( .A(n6068), .B(n6069), .Z(n5963) );
  XNOR U5953 ( .A(n6070), .B(n6071), .Z(n6069) );
  IV U5954 ( .A(n6066), .Z(n5965) );
  NOR U5955 ( .A(n2972), .B(n2707), .Z(n6066) );
  AND U5956 ( .A(n6072), .B(n6073), .Z(n5966) );
  NANDN U5957 ( .A(n5971), .B(n5973), .Z(n6073) );
  NANDN U5958 ( .A(n5974), .B(n6074), .Z(n6072) );
  NANDN U5959 ( .A(n5973), .B(n5971), .Z(n6074) );
  XNOR U5960 ( .A(n6075), .B(n6076), .Z(n5971) );
  XNOR U5961 ( .A(n6077), .B(n6078), .Z(n6076) );
  AND U5962 ( .A(\stack[1][15] ), .B(\stack[0][3] ), .Z(n5973) );
  AND U5963 ( .A(n6079), .B(n6080), .Z(n5974) );
  NANDN U5964 ( .A(n5978), .B(n5980), .Z(n6080) );
  NAND U5965 ( .A(n6081), .B(n5981), .Z(n6079) );
  ANDN U5966 ( .B(n6082), .A(n5986), .Z(n5981) );
  NAND U5967 ( .A(\stack[1][15] ), .B(\stack[0][1] ), .Z(n5986) );
  AND U5968 ( .A(\stack[0][0] ), .B(\stack[1][16] ), .Z(n6082) );
  NANDN U5969 ( .A(n5980), .B(n5978), .Z(n6081) );
  XNOR U5970 ( .A(n6083), .B(n6084), .Z(n5978) );
  NAND U5971 ( .A(\stack[0][0] ), .B(\stack[1][17] ), .Z(n6084) );
  AND U5972 ( .A(\stack[1][15] ), .B(\stack[0][2] ), .Z(n5980) );
  NOR U5973 ( .A(n2972), .B(n2971), .Z(n3421) );
  IV U5974 ( .A(\stack[0][15] ), .Z(n2971) );
  IV U5975 ( .A(\stack[1][15] ), .Z(n2972) );
  XNOR U5976 ( .A(n3533), .B(n6085), .Z(n3422) );
  XNOR U5977 ( .A(n3534), .B(n3535), .Z(n6085) );
  AND U5978 ( .A(n6086), .B(n6087), .Z(n3535) );
  NANDN U5979 ( .A(n5993), .B(n5995), .Z(n6087) );
  NANDN U5980 ( .A(n5996), .B(n6088), .Z(n6086) );
  NANDN U5981 ( .A(n5995), .B(n5993), .Z(n6088) );
  XOR U5982 ( .A(n6089), .B(n6090), .Z(n5993) );
  XOR U5983 ( .A(n6091), .B(n6092), .Z(n6090) );
  AND U5984 ( .A(\stack[1][16] ), .B(\stack[0][13] ), .Z(n5995) );
  AND U5985 ( .A(n6093), .B(n6094), .Z(n5996) );
  NANDN U5986 ( .A(n6000), .B(n6095), .Z(n6094) );
  NANDN U5987 ( .A(n6003), .B(n6096), .Z(n6093) );
  NAND U5988 ( .A(n6002), .B(n6000), .Z(n6096) );
  XOR U5989 ( .A(n6097), .B(n6098), .Z(n6000) );
  XNOR U5990 ( .A(n6099), .B(n6100), .Z(n6098) );
  IV U5991 ( .A(n6095), .Z(n6002) );
  NOR U5992 ( .A(n2996), .B(n2899), .Z(n6095) );
  AND U5993 ( .A(n6101), .B(n6102), .Z(n6003) );
  NANDN U5994 ( .A(n6008), .B(n6010), .Z(n6102) );
  NANDN U5995 ( .A(n6011), .B(n6103), .Z(n6101) );
  NANDN U5996 ( .A(n6010), .B(n6008), .Z(n6103) );
  XOR U5997 ( .A(n6104), .B(n6105), .Z(n6008) );
  XOR U5998 ( .A(n6106), .B(n6107), .Z(n6105) );
  AND U5999 ( .A(\stack[1][16] ), .B(\stack[0][11] ), .Z(n6010) );
  AND U6000 ( .A(n6108), .B(n6109), .Z(n6011) );
  NANDN U6001 ( .A(n6015), .B(n6110), .Z(n6109) );
  NANDN U6002 ( .A(n6018), .B(n6111), .Z(n6108) );
  NAND U6003 ( .A(n6017), .B(n6015), .Z(n6111) );
  XOR U6004 ( .A(n6112), .B(n6113), .Z(n6015) );
  XNOR U6005 ( .A(n6114), .B(n6115), .Z(n6113) );
  IV U6006 ( .A(n6110), .Z(n6017) );
  NOR U6007 ( .A(n2996), .B(n2851), .Z(n6110) );
  AND U6008 ( .A(n6116), .B(n6117), .Z(n6018) );
  NANDN U6009 ( .A(n6023), .B(n6025), .Z(n6117) );
  NANDN U6010 ( .A(n6026), .B(n6118), .Z(n6116) );
  NANDN U6011 ( .A(n6025), .B(n6023), .Z(n6118) );
  XOR U6012 ( .A(n6119), .B(n6120), .Z(n6023) );
  XOR U6013 ( .A(n6121), .B(n6122), .Z(n6120) );
  AND U6014 ( .A(\stack[1][16] ), .B(\stack[0][9] ), .Z(n6025) );
  AND U6015 ( .A(n6123), .B(n6124), .Z(n6026) );
  NANDN U6016 ( .A(n6030), .B(n6125), .Z(n6124) );
  NANDN U6017 ( .A(n6033), .B(n6126), .Z(n6123) );
  NAND U6018 ( .A(n6032), .B(n6030), .Z(n6126) );
  XOR U6019 ( .A(n6127), .B(n6128), .Z(n6030) );
  XNOR U6020 ( .A(n6129), .B(n6130), .Z(n6128) );
  IV U6021 ( .A(n6125), .Z(n6032) );
  NOR U6022 ( .A(n2996), .B(n2803), .Z(n6125) );
  AND U6023 ( .A(n6131), .B(n6132), .Z(n6033) );
  NANDN U6024 ( .A(n6038), .B(n6040), .Z(n6132) );
  NANDN U6025 ( .A(n6041), .B(n6133), .Z(n6131) );
  NANDN U6026 ( .A(n6040), .B(n6038), .Z(n6133) );
  XOR U6027 ( .A(n6134), .B(n6135), .Z(n6038) );
  XOR U6028 ( .A(n6136), .B(n6137), .Z(n6135) );
  AND U6029 ( .A(\stack[1][16] ), .B(\stack[0][7] ), .Z(n6040) );
  AND U6030 ( .A(n6138), .B(n6139), .Z(n6041) );
  NANDN U6031 ( .A(n6045), .B(n6140), .Z(n6139) );
  NANDN U6032 ( .A(n6048), .B(n6141), .Z(n6138) );
  NAND U6033 ( .A(n6047), .B(n6045), .Z(n6141) );
  XOR U6034 ( .A(n6142), .B(n6143), .Z(n6045) );
  XNOR U6035 ( .A(n6144), .B(n6145), .Z(n6143) );
  IV U6036 ( .A(n6140), .Z(n6047) );
  NOR U6037 ( .A(n2996), .B(n2755), .Z(n6140) );
  AND U6038 ( .A(n6146), .B(n6147), .Z(n6048) );
  NANDN U6039 ( .A(n6053), .B(n6055), .Z(n6147) );
  NANDN U6040 ( .A(n6056), .B(n6148), .Z(n6146) );
  NANDN U6041 ( .A(n6055), .B(n6053), .Z(n6148) );
  XOR U6042 ( .A(n6149), .B(n6150), .Z(n6053) );
  XOR U6043 ( .A(n6151), .B(n6152), .Z(n6150) );
  AND U6044 ( .A(\stack[1][16] ), .B(\stack[0][5] ), .Z(n6055) );
  AND U6045 ( .A(n6153), .B(n6154), .Z(n6056) );
  NANDN U6046 ( .A(n6060), .B(n6155), .Z(n6154) );
  NANDN U6047 ( .A(n6063), .B(n6156), .Z(n6153) );
  NAND U6048 ( .A(n6062), .B(n6060), .Z(n6156) );
  XOR U6049 ( .A(n6157), .B(n6158), .Z(n6060) );
  XNOR U6050 ( .A(n6159), .B(n6160), .Z(n6158) );
  IV U6051 ( .A(n6155), .Z(n6062) );
  NOR U6052 ( .A(n2996), .B(n2707), .Z(n6155) );
  AND U6053 ( .A(n6161), .B(n6162), .Z(n6063) );
  NANDN U6054 ( .A(n6068), .B(n6070), .Z(n6162) );
  NANDN U6055 ( .A(n6071), .B(n6163), .Z(n6161) );
  NANDN U6056 ( .A(n6070), .B(n6068), .Z(n6163) );
  XNOR U6057 ( .A(n6164), .B(n6165), .Z(n6068) );
  XNOR U6058 ( .A(n6166), .B(n6167), .Z(n6165) );
  AND U6059 ( .A(\stack[1][16] ), .B(\stack[0][3] ), .Z(n6070) );
  AND U6060 ( .A(n6168), .B(n6169), .Z(n6071) );
  NANDN U6061 ( .A(n6075), .B(n6077), .Z(n6169) );
  NAND U6062 ( .A(n6170), .B(n6078), .Z(n6168) );
  ANDN U6063 ( .B(n6171), .A(n6083), .Z(n6078) );
  NAND U6064 ( .A(\stack[1][16] ), .B(\stack[0][1] ), .Z(n6083) );
  AND U6065 ( .A(\stack[0][0] ), .B(\stack[1][17] ), .Z(n6171) );
  NANDN U6066 ( .A(n6077), .B(n6075), .Z(n6170) );
  XNOR U6067 ( .A(n6172), .B(n6173), .Z(n6075) );
  NAND U6068 ( .A(\stack[0][0] ), .B(\stack[1][18] ), .Z(n6173) );
  AND U6069 ( .A(\stack[1][16] ), .B(\stack[0][2] ), .Z(n6077) );
  ANDN U6070 ( .B(\stack[0][14] ), .A(n2996), .Z(n3534) );
  IV U6071 ( .A(\stack[1][16] ), .Z(n2996) );
  XNOR U6072 ( .A(n3544), .B(n6174), .Z(n3533) );
  XNOR U6073 ( .A(n3543), .B(n3545), .Z(n6174) );
  AND U6074 ( .A(n6175), .B(n6176), .Z(n3545) );
  NANDN U6075 ( .A(n6089), .B(n6177), .Z(n6176) );
  NANDN U6076 ( .A(n6092), .B(n6178), .Z(n6175) );
  NAND U6077 ( .A(n6091), .B(n6089), .Z(n6178) );
  XOR U6078 ( .A(n6179), .B(n6180), .Z(n6089) );
  XNOR U6079 ( .A(n6181), .B(n6182), .Z(n6180) );
  IV U6080 ( .A(n6177), .Z(n6091) );
  NOR U6081 ( .A(n3020), .B(n2899), .Z(n6177) );
  IV U6082 ( .A(\stack[0][12] ), .Z(n2899) );
  AND U6083 ( .A(n6183), .B(n6184), .Z(n6092) );
  NANDN U6084 ( .A(n6097), .B(n6099), .Z(n6184) );
  NANDN U6085 ( .A(n6100), .B(n6185), .Z(n6183) );
  NANDN U6086 ( .A(n6099), .B(n6097), .Z(n6185) );
  XOR U6087 ( .A(n6186), .B(n6187), .Z(n6097) );
  XOR U6088 ( .A(n6188), .B(n6189), .Z(n6187) );
  AND U6089 ( .A(\stack[1][17] ), .B(\stack[0][11] ), .Z(n6099) );
  AND U6090 ( .A(n6190), .B(n6191), .Z(n6100) );
  NANDN U6091 ( .A(n6104), .B(n6192), .Z(n6191) );
  NANDN U6092 ( .A(n6107), .B(n6193), .Z(n6190) );
  NAND U6093 ( .A(n6106), .B(n6104), .Z(n6193) );
  XOR U6094 ( .A(n6194), .B(n6195), .Z(n6104) );
  XNOR U6095 ( .A(n6196), .B(n6197), .Z(n6195) );
  IV U6096 ( .A(n6192), .Z(n6106) );
  NOR U6097 ( .A(n3020), .B(n2851), .Z(n6192) );
  AND U6098 ( .A(n6198), .B(n6199), .Z(n6107) );
  NANDN U6099 ( .A(n6112), .B(n6114), .Z(n6199) );
  NANDN U6100 ( .A(n6115), .B(n6200), .Z(n6198) );
  NANDN U6101 ( .A(n6114), .B(n6112), .Z(n6200) );
  XOR U6102 ( .A(n6201), .B(n6202), .Z(n6112) );
  XOR U6103 ( .A(n6203), .B(n6204), .Z(n6202) );
  AND U6104 ( .A(\stack[1][17] ), .B(\stack[0][9] ), .Z(n6114) );
  AND U6105 ( .A(n6205), .B(n6206), .Z(n6115) );
  NANDN U6106 ( .A(n6119), .B(n6207), .Z(n6206) );
  NANDN U6107 ( .A(n6122), .B(n6208), .Z(n6205) );
  NAND U6108 ( .A(n6121), .B(n6119), .Z(n6208) );
  XOR U6109 ( .A(n6209), .B(n6210), .Z(n6119) );
  XNOR U6110 ( .A(n6211), .B(n6212), .Z(n6210) );
  IV U6111 ( .A(n6207), .Z(n6121) );
  NOR U6112 ( .A(n3020), .B(n2803), .Z(n6207) );
  AND U6113 ( .A(n6213), .B(n6214), .Z(n6122) );
  NANDN U6114 ( .A(n6127), .B(n6129), .Z(n6214) );
  NANDN U6115 ( .A(n6130), .B(n6215), .Z(n6213) );
  NANDN U6116 ( .A(n6129), .B(n6127), .Z(n6215) );
  XOR U6117 ( .A(n6216), .B(n6217), .Z(n6127) );
  XOR U6118 ( .A(n6218), .B(n6219), .Z(n6217) );
  AND U6119 ( .A(\stack[1][17] ), .B(\stack[0][7] ), .Z(n6129) );
  AND U6120 ( .A(n6220), .B(n6221), .Z(n6130) );
  NANDN U6121 ( .A(n6134), .B(n6222), .Z(n6221) );
  NANDN U6122 ( .A(n6137), .B(n6223), .Z(n6220) );
  NAND U6123 ( .A(n6136), .B(n6134), .Z(n6223) );
  XOR U6124 ( .A(n6224), .B(n6225), .Z(n6134) );
  XNOR U6125 ( .A(n6226), .B(n6227), .Z(n6225) );
  IV U6126 ( .A(n6222), .Z(n6136) );
  NOR U6127 ( .A(n3020), .B(n2755), .Z(n6222) );
  AND U6128 ( .A(n6228), .B(n6229), .Z(n6137) );
  NANDN U6129 ( .A(n6142), .B(n6144), .Z(n6229) );
  NANDN U6130 ( .A(n6145), .B(n6230), .Z(n6228) );
  NANDN U6131 ( .A(n6144), .B(n6142), .Z(n6230) );
  XOR U6132 ( .A(n6231), .B(n6232), .Z(n6142) );
  XOR U6133 ( .A(n6233), .B(n6234), .Z(n6232) );
  AND U6134 ( .A(\stack[1][17] ), .B(\stack[0][5] ), .Z(n6144) );
  AND U6135 ( .A(n6235), .B(n6236), .Z(n6145) );
  NANDN U6136 ( .A(n6149), .B(n6237), .Z(n6236) );
  NANDN U6137 ( .A(n6152), .B(n6238), .Z(n6235) );
  NAND U6138 ( .A(n6151), .B(n6149), .Z(n6238) );
  XOR U6139 ( .A(n6239), .B(n6240), .Z(n6149) );
  XNOR U6140 ( .A(n6241), .B(n6242), .Z(n6240) );
  IV U6141 ( .A(n6237), .Z(n6151) );
  NOR U6142 ( .A(n3020), .B(n2707), .Z(n6237) );
  AND U6143 ( .A(n6243), .B(n6244), .Z(n6152) );
  NANDN U6144 ( .A(n6157), .B(n6159), .Z(n6244) );
  NANDN U6145 ( .A(n6160), .B(n6245), .Z(n6243) );
  NANDN U6146 ( .A(n6159), .B(n6157), .Z(n6245) );
  XNOR U6147 ( .A(n6246), .B(n6247), .Z(n6157) );
  XNOR U6148 ( .A(n6248), .B(n6249), .Z(n6247) );
  AND U6149 ( .A(\stack[1][17] ), .B(\stack[0][3] ), .Z(n6159) );
  AND U6150 ( .A(n6250), .B(n6251), .Z(n6160) );
  NANDN U6151 ( .A(n6164), .B(n6166), .Z(n6251) );
  NAND U6152 ( .A(n6252), .B(n6167), .Z(n6250) );
  ANDN U6153 ( .B(n6253), .A(n6172), .Z(n6167) );
  NAND U6154 ( .A(\stack[1][17] ), .B(\stack[0][1] ), .Z(n6172) );
  AND U6155 ( .A(\stack[0][0] ), .B(\stack[1][18] ), .Z(n6253) );
  NANDN U6156 ( .A(n6166), .B(n6164), .Z(n6252) );
  XNOR U6157 ( .A(n6254), .B(n6255), .Z(n6164) );
  NAND U6158 ( .A(\stack[0][0] ), .B(\stack[1][19] ), .Z(n6255) );
  AND U6159 ( .A(\stack[1][17] ), .B(\stack[0][2] ), .Z(n6166) );
  NOR U6160 ( .A(n3020), .B(n2923), .Z(n3543) );
  IV U6161 ( .A(\stack[0][13] ), .Z(n2923) );
  IV U6162 ( .A(\stack[1][17] ), .Z(n3020) );
  XNOR U6163 ( .A(n3551), .B(n6256), .Z(n3544) );
  XNOR U6164 ( .A(n3552), .B(n3553), .Z(n6256) );
  AND U6165 ( .A(n6257), .B(n6258), .Z(n3553) );
  NANDN U6166 ( .A(n6179), .B(n6181), .Z(n6258) );
  NANDN U6167 ( .A(n6182), .B(n6259), .Z(n6257) );
  NANDN U6168 ( .A(n6181), .B(n6179), .Z(n6259) );
  XOR U6169 ( .A(n6260), .B(n6261), .Z(n6179) );
  XOR U6170 ( .A(n6262), .B(n6263), .Z(n6261) );
  AND U6171 ( .A(\stack[1][18] ), .B(\stack[0][11] ), .Z(n6181) );
  AND U6172 ( .A(n6264), .B(n6265), .Z(n6182) );
  NANDN U6173 ( .A(n6186), .B(n6266), .Z(n6265) );
  NANDN U6174 ( .A(n6189), .B(n6267), .Z(n6264) );
  NAND U6175 ( .A(n6188), .B(n6186), .Z(n6267) );
  XOR U6176 ( .A(n6268), .B(n6269), .Z(n6186) );
  XNOR U6177 ( .A(n6270), .B(n6271), .Z(n6269) );
  IV U6178 ( .A(n6266), .Z(n6188) );
  NOR U6179 ( .A(n3044), .B(n2851), .Z(n6266) );
  AND U6180 ( .A(n6272), .B(n6273), .Z(n6189) );
  NANDN U6181 ( .A(n6194), .B(n6196), .Z(n6273) );
  NANDN U6182 ( .A(n6197), .B(n6274), .Z(n6272) );
  NANDN U6183 ( .A(n6196), .B(n6194), .Z(n6274) );
  XOR U6184 ( .A(n6275), .B(n6276), .Z(n6194) );
  XOR U6185 ( .A(n6277), .B(n6278), .Z(n6276) );
  AND U6186 ( .A(\stack[1][18] ), .B(\stack[0][9] ), .Z(n6196) );
  AND U6187 ( .A(n6279), .B(n6280), .Z(n6197) );
  NANDN U6188 ( .A(n6201), .B(n6281), .Z(n6280) );
  NANDN U6189 ( .A(n6204), .B(n6282), .Z(n6279) );
  NAND U6190 ( .A(n6203), .B(n6201), .Z(n6282) );
  XOR U6191 ( .A(n6283), .B(n6284), .Z(n6201) );
  XNOR U6192 ( .A(n6285), .B(n6286), .Z(n6284) );
  IV U6193 ( .A(n6281), .Z(n6203) );
  NOR U6194 ( .A(n3044), .B(n2803), .Z(n6281) );
  AND U6195 ( .A(n6287), .B(n6288), .Z(n6204) );
  NANDN U6196 ( .A(n6209), .B(n6211), .Z(n6288) );
  NANDN U6197 ( .A(n6212), .B(n6289), .Z(n6287) );
  NANDN U6198 ( .A(n6211), .B(n6209), .Z(n6289) );
  XOR U6199 ( .A(n6290), .B(n6291), .Z(n6209) );
  XOR U6200 ( .A(n6292), .B(n6293), .Z(n6291) );
  AND U6201 ( .A(\stack[1][18] ), .B(\stack[0][7] ), .Z(n6211) );
  AND U6202 ( .A(n6294), .B(n6295), .Z(n6212) );
  NANDN U6203 ( .A(n6216), .B(n6296), .Z(n6295) );
  NANDN U6204 ( .A(n6219), .B(n6297), .Z(n6294) );
  NAND U6205 ( .A(n6218), .B(n6216), .Z(n6297) );
  XOR U6206 ( .A(n6298), .B(n6299), .Z(n6216) );
  XNOR U6207 ( .A(n6300), .B(n6301), .Z(n6299) );
  IV U6208 ( .A(n6296), .Z(n6218) );
  NOR U6209 ( .A(n3044), .B(n2755), .Z(n6296) );
  AND U6210 ( .A(n6302), .B(n6303), .Z(n6219) );
  NANDN U6211 ( .A(n6224), .B(n6226), .Z(n6303) );
  NANDN U6212 ( .A(n6227), .B(n6304), .Z(n6302) );
  NANDN U6213 ( .A(n6226), .B(n6224), .Z(n6304) );
  XOR U6214 ( .A(n6305), .B(n6306), .Z(n6224) );
  XOR U6215 ( .A(n6307), .B(n6308), .Z(n6306) );
  AND U6216 ( .A(\stack[1][18] ), .B(\stack[0][5] ), .Z(n6226) );
  AND U6217 ( .A(n6309), .B(n6310), .Z(n6227) );
  NANDN U6218 ( .A(n6231), .B(n6311), .Z(n6310) );
  NANDN U6219 ( .A(n6234), .B(n6312), .Z(n6309) );
  NAND U6220 ( .A(n6233), .B(n6231), .Z(n6312) );
  XOR U6221 ( .A(n6313), .B(n6314), .Z(n6231) );
  XNOR U6222 ( .A(n6315), .B(n6316), .Z(n6314) );
  IV U6223 ( .A(n6311), .Z(n6233) );
  NOR U6224 ( .A(n3044), .B(n2707), .Z(n6311) );
  AND U6225 ( .A(n6317), .B(n6318), .Z(n6234) );
  NANDN U6226 ( .A(n6239), .B(n6241), .Z(n6318) );
  NANDN U6227 ( .A(n6242), .B(n6319), .Z(n6317) );
  NANDN U6228 ( .A(n6241), .B(n6239), .Z(n6319) );
  XNOR U6229 ( .A(n6320), .B(n6321), .Z(n6239) );
  XNOR U6230 ( .A(n6322), .B(n6323), .Z(n6321) );
  AND U6231 ( .A(\stack[1][18] ), .B(\stack[0][3] ), .Z(n6241) );
  AND U6232 ( .A(n6324), .B(n6325), .Z(n6242) );
  NANDN U6233 ( .A(n6246), .B(n6248), .Z(n6325) );
  NAND U6234 ( .A(n6326), .B(n6249), .Z(n6324) );
  ANDN U6235 ( .B(n6327), .A(n6254), .Z(n6249) );
  NAND U6236 ( .A(\stack[1][18] ), .B(\stack[0][1] ), .Z(n6254) );
  AND U6237 ( .A(\stack[0][0] ), .B(\stack[1][19] ), .Z(n6327) );
  NANDN U6238 ( .A(n6248), .B(n6246), .Z(n6326) );
  XNOR U6239 ( .A(n6328), .B(n6329), .Z(n6246) );
  NAND U6240 ( .A(\stack[0][0] ), .B(\stack[1][20] ), .Z(n6329) );
  AND U6241 ( .A(\stack[1][18] ), .B(\stack[0][2] ), .Z(n6248) );
  ANDN U6242 ( .B(\stack[0][12] ), .A(n3044), .Z(n3552) );
  IV U6243 ( .A(\stack[1][18] ), .Z(n3044) );
  XNOR U6244 ( .A(n3434), .B(n6330), .Z(n3551) );
  XNOR U6245 ( .A(n3433), .B(n3435), .Z(n6330) );
  AND U6246 ( .A(n6331), .B(n6332), .Z(n3435) );
  NANDN U6247 ( .A(n6260), .B(n6333), .Z(n6332) );
  NANDN U6248 ( .A(n6263), .B(n6334), .Z(n6331) );
  NAND U6249 ( .A(n6262), .B(n6260), .Z(n6334) );
  XOR U6250 ( .A(n6335), .B(n6336), .Z(n6260) );
  XNOR U6251 ( .A(n6337), .B(n6338), .Z(n6336) );
  IV U6252 ( .A(n6333), .Z(n6262) );
  NOR U6253 ( .A(n3068), .B(n2851), .Z(n6333) );
  IV U6254 ( .A(\stack[0][10] ), .Z(n2851) );
  AND U6255 ( .A(n6339), .B(n6340), .Z(n6263) );
  NANDN U6256 ( .A(n6268), .B(n6270), .Z(n6340) );
  NANDN U6257 ( .A(n6271), .B(n6341), .Z(n6339) );
  NANDN U6258 ( .A(n6270), .B(n6268), .Z(n6341) );
  XOR U6259 ( .A(n6342), .B(n6343), .Z(n6268) );
  XOR U6260 ( .A(n6344), .B(n6345), .Z(n6343) );
  AND U6261 ( .A(\stack[1][19] ), .B(\stack[0][9] ), .Z(n6270) );
  AND U6262 ( .A(n6346), .B(n6347), .Z(n6271) );
  NANDN U6263 ( .A(n6275), .B(n6348), .Z(n6347) );
  NANDN U6264 ( .A(n6278), .B(n6349), .Z(n6346) );
  NAND U6265 ( .A(n6277), .B(n6275), .Z(n6349) );
  XOR U6266 ( .A(n6350), .B(n6351), .Z(n6275) );
  XNOR U6267 ( .A(n6352), .B(n6353), .Z(n6351) );
  IV U6268 ( .A(n6348), .Z(n6277) );
  NOR U6269 ( .A(n3068), .B(n2803), .Z(n6348) );
  AND U6270 ( .A(n6354), .B(n6355), .Z(n6278) );
  NANDN U6271 ( .A(n6283), .B(n6285), .Z(n6355) );
  NANDN U6272 ( .A(n6286), .B(n6356), .Z(n6354) );
  NANDN U6273 ( .A(n6285), .B(n6283), .Z(n6356) );
  XOR U6274 ( .A(n6357), .B(n6358), .Z(n6283) );
  XOR U6275 ( .A(n6359), .B(n6360), .Z(n6358) );
  AND U6276 ( .A(\stack[1][19] ), .B(\stack[0][7] ), .Z(n6285) );
  AND U6277 ( .A(n6361), .B(n6362), .Z(n6286) );
  NANDN U6278 ( .A(n6290), .B(n6363), .Z(n6362) );
  NANDN U6279 ( .A(n6293), .B(n6364), .Z(n6361) );
  NAND U6280 ( .A(n6292), .B(n6290), .Z(n6364) );
  XOR U6281 ( .A(n6365), .B(n6366), .Z(n6290) );
  XNOR U6282 ( .A(n6367), .B(n6368), .Z(n6366) );
  IV U6283 ( .A(n6363), .Z(n6292) );
  NOR U6284 ( .A(n3068), .B(n2755), .Z(n6363) );
  AND U6285 ( .A(n6369), .B(n6370), .Z(n6293) );
  NANDN U6286 ( .A(n6298), .B(n6300), .Z(n6370) );
  NANDN U6287 ( .A(n6301), .B(n6371), .Z(n6369) );
  NANDN U6288 ( .A(n6300), .B(n6298), .Z(n6371) );
  XOR U6289 ( .A(n6372), .B(n6373), .Z(n6298) );
  XOR U6290 ( .A(n6374), .B(n6375), .Z(n6373) );
  AND U6291 ( .A(\stack[1][19] ), .B(\stack[0][5] ), .Z(n6300) );
  AND U6292 ( .A(n6376), .B(n6377), .Z(n6301) );
  NANDN U6293 ( .A(n6305), .B(n6378), .Z(n6377) );
  NANDN U6294 ( .A(n6308), .B(n6379), .Z(n6376) );
  NAND U6295 ( .A(n6307), .B(n6305), .Z(n6379) );
  XOR U6296 ( .A(n6380), .B(n6381), .Z(n6305) );
  XNOR U6297 ( .A(n6382), .B(n6383), .Z(n6381) );
  IV U6298 ( .A(n6378), .Z(n6307) );
  NOR U6299 ( .A(n3068), .B(n2707), .Z(n6378) );
  AND U6300 ( .A(n6384), .B(n6385), .Z(n6308) );
  NANDN U6301 ( .A(n6313), .B(n6315), .Z(n6385) );
  NANDN U6302 ( .A(n6316), .B(n6386), .Z(n6384) );
  NANDN U6303 ( .A(n6315), .B(n6313), .Z(n6386) );
  XNOR U6304 ( .A(n6387), .B(n6388), .Z(n6313) );
  XNOR U6305 ( .A(n6389), .B(n6390), .Z(n6388) );
  AND U6306 ( .A(\stack[1][19] ), .B(\stack[0][3] ), .Z(n6315) );
  AND U6307 ( .A(n6391), .B(n6392), .Z(n6316) );
  NANDN U6308 ( .A(n6320), .B(n6322), .Z(n6392) );
  NAND U6309 ( .A(n6393), .B(n6323), .Z(n6391) );
  ANDN U6310 ( .B(n6394), .A(n6328), .Z(n6323) );
  NAND U6311 ( .A(\stack[1][19] ), .B(\stack[0][1] ), .Z(n6328) );
  AND U6312 ( .A(\stack[0][0] ), .B(\stack[1][20] ), .Z(n6394) );
  NANDN U6313 ( .A(n6322), .B(n6320), .Z(n6393) );
  XNOR U6314 ( .A(n6395), .B(n6396), .Z(n6320) );
  NAND U6315 ( .A(\stack[0][0] ), .B(\stack[1][21] ), .Z(n6396) );
  AND U6316 ( .A(\stack[1][19] ), .B(\stack[0][2] ), .Z(n6322) );
  NOR U6317 ( .A(n3068), .B(n2875), .Z(n3433) );
  IV U6318 ( .A(\stack[0][11] ), .Z(n2875) );
  IV U6319 ( .A(\stack[1][19] ), .Z(n3068) );
  XNOR U6320 ( .A(n3507), .B(n6397), .Z(n3434) );
  XNOR U6321 ( .A(n3508), .B(n3509), .Z(n6397) );
  AND U6322 ( .A(n6398), .B(n6399), .Z(n3509) );
  NANDN U6323 ( .A(n6335), .B(n6337), .Z(n6399) );
  NANDN U6324 ( .A(n6338), .B(n6400), .Z(n6398) );
  NANDN U6325 ( .A(n6337), .B(n6335), .Z(n6400) );
  XOR U6326 ( .A(n6401), .B(n6402), .Z(n6335) );
  XOR U6327 ( .A(n6403), .B(n6404), .Z(n6402) );
  AND U6328 ( .A(\stack[1][20] ), .B(\stack[0][9] ), .Z(n6337) );
  AND U6329 ( .A(n6405), .B(n6406), .Z(n6338) );
  NANDN U6330 ( .A(n6342), .B(n6407), .Z(n6406) );
  NANDN U6331 ( .A(n6345), .B(n6408), .Z(n6405) );
  NAND U6332 ( .A(n6344), .B(n6342), .Z(n6408) );
  XOR U6333 ( .A(n6409), .B(n6410), .Z(n6342) );
  XNOR U6334 ( .A(n6411), .B(n6412), .Z(n6410) );
  IV U6335 ( .A(n6407), .Z(n6344) );
  NOR U6336 ( .A(n3092), .B(n2803), .Z(n6407) );
  AND U6337 ( .A(n6413), .B(n6414), .Z(n6345) );
  NANDN U6338 ( .A(n6350), .B(n6352), .Z(n6414) );
  NANDN U6339 ( .A(n6353), .B(n6415), .Z(n6413) );
  NANDN U6340 ( .A(n6352), .B(n6350), .Z(n6415) );
  XOR U6341 ( .A(n6416), .B(n6417), .Z(n6350) );
  XOR U6342 ( .A(n6418), .B(n6419), .Z(n6417) );
  AND U6343 ( .A(\stack[1][20] ), .B(\stack[0][7] ), .Z(n6352) );
  AND U6344 ( .A(n6420), .B(n6421), .Z(n6353) );
  NANDN U6345 ( .A(n6357), .B(n6422), .Z(n6421) );
  NANDN U6346 ( .A(n6360), .B(n6423), .Z(n6420) );
  NAND U6347 ( .A(n6359), .B(n6357), .Z(n6423) );
  XOR U6348 ( .A(n6424), .B(n6425), .Z(n6357) );
  XNOR U6349 ( .A(n6426), .B(n6427), .Z(n6425) );
  IV U6350 ( .A(n6422), .Z(n6359) );
  NOR U6351 ( .A(n3092), .B(n2755), .Z(n6422) );
  AND U6352 ( .A(n6428), .B(n6429), .Z(n6360) );
  NANDN U6353 ( .A(n6365), .B(n6367), .Z(n6429) );
  NANDN U6354 ( .A(n6368), .B(n6430), .Z(n6428) );
  NANDN U6355 ( .A(n6367), .B(n6365), .Z(n6430) );
  XOR U6356 ( .A(n6431), .B(n6432), .Z(n6365) );
  XOR U6357 ( .A(n6433), .B(n6434), .Z(n6432) );
  AND U6358 ( .A(\stack[1][20] ), .B(\stack[0][5] ), .Z(n6367) );
  AND U6359 ( .A(n6435), .B(n6436), .Z(n6368) );
  NANDN U6360 ( .A(n6372), .B(n6437), .Z(n6436) );
  NANDN U6361 ( .A(n6375), .B(n6438), .Z(n6435) );
  NAND U6362 ( .A(n6374), .B(n6372), .Z(n6438) );
  XOR U6363 ( .A(n6439), .B(n6440), .Z(n6372) );
  XNOR U6364 ( .A(n6441), .B(n6442), .Z(n6440) );
  IV U6365 ( .A(n6437), .Z(n6374) );
  NOR U6366 ( .A(n3092), .B(n2707), .Z(n6437) );
  AND U6367 ( .A(n6443), .B(n6444), .Z(n6375) );
  NANDN U6368 ( .A(n6380), .B(n6382), .Z(n6444) );
  NANDN U6369 ( .A(n6383), .B(n6445), .Z(n6443) );
  NANDN U6370 ( .A(n6382), .B(n6380), .Z(n6445) );
  XNOR U6371 ( .A(n6446), .B(n6447), .Z(n6380) );
  XNOR U6372 ( .A(n6448), .B(n6449), .Z(n6447) );
  AND U6373 ( .A(\stack[1][20] ), .B(\stack[0][3] ), .Z(n6382) );
  AND U6374 ( .A(n6450), .B(n6451), .Z(n6383) );
  NANDN U6375 ( .A(n6387), .B(n6389), .Z(n6451) );
  NAND U6376 ( .A(n6452), .B(n6390), .Z(n6450) );
  ANDN U6377 ( .B(n6453), .A(n6395), .Z(n6390) );
  NAND U6378 ( .A(\stack[1][20] ), .B(\stack[0][1] ), .Z(n6395) );
  AND U6379 ( .A(\stack[0][0] ), .B(\stack[1][21] ), .Z(n6453) );
  NANDN U6380 ( .A(n6389), .B(n6387), .Z(n6452) );
  XNOR U6381 ( .A(n6454), .B(n6455), .Z(n6387) );
  NAND U6382 ( .A(\stack[0][0] ), .B(\stack[1][22] ), .Z(n6455) );
  AND U6383 ( .A(\stack[1][20] ), .B(\stack[0][2] ), .Z(n6389) );
  ANDN U6384 ( .B(\stack[0][10] ), .A(n3092), .Z(n3508) );
  IV U6385 ( .A(\stack[1][20] ), .Z(n3092) );
  XNOR U6386 ( .A(n3518), .B(n6456), .Z(n3507) );
  XNOR U6387 ( .A(n3517), .B(n3519), .Z(n6456) );
  AND U6388 ( .A(n6457), .B(n6458), .Z(n3519) );
  NANDN U6389 ( .A(n6401), .B(n6459), .Z(n6458) );
  NANDN U6390 ( .A(n6404), .B(n6460), .Z(n6457) );
  NAND U6391 ( .A(n6403), .B(n6401), .Z(n6460) );
  XOR U6392 ( .A(n6461), .B(n6462), .Z(n6401) );
  XNOR U6393 ( .A(n6463), .B(n6464), .Z(n6462) );
  IV U6394 ( .A(n6459), .Z(n6403) );
  NOR U6395 ( .A(n3116), .B(n2803), .Z(n6459) );
  IV U6396 ( .A(\stack[0][8] ), .Z(n2803) );
  AND U6397 ( .A(n6465), .B(n6466), .Z(n6404) );
  NANDN U6398 ( .A(n6409), .B(n6411), .Z(n6466) );
  NANDN U6399 ( .A(n6412), .B(n6467), .Z(n6465) );
  NANDN U6400 ( .A(n6411), .B(n6409), .Z(n6467) );
  XOR U6401 ( .A(n6468), .B(n6469), .Z(n6409) );
  XOR U6402 ( .A(n6470), .B(n6471), .Z(n6469) );
  AND U6403 ( .A(\stack[1][21] ), .B(\stack[0][7] ), .Z(n6411) );
  AND U6404 ( .A(n6472), .B(n6473), .Z(n6412) );
  NANDN U6405 ( .A(n6416), .B(n6474), .Z(n6473) );
  NANDN U6406 ( .A(n6419), .B(n6475), .Z(n6472) );
  NAND U6407 ( .A(n6418), .B(n6416), .Z(n6475) );
  XOR U6408 ( .A(n6476), .B(n6477), .Z(n6416) );
  XNOR U6409 ( .A(n6478), .B(n6479), .Z(n6477) );
  IV U6410 ( .A(n6474), .Z(n6418) );
  NOR U6411 ( .A(n3116), .B(n2755), .Z(n6474) );
  AND U6412 ( .A(n6480), .B(n6481), .Z(n6419) );
  NANDN U6413 ( .A(n6424), .B(n6426), .Z(n6481) );
  NANDN U6414 ( .A(n6427), .B(n6482), .Z(n6480) );
  NANDN U6415 ( .A(n6426), .B(n6424), .Z(n6482) );
  XOR U6416 ( .A(n6483), .B(n6484), .Z(n6424) );
  XOR U6417 ( .A(n6485), .B(n6486), .Z(n6484) );
  AND U6418 ( .A(\stack[1][21] ), .B(\stack[0][5] ), .Z(n6426) );
  AND U6419 ( .A(n6487), .B(n6488), .Z(n6427) );
  NANDN U6420 ( .A(n6431), .B(n6489), .Z(n6488) );
  NANDN U6421 ( .A(n6434), .B(n6490), .Z(n6487) );
  NAND U6422 ( .A(n6433), .B(n6431), .Z(n6490) );
  XOR U6423 ( .A(n6491), .B(n6492), .Z(n6431) );
  XNOR U6424 ( .A(n6493), .B(n6494), .Z(n6492) );
  IV U6425 ( .A(n6489), .Z(n6433) );
  NOR U6426 ( .A(n3116), .B(n2707), .Z(n6489) );
  AND U6427 ( .A(n6495), .B(n6496), .Z(n6434) );
  NANDN U6428 ( .A(n6439), .B(n6441), .Z(n6496) );
  NANDN U6429 ( .A(n6442), .B(n6497), .Z(n6495) );
  NANDN U6430 ( .A(n6441), .B(n6439), .Z(n6497) );
  XNOR U6431 ( .A(n6498), .B(n6499), .Z(n6439) );
  XNOR U6432 ( .A(n6500), .B(n6501), .Z(n6499) );
  AND U6433 ( .A(\stack[1][21] ), .B(\stack[0][3] ), .Z(n6441) );
  AND U6434 ( .A(n6502), .B(n6503), .Z(n6442) );
  NANDN U6435 ( .A(n6446), .B(n6448), .Z(n6503) );
  NAND U6436 ( .A(n6504), .B(n6449), .Z(n6502) );
  ANDN U6437 ( .B(n6505), .A(n6454), .Z(n6449) );
  NAND U6438 ( .A(\stack[1][21] ), .B(\stack[0][1] ), .Z(n6454) );
  AND U6439 ( .A(\stack[0][0] ), .B(\stack[1][22] ), .Z(n6505) );
  NANDN U6440 ( .A(n6448), .B(n6446), .Z(n6504) );
  XNOR U6441 ( .A(n6506), .B(n6507), .Z(n6446) );
  NAND U6442 ( .A(\stack[0][0] ), .B(\stack[1][23] ), .Z(n6507) );
  AND U6443 ( .A(\stack[1][21] ), .B(\stack[0][2] ), .Z(n6448) );
  NOR U6444 ( .A(n3116), .B(n2827), .Z(n3517) );
  IV U6445 ( .A(\stack[0][9] ), .Z(n2827) );
  IV U6446 ( .A(\stack[1][21] ), .Z(n3116) );
  XNOR U6447 ( .A(n3525), .B(n6508), .Z(n3518) );
  XNOR U6448 ( .A(n3526), .B(n3527), .Z(n6508) );
  AND U6449 ( .A(n6509), .B(n6510), .Z(n3527) );
  NANDN U6450 ( .A(n6461), .B(n6463), .Z(n6510) );
  NANDN U6451 ( .A(n6464), .B(n6511), .Z(n6509) );
  NANDN U6452 ( .A(n6463), .B(n6461), .Z(n6511) );
  XOR U6453 ( .A(n6512), .B(n6513), .Z(n6461) );
  XOR U6454 ( .A(n6514), .B(n6515), .Z(n6513) );
  AND U6455 ( .A(\stack[1][22] ), .B(\stack[0][7] ), .Z(n6463) );
  AND U6456 ( .A(n6516), .B(n6517), .Z(n6464) );
  NANDN U6457 ( .A(n6468), .B(n6518), .Z(n6517) );
  NANDN U6458 ( .A(n6471), .B(n6519), .Z(n6516) );
  NAND U6459 ( .A(n6470), .B(n6468), .Z(n6519) );
  XOR U6460 ( .A(n6520), .B(n6521), .Z(n6468) );
  XNOR U6461 ( .A(n6522), .B(n6523), .Z(n6521) );
  IV U6462 ( .A(n6518), .Z(n6470) );
  NOR U6463 ( .A(n3140), .B(n2755), .Z(n6518) );
  AND U6464 ( .A(n6524), .B(n6525), .Z(n6471) );
  NANDN U6465 ( .A(n6476), .B(n6478), .Z(n6525) );
  NANDN U6466 ( .A(n6479), .B(n6526), .Z(n6524) );
  NANDN U6467 ( .A(n6478), .B(n6476), .Z(n6526) );
  XOR U6468 ( .A(n6527), .B(n6528), .Z(n6476) );
  XOR U6469 ( .A(n6529), .B(n6530), .Z(n6528) );
  AND U6470 ( .A(\stack[1][22] ), .B(\stack[0][5] ), .Z(n6478) );
  AND U6471 ( .A(n6531), .B(n6532), .Z(n6479) );
  NANDN U6472 ( .A(n6483), .B(n6533), .Z(n6532) );
  NANDN U6473 ( .A(n6486), .B(n6534), .Z(n6531) );
  NAND U6474 ( .A(n6485), .B(n6483), .Z(n6534) );
  XOR U6475 ( .A(n6535), .B(n6536), .Z(n6483) );
  XNOR U6476 ( .A(n6537), .B(n6538), .Z(n6536) );
  IV U6477 ( .A(n6533), .Z(n6485) );
  NOR U6478 ( .A(n3140), .B(n2707), .Z(n6533) );
  AND U6479 ( .A(n6539), .B(n6540), .Z(n6486) );
  NANDN U6480 ( .A(n6491), .B(n6493), .Z(n6540) );
  NANDN U6481 ( .A(n6494), .B(n6541), .Z(n6539) );
  NANDN U6482 ( .A(n6493), .B(n6491), .Z(n6541) );
  XNOR U6483 ( .A(n6542), .B(n6543), .Z(n6491) );
  XNOR U6484 ( .A(n6544), .B(n6545), .Z(n6543) );
  AND U6485 ( .A(\stack[1][22] ), .B(\stack[0][3] ), .Z(n6493) );
  AND U6486 ( .A(n6546), .B(n6547), .Z(n6494) );
  NANDN U6487 ( .A(n6498), .B(n6500), .Z(n6547) );
  NAND U6488 ( .A(n6548), .B(n6501), .Z(n6546) );
  ANDN U6489 ( .B(n6549), .A(n6506), .Z(n6501) );
  NAND U6490 ( .A(\stack[1][22] ), .B(\stack[0][1] ), .Z(n6506) );
  AND U6491 ( .A(\stack[0][0] ), .B(\stack[1][23] ), .Z(n6549) );
  NANDN U6492 ( .A(n6500), .B(n6498), .Z(n6548) );
  XNOR U6493 ( .A(n6550), .B(n6551), .Z(n6498) );
  NAND U6494 ( .A(\stack[0][0] ), .B(\stack[1][24] ), .Z(n6551) );
  AND U6495 ( .A(\stack[1][22] ), .B(\stack[0][2] ), .Z(n6500) );
  ANDN U6496 ( .B(\stack[0][8] ), .A(n3140), .Z(n3526) );
  IV U6497 ( .A(\stack[1][22] ), .Z(n3140) );
  XNOR U6498 ( .A(n3472), .B(n6552), .Z(n3525) );
  XNOR U6499 ( .A(n3471), .B(n3473), .Z(n6552) );
  AND U6500 ( .A(n6553), .B(n6554), .Z(n3473) );
  NANDN U6501 ( .A(n6512), .B(n6555), .Z(n6554) );
  NANDN U6502 ( .A(n6515), .B(n6556), .Z(n6553) );
  NAND U6503 ( .A(n6514), .B(n6512), .Z(n6556) );
  XOR U6504 ( .A(n6557), .B(n6558), .Z(n6512) );
  XNOR U6505 ( .A(n6559), .B(n6560), .Z(n6558) );
  IV U6506 ( .A(n6555), .Z(n6514) );
  NOR U6507 ( .A(n3164), .B(n2755), .Z(n6555) );
  IV U6508 ( .A(\stack[0][6] ), .Z(n2755) );
  AND U6509 ( .A(n6561), .B(n6562), .Z(n6515) );
  NANDN U6510 ( .A(n6520), .B(n6522), .Z(n6562) );
  NANDN U6511 ( .A(n6523), .B(n6563), .Z(n6561) );
  NANDN U6512 ( .A(n6522), .B(n6520), .Z(n6563) );
  XOR U6513 ( .A(n6564), .B(n6565), .Z(n6520) );
  XOR U6514 ( .A(n6566), .B(n6567), .Z(n6565) );
  AND U6515 ( .A(\stack[1][23] ), .B(\stack[0][5] ), .Z(n6522) );
  AND U6516 ( .A(n6568), .B(n6569), .Z(n6523) );
  NANDN U6517 ( .A(n6527), .B(n6570), .Z(n6569) );
  NANDN U6518 ( .A(n6530), .B(n6571), .Z(n6568) );
  NAND U6519 ( .A(n6529), .B(n6527), .Z(n6571) );
  XOR U6520 ( .A(n6572), .B(n6573), .Z(n6527) );
  XNOR U6521 ( .A(n6574), .B(n6575), .Z(n6573) );
  IV U6522 ( .A(n6570), .Z(n6529) );
  NOR U6523 ( .A(n3164), .B(n2707), .Z(n6570) );
  AND U6524 ( .A(n6576), .B(n6577), .Z(n6530) );
  NANDN U6525 ( .A(n6535), .B(n6537), .Z(n6577) );
  NANDN U6526 ( .A(n6538), .B(n6578), .Z(n6576) );
  NANDN U6527 ( .A(n6537), .B(n6535), .Z(n6578) );
  XNOR U6528 ( .A(n6579), .B(n6580), .Z(n6535) );
  XNOR U6529 ( .A(n6581), .B(n6582), .Z(n6580) );
  AND U6530 ( .A(\stack[1][23] ), .B(\stack[0][3] ), .Z(n6537) );
  AND U6531 ( .A(n6583), .B(n6584), .Z(n6538) );
  NANDN U6532 ( .A(n6542), .B(n6544), .Z(n6584) );
  NAND U6533 ( .A(n6585), .B(n6545), .Z(n6583) );
  ANDN U6534 ( .B(n6586), .A(n6550), .Z(n6545) );
  NAND U6535 ( .A(\stack[1][23] ), .B(\stack[0][1] ), .Z(n6550) );
  AND U6536 ( .A(\stack[0][0] ), .B(\stack[1][24] ), .Z(n6586) );
  NANDN U6537 ( .A(n6544), .B(n6542), .Z(n6585) );
  XNOR U6538 ( .A(n6587), .B(n6588), .Z(n6542) );
  NAND U6539 ( .A(\stack[0][0] ), .B(\stack[1][25] ), .Z(n6588) );
  AND U6540 ( .A(\stack[1][23] ), .B(\stack[0][2] ), .Z(n6544) );
  NOR U6541 ( .A(n3164), .B(n2779), .Z(n3471) );
  IV U6542 ( .A(\stack[0][7] ), .Z(n2779) );
  IV U6543 ( .A(\stack[1][23] ), .Z(n3164) );
  XNOR U6544 ( .A(n3481), .B(n6589), .Z(n3472) );
  XNOR U6545 ( .A(n3482), .B(n3483), .Z(n6589) );
  AND U6546 ( .A(n6590), .B(n6591), .Z(n3483) );
  NANDN U6547 ( .A(n6557), .B(n6559), .Z(n6591) );
  NANDN U6548 ( .A(n6560), .B(n6592), .Z(n6590) );
  NANDN U6549 ( .A(n6559), .B(n6557), .Z(n6592) );
  XOR U6550 ( .A(n6593), .B(n6594), .Z(n6557) );
  XOR U6551 ( .A(n6595), .B(n6596), .Z(n6594) );
  AND U6552 ( .A(\stack[1][24] ), .B(\stack[0][5] ), .Z(n6559) );
  AND U6553 ( .A(n6597), .B(n6598), .Z(n6560) );
  NANDN U6554 ( .A(n6564), .B(n6599), .Z(n6598) );
  NANDN U6555 ( .A(n6567), .B(n6600), .Z(n6597) );
  NAND U6556 ( .A(n6566), .B(n6564), .Z(n6600) );
  XOR U6557 ( .A(n6601), .B(n6602), .Z(n6564) );
  XNOR U6558 ( .A(n6603), .B(n6604), .Z(n6602) );
  IV U6559 ( .A(n6599), .Z(n6566) );
  NOR U6560 ( .A(n3188), .B(n2707), .Z(n6599) );
  AND U6561 ( .A(n6605), .B(n6606), .Z(n6567) );
  NANDN U6562 ( .A(n6572), .B(n6574), .Z(n6606) );
  NANDN U6563 ( .A(n6575), .B(n6607), .Z(n6605) );
  NANDN U6564 ( .A(n6574), .B(n6572), .Z(n6607) );
  XNOR U6565 ( .A(n6608), .B(n6609), .Z(n6572) );
  XNOR U6566 ( .A(n6610), .B(n6611), .Z(n6609) );
  AND U6567 ( .A(\stack[1][24] ), .B(\stack[0][3] ), .Z(n6574) );
  AND U6568 ( .A(n6612), .B(n6613), .Z(n6575) );
  NANDN U6569 ( .A(n6579), .B(n6581), .Z(n6613) );
  NAND U6570 ( .A(n6614), .B(n6582), .Z(n6612) );
  ANDN U6571 ( .B(n6615), .A(n6587), .Z(n6582) );
  NAND U6572 ( .A(\stack[1][24] ), .B(\stack[0][1] ), .Z(n6587) );
  AND U6573 ( .A(\stack[0][0] ), .B(\stack[1][25] ), .Z(n6615) );
  NANDN U6574 ( .A(n6581), .B(n6579), .Z(n6614) );
  XNOR U6575 ( .A(n6616), .B(n6617), .Z(n6579) );
  NAND U6576 ( .A(\stack[0][0] ), .B(\stack[1][26] ), .Z(n6617) );
  AND U6577 ( .A(\stack[1][24] ), .B(\stack[0][2] ), .Z(n6581) );
  ANDN U6578 ( .B(\stack[0][6] ), .A(n3188), .Z(n3482) );
  IV U6579 ( .A(\stack[1][24] ), .Z(n3188) );
  XNOR U6580 ( .A(n3492), .B(n6618), .Z(n3481) );
  XNOR U6581 ( .A(n3491), .B(n3493), .Z(n6618) );
  AND U6582 ( .A(n6619), .B(n6620), .Z(n3493) );
  NANDN U6583 ( .A(n6593), .B(n6621), .Z(n6620) );
  NANDN U6584 ( .A(n6596), .B(n6622), .Z(n6619) );
  NAND U6585 ( .A(n6595), .B(n6593), .Z(n6622) );
  XOR U6586 ( .A(n6623), .B(n6624), .Z(n6593) );
  XNOR U6587 ( .A(n6625), .B(n6626), .Z(n6624) );
  IV U6588 ( .A(n6621), .Z(n6595) );
  NOR U6589 ( .A(n3212), .B(n2707), .Z(n6621) );
  IV U6590 ( .A(\stack[0][4] ), .Z(n2707) );
  AND U6591 ( .A(n6627), .B(n6628), .Z(n6596) );
  NANDN U6592 ( .A(n6601), .B(n6603), .Z(n6628) );
  NANDN U6593 ( .A(n6604), .B(n6629), .Z(n6627) );
  NANDN U6594 ( .A(n6603), .B(n6601), .Z(n6629) );
  XNOR U6595 ( .A(n6630), .B(n6631), .Z(n6601) );
  XNOR U6596 ( .A(n6632), .B(n6633), .Z(n6631) );
  AND U6597 ( .A(\stack[1][25] ), .B(\stack[0][3] ), .Z(n6603) );
  AND U6598 ( .A(n6634), .B(n6635), .Z(n6604) );
  NANDN U6599 ( .A(n6608), .B(n6610), .Z(n6635) );
  NAND U6600 ( .A(n6636), .B(n6611), .Z(n6634) );
  ANDN U6601 ( .B(n6637), .A(n6616), .Z(n6611) );
  NAND U6602 ( .A(\stack[1][25] ), .B(\stack[0][1] ), .Z(n6616) );
  AND U6603 ( .A(\stack[0][0] ), .B(\stack[1][26] ), .Z(n6637) );
  NANDN U6604 ( .A(n6610), .B(n6608), .Z(n6636) );
  XNOR U6605 ( .A(n6638), .B(n6639), .Z(n6608) );
  NAND U6606 ( .A(\stack[0][0] ), .B(\stack[1][27] ), .Z(n6639) );
  AND U6607 ( .A(\stack[1][25] ), .B(\stack[0][2] ), .Z(n6610) );
  NOR U6608 ( .A(n3212), .B(n2731), .Z(n3491) );
  IV U6609 ( .A(\stack[0][5] ), .Z(n2731) );
  IV U6610 ( .A(\stack[1][25] ), .Z(n3212) );
  XNOR U6611 ( .A(n3499), .B(n6640), .Z(n3492) );
  XNOR U6612 ( .A(n3500), .B(n3501), .Z(n6640) );
  AND U6613 ( .A(n6641), .B(n6642), .Z(n3501) );
  NANDN U6614 ( .A(n6623), .B(n6625), .Z(n6642) );
  NANDN U6615 ( .A(n6626), .B(n6643), .Z(n6641) );
  NANDN U6616 ( .A(n6625), .B(n6623), .Z(n6643) );
  XNOR U6617 ( .A(n6644), .B(n6645), .Z(n6623) );
  XNOR U6618 ( .A(n6646), .B(n6647), .Z(n6645) );
  AND U6619 ( .A(\stack[1][26] ), .B(\stack[0][3] ), .Z(n6625) );
  AND U6620 ( .A(n6648), .B(n6649), .Z(n6626) );
  NANDN U6621 ( .A(n6630), .B(n6632), .Z(n6649) );
  NAND U6622 ( .A(n6650), .B(n6633), .Z(n6648) );
  ANDN U6623 ( .B(n6651), .A(n6638), .Z(n6633) );
  NAND U6624 ( .A(\stack[1][26] ), .B(\stack[0][1] ), .Z(n6638) );
  AND U6625 ( .A(\stack[0][0] ), .B(\stack[1][27] ), .Z(n6651) );
  NANDN U6626 ( .A(n6632), .B(n6630), .Z(n6650) );
  XNOR U6627 ( .A(n6652), .B(n6653), .Z(n6630) );
  NAND U6628 ( .A(\stack[0][0] ), .B(\stack[1][28] ), .Z(n6653) );
  AND U6629 ( .A(\stack[1][26] ), .B(\stack[0][2] ), .Z(n6632) );
  ANDN U6630 ( .B(\stack[0][4] ), .A(n3236), .Z(n3500) );
  IV U6631 ( .A(\stack[1][26] ), .Z(n3236) );
  XNOR U6632 ( .A(n3458), .B(n6654), .Z(n3499) );
  XNOR U6633 ( .A(n3457), .B(n3459), .Z(n6654) );
  AND U6634 ( .A(n6655), .B(n6656), .Z(n3459) );
  NANDN U6635 ( .A(n6644), .B(n6646), .Z(n6656) );
  NAND U6636 ( .A(n6657), .B(n6647), .Z(n6655) );
  ANDN U6637 ( .B(n6658), .A(n6652), .Z(n6647) );
  NAND U6638 ( .A(\stack[1][27] ), .B(\stack[0][1] ), .Z(n6652) );
  AND U6639 ( .A(\stack[0][0] ), .B(\stack[1][28] ), .Z(n6658) );
  NANDN U6640 ( .A(n6646), .B(n6644), .Z(n6657) );
  XNOR U6641 ( .A(n6659), .B(n6660), .Z(n6644) );
  NAND U6642 ( .A(\stack[0][0] ), .B(\stack[1][29] ), .Z(n6660) );
  AND U6643 ( .A(\stack[1][27] ), .B(\stack[0][2] ), .Z(n6646) );
  NOR U6644 ( .A(n3260), .B(n2683), .Z(n3457) );
  IV U6645 ( .A(\stack[0][3] ), .Z(n2683) );
  IV U6646 ( .A(\stack[1][27] ), .Z(n3260) );
  XNOR U6647 ( .A(n3465), .B(n6661), .Z(n3458) );
  XOR U6648 ( .A(n3467), .B(n3466), .Z(n6661) );
  AND U6649 ( .A(\stack[1][28] ), .B(\stack[0][2] ), .Z(n3466) );
  NANDN U6650 ( .A(n6659), .B(n6662), .Z(n3467) );
  AND U6651 ( .A(\stack[0][0] ), .B(\stack[1][29] ), .Z(n6662) );
  NAND U6652 ( .A(\stack[1][28] ), .B(\stack[0][1] ), .Z(n6659) );
  XOR U6653 ( .A(n3448), .B(n6663), .Z(n3465) );
  NAND U6654 ( .A(\stack[0][0] ), .B(\stack[1][30] ), .Z(n6663) );
  NAND U6655 ( .A(\stack[1][29] ), .B(\stack[0][1] ), .Z(n3448) );
  XOR U6656 ( .A(\stack[1][31] ), .B(\stack[0][31] ), .Z(n3350) );
  AND U6657 ( .A(n6664), .B(n6665), .Z(n3343) );
  NAND U6658 ( .A(\stack[1][31] ), .B(n6666), .Z(n6665) );
  ANDN U6659 ( .B(\stack[0][31] ), .A(n2611), .Z(n6666) );
  NAND U6660 ( .A(n6667), .B(opcode[2]), .Z(n2611) );
  NAND U6661 ( .A(n6668), .B(n2613), .Z(n6664) );
  ANDN U6662 ( .B(opcode[0]), .A(n6669), .Z(n2613) );
  AND U6663 ( .A(n6670), .B(n6671), .Z(n3341) );
  NAND U6664 ( .A(\stack[0][31] ), .B(n2618), .Z(n6671) );
  ANDN U6665 ( .B(n6672), .A(opcode[0]), .Z(n2618) );
  XOR U6666 ( .A(n6673), .B(n6674), .Z(n6670) );
  XOR U6667 ( .A(n6675), .B(n6676), .Z(n6674) );
  NAND U6668 ( .A(n6677), .B(n6678), .Z(n6676) );
  NANDN U6669 ( .A(n3334), .B(n6679), .Z(n6678) );
  OR U6670 ( .A(n3333), .B(n3331), .Z(n6679) );
  AND U6671 ( .A(n6680), .B(n6681), .Z(n3334) );
  NAND U6672 ( .A(\stack[0][30] ), .B(n6682), .Z(n6681) );
  NAND U6673 ( .A(\stack[0][30] ), .B(n6683), .Z(n6680) );
  NAND U6674 ( .A(n3333), .B(n3331), .Z(n6677) );
  XOR U6675 ( .A(n6684), .B(n6685), .Z(n3331) );
  NAND U6676 ( .A(n6686), .B(n6687), .Z(n6685) );
  NAND U6677 ( .A(\stack[1][30] ), .B(n6683), .Z(n6687) );
  AND U6678 ( .A(n6688), .B(n6689), .Z(n6686) );
  NAND U6679 ( .A(\stack[0][30] ), .B(n3339), .Z(n6689) );
  NAND U6680 ( .A(\stack[1][30] ), .B(n6682), .Z(n6688) );
  NAND U6681 ( .A(n6690), .B(n6691), .Z(n3333) );
  NANDN U6682 ( .A(n3311), .B(n6692), .Z(n6691) );
  NANDN U6683 ( .A(n3312), .B(n6693), .Z(n6690) );
  NAND U6684 ( .A(n3309), .B(n3311), .Z(n6693) );
  AND U6685 ( .A(n6694), .B(n6695), .Z(n3311) );
  NANDN U6686 ( .A(n3288), .B(n6696), .Z(n6695) );
  NANDN U6687 ( .A(n3289), .B(n6697), .Z(n6694) );
  NAND U6688 ( .A(n3286), .B(n3288), .Z(n6697) );
  AND U6689 ( .A(n6698), .B(n6699), .Z(n3288) );
  NANDN U6690 ( .A(n3265), .B(n6700), .Z(n6699) );
  NANDN U6691 ( .A(n3266), .B(n6701), .Z(n6698) );
  NAND U6692 ( .A(n3263), .B(n3265), .Z(n6701) );
  AND U6693 ( .A(n6702), .B(n6703), .Z(n3265) );
  NANDN U6694 ( .A(n3241), .B(n6704), .Z(n6703) );
  NANDN U6695 ( .A(n3242), .B(n6705), .Z(n6702) );
  NAND U6696 ( .A(n3239), .B(n3241), .Z(n6705) );
  AND U6697 ( .A(n6706), .B(n6707), .Z(n3241) );
  NANDN U6698 ( .A(n3217), .B(n6708), .Z(n6707) );
  NANDN U6699 ( .A(n3218), .B(n6709), .Z(n6706) );
  NAND U6700 ( .A(n3215), .B(n3217), .Z(n6709) );
  AND U6701 ( .A(n6710), .B(n6711), .Z(n3217) );
  NANDN U6702 ( .A(n3193), .B(n6712), .Z(n6711) );
  NANDN U6703 ( .A(n3194), .B(n6713), .Z(n6710) );
  NAND U6704 ( .A(n3191), .B(n3193), .Z(n6713) );
  AND U6705 ( .A(n6714), .B(n6715), .Z(n3193) );
  NANDN U6706 ( .A(n3169), .B(n6716), .Z(n6715) );
  NANDN U6707 ( .A(n3170), .B(n6717), .Z(n6714) );
  NAND U6708 ( .A(n3167), .B(n3169), .Z(n6717) );
  AND U6709 ( .A(n6718), .B(n6719), .Z(n3169) );
  NANDN U6710 ( .A(n3145), .B(n6720), .Z(n6719) );
  NANDN U6711 ( .A(n3146), .B(n6721), .Z(n6718) );
  NAND U6712 ( .A(n3143), .B(n3145), .Z(n6721) );
  AND U6713 ( .A(n6722), .B(n6723), .Z(n3145) );
  NANDN U6714 ( .A(n3121), .B(n6724), .Z(n6723) );
  NANDN U6715 ( .A(n3122), .B(n6725), .Z(n6722) );
  NAND U6716 ( .A(n3119), .B(n3121), .Z(n6725) );
  AND U6717 ( .A(n6726), .B(n6727), .Z(n3121) );
  NANDN U6718 ( .A(n3097), .B(n6728), .Z(n6727) );
  NANDN U6719 ( .A(n3098), .B(n6729), .Z(n6726) );
  NAND U6720 ( .A(n3095), .B(n3097), .Z(n6729) );
  AND U6721 ( .A(n6730), .B(n6731), .Z(n3097) );
  NANDN U6722 ( .A(n3073), .B(n6732), .Z(n6731) );
  NANDN U6723 ( .A(n3074), .B(n6733), .Z(n6730) );
  NAND U6724 ( .A(n3071), .B(n3073), .Z(n6733) );
  AND U6725 ( .A(n6734), .B(n6735), .Z(n3073) );
  NANDN U6726 ( .A(n3049), .B(n6736), .Z(n6735) );
  NANDN U6727 ( .A(n3050), .B(n6737), .Z(n6734) );
  NAND U6728 ( .A(n3047), .B(n3049), .Z(n6737) );
  AND U6729 ( .A(n6738), .B(n6739), .Z(n3049) );
  NANDN U6730 ( .A(n3025), .B(n6740), .Z(n6739) );
  NANDN U6731 ( .A(n3026), .B(n6741), .Z(n6738) );
  NAND U6732 ( .A(n3023), .B(n3025), .Z(n6741) );
  AND U6733 ( .A(n6742), .B(n6743), .Z(n3025) );
  NANDN U6734 ( .A(n3001), .B(n6744), .Z(n6743) );
  NANDN U6735 ( .A(n3002), .B(n6745), .Z(n6742) );
  NAND U6736 ( .A(n2999), .B(n3001), .Z(n6745) );
  AND U6737 ( .A(n6746), .B(n6747), .Z(n3001) );
  NANDN U6738 ( .A(n2977), .B(n6748), .Z(n6747) );
  NANDN U6739 ( .A(n2978), .B(n6749), .Z(n6746) );
  NAND U6740 ( .A(n2975), .B(n2977), .Z(n6749) );
  AND U6741 ( .A(n6750), .B(n6751), .Z(n2977) );
  NANDN U6742 ( .A(n2953), .B(n6752), .Z(n6751) );
  NANDN U6743 ( .A(n2954), .B(n6753), .Z(n6750) );
  NAND U6744 ( .A(n2951), .B(n2953), .Z(n6753) );
  AND U6745 ( .A(n6754), .B(n6755), .Z(n2953) );
  NANDN U6746 ( .A(n2929), .B(n6756), .Z(n6755) );
  NANDN U6747 ( .A(n2930), .B(n6757), .Z(n6754) );
  NAND U6748 ( .A(n2927), .B(n2929), .Z(n6757) );
  AND U6749 ( .A(n6758), .B(n6759), .Z(n2929) );
  NANDN U6750 ( .A(n2905), .B(n6760), .Z(n6759) );
  NANDN U6751 ( .A(n2906), .B(n6761), .Z(n6758) );
  NAND U6752 ( .A(n2903), .B(n2905), .Z(n6761) );
  AND U6753 ( .A(n6762), .B(n6763), .Z(n2905) );
  NANDN U6754 ( .A(n2881), .B(n6764), .Z(n6763) );
  NANDN U6755 ( .A(n2882), .B(n6765), .Z(n6762) );
  NAND U6756 ( .A(n2879), .B(n2881), .Z(n6765) );
  AND U6757 ( .A(n6766), .B(n6767), .Z(n2881) );
  NANDN U6758 ( .A(n2857), .B(n6768), .Z(n6767) );
  NANDN U6759 ( .A(n2858), .B(n6769), .Z(n6766) );
  NAND U6760 ( .A(n2855), .B(n2857), .Z(n6769) );
  AND U6761 ( .A(n6770), .B(n6771), .Z(n2857) );
  NANDN U6762 ( .A(n2833), .B(n2831), .Z(n6771) );
  NANDN U6763 ( .A(n2834), .B(n6772), .Z(n6770) );
  AND U6764 ( .A(n6773), .B(n6774), .Z(n2833) );
  NANDN U6765 ( .A(n2809), .B(n6775), .Z(n6774) );
  NANDN U6766 ( .A(n2810), .B(n6776), .Z(n6773) );
  NAND U6767 ( .A(n2807), .B(n2809), .Z(n6776) );
  AND U6768 ( .A(n6777), .B(n6778), .Z(n2809) );
  NANDN U6769 ( .A(n2785), .B(n6779), .Z(n6778) );
  NANDN U6770 ( .A(n2786), .B(n6780), .Z(n6777) );
  NAND U6771 ( .A(n2783), .B(n2785), .Z(n6780) );
  AND U6772 ( .A(n6781), .B(n6782), .Z(n2785) );
  NANDN U6773 ( .A(n2761), .B(n6783), .Z(n6782) );
  NANDN U6774 ( .A(n2762), .B(n6784), .Z(n6781) );
  NAND U6775 ( .A(n2759), .B(n2761), .Z(n6784) );
  AND U6776 ( .A(n6785), .B(n6786), .Z(n2761) );
  NANDN U6777 ( .A(n2737), .B(n6787), .Z(n6786) );
  NANDN U6778 ( .A(n2738), .B(n6788), .Z(n6785) );
  NAND U6779 ( .A(n2735), .B(n2737), .Z(n6788) );
  AND U6780 ( .A(n6789), .B(n6790), .Z(n2737) );
  NANDN U6781 ( .A(n2713), .B(n6791), .Z(n6790) );
  NANDN U6782 ( .A(n2714), .B(n6792), .Z(n6789) );
  NAND U6783 ( .A(n2711), .B(n2713), .Z(n6792) );
  AND U6784 ( .A(n6793), .B(n6794), .Z(n2713) );
  NANDN U6785 ( .A(n2689), .B(n6795), .Z(n6794) );
  NANDN U6786 ( .A(n2690), .B(n6796), .Z(n6793) );
  NAND U6787 ( .A(n2687), .B(n2689), .Z(n6796) );
  AND U6788 ( .A(n6797), .B(n6798), .Z(n2689) );
  NANDN U6789 ( .A(n2665), .B(n6799), .Z(n6798) );
  NANDN U6790 ( .A(n2666), .B(n6800), .Z(n6797) );
  NAND U6791 ( .A(n2663), .B(n2665), .Z(n6800) );
  AND U6792 ( .A(n6801), .B(n6802), .Z(n2665) );
  NANDN U6793 ( .A(n2642), .B(n6803), .Z(n6802) );
  NANDN U6794 ( .A(n2643), .B(n6804), .Z(n6801) );
  NAND U6795 ( .A(n2640), .B(n2642), .Z(n6804) );
  AND U6796 ( .A(n6805), .B(n6806), .Z(n2642) );
  NAND U6797 ( .A(n6684), .B(n2619), .Z(n6806) );
  NANDN U6798 ( .A(n2622), .B(n6807), .Z(n6805) );
  XOR U6799 ( .A(n6684), .B(n6808), .Z(n2619) );
  NAND U6800 ( .A(n6809), .B(n6810), .Z(n6808) );
  NAND U6801 ( .A(\stack[1][0] ), .B(n6683), .Z(n6810) );
  AND U6802 ( .A(n6811), .B(n6812), .Z(n6809) );
  NAND U6803 ( .A(\stack[0][0] ), .B(n3339), .Z(n6812) );
  NAND U6804 ( .A(\stack[1][0] ), .B(n6682), .Z(n6811) );
  AND U6805 ( .A(n6813), .B(n6814), .Z(n2622) );
  NAND U6806 ( .A(\stack[0][0] ), .B(n6682), .Z(n6814) );
  NAND U6807 ( .A(\stack[0][0] ), .B(n6683), .Z(n6813) );
  IV U6808 ( .A(n6803), .Z(n2640) );
  XOR U6809 ( .A(n6684), .B(n6815), .Z(n6803) );
  NAND U6810 ( .A(n6816), .B(n6817), .Z(n6815) );
  NAND U6811 ( .A(\stack[1][1] ), .B(n6683), .Z(n6817) );
  AND U6812 ( .A(n6818), .B(n6819), .Z(n6816) );
  NAND U6813 ( .A(\stack[0][1] ), .B(n3339), .Z(n6819) );
  NAND U6814 ( .A(\stack[1][1] ), .B(n6682), .Z(n6818) );
  AND U6815 ( .A(n6820), .B(n6821), .Z(n2643) );
  NAND U6816 ( .A(\stack[0][1] ), .B(n6682), .Z(n6821) );
  NAND U6817 ( .A(\stack[0][1] ), .B(n6683), .Z(n6820) );
  IV U6818 ( .A(n6799), .Z(n2663) );
  XOR U6819 ( .A(n6684), .B(n6822), .Z(n6799) );
  NAND U6820 ( .A(n6823), .B(n6824), .Z(n6822) );
  NAND U6821 ( .A(\stack[1][2] ), .B(n6683), .Z(n6824) );
  AND U6822 ( .A(n6825), .B(n6826), .Z(n6823) );
  NAND U6823 ( .A(\stack[0][2] ), .B(n3339), .Z(n6826) );
  NAND U6824 ( .A(\stack[1][2] ), .B(n6682), .Z(n6825) );
  AND U6825 ( .A(n6827), .B(n6828), .Z(n2666) );
  NAND U6826 ( .A(\stack[0][2] ), .B(n6682), .Z(n6828) );
  NAND U6827 ( .A(\stack[0][2] ), .B(n6683), .Z(n6827) );
  IV U6828 ( .A(n6795), .Z(n2687) );
  XOR U6829 ( .A(n6684), .B(n6829), .Z(n6795) );
  NAND U6830 ( .A(n6830), .B(n6831), .Z(n6829) );
  NAND U6831 ( .A(\stack[1][3] ), .B(n6683), .Z(n6831) );
  AND U6832 ( .A(n6832), .B(n6833), .Z(n6830) );
  NAND U6833 ( .A(\stack[0][3] ), .B(n3339), .Z(n6833) );
  NAND U6834 ( .A(\stack[1][3] ), .B(n6682), .Z(n6832) );
  AND U6835 ( .A(n6834), .B(n6835), .Z(n2690) );
  NAND U6836 ( .A(\stack[0][3] ), .B(n6682), .Z(n6835) );
  NAND U6837 ( .A(\stack[0][3] ), .B(n6683), .Z(n6834) );
  IV U6838 ( .A(n6791), .Z(n2711) );
  XOR U6839 ( .A(n6684), .B(n6836), .Z(n6791) );
  NAND U6840 ( .A(n6837), .B(n6838), .Z(n6836) );
  NAND U6841 ( .A(\stack[1][4] ), .B(n6683), .Z(n6838) );
  AND U6842 ( .A(n6839), .B(n6840), .Z(n6837) );
  NAND U6843 ( .A(\stack[0][4] ), .B(n3339), .Z(n6840) );
  NAND U6844 ( .A(\stack[1][4] ), .B(n6682), .Z(n6839) );
  AND U6845 ( .A(n6841), .B(n6842), .Z(n2714) );
  NAND U6846 ( .A(\stack[0][4] ), .B(n6682), .Z(n6842) );
  NAND U6847 ( .A(\stack[0][4] ), .B(n6683), .Z(n6841) );
  IV U6848 ( .A(n6787), .Z(n2735) );
  XOR U6849 ( .A(n6684), .B(n6843), .Z(n6787) );
  NAND U6850 ( .A(n6844), .B(n6845), .Z(n6843) );
  NAND U6851 ( .A(\stack[1][5] ), .B(n6683), .Z(n6845) );
  AND U6852 ( .A(n6846), .B(n6847), .Z(n6844) );
  NAND U6853 ( .A(\stack[0][5] ), .B(n3339), .Z(n6847) );
  NAND U6854 ( .A(\stack[1][5] ), .B(n6682), .Z(n6846) );
  AND U6855 ( .A(n6848), .B(n6849), .Z(n2738) );
  NAND U6856 ( .A(\stack[0][5] ), .B(n6682), .Z(n6849) );
  NAND U6857 ( .A(\stack[0][5] ), .B(n6683), .Z(n6848) );
  IV U6858 ( .A(n6783), .Z(n2759) );
  XOR U6859 ( .A(n6684), .B(n6850), .Z(n6783) );
  NAND U6860 ( .A(n6851), .B(n6852), .Z(n6850) );
  NAND U6861 ( .A(\stack[1][6] ), .B(n6683), .Z(n6852) );
  AND U6862 ( .A(n6853), .B(n6854), .Z(n6851) );
  NAND U6863 ( .A(\stack[0][6] ), .B(n3339), .Z(n6854) );
  NAND U6864 ( .A(\stack[1][6] ), .B(n6682), .Z(n6853) );
  AND U6865 ( .A(n6855), .B(n6856), .Z(n2762) );
  NAND U6866 ( .A(\stack[0][6] ), .B(n6682), .Z(n6856) );
  NAND U6867 ( .A(\stack[0][6] ), .B(n6683), .Z(n6855) );
  IV U6868 ( .A(n6779), .Z(n2783) );
  XOR U6869 ( .A(n6684), .B(n6857), .Z(n6779) );
  NAND U6870 ( .A(n6858), .B(n6859), .Z(n6857) );
  NAND U6871 ( .A(\stack[1][7] ), .B(n6683), .Z(n6859) );
  AND U6872 ( .A(n6860), .B(n6861), .Z(n6858) );
  NAND U6873 ( .A(\stack[0][7] ), .B(n3339), .Z(n6861) );
  NAND U6874 ( .A(\stack[1][7] ), .B(n6682), .Z(n6860) );
  AND U6875 ( .A(n6862), .B(n6863), .Z(n2786) );
  NAND U6876 ( .A(\stack[0][7] ), .B(n6682), .Z(n6863) );
  NAND U6877 ( .A(\stack[0][7] ), .B(n6683), .Z(n6862) );
  IV U6878 ( .A(n6775), .Z(n2807) );
  XOR U6879 ( .A(n6684), .B(n6864), .Z(n6775) );
  NAND U6880 ( .A(n6865), .B(n6866), .Z(n6864) );
  NAND U6881 ( .A(\stack[1][8] ), .B(n6683), .Z(n6866) );
  AND U6882 ( .A(n6867), .B(n6868), .Z(n6865) );
  NAND U6883 ( .A(\stack[0][8] ), .B(n3339), .Z(n6868) );
  NAND U6884 ( .A(\stack[1][8] ), .B(n6682), .Z(n6867) );
  AND U6885 ( .A(n6869), .B(n6870), .Z(n2810) );
  NAND U6886 ( .A(\stack[0][8] ), .B(n6682), .Z(n6870) );
  NAND U6887 ( .A(\stack[0][8] ), .B(n6683), .Z(n6869) );
  XOR U6888 ( .A(n6871), .B(n2621), .Z(n2831) );
  AND U6889 ( .A(n6872), .B(n6873), .Z(n6871) );
  NAND U6890 ( .A(\stack[1][9] ), .B(n6683), .Z(n6873) );
  AND U6891 ( .A(n6874), .B(n6875), .Z(n6872) );
  NAND U6892 ( .A(\stack[0][9] ), .B(n3339), .Z(n6875) );
  NAND U6893 ( .A(\stack[1][9] ), .B(n6682), .Z(n6874) );
  AND U6894 ( .A(n6876), .B(n6877), .Z(n2834) );
  NAND U6895 ( .A(\stack[0][9] ), .B(n6682), .Z(n6877) );
  NAND U6896 ( .A(\stack[0][9] ), .B(n6683), .Z(n6876) );
  IV U6897 ( .A(n6768), .Z(n2855) );
  XOR U6898 ( .A(n6684), .B(n6878), .Z(n6768) );
  NAND U6899 ( .A(n6879), .B(n6880), .Z(n6878) );
  NAND U6900 ( .A(\stack[1][10] ), .B(n6683), .Z(n6880) );
  AND U6901 ( .A(n6881), .B(n6882), .Z(n6879) );
  NAND U6902 ( .A(\stack[0][10] ), .B(n3339), .Z(n6882) );
  NAND U6903 ( .A(\stack[1][10] ), .B(n6682), .Z(n6881) );
  AND U6904 ( .A(n6883), .B(n6884), .Z(n2858) );
  NAND U6905 ( .A(\stack[0][10] ), .B(n6682), .Z(n6884) );
  NAND U6906 ( .A(\stack[0][10] ), .B(n6683), .Z(n6883) );
  IV U6907 ( .A(n6764), .Z(n2879) );
  XOR U6908 ( .A(n6684), .B(n6885), .Z(n6764) );
  NAND U6909 ( .A(n6886), .B(n6887), .Z(n6885) );
  NAND U6910 ( .A(\stack[1][11] ), .B(n6683), .Z(n6887) );
  AND U6911 ( .A(n6888), .B(n6889), .Z(n6886) );
  NAND U6912 ( .A(\stack[0][11] ), .B(n3339), .Z(n6889) );
  NAND U6913 ( .A(\stack[1][11] ), .B(n6682), .Z(n6888) );
  AND U6914 ( .A(n6890), .B(n6891), .Z(n2882) );
  NAND U6915 ( .A(\stack[0][11] ), .B(n6682), .Z(n6891) );
  NAND U6916 ( .A(\stack[0][11] ), .B(n6683), .Z(n6890) );
  IV U6917 ( .A(n6760), .Z(n2903) );
  XOR U6918 ( .A(n6684), .B(n6892), .Z(n6760) );
  NAND U6919 ( .A(n6893), .B(n6894), .Z(n6892) );
  NAND U6920 ( .A(\stack[1][12] ), .B(n6683), .Z(n6894) );
  AND U6921 ( .A(n6895), .B(n6896), .Z(n6893) );
  NAND U6922 ( .A(\stack[0][12] ), .B(n3339), .Z(n6896) );
  NAND U6923 ( .A(\stack[1][12] ), .B(n6682), .Z(n6895) );
  AND U6924 ( .A(n6897), .B(n6898), .Z(n2906) );
  NAND U6925 ( .A(\stack[0][12] ), .B(n6682), .Z(n6898) );
  NAND U6926 ( .A(\stack[0][12] ), .B(n6683), .Z(n6897) );
  IV U6927 ( .A(n6756), .Z(n2927) );
  XOR U6928 ( .A(n6684), .B(n6899), .Z(n6756) );
  NAND U6929 ( .A(n6900), .B(n6901), .Z(n6899) );
  NAND U6930 ( .A(\stack[1][13] ), .B(n6683), .Z(n6901) );
  AND U6931 ( .A(n6902), .B(n6903), .Z(n6900) );
  NAND U6932 ( .A(\stack[0][13] ), .B(n3339), .Z(n6903) );
  NAND U6933 ( .A(\stack[1][13] ), .B(n6682), .Z(n6902) );
  AND U6934 ( .A(n6904), .B(n6905), .Z(n2930) );
  NAND U6935 ( .A(\stack[0][13] ), .B(n6682), .Z(n6905) );
  NAND U6936 ( .A(\stack[0][13] ), .B(n6683), .Z(n6904) );
  IV U6937 ( .A(n6752), .Z(n2951) );
  XOR U6938 ( .A(n6684), .B(n6906), .Z(n6752) );
  NAND U6939 ( .A(n6907), .B(n6908), .Z(n6906) );
  NAND U6940 ( .A(\stack[1][14] ), .B(n6683), .Z(n6908) );
  AND U6941 ( .A(n6909), .B(n6910), .Z(n6907) );
  NAND U6942 ( .A(\stack[0][14] ), .B(n3339), .Z(n6910) );
  NAND U6943 ( .A(\stack[1][14] ), .B(n6682), .Z(n6909) );
  AND U6944 ( .A(n6911), .B(n6912), .Z(n2954) );
  NAND U6945 ( .A(\stack[0][14] ), .B(n6682), .Z(n6912) );
  NAND U6946 ( .A(\stack[0][14] ), .B(n6683), .Z(n6911) );
  IV U6947 ( .A(n6748), .Z(n2975) );
  XOR U6948 ( .A(n6684), .B(n6913), .Z(n6748) );
  NAND U6949 ( .A(n6914), .B(n6915), .Z(n6913) );
  NAND U6950 ( .A(\stack[1][15] ), .B(n6683), .Z(n6915) );
  AND U6951 ( .A(n6916), .B(n6917), .Z(n6914) );
  NAND U6952 ( .A(\stack[0][15] ), .B(n3339), .Z(n6917) );
  NAND U6953 ( .A(\stack[1][15] ), .B(n6682), .Z(n6916) );
  AND U6954 ( .A(n6918), .B(n6919), .Z(n2978) );
  NAND U6955 ( .A(\stack[0][15] ), .B(n6682), .Z(n6919) );
  NAND U6956 ( .A(\stack[0][15] ), .B(n6683), .Z(n6918) );
  IV U6957 ( .A(n6744), .Z(n2999) );
  XOR U6958 ( .A(n6684), .B(n6920), .Z(n6744) );
  NAND U6959 ( .A(n6921), .B(n6922), .Z(n6920) );
  NAND U6960 ( .A(\stack[1][16] ), .B(n6683), .Z(n6922) );
  AND U6961 ( .A(n6923), .B(n6924), .Z(n6921) );
  NAND U6962 ( .A(\stack[0][16] ), .B(n3339), .Z(n6924) );
  NAND U6963 ( .A(\stack[1][16] ), .B(n6682), .Z(n6923) );
  AND U6964 ( .A(n6925), .B(n6926), .Z(n3002) );
  NAND U6965 ( .A(\stack[0][16] ), .B(n6682), .Z(n6926) );
  NAND U6966 ( .A(\stack[0][16] ), .B(n6683), .Z(n6925) );
  IV U6967 ( .A(n6740), .Z(n3023) );
  XOR U6968 ( .A(n6684), .B(n6927), .Z(n6740) );
  NAND U6969 ( .A(n6928), .B(n6929), .Z(n6927) );
  NAND U6970 ( .A(\stack[1][17] ), .B(n6683), .Z(n6929) );
  AND U6971 ( .A(n6930), .B(n6931), .Z(n6928) );
  NAND U6972 ( .A(\stack[0][17] ), .B(n3339), .Z(n6931) );
  NAND U6973 ( .A(\stack[1][17] ), .B(n6682), .Z(n6930) );
  AND U6974 ( .A(n6932), .B(n6933), .Z(n3026) );
  NAND U6975 ( .A(\stack[0][17] ), .B(n6682), .Z(n6933) );
  NAND U6976 ( .A(\stack[0][17] ), .B(n6683), .Z(n6932) );
  IV U6977 ( .A(n6736), .Z(n3047) );
  XOR U6978 ( .A(n6684), .B(n6934), .Z(n6736) );
  NAND U6979 ( .A(n6935), .B(n6936), .Z(n6934) );
  NAND U6980 ( .A(\stack[1][18] ), .B(n6683), .Z(n6936) );
  AND U6981 ( .A(n6937), .B(n6938), .Z(n6935) );
  NAND U6982 ( .A(\stack[0][18] ), .B(n3339), .Z(n6938) );
  NAND U6983 ( .A(\stack[1][18] ), .B(n6682), .Z(n6937) );
  AND U6984 ( .A(n6939), .B(n6940), .Z(n3050) );
  NAND U6985 ( .A(\stack[0][18] ), .B(n6682), .Z(n6940) );
  NAND U6986 ( .A(\stack[0][18] ), .B(n6683), .Z(n6939) );
  IV U6987 ( .A(n6732), .Z(n3071) );
  XOR U6988 ( .A(n6684), .B(n6941), .Z(n6732) );
  NAND U6989 ( .A(n6942), .B(n6943), .Z(n6941) );
  NAND U6990 ( .A(\stack[1][19] ), .B(n6683), .Z(n6943) );
  AND U6991 ( .A(n6944), .B(n6945), .Z(n6942) );
  NAND U6992 ( .A(\stack[0][19] ), .B(n3339), .Z(n6945) );
  NAND U6993 ( .A(\stack[1][19] ), .B(n6682), .Z(n6944) );
  AND U6994 ( .A(n6946), .B(n6947), .Z(n3074) );
  NAND U6995 ( .A(\stack[0][19] ), .B(n6682), .Z(n6947) );
  NAND U6996 ( .A(\stack[0][19] ), .B(n6683), .Z(n6946) );
  IV U6997 ( .A(n6728), .Z(n3095) );
  XOR U6998 ( .A(n6684), .B(n6948), .Z(n6728) );
  NAND U6999 ( .A(n6949), .B(n6950), .Z(n6948) );
  NAND U7000 ( .A(\stack[1][20] ), .B(n6683), .Z(n6950) );
  AND U7001 ( .A(n6951), .B(n6952), .Z(n6949) );
  NAND U7002 ( .A(\stack[0][20] ), .B(n3339), .Z(n6952) );
  NAND U7003 ( .A(\stack[1][20] ), .B(n6682), .Z(n6951) );
  AND U7004 ( .A(n6953), .B(n6954), .Z(n3098) );
  NAND U7005 ( .A(\stack[0][20] ), .B(n6682), .Z(n6954) );
  NAND U7006 ( .A(\stack[0][20] ), .B(n6683), .Z(n6953) );
  IV U7007 ( .A(n6724), .Z(n3119) );
  XOR U7008 ( .A(n6684), .B(n6955), .Z(n6724) );
  NAND U7009 ( .A(n6956), .B(n6957), .Z(n6955) );
  NAND U7010 ( .A(\stack[1][21] ), .B(n6683), .Z(n6957) );
  AND U7011 ( .A(n6958), .B(n6959), .Z(n6956) );
  NAND U7012 ( .A(\stack[0][21] ), .B(n3339), .Z(n6959) );
  NAND U7013 ( .A(\stack[1][21] ), .B(n6682), .Z(n6958) );
  AND U7014 ( .A(n6960), .B(n6961), .Z(n3122) );
  NAND U7015 ( .A(\stack[0][21] ), .B(n6682), .Z(n6961) );
  NAND U7016 ( .A(\stack[0][21] ), .B(n6683), .Z(n6960) );
  IV U7017 ( .A(n6720), .Z(n3143) );
  XOR U7018 ( .A(n6684), .B(n6962), .Z(n6720) );
  NAND U7019 ( .A(n6963), .B(n6964), .Z(n6962) );
  NAND U7020 ( .A(\stack[1][22] ), .B(n6683), .Z(n6964) );
  AND U7021 ( .A(n6965), .B(n6966), .Z(n6963) );
  NAND U7022 ( .A(\stack[0][22] ), .B(n3339), .Z(n6966) );
  NAND U7023 ( .A(\stack[1][22] ), .B(n6682), .Z(n6965) );
  AND U7024 ( .A(n6967), .B(n6968), .Z(n3146) );
  NAND U7025 ( .A(\stack[0][22] ), .B(n6682), .Z(n6968) );
  NAND U7026 ( .A(\stack[0][22] ), .B(n6683), .Z(n6967) );
  IV U7027 ( .A(n6716), .Z(n3167) );
  XOR U7028 ( .A(n6684), .B(n6969), .Z(n6716) );
  NAND U7029 ( .A(n6970), .B(n6971), .Z(n6969) );
  NAND U7030 ( .A(\stack[1][23] ), .B(n6683), .Z(n6971) );
  AND U7031 ( .A(n6972), .B(n6973), .Z(n6970) );
  NAND U7032 ( .A(\stack[0][23] ), .B(n3339), .Z(n6973) );
  NAND U7033 ( .A(\stack[1][23] ), .B(n6682), .Z(n6972) );
  AND U7034 ( .A(n6974), .B(n6975), .Z(n3170) );
  NAND U7035 ( .A(\stack[0][23] ), .B(n6682), .Z(n6975) );
  NAND U7036 ( .A(\stack[0][23] ), .B(n6683), .Z(n6974) );
  IV U7037 ( .A(n6712), .Z(n3191) );
  XOR U7038 ( .A(n6684), .B(n6976), .Z(n6712) );
  NAND U7039 ( .A(n6977), .B(n6978), .Z(n6976) );
  NAND U7040 ( .A(\stack[1][24] ), .B(n6683), .Z(n6978) );
  AND U7041 ( .A(n6979), .B(n6980), .Z(n6977) );
  NAND U7042 ( .A(\stack[0][24] ), .B(n3339), .Z(n6980) );
  NAND U7043 ( .A(\stack[1][24] ), .B(n6682), .Z(n6979) );
  AND U7044 ( .A(n6981), .B(n6982), .Z(n3194) );
  NAND U7045 ( .A(\stack[0][24] ), .B(n6682), .Z(n6982) );
  NAND U7046 ( .A(\stack[0][24] ), .B(n6683), .Z(n6981) );
  IV U7047 ( .A(n6708), .Z(n3215) );
  XOR U7048 ( .A(n6684), .B(n6983), .Z(n6708) );
  NAND U7049 ( .A(n6984), .B(n6985), .Z(n6983) );
  NAND U7050 ( .A(\stack[1][25] ), .B(n6683), .Z(n6985) );
  AND U7051 ( .A(n6986), .B(n6987), .Z(n6984) );
  NAND U7052 ( .A(\stack[0][25] ), .B(n3339), .Z(n6987) );
  NAND U7053 ( .A(\stack[1][25] ), .B(n6682), .Z(n6986) );
  AND U7054 ( .A(n6988), .B(n6989), .Z(n3218) );
  NAND U7055 ( .A(\stack[0][25] ), .B(n6682), .Z(n6989) );
  NAND U7056 ( .A(\stack[0][25] ), .B(n6683), .Z(n6988) );
  IV U7057 ( .A(n6704), .Z(n3239) );
  XOR U7058 ( .A(n6684), .B(n6990), .Z(n6704) );
  NAND U7059 ( .A(n6991), .B(n6992), .Z(n6990) );
  NAND U7060 ( .A(\stack[1][26] ), .B(n6683), .Z(n6992) );
  AND U7061 ( .A(n6993), .B(n6994), .Z(n6991) );
  NAND U7062 ( .A(\stack[0][26] ), .B(n3339), .Z(n6994) );
  NAND U7063 ( .A(\stack[1][26] ), .B(n6682), .Z(n6993) );
  AND U7064 ( .A(n6995), .B(n6996), .Z(n3242) );
  NAND U7065 ( .A(\stack[0][26] ), .B(n6682), .Z(n6996) );
  NAND U7066 ( .A(\stack[0][26] ), .B(n6683), .Z(n6995) );
  IV U7067 ( .A(n6700), .Z(n3263) );
  XOR U7068 ( .A(n6684), .B(n6997), .Z(n6700) );
  NAND U7069 ( .A(n6998), .B(n6999), .Z(n6997) );
  NAND U7070 ( .A(\stack[1][27] ), .B(n6683), .Z(n6999) );
  AND U7071 ( .A(n7000), .B(n7001), .Z(n6998) );
  NAND U7072 ( .A(\stack[0][27] ), .B(n3339), .Z(n7001) );
  NAND U7073 ( .A(\stack[1][27] ), .B(n6682), .Z(n7000) );
  AND U7074 ( .A(n7002), .B(n7003), .Z(n3266) );
  NAND U7075 ( .A(\stack[0][27] ), .B(n6682), .Z(n7003) );
  NAND U7076 ( .A(\stack[0][27] ), .B(n6683), .Z(n7002) );
  IV U7077 ( .A(n6696), .Z(n3286) );
  XOR U7078 ( .A(n6684), .B(n7004), .Z(n6696) );
  NAND U7079 ( .A(n7005), .B(n7006), .Z(n7004) );
  NAND U7080 ( .A(\stack[1][28] ), .B(n6683), .Z(n7006) );
  AND U7081 ( .A(n7007), .B(n7008), .Z(n7005) );
  NAND U7082 ( .A(\stack[0][28] ), .B(n3339), .Z(n7008) );
  NAND U7083 ( .A(\stack[1][28] ), .B(n6682), .Z(n7007) );
  AND U7084 ( .A(n7009), .B(n7010), .Z(n3289) );
  NAND U7085 ( .A(\stack[0][28] ), .B(n6682), .Z(n7010) );
  NAND U7086 ( .A(\stack[0][28] ), .B(n6683), .Z(n7009) );
  IV U7087 ( .A(n6692), .Z(n3309) );
  XOR U7088 ( .A(n6684), .B(n7011), .Z(n6692) );
  NAND U7089 ( .A(n7012), .B(n7013), .Z(n7011) );
  NAND U7090 ( .A(\stack[1][29] ), .B(n6683), .Z(n7013) );
  AND U7091 ( .A(n7014), .B(n7015), .Z(n7012) );
  NAND U7092 ( .A(\stack[0][29] ), .B(n3339), .Z(n7015) );
  NAND U7093 ( .A(\stack[1][29] ), .B(n6682), .Z(n7014) );
  IV U7094 ( .A(n2621), .Z(n6684) );
  AND U7095 ( .A(n7016), .B(n7017), .Z(n3312) );
  NAND U7096 ( .A(\stack[0][29] ), .B(n6682), .Z(n7017) );
  NAND U7097 ( .A(\stack[0][29] ), .B(n6683), .Z(n7016) );
  AND U7098 ( .A(n7018), .B(n7019), .Z(n6675) );
  NAND U7099 ( .A(\stack[0][31] ), .B(n6682), .Z(n7019) );
  NAND U7100 ( .A(\stack[0][31] ), .B(n6683), .Z(n7018) );
  XOR U7101 ( .A(n2621), .B(n7020), .Z(n6673) );
  AND U7102 ( .A(n7021), .B(n7022), .Z(n7020) );
  NAND U7103 ( .A(\stack[1][31] ), .B(n6683), .Z(n7022) );
  AND U7104 ( .A(n7023), .B(n7024), .Z(n7021) );
  NAND U7105 ( .A(\stack[0][31] ), .B(n3339), .Z(n7024) );
  NAND U7106 ( .A(\stack[1][31] ), .B(n6682), .Z(n7023) );
  NOR U7107 ( .A(n3339), .B(n6683), .Z(n2621) );
  ANDN U7108 ( .B(n7025), .A(n6667), .Z(n3339) );
  AND U7109 ( .A(n6672), .B(opcode[2]), .Z(n7025) );
  NAND U7110 ( .A(n7026), .B(n7027), .Z(n2467) );
  NAND U7111 ( .A(\stack[1][0] ), .B(n7028), .Z(n7027) );
  NAND U7112 ( .A(n7029), .B(n7030), .Z(n7026) );
  NAND U7113 ( .A(n7031), .B(n7032), .Z(n7030) );
  NAND U7114 ( .A(n2503), .B(\stack[2][0] ), .Z(n7032) );
  NAND U7115 ( .A(\stack[0][0] ), .B(n7033), .Z(n7031) );
  NAND U7116 ( .A(n7034), .B(n7035), .Z(n2466) );
  NAND U7117 ( .A(\stack[1][1] ), .B(n7028), .Z(n7035) );
  NAND U7118 ( .A(n7029), .B(n7036), .Z(n7034) );
  NAND U7119 ( .A(n7037), .B(n7038), .Z(n7036) );
  NAND U7120 ( .A(n2503), .B(\stack[2][1] ), .Z(n7038) );
  NAND U7121 ( .A(n7033), .B(\stack[0][1] ), .Z(n7037) );
  NAND U7122 ( .A(n7039), .B(n7040), .Z(n2465) );
  NAND U7123 ( .A(\stack[1][2] ), .B(n7028), .Z(n7040) );
  NAND U7124 ( .A(n7029), .B(n7041), .Z(n7039) );
  NAND U7125 ( .A(n7042), .B(n7043), .Z(n7041) );
  NAND U7126 ( .A(n2503), .B(\stack[2][2] ), .Z(n7043) );
  NAND U7127 ( .A(\stack[0][2] ), .B(n7033), .Z(n7042) );
  NAND U7128 ( .A(n7044), .B(n7045), .Z(n2464) );
  NAND U7129 ( .A(\stack[1][3] ), .B(n7028), .Z(n7045) );
  NAND U7130 ( .A(n7029), .B(n7046), .Z(n7044) );
  NAND U7131 ( .A(n7047), .B(n7048), .Z(n7046) );
  NAND U7132 ( .A(n2503), .B(\stack[2][3] ), .Z(n7048) );
  NAND U7133 ( .A(\stack[0][3] ), .B(n7033), .Z(n7047) );
  NAND U7134 ( .A(n7049), .B(n7050), .Z(n2463) );
  NAND U7135 ( .A(\stack[1][4] ), .B(n7028), .Z(n7050) );
  NAND U7136 ( .A(n7029), .B(n7051), .Z(n7049) );
  NAND U7137 ( .A(n7052), .B(n7053), .Z(n7051) );
  NAND U7138 ( .A(n2503), .B(\stack[2][4] ), .Z(n7053) );
  NAND U7139 ( .A(\stack[0][4] ), .B(n7033), .Z(n7052) );
  NAND U7140 ( .A(n7054), .B(n7055), .Z(n2462) );
  NAND U7141 ( .A(\stack[1][5] ), .B(n7028), .Z(n7055) );
  NAND U7142 ( .A(n7029), .B(n7056), .Z(n7054) );
  NAND U7143 ( .A(n7057), .B(n7058), .Z(n7056) );
  NAND U7144 ( .A(n2503), .B(\stack[2][5] ), .Z(n7058) );
  NAND U7145 ( .A(\stack[0][5] ), .B(n7033), .Z(n7057) );
  NAND U7146 ( .A(n7059), .B(n7060), .Z(n2461) );
  NAND U7147 ( .A(\stack[1][6] ), .B(n7028), .Z(n7060) );
  NAND U7148 ( .A(n7029), .B(n7061), .Z(n7059) );
  NAND U7149 ( .A(n7062), .B(n7063), .Z(n7061) );
  NAND U7150 ( .A(n2503), .B(\stack[2][6] ), .Z(n7063) );
  NAND U7151 ( .A(\stack[0][6] ), .B(n7033), .Z(n7062) );
  NAND U7152 ( .A(n7064), .B(n7065), .Z(n2460) );
  NAND U7153 ( .A(\stack[1][7] ), .B(n7028), .Z(n7065) );
  NAND U7154 ( .A(n7029), .B(n7066), .Z(n7064) );
  NAND U7155 ( .A(n7067), .B(n7068), .Z(n7066) );
  NAND U7156 ( .A(n2503), .B(\stack[2][7] ), .Z(n7068) );
  NAND U7157 ( .A(\stack[0][7] ), .B(n7033), .Z(n7067) );
  NAND U7158 ( .A(n7069), .B(n7070), .Z(n2459) );
  NAND U7159 ( .A(\stack[1][8] ), .B(n7028), .Z(n7070) );
  NAND U7160 ( .A(n7029), .B(n7071), .Z(n7069) );
  NAND U7161 ( .A(n7072), .B(n7073), .Z(n7071) );
  NAND U7162 ( .A(n2503), .B(\stack[2][8] ), .Z(n7073) );
  NAND U7163 ( .A(\stack[0][8] ), .B(n7033), .Z(n7072) );
  NAND U7164 ( .A(n7074), .B(n7075), .Z(n2458) );
  NAND U7165 ( .A(\stack[1][9] ), .B(n7028), .Z(n7075) );
  NAND U7166 ( .A(n7029), .B(n7076), .Z(n7074) );
  NAND U7167 ( .A(n7077), .B(n7078), .Z(n7076) );
  NAND U7168 ( .A(n2503), .B(\stack[2][9] ), .Z(n7078) );
  NAND U7169 ( .A(\stack[0][9] ), .B(n7033), .Z(n7077) );
  NAND U7170 ( .A(n7079), .B(n7080), .Z(n2457) );
  NAND U7171 ( .A(\stack[1][10] ), .B(n7028), .Z(n7080) );
  NAND U7172 ( .A(n7029), .B(n7081), .Z(n7079) );
  NAND U7173 ( .A(n7082), .B(n7083), .Z(n7081) );
  NAND U7174 ( .A(n2503), .B(\stack[2][10] ), .Z(n7083) );
  NAND U7175 ( .A(n7033), .B(\stack[0][10] ), .Z(n7082) );
  NAND U7176 ( .A(n7084), .B(n7085), .Z(n2456) );
  NAND U7177 ( .A(\stack[1][11] ), .B(n7028), .Z(n7085) );
  NAND U7178 ( .A(n7029), .B(n7086), .Z(n7084) );
  NAND U7179 ( .A(n7087), .B(n7088), .Z(n7086) );
  NAND U7180 ( .A(n2503), .B(\stack[2][11] ), .Z(n7088) );
  NAND U7181 ( .A(n7033), .B(\stack[0][11] ), .Z(n7087) );
  NAND U7182 ( .A(n7089), .B(n7090), .Z(n2455) );
  NAND U7183 ( .A(\stack[1][12] ), .B(n7028), .Z(n7090) );
  NAND U7184 ( .A(n7029), .B(n7091), .Z(n7089) );
  NAND U7185 ( .A(n7092), .B(n7093), .Z(n7091) );
  NAND U7186 ( .A(n2503), .B(\stack[2][12] ), .Z(n7093) );
  NAND U7187 ( .A(n7033), .B(\stack[0][12] ), .Z(n7092) );
  NAND U7188 ( .A(n7094), .B(n7095), .Z(n2454) );
  NAND U7189 ( .A(\stack[1][13] ), .B(n7028), .Z(n7095) );
  NAND U7190 ( .A(n7029), .B(n7096), .Z(n7094) );
  NAND U7191 ( .A(n7097), .B(n7098), .Z(n7096) );
  NAND U7192 ( .A(n2503), .B(\stack[2][13] ), .Z(n7098) );
  NAND U7193 ( .A(n7033), .B(\stack[0][13] ), .Z(n7097) );
  NAND U7194 ( .A(n7099), .B(n7100), .Z(n2453) );
  NAND U7195 ( .A(\stack[1][14] ), .B(n7028), .Z(n7100) );
  NAND U7196 ( .A(n7029), .B(n7101), .Z(n7099) );
  NAND U7197 ( .A(n7102), .B(n7103), .Z(n7101) );
  NAND U7198 ( .A(n2503), .B(\stack[2][14] ), .Z(n7103) );
  NAND U7199 ( .A(n7033), .B(\stack[0][14] ), .Z(n7102) );
  NAND U7200 ( .A(n7104), .B(n7105), .Z(n2452) );
  NAND U7201 ( .A(\stack[1][15] ), .B(n7028), .Z(n7105) );
  NAND U7202 ( .A(n7029), .B(n7106), .Z(n7104) );
  NAND U7203 ( .A(n7107), .B(n7108), .Z(n7106) );
  NAND U7204 ( .A(n2503), .B(\stack[2][15] ), .Z(n7108) );
  NAND U7205 ( .A(n7033), .B(\stack[0][15] ), .Z(n7107) );
  NAND U7206 ( .A(n7109), .B(n7110), .Z(n2451) );
  NAND U7207 ( .A(\stack[1][16] ), .B(n7028), .Z(n7110) );
  NAND U7208 ( .A(n7029), .B(n7111), .Z(n7109) );
  NAND U7209 ( .A(n7112), .B(n7113), .Z(n7111) );
  NAND U7210 ( .A(n2503), .B(\stack[2][16] ), .Z(n7113) );
  NAND U7211 ( .A(n7033), .B(\stack[0][16] ), .Z(n7112) );
  NAND U7212 ( .A(n7114), .B(n7115), .Z(n2450) );
  NAND U7213 ( .A(\stack[1][17] ), .B(n7028), .Z(n7115) );
  NAND U7214 ( .A(n7029), .B(n7116), .Z(n7114) );
  NAND U7215 ( .A(n7117), .B(n7118), .Z(n7116) );
  NAND U7216 ( .A(n2503), .B(\stack[2][17] ), .Z(n7118) );
  NAND U7217 ( .A(n7033), .B(\stack[0][17] ), .Z(n7117) );
  NAND U7218 ( .A(n7119), .B(n7120), .Z(n2449) );
  NAND U7219 ( .A(\stack[1][18] ), .B(n7028), .Z(n7120) );
  NAND U7220 ( .A(n7029), .B(n7121), .Z(n7119) );
  NAND U7221 ( .A(n7122), .B(n7123), .Z(n7121) );
  NAND U7222 ( .A(n2503), .B(\stack[2][18] ), .Z(n7123) );
  NAND U7223 ( .A(n7033), .B(\stack[0][18] ), .Z(n7122) );
  NAND U7224 ( .A(n7124), .B(n7125), .Z(n2448) );
  NAND U7225 ( .A(\stack[1][19] ), .B(n7028), .Z(n7125) );
  NAND U7226 ( .A(n7029), .B(n7126), .Z(n7124) );
  NAND U7227 ( .A(n7127), .B(n7128), .Z(n7126) );
  NAND U7228 ( .A(n2503), .B(\stack[2][19] ), .Z(n7128) );
  NAND U7229 ( .A(n7033), .B(\stack[0][19] ), .Z(n7127) );
  NAND U7230 ( .A(n7129), .B(n7130), .Z(n2447) );
  NAND U7231 ( .A(\stack[1][20] ), .B(n7028), .Z(n7130) );
  NAND U7232 ( .A(n7029), .B(n7131), .Z(n7129) );
  NAND U7233 ( .A(n7132), .B(n7133), .Z(n7131) );
  NAND U7234 ( .A(n2503), .B(\stack[2][20] ), .Z(n7133) );
  NAND U7235 ( .A(n7033), .B(\stack[0][20] ), .Z(n7132) );
  NAND U7236 ( .A(n7134), .B(n7135), .Z(n2446) );
  NAND U7237 ( .A(\stack[1][21] ), .B(n7028), .Z(n7135) );
  NAND U7238 ( .A(n7029), .B(n7136), .Z(n7134) );
  NAND U7239 ( .A(n7137), .B(n7138), .Z(n7136) );
  NAND U7240 ( .A(n2503), .B(\stack[2][21] ), .Z(n7138) );
  NAND U7241 ( .A(n7033), .B(\stack[0][21] ), .Z(n7137) );
  NAND U7242 ( .A(n7139), .B(n7140), .Z(n2445) );
  NAND U7243 ( .A(\stack[1][22] ), .B(n7028), .Z(n7140) );
  NAND U7244 ( .A(n7029), .B(n7141), .Z(n7139) );
  NAND U7245 ( .A(n7142), .B(n7143), .Z(n7141) );
  NAND U7246 ( .A(n2503), .B(\stack[2][22] ), .Z(n7143) );
  NAND U7247 ( .A(n7033), .B(\stack[0][22] ), .Z(n7142) );
  NAND U7248 ( .A(n7144), .B(n7145), .Z(n2444) );
  NAND U7249 ( .A(\stack[1][23] ), .B(n7028), .Z(n7145) );
  NAND U7250 ( .A(n7029), .B(n7146), .Z(n7144) );
  NAND U7251 ( .A(n7147), .B(n7148), .Z(n7146) );
  NAND U7252 ( .A(n2503), .B(\stack[2][23] ), .Z(n7148) );
  NAND U7253 ( .A(n7033), .B(\stack[0][23] ), .Z(n7147) );
  NAND U7254 ( .A(n7149), .B(n7150), .Z(n2443) );
  NAND U7255 ( .A(\stack[1][24] ), .B(n7028), .Z(n7150) );
  NAND U7256 ( .A(n7029), .B(n7151), .Z(n7149) );
  NAND U7257 ( .A(n7152), .B(n7153), .Z(n7151) );
  NAND U7258 ( .A(n2503), .B(\stack[2][24] ), .Z(n7153) );
  NAND U7259 ( .A(n7033), .B(\stack[0][24] ), .Z(n7152) );
  NAND U7260 ( .A(n7154), .B(n7155), .Z(n2442) );
  NAND U7261 ( .A(\stack[1][25] ), .B(n7028), .Z(n7155) );
  NAND U7262 ( .A(n7029), .B(n7156), .Z(n7154) );
  NAND U7263 ( .A(n7157), .B(n7158), .Z(n7156) );
  NAND U7264 ( .A(n2503), .B(\stack[2][25] ), .Z(n7158) );
  NAND U7265 ( .A(n7033), .B(\stack[0][25] ), .Z(n7157) );
  NAND U7266 ( .A(n7159), .B(n7160), .Z(n2441) );
  NAND U7267 ( .A(\stack[1][26] ), .B(n7028), .Z(n7160) );
  NAND U7268 ( .A(n7029), .B(n7161), .Z(n7159) );
  NAND U7269 ( .A(n7162), .B(n7163), .Z(n7161) );
  NAND U7270 ( .A(n2503), .B(\stack[2][26] ), .Z(n7163) );
  NAND U7271 ( .A(n7033), .B(\stack[0][26] ), .Z(n7162) );
  NAND U7272 ( .A(n7164), .B(n7165), .Z(n2440) );
  NAND U7273 ( .A(\stack[1][27] ), .B(n7028), .Z(n7165) );
  NAND U7274 ( .A(n7029), .B(n7166), .Z(n7164) );
  NAND U7275 ( .A(n7167), .B(n7168), .Z(n7166) );
  NAND U7276 ( .A(n2503), .B(\stack[2][27] ), .Z(n7168) );
  NAND U7277 ( .A(n7033), .B(\stack[0][27] ), .Z(n7167) );
  NAND U7278 ( .A(n7169), .B(n7170), .Z(n2439) );
  NAND U7279 ( .A(\stack[1][28] ), .B(n7028), .Z(n7170) );
  NAND U7280 ( .A(n7029), .B(n7171), .Z(n7169) );
  NAND U7281 ( .A(n7172), .B(n7173), .Z(n7171) );
  NAND U7282 ( .A(n2503), .B(\stack[2][28] ), .Z(n7173) );
  NAND U7283 ( .A(n7033), .B(\stack[0][28] ), .Z(n7172) );
  NAND U7284 ( .A(n7174), .B(n7175), .Z(n2438) );
  NAND U7285 ( .A(\stack[1][29] ), .B(n7028), .Z(n7175) );
  NAND U7286 ( .A(n7029), .B(n7176), .Z(n7174) );
  NAND U7287 ( .A(n7177), .B(n7178), .Z(n7176) );
  NAND U7288 ( .A(n2503), .B(\stack[2][29] ), .Z(n7178) );
  NAND U7289 ( .A(n7033), .B(\stack[0][29] ), .Z(n7177) );
  NAND U7290 ( .A(n7179), .B(n7180), .Z(n2437) );
  NAND U7291 ( .A(\stack[1][30] ), .B(n7028), .Z(n7180) );
  NAND U7292 ( .A(n7029), .B(n7181), .Z(n7179) );
  NAND U7293 ( .A(n7182), .B(n7183), .Z(n7181) );
  NAND U7294 ( .A(n2503), .B(\stack[2][30] ), .Z(n7183) );
  NAND U7295 ( .A(n7033), .B(\stack[0][30] ), .Z(n7182) );
  NAND U7296 ( .A(n7184), .B(n7185), .Z(n2436) );
  NAND U7297 ( .A(\stack[1][31] ), .B(n7028), .Z(n7185) );
  NAND U7298 ( .A(n7029), .B(n7186), .Z(n7184) );
  NAND U7299 ( .A(n7187), .B(n7188), .Z(n7186) );
  NAND U7300 ( .A(n2503), .B(\stack[2][31] ), .Z(n7188) );
  NAND U7301 ( .A(n7033), .B(\stack[0][31] ), .Z(n7187) );
  NAND U7302 ( .A(n7189), .B(n7190), .Z(n2435) );
  NAND U7303 ( .A(n7028), .B(\stack[2][0] ), .Z(n7190) );
  NAND U7304 ( .A(n7029), .B(n7191), .Z(n7189) );
  NAND U7305 ( .A(n7192), .B(n7193), .Z(n7191) );
  NAND U7306 ( .A(n2503), .B(\stack[3][0] ), .Z(n7193) );
  NAND U7307 ( .A(\stack[1][0] ), .B(n7033), .Z(n7192) );
  NAND U7308 ( .A(n7194), .B(n7195), .Z(n2434) );
  NAND U7309 ( .A(n7028), .B(\stack[2][1] ), .Z(n7195) );
  NAND U7310 ( .A(n7029), .B(n7196), .Z(n7194) );
  NAND U7311 ( .A(n7197), .B(n7198), .Z(n7196) );
  NAND U7312 ( .A(n2503), .B(\stack[3][1] ), .Z(n7198) );
  NAND U7313 ( .A(\stack[1][1] ), .B(n7033), .Z(n7197) );
  NAND U7314 ( .A(n7199), .B(n7200), .Z(n2433) );
  NAND U7315 ( .A(n7028), .B(\stack[2][2] ), .Z(n7200) );
  NAND U7316 ( .A(n7029), .B(n7201), .Z(n7199) );
  NAND U7317 ( .A(n7202), .B(n7203), .Z(n7201) );
  NAND U7318 ( .A(n2503), .B(\stack[3][2] ), .Z(n7203) );
  NAND U7319 ( .A(\stack[1][2] ), .B(n7033), .Z(n7202) );
  NAND U7320 ( .A(n7204), .B(n7205), .Z(n2432) );
  NAND U7321 ( .A(n7028), .B(\stack[2][3] ), .Z(n7205) );
  NAND U7322 ( .A(n7029), .B(n7206), .Z(n7204) );
  NAND U7323 ( .A(n7207), .B(n7208), .Z(n7206) );
  NAND U7324 ( .A(n2503), .B(\stack[3][3] ), .Z(n7208) );
  NAND U7325 ( .A(\stack[1][3] ), .B(n7033), .Z(n7207) );
  NAND U7326 ( .A(n7209), .B(n7210), .Z(n2431) );
  NAND U7327 ( .A(n7028), .B(\stack[2][4] ), .Z(n7210) );
  NAND U7328 ( .A(n7029), .B(n7211), .Z(n7209) );
  NAND U7329 ( .A(n7212), .B(n7213), .Z(n7211) );
  NAND U7330 ( .A(n2503), .B(\stack[3][4] ), .Z(n7213) );
  NAND U7331 ( .A(\stack[1][4] ), .B(n7033), .Z(n7212) );
  NAND U7332 ( .A(n7214), .B(n7215), .Z(n2430) );
  NAND U7333 ( .A(n7028), .B(\stack[2][5] ), .Z(n7215) );
  NAND U7334 ( .A(n7029), .B(n7216), .Z(n7214) );
  NAND U7335 ( .A(n7217), .B(n7218), .Z(n7216) );
  NAND U7336 ( .A(n2503), .B(\stack[3][5] ), .Z(n7218) );
  NAND U7337 ( .A(\stack[1][5] ), .B(n7033), .Z(n7217) );
  NAND U7338 ( .A(n7219), .B(n7220), .Z(n2429) );
  NAND U7339 ( .A(n7028), .B(\stack[2][6] ), .Z(n7220) );
  NAND U7340 ( .A(n7029), .B(n7221), .Z(n7219) );
  NAND U7341 ( .A(n7222), .B(n7223), .Z(n7221) );
  NAND U7342 ( .A(n2503), .B(\stack[3][6] ), .Z(n7223) );
  NAND U7343 ( .A(\stack[1][6] ), .B(n7033), .Z(n7222) );
  NAND U7344 ( .A(n7224), .B(n7225), .Z(n2428) );
  NAND U7345 ( .A(n7028), .B(\stack[2][7] ), .Z(n7225) );
  NAND U7346 ( .A(n7029), .B(n7226), .Z(n7224) );
  NAND U7347 ( .A(n7227), .B(n7228), .Z(n7226) );
  NAND U7348 ( .A(n2503), .B(\stack[3][7] ), .Z(n7228) );
  NAND U7349 ( .A(\stack[1][7] ), .B(n7033), .Z(n7227) );
  NAND U7350 ( .A(n7229), .B(n7230), .Z(n2427) );
  NAND U7351 ( .A(n7028), .B(\stack[2][8] ), .Z(n7230) );
  NAND U7352 ( .A(n7029), .B(n7231), .Z(n7229) );
  NAND U7353 ( .A(n7232), .B(n7233), .Z(n7231) );
  NAND U7354 ( .A(n2503), .B(\stack[3][8] ), .Z(n7233) );
  NAND U7355 ( .A(\stack[1][8] ), .B(n7033), .Z(n7232) );
  NAND U7356 ( .A(n7234), .B(n7235), .Z(n2426) );
  NAND U7357 ( .A(n7028), .B(\stack[2][9] ), .Z(n7235) );
  NAND U7358 ( .A(n7029), .B(n7236), .Z(n7234) );
  NAND U7359 ( .A(n7237), .B(n7238), .Z(n7236) );
  NAND U7360 ( .A(n2503), .B(\stack[3][9] ), .Z(n7238) );
  NAND U7361 ( .A(\stack[1][9] ), .B(n7033), .Z(n7237) );
  NAND U7362 ( .A(n7239), .B(n7240), .Z(n2425) );
  NAND U7363 ( .A(n7028), .B(\stack[2][10] ), .Z(n7240) );
  NAND U7364 ( .A(n7029), .B(n7241), .Z(n7239) );
  NAND U7365 ( .A(n7242), .B(n7243), .Z(n7241) );
  NAND U7366 ( .A(n2503), .B(\stack[3][10] ), .Z(n7243) );
  NAND U7367 ( .A(n7033), .B(\stack[1][10] ), .Z(n7242) );
  NAND U7368 ( .A(n7244), .B(n7245), .Z(n2424) );
  NAND U7369 ( .A(n7028), .B(\stack[2][11] ), .Z(n7245) );
  NAND U7370 ( .A(n7029), .B(n7246), .Z(n7244) );
  NAND U7371 ( .A(n7247), .B(n7248), .Z(n7246) );
  NAND U7372 ( .A(n2503), .B(\stack[3][11] ), .Z(n7248) );
  NAND U7373 ( .A(n7033), .B(\stack[1][11] ), .Z(n7247) );
  NAND U7374 ( .A(n7249), .B(n7250), .Z(n2423) );
  NAND U7375 ( .A(n7028), .B(\stack[2][12] ), .Z(n7250) );
  NAND U7376 ( .A(n7029), .B(n7251), .Z(n7249) );
  NAND U7377 ( .A(n7252), .B(n7253), .Z(n7251) );
  NAND U7378 ( .A(n2503), .B(\stack[3][12] ), .Z(n7253) );
  NAND U7379 ( .A(n7033), .B(\stack[1][12] ), .Z(n7252) );
  NAND U7380 ( .A(n7254), .B(n7255), .Z(n2422) );
  NAND U7381 ( .A(n7028), .B(\stack[2][13] ), .Z(n7255) );
  NAND U7382 ( .A(n7029), .B(n7256), .Z(n7254) );
  NAND U7383 ( .A(n7257), .B(n7258), .Z(n7256) );
  NAND U7384 ( .A(n2503), .B(\stack[3][13] ), .Z(n7258) );
  NAND U7385 ( .A(n7033), .B(\stack[1][13] ), .Z(n7257) );
  NAND U7386 ( .A(n7259), .B(n7260), .Z(n2421) );
  NAND U7387 ( .A(n7028), .B(\stack[2][14] ), .Z(n7260) );
  NAND U7388 ( .A(n7029), .B(n7261), .Z(n7259) );
  NAND U7389 ( .A(n7262), .B(n7263), .Z(n7261) );
  NAND U7390 ( .A(n2503), .B(\stack[3][14] ), .Z(n7263) );
  NAND U7391 ( .A(n7033), .B(\stack[1][14] ), .Z(n7262) );
  NAND U7392 ( .A(n7264), .B(n7265), .Z(n2420) );
  NAND U7393 ( .A(n7028), .B(\stack[2][15] ), .Z(n7265) );
  NAND U7394 ( .A(n7029), .B(n7266), .Z(n7264) );
  NAND U7395 ( .A(n7267), .B(n7268), .Z(n7266) );
  NAND U7396 ( .A(n2503), .B(\stack[3][15] ), .Z(n7268) );
  NAND U7397 ( .A(n7033), .B(\stack[1][15] ), .Z(n7267) );
  NAND U7398 ( .A(n7269), .B(n7270), .Z(n2419) );
  NAND U7399 ( .A(n7028), .B(\stack[2][16] ), .Z(n7270) );
  NAND U7400 ( .A(n7029), .B(n7271), .Z(n7269) );
  NAND U7401 ( .A(n7272), .B(n7273), .Z(n7271) );
  NAND U7402 ( .A(n2503), .B(\stack[3][16] ), .Z(n7273) );
  NAND U7403 ( .A(n7033), .B(\stack[1][16] ), .Z(n7272) );
  NAND U7404 ( .A(n7274), .B(n7275), .Z(n2418) );
  NAND U7405 ( .A(n7028), .B(\stack[2][17] ), .Z(n7275) );
  NAND U7406 ( .A(n7029), .B(n7276), .Z(n7274) );
  NAND U7407 ( .A(n7277), .B(n7278), .Z(n7276) );
  NAND U7408 ( .A(n2503), .B(\stack[3][17] ), .Z(n7278) );
  NAND U7409 ( .A(n7033), .B(\stack[1][17] ), .Z(n7277) );
  NAND U7410 ( .A(n7279), .B(n7280), .Z(n2417) );
  NAND U7411 ( .A(n7028), .B(\stack[2][18] ), .Z(n7280) );
  NAND U7412 ( .A(n7029), .B(n7281), .Z(n7279) );
  NAND U7413 ( .A(n7282), .B(n7283), .Z(n7281) );
  NAND U7414 ( .A(n2503), .B(\stack[3][18] ), .Z(n7283) );
  NAND U7415 ( .A(n7033), .B(\stack[1][18] ), .Z(n7282) );
  NAND U7416 ( .A(n7284), .B(n7285), .Z(n2416) );
  NAND U7417 ( .A(n7028), .B(\stack[2][19] ), .Z(n7285) );
  NAND U7418 ( .A(n7029), .B(n7286), .Z(n7284) );
  NAND U7419 ( .A(n7287), .B(n7288), .Z(n7286) );
  NAND U7420 ( .A(n2503), .B(\stack[3][19] ), .Z(n7288) );
  NAND U7421 ( .A(n7033), .B(\stack[1][19] ), .Z(n7287) );
  NAND U7422 ( .A(n7289), .B(n7290), .Z(n2415) );
  NAND U7423 ( .A(n7028), .B(\stack[2][20] ), .Z(n7290) );
  NAND U7424 ( .A(n7029), .B(n7291), .Z(n7289) );
  NAND U7425 ( .A(n7292), .B(n7293), .Z(n7291) );
  NAND U7426 ( .A(n2503), .B(\stack[3][20] ), .Z(n7293) );
  NAND U7427 ( .A(n7033), .B(\stack[1][20] ), .Z(n7292) );
  NAND U7428 ( .A(n7294), .B(n7295), .Z(n2414) );
  NAND U7429 ( .A(n7028), .B(\stack[2][21] ), .Z(n7295) );
  NAND U7430 ( .A(n7029), .B(n7296), .Z(n7294) );
  NAND U7431 ( .A(n7297), .B(n7298), .Z(n7296) );
  NAND U7432 ( .A(n2503), .B(\stack[3][21] ), .Z(n7298) );
  NAND U7433 ( .A(n7033), .B(\stack[1][21] ), .Z(n7297) );
  NAND U7434 ( .A(n7299), .B(n7300), .Z(n2413) );
  NAND U7435 ( .A(n7028), .B(\stack[2][22] ), .Z(n7300) );
  NAND U7436 ( .A(n7029), .B(n7301), .Z(n7299) );
  NAND U7437 ( .A(n7302), .B(n7303), .Z(n7301) );
  NAND U7438 ( .A(n2503), .B(\stack[3][22] ), .Z(n7303) );
  NAND U7439 ( .A(n7033), .B(\stack[1][22] ), .Z(n7302) );
  NAND U7440 ( .A(n7304), .B(n7305), .Z(n2412) );
  NAND U7441 ( .A(n7028), .B(\stack[2][23] ), .Z(n7305) );
  NAND U7442 ( .A(n7029), .B(n7306), .Z(n7304) );
  NAND U7443 ( .A(n7307), .B(n7308), .Z(n7306) );
  NAND U7444 ( .A(n2503), .B(\stack[3][23] ), .Z(n7308) );
  NAND U7445 ( .A(n7033), .B(\stack[1][23] ), .Z(n7307) );
  NAND U7446 ( .A(n7309), .B(n7310), .Z(n2411) );
  NAND U7447 ( .A(n7028), .B(\stack[2][24] ), .Z(n7310) );
  NAND U7448 ( .A(n7029), .B(n7311), .Z(n7309) );
  NAND U7449 ( .A(n7312), .B(n7313), .Z(n7311) );
  NAND U7450 ( .A(n2503), .B(\stack[3][24] ), .Z(n7313) );
  NAND U7451 ( .A(n7033), .B(\stack[1][24] ), .Z(n7312) );
  NAND U7452 ( .A(n7314), .B(n7315), .Z(n2410) );
  NAND U7453 ( .A(n7028), .B(\stack[2][25] ), .Z(n7315) );
  NAND U7454 ( .A(n7029), .B(n7316), .Z(n7314) );
  NAND U7455 ( .A(n7317), .B(n7318), .Z(n7316) );
  NAND U7456 ( .A(n2503), .B(\stack[3][25] ), .Z(n7318) );
  NAND U7457 ( .A(n7033), .B(\stack[1][25] ), .Z(n7317) );
  NAND U7458 ( .A(n7319), .B(n7320), .Z(n2409) );
  NAND U7459 ( .A(n7028), .B(\stack[2][26] ), .Z(n7320) );
  NAND U7460 ( .A(n7029), .B(n7321), .Z(n7319) );
  NAND U7461 ( .A(n7322), .B(n7323), .Z(n7321) );
  NAND U7462 ( .A(n2503), .B(\stack[3][26] ), .Z(n7323) );
  NAND U7463 ( .A(n7033), .B(\stack[1][26] ), .Z(n7322) );
  NAND U7464 ( .A(n7324), .B(n7325), .Z(n2408) );
  NAND U7465 ( .A(n7028), .B(\stack[2][27] ), .Z(n7325) );
  NAND U7466 ( .A(n7029), .B(n7326), .Z(n7324) );
  NAND U7467 ( .A(n7327), .B(n7328), .Z(n7326) );
  NAND U7468 ( .A(n2503), .B(\stack[3][27] ), .Z(n7328) );
  NAND U7469 ( .A(n7033), .B(\stack[1][27] ), .Z(n7327) );
  NAND U7470 ( .A(n7329), .B(n7330), .Z(n2407) );
  NAND U7471 ( .A(n7028), .B(\stack[2][28] ), .Z(n7330) );
  NAND U7472 ( .A(n7029), .B(n7331), .Z(n7329) );
  NAND U7473 ( .A(n7332), .B(n7333), .Z(n7331) );
  NAND U7474 ( .A(n2503), .B(\stack[3][28] ), .Z(n7333) );
  NAND U7475 ( .A(n7033), .B(\stack[1][28] ), .Z(n7332) );
  NAND U7476 ( .A(n7334), .B(n7335), .Z(n2406) );
  NAND U7477 ( .A(n7028), .B(\stack[2][29] ), .Z(n7335) );
  NAND U7478 ( .A(n7029), .B(n7336), .Z(n7334) );
  NAND U7479 ( .A(n7337), .B(n7338), .Z(n7336) );
  NAND U7480 ( .A(n2503), .B(\stack[3][29] ), .Z(n7338) );
  NAND U7481 ( .A(n7033), .B(\stack[1][29] ), .Z(n7337) );
  NAND U7482 ( .A(n7339), .B(n7340), .Z(n2405) );
  NAND U7483 ( .A(n7028), .B(\stack[2][30] ), .Z(n7340) );
  NAND U7484 ( .A(n7029), .B(n7341), .Z(n7339) );
  NAND U7485 ( .A(n7342), .B(n7343), .Z(n7341) );
  NAND U7486 ( .A(n2503), .B(\stack[3][30] ), .Z(n7343) );
  NAND U7487 ( .A(n7033), .B(\stack[1][30] ), .Z(n7342) );
  NAND U7488 ( .A(n7344), .B(n7345), .Z(n2404) );
  NAND U7489 ( .A(n7028), .B(\stack[2][31] ), .Z(n7345) );
  NAND U7490 ( .A(n7029), .B(n7346), .Z(n7344) );
  NAND U7491 ( .A(n7347), .B(n7348), .Z(n7346) );
  NAND U7492 ( .A(n2503), .B(\stack[3][31] ), .Z(n7348) );
  NAND U7493 ( .A(n7033), .B(\stack[1][31] ), .Z(n7347) );
  NAND U7494 ( .A(n7349), .B(n7350), .Z(n2403) );
  NAND U7495 ( .A(n7028), .B(\stack[3][0] ), .Z(n7350) );
  NAND U7496 ( .A(n7029), .B(n7351), .Z(n7349) );
  NAND U7497 ( .A(n7352), .B(n7353), .Z(n7351) );
  NAND U7498 ( .A(n2503), .B(\stack[4][0] ), .Z(n7353) );
  NAND U7499 ( .A(n7033), .B(\stack[2][0] ), .Z(n7352) );
  NAND U7500 ( .A(n7354), .B(n7355), .Z(n2402) );
  NAND U7501 ( .A(n7028), .B(\stack[3][1] ), .Z(n7355) );
  NAND U7502 ( .A(n7029), .B(n7356), .Z(n7354) );
  NAND U7503 ( .A(n7357), .B(n7358), .Z(n7356) );
  NAND U7504 ( .A(n2503), .B(\stack[4][1] ), .Z(n7358) );
  NAND U7505 ( .A(n7033), .B(\stack[2][1] ), .Z(n7357) );
  NAND U7506 ( .A(n7359), .B(n7360), .Z(n2401) );
  NAND U7507 ( .A(n7028), .B(\stack[3][2] ), .Z(n7360) );
  NAND U7508 ( .A(n7029), .B(n7361), .Z(n7359) );
  NAND U7509 ( .A(n7362), .B(n7363), .Z(n7361) );
  NAND U7510 ( .A(n2503), .B(\stack[4][2] ), .Z(n7363) );
  NAND U7511 ( .A(n7033), .B(\stack[2][2] ), .Z(n7362) );
  NAND U7512 ( .A(n7364), .B(n7365), .Z(n2400) );
  NAND U7513 ( .A(n7028), .B(\stack[3][3] ), .Z(n7365) );
  NAND U7514 ( .A(n7029), .B(n7366), .Z(n7364) );
  NAND U7515 ( .A(n7367), .B(n7368), .Z(n7366) );
  NAND U7516 ( .A(n2503), .B(\stack[4][3] ), .Z(n7368) );
  NAND U7517 ( .A(n7033), .B(\stack[2][3] ), .Z(n7367) );
  NAND U7518 ( .A(n7369), .B(n7370), .Z(n2399) );
  NAND U7519 ( .A(n7028), .B(\stack[3][4] ), .Z(n7370) );
  NAND U7520 ( .A(n7029), .B(n7371), .Z(n7369) );
  NAND U7521 ( .A(n7372), .B(n7373), .Z(n7371) );
  NAND U7522 ( .A(n2503), .B(\stack[4][4] ), .Z(n7373) );
  NAND U7523 ( .A(n7033), .B(\stack[2][4] ), .Z(n7372) );
  NAND U7524 ( .A(n7374), .B(n7375), .Z(n2398) );
  NAND U7525 ( .A(n7028), .B(\stack[3][5] ), .Z(n7375) );
  NAND U7526 ( .A(n7029), .B(n7376), .Z(n7374) );
  NAND U7527 ( .A(n7377), .B(n7378), .Z(n7376) );
  NAND U7528 ( .A(n2503), .B(\stack[4][5] ), .Z(n7378) );
  NAND U7529 ( .A(n7033), .B(\stack[2][5] ), .Z(n7377) );
  NAND U7530 ( .A(n7379), .B(n7380), .Z(n2397) );
  NAND U7531 ( .A(n7028), .B(\stack[3][6] ), .Z(n7380) );
  NAND U7532 ( .A(n7029), .B(n7381), .Z(n7379) );
  NAND U7533 ( .A(n7382), .B(n7383), .Z(n7381) );
  NAND U7534 ( .A(n2503), .B(\stack[4][6] ), .Z(n7383) );
  NAND U7535 ( .A(n7033), .B(\stack[2][6] ), .Z(n7382) );
  NAND U7536 ( .A(n7384), .B(n7385), .Z(n2396) );
  NAND U7537 ( .A(n7028), .B(\stack[3][7] ), .Z(n7385) );
  NAND U7538 ( .A(n7029), .B(n7386), .Z(n7384) );
  NAND U7539 ( .A(n7387), .B(n7388), .Z(n7386) );
  NAND U7540 ( .A(n2503), .B(\stack[4][7] ), .Z(n7388) );
  NAND U7541 ( .A(n7033), .B(\stack[2][7] ), .Z(n7387) );
  NAND U7542 ( .A(n7389), .B(n7390), .Z(n2395) );
  NAND U7543 ( .A(n7028), .B(\stack[3][8] ), .Z(n7390) );
  NAND U7544 ( .A(n7029), .B(n7391), .Z(n7389) );
  NAND U7545 ( .A(n7392), .B(n7393), .Z(n7391) );
  NAND U7546 ( .A(n2503), .B(\stack[4][8] ), .Z(n7393) );
  NAND U7547 ( .A(n7033), .B(\stack[2][8] ), .Z(n7392) );
  NAND U7548 ( .A(n7394), .B(n7395), .Z(n2394) );
  NAND U7549 ( .A(n7028), .B(\stack[3][9] ), .Z(n7395) );
  NAND U7550 ( .A(n7029), .B(n7396), .Z(n7394) );
  NAND U7551 ( .A(n7397), .B(n7398), .Z(n7396) );
  NAND U7552 ( .A(n2503), .B(\stack[4][9] ), .Z(n7398) );
  NAND U7553 ( .A(n7033), .B(\stack[2][9] ), .Z(n7397) );
  NAND U7554 ( .A(n7399), .B(n7400), .Z(n2393) );
  NAND U7555 ( .A(n7028), .B(\stack[3][10] ), .Z(n7400) );
  NAND U7556 ( .A(n7029), .B(n7401), .Z(n7399) );
  NAND U7557 ( .A(n7402), .B(n7403), .Z(n7401) );
  NAND U7558 ( .A(n2503), .B(\stack[4][10] ), .Z(n7403) );
  NAND U7559 ( .A(n7033), .B(\stack[2][10] ), .Z(n7402) );
  NAND U7560 ( .A(n7404), .B(n7405), .Z(n2392) );
  NAND U7561 ( .A(n7028), .B(\stack[3][11] ), .Z(n7405) );
  NAND U7562 ( .A(n7029), .B(n7406), .Z(n7404) );
  NAND U7563 ( .A(n7407), .B(n7408), .Z(n7406) );
  NAND U7564 ( .A(n2503), .B(\stack[4][11] ), .Z(n7408) );
  NAND U7565 ( .A(n7033), .B(\stack[2][11] ), .Z(n7407) );
  NAND U7566 ( .A(n7409), .B(n7410), .Z(n2391) );
  NAND U7567 ( .A(n7028), .B(\stack[3][12] ), .Z(n7410) );
  NAND U7568 ( .A(n7029), .B(n7411), .Z(n7409) );
  NAND U7569 ( .A(n7412), .B(n7413), .Z(n7411) );
  NAND U7570 ( .A(n2503), .B(\stack[4][12] ), .Z(n7413) );
  NAND U7571 ( .A(n7033), .B(\stack[2][12] ), .Z(n7412) );
  NAND U7572 ( .A(n7414), .B(n7415), .Z(n2390) );
  NAND U7573 ( .A(n7028), .B(\stack[3][13] ), .Z(n7415) );
  NAND U7574 ( .A(n7029), .B(n7416), .Z(n7414) );
  NAND U7575 ( .A(n7417), .B(n7418), .Z(n7416) );
  NAND U7576 ( .A(n2503), .B(\stack[4][13] ), .Z(n7418) );
  NAND U7577 ( .A(n7033), .B(\stack[2][13] ), .Z(n7417) );
  NAND U7578 ( .A(n7419), .B(n7420), .Z(n2389) );
  NAND U7579 ( .A(n7028), .B(\stack[3][14] ), .Z(n7420) );
  NAND U7580 ( .A(n7029), .B(n7421), .Z(n7419) );
  NAND U7581 ( .A(n7422), .B(n7423), .Z(n7421) );
  NAND U7582 ( .A(n2503), .B(\stack[4][14] ), .Z(n7423) );
  NAND U7583 ( .A(n7033), .B(\stack[2][14] ), .Z(n7422) );
  NAND U7584 ( .A(n7424), .B(n7425), .Z(n2388) );
  NAND U7585 ( .A(n7028), .B(\stack[3][15] ), .Z(n7425) );
  NAND U7586 ( .A(n7029), .B(n7426), .Z(n7424) );
  NAND U7587 ( .A(n7427), .B(n7428), .Z(n7426) );
  NAND U7588 ( .A(n2503), .B(\stack[4][15] ), .Z(n7428) );
  NAND U7589 ( .A(n7033), .B(\stack[2][15] ), .Z(n7427) );
  NAND U7590 ( .A(n7429), .B(n7430), .Z(n2387) );
  NAND U7591 ( .A(n7028), .B(\stack[3][16] ), .Z(n7430) );
  NAND U7592 ( .A(n7029), .B(n7431), .Z(n7429) );
  NAND U7593 ( .A(n7432), .B(n7433), .Z(n7431) );
  NAND U7594 ( .A(n2503), .B(\stack[4][16] ), .Z(n7433) );
  NAND U7595 ( .A(n7033), .B(\stack[2][16] ), .Z(n7432) );
  NAND U7596 ( .A(n7434), .B(n7435), .Z(n2386) );
  NAND U7597 ( .A(n7028), .B(\stack[3][17] ), .Z(n7435) );
  NAND U7598 ( .A(n7029), .B(n7436), .Z(n7434) );
  NAND U7599 ( .A(n7437), .B(n7438), .Z(n7436) );
  NAND U7600 ( .A(n2503), .B(\stack[4][17] ), .Z(n7438) );
  NAND U7601 ( .A(n7033), .B(\stack[2][17] ), .Z(n7437) );
  NAND U7602 ( .A(n7439), .B(n7440), .Z(n2385) );
  NAND U7603 ( .A(n7028), .B(\stack[3][18] ), .Z(n7440) );
  NAND U7604 ( .A(n7029), .B(n7441), .Z(n7439) );
  NAND U7605 ( .A(n7442), .B(n7443), .Z(n7441) );
  NAND U7606 ( .A(n2503), .B(\stack[4][18] ), .Z(n7443) );
  NAND U7607 ( .A(n7033), .B(\stack[2][18] ), .Z(n7442) );
  NAND U7608 ( .A(n7444), .B(n7445), .Z(n2384) );
  NAND U7609 ( .A(n7028), .B(\stack[3][19] ), .Z(n7445) );
  NAND U7610 ( .A(n7029), .B(n7446), .Z(n7444) );
  NAND U7611 ( .A(n7447), .B(n7448), .Z(n7446) );
  NAND U7612 ( .A(n2503), .B(\stack[4][19] ), .Z(n7448) );
  NAND U7613 ( .A(n7033), .B(\stack[2][19] ), .Z(n7447) );
  NAND U7614 ( .A(n7449), .B(n7450), .Z(n2383) );
  NAND U7615 ( .A(n7028), .B(\stack[3][20] ), .Z(n7450) );
  NAND U7616 ( .A(n7029), .B(n7451), .Z(n7449) );
  NAND U7617 ( .A(n7452), .B(n7453), .Z(n7451) );
  NAND U7618 ( .A(n2503), .B(\stack[4][20] ), .Z(n7453) );
  NAND U7619 ( .A(n7033), .B(\stack[2][20] ), .Z(n7452) );
  NAND U7620 ( .A(n7454), .B(n7455), .Z(n2382) );
  NAND U7621 ( .A(n7028), .B(\stack[3][21] ), .Z(n7455) );
  NAND U7622 ( .A(n7029), .B(n7456), .Z(n7454) );
  NAND U7623 ( .A(n7457), .B(n7458), .Z(n7456) );
  NAND U7624 ( .A(n2503), .B(\stack[4][21] ), .Z(n7458) );
  NAND U7625 ( .A(n7033), .B(\stack[2][21] ), .Z(n7457) );
  NAND U7626 ( .A(n7459), .B(n7460), .Z(n2381) );
  NAND U7627 ( .A(n7028), .B(\stack[3][22] ), .Z(n7460) );
  NAND U7628 ( .A(n7029), .B(n7461), .Z(n7459) );
  NAND U7629 ( .A(n7462), .B(n7463), .Z(n7461) );
  NAND U7630 ( .A(n2503), .B(\stack[4][22] ), .Z(n7463) );
  NAND U7631 ( .A(n7033), .B(\stack[2][22] ), .Z(n7462) );
  NAND U7632 ( .A(n7464), .B(n7465), .Z(n2380) );
  NAND U7633 ( .A(n7028), .B(\stack[3][23] ), .Z(n7465) );
  NAND U7634 ( .A(n7029), .B(n7466), .Z(n7464) );
  NAND U7635 ( .A(n7467), .B(n7468), .Z(n7466) );
  NAND U7636 ( .A(n2503), .B(\stack[4][23] ), .Z(n7468) );
  NAND U7637 ( .A(n7033), .B(\stack[2][23] ), .Z(n7467) );
  NAND U7638 ( .A(n7469), .B(n7470), .Z(n2379) );
  NAND U7639 ( .A(n7028), .B(\stack[3][24] ), .Z(n7470) );
  NAND U7640 ( .A(n7029), .B(n7471), .Z(n7469) );
  NAND U7641 ( .A(n7472), .B(n7473), .Z(n7471) );
  NAND U7642 ( .A(n2503), .B(\stack[4][24] ), .Z(n7473) );
  NAND U7643 ( .A(n7033), .B(\stack[2][24] ), .Z(n7472) );
  NAND U7644 ( .A(n7474), .B(n7475), .Z(n2378) );
  NAND U7645 ( .A(n7028), .B(\stack[3][25] ), .Z(n7475) );
  NAND U7646 ( .A(n7029), .B(n7476), .Z(n7474) );
  NAND U7647 ( .A(n7477), .B(n7478), .Z(n7476) );
  NAND U7648 ( .A(n2503), .B(\stack[4][25] ), .Z(n7478) );
  NAND U7649 ( .A(n7033), .B(\stack[2][25] ), .Z(n7477) );
  NAND U7650 ( .A(n7479), .B(n7480), .Z(n2377) );
  NAND U7651 ( .A(n7028), .B(\stack[3][26] ), .Z(n7480) );
  NAND U7652 ( .A(n7029), .B(n7481), .Z(n7479) );
  NAND U7653 ( .A(n7482), .B(n7483), .Z(n7481) );
  NAND U7654 ( .A(n2503), .B(\stack[4][26] ), .Z(n7483) );
  NAND U7655 ( .A(n7033), .B(\stack[2][26] ), .Z(n7482) );
  NAND U7656 ( .A(n7484), .B(n7485), .Z(n2376) );
  NAND U7657 ( .A(n7028), .B(\stack[3][27] ), .Z(n7485) );
  NAND U7658 ( .A(n7029), .B(n7486), .Z(n7484) );
  NAND U7659 ( .A(n7487), .B(n7488), .Z(n7486) );
  NAND U7660 ( .A(n2503), .B(\stack[4][27] ), .Z(n7488) );
  NAND U7661 ( .A(n7033), .B(\stack[2][27] ), .Z(n7487) );
  NAND U7662 ( .A(n7489), .B(n7490), .Z(n2375) );
  NAND U7663 ( .A(n7028), .B(\stack[3][28] ), .Z(n7490) );
  NAND U7664 ( .A(n7029), .B(n7491), .Z(n7489) );
  NAND U7665 ( .A(n7492), .B(n7493), .Z(n7491) );
  NAND U7666 ( .A(n2503), .B(\stack[4][28] ), .Z(n7493) );
  NAND U7667 ( .A(n7033), .B(\stack[2][28] ), .Z(n7492) );
  NAND U7668 ( .A(n7494), .B(n7495), .Z(n2374) );
  NAND U7669 ( .A(n7028), .B(\stack[3][29] ), .Z(n7495) );
  NAND U7670 ( .A(n7029), .B(n7496), .Z(n7494) );
  NAND U7671 ( .A(n7497), .B(n7498), .Z(n7496) );
  NAND U7672 ( .A(n2503), .B(\stack[4][29] ), .Z(n7498) );
  NAND U7673 ( .A(n7033), .B(\stack[2][29] ), .Z(n7497) );
  NAND U7674 ( .A(n7499), .B(n7500), .Z(n2373) );
  NAND U7675 ( .A(n7028), .B(\stack[3][30] ), .Z(n7500) );
  NAND U7676 ( .A(n7029), .B(n7501), .Z(n7499) );
  NAND U7677 ( .A(n7502), .B(n7503), .Z(n7501) );
  NAND U7678 ( .A(n2503), .B(\stack[4][30] ), .Z(n7503) );
  NAND U7679 ( .A(n7033), .B(\stack[2][30] ), .Z(n7502) );
  NAND U7680 ( .A(n7504), .B(n7505), .Z(n2372) );
  NAND U7681 ( .A(n7028), .B(\stack[3][31] ), .Z(n7505) );
  NAND U7682 ( .A(n7029), .B(n7506), .Z(n7504) );
  NAND U7683 ( .A(n7507), .B(n7508), .Z(n7506) );
  NAND U7684 ( .A(n2503), .B(\stack[4][31] ), .Z(n7508) );
  NAND U7685 ( .A(n7033), .B(\stack[2][31] ), .Z(n7507) );
  NAND U7686 ( .A(n7509), .B(n7510), .Z(n2371) );
  NAND U7687 ( .A(n7028), .B(\stack[4][0] ), .Z(n7510) );
  NAND U7688 ( .A(n7029), .B(n7511), .Z(n7509) );
  NAND U7689 ( .A(n7512), .B(n7513), .Z(n7511) );
  NAND U7690 ( .A(n2503), .B(\stack[5][0] ), .Z(n7513) );
  NAND U7691 ( .A(n7033), .B(\stack[3][0] ), .Z(n7512) );
  NAND U7692 ( .A(n7514), .B(n7515), .Z(n2370) );
  NAND U7693 ( .A(n7028), .B(\stack[4][1] ), .Z(n7515) );
  NAND U7694 ( .A(n7029), .B(n7516), .Z(n7514) );
  NAND U7695 ( .A(n7517), .B(n7518), .Z(n7516) );
  NAND U7696 ( .A(n2503), .B(\stack[5][1] ), .Z(n7518) );
  NAND U7697 ( .A(n7033), .B(\stack[3][1] ), .Z(n7517) );
  NAND U7698 ( .A(n7519), .B(n7520), .Z(n2369) );
  NAND U7699 ( .A(n7028), .B(\stack[4][2] ), .Z(n7520) );
  NAND U7700 ( .A(n7029), .B(n7521), .Z(n7519) );
  NAND U7701 ( .A(n7522), .B(n7523), .Z(n7521) );
  NAND U7702 ( .A(n2503), .B(\stack[5][2] ), .Z(n7523) );
  NAND U7703 ( .A(n7033), .B(\stack[3][2] ), .Z(n7522) );
  NAND U7704 ( .A(n7524), .B(n7525), .Z(n2368) );
  NAND U7705 ( .A(n7028), .B(\stack[4][3] ), .Z(n7525) );
  NAND U7706 ( .A(n7029), .B(n7526), .Z(n7524) );
  NAND U7707 ( .A(n7527), .B(n7528), .Z(n7526) );
  NAND U7708 ( .A(n2503), .B(\stack[5][3] ), .Z(n7528) );
  NAND U7709 ( .A(n7033), .B(\stack[3][3] ), .Z(n7527) );
  NAND U7710 ( .A(n7529), .B(n7530), .Z(n2367) );
  NAND U7711 ( .A(n7028), .B(\stack[4][4] ), .Z(n7530) );
  NAND U7712 ( .A(n7029), .B(n7531), .Z(n7529) );
  NAND U7713 ( .A(n7532), .B(n7533), .Z(n7531) );
  NAND U7714 ( .A(n2503), .B(\stack[5][4] ), .Z(n7533) );
  NAND U7715 ( .A(n7033), .B(\stack[3][4] ), .Z(n7532) );
  NAND U7716 ( .A(n7534), .B(n7535), .Z(n2366) );
  NAND U7717 ( .A(n7028), .B(\stack[4][5] ), .Z(n7535) );
  NAND U7718 ( .A(n7029), .B(n7536), .Z(n7534) );
  NAND U7719 ( .A(n7537), .B(n7538), .Z(n7536) );
  NAND U7720 ( .A(n2503), .B(\stack[5][5] ), .Z(n7538) );
  NAND U7721 ( .A(n7033), .B(\stack[3][5] ), .Z(n7537) );
  NAND U7722 ( .A(n7539), .B(n7540), .Z(n2365) );
  NAND U7723 ( .A(n7028), .B(\stack[4][6] ), .Z(n7540) );
  NAND U7724 ( .A(n7029), .B(n7541), .Z(n7539) );
  NAND U7725 ( .A(n7542), .B(n7543), .Z(n7541) );
  NAND U7726 ( .A(n2503), .B(\stack[5][6] ), .Z(n7543) );
  NAND U7727 ( .A(n7033), .B(\stack[3][6] ), .Z(n7542) );
  NAND U7728 ( .A(n7544), .B(n7545), .Z(n2364) );
  NAND U7729 ( .A(n7028), .B(\stack[4][7] ), .Z(n7545) );
  NAND U7730 ( .A(n7029), .B(n7546), .Z(n7544) );
  NAND U7731 ( .A(n7547), .B(n7548), .Z(n7546) );
  NAND U7732 ( .A(n2503), .B(\stack[5][7] ), .Z(n7548) );
  NAND U7733 ( .A(n7033), .B(\stack[3][7] ), .Z(n7547) );
  NAND U7734 ( .A(n7549), .B(n7550), .Z(n2363) );
  NAND U7735 ( .A(n7028), .B(\stack[4][8] ), .Z(n7550) );
  NAND U7736 ( .A(n7029), .B(n7551), .Z(n7549) );
  NAND U7737 ( .A(n7552), .B(n7553), .Z(n7551) );
  NAND U7738 ( .A(n2503), .B(\stack[5][8] ), .Z(n7553) );
  NAND U7739 ( .A(n7033), .B(\stack[3][8] ), .Z(n7552) );
  NAND U7740 ( .A(n7554), .B(n7555), .Z(n2362) );
  NAND U7741 ( .A(n7028), .B(\stack[4][9] ), .Z(n7555) );
  NAND U7742 ( .A(n7029), .B(n7556), .Z(n7554) );
  NAND U7743 ( .A(n7557), .B(n7558), .Z(n7556) );
  NAND U7744 ( .A(n2503), .B(\stack[5][9] ), .Z(n7558) );
  NAND U7745 ( .A(n7033), .B(\stack[3][9] ), .Z(n7557) );
  NAND U7746 ( .A(n7559), .B(n7560), .Z(n2361) );
  NAND U7747 ( .A(n7028), .B(\stack[4][10] ), .Z(n7560) );
  NAND U7748 ( .A(n7029), .B(n7561), .Z(n7559) );
  NAND U7749 ( .A(n7562), .B(n7563), .Z(n7561) );
  NAND U7750 ( .A(n2503), .B(\stack[5][10] ), .Z(n7563) );
  NAND U7751 ( .A(n7033), .B(\stack[3][10] ), .Z(n7562) );
  NAND U7752 ( .A(n7564), .B(n7565), .Z(n2360) );
  NAND U7753 ( .A(n7028), .B(\stack[4][11] ), .Z(n7565) );
  NAND U7754 ( .A(n7029), .B(n7566), .Z(n7564) );
  NAND U7755 ( .A(n7567), .B(n7568), .Z(n7566) );
  NAND U7756 ( .A(n2503), .B(\stack[5][11] ), .Z(n7568) );
  NAND U7757 ( .A(n7033), .B(\stack[3][11] ), .Z(n7567) );
  NAND U7758 ( .A(n7569), .B(n7570), .Z(n2359) );
  NAND U7759 ( .A(n7028), .B(\stack[4][12] ), .Z(n7570) );
  NAND U7760 ( .A(n7029), .B(n7571), .Z(n7569) );
  NAND U7761 ( .A(n7572), .B(n7573), .Z(n7571) );
  NAND U7762 ( .A(n2503), .B(\stack[5][12] ), .Z(n7573) );
  NAND U7763 ( .A(n7033), .B(\stack[3][12] ), .Z(n7572) );
  NAND U7764 ( .A(n7574), .B(n7575), .Z(n2358) );
  NAND U7765 ( .A(n7028), .B(\stack[4][13] ), .Z(n7575) );
  NAND U7766 ( .A(n7029), .B(n7576), .Z(n7574) );
  NAND U7767 ( .A(n7577), .B(n7578), .Z(n7576) );
  NAND U7768 ( .A(n2503), .B(\stack[5][13] ), .Z(n7578) );
  NAND U7769 ( .A(n7033), .B(\stack[3][13] ), .Z(n7577) );
  NAND U7770 ( .A(n7579), .B(n7580), .Z(n2357) );
  NAND U7771 ( .A(n7028), .B(\stack[4][14] ), .Z(n7580) );
  NAND U7772 ( .A(n7029), .B(n7581), .Z(n7579) );
  NAND U7773 ( .A(n7582), .B(n7583), .Z(n7581) );
  NAND U7774 ( .A(n2503), .B(\stack[5][14] ), .Z(n7583) );
  NAND U7775 ( .A(n7033), .B(\stack[3][14] ), .Z(n7582) );
  NAND U7776 ( .A(n7584), .B(n7585), .Z(n2356) );
  NAND U7777 ( .A(n7028), .B(\stack[4][15] ), .Z(n7585) );
  NAND U7778 ( .A(n7029), .B(n7586), .Z(n7584) );
  NAND U7779 ( .A(n7587), .B(n7588), .Z(n7586) );
  NAND U7780 ( .A(n2503), .B(\stack[5][15] ), .Z(n7588) );
  NAND U7781 ( .A(n7033), .B(\stack[3][15] ), .Z(n7587) );
  NAND U7782 ( .A(n7589), .B(n7590), .Z(n2355) );
  NAND U7783 ( .A(n7028), .B(\stack[4][16] ), .Z(n7590) );
  NAND U7784 ( .A(n7029), .B(n7591), .Z(n7589) );
  NAND U7785 ( .A(n7592), .B(n7593), .Z(n7591) );
  NAND U7786 ( .A(n2503), .B(\stack[5][16] ), .Z(n7593) );
  NAND U7787 ( .A(n7033), .B(\stack[3][16] ), .Z(n7592) );
  NAND U7788 ( .A(n7594), .B(n7595), .Z(n2354) );
  NAND U7789 ( .A(n7028), .B(\stack[4][17] ), .Z(n7595) );
  NAND U7790 ( .A(n7029), .B(n7596), .Z(n7594) );
  NAND U7791 ( .A(n7597), .B(n7598), .Z(n7596) );
  NAND U7792 ( .A(n2503), .B(\stack[5][17] ), .Z(n7598) );
  NAND U7793 ( .A(n7033), .B(\stack[3][17] ), .Z(n7597) );
  NAND U7794 ( .A(n7599), .B(n7600), .Z(n2353) );
  NAND U7795 ( .A(n7028), .B(\stack[4][18] ), .Z(n7600) );
  NAND U7796 ( .A(n7029), .B(n7601), .Z(n7599) );
  NAND U7797 ( .A(n7602), .B(n7603), .Z(n7601) );
  NAND U7798 ( .A(n2503), .B(\stack[5][18] ), .Z(n7603) );
  NAND U7799 ( .A(n7033), .B(\stack[3][18] ), .Z(n7602) );
  NAND U7800 ( .A(n7604), .B(n7605), .Z(n2352) );
  NAND U7801 ( .A(n7028), .B(\stack[4][19] ), .Z(n7605) );
  NAND U7802 ( .A(n7029), .B(n7606), .Z(n7604) );
  NAND U7803 ( .A(n7607), .B(n7608), .Z(n7606) );
  NAND U7804 ( .A(n2503), .B(\stack[5][19] ), .Z(n7608) );
  NAND U7805 ( .A(n7033), .B(\stack[3][19] ), .Z(n7607) );
  NAND U7806 ( .A(n7609), .B(n7610), .Z(n2351) );
  NAND U7807 ( .A(n7028), .B(\stack[4][20] ), .Z(n7610) );
  NAND U7808 ( .A(n7029), .B(n7611), .Z(n7609) );
  NAND U7809 ( .A(n7612), .B(n7613), .Z(n7611) );
  NAND U7810 ( .A(n2503), .B(\stack[5][20] ), .Z(n7613) );
  NAND U7811 ( .A(n7033), .B(\stack[3][20] ), .Z(n7612) );
  NAND U7812 ( .A(n7614), .B(n7615), .Z(n2350) );
  NAND U7813 ( .A(n7028), .B(\stack[4][21] ), .Z(n7615) );
  NAND U7814 ( .A(n7029), .B(n7616), .Z(n7614) );
  NAND U7815 ( .A(n7617), .B(n7618), .Z(n7616) );
  NAND U7816 ( .A(n2503), .B(\stack[5][21] ), .Z(n7618) );
  NAND U7817 ( .A(n7033), .B(\stack[3][21] ), .Z(n7617) );
  NAND U7818 ( .A(n7619), .B(n7620), .Z(n2349) );
  NAND U7819 ( .A(n7028), .B(\stack[4][22] ), .Z(n7620) );
  NAND U7820 ( .A(n7029), .B(n7621), .Z(n7619) );
  NAND U7821 ( .A(n7622), .B(n7623), .Z(n7621) );
  NAND U7822 ( .A(n2503), .B(\stack[5][22] ), .Z(n7623) );
  NAND U7823 ( .A(n7033), .B(\stack[3][22] ), .Z(n7622) );
  NAND U7824 ( .A(n7624), .B(n7625), .Z(n2348) );
  NAND U7825 ( .A(n7028), .B(\stack[4][23] ), .Z(n7625) );
  NAND U7826 ( .A(n7029), .B(n7626), .Z(n7624) );
  NAND U7827 ( .A(n7627), .B(n7628), .Z(n7626) );
  NAND U7828 ( .A(n2503), .B(\stack[5][23] ), .Z(n7628) );
  NAND U7829 ( .A(n7033), .B(\stack[3][23] ), .Z(n7627) );
  NAND U7830 ( .A(n7629), .B(n7630), .Z(n2347) );
  NAND U7831 ( .A(n7028), .B(\stack[4][24] ), .Z(n7630) );
  NAND U7832 ( .A(n7029), .B(n7631), .Z(n7629) );
  NAND U7833 ( .A(n7632), .B(n7633), .Z(n7631) );
  NAND U7834 ( .A(n2503), .B(\stack[5][24] ), .Z(n7633) );
  NAND U7835 ( .A(n7033), .B(\stack[3][24] ), .Z(n7632) );
  NAND U7836 ( .A(n7634), .B(n7635), .Z(n2346) );
  NAND U7837 ( .A(n7028), .B(\stack[4][25] ), .Z(n7635) );
  NAND U7838 ( .A(n7029), .B(n7636), .Z(n7634) );
  NAND U7839 ( .A(n7637), .B(n7638), .Z(n7636) );
  NAND U7840 ( .A(n2503), .B(\stack[5][25] ), .Z(n7638) );
  NAND U7841 ( .A(n7033), .B(\stack[3][25] ), .Z(n7637) );
  NAND U7842 ( .A(n7639), .B(n7640), .Z(n2345) );
  NAND U7843 ( .A(n7028), .B(\stack[4][26] ), .Z(n7640) );
  NAND U7844 ( .A(n7029), .B(n7641), .Z(n7639) );
  NAND U7845 ( .A(n7642), .B(n7643), .Z(n7641) );
  NAND U7846 ( .A(n2503), .B(\stack[5][26] ), .Z(n7643) );
  NAND U7847 ( .A(n7033), .B(\stack[3][26] ), .Z(n7642) );
  NAND U7848 ( .A(n7644), .B(n7645), .Z(n2344) );
  NAND U7849 ( .A(n7028), .B(\stack[4][27] ), .Z(n7645) );
  NAND U7850 ( .A(n7029), .B(n7646), .Z(n7644) );
  NAND U7851 ( .A(n7647), .B(n7648), .Z(n7646) );
  NAND U7852 ( .A(n2503), .B(\stack[5][27] ), .Z(n7648) );
  NAND U7853 ( .A(n7033), .B(\stack[3][27] ), .Z(n7647) );
  NAND U7854 ( .A(n7649), .B(n7650), .Z(n2343) );
  NAND U7855 ( .A(n7028), .B(\stack[4][28] ), .Z(n7650) );
  NAND U7856 ( .A(n7029), .B(n7651), .Z(n7649) );
  NAND U7857 ( .A(n7652), .B(n7653), .Z(n7651) );
  NAND U7858 ( .A(n2503), .B(\stack[5][28] ), .Z(n7653) );
  NAND U7859 ( .A(n7033), .B(\stack[3][28] ), .Z(n7652) );
  NAND U7860 ( .A(n7654), .B(n7655), .Z(n2342) );
  NAND U7861 ( .A(n7028), .B(\stack[4][29] ), .Z(n7655) );
  NAND U7862 ( .A(n7029), .B(n7656), .Z(n7654) );
  NAND U7863 ( .A(n7657), .B(n7658), .Z(n7656) );
  NAND U7864 ( .A(n2503), .B(\stack[5][29] ), .Z(n7658) );
  NAND U7865 ( .A(n7033), .B(\stack[3][29] ), .Z(n7657) );
  NAND U7866 ( .A(n7659), .B(n7660), .Z(n2341) );
  NAND U7867 ( .A(n7028), .B(\stack[4][30] ), .Z(n7660) );
  NAND U7868 ( .A(n7029), .B(n7661), .Z(n7659) );
  NAND U7869 ( .A(n7662), .B(n7663), .Z(n7661) );
  NAND U7870 ( .A(n2503), .B(\stack[5][30] ), .Z(n7663) );
  NAND U7871 ( .A(n7033), .B(\stack[3][30] ), .Z(n7662) );
  NAND U7872 ( .A(n7664), .B(n7665), .Z(n2340) );
  NAND U7873 ( .A(n7028), .B(\stack[4][31] ), .Z(n7665) );
  NAND U7874 ( .A(n7029), .B(n7666), .Z(n7664) );
  NAND U7875 ( .A(n7667), .B(n7668), .Z(n7666) );
  NAND U7876 ( .A(n2503), .B(\stack[5][31] ), .Z(n7668) );
  NAND U7877 ( .A(n7033), .B(\stack[3][31] ), .Z(n7667) );
  NAND U7878 ( .A(n7669), .B(n7670), .Z(n2339) );
  NAND U7879 ( .A(n7028), .B(\stack[5][0] ), .Z(n7670) );
  NAND U7880 ( .A(n7029), .B(n7671), .Z(n7669) );
  NAND U7881 ( .A(n7672), .B(n7673), .Z(n7671) );
  NAND U7882 ( .A(n2503), .B(\stack[6][0] ), .Z(n7673) );
  NAND U7883 ( .A(n7033), .B(\stack[4][0] ), .Z(n7672) );
  NAND U7884 ( .A(n7674), .B(n7675), .Z(n2338) );
  NAND U7885 ( .A(n7028), .B(\stack[5][1] ), .Z(n7675) );
  NAND U7886 ( .A(n7029), .B(n7676), .Z(n7674) );
  NAND U7887 ( .A(n7677), .B(n7678), .Z(n7676) );
  NAND U7888 ( .A(n2503), .B(\stack[6][1] ), .Z(n7678) );
  NAND U7889 ( .A(n7033), .B(\stack[4][1] ), .Z(n7677) );
  NAND U7890 ( .A(n7679), .B(n7680), .Z(n2337) );
  NAND U7891 ( .A(n7028), .B(\stack[5][2] ), .Z(n7680) );
  NAND U7892 ( .A(n7029), .B(n7681), .Z(n7679) );
  NAND U7893 ( .A(n7682), .B(n7683), .Z(n7681) );
  NAND U7894 ( .A(n2503), .B(\stack[6][2] ), .Z(n7683) );
  NAND U7895 ( .A(n7033), .B(\stack[4][2] ), .Z(n7682) );
  NAND U7896 ( .A(n7684), .B(n7685), .Z(n2336) );
  NAND U7897 ( .A(n7028), .B(\stack[5][3] ), .Z(n7685) );
  NAND U7898 ( .A(n7029), .B(n7686), .Z(n7684) );
  NAND U7899 ( .A(n7687), .B(n7688), .Z(n7686) );
  NAND U7900 ( .A(n2503), .B(\stack[6][3] ), .Z(n7688) );
  NAND U7901 ( .A(n7033), .B(\stack[4][3] ), .Z(n7687) );
  NAND U7902 ( .A(n7689), .B(n7690), .Z(n2335) );
  NAND U7903 ( .A(n7028), .B(\stack[5][4] ), .Z(n7690) );
  NAND U7904 ( .A(n7029), .B(n7691), .Z(n7689) );
  NAND U7905 ( .A(n7692), .B(n7693), .Z(n7691) );
  NAND U7906 ( .A(n2503), .B(\stack[6][4] ), .Z(n7693) );
  NAND U7907 ( .A(n7033), .B(\stack[4][4] ), .Z(n7692) );
  NAND U7908 ( .A(n7694), .B(n7695), .Z(n2334) );
  NAND U7909 ( .A(n7028), .B(\stack[5][5] ), .Z(n7695) );
  NAND U7910 ( .A(n7029), .B(n7696), .Z(n7694) );
  NAND U7911 ( .A(n7697), .B(n7698), .Z(n7696) );
  NAND U7912 ( .A(n2503), .B(\stack[6][5] ), .Z(n7698) );
  NAND U7913 ( .A(n7033), .B(\stack[4][5] ), .Z(n7697) );
  NAND U7914 ( .A(n7699), .B(n7700), .Z(n2333) );
  NAND U7915 ( .A(n7028), .B(\stack[5][6] ), .Z(n7700) );
  NAND U7916 ( .A(n7029), .B(n7701), .Z(n7699) );
  NAND U7917 ( .A(n7702), .B(n7703), .Z(n7701) );
  NAND U7918 ( .A(n2503), .B(\stack[6][6] ), .Z(n7703) );
  NAND U7919 ( .A(n7033), .B(\stack[4][6] ), .Z(n7702) );
  NAND U7920 ( .A(n7704), .B(n7705), .Z(n2332) );
  NAND U7921 ( .A(n7028), .B(\stack[5][7] ), .Z(n7705) );
  NAND U7922 ( .A(n7029), .B(n7706), .Z(n7704) );
  NAND U7923 ( .A(n7707), .B(n7708), .Z(n7706) );
  NAND U7924 ( .A(n2503), .B(\stack[6][7] ), .Z(n7708) );
  NAND U7925 ( .A(n7033), .B(\stack[4][7] ), .Z(n7707) );
  NAND U7926 ( .A(n7709), .B(n7710), .Z(n2331) );
  NAND U7927 ( .A(n7028), .B(\stack[5][8] ), .Z(n7710) );
  NAND U7928 ( .A(n7029), .B(n7711), .Z(n7709) );
  NAND U7929 ( .A(n7712), .B(n7713), .Z(n7711) );
  NAND U7930 ( .A(n2503), .B(\stack[6][8] ), .Z(n7713) );
  NAND U7931 ( .A(n7033), .B(\stack[4][8] ), .Z(n7712) );
  NAND U7932 ( .A(n7714), .B(n7715), .Z(n2330) );
  NAND U7933 ( .A(n7028), .B(\stack[5][9] ), .Z(n7715) );
  NAND U7934 ( .A(n7029), .B(n7716), .Z(n7714) );
  NAND U7935 ( .A(n7717), .B(n7718), .Z(n7716) );
  NAND U7936 ( .A(n2503), .B(\stack[6][9] ), .Z(n7718) );
  NAND U7937 ( .A(n7033), .B(\stack[4][9] ), .Z(n7717) );
  NAND U7938 ( .A(n7719), .B(n7720), .Z(n2329) );
  NAND U7939 ( .A(n7028), .B(\stack[5][10] ), .Z(n7720) );
  NAND U7940 ( .A(n7029), .B(n7721), .Z(n7719) );
  NAND U7941 ( .A(n7722), .B(n7723), .Z(n7721) );
  NAND U7942 ( .A(n2503), .B(\stack[6][10] ), .Z(n7723) );
  NAND U7943 ( .A(n7033), .B(\stack[4][10] ), .Z(n7722) );
  NAND U7944 ( .A(n7724), .B(n7725), .Z(n2328) );
  NAND U7945 ( .A(n7028), .B(\stack[5][11] ), .Z(n7725) );
  NAND U7946 ( .A(n7029), .B(n7726), .Z(n7724) );
  NAND U7947 ( .A(n7727), .B(n7728), .Z(n7726) );
  NAND U7948 ( .A(n2503), .B(\stack[6][11] ), .Z(n7728) );
  NAND U7949 ( .A(n7033), .B(\stack[4][11] ), .Z(n7727) );
  NAND U7950 ( .A(n7729), .B(n7730), .Z(n2327) );
  NAND U7951 ( .A(n7028), .B(\stack[5][12] ), .Z(n7730) );
  NAND U7952 ( .A(n7029), .B(n7731), .Z(n7729) );
  NAND U7953 ( .A(n7732), .B(n7733), .Z(n7731) );
  NAND U7954 ( .A(n2503), .B(\stack[6][12] ), .Z(n7733) );
  NAND U7955 ( .A(n7033), .B(\stack[4][12] ), .Z(n7732) );
  NAND U7956 ( .A(n7734), .B(n7735), .Z(n2326) );
  NAND U7957 ( .A(n7028), .B(\stack[5][13] ), .Z(n7735) );
  NAND U7958 ( .A(n7029), .B(n7736), .Z(n7734) );
  NAND U7959 ( .A(n7737), .B(n7738), .Z(n7736) );
  NAND U7960 ( .A(n2503), .B(\stack[6][13] ), .Z(n7738) );
  NAND U7961 ( .A(n7033), .B(\stack[4][13] ), .Z(n7737) );
  NAND U7962 ( .A(n7739), .B(n7740), .Z(n2325) );
  NAND U7963 ( .A(n7028), .B(\stack[5][14] ), .Z(n7740) );
  NAND U7964 ( .A(n7029), .B(n7741), .Z(n7739) );
  NAND U7965 ( .A(n7742), .B(n7743), .Z(n7741) );
  NAND U7966 ( .A(n2503), .B(\stack[6][14] ), .Z(n7743) );
  NAND U7967 ( .A(n7033), .B(\stack[4][14] ), .Z(n7742) );
  NAND U7968 ( .A(n7744), .B(n7745), .Z(n2324) );
  NAND U7969 ( .A(n7028), .B(\stack[5][15] ), .Z(n7745) );
  NAND U7970 ( .A(n7029), .B(n7746), .Z(n7744) );
  NAND U7971 ( .A(n7747), .B(n7748), .Z(n7746) );
  NAND U7972 ( .A(n2503), .B(\stack[6][15] ), .Z(n7748) );
  NAND U7973 ( .A(n7033), .B(\stack[4][15] ), .Z(n7747) );
  NAND U7974 ( .A(n7749), .B(n7750), .Z(n2323) );
  NAND U7975 ( .A(n7028), .B(\stack[5][16] ), .Z(n7750) );
  NAND U7976 ( .A(n7029), .B(n7751), .Z(n7749) );
  NAND U7977 ( .A(n7752), .B(n7753), .Z(n7751) );
  NAND U7978 ( .A(n2503), .B(\stack[6][16] ), .Z(n7753) );
  NAND U7979 ( .A(n7033), .B(\stack[4][16] ), .Z(n7752) );
  NAND U7980 ( .A(n7754), .B(n7755), .Z(n2322) );
  NAND U7981 ( .A(n7028), .B(\stack[5][17] ), .Z(n7755) );
  NAND U7982 ( .A(n7029), .B(n7756), .Z(n7754) );
  NAND U7983 ( .A(n7757), .B(n7758), .Z(n7756) );
  NAND U7984 ( .A(n2503), .B(\stack[6][17] ), .Z(n7758) );
  NAND U7985 ( .A(n7033), .B(\stack[4][17] ), .Z(n7757) );
  NAND U7986 ( .A(n7759), .B(n7760), .Z(n2321) );
  NAND U7987 ( .A(n7028), .B(\stack[5][18] ), .Z(n7760) );
  NAND U7988 ( .A(n7029), .B(n7761), .Z(n7759) );
  NAND U7989 ( .A(n7762), .B(n7763), .Z(n7761) );
  NAND U7990 ( .A(n2503), .B(\stack[6][18] ), .Z(n7763) );
  NAND U7991 ( .A(n7033), .B(\stack[4][18] ), .Z(n7762) );
  NAND U7992 ( .A(n7764), .B(n7765), .Z(n2320) );
  NAND U7993 ( .A(n7028), .B(\stack[5][19] ), .Z(n7765) );
  NAND U7994 ( .A(n7029), .B(n7766), .Z(n7764) );
  NAND U7995 ( .A(n7767), .B(n7768), .Z(n7766) );
  NAND U7996 ( .A(n2503), .B(\stack[6][19] ), .Z(n7768) );
  NAND U7997 ( .A(n7033), .B(\stack[4][19] ), .Z(n7767) );
  NAND U7998 ( .A(n7769), .B(n7770), .Z(n2319) );
  NAND U7999 ( .A(n7028), .B(\stack[5][20] ), .Z(n7770) );
  NAND U8000 ( .A(n7029), .B(n7771), .Z(n7769) );
  NAND U8001 ( .A(n7772), .B(n7773), .Z(n7771) );
  NAND U8002 ( .A(n2503), .B(\stack[6][20] ), .Z(n7773) );
  NAND U8003 ( .A(n7033), .B(\stack[4][20] ), .Z(n7772) );
  NAND U8004 ( .A(n7774), .B(n7775), .Z(n2318) );
  NAND U8005 ( .A(n7028), .B(\stack[5][21] ), .Z(n7775) );
  NAND U8006 ( .A(n7029), .B(n7776), .Z(n7774) );
  NAND U8007 ( .A(n7777), .B(n7778), .Z(n7776) );
  NAND U8008 ( .A(n2503), .B(\stack[6][21] ), .Z(n7778) );
  NAND U8009 ( .A(n7033), .B(\stack[4][21] ), .Z(n7777) );
  NAND U8010 ( .A(n7779), .B(n7780), .Z(n2317) );
  NAND U8011 ( .A(n7028), .B(\stack[5][22] ), .Z(n7780) );
  NAND U8012 ( .A(n7029), .B(n7781), .Z(n7779) );
  NAND U8013 ( .A(n7782), .B(n7783), .Z(n7781) );
  NAND U8014 ( .A(n2503), .B(\stack[6][22] ), .Z(n7783) );
  NAND U8015 ( .A(n7033), .B(\stack[4][22] ), .Z(n7782) );
  NAND U8016 ( .A(n7784), .B(n7785), .Z(n2316) );
  NAND U8017 ( .A(n7028), .B(\stack[5][23] ), .Z(n7785) );
  NAND U8018 ( .A(n7029), .B(n7786), .Z(n7784) );
  NAND U8019 ( .A(n7787), .B(n7788), .Z(n7786) );
  NAND U8020 ( .A(n2503), .B(\stack[6][23] ), .Z(n7788) );
  NAND U8021 ( .A(n7033), .B(\stack[4][23] ), .Z(n7787) );
  NAND U8022 ( .A(n7789), .B(n7790), .Z(n2315) );
  NAND U8023 ( .A(n7028), .B(\stack[5][24] ), .Z(n7790) );
  NAND U8024 ( .A(n7029), .B(n7791), .Z(n7789) );
  NAND U8025 ( .A(n7792), .B(n7793), .Z(n7791) );
  NAND U8026 ( .A(n2503), .B(\stack[6][24] ), .Z(n7793) );
  NAND U8027 ( .A(n7033), .B(\stack[4][24] ), .Z(n7792) );
  NAND U8028 ( .A(n7794), .B(n7795), .Z(n2314) );
  NAND U8029 ( .A(n7028), .B(\stack[5][25] ), .Z(n7795) );
  NAND U8030 ( .A(n7029), .B(n7796), .Z(n7794) );
  NAND U8031 ( .A(n7797), .B(n7798), .Z(n7796) );
  NAND U8032 ( .A(n2503), .B(\stack[6][25] ), .Z(n7798) );
  NAND U8033 ( .A(n7033), .B(\stack[4][25] ), .Z(n7797) );
  NAND U8034 ( .A(n7799), .B(n7800), .Z(n2313) );
  NAND U8035 ( .A(n7028), .B(\stack[5][26] ), .Z(n7800) );
  NAND U8036 ( .A(n7029), .B(n7801), .Z(n7799) );
  NAND U8037 ( .A(n7802), .B(n7803), .Z(n7801) );
  NAND U8038 ( .A(n2503), .B(\stack[6][26] ), .Z(n7803) );
  NAND U8039 ( .A(n7033), .B(\stack[4][26] ), .Z(n7802) );
  NAND U8040 ( .A(n7804), .B(n7805), .Z(n2312) );
  NAND U8041 ( .A(n7028), .B(\stack[5][27] ), .Z(n7805) );
  NAND U8042 ( .A(n7029), .B(n7806), .Z(n7804) );
  NAND U8043 ( .A(n7807), .B(n7808), .Z(n7806) );
  NAND U8044 ( .A(n2503), .B(\stack[6][27] ), .Z(n7808) );
  NAND U8045 ( .A(n7033), .B(\stack[4][27] ), .Z(n7807) );
  NAND U8046 ( .A(n7809), .B(n7810), .Z(n2311) );
  NAND U8047 ( .A(n7028), .B(\stack[5][28] ), .Z(n7810) );
  NAND U8048 ( .A(n7029), .B(n7811), .Z(n7809) );
  NAND U8049 ( .A(n7812), .B(n7813), .Z(n7811) );
  NAND U8050 ( .A(n2503), .B(\stack[6][28] ), .Z(n7813) );
  NAND U8051 ( .A(n7033), .B(\stack[4][28] ), .Z(n7812) );
  NAND U8052 ( .A(n7814), .B(n7815), .Z(n2310) );
  NAND U8053 ( .A(n7028), .B(\stack[5][29] ), .Z(n7815) );
  NAND U8054 ( .A(n7029), .B(n7816), .Z(n7814) );
  NAND U8055 ( .A(n7817), .B(n7818), .Z(n7816) );
  NAND U8056 ( .A(n2503), .B(\stack[6][29] ), .Z(n7818) );
  NAND U8057 ( .A(n7033), .B(\stack[4][29] ), .Z(n7817) );
  NAND U8058 ( .A(n7819), .B(n7820), .Z(n2309) );
  NAND U8059 ( .A(n7028), .B(\stack[5][30] ), .Z(n7820) );
  NAND U8060 ( .A(n7029), .B(n7821), .Z(n7819) );
  NAND U8061 ( .A(n7822), .B(n7823), .Z(n7821) );
  NAND U8062 ( .A(n2503), .B(\stack[6][30] ), .Z(n7823) );
  NAND U8063 ( .A(n7033), .B(\stack[4][30] ), .Z(n7822) );
  NAND U8064 ( .A(n7824), .B(n7825), .Z(n2308) );
  NAND U8065 ( .A(n7028), .B(\stack[5][31] ), .Z(n7825) );
  NAND U8066 ( .A(n7029), .B(n7826), .Z(n7824) );
  NAND U8067 ( .A(n7827), .B(n7828), .Z(n7826) );
  NAND U8068 ( .A(n2503), .B(\stack[6][31] ), .Z(n7828) );
  NAND U8069 ( .A(n7033), .B(\stack[4][31] ), .Z(n7827) );
  NAND U8070 ( .A(n7829), .B(n7830), .Z(n2307) );
  NAND U8071 ( .A(n7028), .B(\stack[6][0] ), .Z(n7830) );
  NAND U8072 ( .A(n7029), .B(n7831), .Z(n7829) );
  NANDN U8073 ( .A(n7832), .B(n7833), .Z(n7831) );
  NAND U8074 ( .A(n7033), .B(\stack[5][0] ), .Z(n7833) );
  NAND U8075 ( .A(n7834), .B(n7835), .Z(n2306) );
  NAND U8076 ( .A(n7028), .B(\stack[6][1] ), .Z(n7835) );
  NAND U8077 ( .A(n7029), .B(n7836), .Z(n7834) );
  NANDN U8078 ( .A(n7837), .B(n7838), .Z(n7836) );
  NAND U8079 ( .A(n7033), .B(\stack[5][1] ), .Z(n7838) );
  NAND U8080 ( .A(n7839), .B(n7840), .Z(n2305) );
  NAND U8081 ( .A(n7028), .B(\stack[6][2] ), .Z(n7840) );
  NAND U8082 ( .A(n7029), .B(n7841), .Z(n7839) );
  NANDN U8083 ( .A(n7842), .B(n7843), .Z(n7841) );
  NAND U8084 ( .A(n7033), .B(\stack[5][2] ), .Z(n7843) );
  NAND U8085 ( .A(n7844), .B(n7845), .Z(n2304) );
  NAND U8086 ( .A(n7028), .B(\stack[6][3] ), .Z(n7845) );
  NAND U8087 ( .A(n7029), .B(n7846), .Z(n7844) );
  NANDN U8088 ( .A(n7847), .B(n7848), .Z(n7846) );
  NAND U8089 ( .A(n7033), .B(\stack[5][3] ), .Z(n7848) );
  NAND U8090 ( .A(n7849), .B(n7850), .Z(n2303) );
  NAND U8091 ( .A(n7028), .B(\stack[6][4] ), .Z(n7850) );
  NAND U8092 ( .A(n7029), .B(n7851), .Z(n7849) );
  NANDN U8093 ( .A(n7852), .B(n7853), .Z(n7851) );
  NAND U8094 ( .A(n7033), .B(\stack[5][4] ), .Z(n7853) );
  NAND U8095 ( .A(n7854), .B(n7855), .Z(n2302) );
  NAND U8096 ( .A(n7028), .B(\stack[6][5] ), .Z(n7855) );
  NAND U8097 ( .A(n7029), .B(n7856), .Z(n7854) );
  NANDN U8098 ( .A(n7857), .B(n7858), .Z(n7856) );
  NAND U8099 ( .A(n7033), .B(\stack[5][5] ), .Z(n7858) );
  NAND U8100 ( .A(n7859), .B(n7860), .Z(n2301) );
  NAND U8101 ( .A(n7028), .B(\stack[6][6] ), .Z(n7860) );
  NAND U8102 ( .A(n7029), .B(n7861), .Z(n7859) );
  NANDN U8103 ( .A(n7862), .B(n7863), .Z(n7861) );
  NAND U8104 ( .A(n7033), .B(\stack[5][6] ), .Z(n7863) );
  NAND U8105 ( .A(n7864), .B(n7865), .Z(n2300) );
  NAND U8106 ( .A(n7028), .B(\stack[6][7] ), .Z(n7865) );
  NAND U8107 ( .A(n7029), .B(n7866), .Z(n7864) );
  NANDN U8108 ( .A(n7867), .B(n7868), .Z(n7866) );
  NAND U8109 ( .A(n7033), .B(\stack[5][7] ), .Z(n7868) );
  NAND U8110 ( .A(n7869), .B(n7870), .Z(n2299) );
  NAND U8111 ( .A(n7028), .B(\stack[6][8] ), .Z(n7870) );
  NAND U8112 ( .A(n7029), .B(n7871), .Z(n7869) );
  NANDN U8113 ( .A(n7872), .B(n7873), .Z(n7871) );
  NAND U8114 ( .A(n7033), .B(\stack[5][8] ), .Z(n7873) );
  NAND U8115 ( .A(n7874), .B(n7875), .Z(n2298) );
  NAND U8116 ( .A(n7028), .B(\stack[6][9] ), .Z(n7875) );
  NAND U8117 ( .A(n7029), .B(n7876), .Z(n7874) );
  NANDN U8118 ( .A(n7877), .B(n7878), .Z(n7876) );
  NAND U8119 ( .A(n7033), .B(\stack[5][9] ), .Z(n7878) );
  NAND U8120 ( .A(n7879), .B(n7880), .Z(n2297) );
  NAND U8121 ( .A(n7028), .B(\stack[6][10] ), .Z(n7880) );
  NAND U8122 ( .A(n7029), .B(n7881), .Z(n7879) );
  NANDN U8123 ( .A(n7882), .B(n7883), .Z(n7881) );
  NAND U8124 ( .A(n7033), .B(\stack[5][10] ), .Z(n7883) );
  NAND U8125 ( .A(n7884), .B(n7885), .Z(n2296) );
  NAND U8126 ( .A(n7028), .B(\stack[6][11] ), .Z(n7885) );
  NAND U8127 ( .A(n7029), .B(n7886), .Z(n7884) );
  NANDN U8128 ( .A(n7887), .B(n7888), .Z(n7886) );
  NAND U8129 ( .A(n7033), .B(\stack[5][11] ), .Z(n7888) );
  NAND U8130 ( .A(n7889), .B(n7890), .Z(n2295) );
  NAND U8131 ( .A(n7028), .B(\stack[6][12] ), .Z(n7890) );
  NAND U8132 ( .A(n7029), .B(n7891), .Z(n7889) );
  NANDN U8133 ( .A(n7892), .B(n7893), .Z(n7891) );
  NAND U8134 ( .A(n7033), .B(\stack[5][12] ), .Z(n7893) );
  NAND U8135 ( .A(n7894), .B(n7895), .Z(n2294) );
  NAND U8136 ( .A(n7028), .B(\stack[6][13] ), .Z(n7895) );
  NAND U8137 ( .A(n7029), .B(n7896), .Z(n7894) );
  NANDN U8138 ( .A(n7897), .B(n7898), .Z(n7896) );
  NAND U8139 ( .A(n7033), .B(\stack[5][13] ), .Z(n7898) );
  NAND U8140 ( .A(n7899), .B(n7900), .Z(n2293) );
  NAND U8141 ( .A(n7028), .B(\stack[6][14] ), .Z(n7900) );
  NAND U8142 ( .A(n7029), .B(n7901), .Z(n7899) );
  NANDN U8143 ( .A(n7902), .B(n7903), .Z(n7901) );
  NAND U8144 ( .A(n7033), .B(\stack[5][14] ), .Z(n7903) );
  NAND U8145 ( .A(n7904), .B(n7905), .Z(n2292) );
  NAND U8146 ( .A(n7028), .B(\stack[6][15] ), .Z(n7905) );
  NAND U8147 ( .A(n7029), .B(n7906), .Z(n7904) );
  NANDN U8148 ( .A(n7907), .B(n7908), .Z(n7906) );
  NAND U8149 ( .A(n7033), .B(\stack[5][15] ), .Z(n7908) );
  NAND U8150 ( .A(n7909), .B(n7910), .Z(n2291) );
  NAND U8151 ( .A(n7028), .B(\stack[6][16] ), .Z(n7910) );
  NAND U8152 ( .A(n7029), .B(n7911), .Z(n7909) );
  NANDN U8153 ( .A(n7912), .B(n7913), .Z(n7911) );
  NAND U8154 ( .A(n7033), .B(\stack[5][16] ), .Z(n7913) );
  NAND U8155 ( .A(n7914), .B(n7915), .Z(n2290) );
  NAND U8156 ( .A(n7028), .B(\stack[6][17] ), .Z(n7915) );
  NAND U8157 ( .A(n7029), .B(n7916), .Z(n7914) );
  NANDN U8158 ( .A(n7917), .B(n7918), .Z(n7916) );
  NAND U8159 ( .A(n7033), .B(\stack[5][17] ), .Z(n7918) );
  NAND U8160 ( .A(n7919), .B(n7920), .Z(n2289) );
  NAND U8161 ( .A(n7028), .B(\stack[6][18] ), .Z(n7920) );
  NAND U8162 ( .A(n7029), .B(n7921), .Z(n7919) );
  NANDN U8163 ( .A(n7922), .B(n7923), .Z(n7921) );
  NAND U8164 ( .A(n7033), .B(\stack[5][18] ), .Z(n7923) );
  NAND U8165 ( .A(n7924), .B(n7925), .Z(n2288) );
  NAND U8166 ( .A(n7028), .B(\stack[6][19] ), .Z(n7925) );
  NAND U8167 ( .A(n7029), .B(n7926), .Z(n7924) );
  NANDN U8168 ( .A(n7927), .B(n7928), .Z(n7926) );
  NAND U8169 ( .A(n7033), .B(\stack[5][19] ), .Z(n7928) );
  NAND U8170 ( .A(n7929), .B(n7930), .Z(n2287) );
  NAND U8171 ( .A(n7028), .B(\stack[6][20] ), .Z(n7930) );
  NAND U8172 ( .A(n7029), .B(n7931), .Z(n7929) );
  NANDN U8173 ( .A(n7932), .B(n7933), .Z(n7931) );
  NAND U8174 ( .A(n7033), .B(\stack[5][20] ), .Z(n7933) );
  NAND U8175 ( .A(n7934), .B(n7935), .Z(n2286) );
  NAND U8176 ( .A(n7028), .B(\stack[6][21] ), .Z(n7935) );
  NAND U8177 ( .A(n7029), .B(n7936), .Z(n7934) );
  NANDN U8178 ( .A(n7937), .B(n7938), .Z(n7936) );
  NAND U8179 ( .A(n7033), .B(\stack[5][21] ), .Z(n7938) );
  NAND U8180 ( .A(n7939), .B(n7940), .Z(n2285) );
  NAND U8181 ( .A(n7028), .B(\stack[6][22] ), .Z(n7940) );
  NAND U8182 ( .A(n7029), .B(n7941), .Z(n7939) );
  NANDN U8183 ( .A(n7942), .B(n7943), .Z(n7941) );
  NAND U8184 ( .A(n7033), .B(\stack[5][22] ), .Z(n7943) );
  NAND U8185 ( .A(n7944), .B(n7945), .Z(n2284) );
  NAND U8186 ( .A(n7028), .B(\stack[6][23] ), .Z(n7945) );
  NAND U8187 ( .A(n7029), .B(n7946), .Z(n7944) );
  NANDN U8188 ( .A(n7947), .B(n7948), .Z(n7946) );
  NAND U8189 ( .A(n7033), .B(\stack[5][23] ), .Z(n7948) );
  NAND U8190 ( .A(n7949), .B(n7950), .Z(n2283) );
  NAND U8191 ( .A(n7028), .B(\stack[6][24] ), .Z(n7950) );
  NAND U8192 ( .A(n7029), .B(n7951), .Z(n7949) );
  NANDN U8193 ( .A(n7952), .B(n7953), .Z(n7951) );
  NAND U8194 ( .A(n7033), .B(\stack[5][24] ), .Z(n7953) );
  NAND U8195 ( .A(n7954), .B(n7955), .Z(n2282) );
  NAND U8196 ( .A(n7028), .B(\stack[6][25] ), .Z(n7955) );
  NAND U8197 ( .A(n7029), .B(n7956), .Z(n7954) );
  NANDN U8198 ( .A(n7957), .B(n7958), .Z(n7956) );
  NAND U8199 ( .A(n7033), .B(\stack[5][25] ), .Z(n7958) );
  NAND U8200 ( .A(n7959), .B(n7960), .Z(n2281) );
  NAND U8201 ( .A(n7028), .B(\stack[6][26] ), .Z(n7960) );
  NAND U8202 ( .A(n7029), .B(n7961), .Z(n7959) );
  NANDN U8203 ( .A(n7962), .B(n7963), .Z(n7961) );
  NAND U8204 ( .A(n7033), .B(\stack[5][26] ), .Z(n7963) );
  NAND U8205 ( .A(n7964), .B(n7965), .Z(n2280) );
  NAND U8206 ( .A(n7028), .B(\stack[6][27] ), .Z(n7965) );
  NAND U8207 ( .A(n7029), .B(n7966), .Z(n7964) );
  NANDN U8208 ( .A(n7967), .B(n7968), .Z(n7966) );
  NAND U8209 ( .A(n7033), .B(\stack[5][27] ), .Z(n7968) );
  NAND U8210 ( .A(n7969), .B(n7970), .Z(n2279) );
  NAND U8211 ( .A(n7028), .B(\stack[6][28] ), .Z(n7970) );
  NAND U8212 ( .A(n7029), .B(n7971), .Z(n7969) );
  NANDN U8213 ( .A(n7972), .B(n7973), .Z(n7971) );
  NAND U8214 ( .A(n7033), .B(\stack[5][28] ), .Z(n7973) );
  NAND U8215 ( .A(n7974), .B(n7975), .Z(n2278) );
  NAND U8216 ( .A(n7028), .B(\stack[6][29] ), .Z(n7975) );
  NAND U8217 ( .A(n7029), .B(n7976), .Z(n7974) );
  NANDN U8218 ( .A(n7977), .B(n7978), .Z(n7976) );
  NAND U8219 ( .A(n7033), .B(\stack[5][29] ), .Z(n7978) );
  NAND U8220 ( .A(n7979), .B(n7980), .Z(n2277) );
  NAND U8221 ( .A(n7028), .B(\stack[6][30] ), .Z(n7980) );
  NAND U8222 ( .A(n7029), .B(n7981), .Z(n7979) );
  NANDN U8223 ( .A(n7982), .B(n7983), .Z(n7981) );
  NAND U8224 ( .A(n7033), .B(\stack[5][30] ), .Z(n7983) );
  NAND U8225 ( .A(n7984), .B(n7985), .Z(n2276) );
  NAND U8226 ( .A(n7028), .B(\stack[6][31] ), .Z(n7985) );
  NAND U8227 ( .A(n7029), .B(n7986), .Z(n7984) );
  NANDN U8228 ( .A(n7987), .B(n7988), .Z(n7986) );
  NAND U8229 ( .A(n7033), .B(\stack[5][31] ), .Z(n7988) );
  IV U8230 ( .A(n7028), .Z(n7029) );
  ANDN U8231 ( .B(n2503), .A(n3337), .Z(n7028) );
  NAND U8232 ( .A(n7989), .B(n7990), .Z(n3337) );
  NOR U8233 ( .A(n2607), .B(n6683), .Z(n7990) );
  NOR U8234 ( .A(opcode[0]), .B(n7991), .Z(n6683) );
  ANDN U8235 ( .B(opcode[0]), .A(n7991), .Z(n2607) );
  NAND U8236 ( .A(n7992), .B(opcode[1]), .Z(n7991) );
  ANDN U8237 ( .B(n6669), .A(n6682), .Z(n7989) );
  ANDN U8238 ( .B(n7993), .A(n6667), .Z(n6682) );
  AND U8239 ( .A(n6672), .B(n7992), .Z(n7993) );
  NAND U8240 ( .A(opcode[2]), .B(opcode[1]), .Z(n6669) );
  IV U8241 ( .A(n7033), .Z(n2503) );
  NANDN U8242 ( .A(n7837), .B(n7994), .Z(n2264) );
  NAND U8243 ( .A(n7033), .B(\stack[6][1] ), .Z(n7994) );
  ANDN U8244 ( .B(\stack[7][1] ), .A(n7033), .Z(n7837) );
  NANDN U8245 ( .A(n7842), .B(n7995), .Z(n2255) );
  NAND U8246 ( .A(n7033), .B(\stack[6][2] ), .Z(n7995) );
  ANDN U8247 ( .B(\stack[7][2] ), .A(n7033), .Z(n7842) );
  NANDN U8248 ( .A(n7847), .B(n7996), .Z(n2246) );
  NAND U8249 ( .A(n7033), .B(\stack[6][3] ), .Z(n7996) );
  ANDN U8250 ( .B(\stack[7][3] ), .A(n7033), .Z(n7847) );
  NANDN U8251 ( .A(n7852), .B(n7997), .Z(n2237) );
  NAND U8252 ( .A(n7033), .B(\stack[6][4] ), .Z(n7997) );
  ANDN U8253 ( .B(\stack[7][4] ), .A(n7033), .Z(n7852) );
  NANDN U8254 ( .A(n7857), .B(n7998), .Z(n2228) );
  NAND U8255 ( .A(n7033), .B(\stack[6][5] ), .Z(n7998) );
  ANDN U8256 ( .B(\stack[7][5] ), .A(n7033), .Z(n7857) );
  NANDN U8257 ( .A(n7862), .B(n7999), .Z(n2219) );
  NAND U8258 ( .A(n7033), .B(\stack[6][6] ), .Z(n7999) );
  ANDN U8259 ( .B(\stack[7][6] ), .A(n7033), .Z(n7862) );
  NANDN U8260 ( .A(n7867), .B(n8000), .Z(n2210) );
  NAND U8261 ( .A(n7033), .B(\stack[6][7] ), .Z(n8000) );
  ANDN U8262 ( .B(\stack[7][7] ), .A(n7033), .Z(n7867) );
  NANDN U8263 ( .A(n7872), .B(n8001), .Z(n2201) );
  NAND U8264 ( .A(n7033), .B(\stack[6][8] ), .Z(n8001) );
  ANDN U8265 ( .B(\stack[7][8] ), .A(n7033), .Z(n7872) );
  NANDN U8266 ( .A(n7877), .B(n8002), .Z(n2192) );
  NAND U8267 ( .A(n7033), .B(\stack[6][9] ), .Z(n8002) );
  ANDN U8268 ( .B(\stack[7][9] ), .A(n7033), .Z(n7877) );
  NANDN U8269 ( .A(n7882), .B(n8003), .Z(n2183) );
  NAND U8270 ( .A(n7033), .B(\stack[6][10] ), .Z(n8003) );
  ANDN U8271 ( .B(\stack[7][10] ), .A(n7033), .Z(n7882) );
  NANDN U8272 ( .A(n7887), .B(n8004), .Z(n2174) );
  NAND U8273 ( .A(n7033), .B(\stack[6][11] ), .Z(n8004) );
  ANDN U8274 ( .B(\stack[7][11] ), .A(n7033), .Z(n7887) );
  NANDN U8275 ( .A(n7892), .B(n8005), .Z(n2165) );
  NAND U8276 ( .A(n7033), .B(\stack[6][12] ), .Z(n8005) );
  ANDN U8277 ( .B(\stack[7][12] ), .A(n7033), .Z(n7892) );
  NANDN U8278 ( .A(n7897), .B(n8006), .Z(n2156) );
  NAND U8279 ( .A(n7033), .B(\stack[6][13] ), .Z(n8006) );
  ANDN U8280 ( .B(\stack[7][13] ), .A(n7033), .Z(n7897) );
  NANDN U8281 ( .A(n7902), .B(n8007), .Z(n2147) );
  NAND U8282 ( .A(n7033), .B(\stack[6][14] ), .Z(n8007) );
  ANDN U8283 ( .B(\stack[7][14] ), .A(n7033), .Z(n7902) );
  NANDN U8284 ( .A(n7907), .B(n8008), .Z(n2138) );
  NAND U8285 ( .A(n7033), .B(\stack[6][15] ), .Z(n8008) );
  ANDN U8286 ( .B(\stack[7][15] ), .A(n7033), .Z(n7907) );
  NANDN U8287 ( .A(n7912), .B(n8009), .Z(n2129) );
  NAND U8288 ( .A(n7033), .B(\stack[6][16] ), .Z(n8009) );
  ANDN U8289 ( .B(\stack[7][16] ), .A(n7033), .Z(n7912) );
  NANDN U8290 ( .A(n7917), .B(n8010), .Z(n2120) );
  NAND U8291 ( .A(n7033), .B(\stack[6][17] ), .Z(n8010) );
  ANDN U8292 ( .B(\stack[7][17] ), .A(n7033), .Z(n7917) );
  NANDN U8293 ( .A(n7922), .B(n8011), .Z(n2111) );
  NAND U8294 ( .A(n7033), .B(\stack[6][18] ), .Z(n8011) );
  ANDN U8295 ( .B(\stack[7][18] ), .A(n7033), .Z(n7922) );
  NANDN U8296 ( .A(n7927), .B(n8012), .Z(n2102) );
  NAND U8297 ( .A(n7033), .B(\stack[6][19] ), .Z(n8012) );
  ANDN U8298 ( .B(\stack[7][19] ), .A(n7033), .Z(n7927) );
  NANDN U8299 ( .A(n7932), .B(n8013), .Z(n2093) );
  NAND U8300 ( .A(n7033), .B(\stack[6][20] ), .Z(n8013) );
  ANDN U8301 ( .B(\stack[7][20] ), .A(n7033), .Z(n7932) );
  NANDN U8302 ( .A(n7937), .B(n8014), .Z(n2084) );
  NAND U8303 ( .A(n7033), .B(\stack[6][21] ), .Z(n8014) );
  ANDN U8304 ( .B(\stack[7][21] ), .A(n7033), .Z(n7937) );
  NANDN U8305 ( .A(n7942), .B(n8015), .Z(n2075) );
  NAND U8306 ( .A(n7033), .B(\stack[6][22] ), .Z(n8015) );
  ANDN U8307 ( .B(\stack[7][22] ), .A(n7033), .Z(n7942) );
  NANDN U8308 ( .A(n7947), .B(n8016), .Z(n2066) );
  NAND U8309 ( .A(n7033), .B(\stack[6][23] ), .Z(n8016) );
  ANDN U8310 ( .B(\stack[7][23] ), .A(n7033), .Z(n7947) );
  NANDN U8311 ( .A(n7952), .B(n8017), .Z(n2057) );
  NAND U8312 ( .A(n7033), .B(\stack[6][24] ), .Z(n8017) );
  ANDN U8313 ( .B(\stack[7][24] ), .A(n7033), .Z(n7952) );
  NANDN U8314 ( .A(n7957), .B(n8018), .Z(n2048) );
  NAND U8315 ( .A(n7033), .B(\stack[6][25] ), .Z(n8018) );
  ANDN U8316 ( .B(\stack[7][25] ), .A(n7033), .Z(n7957) );
  NANDN U8317 ( .A(n7962), .B(n8019), .Z(n2039) );
  NAND U8318 ( .A(n7033), .B(\stack[6][26] ), .Z(n8019) );
  ANDN U8319 ( .B(\stack[7][26] ), .A(n7033), .Z(n7962) );
  NANDN U8320 ( .A(n7967), .B(n8020), .Z(n2030) );
  NAND U8321 ( .A(n7033), .B(\stack[6][27] ), .Z(n8020) );
  ANDN U8322 ( .B(\stack[7][27] ), .A(n7033), .Z(n7967) );
  NANDN U8323 ( .A(n7972), .B(n8021), .Z(n2021) );
  NAND U8324 ( .A(n7033), .B(\stack[6][28] ), .Z(n8021) );
  ANDN U8325 ( .B(\stack[7][28] ), .A(n7033), .Z(n7972) );
  NANDN U8326 ( .A(n7977), .B(n8022), .Z(n2012) );
  NAND U8327 ( .A(n7033), .B(\stack[6][29] ), .Z(n8022) );
  ANDN U8328 ( .B(\stack[7][29] ), .A(n7033), .Z(n7977) );
  NANDN U8329 ( .A(n7982), .B(n8023), .Z(n2003) );
  NAND U8330 ( .A(n7033), .B(\stack[6][30] ), .Z(n8023) );
  ANDN U8331 ( .B(\stack[7][30] ), .A(n7033), .Z(n7982) );
  NANDN U8332 ( .A(n7987), .B(n8024), .Z(n1996) );
  NAND U8333 ( .A(n7033), .B(\stack[6][31] ), .Z(n8024) );
  ANDN U8334 ( .B(\stack[7][31] ), .A(n7033), .Z(n7987) );
  NANDN U8335 ( .A(n7832), .B(n8025), .Z(n1989) );
  NAND U8336 ( .A(n7033), .B(\stack[6][0] ), .Z(n8025) );
  ANDN U8337 ( .B(\stack[7][0] ), .A(n7033), .Z(n7832) );
  ANDN U8338 ( .B(n8026), .A(n7992), .Z(n7033) );
  IV U8339 ( .A(opcode[2]), .Z(n7992) );
  AND U8340 ( .A(n6667), .B(n6672), .Z(n8026) );
  IV U8341 ( .A(opcode[1]), .Z(n6672) );
  IV U8342 ( .A(opcode[0]), .Z(n6667) );
endmodule

