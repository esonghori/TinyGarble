
module compare_N16384_CC16 ( clk, rst, x, y, g, e );
  input [1023:0] x;
  input [1023:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NANDN U10 ( .A(x[266]), .B(y[266]), .Z(n8) );
  NAND U11 ( .A(n8), .B(n509), .Z(n4811) );
  NANDN U12 ( .A(x[758]), .B(y[758]), .Z(n9) );
  NAND U13 ( .A(n9), .B(n2338), .Z(n5810) );
  NANDN U14 ( .A(x[86]), .B(y[86]), .Z(n10) );
  NAND U15 ( .A(n10), .B(n614), .Z(n4420) );
  NANDN U16 ( .A(x[128]), .B(y[128]), .Z(n11) );
  NANDN U17 ( .A(n582), .B(n11), .Z(n3221) );
  NANDN U18 ( .A(n4839), .B(n4838), .Z(n12) );
  NAND U19 ( .A(n12), .B(n4840), .Z(n13) );
  NANDN U20 ( .A(n4841), .B(n13), .Z(n14) );
  NAND U21 ( .A(n14), .B(n4842), .Z(n15) );
  NANDN U22 ( .A(n4843), .B(n15), .Z(n16) );
  AND U23 ( .A(n4844), .B(n16), .Z(n17) );
  OR U24 ( .A(n4845), .B(n17), .Z(n18) );
  ANDN U25 ( .B(n18), .A(n4846), .Z(n19) );
  NANDN U26 ( .A(y[286]), .B(x[286]), .Z(n20) );
  NANDN U27 ( .A(n19), .B(n20), .Z(n21) );
  ANDN U28 ( .B(n21), .A(n4847), .Z(n22) );
  OR U29 ( .A(n4848), .B(n22), .Z(n23) );
  NAND U30 ( .A(n23), .B(n4849), .Z(n24) );
  ANDN U31 ( .B(n24), .A(n4850), .Z(n25) );
  NANDN U32 ( .A(n25), .B(n4851), .Z(n26) );
  ANDN U33 ( .B(n26), .A(n4852), .Z(n27) );
  NANDN U34 ( .A(n27), .B(n4853), .Z(n28) );
  NANDN U35 ( .A(n4854), .B(n28), .Z(n29) );
  NAND U36 ( .A(n29), .B(n4369), .Z(n4855) );
  NANDN U37 ( .A(x[448]), .B(y[448]), .Z(n30) );
  NAND U38 ( .A(n30), .B(n1636), .Z(n3626) );
  NANDN U39 ( .A(x[462]), .B(y[462]), .Z(n31) );
  NAND U40 ( .A(n31), .B(n1661), .Z(n5200) );
  NANDN U41 ( .A(x[746]), .B(y[746]), .Z(n32) );
  NAND U42 ( .A(n32), .B(n2315), .Z(n5779) );
  NANDN U43 ( .A(x[771]), .B(y[771]), .Z(n33) );
  XNOR U44 ( .A(x[771]), .B(y[771]), .Z(n34) );
  NANDN U45 ( .A(y[770]), .B(x[770]), .Z(n35) );
  NAND U46 ( .A(n34), .B(n35), .Z(n36) );
  NAND U47 ( .A(n33), .B(n36), .Z(n5835) );
  NANDN U48 ( .A(x[802]), .B(y[802]), .Z(n37) );
  NAND U49 ( .A(n37), .B(n2434), .Z(n4035) );
  NANDN U50 ( .A(x[781]), .B(y[781]), .Z(n38) );
  XNOR U51 ( .A(x[781]), .B(y[781]), .Z(n39) );
  NANDN U52 ( .A(y[780]), .B(x[780]), .Z(n40) );
  NAND U53 ( .A(n39), .B(n40), .Z(n41) );
  NAND U54 ( .A(n38), .B(n41), .Z(n5859) );
  NANDN U55 ( .A(x[806]), .B(y[806]), .Z(n42) );
  NAND U56 ( .A(n42), .B(n2440), .Z(n5916) );
  NANDN U57 ( .A(x[1]), .B(y[1]), .Z(n2986) );
  NANDN U58 ( .A(x[68]), .B(y[68]), .Z(n43) );
  AND U59 ( .A(n627), .B(n43), .Z(n4379) );
  NANDN U60 ( .A(x[100]), .B(y[100]), .Z(n44) );
  NAND U61 ( .A(n44), .B(n881), .Z(n4452) );
  NANDN U62 ( .A(x[112]), .B(y[112]), .Z(n45) );
  NAND U63 ( .A(n45), .B(n591), .Z(n4478) );
  NANDN U64 ( .A(x[124]), .B(y[124]), .Z(n46) );
  NAND U65 ( .A(n46), .B(n925), .Z(n4506) );
  NANDN U66 ( .A(x[140]), .B(y[140]), .Z(n47) );
  NAND U67 ( .A(n47), .B(n574), .Z(n3241) );
  NANDN U68 ( .A(x[162]), .B(y[162]), .Z(n48) );
  NANDN U69 ( .A(n996), .B(n48), .Z(n3272) );
  NANDN U70 ( .A(x[178]), .B(y[178]), .Z(n49) );
  NAND U71 ( .A(n49), .B(n557), .Z(n3297) );
  NANDN U72 ( .A(x[200]), .B(y[200]), .Z(n50) );
  NANDN U73 ( .A(n1089), .B(n50), .Z(n3325) );
  NANDN U74 ( .A(x[230]), .B(y[230]), .Z(n51) );
  NAND U75 ( .A(n51), .B(n534), .Z(n4735) );
  NANDN U76 ( .A(x[242]), .B(y[242]), .Z(n52) );
  NANDN U77 ( .A(n526), .B(n52), .Z(n3375) );
  NANDN U78 ( .A(x[286]), .B(y[286]), .Z(n53) );
  NAND U79 ( .A(n53), .B(n495), .Z(n4847) );
  NANDN U80 ( .A(x[274]), .B(y[274]), .Z(n54) );
  NAND U81 ( .A(n54), .B(n503), .Z(n4371) );
  NANDN U82 ( .A(x[312]), .B(y[312]), .Z(n55) );
  NAND U83 ( .A(n55), .B(n1319), .Z(n3466) );
  NANDN U84 ( .A(x[330]), .B(y[330]), .Z(n56) );
  NAND U85 ( .A(n56), .B(n464), .Z(n3488) );
  NANDN U86 ( .A(x[294]), .B(y[294]), .Z(n57) );
  AND U87 ( .A(n4369), .B(n57), .Z(n3434) );
  NANDN U88 ( .A(x[350]), .B(y[350]), .Z(n58) );
  NAND U89 ( .A(n58), .B(n1407), .Z(n4972) );
  NANDN U90 ( .A(x[358]), .B(y[358]), .Z(n59) );
  NAND U91 ( .A(n59), .B(n446), .Z(n4992) );
  NANDN U92 ( .A(x[406]), .B(y[406]), .Z(n60) );
  NAND U93 ( .A(n60), .B(n1527), .Z(n3578) );
  NANDN U94 ( .A(x[455]), .B(y[455]), .Z(n61) );
  XNOR U95 ( .A(x[455]), .B(y[455]), .Z(n62) );
  NANDN U96 ( .A(y[454]), .B(x[454]), .Z(n63) );
  NAND U97 ( .A(n62), .B(n63), .Z(n64) );
  NAND U98 ( .A(n61), .B(n64), .Z(n5185) );
  NANDN U99 ( .A(x[532]), .B(y[532]), .Z(n65) );
  NAND U100 ( .A(n65), .B(n345), .Z(n5344) );
  NANDN U101 ( .A(x[556]), .B(y[556]), .Z(n66) );
  NAND U102 ( .A(n66), .B(n329), .Z(n5396) );
  NANDN U103 ( .A(x[569]), .B(y[569]), .Z(n67) );
  XNOR U104 ( .A(x[569]), .B(y[569]), .Z(n68) );
  NANDN U105 ( .A(y[568]), .B(x[568]), .Z(n69) );
  NAND U106 ( .A(n68), .B(n69), .Z(n70) );
  NAND U107 ( .A(n67), .B(n70), .Z(n5417) );
  NANDN U108 ( .A(x[588]), .B(y[588]), .Z(n71) );
  NAND U109 ( .A(n71), .B(n306), .Z(n5460) );
  NANDN U110 ( .A(x[676]), .B(y[676]), .Z(n72) );
  NAND U111 ( .A(n72), .B(n2151), .Z(n3891) );
  NANDN U112 ( .A(x[720]), .B(y[720]), .Z(n73) );
  NAND U113 ( .A(n73), .B(n2264), .Z(n5726) );
  NANDN U114 ( .A(y[730]), .B(x[730]), .Z(n74) );
  NANDN U115 ( .A(x[731]), .B(y[731]), .Z(n75) );
  XNOR U116 ( .A(x[731]), .B(y[731]), .Z(n76) );
  NAND U117 ( .A(n76), .B(n74), .Z(n77) );
  NAND U118 ( .A(n75), .B(n77), .Z(n5743) );
  NANDN U119 ( .A(x[754]), .B(y[754]), .Z(n78) );
  NAND U120 ( .A(n78), .B(n221), .Z(n5798) );
  NANDN U121 ( .A(x[772]), .B(y[772]), .Z(n79) );
  AND U122 ( .A(n2369), .B(n79), .Z(n5839) );
  NANDN U123 ( .A(x[782]), .B(y[782]), .Z(n80) );
  AND U124 ( .A(n202), .B(n80), .Z(n5861) );
  NANDN U125 ( .A(x[808]), .B(y[808]), .Z(n81) );
  AND U126 ( .A(n2443), .B(n81), .Z(n5913) );
  OR U127 ( .A(x[862]), .B(n2920), .Z(n4114) );
  NANDN U128 ( .A(y[870]), .B(x[870]), .Z(n82) );
  AND U129 ( .A(n167), .B(n82), .Z(n6055) );
  NANDN U130 ( .A(y[882]), .B(x[882]), .Z(n83) );
  AND U131 ( .A(n2617), .B(n83), .Z(n6083) );
  NANDN U132 ( .A(x[990]), .B(y[990]), .Z(n4361) );
  IV U133 ( .A(ebreg), .Z(e) );
  NANDN U134 ( .A(x[1023]), .B(y[1023]), .Z(n6426) );
  NANDN U135 ( .A(x[1019]), .B(y[1019]), .Z(n85) );
  NANDN U136 ( .A(x[1020]), .B(y[1020]), .Z(n84) );
  NAND U137 ( .A(n85), .B(n84), .Z(n6418) );
  NANDN U138 ( .A(y[1014]), .B(x[1014]), .Z(n2898) );
  NANDN U139 ( .A(y[1016]), .B(x[1016]), .Z(n87) );
  NANDN U140 ( .A(y[1017]), .B(x[1017]), .Z(n86) );
  NAND U141 ( .A(n87), .B(n86), .Z(n6412) );
  NANDN U142 ( .A(x[1015]), .B(y[1015]), .Z(n89) );
  NANDN U143 ( .A(x[1016]), .B(y[1016]), .Z(n88) );
  NAND U144 ( .A(n89), .B(n88), .Z(n6409) );
  NOR U145 ( .A(n6412), .B(n6409), .Z(n90) );
  AND U146 ( .A(n2898), .B(n90), .Z(n91) );
  NANDN U147 ( .A(n6418), .B(n91), .Z(n94) );
  NANDN U148 ( .A(x[1021]), .B(y[1021]), .Z(n93) );
  NANDN U149 ( .A(x[1022]), .B(y[1022]), .Z(n92) );
  NAND U150 ( .A(n93), .B(n92), .Z(n6421) );
  NOR U151 ( .A(n94), .B(n6421), .Z(n95) );
  AND U152 ( .A(n6426), .B(n95), .Z(n96) );
  NANDN U153 ( .A(y[1015]), .B(x[1015]), .Z(n2899) );
  NAND U154 ( .A(n96), .B(n2899), .Z(n108) );
  NANDN U155 ( .A(y[1022]), .B(x[1022]), .Z(n98) );
  NANDN U156 ( .A(y[1023]), .B(x[1023]), .Z(n97) );
  NAND U157 ( .A(n98), .B(n97), .Z(n6424) );
  NANDN U158 ( .A(x[1017]), .B(y[1017]), .Z(n100) );
  NANDN U159 ( .A(x[1018]), .B(y[1018]), .Z(n99) );
  NAND U160 ( .A(n100), .B(n99), .Z(n6414) );
  NANDN U161 ( .A(y[1018]), .B(x[1018]), .Z(n102) );
  NANDN U162 ( .A(y[1019]), .B(x[1019]), .Z(n101) );
  NAND U163 ( .A(n102), .B(n101), .Z(n6416) );
  NOR U164 ( .A(n6414), .B(n6416), .Z(n105) );
  NANDN U165 ( .A(y[1020]), .B(x[1020]), .Z(n104) );
  NANDN U166 ( .A(y[1021]), .B(x[1021]), .Z(n103) );
  NAND U167 ( .A(n104), .B(n103), .Z(n6420) );
  ANDN U168 ( .B(n105), .A(n6420), .Z(n106) );
  NANDN U169 ( .A(n6424), .B(n106), .Z(n107) );
  NOR U170 ( .A(n108), .B(n107), .Z(n2902) );
  NANDN U171 ( .A(y[1010]), .B(x[1010]), .Z(n110) );
  NANDN U172 ( .A(y[1011]), .B(x[1011]), .Z(n109) );
  AND U173 ( .A(n110), .B(n109), .Z(n6399) );
  NANDN U174 ( .A(x[1008]), .B(y[1008]), .Z(n6393) );
  NANDN U175 ( .A(x[1004]), .B(y[1004]), .Z(n6381) );
  NANDN U176 ( .A(x[1005]), .B(y[1005]), .Z(n6386) );
  NAND U177 ( .A(n6381), .B(n6386), .Z(n2879) );
  ANDN U178 ( .B(y[1002]), .A(x[1002]), .Z(n6373) );
  ANDN U179 ( .B(y[1003]), .A(x[1003]), .Z(n6379) );
  OR U180 ( .A(n6373), .B(n6379), .Z(n4331) );
  NANDN U181 ( .A(y[999]), .B(x[999]), .Z(n112) );
  NANDN U182 ( .A(y[998]), .B(x[998]), .Z(n111) );
  NAND U183 ( .A(n112), .B(n111), .Z(n6368) );
  NANDN U184 ( .A(x[994]), .B(y[994]), .Z(n4318) );
  NANDN U185 ( .A(x[995]), .B(y[995]), .Z(n4321) );
  NAND U186 ( .A(n4318), .B(n4321), .Z(n6358) );
  NANDN U187 ( .A(x[992]), .B(y[992]), .Z(n113) );
  NANDN U188 ( .A(x[993]), .B(y[993]), .Z(n2908) );
  NAND U189 ( .A(n113), .B(n2908), .Z(n4310) );
  NANDN U190 ( .A(y[992]), .B(x[992]), .Z(n2907) );
  ANDN U191 ( .B(y[991]), .A(x[991]), .Z(n4311) );
  ANDN U192 ( .B(n4361), .A(n4311), .Z(n2856) );
  NANDN U193 ( .A(x[989]), .B(y[989]), .Z(n4303) );
  IV U194 ( .A(n4303), .Z(n4360) );
  NANDN U195 ( .A(x[986]), .B(y[986]), .Z(n115) );
  NANDN U196 ( .A(x[985]), .B(y[985]), .Z(n114) );
  NAND U197 ( .A(n115), .B(n114), .Z(n6340) );
  ANDN U198 ( .B(y[983]), .A(x[983]), .Z(n4295) );
  ANDN U199 ( .B(y[982]), .A(x[982]), .Z(n4290) );
  NOR U200 ( .A(n4295), .B(n4290), .Z(n6331) );
  NANDN U201 ( .A(y[981]), .B(x[981]), .Z(n116) );
  NANDN U202 ( .A(y[982]), .B(x[982]), .Z(n4293) );
  NAND U203 ( .A(n116), .B(n4293), .Z(n6330) );
  NANDN U204 ( .A(x[980]), .B(y[980]), .Z(n4282) );
  NANDN U205 ( .A(x[981]), .B(y[981]), .Z(n117) );
  NAND U206 ( .A(n4282), .B(n117), .Z(n6328) );
  ANDN U207 ( .B(y[979]), .A(x[979]), .Z(n6324) );
  ANDN U208 ( .B(x[979]), .A(y[979]), .Z(n2830) );
  ANDN U209 ( .B(y[978]), .A(x[978]), .Z(n6320) );
  NANDN U210 ( .A(n2830), .B(n6320), .Z(n118) );
  NANDN U211 ( .A(n6324), .B(n118), .Z(n4284) );
  NANDN U212 ( .A(x[977]), .B(y[977]), .Z(n6318) );
  NANDN U213 ( .A(x[972]), .B(y[972]), .Z(n6305) );
  NANDN U214 ( .A(x[966]), .B(y[966]), .Z(n120) );
  NANDN U215 ( .A(x[967]), .B(y[967]), .Z(n119) );
  AND U216 ( .A(n120), .B(n119), .Z(n6293) );
  NANDN U217 ( .A(x[961]), .B(y[961]), .Z(n122) );
  NANDN U218 ( .A(x[962]), .B(y[962]), .Z(n121) );
  AND U219 ( .A(n122), .B(n121), .Z(n6281) );
  NANDN U220 ( .A(x[956]), .B(y[956]), .Z(n124) );
  NANDN U221 ( .A(x[957]), .B(y[957]), .Z(n123) );
  AND U222 ( .A(n124), .B(n123), .Z(n6269) );
  NANDN U223 ( .A(x[951]), .B(y[951]), .Z(n126) );
  NANDN U224 ( .A(x[952]), .B(y[952]), .Z(n125) );
  AND U225 ( .A(n126), .B(n125), .Z(n6257) );
  NANDN U226 ( .A(y[945]), .B(x[945]), .Z(n4237) );
  IV U227 ( .A(x[946]), .Z(n2913) );
  IV U228 ( .A(y[946]), .Z(n2912) );
  NANDN U229 ( .A(n2913), .B(n2912), .Z(n127) );
  NAND U230 ( .A(n4237), .B(n127), .Z(n6244) );
  NANDN U231 ( .A(x[944]), .B(y[944]), .Z(n129) );
  NANDN U232 ( .A(x[943]), .B(y[943]), .Z(n128) );
  NAND U233 ( .A(n129), .B(n128), .Z(n6238) );
  ANDN U234 ( .B(x[943]), .A(y[943]), .Z(n2743) );
  ANDN U235 ( .B(y[942]), .A(x[942]), .Z(n6231) );
  NANDN U236 ( .A(n2743), .B(n6231), .Z(n130) );
  NANDN U237 ( .A(n6238), .B(n130), .Z(n4234) );
  NANDN U238 ( .A(x[941]), .B(y[941]), .Z(n6232) );
  NANDN U239 ( .A(x[940]), .B(y[940]), .Z(n132) );
  NANDN U240 ( .A(x[939]), .B(y[939]), .Z(n131) );
  NAND U241 ( .A(n132), .B(n131), .Z(n6228) );
  NANDN U242 ( .A(x[938]), .B(y[938]), .Z(n134) );
  NANDN U243 ( .A(x[937]), .B(y[937]), .Z(n133) );
  NAND U244 ( .A(n134), .B(n133), .Z(n6224) );
  NANDN U245 ( .A(x[936]), .B(y[936]), .Z(n6219) );
  NANDN U246 ( .A(y[933]), .B(x[933]), .Z(n2914) );
  NANDN U247 ( .A(x[932]), .B(y[932]), .Z(n6207) );
  NANDN U248 ( .A(x[933]), .B(y[933]), .Z(n6211) );
  AND U249 ( .A(n6207), .B(n6211), .Z(n2725) );
  NANDN U250 ( .A(x[931]), .B(y[931]), .Z(n6203) );
  NANDN U251 ( .A(x[930]), .B(y[930]), .Z(n135) );
  NAND U252 ( .A(n6203), .B(n135), .Z(n6199) );
  ANDN U253 ( .B(x[931]), .A(y[931]), .Z(n2719) );
  ANDN U254 ( .B(n6199), .A(n2719), .Z(n4217) );
  NANDN U255 ( .A(x[929]), .B(y[929]), .Z(n6201) );
  NANDN U256 ( .A(y[925]), .B(x[925]), .Z(n137) );
  NANDN U257 ( .A(y[924]), .B(x[924]), .Z(n136) );
  NAND U258 ( .A(n137), .B(n136), .Z(n6189) );
  NANDN U259 ( .A(x[922]), .B(y[922]), .Z(n4202) );
  NANDN U260 ( .A(x[923]), .B(y[923]), .Z(n4206) );
  NAND U261 ( .A(n4202), .B(n4206), .Z(n6184) );
  ANDN U262 ( .B(x[920]), .A(y[920]), .Z(n6177) );
  NANDN U263 ( .A(y[919]), .B(x[919]), .Z(n138) );
  NANDN U264 ( .A(n6177), .B(n138), .Z(n4199) );
  NANDN U265 ( .A(y[916]), .B(x[916]), .Z(n140) );
  NANDN U266 ( .A(y[917]), .B(x[917]), .Z(n139) );
  AND U267 ( .A(n140), .B(n139), .Z(n6165) );
  NANDN U268 ( .A(y[911]), .B(x[911]), .Z(n6153) );
  NANDN U269 ( .A(y[907]), .B(x[907]), .Z(n141) );
  NANDN U270 ( .A(y[908]), .B(x[908]), .Z(n6144) );
  NAND U271 ( .A(n141), .B(n6144), .Z(n2666) );
  NANDN U272 ( .A(y[906]), .B(x[906]), .Z(n142) );
  NANDN U273 ( .A(n2666), .B(n142), .Z(n6142) );
  NANDN U274 ( .A(y[903]), .B(x[903]), .Z(n144) );
  NANDN U275 ( .A(y[902]), .B(x[902]), .Z(n143) );
  NAND U276 ( .A(n144), .B(n143), .Z(n6132) );
  NANDN U277 ( .A(y[901]), .B(x[901]), .Z(n146) );
  NANDN U278 ( .A(y[900]), .B(x[900]), .Z(n145) );
  NAND U279 ( .A(n146), .B(n145), .Z(n6127) );
  NANDN U280 ( .A(y[899]), .B(x[899]), .Z(n6123) );
  NANDN U281 ( .A(y[898]), .B(x[898]), .Z(n148) );
  NANDN U282 ( .A(y[897]), .B(x[897]), .Z(n147) );
  NAND U283 ( .A(n148), .B(n147), .Z(n6120) );
  NANDN U284 ( .A(y[896]), .B(x[896]), .Z(n150) );
  NANDN U285 ( .A(y[895]), .B(x[895]), .Z(n149) );
  NAND U286 ( .A(n150), .B(n149), .Z(n6115) );
  NANDN U287 ( .A(y[894]), .B(x[894]), .Z(n6111) );
  NANDN U288 ( .A(y[892]), .B(x[892]), .Z(n152) );
  NANDN U289 ( .A(y[893]), .B(x[893]), .Z(n151) );
  NAND U290 ( .A(n152), .B(n151), .Z(n6108) );
  NANDN U291 ( .A(x[891]), .B(y[891]), .Z(n154) );
  NANDN U292 ( .A(x[892]), .B(y[892]), .Z(n153) );
  AND U293 ( .A(n154), .B(n153), .Z(n6105) );
  NANDN U294 ( .A(x[886]), .B(y[886]), .Z(n155) );
  NANDN U295 ( .A(x[887]), .B(y[887]), .Z(n2918) );
  AND U296 ( .A(n155), .B(n2918), .Z(n6093) );
  NANDN U297 ( .A(y[885]), .B(x[885]), .Z(n156) );
  NANDN U298 ( .A(y[886]), .B(x[886]), .Z(n2916) );
  NAND U299 ( .A(n156), .B(n2916), .Z(n6092) );
  NANDN U300 ( .A(x[884]), .B(y[884]), .Z(n4150) );
  IV U301 ( .A(y[885]), .Z(n4153) );
  OR U302 ( .A(x[885]), .B(n4153), .Z(n157) );
  NAND U303 ( .A(n4150), .B(n157), .Z(n6090) );
  ANDN U304 ( .B(y[883]), .A(x[883]), .Z(n6085) );
  NANDN U305 ( .A(x[882]), .B(y[882]), .Z(n6080) );
  NANDN U306 ( .A(n6085), .B(n6080), .Z(n158) );
  NANDN U307 ( .A(y[883]), .B(x[883]), .Z(n2617) );
  AND U308 ( .A(n158), .B(n2617), .Z(n4149) );
  NANDN U309 ( .A(x[881]), .B(y[881]), .Z(n6081) );
  NANDN U310 ( .A(x[876]), .B(y[876]), .Z(n6068) );
  ANDN U311 ( .B(x[875]), .A(y[875]), .Z(n163) );
  IV U312 ( .A(y[875]), .Z(n4135) );
  IV U313 ( .A(x[875]), .Z(n4132) );
  NANDN U314 ( .A(n4135), .B(n4132), .Z(n160) );
  NANDN U315 ( .A(x[874]), .B(y[874]), .Z(n159) );
  NAND U316 ( .A(n160), .B(n159), .Z(n165) );
  ANDN U317 ( .B(x[874]), .A(y[874]), .Z(n4133) );
  NANDN U318 ( .A(y[873]), .B(x[873]), .Z(n2919) );
  NANDN U319 ( .A(n4133), .B(n2919), .Z(n161) );
  NANDN U320 ( .A(n165), .B(n161), .Z(n162) );
  NANDN U321 ( .A(n163), .B(n162), .Z(n6066) );
  NANDN U322 ( .A(x[873]), .B(y[873]), .Z(n164) );
  NANDN U323 ( .A(n165), .B(n164), .Z(n6064) );
  NANDN U324 ( .A(x[872]), .B(y[872]), .Z(n6059) );
  ANDN U325 ( .B(y[870]), .A(x[870]), .Z(n6051) );
  NANDN U326 ( .A(x[871]), .B(y[871]), .Z(n6057) );
  NANDN U327 ( .A(n6051), .B(n6057), .Z(n166) );
  NANDN U328 ( .A(y[871]), .B(x[871]), .Z(n167) );
  AND U329 ( .A(n166), .B(n167), .Z(n4128) );
  NANDN U330 ( .A(y[869]), .B(x[869]), .Z(n169) );
  NANDN U331 ( .A(y[868]), .B(x[868]), .Z(n168) );
  NAND U332 ( .A(n169), .B(n168), .Z(n6050) );
  NANDN U333 ( .A(y[867]), .B(x[867]), .Z(n171) );
  NANDN U334 ( .A(y[866]), .B(x[866]), .Z(n170) );
  NAND U335 ( .A(n171), .B(n170), .Z(n6046) );
  IV U336 ( .A(y[862]), .Z(n2920) );
  NANDN U337 ( .A(x[863]), .B(y[863]), .Z(n4117) );
  NAND U338 ( .A(n4114), .B(n4117), .Z(n6036) );
  NANDN U339 ( .A(y[861]), .B(x[861]), .Z(n4108) );
  NANDN U340 ( .A(y[862]), .B(x[862]), .Z(n172) );
  NAND U341 ( .A(n4108), .B(n172), .Z(n6034) );
  NANDN U342 ( .A(y[860]), .B(x[860]), .Z(n6029) );
  NANDN U343 ( .A(y[859]), .B(x[859]), .Z(n2572) );
  NANDN U344 ( .A(y[858]), .B(x[858]), .Z(n173) );
  NAND U345 ( .A(n2572), .B(n173), .Z(n6026) );
  NANDN U346 ( .A(y[854]), .B(x[854]), .Z(n175) );
  NANDN U347 ( .A(y[855]), .B(x[855]), .Z(n174) );
  AND U348 ( .A(n175), .B(n174), .Z(n6015) );
  NANDN U349 ( .A(y[844]), .B(x[844]), .Z(n177) );
  NANDN U350 ( .A(y[845]), .B(x[845]), .Z(n176) );
  AND U351 ( .A(n177), .B(n176), .Z(n5991) );
  NANDN U352 ( .A(y[838]), .B(x[838]), .Z(n179) );
  NANDN U353 ( .A(y[839]), .B(x[839]), .Z(n178) );
  AND U354 ( .A(n179), .B(n178), .Z(n5979) );
  NANDN U355 ( .A(y[832]), .B(x[832]), .Z(n181) );
  NANDN U356 ( .A(y[833]), .B(x[833]), .Z(n180) );
  AND U357 ( .A(n181), .B(n180), .Z(n5967) );
  NANDN U358 ( .A(y[826]), .B(x[826]), .Z(n183) );
  NANDN U359 ( .A(y[827]), .B(x[827]), .Z(n182) );
  AND U360 ( .A(n183), .B(n182), .Z(n5955) );
  NANDN U361 ( .A(y[820]), .B(x[820]), .Z(n185) );
  NANDN U362 ( .A(y[821]), .B(x[821]), .Z(n184) );
  AND U363 ( .A(n185), .B(n184), .Z(n5943) );
  NANDN U364 ( .A(y[814]), .B(x[814]), .Z(n187) );
  NANDN U365 ( .A(y[815]), .B(x[815]), .Z(n186) );
  AND U366 ( .A(n187), .B(n186), .Z(n5931) );
  NANDN U367 ( .A(x[809]), .B(y[809]), .Z(n2443) );
  NANDN U368 ( .A(y[809]), .B(x[809]), .Z(n4047) );
  NANDN U369 ( .A(y[808]), .B(x[808]), .Z(n188) );
  AND U370 ( .A(n4047), .B(n188), .Z(n189) );
  ANDN U371 ( .B(n2443), .A(n189), .Z(n5920) );
  NANDN U372 ( .A(y[807]), .B(x[807]), .Z(n5915) );
  NANDN U373 ( .A(y[806]), .B(x[806]), .Z(n190) );
  NAND U374 ( .A(n5915), .B(n190), .Z(n5912) );
  NANDN U375 ( .A(x[807]), .B(y[807]), .Z(n2440) );
  AND U376 ( .A(n5912), .B(n2440), .Z(n4043) );
  NANDN U377 ( .A(x[798]), .B(y[798]), .Z(n192) );
  NANDN U378 ( .A(x[797]), .B(y[797]), .Z(n191) );
  NAND U379 ( .A(n192), .B(n191), .Z(n5894) );
  NANDN U380 ( .A(x[796]), .B(y[796]), .Z(n194) );
  NANDN U381 ( .A(x[795]), .B(y[795]), .Z(n193) );
  NAND U382 ( .A(n194), .B(n193), .Z(n5890) );
  NANDN U383 ( .A(x[792]), .B(y[792]), .Z(n196) );
  NANDN U384 ( .A(x[791]), .B(y[791]), .Z(n195) );
  NAND U385 ( .A(n196), .B(n195), .Z(n5882) );
  NANDN U386 ( .A(x[790]), .B(y[790]), .Z(n198) );
  NANDN U387 ( .A(x[789]), .B(y[789]), .Z(n197) );
  NAND U388 ( .A(n198), .B(n197), .Z(n5878) );
  NANDN U389 ( .A(x[786]), .B(y[786]), .Z(n200) );
  NANDN U390 ( .A(x[785]), .B(y[785]), .Z(n199) );
  NAND U391 ( .A(n200), .B(n199), .Z(n5870) );
  ANDN U392 ( .B(x[782]), .A(y[782]), .Z(n5857) );
  NANDN U393 ( .A(y[783]), .B(x[783]), .Z(n5863) );
  NANDN U394 ( .A(n5857), .B(n5863), .Z(n201) );
  NANDN U395 ( .A(x[783]), .B(y[783]), .Z(n202) );
  AND U396 ( .A(n201), .B(n202), .Z(n4011) );
  NANDN U397 ( .A(x[780]), .B(y[780]), .Z(n204) );
  NANDN U398 ( .A(x[779]), .B(y[779]), .Z(n203) );
  AND U399 ( .A(n204), .B(n203), .Z(n206) );
  NANDN U400 ( .A(x[781]), .B(y[781]), .Z(n205) );
  NAND U401 ( .A(n206), .B(n205), .Z(n5856) );
  NANDN U402 ( .A(x[778]), .B(y[778]), .Z(n208) );
  NANDN U403 ( .A(x[777]), .B(y[777]), .Z(n207) );
  NAND U404 ( .A(n208), .B(n207), .Z(n5852) );
  NANDN U405 ( .A(x[773]), .B(y[773]), .Z(n2369) );
  NANDN U406 ( .A(y[772]), .B(x[772]), .Z(n209) );
  ANDN U407 ( .B(x[773]), .A(y[773]), .Z(n5842) );
  ANDN U408 ( .B(n209), .A(n5842), .Z(n210) );
  ANDN U409 ( .B(n2369), .A(n210), .Z(n4000) );
  NANDN U410 ( .A(x[768]), .B(y[768]), .Z(n212) );
  NANDN U411 ( .A(x[767]), .B(y[767]), .Z(n211) );
  NAND U412 ( .A(n212), .B(n211), .Z(n5829) );
  NANDN U413 ( .A(x[766]), .B(y[766]), .Z(n214) );
  NANDN U414 ( .A(x[765]), .B(y[765]), .Z(n213) );
  NAND U415 ( .A(n214), .B(n213), .Z(n5826) );
  NANDN U416 ( .A(x[762]), .B(y[762]), .Z(n216) );
  NANDN U417 ( .A(x[761]), .B(y[761]), .Z(n215) );
  NAND U418 ( .A(n216), .B(n215), .Z(n5817) );
  NANDN U419 ( .A(x[759]), .B(y[759]), .Z(n2338) );
  NANDN U420 ( .A(y[758]), .B(x[758]), .Z(n217) );
  ANDN U421 ( .B(x[759]), .A(y[759]), .Z(n5812) );
  ANDN U422 ( .B(n217), .A(n5812), .Z(n218) );
  ANDN U423 ( .B(n2338), .A(n218), .Z(n3985) );
  NANDN U424 ( .A(x[755]), .B(y[755]), .Z(n221) );
  NANDN U425 ( .A(y[754]), .B(x[754]), .Z(n219) );
  ANDN U426 ( .B(x[755]), .A(y[755]), .Z(n5800) );
  ANDN U427 ( .B(n219), .A(n5800), .Z(n220) );
  ANDN U428 ( .B(n221), .A(n220), .Z(n3979) );
  ANDN U429 ( .B(y[753]), .A(x[753]), .Z(n5793) );
  OR U430 ( .A(n5798), .B(n5793), .Z(n3977) );
  NANDN U431 ( .A(x[750]), .B(y[750]), .Z(n223) );
  NANDN U432 ( .A(x[749]), .B(y[749]), .Z(n222) );
  NAND U433 ( .A(n223), .B(n222), .Z(n5786) );
  ANDN U434 ( .B(x[747]), .A(y[747]), .Z(n5780) );
  NANDN U435 ( .A(y[746]), .B(x[746]), .Z(n224) );
  NANDN U436 ( .A(n5780), .B(n224), .Z(n5776) );
  NANDN U437 ( .A(x[747]), .B(y[747]), .Z(n2315) );
  AND U438 ( .A(n5776), .B(n2315), .Z(n3969) );
  NANDN U439 ( .A(x[744]), .B(y[744]), .Z(n226) );
  NANDN U440 ( .A(x[743]), .B(y[743]), .Z(n225) );
  NAND U441 ( .A(n226), .B(n225), .Z(n5769) );
  NANDN U442 ( .A(x[742]), .B(y[742]), .Z(n228) );
  NANDN U443 ( .A(x[741]), .B(y[741]), .Z(n227) );
  NAND U444 ( .A(n228), .B(n227), .Z(n5766) );
  NANDN U445 ( .A(x[738]), .B(y[738]), .Z(n230) );
  NANDN U446 ( .A(x[737]), .B(y[737]), .Z(n229) );
  NAND U447 ( .A(n230), .B(n229), .Z(n5757) );
  NANDN U448 ( .A(x[736]), .B(y[736]), .Z(n232) );
  NANDN U449 ( .A(x[735]), .B(y[735]), .Z(n231) );
  NAND U450 ( .A(n232), .B(n231), .Z(n5754) );
  NANDN U451 ( .A(x[731]), .B(y[731]), .Z(n234) );
  NANDN U452 ( .A(x[730]), .B(y[730]), .Z(n233) );
  AND U453 ( .A(n234), .B(n233), .Z(n240) );
  NANDN U454 ( .A(x[728]), .B(y[728]), .Z(n235) );
  NANDN U455 ( .A(y[729]), .B(n235), .Z(n238) );
  XNOR U456 ( .A(n235), .B(y[729]), .Z(n236) );
  NAND U457 ( .A(n236), .B(x[729]), .Z(n237) );
  NAND U458 ( .A(n238), .B(n237), .Z(n239) );
  NAND U459 ( .A(n240), .B(n239), .Z(n5742) );
  NANDN U460 ( .A(y[729]), .B(x[729]), .Z(n242) );
  NANDN U461 ( .A(y[728]), .B(x[728]), .Z(n241) );
  AND U462 ( .A(n242), .B(n241), .Z(n248) );
  NANDN U463 ( .A(y[726]), .B(x[726]), .Z(n243) );
  NANDN U464 ( .A(x[727]), .B(n243), .Z(n246) );
  XNOR U465 ( .A(n243), .B(x[727]), .Z(n244) );
  NAND U466 ( .A(n244), .B(y[727]), .Z(n245) );
  NAND U467 ( .A(n246), .B(n245), .Z(n247) );
  NAND U468 ( .A(n248), .B(n247), .Z(n5740) );
  NANDN U469 ( .A(x[724]), .B(y[724]), .Z(n250) );
  NANDN U470 ( .A(x[723]), .B(y[723]), .Z(n249) );
  NAND U471 ( .A(n250), .B(n249), .Z(n5733) );
  NANDN U472 ( .A(x[721]), .B(y[721]), .Z(n2264) );
  NANDN U473 ( .A(y[720]), .B(x[720]), .Z(n5724) );
  ANDN U474 ( .B(x[721]), .A(y[721]), .Z(n5727) );
  ANDN U475 ( .B(n5724), .A(n5727), .Z(n251) );
  ANDN U476 ( .B(n2264), .A(n251), .Z(n3943) );
  NANDN U477 ( .A(x[718]), .B(y[718]), .Z(n253) );
  NANDN U478 ( .A(x[717]), .B(y[717]), .Z(n252) );
  NAND U479 ( .A(n253), .B(n252), .Z(n5718) );
  NANDN U480 ( .A(x[716]), .B(y[716]), .Z(n255) );
  NANDN U481 ( .A(x[715]), .B(y[715]), .Z(n254) );
  NAND U482 ( .A(n255), .B(n254), .Z(n5714) );
  NANDN U483 ( .A(x[712]), .B(y[712]), .Z(n261) );
  ANDN U484 ( .B(y[710]), .A(x[710]), .Z(n256) );
  OR U485 ( .A(n256), .B(y[711]), .Z(n259) );
  XOR U486 ( .A(y[711]), .B(n256), .Z(n257) );
  NAND U487 ( .A(n257), .B(x[711]), .Z(n258) );
  NAND U488 ( .A(n259), .B(n258), .Z(n260) );
  NAND U489 ( .A(n261), .B(n260), .Z(n5706) );
  NANDN U490 ( .A(y[702]), .B(x[702]), .Z(n263) );
  NANDN U491 ( .A(y[703]), .B(x[703]), .Z(n262) );
  AND U492 ( .A(n263), .B(n262), .Z(n5691) );
  NANDN U493 ( .A(y[690]), .B(x[690]), .Z(n265) );
  NANDN U494 ( .A(y[691]), .B(x[691]), .Z(n264) );
  AND U495 ( .A(n265), .B(n264), .Z(n5667) );
  NANDN U496 ( .A(y[684]), .B(x[684]), .Z(n267) );
  NANDN U497 ( .A(y[685]), .B(x[685]), .Z(n266) );
  AND U498 ( .A(n267), .B(n266), .Z(n5655) );
  NANDN U499 ( .A(y[678]), .B(x[678]), .Z(n269) );
  NANDN U500 ( .A(y[679]), .B(x[679]), .Z(n268) );
  AND U501 ( .A(n269), .B(n268), .Z(n5643) );
  NANDN U502 ( .A(x[677]), .B(y[677]), .Z(n2151) );
  NANDN U503 ( .A(y[676]), .B(x[676]), .Z(n270) );
  ANDN U504 ( .B(x[677]), .A(y[677]), .Z(n3892) );
  ANDN U505 ( .B(n270), .A(n3892), .Z(n3888) );
  ANDN U506 ( .B(n2151), .A(n3888), .Z(n5640) );
  NANDN U507 ( .A(y[672]), .B(x[672]), .Z(n272) );
  NANDN U508 ( .A(y[673]), .B(x[673]), .Z(n271) );
  AND U509 ( .A(n272), .B(n271), .Z(n5631) );
  NANDN U510 ( .A(y[666]), .B(x[666]), .Z(n274) );
  NANDN U511 ( .A(y[667]), .B(x[667]), .Z(n273) );
  AND U512 ( .A(n274), .B(n273), .Z(n5619) );
  NANDN U513 ( .A(y[660]), .B(x[660]), .Z(n276) );
  NANDN U514 ( .A(y[661]), .B(x[661]), .Z(n275) );
  AND U515 ( .A(n276), .B(n275), .Z(n5607) );
  NANDN U516 ( .A(y[654]), .B(x[654]), .Z(n278) );
  NANDN U517 ( .A(y[655]), .B(x[655]), .Z(n277) );
  AND U518 ( .A(n278), .B(n277), .Z(n5595) );
  NANDN U519 ( .A(y[648]), .B(x[648]), .Z(n280) );
  NANDN U520 ( .A(y[649]), .B(x[649]), .Z(n279) );
  AND U521 ( .A(n280), .B(n279), .Z(n5583) );
  NANDN U522 ( .A(y[642]), .B(x[642]), .Z(n282) );
  NANDN U523 ( .A(y[643]), .B(x[643]), .Z(n281) );
  AND U524 ( .A(n282), .B(n281), .Z(n5571) );
  NANDN U525 ( .A(y[636]), .B(x[636]), .Z(n284) );
  NANDN U526 ( .A(y[637]), .B(x[637]), .Z(n283) );
  AND U527 ( .A(n284), .B(n283), .Z(n5559) );
  NANDN U528 ( .A(y[630]), .B(x[630]), .Z(n286) );
  NANDN U529 ( .A(y[631]), .B(x[631]), .Z(n285) );
  AND U530 ( .A(n286), .B(n285), .Z(n5547) );
  ANDN U531 ( .B(x[629]), .A(y[629]), .Z(n4364) );
  NANDN U532 ( .A(y[628]), .B(x[628]), .Z(n4365) );
  NANDN U533 ( .A(n4364), .B(n4365), .Z(n3836) );
  NANDN U534 ( .A(x[622]), .B(y[622]), .Z(n288) );
  NANDN U535 ( .A(x[621]), .B(y[621]), .Z(n287) );
  NAND U536 ( .A(n288), .B(n287), .Z(n5527) );
  NANDN U537 ( .A(y[616]), .B(x[616]), .Z(n289) );
  ANDN U538 ( .B(x[617]), .A(y[617]), .Z(n2934) );
  ANDN U539 ( .B(n289), .A(n2934), .Z(n3819) );
  ANDN U540 ( .B(y[617]), .A(x[617]), .Z(n291) );
  NOR U541 ( .A(n3819), .B(n291), .Z(n5518) );
  NANDN U542 ( .A(x[616]), .B(y[616]), .Z(n290) );
  NANDN U543 ( .A(n291), .B(n290), .Z(n2933) );
  NANDN U544 ( .A(x[615]), .B(y[615]), .Z(n3817) );
  NANDN U545 ( .A(n2933), .B(n3817), .Z(n5515) );
  NANDN U546 ( .A(x[612]), .B(y[612]), .Z(n2936) );
  NANDN U547 ( .A(x[610]), .B(y[610]), .Z(n293) );
  NANDN U548 ( .A(x[609]), .B(y[609]), .Z(n292) );
  NAND U549 ( .A(n293), .B(n292), .Z(n5503) );
  NANDN U550 ( .A(x[608]), .B(y[608]), .Z(n295) );
  NANDN U551 ( .A(x[607]), .B(y[607]), .Z(n294) );
  NAND U552 ( .A(n295), .B(n294), .Z(n2942) );
  NANDN U553 ( .A(x[606]), .B(y[606]), .Z(n2940) );
  NANDN U554 ( .A(x[605]), .B(y[605]), .Z(n2945) );
  AND U555 ( .A(n2940), .B(n2945), .Z(n1981) );
  NANDN U556 ( .A(y[605]), .B(x[605]), .Z(n2944) );
  NANDN U557 ( .A(y[604]), .B(x[604]), .Z(n296) );
  NAND U558 ( .A(n2944), .B(n296), .Z(n5494) );
  NANDN U559 ( .A(x[603]), .B(y[603]), .Z(n5492) );
  ANDN U560 ( .B(y[604]), .A(x[604]), .Z(n2943) );
  ANDN U561 ( .B(n5492), .A(n2943), .Z(n1978) );
  NANDN U562 ( .A(x[600]), .B(y[600]), .Z(n298) );
  NANDN U563 ( .A(x[599]), .B(y[599]), .Z(n297) );
  NAND U564 ( .A(n298), .B(n297), .Z(n5484) );
  NANDN U565 ( .A(x[598]), .B(y[598]), .Z(n300) );
  NANDN U566 ( .A(x[597]), .B(y[597]), .Z(n299) );
  NAND U567 ( .A(n300), .B(n299), .Z(n5479) );
  NANDN U568 ( .A(x[594]), .B(y[594]), .Z(n302) );
  NANDN U569 ( .A(x[593]), .B(y[593]), .Z(n301) );
  NAND U570 ( .A(n302), .B(n301), .Z(n5472) );
  NANDN U571 ( .A(x[592]), .B(y[592]), .Z(n304) );
  NANDN U572 ( .A(x[591]), .B(y[591]), .Z(n303) );
  NAND U573 ( .A(n304), .B(n303), .Z(n5468) );
  NANDN U574 ( .A(x[590]), .B(y[590]), .Z(n5463) );
  NANDN U575 ( .A(x[589]), .B(y[589]), .Z(n306) );
  NANDN U576 ( .A(y[588]), .B(x[588]), .Z(n5457) );
  ANDN U577 ( .B(x[589]), .A(y[589]), .Z(n5461) );
  ANDN U578 ( .B(n5457), .A(n5461), .Z(n305) );
  ANDN U579 ( .B(n306), .A(n305), .Z(n3790) );
  ANDN U580 ( .B(y[587]), .A(x[587]), .Z(n5456) );
  OR U581 ( .A(n5460), .B(n5456), .Z(n3788) );
  NANDN U582 ( .A(x[586]), .B(y[586]), .Z(n308) );
  NANDN U583 ( .A(x[585]), .B(y[585]), .Z(n307) );
  NAND U584 ( .A(n308), .B(n307), .Z(n5452) );
  NANDN U585 ( .A(y[583]), .B(x[583]), .Z(n2948) );
  IV U586 ( .A(x[582]), .Z(n2950) );
  IV U587 ( .A(y[582]), .Z(n2949) );
  NANDN U588 ( .A(n2950), .B(n2949), .Z(n309) );
  NAND U589 ( .A(n2948), .B(n309), .Z(n5445) );
  NANDN U590 ( .A(x[580]), .B(y[580]), .Z(n311) );
  NANDN U591 ( .A(x[579]), .B(y[579]), .Z(n310) );
  NAND U592 ( .A(n311), .B(n310), .Z(n5440) );
  NANDN U593 ( .A(x[576]), .B(y[576]), .Z(n313) );
  NANDN U594 ( .A(x[575]), .B(y[575]), .Z(n312) );
  NAND U595 ( .A(n313), .B(n312), .Z(n5432) );
  NANDN U596 ( .A(x[574]), .B(y[574]), .Z(n315) );
  NANDN U597 ( .A(x[573]), .B(y[573]), .Z(n314) );
  NAND U598 ( .A(n315), .B(n314), .Z(n5428) );
  NANDN U599 ( .A(x[569]), .B(y[569]), .Z(n317) );
  NANDN U600 ( .A(x[568]), .B(y[568]), .Z(n316) );
  AND U601 ( .A(n317), .B(n316), .Z(n323) );
  NANDN U602 ( .A(x[566]), .B(y[566]), .Z(n318) );
  NANDN U603 ( .A(y[567]), .B(n318), .Z(n321) );
  XNOR U604 ( .A(n318), .B(y[567]), .Z(n319) );
  NAND U605 ( .A(n319), .B(x[567]), .Z(n320) );
  NAND U606 ( .A(n321), .B(n320), .Z(n322) );
  NAND U607 ( .A(n323), .B(n322), .Z(n5416) );
  NANDN U608 ( .A(x[562]), .B(y[562]), .Z(n325) );
  NANDN U609 ( .A(x[561]), .B(y[561]), .Z(n324) );
  NAND U610 ( .A(n325), .B(n324), .Z(n5408) );
  NANDN U611 ( .A(x[560]), .B(y[560]), .Z(n327) );
  NANDN U612 ( .A(x[559]), .B(y[559]), .Z(n326) );
  NAND U613 ( .A(n327), .B(n326), .Z(n5404) );
  NANDN U614 ( .A(x[558]), .B(y[558]), .Z(n5399) );
  NANDN U615 ( .A(x[557]), .B(y[557]), .Z(n329) );
  NANDN U616 ( .A(y[556]), .B(x[556]), .Z(n5393) );
  ANDN U617 ( .B(x[557]), .A(y[557]), .Z(n5397) );
  ANDN U618 ( .B(n5393), .A(n5397), .Z(n328) );
  ANDN U619 ( .B(n329), .A(n328), .Z(n3754) );
  ANDN U620 ( .B(y[555]), .A(x[555]), .Z(n5392) );
  OR U621 ( .A(n5396), .B(n5392), .Z(n3752) );
  NANDN U622 ( .A(x[554]), .B(y[554]), .Z(n331) );
  NANDN U623 ( .A(x[553]), .B(y[553]), .Z(n330) );
  NAND U624 ( .A(n331), .B(n330), .Z(n5388) );
  NANDN U625 ( .A(x[550]), .B(y[550]), .Z(n333) );
  NANDN U626 ( .A(x[549]), .B(y[549]), .Z(n332) );
  NAND U627 ( .A(n333), .B(n332), .Z(n5380) );
  NANDN U628 ( .A(x[548]), .B(y[548]), .Z(n335) );
  NANDN U629 ( .A(x[547]), .B(y[547]), .Z(n334) );
  NAND U630 ( .A(n335), .B(n334), .Z(n5376) );
  NANDN U631 ( .A(x[544]), .B(y[544]), .Z(n337) );
  NANDN U632 ( .A(x[543]), .B(y[543]), .Z(n336) );
  NAND U633 ( .A(n337), .B(n336), .Z(n5368) );
  NANDN U634 ( .A(x[542]), .B(y[542]), .Z(n339) );
  NANDN U635 ( .A(x[541]), .B(y[541]), .Z(n338) );
  NAND U636 ( .A(n339), .B(n338), .Z(n5364) );
  NANDN U637 ( .A(x[538]), .B(y[538]), .Z(n341) );
  NANDN U638 ( .A(x[537]), .B(y[537]), .Z(n340) );
  NAND U639 ( .A(n341), .B(n340), .Z(n5356) );
  NANDN U640 ( .A(x[536]), .B(y[536]), .Z(n343) );
  NANDN U641 ( .A(x[535]), .B(y[535]), .Z(n342) );
  NAND U642 ( .A(n343), .B(n342), .Z(n5352) );
  NANDN U643 ( .A(x[534]), .B(y[534]), .Z(n5347) );
  NANDN U644 ( .A(x[533]), .B(y[533]), .Z(n345) );
  NANDN U645 ( .A(y[532]), .B(x[532]), .Z(n5341) );
  ANDN U646 ( .B(x[533]), .A(y[533]), .Z(n5345) );
  ANDN U647 ( .B(n5341), .A(n5345), .Z(n344) );
  ANDN U648 ( .B(n345), .A(n344), .Z(n3728) );
  ANDN U649 ( .B(y[531]), .A(x[531]), .Z(n5340) );
  OR U650 ( .A(n5344), .B(n5340), .Z(n3726) );
  NANDN U651 ( .A(x[530]), .B(y[530]), .Z(n347) );
  NANDN U652 ( .A(x[529]), .B(y[529]), .Z(n346) );
  NAND U653 ( .A(n347), .B(n346), .Z(n5336) );
  NANDN U654 ( .A(x[526]), .B(y[526]), .Z(n349) );
  NANDN U655 ( .A(x[525]), .B(y[525]), .Z(n348) );
  NAND U656 ( .A(n349), .B(n348), .Z(n5328) );
  NANDN U657 ( .A(x[524]), .B(y[524]), .Z(n351) );
  NANDN U658 ( .A(x[523]), .B(y[523]), .Z(n350) );
  NAND U659 ( .A(n351), .B(n350), .Z(n5324) );
  NANDN U660 ( .A(x[520]), .B(y[520]), .Z(n353) );
  NANDN U661 ( .A(x[519]), .B(y[519]), .Z(n352) );
  NAND U662 ( .A(n353), .B(n352), .Z(n5316) );
  NANDN U663 ( .A(x[518]), .B(y[518]), .Z(n355) );
  NANDN U664 ( .A(x[517]), .B(y[517]), .Z(n354) );
  NAND U665 ( .A(n355), .B(n354), .Z(n5312) );
  NANDN U666 ( .A(x[514]), .B(y[514]), .Z(n357) );
  NANDN U667 ( .A(x[513]), .B(y[513]), .Z(n356) );
  NAND U668 ( .A(n357), .B(n356), .Z(n5304) );
  NANDN U669 ( .A(x[512]), .B(y[512]), .Z(n359) );
  NANDN U670 ( .A(x[511]), .B(y[511]), .Z(n358) );
  NAND U671 ( .A(n359), .B(n358), .Z(n5300) );
  NANDN U672 ( .A(x[508]), .B(y[508]), .Z(n361) );
  NANDN U673 ( .A(x[507]), .B(y[507]), .Z(n360) );
  NAND U674 ( .A(n361), .B(n360), .Z(n5292) );
  ANDN U675 ( .B(y[503]), .A(x[503]), .Z(n3692) );
  NANDN U676 ( .A(x[505]), .B(y[505]), .Z(n1758) );
  NANDN U677 ( .A(x[504]), .B(y[504]), .Z(n362) );
  NAND U678 ( .A(n1758), .B(n362), .Z(n3696) );
  NOR U679 ( .A(n3692), .B(n3696), .Z(n5283) );
  NANDN U680 ( .A(x[502]), .B(y[502]), .Z(n364) );
  NANDN U681 ( .A(x[501]), .B(y[501]), .Z(n363) );
  NAND U682 ( .A(n364), .B(n363), .Z(n5280) );
  NANDN U683 ( .A(x[500]), .B(y[500]), .Z(n366) );
  NANDN U684 ( .A(x[499]), .B(y[499]), .Z(n365) );
  NAND U685 ( .A(n366), .B(n365), .Z(n5276) );
  NANDN U686 ( .A(x[496]), .B(y[496]), .Z(n368) );
  NANDN U687 ( .A(x[495]), .B(y[495]), .Z(n367) );
  NAND U688 ( .A(n368), .B(n367), .Z(n5268) );
  NANDN U689 ( .A(x[494]), .B(y[494]), .Z(n370) );
  NANDN U690 ( .A(x[493]), .B(y[493]), .Z(n369) );
  NAND U691 ( .A(n370), .B(n369), .Z(n5264) );
  NANDN U692 ( .A(x[490]), .B(y[490]), .Z(n372) );
  NANDN U693 ( .A(x[489]), .B(y[489]), .Z(n371) );
  NAND U694 ( .A(n372), .B(n371), .Z(n5256) );
  NANDN U695 ( .A(x[488]), .B(y[488]), .Z(n374) );
  NANDN U696 ( .A(x[487]), .B(y[487]), .Z(n373) );
  NAND U697 ( .A(n374), .B(n373), .Z(n5252) );
  NANDN U698 ( .A(x[484]), .B(y[484]), .Z(n376) );
  NANDN U699 ( .A(x[483]), .B(y[483]), .Z(n375) );
  NAND U700 ( .A(n376), .B(n375), .Z(n5244) );
  NANDN U701 ( .A(x[482]), .B(y[482]), .Z(n378) );
  NANDN U702 ( .A(x[481]), .B(y[481]), .Z(n377) );
  NAND U703 ( .A(n378), .B(n377), .Z(n5240) );
  NANDN U704 ( .A(x[478]), .B(y[478]), .Z(n380) );
  NANDN U705 ( .A(x[477]), .B(y[477]), .Z(n379) );
  NAND U706 ( .A(n380), .B(n379), .Z(n5232) );
  NANDN U707 ( .A(x[476]), .B(y[476]), .Z(n382) );
  NANDN U708 ( .A(x[475]), .B(y[475]), .Z(n381) );
  NAND U709 ( .A(n382), .B(n381), .Z(n5228) );
  NANDN U710 ( .A(x[472]), .B(y[472]), .Z(n384) );
  NANDN U711 ( .A(x[471]), .B(y[471]), .Z(n383) );
  NAND U712 ( .A(n384), .B(n383), .Z(n5220) );
  NANDN U713 ( .A(x[470]), .B(y[470]), .Z(n386) );
  NANDN U714 ( .A(x[469]), .B(y[469]), .Z(n385) );
  NAND U715 ( .A(n386), .B(n385), .Z(n5216) );
  NANDN U716 ( .A(x[466]), .B(y[466]), .Z(n388) );
  NANDN U717 ( .A(x[465]), .B(y[465]), .Z(n387) );
  NAND U718 ( .A(n388), .B(n387), .Z(n5208) );
  NANDN U719 ( .A(x[463]), .B(y[463]), .Z(n1661) );
  NANDN U720 ( .A(y[462]), .B(x[462]), .Z(n5197) );
  ANDN U721 ( .B(x[463]), .A(y[463]), .Z(n5201) );
  ANDN U722 ( .B(n5197), .A(n5201), .Z(n389) );
  ANDN U723 ( .B(n1661), .A(n389), .Z(n3650) );
  NANDN U724 ( .A(y[461]), .B(x[461]), .Z(n1660) );
  NANDN U725 ( .A(y[460]), .B(x[460]), .Z(n390) );
  NAND U726 ( .A(n1660), .B(n390), .Z(n3646) );
  NANDN U727 ( .A(y[459]), .B(x[459]), .Z(n3643) );
  NANDN U728 ( .A(y[458]), .B(x[458]), .Z(n391) );
  AND U729 ( .A(n3643), .B(n391), .Z(n392) );
  NANDN U730 ( .A(x[459]), .B(y[459]), .Z(n395) );
  NANDN U731 ( .A(n392), .B(n395), .Z(n393) );
  NANDN U732 ( .A(n3646), .B(n393), .Z(n5194) );
  NANDN U733 ( .A(x[458]), .B(y[458]), .Z(n394) );
  NAND U734 ( .A(n395), .B(n394), .Z(n5192) );
  ANDN U735 ( .B(x[457]), .A(y[457]), .Z(n3639) );
  NANDN U736 ( .A(y[456]), .B(x[456]), .Z(n3635) );
  NANDN U737 ( .A(n3639), .B(n3635), .Z(n396) );
  ANDN U738 ( .B(y[457]), .A(x[457]), .Z(n398) );
  ANDN U739 ( .B(n396), .A(n398), .Z(n5190) );
  NANDN U740 ( .A(x[456]), .B(y[456]), .Z(n397) );
  NANDN U741 ( .A(n398), .B(n397), .Z(n5187) );
  NANDN U742 ( .A(x[452]), .B(y[452]), .Z(n400) );
  NANDN U743 ( .A(x[451]), .B(y[451]), .Z(n399) );
  NAND U744 ( .A(n400), .B(n399), .Z(n5180) );
  NANDN U745 ( .A(x[449]), .B(y[449]), .Z(n1636) );
  NANDN U746 ( .A(y[448]), .B(x[448]), .Z(n3624) );
  ANDN U747 ( .B(x[449]), .A(y[449]), .Z(n3627) );
  ANDN U748 ( .B(n3624), .A(n3627), .Z(n401) );
  ANDN U749 ( .B(n1636), .A(n401), .Z(n5174) );
  NANDN U750 ( .A(x[441]), .B(y[441]), .Z(n403) );
  NANDN U751 ( .A(x[442]), .B(y[442]), .Z(n402) );
  AND U752 ( .A(n403), .B(n402), .Z(n5159) );
  NANDN U753 ( .A(x[435]), .B(y[435]), .Z(n405) );
  NANDN U754 ( .A(x[436]), .B(y[436]), .Z(n404) );
  AND U755 ( .A(n405), .B(n404), .Z(n5147) );
  NANDN U756 ( .A(x[429]), .B(y[429]), .Z(n407) );
  NANDN U757 ( .A(x[430]), .B(y[430]), .Z(n406) );
  AND U758 ( .A(n407), .B(n406), .Z(n5135) );
  NANDN U759 ( .A(x[423]), .B(y[423]), .Z(n409) );
  NANDN U760 ( .A(x[424]), .B(y[424]), .Z(n408) );
  AND U761 ( .A(n409), .B(n408), .Z(n5123) );
  NANDN U762 ( .A(x[417]), .B(y[417]), .Z(n411) );
  NANDN U763 ( .A(x[418]), .B(y[418]), .Z(n410) );
  AND U764 ( .A(n411), .B(n410), .Z(n5111) );
  NANDN U765 ( .A(x[411]), .B(y[411]), .Z(n413) );
  NANDN U766 ( .A(x[412]), .B(y[412]), .Z(n412) );
  AND U767 ( .A(n413), .B(n412), .Z(n5099) );
  NANDN U768 ( .A(x[407]), .B(y[407]), .Z(n1527) );
  NANDN U769 ( .A(y[406]), .B(x[406]), .Z(n3576) );
  ANDN U770 ( .B(x[407]), .A(y[407]), .Z(n3579) );
  ANDN U771 ( .B(n3576), .A(n3579), .Z(n414) );
  ANDN U772 ( .B(n1527), .A(n414), .Z(n5090) );
  NANDN U773 ( .A(x[399]), .B(y[399]), .Z(n416) );
  NANDN U774 ( .A(x[400]), .B(y[400]), .Z(n415) );
  AND U775 ( .A(n416), .B(n415), .Z(n5075) );
  NANDN U776 ( .A(x[393]), .B(y[393]), .Z(n418) );
  NANDN U777 ( .A(x[394]), .B(y[394]), .Z(n417) );
  AND U778 ( .A(n418), .B(n417), .Z(n5063) );
  NANDN U779 ( .A(x[388]), .B(y[388]), .Z(n5051) );
  NANDN U780 ( .A(x[386]), .B(y[386]), .Z(n420) );
  NANDN U781 ( .A(x[385]), .B(y[385]), .Z(n419) );
  AND U782 ( .A(n420), .B(n419), .Z(n421) );
  NANDN U783 ( .A(x[387]), .B(y[387]), .Z(n1477) );
  NAND U784 ( .A(n421), .B(n1477), .Z(n2954) );
  NANDN U785 ( .A(y[385]), .B(x[385]), .Z(n2951) );
  NANDN U786 ( .A(y[384]), .B(x[384]), .Z(n422) );
  NAND U787 ( .A(n2951), .B(n422), .Z(n5046) );
  NANDN U788 ( .A(x[383]), .B(y[383]), .Z(n3550) );
  NANDN U789 ( .A(x[382]), .B(y[382]), .Z(n3547) );
  NANDN U790 ( .A(y[383]), .B(x[383]), .Z(n1468) );
  NANDN U791 ( .A(n3547), .B(n1468), .Z(n423) );
  NAND U792 ( .A(n3550), .B(n423), .Z(n5044) );
  NANDN U793 ( .A(x[384]), .B(y[384]), .Z(n2952) );
  NANDN U794 ( .A(y[381]), .B(x[381]), .Z(n425) );
  NANDN U795 ( .A(y[380]), .B(x[380]), .Z(n424) );
  NAND U796 ( .A(n425), .B(n424), .Z(n5037) );
  NANDN U797 ( .A(y[379]), .B(x[379]), .Z(n427) );
  NANDN U798 ( .A(y[378]), .B(x[378]), .Z(n426) );
  NAND U799 ( .A(n427), .B(n426), .Z(n5034) );
  NANDN U800 ( .A(y[375]), .B(x[375]), .Z(n429) );
  NANDN U801 ( .A(y[374]), .B(x[374]), .Z(n428) );
  NAND U802 ( .A(n429), .B(n428), .Z(n5025) );
  NANDN U803 ( .A(y[373]), .B(x[373]), .Z(n431) );
  NANDN U804 ( .A(y[372]), .B(x[372]), .Z(n430) );
  NAND U805 ( .A(n431), .B(n430), .Z(n5022) );
  ANDN U806 ( .B(x[369]), .A(y[369]), .Z(n4366) );
  NANDN U807 ( .A(y[368]), .B(x[368]), .Z(n4367) );
  NANDN U808 ( .A(n4366), .B(n4367), .Z(n3532) );
  NANDN U809 ( .A(y[367]), .B(x[367]), .Z(n438) );
  XNOR U810 ( .A(y[367]), .B(x[367]), .Z(n433) );
  NANDN U811 ( .A(x[366]), .B(y[366]), .Z(n432) );
  NAND U812 ( .A(n433), .B(n432), .Z(n434) );
  AND U813 ( .A(n438), .B(n434), .Z(n5009) );
  IV U814 ( .A(y[368]), .Z(n4368) );
  OR U815 ( .A(x[368]), .B(n4368), .Z(n435) );
  NANDN U816 ( .A(n5009), .B(n435), .Z(n3531) );
  NANDN U817 ( .A(y[366]), .B(x[366]), .Z(n437) );
  NANDN U818 ( .A(y[365]), .B(x[365]), .Z(n436) );
  AND U819 ( .A(n437), .B(n436), .Z(n439) );
  NAND U820 ( .A(n439), .B(n438), .Z(n5007) );
  NANDN U821 ( .A(x[365]), .B(y[365]), .Z(n442) );
  ANDN U822 ( .B(x[364]), .A(y[364]), .Z(n5002) );
  NAND U823 ( .A(n442), .B(n5002), .Z(n440) );
  NANDN U824 ( .A(n5007), .B(n440), .Z(n3529) );
  NANDN U825 ( .A(x[364]), .B(y[364]), .Z(n441) );
  NAND U826 ( .A(n442), .B(n441), .Z(n5005) );
  NANDN U827 ( .A(y[361]), .B(x[361]), .Z(n444) );
  NANDN U828 ( .A(y[360]), .B(x[360]), .Z(n443) );
  NAND U829 ( .A(n444), .B(n443), .Z(n4998) );
  NANDN U830 ( .A(x[359]), .B(y[359]), .Z(n446) );
  NANDN U831 ( .A(y[358]), .B(x[358]), .Z(n4989) );
  ANDN U832 ( .B(x[359]), .A(y[359]), .Z(n4993) );
  ANDN U833 ( .B(n4989), .A(n4993), .Z(n445) );
  ANDN U834 ( .B(n446), .A(n445), .Z(n3522) );
  ANDN U835 ( .B(y[357]), .A(x[357]), .Z(n4988) );
  OR U836 ( .A(n4992), .B(n4988), .Z(n3520) );
  NANDN U837 ( .A(y[355]), .B(x[355]), .Z(n448) );
  NANDN U838 ( .A(y[354]), .B(x[354]), .Z(n447) );
  NAND U839 ( .A(n448), .B(n447), .Z(n4982) );
  NANDN U840 ( .A(y[353]), .B(x[353]), .Z(n450) );
  NANDN U841 ( .A(y[352]), .B(x[352]), .Z(n449) );
  NAND U842 ( .A(n450), .B(n449), .Z(n4978) );
  NANDN U843 ( .A(x[351]), .B(y[351]), .Z(n1407) );
  ANDN U844 ( .B(y[349]), .A(x[349]), .Z(n4968) );
  OR U845 ( .A(n4972), .B(n4968), .Z(n3510) );
  NANDN U846 ( .A(y[349]), .B(x[349]), .Z(n452) );
  NANDN U847 ( .A(y[348]), .B(x[348]), .Z(n451) );
  NAND U848 ( .A(n452), .B(n451), .Z(n4966) );
  NANDN U849 ( .A(y[347]), .B(x[347]), .Z(n454) );
  NANDN U850 ( .A(y[346]), .B(x[346]), .Z(n453) );
  NAND U851 ( .A(n454), .B(n453), .Z(n4962) );
  NANDN U852 ( .A(y[343]), .B(x[343]), .Z(n456) );
  NANDN U853 ( .A(y[342]), .B(x[342]), .Z(n455) );
  NAND U854 ( .A(n456), .B(n455), .Z(n4954) );
  NANDN U855 ( .A(y[341]), .B(x[341]), .Z(n458) );
  NANDN U856 ( .A(y[340]), .B(x[340]), .Z(n457) );
  NAND U857 ( .A(n458), .B(n457), .Z(n4950) );
  NANDN U858 ( .A(y[337]), .B(x[337]), .Z(n460) );
  NANDN U859 ( .A(y[336]), .B(x[336]), .Z(n459) );
  NAND U860 ( .A(n460), .B(n459), .Z(n4942) );
  NANDN U861 ( .A(y[335]), .B(x[335]), .Z(n462) );
  NANDN U862 ( .A(y[334]), .B(x[334]), .Z(n461) );
  NAND U863 ( .A(n462), .B(n461), .Z(n4938) );
  NANDN U864 ( .A(x[331]), .B(y[331]), .Z(n464) );
  NANDN U865 ( .A(y[330]), .B(x[330]), .Z(n3486) );
  ANDN U866 ( .B(x[331]), .A(y[331]), .Z(n3489) );
  ANDN U867 ( .B(n3486), .A(n3489), .Z(n463) );
  ANDN U868 ( .B(n464), .A(n463), .Z(n4930) );
  NANDN U869 ( .A(x[329]), .B(y[329]), .Z(n3483) );
  NANDN U870 ( .A(n3488), .B(n3483), .Z(n4928) );
  NANDN U871 ( .A(y[329]), .B(x[329]), .Z(n466) );
  NANDN U872 ( .A(y[328]), .B(x[328]), .Z(n465) );
  NAND U873 ( .A(n466), .B(n465), .Z(n4926) );
  NANDN U874 ( .A(y[323]), .B(x[323]), .Z(n468) );
  NANDN U875 ( .A(y[322]), .B(x[322]), .Z(n467) );
  NAND U876 ( .A(n468), .B(n467), .Z(n4918) );
  NANDN U877 ( .A(y[321]), .B(x[321]), .Z(n470) );
  NANDN U878 ( .A(y[320]), .B(x[320]), .Z(n469) );
  NAND U879 ( .A(n470), .B(n469), .Z(n4914) );
  NANDN U880 ( .A(y[317]), .B(x[317]), .Z(n472) );
  NANDN U881 ( .A(y[316]), .B(x[316]), .Z(n471) );
  NAND U882 ( .A(n472), .B(n471), .Z(n4906) );
  NANDN U883 ( .A(y[315]), .B(x[315]), .Z(n474) );
  NANDN U884 ( .A(y[314]), .B(x[314]), .Z(n473) );
  NAND U885 ( .A(n474), .B(n473), .Z(n4902) );
  NANDN U886 ( .A(x[313]), .B(y[313]), .Z(n1319) );
  NANDN U887 ( .A(x[311]), .B(y[311]), .Z(n3461) );
  NANDN U888 ( .A(n3466), .B(n3461), .Z(n4896) );
  NANDN U889 ( .A(y[311]), .B(x[311]), .Z(n476) );
  NANDN U890 ( .A(y[310]), .B(x[310]), .Z(n475) );
  NAND U891 ( .A(n476), .B(n475), .Z(n4894) );
  NANDN U892 ( .A(y[309]), .B(x[309]), .Z(n478) );
  NANDN U893 ( .A(y[308]), .B(x[308]), .Z(n477) );
  NAND U894 ( .A(n478), .B(n477), .Z(n4890) );
  NANDN U895 ( .A(y[305]), .B(x[305]), .Z(n480) );
  NANDN U896 ( .A(y[304]), .B(x[304]), .Z(n479) );
  NAND U897 ( .A(n480), .B(n479), .Z(n4882) );
  ANDN U898 ( .B(y[303]), .A(x[303]), .Z(n483) );
  NANDN U899 ( .A(y[302]), .B(x[302]), .Z(n481) );
  ANDN U900 ( .B(x[303]), .A(y[303]), .Z(n3451) );
  ANDN U901 ( .B(n481), .A(n3451), .Z(n3448) );
  NOR U902 ( .A(n483), .B(n3448), .Z(n4878) );
  NANDN U903 ( .A(x[302]), .B(y[302]), .Z(n482) );
  NANDN U904 ( .A(n483), .B(n482), .Z(n3450) );
  NANDN U905 ( .A(x[301]), .B(y[301]), .Z(n3445) );
  NANDN U906 ( .A(n3450), .B(n3445), .Z(n4875) );
  NANDN U907 ( .A(y[299]), .B(x[299]), .Z(n485) );
  NANDN U908 ( .A(y[298]), .B(x[298]), .Z(n484) );
  NAND U909 ( .A(n485), .B(n484), .Z(n4870) );
  NANDN U910 ( .A(y[297]), .B(x[297]), .Z(n487) );
  NANDN U911 ( .A(y[296]), .B(x[296]), .Z(n486) );
  NAND U912 ( .A(n487), .B(n486), .Z(n4866) );
  ANDN U913 ( .B(y[296]), .A(x[296]), .Z(n4863) );
  NANDN U914 ( .A(x[295]), .B(y[295]), .Z(n488) );
  NANDN U915 ( .A(n4863), .B(n488), .Z(n3439) );
  NANDN U916 ( .A(y[293]), .B(x[293]), .Z(n490) );
  NANDN U917 ( .A(y[292]), .B(x[292]), .Z(n489) );
  NAND U918 ( .A(n490), .B(n489), .Z(n4854) );
  NANDN U919 ( .A(y[291]), .B(x[291]), .Z(n492) );
  NANDN U920 ( .A(y[290]), .B(x[290]), .Z(n491) );
  NAND U921 ( .A(n492), .B(n491), .Z(n4852) );
  NANDN U922 ( .A(x[287]), .B(y[287]), .Z(n495) );
  NANDN U923 ( .A(y[286]), .B(x[286]), .Z(n493) );
  ANDN U924 ( .B(x[287]), .A(y[287]), .Z(n4848) );
  ANDN U925 ( .B(n493), .A(n4848), .Z(n494) );
  ANDN U926 ( .B(n495), .A(n494), .Z(n3427) );
  ANDN U927 ( .B(y[285]), .A(x[285]), .Z(n4846) );
  OR U928 ( .A(n4847), .B(n4846), .Z(n3425) );
  NANDN U929 ( .A(y[285]), .B(x[285]), .Z(n497) );
  NANDN U930 ( .A(y[284]), .B(x[284]), .Z(n496) );
  NAND U931 ( .A(n497), .B(n496), .Z(n4845) );
  NANDN U932 ( .A(y[281]), .B(x[281]), .Z(n499) );
  NANDN U933 ( .A(y[280]), .B(x[280]), .Z(n498) );
  NAND U934 ( .A(n499), .B(n498), .Z(n4841) );
  NANDN U935 ( .A(y[279]), .B(x[279]), .Z(n501) );
  NANDN U936 ( .A(y[278]), .B(x[278]), .Z(n500) );
  NAND U937 ( .A(n501), .B(n500), .Z(n4839) );
  NANDN U938 ( .A(y[275]), .B(x[275]), .Z(n4370) );
  NANDN U939 ( .A(y[274]), .B(x[274]), .Z(n502) );
  NAND U940 ( .A(n4370), .B(n502), .Z(n4829) );
  NANDN U941 ( .A(x[275]), .B(y[275]), .Z(n503) );
  AND U942 ( .A(n4829), .B(n503), .Z(n3413) );
  ANDN U943 ( .B(y[273]), .A(x[273]), .Z(n4827) );
  OR U944 ( .A(n4827), .B(n4371), .Z(n3411) );
  NANDN U945 ( .A(y[273]), .B(x[273]), .Z(n505) );
  NANDN U946 ( .A(y[272]), .B(x[272]), .Z(n504) );
  NAND U947 ( .A(n505), .B(n504), .Z(n4825) );
  NANDN U948 ( .A(y[269]), .B(x[269]), .Z(n507) );
  NANDN U949 ( .A(y[268]), .B(x[268]), .Z(n506) );
  NAND U950 ( .A(n507), .B(n506), .Z(n4817) );
  NANDN U951 ( .A(x[267]), .B(y[267]), .Z(n509) );
  NANDN U952 ( .A(y[266]), .B(x[266]), .Z(n4808) );
  ANDN U953 ( .B(x[267]), .A(y[267]), .Z(n4812) );
  ANDN U954 ( .B(n4808), .A(n4812), .Z(n508) );
  ANDN U955 ( .B(n509), .A(n508), .Z(n3402) );
  ANDN U956 ( .B(y[265]), .A(x[265]), .Z(n4807) );
  OR U957 ( .A(n4811), .B(n4807), .Z(n3401) );
  NANDN U958 ( .A(y[263]), .B(x[263]), .Z(n511) );
  NANDN U959 ( .A(y[262]), .B(x[262]), .Z(n510) );
  NAND U960 ( .A(n511), .B(n510), .Z(n4800) );
  NANDN U961 ( .A(y[261]), .B(x[261]), .Z(n513) );
  NANDN U962 ( .A(y[260]), .B(x[260]), .Z(n512) );
  NAND U963 ( .A(n513), .B(n512), .Z(n4796) );
  NANDN U964 ( .A(y[257]), .B(x[257]), .Z(n515) );
  NANDN U965 ( .A(y[256]), .B(x[256]), .Z(n514) );
  NAND U966 ( .A(n515), .B(n514), .Z(n4789) );
  NANDN U967 ( .A(y[255]), .B(x[255]), .Z(n517) );
  NANDN U968 ( .A(y[254]), .B(x[254]), .Z(n516) );
  NAND U969 ( .A(n517), .B(n516), .Z(n4784) );
  NANDN U970 ( .A(x[251]), .B(y[251]), .Z(n1196) );
  XNOR U971 ( .A(x[251]), .B(y[251]), .Z(n519) );
  NANDN U972 ( .A(y[250]), .B(x[250]), .Z(n518) );
  NAND U973 ( .A(n519), .B(n518), .Z(n520) );
  AND U974 ( .A(n1196), .B(n520), .Z(n4777) );
  NANDN U975 ( .A(y[249]), .B(x[249]), .Z(n522) );
  NANDN U976 ( .A(y[248]), .B(x[248]), .Z(n521) );
  NAND U977 ( .A(n522), .B(n521), .Z(n4772) );
  NANDN U978 ( .A(y[245]), .B(x[245]), .Z(n524) );
  NANDN U979 ( .A(y[244]), .B(x[244]), .Z(n523) );
  NAND U980 ( .A(n524), .B(n523), .Z(n4765) );
  ANDN U981 ( .B(y[243]), .A(x[243]), .Z(n526) );
  NANDN U982 ( .A(y[242]), .B(x[242]), .Z(n3373) );
  ANDN U983 ( .B(x[243]), .A(y[243]), .Z(n3376) );
  ANDN U984 ( .B(n3373), .A(n3376), .Z(n525) );
  NOR U985 ( .A(n526), .B(n525), .Z(n4760) );
  NANDN U986 ( .A(x[241]), .B(y[241]), .Z(n3370) );
  NANDN U987 ( .A(n3375), .B(n3370), .Z(n4759) );
  NANDN U988 ( .A(y[239]), .B(x[239]), .Z(n528) );
  NANDN U989 ( .A(y[238]), .B(x[238]), .Z(n527) );
  NAND U990 ( .A(n528), .B(n527), .Z(n4753) );
  NANDN U991 ( .A(y[237]), .B(x[237]), .Z(n530) );
  NANDN U992 ( .A(y[236]), .B(x[236]), .Z(n529) );
  NAND U993 ( .A(n530), .B(n529), .Z(n4748) );
  NANDN U994 ( .A(y[233]), .B(x[233]), .Z(n532) );
  NANDN U995 ( .A(y[232]), .B(x[232]), .Z(n531) );
  NAND U996 ( .A(n532), .B(n531), .Z(n4741) );
  NANDN U997 ( .A(x[231]), .B(y[231]), .Z(n534) );
  NANDN U998 ( .A(y[230]), .B(x[230]), .Z(n4732) );
  ANDN U999 ( .B(x[231]), .A(y[231]), .Z(n4736) );
  ANDN U1000 ( .B(n4732), .A(n4736), .Z(n533) );
  ANDN U1001 ( .B(n534), .A(n533), .Z(n3358) );
  ANDN U1002 ( .B(y[229]), .A(x[229]), .Z(n4731) );
  OR U1003 ( .A(n4735), .B(n4731), .Z(n3357) );
  NANDN U1004 ( .A(y[227]), .B(x[227]), .Z(n536) );
  NANDN U1005 ( .A(y[226]), .B(x[226]), .Z(n535) );
  NAND U1006 ( .A(n536), .B(n535), .Z(n4724) );
  NANDN U1007 ( .A(y[225]), .B(x[225]), .Z(n538) );
  NANDN U1008 ( .A(y[224]), .B(x[224]), .Z(n537) );
  NAND U1009 ( .A(n538), .B(n537), .Z(n4720) );
  NANDN U1010 ( .A(y[221]), .B(x[221]), .Z(n540) );
  NANDN U1011 ( .A(y[220]), .B(x[220]), .Z(n539) );
  NAND U1012 ( .A(n540), .B(n539), .Z(n4713) );
  NANDN U1013 ( .A(y[219]), .B(x[219]), .Z(n542) );
  NANDN U1014 ( .A(y[218]), .B(x[218]), .Z(n541) );
  NAND U1015 ( .A(n542), .B(n541), .Z(n4708) );
  NANDN U1016 ( .A(x[218]), .B(y[218]), .Z(n544) );
  NANDN U1017 ( .A(x[217]), .B(y[217]), .Z(n543) );
  NAND U1018 ( .A(n544), .B(n543), .Z(n2958) );
  NANDN U1019 ( .A(y[217]), .B(x[217]), .Z(n2955) );
  NANDN U1020 ( .A(y[216]), .B(x[216]), .Z(n545) );
  NAND U1021 ( .A(n2955), .B(n545), .Z(n4705) );
  NANDN U1022 ( .A(x[216]), .B(y[216]), .Z(n2956) );
  NANDN U1023 ( .A(x[211]), .B(y[211]), .Z(n547) );
  NANDN U1024 ( .A(x[212]), .B(y[212]), .Z(n546) );
  AND U1025 ( .A(n547), .B(n546), .Z(n4694) );
  NANDN U1026 ( .A(x[205]), .B(y[205]), .Z(n549) );
  NANDN U1027 ( .A(x[206]), .B(y[206]), .Z(n548) );
  AND U1028 ( .A(n549), .B(n548), .Z(n4682) );
  NANDN U1029 ( .A(x[193]), .B(y[193]), .Z(n551) );
  NANDN U1030 ( .A(x[194]), .B(y[194]), .Z(n550) );
  AND U1031 ( .A(n551), .B(n550), .Z(n4658) );
  NANDN U1032 ( .A(x[187]), .B(y[187]), .Z(n553) );
  NANDN U1033 ( .A(x[188]), .B(y[188]), .Z(n552) );
  AND U1034 ( .A(n553), .B(n552), .Z(n4646) );
  NANDN U1035 ( .A(x[181]), .B(y[181]), .Z(n555) );
  NANDN U1036 ( .A(x[182]), .B(y[182]), .Z(n554) );
  AND U1037 ( .A(n555), .B(n554), .Z(n4634) );
  NANDN U1038 ( .A(x[179]), .B(y[179]), .Z(n557) );
  NANDN U1039 ( .A(y[178]), .B(x[178]), .Z(n3295) );
  ANDN U1040 ( .B(x[179]), .A(y[179]), .Z(n3298) );
  ANDN U1041 ( .B(n3295), .A(n3298), .Z(n556) );
  ANDN U1042 ( .B(n557), .A(n556), .Z(n4629) );
  NANDN U1043 ( .A(x[177]), .B(y[177]), .Z(n3292) );
  NANDN U1044 ( .A(n3297), .B(n3292), .Z(n4627) );
  NANDN U1045 ( .A(y[175]), .B(x[175]), .Z(n2959) );
  NANDN U1046 ( .A(y[174]), .B(x[174]), .Z(n558) );
  NAND U1047 ( .A(n2959), .B(n558), .Z(n4621) );
  NANDN U1048 ( .A(x[174]), .B(y[174]), .Z(n2960) );
  ANDN U1049 ( .B(y[165]), .A(x[165]), .Z(n4596) );
  NANDN U1050 ( .A(x[166]), .B(y[166]), .Z(n4600) );
  NANDN U1051 ( .A(n4596), .B(n4600), .Z(n3278) );
  NANDN U1052 ( .A(y[162]), .B(x[162]), .Z(n3270) );
  ANDN U1053 ( .B(x[163]), .A(y[163]), .Z(n3273) );
  ANDN U1054 ( .B(n3270), .A(n3273), .Z(n559) );
  ANDN U1055 ( .B(y[163]), .A(x[163]), .Z(n996) );
  NOR U1056 ( .A(n559), .B(n996), .Z(n4590) );
  NANDN U1057 ( .A(x[160]), .B(y[160]), .Z(n561) );
  NANDN U1058 ( .A(x[159]), .B(y[159]), .Z(n560) );
  NAND U1059 ( .A(n561), .B(n560), .Z(n2966) );
  NANDN U1060 ( .A(x[158]), .B(y[158]), .Z(n2964) );
  NANDN U1061 ( .A(y[155]), .B(x[155]), .Z(n563) );
  NANDN U1062 ( .A(y[154]), .B(x[154]), .Z(n562) );
  NAND U1063 ( .A(n563), .B(n562), .Z(n4574) );
  NANDN U1064 ( .A(x[153]), .B(y[153]), .Z(n565) );
  NANDN U1065 ( .A(x[154]), .B(y[154]), .Z(n564) );
  AND U1066 ( .A(n565), .B(n564), .Z(n4571) );
  ANDN U1067 ( .B(x[153]), .A(y[153]), .Z(n4373) );
  NANDN U1068 ( .A(y[152]), .B(x[152]), .Z(n4374) );
  NANDN U1069 ( .A(n4373), .B(n4374), .Z(n3257) );
  ANDN U1070 ( .B(y[151]), .A(x[151]), .Z(n4565) );
  NANDN U1071 ( .A(x[152]), .B(y[152]), .Z(n566) );
  NANDN U1072 ( .A(n4565), .B(n566), .Z(n3256) );
  NANDN U1073 ( .A(x[147]), .B(y[147]), .Z(n568) );
  NANDN U1074 ( .A(x[148]), .B(y[148]), .Z(n567) );
  AND U1075 ( .A(n568), .B(n567), .Z(n4557) );
  ANDN U1076 ( .B(x[143]), .A(y[143]), .Z(n4548) );
  ANDN U1077 ( .B(y[143]), .A(x[143]), .Z(n570) );
  ANDN U1078 ( .B(x[142]), .A(y[142]), .Z(n4544) );
  NANDN U1079 ( .A(n570), .B(n4544), .Z(n569) );
  NANDN U1080 ( .A(n4548), .B(n569), .Z(n3246) );
  NANDN U1081 ( .A(x[142]), .B(y[142]), .Z(n571) );
  ANDN U1082 ( .B(n571), .A(n570), .Z(n4545) );
  NANDN U1083 ( .A(x[141]), .B(y[141]), .Z(n574) );
  NANDN U1084 ( .A(y[141]), .B(x[141]), .Z(n3242) );
  NANDN U1085 ( .A(y[140]), .B(x[140]), .Z(n572) );
  AND U1086 ( .A(n3242), .B(n572), .Z(n573) );
  ANDN U1087 ( .B(n574), .A(n573), .Z(n4542) );
  NANDN U1088 ( .A(x[139]), .B(y[139]), .Z(n3237) );
  NANDN U1089 ( .A(n3241), .B(n3237), .Z(n4540) );
  NANDN U1090 ( .A(x[138]), .B(y[138]), .Z(n576) );
  NANDN U1091 ( .A(x[137]), .B(y[137]), .Z(n575) );
  NAND U1092 ( .A(n576), .B(n575), .Z(n4535) );
  ANDN U1093 ( .B(x[135]), .A(y[135]), .Z(n4375) );
  NANDN U1094 ( .A(y[134]), .B(x[134]), .Z(n4376) );
  NANDN U1095 ( .A(n4375), .B(n4376), .Z(n3231) );
  ANDN U1096 ( .B(y[133]), .A(x[133]), .Z(n4525) );
  NANDN U1097 ( .A(x[134]), .B(y[134]), .Z(n577) );
  NANDN U1098 ( .A(n4525), .B(n577), .Z(n3229) );
  NANDN U1099 ( .A(x[132]), .B(y[132]), .Z(n579) );
  NANDN U1100 ( .A(x[131]), .B(y[131]), .Z(n578) );
  NAND U1101 ( .A(n579), .B(n578), .Z(n4522) );
  NANDN U1102 ( .A(x[130]), .B(y[130]), .Z(n4517) );
  NANDN U1103 ( .A(y[129]), .B(x[129]), .Z(n3222) );
  NANDN U1104 ( .A(y[128]), .B(x[128]), .Z(n580) );
  AND U1105 ( .A(n3222), .B(n580), .Z(n581) );
  ANDN U1106 ( .B(y[129]), .A(x[129]), .Z(n582) );
  NOR U1107 ( .A(n581), .B(n582), .Z(n4516) );
  NANDN U1108 ( .A(x[127]), .B(y[127]), .Z(n3217) );
  NANDN U1109 ( .A(n3221), .B(n3217), .Z(n4513) );
  NANDN U1110 ( .A(x[125]), .B(y[125]), .Z(n925) );
  NANDN U1111 ( .A(y[124]), .B(x[124]), .Z(n583) );
  ANDN U1112 ( .B(x[125]), .A(y[125]), .Z(n4508) );
  ANDN U1113 ( .B(n583), .A(n4508), .Z(n584) );
  ANDN U1114 ( .B(n925), .A(n584), .Z(n3213) );
  NANDN U1115 ( .A(x[122]), .B(y[122]), .Z(n586) );
  NANDN U1116 ( .A(x[121]), .B(y[121]), .Z(n585) );
  NAND U1117 ( .A(n586), .B(n585), .Z(n2970) );
  NANDN U1118 ( .A(y[121]), .B(x[121]), .Z(n2967) );
  NANDN U1119 ( .A(y[120]), .B(x[120]), .Z(n587) );
  NAND U1120 ( .A(n2967), .B(n587), .Z(n4496) );
  NANDN U1121 ( .A(x[120]), .B(y[120]), .Z(n2968) );
  NANDN U1122 ( .A(x[118]), .B(y[118]), .Z(n589) );
  NANDN U1123 ( .A(x[117]), .B(y[117]), .Z(n588) );
  NAND U1124 ( .A(n589), .B(n588), .Z(n4490) );
  NANDN U1125 ( .A(x[113]), .B(y[113]), .Z(n591) );
  NANDN U1126 ( .A(y[112]), .B(x[112]), .Z(n4476) );
  ANDN U1127 ( .B(x[113]), .A(y[113]), .Z(n4479) );
  ANDN U1128 ( .B(n4476), .A(n4479), .Z(n590) );
  ANDN U1129 ( .B(n591), .A(n590), .Z(n3199) );
  ANDN U1130 ( .B(y[111]), .A(x[111]), .Z(n4474) );
  OR U1131 ( .A(n4478), .B(n4474), .Z(n3197) );
  NANDN U1132 ( .A(x[108]), .B(y[108]), .Z(n593) );
  NANDN U1133 ( .A(x[107]), .B(y[107]), .Z(n592) );
  NAND U1134 ( .A(n593), .B(n592), .Z(n4465) );
  NANDN U1135 ( .A(x[106]), .B(y[106]), .Z(n595) );
  NANDN U1136 ( .A(x[105]), .B(y[105]), .Z(n594) );
  NAND U1137 ( .A(n595), .B(n594), .Z(n2974) );
  ANDN U1138 ( .B(y[104]), .A(x[104]), .Z(n2971) );
  NANDN U1139 ( .A(y[103]), .B(x[103]), .Z(n600) );
  XNOR U1140 ( .A(y[103]), .B(x[103]), .Z(n597) );
  NANDN U1141 ( .A(x[102]), .B(y[102]), .Z(n596) );
  NAND U1142 ( .A(n597), .B(n596), .Z(n598) );
  AND U1143 ( .A(n600), .B(n598), .Z(n4458) );
  NOR U1144 ( .A(n2971), .B(n4458), .Z(n885) );
  NANDN U1145 ( .A(y[102]), .B(x[102]), .Z(n599) );
  NAND U1146 ( .A(n600), .B(n599), .Z(n4455) );
  NANDN U1147 ( .A(y[100]), .B(x[100]), .Z(n601) );
  ANDN U1148 ( .B(x[101]), .A(y[101]), .Z(n4454) );
  ANDN U1149 ( .B(n601), .A(n4454), .Z(n602) );
  NANDN U1150 ( .A(x[101]), .B(y[101]), .Z(n881) );
  NANDN U1151 ( .A(n602), .B(n881), .Z(n603) );
  NANDN U1152 ( .A(n4455), .B(n603), .Z(n3186) );
  NANDN U1153 ( .A(x[98]), .B(y[98]), .Z(n605) );
  NANDN U1154 ( .A(x[97]), .B(y[97]), .Z(n604) );
  NAND U1155 ( .A(n605), .B(n604), .Z(n4444) );
  NANDN U1156 ( .A(x[96]), .B(y[96]), .Z(n607) );
  NANDN U1157 ( .A(x[95]), .B(y[95]), .Z(n606) );
  NAND U1158 ( .A(n607), .B(n606), .Z(n4439) );
  NANDN U1159 ( .A(x[92]), .B(y[92]), .Z(n609) );
  NANDN U1160 ( .A(x[91]), .B(y[91]), .Z(n608) );
  NAND U1161 ( .A(n609), .B(n608), .Z(n4432) );
  NANDN U1162 ( .A(x[90]), .B(y[90]), .Z(n611) );
  NANDN U1163 ( .A(x[89]), .B(y[89]), .Z(n610) );
  NAND U1164 ( .A(n611), .B(n610), .Z(n4427) );
  NANDN U1165 ( .A(x[88]), .B(y[88]), .Z(n4423) );
  NANDN U1166 ( .A(x[87]), .B(y[87]), .Z(n614) );
  NANDN U1167 ( .A(y[86]), .B(x[86]), .Z(n612) );
  ANDN U1168 ( .B(x[87]), .A(y[87]), .Z(n4422) );
  ANDN U1169 ( .B(n612), .A(n4422), .Z(n613) );
  ANDN U1170 ( .B(n614), .A(n613), .Z(n3171) );
  ANDN U1171 ( .B(y[85]), .A(x[85]), .Z(n4415) );
  OR U1172 ( .A(n4420), .B(n4415), .Z(n3169) );
  NANDN U1173 ( .A(x[84]), .B(y[84]), .Z(n616) );
  NANDN U1174 ( .A(x[83]), .B(y[83]), .Z(n615) );
  NAND U1175 ( .A(n616), .B(n615), .Z(n4411) );
  NANDN U1176 ( .A(x[80]), .B(y[80]), .Z(n618) );
  NANDN U1177 ( .A(x[79]), .B(y[79]), .Z(n617) );
  NAND U1178 ( .A(n618), .B(n617), .Z(n4404) );
  NANDN U1179 ( .A(x[78]), .B(y[78]), .Z(n620) );
  NANDN U1180 ( .A(x[77]), .B(y[77]), .Z(n619) );
  NAND U1181 ( .A(n620), .B(n619), .Z(n4399) );
  NANDN U1182 ( .A(x[74]), .B(y[74]), .Z(n622) );
  NANDN U1183 ( .A(x[73]), .B(y[73]), .Z(n621) );
  NAND U1184 ( .A(n622), .B(n621), .Z(n4392) );
  NANDN U1185 ( .A(x[72]), .B(y[72]), .Z(n624) );
  NANDN U1186 ( .A(x[71]), .B(y[71]), .Z(n623) );
  NAND U1187 ( .A(n624), .B(n623), .Z(n4387) );
  NANDN U1188 ( .A(x[70]), .B(y[70]), .Z(n4383) );
  NANDN U1189 ( .A(x[69]), .B(y[69]), .Z(n627) );
  NANDN U1190 ( .A(y[68]), .B(x[68]), .Z(n625) );
  ANDN U1191 ( .B(x[69]), .A(y[69]), .Z(n4382) );
  ANDN U1192 ( .B(n625), .A(n4382), .Z(n626) );
  ANDN U1193 ( .B(n627), .A(n626), .Z(n3151) );
  NANDN U1194 ( .A(y[67]), .B(x[67]), .Z(n629) );
  NANDN U1195 ( .A(y[66]), .B(x[66]), .Z(n628) );
  NAND U1196 ( .A(n629), .B(n628), .Z(n3147) );
  NANDN U1197 ( .A(x[66]), .B(y[66]), .Z(n631) );
  NANDN U1198 ( .A(x[65]), .B(y[65]), .Z(n630) );
  NAND U1199 ( .A(n631), .B(n630), .Z(n3145) );
  NANDN U1200 ( .A(y[64]), .B(x[64]), .Z(n633) );
  NANDN U1201 ( .A(y[65]), .B(x[65]), .Z(n632) );
  NAND U1202 ( .A(n633), .B(n632), .Z(n3143) );
  NANDN U1203 ( .A(x[64]), .B(y[64]), .Z(n635) );
  NANDN U1204 ( .A(x[63]), .B(y[63]), .Z(n634) );
  NAND U1205 ( .A(n635), .B(n634), .Z(n3140) );
  NANDN U1206 ( .A(y[62]), .B(x[62]), .Z(n637) );
  NANDN U1207 ( .A(y[63]), .B(x[63]), .Z(n636) );
  NAND U1208 ( .A(n637), .B(n636), .Z(n3139) );
  NANDN U1209 ( .A(y[60]), .B(x[60]), .Z(n639) );
  NANDN U1210 ( .A(y[61]), .B(x[61]), .Z(n638) );
  NAND U1211 ( .A(n639), .B(n638), .Z(n3135) );
  NANDN U1212 ( .A(x[60]), .B(y[60]), .Z(n641) );
  NANDN U1213 ( .A(x[59]), .B(y[59]), .Z(n640) );
  NAND U1214 ( .A(n641), .B(n640), .Z(n3133) );
  NANDN U1215 ( .A(y[58]), .B(x[58]), .Z(n643) );
  NANDN U1216 ( .A(y[59]), .B(x[59]), .Z(n642) );
  NAND U1217 ( .A(n643), .B(n642), .Z(n3131) );
  NANDN U1218 ( .A(x[58]), .B(y[58]), .Z(n645) );
  NANDN U1219 ( .A(x[57]), .B(y[57]), .Z(n644) );
  NAND U1220 ( .A(n645), .B(n644), .Z(n3128) );
  NANDN U1221 ( .A(y[56]), .B(x[56]), .Z(n647) );
  NANDN U1222 ( .A(y[57]), .B(x[57]), .Z(n646) );
  NAND U1223 ( .A(n647), .B(n646), .Z(n3127) );
  NANDN U1224 ( .A(y[54]), .B(x[54]), .Z(n649) );
  NANDN U1225 ( .A(y[55]), .B(x[55]), .Z(n648) );
  NAND U1226 ( .A(n649), .B(n648), .Z(n3123) );
  NANDN U1227 ( .A(x[54]), .B(y[54]), .Z(n651) );
  NANDN U1228 ( .A(x[53]), .B(y[53]), .Z(n650) );
  NAND U1229 ( .A(n651), .B(n650), .Z(n3121) );
  NANDN U1230 ( .A(y[52]), .B(x[52]), .Z(n653) );
  NANDN U1231 ( .A(y[53]), .B(x[53]), .Z(n652) );
  NAND U1232 ( .A(n653), .B(n652), .Z(n3119) );
  NANDN U1233 ( .A(x[52]), .B(y[52]), .Z(n655) );
  NANDN U1234 ( .A(x[51]), .B(y[51]), .Z(n654) );
  NAND U1235 ( .A(n655), .B(n654), .Z(n3116) );
  NANDN U1236 ( .A(y[50]), .B(x[50]), .Z(n657) );
  NANDN U1237 ( .A(y[51]), .B(x[51]), .Z(n656) );
  NAND U1238 ( .A(n657), .B(n656), .Z(n3115) );
  NANDN U1239 ( .A(y[48]), .B(x[48]), .Z(n659) );
  NANDN U1240 ( .A(y[49]), .B(x[49]), .Z(n658) );
  NAND U1241 ( .A(n659), .B(n658), .Z(n3111) );
  NANDN U1242 ( .A(x[48]), .B(y[48]), .Z(n661) );
  NANDN U1243 ( .A(x[47]), .B(y[47]), .Z(n660) );
  NAND U1244 ( .A(n661), .B(n660), .Z(n3109) );
  NANDN U1245 ( .A(y[46]), .B(x[46]), .Z(n663) );
  NANDN U1246 ( .A(y[47]), .B(x[47]), .Z(n662) );
  NAND U1247 ( .A(n663), .B(n662), .Z(n3107) );
  NANDN U1248 ( .A(x[46]), .B(y[46]), .Z(n665) );
  NANDN U1249 ( .A(x[45]), .B(y[45]), .Z(n664) );
  NAND U1250 ( .A(n665), .B(n664), .Z(n3104) );
  NANDN U1251 ( .A(y[44]), .B(x[44]), .Z(n667) );
  NANDN U1252 ( .A(y[45]), .B(x[45]), .Z(n666) );
  NAND U1253 ( .A(n667), .B(n666), .Z(n3103) );
  NANDN U1254 ( .A(y[42]), .B(x[42]), .Z(n669) );
  NANDN U1255 ( .A(y[43]), .B(x[43]), .Z(n668) );
  NAND U1256 ( .A(n669), .B(n668), .Z(n3099) );
  NANDN U1257 ( .A(x[42]), .B(y[42]), .Z(n671) );
  NANDN U1258 ( .A(x[41]), .B(y[41]), .Z(n670) );
  NAND U1259 ( .A(n671), .B(n670), .Z(n3097) );
  NANDN U1260 ( .A(y[40]), .B(x[40]), .Z(n673) );
  NANDN U1261 ( .A(y[41]), .B(x[41]), .Z(n672) );
  NAND U1262 ( .A(n673), .B(n672), .Z(n3095) );
  NANDN U1263 ( .A(x[40]), .B(y[40]), .Z(n675) );
  NANDN U1264 ( .A(x[39]), .B(y[39]), .Z(n674) );
  NAND U1265 ( .A(n675), .B(n674), .Z(n3092) );
  NANDN U1266 ( .A(y[38]), .B(x[38]), .Z(n677) );
  NANDN U1267 ( .A(y[39]), .B(x[39]), .Z(n676) );
  NAND U1268 ( .A(n677), .B(n676), .Z(n3091) );
  IV U1269 ( .A(y[36]), .Z(n3083) );
  OR U1270 ( .A(x[36]), .B(n3083), .Z(n769) );
  NANDN U1271 ( .A(y[35]), .B(x[35]), .Z(n679) );
  NANDN U1272 ( .A(y[34]), .B(x[34]), .Z(n678) );
  NAND U1273 ( .A(n679), .B(n678), .Z(n3078) );
  NANDN U1274 ( .A(x[34]), .B(y[34]), .Z(n681) );
  NANDN U1275 ( .A(x[33]), .B(y[33]), .Z(n680) );
  NAND U1276 ( .A(n681), .B(n680), .Z(n3075) );
  NANDN U1277 ( .A(y[32]), .B(x[32]), .Z(n683) );
  NANDN U1278 ( .A(y[33]), .B(x[33]), .Z(n682) );
  NAND U1279 ( .A(n683), .B(n682), .Z(n3074) );
  NANDN U1280 ( .A(x[32]), .B(y[32]), .Z(n685) );
  NANDN U1281 ( .A(x[31]), .B(y[31]), .Z(n684) );
  NAND U1282 ( .A(n685), .B(n684), .Z(n3072) );
  NANDN U1283 ( .A(y[30]), .B(x[30]), .Z(n687) );
  NANDN U1284 ( .A(y[31]), .B(x[31]), .Z(n686) );
  NAND U1285 ( .A(n687), .B(n686), .Z(n3070) );
  NANDN U1286 ( .A(y[28]), .B(x[28]), .Z(n689) );
  NANDN U1287 ( .A(y[29]), .B(x[29]), .Z(n688) );
  NAND U1288 ( .A(n689), .B(n688), .Z(n3066) );
  NANDN U1289 ( .A(x[28]), .B(y[28]), .Z(n691) );
  NANDN U1290 ( .A(x[27]), .B(y[27]), .Z(n690) );
  NAND U1291 ( .A(n691), .B(n690), .Z(n3063) );
  NANDN U1292 ( .A(y[26]), .B(x[26]), .Z(n693) );
  NANDN U1293 ( .A(y[27]), .B(x[27]), .Z(n692) );
  NAND U1294 ( .A(n693), .B(n692), .Z(n3062) );
  NANDN U1295 ( .A(x[26]), .B(y[26]), .Z(n695) );
  NANDN U1296 ( .A(x[25]), .B(y[25]), .Z(n694) );
  NAND U1297 ( .A(n695), .B(n694), .Z(n3060) );
  NANDN U1298 ( .A(y[24]), .B(x[24]), .Z(n697) );
  NANDN U1299 ( .A(y[25]), .B(x[25]), .Z(n696) );
  NAND U1300 ( .A(n697), .B(n696), .Z(n3058) );
  NANDN U1301 ( .A(y[22]), .B(x[22]), .Z(n699) );
  NANDN U1302 ( .A(y[23]), .B(x[23]), .Z(n698) );
  NAND U1303 ( .A(n699), .B(n698), .Z(n3054) );
  NANDN U1304 ( .A(x[22]), .B(y[22]), .Z(n701) );
  NANDN U1305 ( .A(x[21]), .B(y[21]), .Z(n700) );
  NAND U1306 ( .A(n701), .B(n700), .Z(n3051) );
  NANDN U1307 ( .A(y[21]), .B(x[21]), .Z(n3048) );
  ANDN U1308 ( .B(y[18]), .A(x[18]), .Z(n2975) );
  ANDN U1309 ( .B(x[17]), .A(y[17]), .Z(n3034) );
  ANDN U1310 ( .B(y[16]), .A(x[16]), .Z(n2977) );
  NANDN U1311 ( .A(x[17]), .B(y[17]), .Z(n2976) );
  ANDN U1312 ( .B(x[15]), .A(y[15]), .Z(n3027) );
  ANDN U1313 ( .B(x[16]), .A(y[16]), .Z(n3036) );
  ANDN U1314 ( .B(y[14]), .A(x[14]), .Z(n3023) );
  ANDN U1315 ( .B(x[13]), .A(y[13]), .Z(n3022) );
  ANDN U1316 ( .B(y[12]), .A(x[12]), .Z(n3017) );
  NANDN U1317 ( .A(y[9]), .B(x[9]), .Z(n703) );
  NANDN U1318 ( .A(y[10]), .B(x[10]), .Z(n702) );
  NAND U1319 ( .A(n703), .B(n702), .Z(n3012) );
  NANDN U1320 ( .A(x[9]), .B(y[9]), .Z(n705) );
  NANDN U1321 ( .A(x[8]), .B(y[8]), .Z(n704) );
  NAND U1322 ( .A(n705), .B(n704), .Z(n3007) );
  ANDN U1323 ( .B(x[8]), .A(y[8]), .Z(n2980) );
  NANDN U1324 ( .A(y[7]), .B(x[7]), .Z(n706) );
  NANDN U1325 ( .A(n2980), .B(n706), .Z(n3003) );
  ANDN U1326 ( .B(x[5]), .A(y[5]), .Z(n2998) );
  NANDN U1327 ( .A(x[5]), .B(y[5]), .Z(n3001) );
  ANDN U1328 ( .B(x[3]), .A(y[3]), .Z(n2992) );
  NANDN U1329 ( .A(y[1]), .B(x[1]), .Z(n707) );
  ANDN U1330 ( .B(x[2]), .A(y[2]), .Z(n2990) );
  ANDN U1331 ( .B(n707), .A(n2990), .Z(n710) );
  NANDN U1332 ( .A(x[0]), .B(y[0]), .Z(n708) );
  NAND U1333 ( .A(n708), .B(n2986), .Z(n709) );
  AND U1334 ( .A(n710), .B(n709), .Z(n712) );
  NANDN U1335 ( .A(x[2]), .B(y[2]), .Z(n2985) );
  ANDN U1336 ( .B(y[3]), .A(x[3]), .Z(n2981) );
  ANDN U1337 ( .B(n2985), .A(n2981), .Z(n711) );
  NANDN U1338 ( .A(n712), .B(n711), .Z(n713) );
  ANDN U1339 ( .B(x[4]), .A(y[4]), .Z(n2995) );
  ANDN U1340 ( .B(n713), .A(n2995), .Z(n714) );
  NANDN U1341 ( .A(n2992), .B(n714), .Z(n715) );
  AND U1342 ( .A(n3001), .B(n715), .Z(n716) );
  NANDN U1343 ( .A(x[4]), .B(y[4]), .Z(n2982) );
  NAND U1344 ( .A(n716), .B(n2982), .Z(n717) );
  NANDN U1345 ( .A(n2998), .B(n717), .Z(n719) );
  ANDN U1346 ( .B(x[6]), .A(y[6]), .Z(n718) );
  OR U1347 ( .A(n719), .B(n718), .Z(n721) );
  ANDN U1348 ( .B(y[7]), .A(x[7]), .Z(n2979) );
  ANDN U1349 ( .B(y[6]), .A(x[6]), .Z(n2999) );
  NOR U1350 ( .A(n2979), .B(n2999), .Z(n720) );
  NAND U1351 ( .A(n721), .B(n720), .Z(n722) );
  NANDN U1352 ( .A(n3003), .B(n722), .Z(n723) );
  NANDN U1353 ( .A(n3007), .B(n723), .Z(n724) );
  NANDN U1354 ( .A(n3012), .B(n724), .Z(n727) );
  NANDN U1355 ( .A(x[10]), .B(y[10]), .Z(n726) );
  NANDN U1356 ( .A(x[11]), .B(y[11]), .Z(n725) );
  NAND U1357 ( .A(n726), .B(n725), .Z(n3014) );
  ANDN U1358 ( .B(n727), .A(n3014), .Z(n729) );
  ANDN U1359 ( .B(x[11]), .A(y[11]), .Z(n3016) );
  ANDN U1360 ( .B(x[12]), .A(y[12]), .Z(n3019) );
  NOR U1361 ( .A(n3016), .B(n3019), .Z(n728) );
  NANDN U1362 ( .A(n729), .B(n728), .Z(n730) );
  ANDN U1363 ( .B(y[13]), .A(x[13]), .Z(n3026) );
  ANDN U1364 ( .B(n730), .A(n3026), .Z(n731) );
  NANDN U1365 ( .A(n3017), .B(n731), .Z(n732) );
  ANDN U1366 ( .B(x[14]), .A(y[14]), .Z(n3030) );
  ANDN U1367 ( .B(n732), .A(n3030), .Z(n733) );
  NANDN U1368 ( .A(n3022), .B(n733), .Z(n734) );
  NANDN U1369 ( .A(x[15]), .B(y[15]), .Z(n2978) );
  AND U1370 ( .A(n734), .B(n2978), .Z(n735) );
  NANDN U1371 ( .A(n3023), .B(n735), .Z(n736) );
  NANDN U1372 ( .A(n3036), .B(n736), .Z(n737) );
  OR U1373 ( .A(n3027), .B(n737), .Z(n738) );
  AND U1374 ( .A(n2976), .B(n738), .Z(n739) );
  NANDN U1375 ( .A(n2977), .B(n739), .Z(n740) );
  ANDN U1376 ( .B(x[18]), .A(y[18]), .Z(n3039) );
  ANDN U1377 ( .B(n740), .A(n3039), .Z(n741) );
  NANDN U1378 ( .A(n3034), .B(n741), .Z(n742) );
  ANDN U1379 ( .B(y[19]), .A(x[19]), .Z(n3046) );
  ANDN U1380 ( .B(n742), .A(n3046), .Z(n743) );
  NANDN U1381 ( .A(n2975), .B(n743), .Z(n744) );
  ANDN U1382 ( .B(x[19]), .A(y[19]), .Z(n3042) );
  ANDN U1383 ( .B(n744), .A(n3042), .Z(n746) );
  OR U1384 ( .A(n746), .B(y[20]), .Z(n745) );
  AND U1385 ( .A(n3048), .B(n745), .Z(n749) );
  XOR U1386 ( .A(n746), .B(y[20]), .Z(n747) );
  NAND U1387 ( .A(n747), .B(x[20]), .Z(n748) );
  NAND U1388 ( .A(n749), .B(n748), .Z(n750) );
  NANDN U1389 ( .A(n3051), .B(n750), .Z(n751) );
  NANDN U1390 ( .A(n3054), .B(n751), .Z(n754) );
  NANDN U1391 ( .A(x[24]), .B(y[24]), .Z(n753) );
  NANDN U1392 ( .A(x[23]), .B(y[23]), .Z(n752) );
  NAND U1393 ( .A(n753), .B(n752), .Z(n3056) );
  ANDN U1394 ( .B(n754), .A(n3056), .Z(n755) );
  OR U1395 ( .A(n3058), .B(n755), .Z(n756) );
  NANDN U1396 ( .A(n3060), .B(n756), .Z(n757) );
  NANDN U1397 ( .A(n3062), .B(n757), .Z(n758) );
  NANDN U1398 ( .A(n3063), .B(n758), .Z(n759) );
  NANDN U1399 ( .A(n3066), .B(n759), .Z(n762) );
  NANDN U1400 ( .A(x[30]), .B(y[30]), .Z(n761) );
  NANDN U1401 ( .A(x[29]), .B(y[29]), .Z(n760) );
  NAND U1402 ( .A(n761), .B(n760), .Z(n3068) );
  ANDN U1403 ( .B(n762), .A(n3068), .Z(n763) );
  OR U1404 ( .A(n3070), .B(n763), .Z(n764) );
  NANDN U1405 ( .A(n3072), .B(n764), .Z(n765) );
  NANDN U1406 ( .A(n3074), .B(n765), .Z(n766) );
  NANDN U1407 ( .A(n3075), .B(n766), .Z(n767) );
  NANDN U1408 ( .A(n3078), .B(n767), .Z(n768) );
  AND U1409 ( .A(n769), .B(n768), .Z(n770) );
  NANDN U1410 ( .A(x[35]), .B(y[35]), .Z(n3079) );
  NAND U1411 ( .A(n770), .B(n3079), .Z(n773) );
  NANDN U1412 ( .A(y[36]), .B(x[36]), .Z(n771) );
  ANDN U1413 ( .B(x[37]), .A(y[37]), .Z(n3081) );
  ANDN U1414 ( .B(n771), .A(n3081), .Z(n772) );
  NAND U1415 ( .A(n773), .B(n772), .Z(n776) );
  NANDN U1416 ( .A(x[38]), .B(y[38]), .Z(n775) );
  NANDN U1417 ( .A(x[37]), .B(y[37]), .Z(n774) );
  NAND U1418 ( .A(n775), .B(n774), .Z(n3089) );
  ANDN U1419 ( .B(n776), .A(n3089), .Z(n777) );
  OR U1420 ( .A(n3091), .B(n777), .Z(n778) );
  NANDN U1421 ( .A(n3092), .B(n778), .Z(n779) );
  NANDN U1422 ( .A(n3095), .B(n779), .Z(n780) );
  NANDN U1423 ( .A(n3097), .B(n780), .Z(n781) );
  NANDN U1424 ( .A(n3099), .B(n781), .Z(n784) );
  NANDN U1425 ( .A(x[44]), .B(y[44]), .Z(n783) );
  NANDN U1426 ( .A(x[43]), .B(y[43]), .Z(n782) );
  NAND U1427 ( .A(n783), .B(n782), .Z(n3101) );
  ANDN U1428 ( .B(n784), .A(n3101), .Z(n785) );
  OR U1429 ( .A(n3103), .B(n785), .Z(n786) );
  NANDN U1430 ( .A(n3104), .B(n786), .Z(n787) );
  NANDN U1431 ( .A(n3107), .B(n787), .Z(n788) );
  NANDN U1432 ( .A(n3109), .B(n788), .Z(n789) );
  NANDN U1433 ( .A(n3111), .B(n789), .Z(n792) );
  NANDN U1434 ( .A(x[50]), .B(y[50]), .Z(n791) );
  NANDN U1435 ( .A(x[49]), .B(y[49]), .Z(n790) );
  NAND U1436 ( .A(n791), .B(n790), .Z(n3113) );
  ANDN U1437 ( .B(n792), .A(n3113), .Z(n793) );
  OR U1438 ( .A(n3115), .B(n793), .Z(n794) );
  NANDN U1439 ( .A(n3116), .B(n794), .Z(n795) );
  NANDN U1440 ( .A(n3119), .B(n795), .Z(n796) );
  NANDN U1441 ( .A(n3121), .B(n796), .Z(n797) );
  NANDN U1442 ( .A(n3123), .B(n797), .Z(n800) );
  NANDN U1443 ( .A(x[56]), .B(y[56]), .Z(n799) );
  NANDN U1444 ( .A(x[55]), .B(y[55]), .Z(n798) );
  NAND U1445 ( .A(n799), .B(n798), .Z(n3125) );
  ANDN U1446 ( .B(n800), .A(n3125), .Z(n801) );
  OR U1447 ( .A(n3127), .B(n801), .Z(n802) );
  NANDN U1448 ( .A(n3128), .B(n802), .Z(n803) );
  NANDN U1449 ( .A(n3131), .B(n803), .Z(n804) );
  NANDN U1450 ( .A(n3133), .B(n804), .Z(n805) );
  NANDN U1451 ( .A(n3135), .B(n805), .Z(n808) );
  NANDN U1452 ( .A(x[62]), .B(y[62]), .Z(n807) );
  NANDN U1453 ( .A(x[61]), .B(y[61]), .Z(n806) );
  NAND U1454 ( .A(n807), .B(n806), .Z(n3137) );
  ANDN U1455 ( .B(n808), .A(n3137), .Z(n809) );
  OR U1456 ( .A(n3139), .B(n809), .Z(n810) );
  NANDN U1457 ( .A(n3140), .B(n810), .Z(n811) );
  NANDN U1458 ( .A(n3143), .B(n811), .Z(n812) );
  NANDN U1459 ( .A(n3145), .B(n812), .Z(n813) );
  NANDN U1460 ( .A(n3147), .B(n813), .Z(n814) );
  AND U1461 ( .A(n4379), .B(n814), .Z(n815) );
  NANDN U1462 ( .A(x[67]), .B(y[67]), .Z(n3148) );
  NAND U1463 ( .A(n815), .B(n3148), .Z(n816) );
  NANDN U1464 ( .A(n3151), .B(n816), .Z(n817) );
  AND U1465 ( .A(n4383), .B(n817), .Z(n820) );
  NANDN U1466 ( .A(y[70]), .B(x[70]), .Z(n819) );
  NANDN U1467 ( .A(y[71]), .B(x[71]), .Z(n818) );
  AND U1468 ( .A(n819), .B(n818), .Z(n4385) );
  NANDN U1469 ( .A(n820), .B(n4385), .Z(n821) );
  NANDN U1470 ( .A(n4387), .B(n821), .Z(n824) );
  NANDN U1471 ( .A(y[72]), .B(x[72]), .Z(n823) );
  NANDN U1472 ( .A(y[73]), .B(x[73]), .Z(n822) );
  AND U1473 ( .A(n823), .B(n822), .Z(n4389) );
  NAND U1474 ( .A(n824), .B(n4389), .Z(n825) );
  NANDN U1475 ( .A(n4392), .B(n825), .Z(n828) );
  NANDN U1476 ( .A(y[74]), .B(x[74]), .Z(n827) );
  NANDN U1477 ( .A(y[75]), .B(x[75]), .Z(n826) );
  AND U1478 ( .A(n827), .B(n826), .Z(n4393) );
  NAND U1479 ( .A(n828), .B(n4393), .Z(n831) );
  NANDN U1480 ( .A(x[76]), .B(y[76]), .Z(n830) );
  NANDN U1481 ( .A(x[75]), .B(y[75]), .Z(n829) );
  NAND U1482 ( .A(n830), .B(n829), .Z(n4396) );
  ANDN U1483 ( .B(n831), .A(n4396), .Z(n834) );
  NANDN U1484 ( .A(y[76]), .B(x[76]), .Z(n833) );
  NANDN U1485 ( .A(y[77]), .B(x[77]), .Z(n832) );
  AND U1486 ( .A(n833), .B(n832), .Z(n4397) );
  NANDN U1487 ( .A(n834), .B(n4397), .Z(n835) );
  NANDN U1488 ( .A(n4399), .B(n835), .Z(n838) );
  NANDN U1489 ( .A(y[78]), .B(x[78]), .Z(n837) );
  NANDN U1490 ( .A(y[79]), .B(x[79]), .Z(n836) );
  AND U1491 ( .A(n837), .B(n836), .Z(n4401) );
  NAND U1492 ( .A(n838), .B(n4401), .Z(n839) );
  NANDN U1493 ( .A(n4404), .B(n839), .Z(n842) );
  NANDN U1494 ( .A(y[80]), .B(x[80]), .Z(n841) );
  NANDN U1495 ( .A(y[81]), .B(x[81]), .Z(n840) );
  AND U1496 ( .A(n841), .B(n840), .Z(n4405) );
  NAND U1497 ( .A(n842), .B(n4405), .Z(n845) );
  NANDN U1498 ( .A(x[82]), .B(y[82]), .Z(n844) );
  NANDN U1499 ( .A(x[81]), .B(y[81]), .Z(n843) );
  NAND U1500 ( .A(n844), .B(n843), .Z(n4408) );
  ANDN U1501 ( .B(n845), .A(n4408), .Z(n848) );
  NANDN U1502 ( .A(y[82]), .B(x[82]), .Z(n847) );
  NANDN U1503 ( .A(y[83]), .B(x[83]), .Z(n846) );
  AND U1504 ( .A(n847), .B(n846), .Z(n4409) );
  NANDN U1505 ( .A(n848), .B(n4409), .Z(n849) );
  NANDN U1506 ( .A(n4411), .B(n849), .Z(n852) );
  NANDN U1507 ( .A(y[84]), .B(x[84]), .Z(n851) );
  NANDN U1508 ( .A(y[85]), .B(x[85]), .Z(n850) );
  AND U1509 ( .A(n851), .B(n850), .Z(n4413) );
  NAND U1510 ( .A(n852), .B(n4413), .Z(n853) );
  NANDN U1511 ( .A(n3169), .B(n853), .Z(n854) );
  NANDN U1512 ( .A(n3171), .B(n854), .Z(n855) );
  AND U1513 ( .A(n4423), .B(n855), .Z(n858) );
  NANDN U1514 ( .A(y[88]), .B(x[88]), .Z(n857) );
  NANDN U1515 ( .A(y[89]), .B(x[89]), .Z(n856) );
  AND U1516 ( .A(n857), .B(n856), .Z(n4425) );
  NANDN U1517 ( .A(n858), .B(n4425), .Z(n859) );
  NANDN U1518 ( .A(n4427), .B(n859), .Z(n862) );
  NANDN U1519 ( .A(y[90]), .B(x[90]), .Z(n861) );
  NANDN U1520 ( .A(y[91]), .B(x[91]), .Z(n860) );
  AND U1521 ( .A(n861), .B(n860), .Z(n4429) );
  NAND U1522 ( .A(n862), .B(n4429), .Z(n863) );
  NANDN U1523 ( .A(n4432), .B(n863), .Z(n866) );
  NANDN U1524 ( .A(y[92]), .B(x[92]), .Z(n865) );
  NANDN U1525 ( .A(y[93]), .B(x[93]), .Z(n864) );
  AND U1526 ( .A(n865), .B(n864), .Z(n4433) );
  NAND U1527 ( .A(n866), .B(n4433), .Z(n869) );
  NANDN U1528 ( .A(x[94]), .B(y[94]), .Z(n868) );
  NANDN U1529 ( .A(x[93]), .B(y[93]), .Z(n867) );
  NAND U1530 ( .A(n868), .B(n867), .Z(n4436) );
  ANDN U1531 ( .B(n869), .A(n4436), .Z(n872) );
  NANDN U1532 ( .A(y[94]), .B(x[94]), .Z(n871) );
  NANDN U1533 ( .A(y[95]), .B(x[95]), .Z(n870) );
  AND U1534 ( .A(n871), .B(n870), .Z(n4437) );
  NANDN U1535 ( .A(n872), .B(n4437), .Z(n873) );
  NANDN U1536 ( .A(n4439), .B(n873), .Z(n876) );
  NANDN U1537 ( .A(y[96]), .B(x[96]), .Z(n875) );
  NANDN U1538 ( .A(y[97]), .B(x[97]), .Z(n874) );
  AND U1539 ( .A(n875), .B(n874), .Z(n4441) );
  NAND U1540 ( .A(n876), .B(n4441), .Z(n877) );
  NANDN U1541 ( .A(n4444), .B(n877), .Z(n880) );
  NANDN U1542 ( .A(y[99]), .B(x[99]), .Z(n879) );
  NANDN U1543 ( .A(y[98]), .B(x[98]), .Z(n878) );
  AND U1544 ( .A(n879), .B(n878), .Z(n4445) );
  NAND U1545 ( .A(n880), .B(n4445), .Z(n882) );
  ANDN U1546 ( .B(y[99]), .A(x[99]), .Z(n4447) );
  OR U1547 ( .A(n4452), .B(n4447), .Z(n3184) );
  ANDN U1548 ( .B(n882), .A(n3184), .Z(n883) );
  OR U1549 ( .A(n3186), .B(n883), .Z(n884) );
  AND U1550 ( .A(n885), .B(n884), .Z(n887) );
  NANDN U1551 ( .A(y[104]), .B(x[104]), .Z(n886) );
  NANDN U1552 ( .A(y[105]), .B(x[105]), .Z(n2972) );
  AND U1553 ( .A(n886), .B(n2972), .Z(n4459) );
  NANDN U1554 ( .A(n887), .B(n4459), .Z(n888) );
  NANDN U1555 ( .A(n2974), .B(n888), .Z(n891) );
  NANDN U1556 ( .A(y[106]), .B(x[106]), .Z(n890) );
  NANDN U1557 ( .A(y[107]), .B(x[107]), .Z(n889) );
  AND U1558 ( .A(n890), .B(n889), .Z(n4463) );
  NAND U1559 ( .A(n891), .B(n4463), .Z(n892) );
  NANDN U1560 ( .A(n4465), .B(n892), .Z(n895) );
  NANDN U1561 ( .A(y[108]), .B(x[108]), .Z(n894) );
  NANDN U1562 ( .A(y[109]), .B(x[109]), .Z(n893) );
  AND U1563 ( .A(n894), .B(n893), .Z(n4467) );
  NAND U1564 ( .A(n895), .B(n4467), .Z(n898) );
  NANDN U1565 ( .A(x[110]), .B(y[110]), .Z(n897) );
  NANDN U1566 ( .A(x[109]), .B(y[109]), .Z(n896) );
  NAND U1567 ( .A(n897), .B(n896), .Z(n4470) );
  ANDN U1568 ( .B(n898), .A(n4470), .Z(n901) );
  NANDN U1569 ( .A(y[110]), .B(x[110]), .Z(n900) );
  NANDN U1570 ( .A(y[111]), .B(x[111]), .Z(n899) );
  AND U1571 ( .A(n900), .B(n899), .Z(n4471) );
  NANDN U1572 ( .A(n901), .B(n4471), .Z(n902) );
  NANDN U1573 ( .A(n3197), .B(n902), .Z(n903) );
  NANDN U1574 ( .A(n3199), .B(n903), .Z(n904) );
  NANDN U1575 ( .A(x[114]), .B(y[114]), .Z(n4481) );
  NAND U1576 ( .A(n904), .B(n4481), .Z(n907) );
  NANDN U1577 ( .A(y[114]), .B(x[114]), .Z(n906) );
  NANDN U1578 ( .A(y[115]), .B(x[115]), .Z(n905) );
  AND U1579 ( .A(n906), .B(n905), .Z(n4483) );
  NAND U1580 ( .A(n907), .B(n4483), .Z(n910) );
  NANDN U1581 ( .A(x[116]), .B(y[116]), .Z(n909) );
  NANDN U1582 ( .A(x[115]), .B(y[115]), .Z(n908) );
  NAND U1583 ( .A(n909), .B(n908), .Z(n4486) );
  ANDN U1584 ( .B(n910), .A(n4486), .Z(n913) );
  NANDN U1585 ( .A(y[116]), .B(x[116]), .Z(n912) );
  NANDN U1586 ( .A(y[117]), .B(x[117]), .Z(n911) );
  AND U1587 ( .A(n912), .B(n911), .Z(n4487) );
  NANDN U1588 ( .A(n913), .B(n4487), .Z(n914) );
  NANDN U1589 ( .A(n4490), .B(n914), .Z(n917) );
  NANDN U1590 ( .A(y[119]), .B(x[119]), .Z(n916) );
  NANDN U1591 ( .A(y[118]), .B(x[118]), .Z(n915) );
  AND U1592 ( .A(n916), .B(n915), .Z(n4492) );
  NAND U1593 ( .A(n917), .B(n4492), .Z(n918) );
  AND U1594 ( .A(n2968), .B(n918), .Z(n919) );
  NANDN U1595 ( .A(x[119]), .B(y[119]), .Z(n4493) );
  NAND U1596 ( .A(n919), .B(n4493), .Z(n920) );
  NANDN U1597 ( .A(n4496), .B(n920), .Z(n921) );
  NANDN U1598 ( .A(n2970), .B(n921), .Z(n924) );
  NANDN U1599 ( .A(y[122]), .B(x[122]), .Z(n923) );
  NANDN U1600 ( .A(y[123]), .B(x[123]), .Z(n922) );
  AND U1601 ( .A(n923), .B(n922), .Z(n4499) );
  NAND U1602 ( .A(n924), .B(n4499), .Z(n926) );
  ANDN U1603 ( .B(y[123]), .A(x[123]), .Z(n4501) );
  OR U1604 ( .A(n4506), .B(n4501), .Z(n3211) );
  ANDN U1605 ( .B(n926), .A(n3211), .Z(n927) );
  OR U1606 ( .A(n3213), .B(n927), .Z(n928) );
  NANDN U1607 ( .A(x[126]), .B(y[126]), .Z(n4509) );
  NAND U1608 ( .A(n928), .B(n4509), .Z(n931) );
  NANDN U1609 ( .A(y[126]), .B(x[126]), .Z(n930) );
  NANDN U1610 ( .A(y[127]), .B(x[127]), .Z(n929) );
  AND U1611 ( .A(n930), .B(n929), .Z(n4511) );
  NAND U1612 ( .A(n931), .B(n4511), .Z(n932) );
  NANDN U1613 ( .A(n4513), .B(n932), .Z(n933) );
  NANDN U1614 ( .A(n4516), .B(n933), .Z(n934) );
  AND U1615 ( .A(n4517), .B(n934), .Z(n937) );
  NANDN U1616 ( .A(y[130]), .B(x[130]), .Z(n936) );
  NANDN U1617 ( .A(y[131]), .B(x[131]), .Z(n935) );
  AND U1618 ( .A(n936), .B(n935), .Z(n4519) );
  NANDN U1619 ( .A(n937), .B(n4519), .Z(n938) );
  NANDN U1620 ( .A(n4522), .B(n938), .Z(n941) );
  NANDN U1621 ( .A(y[132]), .B(x[132]), .Z(n940) );
  NANDN U1622 ( .A(y[133]), .B(x[133]), .Z(n939) );
  AND U1623 ( .A(n940), .B(n939), .Z(n4523) );
  NAND U1624 ( .A(n941), .B(n4523), .Z(n942) );
  NANDN U1625 ( .A(n3229), .B(n942), .Z(n943) );
  NANDN U1626 ( .A(n3231), .B(n943), .Z(n946) );
  NANDN U1627 ( .A(x[136]), .B(y[136]), .Z(n945) );
  NANDN U1628 ( .A(x[135]), .B(y[135]), .Z(n944) );
  NAND U1629 ( .A(n945), .B(n944), .Z(n4532) );
  ANDN U1630 ( .B(n946), .A(n4532), .Z(n949) );
  NANDN U1631 ( .A(y[136]), .B(x[136]), .Z(n948) );
  NANDN U1632 ( .A(y[137]), .B(x[137]), .Z(n947) );
  AND U1633 ( .A(n948), .B(n947), .Z(n4533) );
  NANDN U1634 ( .A(n949), .B(n4533), .Z(n950) );
  NANDN U1635 ( .A(n4535), .B(n950), .Z(n953) );
  NANDN U1636 ( .A(y[138]), .B(x[138]), .Z(n952) );
  NANDN U1637 ( .A(y[139]), .B(x[139]), .Z(n951) );
  AND U1638 ( .A(n952), .B(n951), .Z(n4537) );
  NAND U1639 ( .A(n953), .B(n4537), .Z(n954) );
  NANDN U1640 ( .A(n4540), .B(n954), .Z(n955) );
  NANDN U1641 ( .A(n4542), .B(n955), .Z(n956) );
  AND U1642 ( .A(n4545), .B(n956), .Z(n957) );
  OR U1643 ( .A(n3246), .B(n957), .Z(n958) );
  NANDN U1644 ( .A(x[144]), .B(y[144]), .Z(n4549) );
  NAND U1645 ( .A(n958), .B(n4549), .Z(n961) );
  NANDN U1646 ( .A(y[145]), .B(x[145]), .Z(n960) );
  NANDN U1647 ( .A(y[144]), .B(x[144]), .Z(n959) );
  AND U1648 ( .A(n960), .B(n959), .Z(n4551) );
  NAND U1649 ( .A(n961), .B(n4551), .Z(n964) );
  NANDN U1650 ( .A(x[145]), .B(y[145]), .Z(n963) );
  NANDN U1651 ( .A(x[146]), .B(y[146]), .Z(n962) );
  AND U1652 ( .A(n963), .B(n962), .Z(n4554) );
  NAND U1653 ( .A(n964), .B(n4554), .Z(n967) );
  NANDN U1654 ( .A(y[147]), .B(x[147]), .Z(n966) );
  NANDN U1655 ( .A(y[146]), .B(x[146]), .Z(n965) );
  AND U1656 ( .A(n966), .B(n965), .Z(n4555) );
  NAND U1657 ( .A(n967), .B(n4555), .Z(n968) );
  AND U1658 ( .A(n4557), .B(n968), .Z(n971) );
  NANDN U1659 ( .A(y[149]), .B(x[149]), .Z(n970) );
  NANDN U1660 ( .A(y[148]), .B(x[148]), .Z(n969) );
  AND U1661 ( .A(n970), .B(n969), .Z(n4559) );
  NANDN U1662 ( .A(n971), .B(n4559), .Z(n974) );
  NANDN U1663 ( .A(x[149]), .B(y[149]), .Z(n973) );
  NANDN U1664 ( .A(x[150]), .B(y[150]), .Z(n972) );
  AND U1665 ( .A(n973), .B(n972), .Z(n4561) );
  NAND U1666 ( .A(n974), .B(n4561), .Z(n977) );
  NANDN U1667 ( .A(y[151]), .B(x[151]), .Z(n976) );
  NANDN U1668 ( .A(y[150]), .B(x[150]), .Z(n975) );
  AND U1669 ( .A(n976), .B(n975), .Z(n4563) );
  NAND U1670 ( .A(n977), .B(n4563), .Z(n978) );
  NANDN U1671 ( .A(n3256), .B(n978), .Z(n979) );
  NANDN U1672 ( .A(n3257), .B(n979), .Z(n980) );
  AND U1673 ( .A(n4571), .B(n980), .Z(n981) );
  OR U1674 ( .A(n4574), .B(n981), .Z(n984) );
  NANDN U1675 ( .A(x[155]), .B(y[155]), .Z(n983) );
  NANDN U1676 ( .A(x[156]), .B(y[156]), .Z(n982) );
  AND U1677 ( .A(n983), .B(n982), .Z(n4576) );
  NAND U1678 ( .A(n984), .B(n4576), .Z(n987) );
  NANDN U1679 ( .A(y[156]), .B(x[156]), .Z(n986) );
  NANDN U1680 ( .A(y[157]), .B(x[157]), .Z(n985) );
  AND U1681 ( .A(n986), .B(n985), .Z(n4577) );
  NAND U1682 ( .A(n987), .B(n4577), .Z(n988) );
  AND U1683 ( .A(n2964), .B(n988), .Z(n989) );
  NANDN U1684 ( .A(x[157]), .B(y[157]), .Z(n4579) );
  NAND U1685 ( .A(n989), .B(n4579), .Z(n991) );
  NANDN U1686 ( .A(y[158]), .B(x[158]), .Z(n990) );
  NANDN U1687 ( .A(y[159]), .B(x[159]), .Z(n2963) );
  AND U1688 ( .A(n990), .B(n2963), .Z(n4581) );
  NAND U1689 ( .A(n991), .B(n4581), .Z(n992) );
  NANDN U1690 ( .A(n2966), .B(n992), .Z(n995) );
  NANDN U1691 ( .A(y[161]), .B(x[161]), .Z(n994) );
  NANDN U1692 ( .A(y[160]), .B(x[160]), .Z(n993) );
  AND U1693 ( .A(n994), .B(n993), .Z(n4585) );
  NAND U1694 ( .A(n995), .B(n4585), .Z(n997) );
  NANDN U1695 ( .A(x[161]), .B(y[161]), .Z(n3267) );
  NANDN U1696 ( .A(n3272), .B(n3267), .Z(n4587) );
  ANDN U1697 ( .B(n997), .A(n4587), .Z(n998) );
  OR U1698 ( .A(n4590), .B(n998), .Z(n999) );
  NANDN U1699 ( .A(x[164]), .B(y[164]), .Z(n4591) );
  NAND U1700 ( .A(n999), .B(n4591), .Z(n1002) );
  NANDN U1701 ( .A(y[164]), .B(x[164]), .Z(n1001) );
  NANDN U1702 ( .A(y[165]), .B(x[165]), .Z(n1000) );
  AND U1703 ( .A(n1001), .B(n1000), .Z(n4593) );
  NAND U1704 ( .A(n1002), .B(n4593), .Z(n1003) );
  NANDN U1705 ( .A(n3278), .B(n1003), .Z(n1006) );
  IV U1706 ( .A(x[167]), .Z(n4604) );
  OR U1707 ( .A(y[167]), .B(n4604), .Z(n1005) );
  IV U1708 ( .A(x[166]), .Z(n4372) );
  OR U1709 ( .A(y[166]), .B(n4372), .Z(n1004) );
  AND U1710 ( .A(n1005), .B(n1004), .Z(n3279) );
  NAND U1711 ( .A(n1006), .B(n3279), .Z(n1008) );
  ANDN U1712 ( .B(y[168]), .A(x[168]), .Z(n4601) );
  NANDN U1713 ( .A(x[167]), .B(y[167]), .Z(n1007) );
  NANDN U1714 ( .A(n4601), .B(n1007), .Z(n3282) );
  ANDN U1715 ( .B(n1008), .A(n3282), .Z(n1011) );
  NANDN U1716 ( .A(y[169]), .B(x[169]), .Z(n1010) );
  NANDN U1717 ( .A(y[168]), .B(x[168]), .Z(n1009) );
  AND U1718 ( .A(n1010), .B(n1009), .Z(n4608) );
  NANDN U1719 ( .A(n1011), .B(n4608), .Z(n1014) );
  NANDN U1720 ( .A(x[169]), .B(y[169]), .Z(n1013) );
  NANDN U1721 ( .A(x[170]), .B(y[170]), .Z(n1012) );
  AND U1722 ( .A(n1013), .B(n1012), .Z(n4610) );
  NAND U1723 ( .A(n1014), .B(n4610), .Z(n1017) );
  NANDN U1724 ( .A(y[171]), .B(x[171]), .Z(n1016) );
  NANDN U1725 ( .A(y[170]), .B(x[170]), .Z(n1015) );
  AND U1726 ( .A(n1016), .B(n1015), .Z(n4613) );
  NAND U1727 ( .A(n1017), .B(n4613), .Z(n1020) );
  NANDN U1728 ( .A(x[171]), .B(y[171]), .Z(n1019) );
  NANDN U1729 ( .A(x[172]), .B(y[172]), .Z(n1018) );
  AND U1730 ( .A(n1019), .B(n1018), .Z(n4614) );
  NAND U1731 ( .A(n1020), .B(n4614), .Z(n1023) );
  NANDN U1732 ( .A(y[172]), .B(x[172]), .Z(n1022) );
  NANDN U1733 ( .A(y[173]), .B(x[173]), .Z(n1021) );
  AND U1734 ( .A(n1022), .B(n1021), .Z(n4616) );
  NAND U1735 ( .A(n1023), .B(n4616), .Z(n1024) );
  AND U1736 ( .A(n2960), .B(n1024), .Z(n1025) );
  NANDN U1737 ( .A(x[173]), .B(y[173]), .Z(n4618) );
  NAND U1738 ( .A(n1025), .B(n4618), .Z(n1026) );
  NANDN U1739 ( .A(n4621), .B(n1026), .Z(n1029) );
  NANDN U1740 ( .A(x[176]), .B(y[176]), .Z(n1028) );
  NANDN U1741 ( .A(x[175]), .B(y[175]), .Z(n1027) );
  NAND U1742 ( .A(n1028), .B(n1027), .Z(n2962) );
  ANDN U1743 ( .B(n1029), .A(n2962), .Z(n1032) );
  NANDN U1744 ( .A(y[177]), .B(x[177]), .Z(n1031) );
  NANDN U1745 ( .A(y[176]), .B(x[176]), .Z(n1030) );
  AND U1746 ( .A(n1031), .B(n1030), .Z(n4625) );
  NANDN U1747 ( .A(n1032), .B(n4625), .Z(n1033) );
  NANDN U1748 ( .A(n4627), .B(n1033), .Z(n1034) );
  NANDN U1749 ( .A(n4629), .B(n1034), .Z(n1035) );
  NANDN U1750 ( .A(x[180]), .B(y[180]), .Z(n4630) );
  NAND U1751 ( .A(n1035), .B(n4630), .Z(n1038) );
  NANDN U1752 ( .A(y[181]), .B(x[181]), .Z(n1037) );
  NANDN U1753 ( .A(y[180]), .B(x[180]), .Z(n1036) );
  AND U1754 ( .A(n1037), .B(n1036), .Z(n4632) );
  NAND U1755 ( .A(n1038), .B(n4632), .Z(n1039) );
  AND U1756 ( .A(n4634), .B(n1039), .Z(n1042) );
  NANDN U1757 ( .A(y[183]), .B(x[183]), .Z(n1041) );
  NANDN U1758 ( .A(y[182]), .B(x[182]), .Z(n1040) );
  AND U1759 ( .A(n1041), .B(n1040), .Z(n4637) );
  NANDN U1760 ( .A(n1042), .B(n4637), .Z(n1045) );
  NANDN U1761 ( .A(x[183]), .B(y[183]), .Z(n1044) );
  NANDN U1762 ( .A(x[184]), .B(y[184]), .Z(n1043) );
  AND U1763 ( .A(n1044), .B(n1043), .Z(n4638) );
  NAND U1764 ( .A(n1045), .B(n4638), .Z(n1048) );
  NANDN U1765 ( .A(y[185]), .B(x[185]), .Z(n1047) );
  NANDN U1766 ( .A(y[184]), .B(x[184]), .Z(n1046) );
  AND U1767 ( .A(n1047), .B(n1046), .Z(n4640) );
  NAND U1768 ( .A(n1048), .B(n4640), .Z(n1051) );
  NANDN U1769 ( .A(x[185]), .B(y[185]), .Z(n1050) );
  NANDN U1770 ( .A(x[186]), .B(y[186]), .Z(n1049) );
  AND U1771 ( .A(n1050), .B(n1049), .Z(n4642) );
  NAND U1772 ( .A(n1051), .B(n4642), .Z(n1054) );
  NANDN U1773 ( .A(y[187]), .B(x[187]), .Z(n1053) );
  NANDN U1774 ( .A(y[186]), .B(x[186]), .Z(n1052) );
  AND U1775 ( .A(n1053), .B(n1052), .Z(n4644) );
  NAND U1776 ( .A(n1054), .B(n4644), .Z(n1055) );
  AND U1777 ( .A(n4646), .B(n1055), .Z(n1058) );
  NANDN U1778 ( .A(y[189]), .B(x[189]), .Z(n1057) );
  NANDN U1779 ( .A(y[188]), .B(x[188]), .Z(n1056) );
  AND U1780 ( .A(n1057), .B(n1056), .Z(n4649) );
  NANDN U1781 ( .A(n1058), .B(n4649), .Z(n1061) );
  NANDN U1782 ( .A(x[189]), .B(y[189]), .Z(n1060) );
  NANDN U1783 ( .A(x[190]), .B(y[190]), .Z(n1059) );
  AND U1784 ( .A(n1060), .B(n1059), .Z(n4650) );
  NAND U1785 ( .A(n1061), .B(n4650), .Z(n1064) );
  NANDN U1786 ( .A(y[191]), .B(x[191]), .Z(n1063) );
  NANDN U1787 ( .A(y[190]), .B(x[190]), .Z(n1062) );
  AND U1788 ( .A(n1063), .B(n1062), .Z(n4652) );
  NAND U1789 ( .A(n1064), .B(n4652), .Z(n1067) );
  NANDN U1790 ( .A(x[191]), .B(y[191]), .Z(n1066) );
  NANDN U1791 ( .A(x[192]), .B(y[192]), .Z(n1065) );
  AND U1792 ( .A(n1066), .B(n1065), .Z(n4654) );
  NAND U1793 ( .A(n1067), .B(n4654), .Z(n1070) );
  NANDN U1794 ( .A(y[193]), .B(x[193]), .Z(n1069) );
  NANDN U1795 ( .A(y[192]), .B(x[192]), .Z(n1068) );
  AND U1796 ( .A(n1069), .B(n1068), .Z(n4656) );
  NAND U1797 ( .A(n1070), .B(n4656), .Z(n1071) );
  AND U1798 ( .A(n4658), .B(n1071), .Z(n1074) );
  NANDN U1799 ( .A(y[195]), .B(x[195]), .Z(n1073) );
  NANDN U1800 ( .A(y[194]), .B(x[194]), .Z(n1072) );
  AND U1801 ( .A(n1073), .B(n1072), .Z(n4661) );
  NANDN U1802 ( .A(n1074), .B(n4661), .Z(n1077) );
  NANDN U1803 ( .A(x[195]), .B(y[195]), .Z(n1076) );
  NANDN U1804 ( .A(x[196]), .B(y[196]), .Z(n1075) );
  AND U1805 ( .A(n1076), .B(n1075), .Z(n4662) );
  NAND U1806 ( .A(n1077), .B(n4662), .Z(n1080) );
  NANDN U1807 ( .A(y[197]), .B(x[197]), .Z(n1079) );
  NANDN U1808 ( .A(y[196]), .B(x[196]), .Z(n1078) );
  AND U1809 ( .A(n1079), .B(n1078), .Z(n4664) );
  NAND U1810 ( .A(n1080), .B(n4664), .Z(n1083) );
  NANDN U1811 ( .A(x[197]), .B(y[197]), .Z(n1082) );
  NANDN U1812 ( .A(x[198]), .B(y[198]), .Z(n1081) );
  AND U1813 ( .A(n1082), .B(n1081), .Z(n4666) );
  NAND U1814 ( .A(n1083), .B(n4666), .Z(n1086) );
  NANDN U1815 ( .A(y[199]), .B(x[199]), .Z(n1085) );
  NANDN U1816 ( .A(y[198]), .B(x[198]), .Z(n1084) );
  AND U1817 ( .A(n1085), .B(n1084), .Z(n4668) );
  NAND U1818 ( .A(n1086), .B(n4668), .Z(n1087) );
  ANDN U1819 ( .B(y[201]), .A(x[201]), .Z(n1089) );
  NANDN U1820 ( .A(x[199]), .B(y[199]), .Z(n3320) );
  NANDN U1821 ( .A(n3325), .B(n3320), .Z(n4671) );
  ANDN U1822 ( .B(n1087), .A(n4671), .Z(n1090) );
  NANDN U1823 ( .A(y[200]), .B(x[200]), .Z(n3323) );
  ANDN U1824 ( .B(x[201]), .A(y[201]), .Z(n3326) );
  ANDN U1825 ( .B(n3323), .A(n3326), .Z(n1088) );
  OR U1826 ( .A(n1089), .B(n1088), .Z(n4673) );
  NANDN U1827 ( .A(n1090), .B(n4673), .Z(n1091) );
  NANDN U1828 ( .A(x[202]), .B(y[202]), .Z(n4674) );
  NAND U1829 ( .A(n1091), .B(n4674), .Z(n1094) );
  NANDN U1830 ( .A(y[203]), .B(x[203]), .Z(n1093) );
  NANDN U1831 ( .A(y[202]), .B(x[202]), .Z(n1092) );
  AND U1832 ( .A(n1093), .B(n1092), .Z(n4676) );
  NAND U1833 ( .A(n1094), .B(n4676), .Z(n1097) );
  NANDN U1834 ( .A(x[203]), .B(y[203]), .Z(n1096) );
  NANDN U1835 ( .A(x[204]), .B(y[204]), .Z(n1095) );
  AND U1836 ( .A(n1096), .B(n1095), .Z(n4678) );
  NAND U1837 ( .A(n1097), .B(n4678), .Z(n1100) );
  NANDN U1838 ( .A(y[205]), .B(x[205]), .Z(n1099) );
  NANDN U1839 ( .A(y[204]), .B(x[204]), .Z(n1098) );
  AND U1840 ( .A(n1099), .B(n1098), .Z(n4680) );
  NAND U1841 ( .A(n1100), .B(n4680), .Z(n1101) );
  AND U1842 ( .A(n4682), .B(n1101), .Z(n1104) );
  NANDN U1843 ( .A(y[207]), .B(x[207]), .Z(n1103) );
  NANDN U1844 ( .A(y[206]), .B(x[206]), .Z(n1102) );
  AND U1845 ( .A(n1103), .B(n1102), .Z(n4685) );
  NANDN U1846 ( .A(n1104), .B(n4685), .Z(n1107) );
  NANDN U1847 ( .A(x[207]), .B(y[207]), .Z(n1106) );
  NANDN U1848 ( .A(x[208]), .B(y[208]), .Z(n1105) );
  AND U1849 ( .A(n1106), .B(n1105), .Z(n4686) );
  NAND U1850 ( .A(n1107), .B(n4686), .Z(n1110) );
  NANDN U1851 ( .A(y[209]), .B(x[209]), .Z(n1109) );
  NANDN U1852 ( .A(y[208]), .B(x[208]), .Z(n1108) );
  AND U1853 ( .A(n1109), .B(n1108), .Z(n4688) );
  NAND U1854 ( .A(n1110), .B(n4688), .Z(n1113) );
  NANDN U1855 ( .A(x[209]), .B(y[209]), .Z(n1112) );
  NANDN U1856 ( .A(x[210]), .B(y[210]), .Z(n1111) );
  AND U1857 ( .A(n1112), .B(n1111), .Z(n4690) );
  NAND U1858 ( .A(n1113), .B(n4690), .Z(n1116) );
  NANDN U1859 ( .A(y[211]), .B(x[211]), .Z(n1115) );
  NANDN U1860 ( .A(y[210]), .B(x[210]), .Z(n1114) );
  AND U1861 ( .A(n1115), .B(n1114), .Z(n4692) );
  NAND U1862 ( .A(n1116), .B(n4692), .Z(n1117) );
  AND U1863 ( .A(n4694), .B(n1117), .Z(n1120) );
  NANDN U1864 ( .A(y[213]), .B(x[213]), .Z(n1119) );
  NANDN U1865 ( .A(y[212]), .B(x[212]), .Z(n1118) );
  AND U1866 ( .A(n1119), .B(n1118), .Z(n4697) );
  NANDN U1867 ( .A(n1120), .B(n4697), .Z(n1123) );
  NANDN U1868 ( .A(x[213]), .B(y[213]), .Z(n1122) );
  NANDN U1869 ( .A(x[214]), .B(y[214]), .Z(n1121) );
  AND U1870 ( .A(n1122), .B(n1121), .Z(n4698) );
  NAND U1871 ( .A(n1123), .B(n4698), .Z(n1126) );
  NANDN U1872 ( .A(y[214]), .B(x[214]), .Z(n1125) );
  NANDN U1873 ( .A(y[215]), .B(x[215]), .Z(n1124) );
  AND U1874 ( .A(n1125), .B(n1124), .Z(n4700) );
  NAND U1875 ( .A(n1126), .B(n4700), .Z(n1127) );
  AND U1876 ( .A(n2956), .B(n1127), .Z(n1128) );
  NANDN U1877 ( .A(x[215]), .B(y[215]), .Z(n4702) );
  NAND U1878 ( .A(n1128), .B(n4702), .Z(n1129) );
  NANDN U1879 ( .A(n4705), .B(n1129), .Z(n1130) );
  NANDN U1880 ( .A(n2958), .B(n1130), .Z(n1131) );
  NANDN U1881 ( .A(n4708), .B(n1131), .Z(n1134) );
  NANDN U1882 ( .A(x[219]), .B(y[219]), .Z(n1133) );
  NANDN U1883 ( .A(x[220]), .B(y[220]), .Z(n1132) );
  AND U1884 ( .A(n1133), .B(n1132), .Z(n4710) );
  NAND U1885 ( .A(n1134), .B(n4710), .Z(n1135) );
  NANDN U1886 ( .A(n4713), .B(n1135), .Z(n1138) );
  NANDN U1887 ( .A(x[221]), .B(y[221]), .Z(n1137) );
  NANDN U1888 ( .A(x[222]), .B(y[222]), .Z(n1136) );
  AND U1889 ( .A(n1137), .B(n1136), .Z(n4714) );
  NAND U1890 ( .A(n1138), .B(n4714), .Z(n1141) );
  NANDN U1891 ( .A(y[223]), .B(x[223]), .Z(n1140) );
  NANDN U1892 ( .A(y[222]), .B(x[222]), .Z(n1139) );
  NAND U1893 ( .A(n1140), .B(n1139), .Z(n4717) );
  ANDN U1894 ( .B(n1141), .A(n4717), .Z(n1144) );
  NANDN U1895 ( .A(x[223]), .B(y[223]), .Z(n1143) );
  NANDN U1896 ( .A(x[224]), .B(y[224]), .Z(n1142) );
  AND U1897 ( .A(n1143), .B(n1142), .Z(n4718) );
  NANDN U1898 ( .A(n1144), .B(n4718), .Z(n1145) );
  NANDN U1899 ( .A(n4720), .B(n1145), .Z(n1148) );
  NANDN U1900 ( .A(x[225]), .B(y[225]), .Z(n1147) );
  NANDN U1901 ( .A(x[226]), .B(y[226]), .Z(n1146) );
  AND U1902 ( .A(n1147), .B(n1146), .Z(n4722) );
  NAND U1903 ( .A(n1148), .B(n4722), .Z(n1149) );
  NANDN U1904 ( .A(n4724), .B(n1149), .Z(n1152) );
  NANDN U1905 ( .A(x[227]), .B(y[227]), .Z(n1151) );
  NANDN U1906 ( .A(x[228]), .B(y[228]), .Z(n1150) );
  AND U1907 ( .A(n1151), .B(n1150), .Z(n4726) );
  NAND U1908 ( .A(n1152), .B(n4726), .Z(n1155) );
  NANDN U1909 ( .A(y[229]), .B(x[229]), .Z(n1154) );
  NANDN U1910 ( .A(y[228]), .B(x[228]), .Z(n1153) );
  NAND U1911 ( .A(n1154), .B(n1153), .Z(n4729) );
  ANDN U1912 ( .B(n1155), .A(n4729), .Z(n1156) );
  OR U1913 ( .A(n3357), .B(n1156), .Z(n1157) );
  NANDN U1914 ( .A(n3358), .B(n1157), .Z(n1158) );
  NANDN U1915 ( .A(x[232]), .B(y[232]), .Z(n4738) );
  NAND U1916 ( .A(n1158), .B(n4738), .Z(n1159) );
  NANDN U1917 ( .A(n4741), .B(n1159), .Z(n1162) );
  NANDN U1918 ( .A(x[233]), .B(y[233]), .Z(n1161) );
  NANDN U1919 ( .A(x[234]), .B(y[234]), .Z(n1160) );
  AND U1920 ( .A(n1161), .B(n1160), .Z(n4742) );
  NAND U1921 ( .A(n1162), .B(n4742), .Z(n1165) );
  NANDN U1922 ( .A(y[235]), .B(x[235]), .Z(n1164) );
  NANDN U1923 ( .A(y[234]), .B(x[234]), .Z(n1163) );
  NAND U1924 ( .A(n1164), .B(n1163), .Z(n4745) );
  ANDN U1925 ( .B(n1165), .A(n4745), .Z(n1168) );
  NANDN U1926 ( .A(x[235]), .B(y[235]), .Z(n1167) );
  NANDN U1927 ( .A(x[236]), .B(y[236]), .Z(n1166) );
  AND U1928 ( .A(n1167), .B(n1166), .Z(n4746) );
  NANDN U1929 ( .A(n1168), .B(n4746), .Z(n1169) );
  NANDN U1930 ( .A(n4748), .B(n1169), .Z(n1172) );
  NANDN U1931 ( .A(x[237]), .B(y[237]), .Z(n1171) );
  NANDN U1932 ( .A(x[238]), .B(y[238]), .Z(n1170) );
  AND U1933 ( .A(n1171), .B(n1170), .Z(n4750) );
  NAND U1934 ( .A(n1172), .B(n4750), .Z(n1173) );
  NANDN U1935 ( .A(n4753), .B(n1173), .Z(n1176) );
  NANDN U1936 ( .A(x[239]), .B(y[239]), .Z(n1175) );
  NANDN U1937 ( .A(x[240]), .B(y[240]), .Z(n1174) );
  AND U1938 ( .A(n1175), .B(n1174), .Z(n4754) );
  NAND U1939 ( .A(n1176), .B(n4754), .Z(n1179) );
  NANDN U1940 ( .A(y[241]), .B(x[241]), .Z(n1178) );
  NANDN U1941 ( .A(y[240]), .B(x[240]), .Z(n1177) );
  NAND U1942 ( .A(n1178), .B(n1177), .Z(n4757) );
  ANDN U1943 ( .B(n1179), .A(n4757), .Z(n1180) );
  OR U1944 ( .A(n4759), .B(n1180), .Z(n1181) );
  NANDN U1945 ( .A(n4760), .B(n1181), .Z(n1182) );
  NANDN U1946 ( .A(x[244]), .B(y[244]), .Z(n4762) );
  NAND U1947 ( .A(n1182), .B(n4762), .Z(n1183) );
  NANDN U1948 ( .A(n4765), .B(n1183), .Z(n1186) );
  NANDN U1949 ( .A(x[245]), .B(y[245]), .Z(n1185) );
  NANDN U1950 ( .A(x[246]), .B(y[246]), .Z(n1184) );
  AND U1951 ( .A(n1185), .B(n1184), .Z(n4766) );
  NAND U1952 ( .A(n1186), .B(n4766), .Z(n1189) );
  NANDN U1953 ( .A(y[247]), .B(x[247]), .Z(n1188) );
  NANDN U1954 ( .A(y[246]), .B(x[246]), .Z(n1187) );
  NAND U1955 ( .A(n1188), .B(n1187), .Z(n4769) );
  ANDN U1956 ( .B(n1189), .A(n4769), .Z(n1192) );
  NANDN U1957 ( .A(x[247]), .B(y[247]), .Z(n1191) );
  NANDN U1958 ( .A(x[248]), .B(y[248]), .Z(n1190) );
  AND U1959 ( .A(n1191), .B(n1190), .Z(n4770) );
  NANDN U1960 ( .A(n1192), .B(n4770), .Z(n1193) );
  NANDN U1961 ( .A(n4772), .B(n1193), .Z(n1198) );
  NANDN U1962 ( .A(x[250]), .B(y[250]), .Z(n1195) );
  NANDN U1963 ( .A(x[249]), .B(y[249]), .Z(n1194) );
  AND U1964 ( .A(n1195), .B(n1194), .Z(n1197) );
  AND U1965 ( .A(n1197), .B(n1196), .Z(n4774) );
  NAND U1966 ( .A(n1198), .B(n4774), .Z(n1199) );
  NANDN U1967 ( .A(n4777), .B(n1199), .Z(n1200) );
  NANDN U1968 ( .A(x[252]), .B(y[252]), .Z(n4778) );
  NAND U1969 ( .A(n1200), .B(n4778), .Z(n1203) );
  NANDN U1970 ( .A(y[253]), .B(x[253]), .Z(n1202) );
  NANDN U1971 ( .A(y[252]), .B(x[252]), .Z(n1201) );
  NAND U1972 ( .A(n1202), .B(n1201), .Z(n4781) );
  ANDN U1973 ( .B(n1203), .A(n4781), .Z(n1206) );
  NANDN U1974 ( .A(x[253]), .B(y[253]), .Z(n1205) );
  NANDN U1975 ( .A(x[254]), .B(y[254]), .Z(n1204) );
  AND U1976 ( .A(n1205), .B(n1204), .Z(n4782) );
  NANDN U1977 ( .A(n1206), .B(n4782), .Z(n1207) );
  NANDN U1978 ( .A(n4784), .B(n1207), .Z(n1210) );
  NANDN U1979 ( .A(x[255]), .B(y[255]), .Z(n1209) );
  NANDN U1980 ( .A(x[256]), .B(y[256]), .Z(n1208) );
  AND U1981 ( .A(n1209), .B(n1208), .Z(n4786) );
  NAND U1982 ( .A(n1210), .B(n4786), .Z(n1211) );
  NANDN U1983 ( .A(n4789), .B(n1211), .Z(n1214) );
  NANDN U1984 ( .A(x[257]), .B(y[257]), .Z(n1213) );
  NANDN U1985 ( .A(x[258]), .B(y[258]), .Z(n1212) );
  AND U1986 ( .A(n1213), .B(n1212), .Z(n4790) );
  NAND U1987 ( .A(n1214), .B(n4790), .Z(n1217) );
  NANDN U1988 ( .A(y[259]), .B(x[259]), .Z(n1216) );
  NANDN U1989 ( .A(y[258]), .B(x[258]), .Z(n1215) );
  NAND U1990 ( .A(n1216), .B(n1215), .Z(n4793) );
  ANDN U1991 ( .B(n1217), .A(n4793), .Z(n1220) );
  NANDN U1992 ( .A(x[259]), .B(y[259]), .Z(n1219) );
  NANDN U1993 ( .A(x[260]), .B(y[260]), .Z(n1218) );
  AND U1994 ( .A(n1219), .B(n1218), .Z(n4794) );
  NANDN U1995 ( .A(n1220), .B(n4794), .Z(n1221) );
  NANDN U1996 ( .A(n4796), .B(n1221), .Z(n1224) );
  NANDN U1997 ( .A(x[261]), .B(y[261]), .Z(n1223) );
  NANDN U1998 ( .A(x[262]), .B(y[262]), .Z(n1222) );
  AND U1999 ( .A(n1223), .B(n1222), .Z(n4798) );
  NAND U2000 ( .A(n1224), .B(n4798), .Z(n1225) );
  NANDN U2001 ( .A(n4800), .B(n1225), .Z(n1228) );
  NANDN U2002 ( .A(x[263]), .B(y[263]), .Z(n1227) );
  NANDN U2003 ( .A(x[264]), .B(y[264]), .Z(n1226) );
  AND U2004 ( .A(n1227), .B(n1226), .Z(n4802) );
  NAND U2005 ( .A(n1228), .B(n4802), .Z(n1231) );
  NANDN U2006 ( .A(y[265]), .B(x[265]), .Z(n1230) );
  NANDN U2007 ( .A(y[264]), .B(x[264]), .Z(n1229) );
  NAND U2008 ( .A(n1230), .B(n1229), .Z(n4805) );
  ANDN U2009 ( .B(n1231), .A(n4805), .Z(n1232) );
  OR U2010 ( .A(n3401), .B(n1232), .Z(n1233) );
  NANDN U2011 ( .A(n3402), .B(n1233), .Z(n1234) );
  NANDN U2012 ( .A(x[268]), .B(y[268]), .Z(n4814) );
  NAND U2013 ( .A(n1234), .B(n4814), .Z(n1235) );
  NANDN U2014 ( .A(n4817), .B(n1235), .Z(n1238) );
  NANDN U2015 ( .A(x[269]), .B(y[269]), .Z(n1237) );
  NANDN U2016 ( .A(x[270]), .B(y[270]), .Z(n1236) );
  AND U2017 ( .A(n1237), .B(n1236), .Z(n4818) );
  NAND U2018 ( .A(n1238), .B(n4818), .Z(n1241) );
  NANDN U2019 ( .A(y[271]), .B(x[271]), .Z(n1240) );
  NANDN U2020 ( .A(y[270]), .B(x[270]), .Z(n1239) );
  NAND U2021 ( .A(n1240), .B(n1239), .Z(n4821) );
  ANDN U2022 ( .B(n1241), .A(n4821), .Z(n1244) );
  NANDN U2023 ( .A(x[271]), .B(y[271]), .Z(n1243) );
  NANDN U2024 ( .A(x[272]), .B(y[272]), .Z(n1242) );
  AND U2025 ( .A(n1243), .B(n1242), .Z(n4822) );
  NANDN U2026 ( .A(n1244), .B(n4822), .Z(n1245) );
  NANDN U2027 ( .A(n4825), .B(n1245), .Z(n1246) );
  NANDN U2028 ( .A(n3411), .B(n1246), .Z(n1247) );
  NANDN U2029 ( .A(n3413), .B(n1247), .Z(n1248) );
  NANDN U2030 ( .A(x[276]), .B(y[276]), .Z(n4831) );
  NAND U2031 ( .A(n1248), .B(n4831), .Z(n1251) );
  NANDN U2032 ( .A(y[277]), .B(x[277]), .Z(n1250) );
  NANDN U2033 ( .A(y[276]), .B(x[276]), .Z(n1249) );
  NAND U2034 ( .A(n1250), .B(n1249), .Z(n4835) );
  ANDN U2035 ( .B(n1251), .A(n4835), .Z(n1254) );
  NANDN U2036 ( .A(x[277]), .B(y[277]), .Z(n1253) );
  NANDN U2037 ( .A(x[278]), .B(y[278]), .Z(n1252) );
  AND U2038 ( .A(n1253), .B(n1252), .Z(n4836) );
  NANDN U2039 ( .A(n1254), .B(n4836), .Z(n1255) );
  NANDN U2040 ( .A(n4839), .B(n1255), .Z(n1258) );
  NANDN U2041 ( .A(x[279]), .B(y[279]), .Z(n1257) );
  NANDN U2042 ( .A(x[280]), .B(y[280]), .Z(n1256) );
  AND U2043 ( .A(n1257), .B(n1256), .Z(n4840) );
  NAND U2044 ( .A(n1258), .B(n4840), .Z(n1259) );
  NANDN U2045 ( .A(n4841), .B(n1259), .Z(n1262) );
  NANDN U2046 ( .A(x[281]), .B(y[281]), .Z(n1261) );
  NANDN U2047 ( .A(x[282]), .B(y[282]), .Z(n1260) );
  AND U2048 ( .A(n1261), .B(n1260), .Z(n4842) );
  NAND U2049 ( .A(n1262), .B(n4842), .Z(n1265) );
  NANDN U2050 ( .A(y[283]), .B(x[283]), .Z(n1264) );
  NANDN U2051 ( .A(y[282]), .B(x[282]), .Z(n1263) );
  NAND U2052 ( .A(n1264), .B(n1263), .Z(n4843) );
  ANDN U2053 ( .B(n1265), .A(n4843), .Z(n1268) );
  NANDN U2054 ( .A(x[283]), .B(y[283]), .Z(n1267) );
  NANDN U2055 ( .A(x[284]), .B(y[284]), .Z(n1266) );
  AND U2056 ( .A(n1267), .B(n1266), .Z(n4844) );
  NANDN U2057 ( .A(n1268), .B(n4844), .Z(n1269) );
  NANDN U2058 ( .A(n4845), .B(n1269), .Z(n1270) );
  NANDN U2059 ( .A(n3425), .B(n1270), .Z(n1271) );
  NANDN U2060 ( .A(n3427), .B(n1271), .Z(n1272) );
  NANDN U2061 ( .A(x[288]), .B(y[288]), .Z(n4849) );
  NAND U2062 ( .A(n1272), .B(n4849), .Z(n1275) );
  NANDN U2063 ( .A(y[289]), .B(x[289]), .Z(n1274) );
  NANDN U2064 ( .A(y[288]), .B(x[288]), .Z(n1273) );
  NAND U2065 ( .A(n1274), .B(n1273), .Z(n4850) );
  ANDN U2066 ( .B(n1275), .A(n4850), .Z(n1278) );
  NANDN U2067 ( .A(x[289]), .B(y[289]), .Z(n1277) );
  NANDN U2068 ( .A(x[290]), .B(y[290]), .Z(n1276) );
  AND U2069 ( .A(n1277), .B(n1276), .Z(n4851) );
  NANDN U2070 ( .A(n1278), .B(n4851), .Z(n1279) );
  NANDN U2071 ( .A(n4852), .B(n1279), .Z(n1282) );
  NANDN U2072 ( .A(x[291]), .B(y[291]), .Z(n1281) );
  NANDN U2073 ( .A(x[292]), .B(y[292]), .Z(n1280) );
  AND U2074 ( .A(n1281), .B(n1280), .Z(n4853) );
  NAND U2075 ( .A(n1282), .B(n4853), .Z(n1283) );
  NANDN U2076 ( .A(n4854), .B(n1283), .Z(n1284) );
  NANDN U2077 ( .A(x[293]), .B(y[293]), .Z(n4369) );
  NAND U2078 ( .A(n1284), .B(n3434), .Z(n1286) );
  NANDN U2079 ( .A(y[295]), .B(x[295]), .Z(n4862) );
  NANDN U2080 ( .A(y[294]), .B(x[294]), .Z(n1285) );
  NAND U2081 ( .A(n4862), .B(n1285), .Z(n3437) );
  ANDN U2082 ( .B(n1286), .A(n3437), .Z(n1287) );
  OR U2083 ( .A(n3439), .B(n1287), .Z(n1288) );
  NANDN U2084 ( .A(n4866), .B(n1288), .Z(n1291) );
  NANDN U2085 ( .A(x[297]), .B(y[297]), .Z(n1290) );
  NANDN U2086 ( .A(x[298]), .B(y[298]), .Z(n1289) );
  AND U2087 ( .A(n1290), .B(n1289), .Z(n4867) );
  NAND U2088 ( .A(n1291), .B(n4867), .Z(n1292) );
  NANDN U2089 ( .A(n4870), .B(n1292), .Z(n1295) );
  NANDN U2090 ( .A(x[299]), .B(y[299]), .Z(n1294) );
  NANDN U2091 ( .A(x[300]), .B(y[300]), .Z(n1293) );
  AND U2092 ( .A(n1294), .B(n1293), .Z(n4871) );
  NAND U2093 ( .A(n1295), .B(n4871), .Z(n1298) );
  NANDN U2094 ( .A(y[301]), .B(x[301]), .Z(n1297) );
  NANDN U2095 ( .A(y[300]), .B(x[300]), .Z(n1296) );
  NAND U2096 ( .A(n1297), .B(n1296), .Z(n4874) );
  ANDN U2097 ( .B(n1298), .A(n4874), .Z(n1299) );
  OR U2098 ( .A(n4875), .B(n1299), .Z(n1300) );
  NANDN U2099 ( .A(n4878), .B(n1300), .Z(n1301) );
  NANDN U2100 ( .A(x[304]), .B(y[304]), .Z(n4879) );
  NAND U2101 ( .A(n1301), .B(n4879), .Z(n1302) );
  NANDN U2102 ( .A(n4882), .B(n1302), .Z(n1305) );
  NANDN U2103 ( .A(x[305]), .B(y[305]), .Z(n1304) );
  NANDN U2104 ( .A(x[306]), .B(y[306]), .Z(n1303) );
  AND U2105 ( .A(n1304), .B(n1303), .Z(n4883) );
  NAND U2106 ( .A(n1305), .B(n4883), .Z(n1308) );
  NANDN U2107 ( .A(y[307]), .B(x[307]), .Z(n1307) );
  NANDN U2108 ( .A(y[306]), .B(x[306]), .Z(n1306) );
  NAND U2109 ( .A(n1307), .B(n1306), .Z(n4886) );
  ANDN U2110 ( .B(n1308), .A(n4886), .Z(n1311) );
  NANDN U2111 ( .A(x[307]), .B(y[307]), .Z(n1310) );
  NANDN U2112 ( .A(x[308]), .B(y[308]), .Z(n1309) );
  AND U2113 ( .A(n1310), .B(n1309), .Z(n4888) );
  NANDN U2114 ( .A(n1311), .B(n4888), .Z(n1312) );
  NANDN U2115 ( .A(n4890), .B(n1312), .Z(n1315) );
  NANDN U2116 ( .A(x[309]), .B(y[309]), .Z(n1314) );
  NANDN U2117 ( .A(x[310]), .B(y[310]), .Z(n1313) );
  AND U2118 ( .A(n1314), .B(n1313), .Z(n4891) );
  NAND U2119 ( .A(n1315), .B(n4891), .Z(n1316) );
  NANDN U2120 ( .A(n4894), .B(n1316), .Z(n1317) );
  NANDN U2121 ( .A(n4896), .B(n1317), .Z(n1320) );
  NANDN U2122 ( .A(y[312]), .B(x[312]), .Z(n3464) );
  ANDN U2123 ( .B(x[313]), .A(y[313]), .Z(n3467) );
  ANDN U2124 ( .B(n3464), .A(n3467), .Z(n1318) );
  ANDN U2125 ( .B(n1319), .A(n1318), .Z(n4898) );
  ANDN U2126 ( .B(n1320), .A(n4898), .Z(n1321) );
  NANDN U2127 ( .A(x[314]), .B(y[314]), .Z(n4900) );
  NANDN U2128 ( .A(n1321), .B(n4900), .Z(n1322) );
  NANDN U2129 ( .A(n4902), .B(n1322), .Z(n1325) );
  NANDN U2130 ( .A(x[315]), .B(y[315]), .Z(n1324) );
  NANDN U2131 ( .A(x[316]), .B(y[316]), .Z(n1323) );
  AND U2132 ( .A(n1324), .B(n1323), .Z(n4903) );
  NAND U2133 ( .A(n1325), .B(n4903), .Z(n1326) );
  NANDN U2134 ( .A(n4906), .B(n1326), .Z(n1329) );
  NANDN U2135 ( .A(x[317]), .B(y[317]), .Z(n1328) );
  NANDN U2136 ( .A(x[318]), .B(y[318]), .Z(n1327) );
  AND U2137 ( .A(n1328), .B(n1327), .Z(n4907) );
  NAND U2138 ( .A(n1329), .B(n4907), .Z(n1332) );
  NANDN U2139 ( .A(y[319]), .B(x[319]), .Z(n1331) );
  NANDN U2140 ( .A(y[318]), .B(x[318]), .Z(n1330) );
  NAND U2141 ( .A(n1331), .B(n1330), .Z(n4910) );
  ANDN U2142 ( .B(n1332), .A(n4910), .Z(n1335) );
  NANDN U2143 ( .A(x[319]), .B(y[319]), .Z(n1334) );
  NANDN U2144 ( .A(x[320]), .B(y[320]), .Z(n1333) );
  AND U2145 ( .A(n1334), .B(n1333), .Z(n4912) );
  NANDN U2146 ( .A(n1335), .B(n4912), .Z(n1336) );
  NANDN U2147 ( .A(n4914), .B(n1336), .Z(n1339) );
  NANDN U2148 ( .A(x[321]), .B(y[321]), .Z(n1338) );
  NANDN U2149 ( .A(x[322]), .B(y[322]), .Z(n1337) );
  AND U2150 ( .A(n1338), .B(n1337), .Z(n4915) );
  NAND U2151 ( .A(n1339), .B(n4915), .Z(n1340) );
  NANDN U2152 ( .A(n4918), .B(n1340), .Z(n1345) );
  NANDN U2153 ( .A(x[324]), .B(y[324]), .Z(n1342) );
  NANDN U2154 ( .A(x[323]), .B(y[323]), .Z(n1341) );
  AND U2155 ( .A(n1342), .B(n1341), .Z(n1344) );
  NANDN U2156 ( .A(x[325]), .B(y[325]), .Z(n1343) );
  AND U2157 ( .A(n1344), .B(n1343), .Z(n4919) );
  NAND U2158 ( .A(n1345), .B(n4919), .Z(n1354) );
  NANDN U2159 ( .A(y[327]), .B(x[327]), .Z(n1347) );
  NANDN U2160 ( .A(y[326]), .B(x[326]), .Z(n1346) );
  AND U2161 ( .A(n1347), .B(n1346), .Z(n1353) );
  NANDN U2162 ( .A(y[324]), .B(x[324]), .Z(n1348) );
  NANDN U2163 ( .A(x[325]), .B(n1348), .Z(n1351) );
  XNOR U2164 ( .A(n1348), .B(x[325]), .Z(n1349) );
  NAND U2165 ( .A(n1349), .B(y[325]), .Z(n1350) );
  NAND U2166 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U2167 ( .A(n1353), .B(n1352), .Z(n4922) );
  ANDN U2168 ( .B(n1354), .A(n4922), .Z(n1361) );
  NANDN U2169 ( .A(x[327]), .B(y[327]), .Z(n1356) );
  ANDN U2170 ( .B(y[328]), .A(x[328]), .Z(n1355) );
  ANDN U2171 ( .B(n1356), .A(n1355), .Z(n1360) );
  XNOR U2172 ( .A(y[327]), .B(x[327]), .Z(n1358) );
  ANDN U2173 ( .B(y[326]), .A(x[326]), .Z(n1357) );
  NAND U2174 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U2175 ( .A(n1360), .B(n1359), .Z(n4924) );
  NANDN U2176 ( .A(n1361), .B(n4924), .Z(n1362) );
  NANDN U2177 ( .A(n4926), .B(n1362), .Z(n1363) );
  NANDN U2178 ( .A(n4928), .B(n1363), .Z(n1364) );
  NANDN U2179 ( .A(n4930), .B(n1364), .Z(n1365) );
  NANDN U2180 ( .A(x[332]), .B(y[332]), .Z(n4931) );
  NAND U2181 ( .A(n1365), .B(n4931), .Z(n1368) );
  NANDN U2182 ( .A(y[333]), .B(x[333]), .Z(n1367) );
  NANDN U2183 ( .A(y[332]), .B(x[332]), .Z(n1366) );
  NAND U2184 ( .A(n1367), .B(n1366), .Z(n4934) );
  ANDN U2185 ( .B(n1368), .A(n4934), .Z(n1371) );
  NANDN U2186 ( .A(x[333]), .B(y[333]), .Z(n1370) );
  NANDN U2187 ( .A(x[334]), .B(y[334]), .Z(n1369) );
  AND U2188 ( .A(n1370), .B(n1369), .Z(n4936) );
  NANDN U2189 ( .A(n1371), .B(n4936), .Z(n1372) );
  NANDN U2190 ( .A(n4938), .B(n1372), .Z(n1375) );
  NANDN U2191 ( .A(x[335]), .B(y[335]), .Z(n1374) );
  NANDN U2192 ( .A(x[336]), .B(y[336]), .Z(n1373) );
  AND U2193 ( .A(n1374), .B(n1373), .Z(n4939) );
  NAND U2194 ( .A(n1375), .B(n4939), .Z(n1376) );
  NANDN U2195 ( .A(n4942), .B(n1376), .Z(n1379) );
  NANDN U2196 ( .A(x[337]), .B(y[337]), .Z(n1378) );
  NANDN U2197 ( .A(x[338]), .B(y[338]), .Z(n1377) );
  AND U2198 ( .A(n1378), .B(n1377), .Z(n4943) );
  NAND U2199 ( .A(n1379), .B(n4943), .Z(n1382) );
  NANDN U2200 ( .A(y[339]), .B(x[339]), .Z(n1381) );
  NANDN U2201 ( .A(y[338]), .B(x[338]), .Z(n1380) );
  NAND U2202 ( .A(n1381), .B(n1380), .Z(n4946) );
  ANDN U2203 ( .B(n1382), .A(n4946), .Z(n1385) );
  NANDN U2204 ( .A(x[339]), .B(y[339]), .Z(n1384) );
  NANDN U2205 ( .A(x[340]), .B(y[340]), .Z(n1383) );
  AND U2206 ( .A(n1384), .B(n1383), .Z(n4948) );
  NANDN U2207 ( .A(n1385), .B(n4948), .Z(n1386) );
  NANDN U2208 ( .A(n4950), .B(n1386), .Z(n1389) );
  NANDN U2209 ( .A(x[341]), .B(y[341]), .Z(n1388) );
  NANDN U2210 ( .A(x[342]), .B(y[342]), .Z(n1387) );
  AND U2211 ( .A(n1388), .B(n1387), .Z(n4951) );
  NAND U2212 ( .A(n1389), .B(n4951), .Z(n1390) );
  NANDN U2213 ( .A(n4954), .B(n1390), .Z(n1393) );
  NANDN U2214 ( .A(x[343]), .B(y[343]), .Z(n1392) );
  NANDN U2215 ( .A(x[344]), .B(y[344]), .Z(n1391) );
  AND U2216 ( .A(n1392), .B(n1391), .Z(n4955) );
  NAND U2217 ( .A(n1393), .B(n4955), .Z(n1396) );
  NANDN U2218 ( .A(y[345]), .B(x[345]), .Z(n1395) );
  NANDN U2219 ( .A(y[344]), .B(x[344]), .Z(n1394) );
  NAND U2220 ( .A(n1395), .B(n1394), .Z(n4958) );
  ANDN U2221 ( .B(n1396), .A(n4958), .Z(n1399) );
  NANDN U2222 ( .A(x[345]), .B(y[345]), .Z(n1398) );
  NANDN U2223 ( .A(x[346]), .B(y[346]), .Z(n1397) );
  AND U2224 ( .A(n1398), .B(n1397), .Z(n4960) );
  NANDN U2225 ( .A(n1399), .B(n4960), .Z(n1400) );
  NANDN U2226 ( .A(n4962), .B(n1400), .Z(n1403) );
  NANDN U2227 ( .A(x[347]), .B(y[347]), .Z(n1402) );
  NANDN U2228 ( .A(x[348]), .B(y[348]), .Z(n1401) );
  AND U2229 ( .A(n1402), .B(n1401), .Z(n4963) );
  NAND U2230 ( .A(n1403), .B(n4963), .Z(n1404) );
  NANDN U2231 ( .A(n4966), .B(n1404), .Z(n1405) );
  NANDN U2232 ( .A(n3510), .B(n1405), .Z(n1408) );
  NANDN U2233 ( .A(y[350]), .B(x[350]), .Z(n4969) );
  ANDN U2234 ( .B(x[351]), .A(y[351]), .Z(n4973) );
  ANDN U2235 ( .B(n4969), .A(n4973), .Z(n1406) );
  ANDN U2236 ( .B(n1407), .A(n1406), .Z(n3512) );
  ANDN U2237 ( .B(n1408), .A(n3512), .Z(n1409) );
  NANDN U2238 ( .A(x[352]), .B(y[352]), .Z(n4975) );
  NANDN U2239 ( .A(n1409), .B(n4975), .Z(n1410) );
  NANDN U2240 ( .A(n4978), .B(n1410), .Z(n1413) );
  NANDN U2241 ( .A(x[353]), .B(y[353]), .Z(n1412) );
  NANDN U2242 ( .A(x[354]), .B(y[354]), .Z(n1411) );
  AND U2243 ( .A(n1412), .B(n1411), .Z(n4980) );
  NAND U2244 ( .A(n1413), .B(n4980), .Z(n1414) );
  NANDN U2245 ( .A(n4982), .B(n1414), .Z(n1417) );
  NANDN U2246 ( .A(x[355]), .B(y[355]), .Z(n1416) );
  NANDN U2247 ( .A(x[356]), .B(y[356]), .Z(n1415) );
  AND U2248 ( .A(n1416), .B(n1415), .Z(n4983) );
  NAND U2249 ( .A(n1417), .B(n4983), .Z(n1420) );
  NANDN U2250 ( .A(y[356]), .B(x[356]), .Z(n1419) );
  NANDN U2251 ( .A(y[357]), .B(x[357]), .Z(n1418) );
  NAND U2252 ( .A(n1419), .B(n1418), .Z(n4986) );
  ANDN U2253 ( .B(n1420), .A(n4986), .Z(n1421) );
  OR U2254 ( .A(n3520), .B(n1421), .Z(n1422) );
  NANDN U2255 ( .A(n3522), .B(n1422), .Z(n1423) );
  NANDN U2256 ( .A(x[360]), .B(y[360]), .Z(n4995) );
  NAND U2257 ( .A(n1423), .B(n4995), .Z(n1424) );
  NANDN U2258 ( .A(n4998), .B(n1424), .Z(n1428) );
  NANDN U2259 ( .A(x[362]), .B(y[362]), .Z(n1426) );
  NANDN U2260 ( .A(x[361]), .B(y[361]), .Z(n1425) );
  AND U2261 ( .A(n1426), .B(n1425), .Z(n1427) );
  NANDN U2262 ( .A(x[363]), .B(y[363]), .Z(n1432) );
  AND U2263 ( .A(n1427), .B(n1432), .Z(n5000) );
  NAND U2264 ( .A(n1428), .B(n5000), .Z(n1433) );
  XNOR U2265 ( .A(x[363]), .B(y[363]), .Z(n1430) );
  NANDN U2266 ( .A(y[362]), .B(x[362]), .Z(n1429) );
  NAND U2267 ( .A(n1430), .B(n1429), .Z(n1431) );
  AND U2268 ( .A(n1432), .B(n1431), .Z(n5001) );
  ANDN U2269 ( .B(n1433), .A(n5001), .Z(n1434) );
  OR U2270 ( .A(n5005), .B(n1434), .Z(n1435) );
  NANDN U2271 ( .A(n3529), .B(n1435), .Z(n1436) );
  NANDN U2272 ( .A(n3531), .B(n1436), .Z(n1437) );
  NANDN U2273 ( .A(n3532), .B(n1437), .Z(n1440) );
  NANDN U2274 ( .A(x[369]), .B(y[369]), .Z(n1439) );
  NANDN U2275 ( .A(x[370]), .B(y[370]), .Z(n1438) );
  AND U2276 ( .A(n1439), .B(n1438), .Z(n5015) );
  NAND U2277 ( .A(n1440), .B(n5015), .Z(n1443) );
  NANDN U2278 ( .A(y[371]), .B(x[371]), .Z(n1442) );
  NANDN U2279 ( .A(y[370]), .B(x[370]), .Z(n1441) );
  NAND U2280 ( .A(n1442), .B(n1441), .Z(n5018) );
  ANDN U2281 ( .B(n1443), .A(n5018), .Z(n1446) );
  NANDN U2282 ( .A(x[371]), .B(y[371]), .Z(n1445) );
  NANDN U2283 ( .A(x[372]), .B(y[372]), .Z(n1444) );
  AND U2284 ( .A(n1445), .B(n1444), .Z(n5019) );
  NANDN U2285 ( .A(n1446), .B(n5019), .Z(n1447) );
  NANDN U2286 ( .A(n5022), .B(n1447), .Z(n1450) );
  NANDN U2287 ( .A(x[373]), .B(y[373]), .Z(n1449) );
  NANDN U2288 ( .A(x[374]), .B(y[374]), .Z(n1448) );
  AND U2289 ( .A(n1449), .B(n1448), .Z(n5023) );
  NAND U2290 ( .A(n1450), .B(n5023), .Z(n1451) );
  NANDN U2291 ( .A(n5025), .B(n1451), .Z(n1454) );
  NANDN U2292 ( .A(x[375]), .B(y[375]), .Z(n1453) );
  NANDN U2293 ( .A(x[376]), .B(y[376]), .Z(n1452) );
  AND U2294 ( .A(n1453), .B(n1452), .Z(n5027) );
  NAND U2295 ( .A(n1454), .B(n5027), .Z(n1457) );
  NANDN U2296 ( .A(y[377]), .B(x[377]), .Z(n1456) );
  NANDN U2297 ( .A(y[376]), .B(x[376]), .Z(n1455) );
  NAND U2298 ( .A(n1456), .B(n1455), .Z(n5030) );
  ANDN U2299 ( .B(n1457), .A(n5030), .Z(n1460) );
  NANDN U2300 ( .A(x[377]), .B(y[377]), .Z(n1459) );
  NANDN U2301 ( .A(x[378]), .B(y[378]), .Z(n1458) );
  AND U2302 ( .A(n1459), .B(n1458), .Z(n5031) );
  NANDN U2303 ( .A(n1460), .B(n5031), .Z(n1461) );
  NANDN U2304 ( .A(n5034), .B(n1461), .Z(n1464) );
  NANDN U2305 ( .A(x[379]), .B(y[379]), .Z(n1463) );
  NANDN U2306 ( .A(x[380]), .B(y[380]), .Z(n1462) );
  AND U2307 ( .A(n1463), .B(n1462), .Z(n5035) );
  NAND U2308 ( .A(n1464), .B(n5035), .Z(n1465) );
  NANDN U2309 ( .A(n5037), .B(n1465), .Z(n1466) );
  NANDN U2310 ( .A(x[381]), .B(y[381]), .Z(n5039) );
  NAND U2311 ( .A(n1466), .B(n5039), .Z(n1469) );
  NANDN U2312 ( .A(y[382]), .B(x[382]), .Z(n1467) );
  NAND U2313 ( .A(n1468), .B(n1467), .Z(n5042) );
  ANDN U2314 ( .B(n1469), .A(n5042), .Z(n1470) );
  ANDN U2315 ( .B(n2952), .A(n1470), .Z(n1471) );
  NANDN U2316 ( .A(n5044), .B(n1471), .Z(n1472) );
  NANDN U2317 ( .A(n5046), .B(n1472), .Z(n1473) );
  NANDN U2318 ( .A(n2954), .B(n1473), .Z(n1478) );
  XNOR U2319 ( .A(x[387]), .B(y[387]), .Z(n1475) );
  NANDN U2320 ( .A(y[386]), .B(x[386]), .Z(n1474) );
  NAND U2321 ( .A(n1475), .B(n1474), .Z(n1476) );
  NAND U2322 ( .A(n1477), .B(n1476), .Z(n5050) );
  NAND U2323 ( .A(n1478), .B(n5050), .Z(n1479) );
  AND U2324 ( .A(n5051), .B(n1479), .Z(n1482) );
  NANDN U2325 ( .A(y[389]), .B(x[389]), .Z(n1481) );
  NANDN U2326 ( .A(y[388]), .B(x[388]), .Z(n1480) );
  AND U2327 ( .A(n1481), .B(n1480), .Z(n5053) );
  NANDN U2328 ( .A(n1482), .B(n5053), .Z(n1485) );
  NANDN U2329 ( .A(x[389]), .B(y[389]), .Z(n1484) );
  NANDN U2330 ( .A(x[390]), .B(y[390]), .Z(n1483) );
  AND U2331 ( .A(n1484), .B(n1483), .Z(n5056) );
  NAND U2332 ( .A(n1485), .B(n5056), .Z(n1488) );
  NANDN U2333 ( .A(y[391]), .B(x[391]), .Z(n1487) );
  NANDN U2334 ( .A(y[390]), .B(x[390]), .Z(n1486) );
  AND U2335 ( .A(n1487), .B(n1486), .Z(n5057) );
  NAND U2336 ( .A(n1488), .B(n5057), .Z(n1491) );
  NANDN U2337 ( .A(x[391]), .B(y[391]), .Z(n1490) );
  NANDN U2338 ( .A(x[392]), .B(y[392]), .Z(n1489) );
  AND U2339 ( .A(n1490), .B(n1489), .Z(n5059) );
  NAND U2340 ( .A(n1491), .B(n5059), .Z(n1494) );
  NANDN U2341 ( .A(y[393]), .B(x[393]), .Z(n1493) );
  NANDN U2342 ( .A(y[392]), .B(x[392]), .Z(n1492) );
  AND U2343 ( .A(n1493), .B(n1492), .Z(n5061) );
  NAND U2344 ( .A(n1494), .B(n5061), .Z(n1495) );
  AND U2345 ( .A(n5063), .B(n1495), .Z(n1498) );
  NANDN U2346 ( .A(y[395]), .B(x[395]), .Z(n1497) );
  NANDN U2347 ( .A(y[394]), .B(x[394]), .Z(n1496) );
  AND U2348 ( .A(n1497), .B(n1496), .Z(n5065) );
  NANDN U2349 ( .A(n1498), .B(n5065), .Z(n1501) );
  NANDN U2350 ( .A(x[395]), .B(y[395]), .Z(n1500) );
  NANDN U2351 ( .A(x[396]), .B(y[396]), .Z(n1499) );
  AND U2352 ( .A(n1500), .B(n1499), .Z(n5068) );
  NAND U2353 ( .A(n1501), .B(n5068), .Z(n1504) );
  NANDN U2354 ( .A(y[397]), .B(x[397]), .Z(n1503) );
  NANDN U2355 ( .A(y[396]), .B(x[396]), .Z(n1502) );
  AND U2356 ( .A(n1503), .B(n1502), .Z(n5069) );
  NAND U2357 ( .A(n1504), .B(n5069), .Z(n1507) );
  NANDN U2358 ( .A(x[397]), .B(y[397]), .Z(n1506) );
  NANDN U2359 ( .A(x[398]), .B(y[398]), .Z(n1505) );
  AND U2360 ( .A(n1506), .B(n1505), .Z(n5071) );
  NAND U2361 ( .A(n1507), .B(n5071), .Z(n1510) );
  NANDN U2362 ( .A(y[399]), .B(x[399]), .Z(n1509) );
  NANDN U2363 ( .A(y[398]), .B(x[398]), .Z(n1508) );
  AND U2364 ( .A(n1509), .B(n1508), .Z(n5073) );
  NAND U2365 ( .A(n1510), .B(n5073), .Z(n1511) );
  AND U2366 ( .A(n5075), .B(n1511), .Z(n1514) );
  NANDN U2367 ( .A(y[401]), .B(x[401]), .Z(n1513) );
  NANDN U2368 ( .A(y[400]), .B(x[400]), .Z(n1512) );
  AND U2369 ( .A(n1513), .B(n1512), .Z(n5077) );
  NANDN U2370 ( .A(n1514), .B(n5077), .Z(n1517) );
  NANDN U2371 ( .A(x[401]), .B(y[401]), .Z(n1516) );
  NANDN U2372 ( .A(x[402]), .B(y[402]), .Z(n1515) );
  AND U2373 ( .A(n1516), .B(n1515), .Z(n5080) );
  NAND U2374 ( .A(n1517), .B(n5080), .Z(n1520) );
  NANDN U2375 ( .A(y[403]), .B(x[403]), .Z(n1519) );
  NANDN U2376 ( .A(y[402]), .B(x[402]), .Z(n1518) );
  AND U2377 ( .A(n1519), .B(n1518), .Z(n5081) );
  NAND U2378 ( .A(n1520), .B(n5081), .Z(n1523) );
  NANDN U2379 ( .A(x[403]), .B(y[403]), .Z(n1522) );
  NANDN U2380 ( .A(x[404]), .B(y[404]), .Z(n1521) );
  AND U2381 ( .A(n1522), .B(n1521), .Z(n5083) );
  NAND U2382 ( .A(n1523), .B(n5083), .Z(n1526) );
  NANDN U2383 ( .A(y[405]), .B(x[405]), .Z(n1525) );
  NANDN U2384 ( .A(y[404]), .B(x[404]), .Z(n1524) );
  AND U2385 ( .A(n1525), .B(n1524), .Z(n5085) );
  NAND U2386 ( .A(n1526), .B(n5085), .Z(n1528) );
  NANDN U2387 ( .A(x[405]), .B(y[405]), .Z(n3573) );
  NANDN U2388 ( .A(n3578), .B(n3573), .Z(n5088) );
  ANDN U2389 ( .B(n1528), .A(n5088), .Z(n1529) );
  OR U2390 ( .A(n5090), .B(n1529), .Z(n1530) );
  NANDN U2391 ( .A(x[408]), .B(y[408]), .Z(n5092) );
  NAND U2392 ( .A(n1530), .B(n5092), .Z(n1533) );
  NANDN U2393 ( .A(y[409]), .B(x[409]), .Z(n1532) );
  NANDN U2394 ( .A(y[408]), .B(x[408]), .Z(n1531) );
  AND U2395 ( .A(n1532), .B(n1531), .Z(n5093) );
  NAND U2396 ( .A(n1533), .B(n5093), .Z(n1536) );
  NANDN U2397 ( .A(x[409]), .B(y[409]), .Z(n1535) );
  NANDN U2398 ( .A(x[410]), .B(y[410]), .Z(n1534) );
  AND U2399 ( .A(n1535), .B(n1534), .Z(n5095) );
  NAND U2400 ( .A(n1536), .B(n5095), .Z(n1539) );
  NANDN U2401 ( .A(y[411]), .B(x[411]), .Z(n1538) );
  NANDN U2402 ( .A(y[410]), .B(x[410]), .Z(n1537) );
  AND U2403 ( .A(n1538), .B(n1537), .Z(n5097) );
  NAND U2404 ( .A(n1539), .B(n5097), .Z(n1540) );
  AND U2405 ( .A(n5099), .B(n1540), .Z(n1543) );
  NANDN U2406 ( .A(y[413]), .B(x[413]), .Z(n1542) );
  NANDN U2407 ( .A(y[412]), .B(x[412]), .Z(n1541) );
  AND U2408 ( .A(n1542), .B(n1541), .Z(n5101) );
  NANDN U2409 ( .A(n1543), .B(n5101), .Z(n1546) );
  NANDN U2410 ( .A(x[413]), .B(y[413]), .Z(n1545) );
  NANDN U2411 ( .A(x[414]), .B(y[414]), .Z(n1544) );
  AND U2412 ( .A(n1545), .B(n1544), .Z(n5104) );
  NAND U2413 ( .A(n1546), .B(n5104), .Z(n1549) );
  NANDN U2414 ( .A(y[415]), .B(x[415]), .Z(n1548) );
  NANDN U2415 ( .A(y[414]), .B(x[414]), .Z(n1547) );
  AND U2416 ( .A(n1548), .B(n1547), .Z(n5105) );
  NAND U2417 ( .A(n1549), .B(n5105), .Z(n1552) );
  NANDN U2418 ( .A(x[415]), .B(y[415]), .Z(n1551) );
  NANDN U2419 ( .A(x[416]), .B(y[416]), .Z(n1550) );
  AND U2420 ( .A(n1551), .B(n1550), .Z(n5107) );
  NAND U2421 ( .A(n1552), .B(n5107), .Z(n1555) );
  NANDN U2422 ( .A(y[417]), .B(x[417]), .Z(n1554) );
  NANDN U2423 ( .A(y[416]), .B(x[416]), .Z(n1553) );
  AND U2424 ( .A(n1554), .B(n1553), .Z(n5109) );
  NAND U2425 ( .A(n1555), .B(n5109), .Z(n1556) );
  AND U2426 ( .A(n5111), .B(n1556), .Z(n1559) );
  NANDN U2427 ( .A(y[419]), .B(x[419]), .Z(n1558) );
  NANDN U2428 ( .A(y[418]), .B(x[418]), .Z(n1557) );
  AND U2429 ( .A(n1558), .B(n1557), .Z(n5113) );
  NANDN U2430 ( .A(n1559), .B(n5113), .Z(n1562) );
  NANDN U2431 ( .A(x[419]), .B(y[419]), .Z(n1561) );
  NANDN U2432 ( .A(x[420]), .B(y[420]), .Z(n1560) );
  AND U2433 ( .A(n1561), .B(n1560), .Z(n5116) );
  NAND U2434 ( .A(n1562), .B(n5116), .Z(n1565) );
  NANDN U2435 ( .A(y[421]), .B(x[421]), .Z(n1564) );
  NANDN U2436 ( .A(y[420]), .B(x[420]), .Z(n1563) );
  AND U2437 ( .A(n1564), .B(n1563), .Z(n5117) );
  NAND U2438 ( .A(n1565), .B(n5117), .Z(n1568) );
  NANDN U2439 ( .A(x[421]), .B(y[421]), .Z(n1567) );
  NANDN U2440 ( .A(x[422]), .B(y[422]), .Z(n1566) );
  AND U2441 ( .A(n1567), .B(n1566), .Z(n5119) );
  NAND U2442 ( .A(n1568), .B(n5119), .Z(n1571) );
  NANDN U2443 ( .A(y[423]), .B(x[423]), .Z(n1570) );
  NANDN U2444 ( .A(y[422]), .B(x[422]), .Z(n1569) );
  AND U2445 ( .A(n1570), .B(n1569), .Z(n5121) );
  NAND U2446 ( .A(n1571), .B(n5121), .Z(n1572) );
  AND U2447 ( .A(n5123), .B(n1572), .Z(n1575) );
  NANDN U2448 ( .A(y[425]), .B(x[425]), .Z(n1574) );
  NANDN U2449 ( .A(y[424]), .B(x[424]), .Z(n1573) );
  AND U2450 ( .A(n1574), .B(n1573), .Z(n5125) );
  NANDN U2451 ( .A(n1575), .B(n5125), .Z(n1578) );
  NANDN U2452 ( .A(x[425]), .B(y[425]), .Z(n1577) );
  NANDN U2453 ( .A(x[426]), .B(y[426]), .Z(n1576) );
  AND U2454 ( .A(n1577), .B(n1576), .Z(n5128) );
  NAND U2455 ( .A(n1578), .B(n5128), .Z(n1581) );
  NANDN U2456 ( .A(y[427]), .B(x[427]), .Z(n1580) );
  NANDN U2457 ( .A(y[426]), .B(x[426]), .Z(n1579) );
  AND U2458 ( .A(n1580), .B(n1579), .Z(n5129) );
  NAND U2459 ( .A(n1581), .B(n5129), .Z(n1584) );
  NANDN U2460 ( .A(x[427]), .B(y[427]), .Z(n1583) );
  NANDN U2461 ( .A(x[428]), .B(y[428]), .Z(n1582) );
  AND U2462 ( .A(n1583), .B(n1582), .Z(n5131) );
  NAND U2463 ( .A(n1584), .B(n5131), .Z(n1587) );
  NANDN U2464 ( .A(y[429]), .B(x[429]), .Z(n1586) );
  NANDN U2465 ( .A(y[428]), .B(x[428]), .Z(n1585) );
  AND U2466 ( .A(n1586), .B(n1585), .Z(n5133) );
  NAND U2467 ( .A(n1587), .B(n5133), .Z(n1588) );
  AND U2468 ( .A(n5135), .B(n1588), .Z(n1591) );
  NANDN U2469 ( .A(y[431]), .B(x[431]), .Z(n1590) );
  NANDN U2470 ( .A(y[430]), .B(x[430]), .Z(n1589) );
  AND U2471 ( .A(n1590), .B(n1589), .Z(n5137) );
  NANDN U2472 ( .A(n1591), .B(n5137), .Z(n1594) );
  NANDN U2473 ( .A(x[431]), .B(y[431]), .Z(n1593) );
  NANDN U2474 ( .A(x[432]), .B(y[432]), .Z(n1592) );
  AND U2475 ( .A(n1593), .B(n1592), .Z(n5140) );
  NAND U2476 ( .A(n1594), .B(n5140), .Z(n1597) );
  NANDN U2477 ( .A(y[433]), .B(x[433]), .Z(n1596) );
  NANDN U2478 ( .A(y[432]), .B(x[432]), .Z(n1595) );
  AND U2479 ( .A(n1596), .B(n1595), .Z(n5141) );
  NAND U2480 ( .A(n1597), .B(n5141), .Z(n1600) );
  NANDN U2481 ( .A(x[433]), .B(y[433]), .Z(n1599) );
  NANDN U2482 ( .A(x[434]), .B(y[434]), .Z(n1598) );
  AND U2483 ( .A(n1599), .B(n1598), .Z(n5143) );
  NAND U2484 ( .A(n1600), .B(n5143), .Z(n1603) );
  NANDN U2485 ( .A(y[435]), .B(x[435]), .Z(n1602) );
  NANDN U2486 ( .A(y[434]), .B(x[434]), .Z(n1601) );
  AND U2487 ( .A(n1602), .B(n1601), .Z(n5145) );
  NAND U2488 ( .A(n1603), .B(n5145), .Z(n1604) );
  AND U2489 ( .A(n5147), .B(n1604), .Z(n1607) );
  NANDN U2490 ( .A(y[437]), .B(x[437]), .Z(n1606) );
  NANDN U2491 ( .A(y[436]), .B(x[436]), .Z(n1605) );
  AND U2492 ( .A(n1606), .B(n1605), .Z(n5149) );
  NANDN U2493 ( .A(n1607), .B(n5149), .Z(n1610) );
  NANDN U2494 ( .A(x[437]), .B(y[437]), .Z(n1609) );
  NANDN U2495 ( .A(x[438]), .B(y[438]), .Z(n1608) );
  AND U2496 ( .A(n1609), .B(n1608), .Z(n5152) );
  NAND U2497 ( .A(n1610), .B(n5152), .Z(n1613) );
  NANDN U2498 ( .A(y[439]), .B(x[439]), .Z(n1612) );
  NANDN U2499 ( .A(y[438]), .B(x[438]), .Z(n1611) );
  AND U2500 ( .A(n1612), .B(n1611), .Z(n5153) );
  NAND U2501 ( .A(n1613), .B(n5153), .Z(n1616) );
  NANDN U2502 ( .A(x[439]), .B(y[439]), .Z(n1615) );
  NANDN U2503 ( .A(x[440]), .B(y[440]), .Z(n1614) );
  AND U2504 ( .A(n1615), .B(n1614), .Z(n5155) );
  NAND U2505 ( .A(n1616), .B(n5155), .Z(n1619) );
  NANDN U2506 ( .A(y[441]), .B(x[441]), .Z(n1618) );
  NANDN U2507 ( .A(y[440]), .B(x[440]), .Z(n1617) );
  AND U2508 ( .A(n1618), .B(n1617), .Z(n5157) );
  NAND U2509 ( .A(n1619), .B(n5157), .Z(n1620) );
  AND U2510 ( .A(n5159), .B(n1620), .Z(n1623) );
  NANDN U2511 ( .A(y[443]), .B(x[443]), .Z(n1622) );
  NANDN U2512 ( .A(y[442]), .B(x[442]), .Z(n1621) );
  AND U2513 ( .A(n1622), .B(n1621), .Z(n5161) );
  NANDN U2514 ( .A(n1623), .B(n5161), .Z(n1626) );
  NANDN U2515 ( .A(x[443]), .B(y[443]), .Z(n1625) );
  NANDN U2516 ( .A(x[444]), .B(y[444]), .Z(n1624) );
  AND U2517 ( .A(n1625), .B(n1624), .Z(n5164) );
  NAND U2518 ( .A(n1626), .B(n5164), .Z(n1629) );
  NANDN U2519 ( .A(y[445]), .B(x[445]), .Z(n1628) );
  NANDN U2520 ( .A(y[444]), .B(x[444]), .Z(n1627) );
  AND U2521 ( .A(n1628), .B(n1627), .Z(n5165) );
  NAND U2522 ( .A(n1629), .B(n5165), .Z(n1632) );
  NANDN U2523 ( .A(x[445]), .B(y[445]), .Z(n1631) );
  NANDN U2524 ( .A(x[446]), .B(y[446]), .Z(n1630) );
  AND U2525 ( .A(n1631), .B(n1630), .Z(n5167) );
  NAND U2526 ( .A(n1632), .B(n5167), .Z(n1635) );
  NANDN U2527 ( .A(y[447]), .B(x[447]), .Z(n1634) );
  NANDN U2528 ( .A(y[446]), .B(x[446]), .Z(n1633) );
  AND U2529 ( .A(n1634), .B(n1633), .Z(n5169) );
  NAND U2530 ( .A(n1635), .B(n5169), .Z(n1637) );
  NANDN U2531 ( .A(x[447]), .B(y[447]), .Z(n3621) );
  NANDN U2532 ( .A(n3626), .B(n3621), .Z(n5172) );
  ANDN U2533 ( .B(n1637), .A(n5172), .Z(n1638) );
  OR U2534 ( .A(n5174), .B(n1638), .Z(n1639) );
  NANDN U2535 ( .A(x[450]), .B(y[450]), .Z(n5176) );
  NAND U2536 ( .A(n1639), .B(n5176), .Z(n1642) );
  NANDN U2537 ( .A(y[450]), .B(x[450]), .Z(n1641) );
  NANDN U2538 ( .A(y[451]), .B(x[451]), .Z(n1640) );
  AND U2539 ( .A(n1641), .B(n1640), .Z(n5177) );
  NAND U2540 ( .A(n1642), .B(n5177), .Z(n1643) );
  NANDN U2541 ( .A(n5180), .B(n1643), .Z(n1646) );
  NANDN U2542 ( .A(y[452]), .B(x[452]), .Z(n1645) );
  NANDN U2543 ( .A(y[453]), .B(x[453]), .Z(n1644) );
  AND U2544 ( .A(n1645), .B(n1644), .Z(n5181) );
  NAND U2545 ( .A(n1646), .B(n5181), .Z(n1651) );
  NANDN U2546 ( .A(x[454]), .B(y[454]), .Z(n1648) );
  NANDN U2547 ( .A(x[453]), .B(y[453]), .Z(n1647) );
  AND U2548 ( .A(n1648), .B(n1647), .Z(n1650) );
  NANDN U2549 ( .A(x[455]), .B(y[455]), .Z(n1649) );
  NAND U2550 ( .A(n1650), .B(n1649), .Z(n5184) );
  ANDN U2551 ( .B(n1651), .A(n5184), .Z(n1652) );
  NANDN U2552 ( .A(n1652), .B(n5185), .Z(n1653) );
  NANDN U2553 ( .A(n5187), .B(n1653), .Z(n1654) );
  NANDN U2554 ( .A(n5190), .B(n1654), .Z(n1655) );
  NANDN U2555 ( .A(n5192), .B(n1655), .Z(n1656) );
  NANDN U2556 ( .A(n5194), .B(n1656), .Z(n1662) );
  XNOR U2557 ( .A(y[461]), .B(x[461]), .Z(n1658) );
  NANDN U2558 ( .A(x[460]), .B(y[460]), .Z(n1657) );
  NAND U2559 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U2560 ( .A(n1660), .B(n1659), .Z(n5196) );
  OR U2561 ( .A(n5196), .B(n5200), .Z(n3648) );
  ANDN U2562 ( .B(n1662), .A(n3648), .Z(n1663) );
  OR U2563 ( .A(n3650), .B(n1663), .Z(n1664) );
  NANDN U2564 ( .A(x[464]), .B(y[464]), .Z(n5203) );
  NAND U2565 ( .A(n1664), .B(n5203), .Z(n1667) );
  NANDN U2566 ( .A(y[464]), .B(x[464]), .Z(n1666) );
  NANDN U2567 ( .A(y[465]), .B(x[465]), .Z(n1665) );
  AND U2568 ( .A(n1666), .B(n1665), .Z(n5205) );
  NAND U2569 ( .A(n1667), .B(n5205), .Z(n1668) );
  NANDN U2570 ( .A(n5208), .B(n1668), .Z(n1671) );
  NANDN U2571 ( .A(y[466]), .B(x[466]), .Z(n1670) );
  NANDN U2572 ( .A(y[467]), .B(x[467]), .Z(n1669) );
  AND U2573 ( .A(n1670), .B(n1669), .Z(n5209) );
  NAND U2574 ( .A(n1671), .B(n5209), .Z(n1674) );
  NANDN U2575 ( .A(x[468]), .B(y[468]), .Z(n1673) );
  NANDN U2576 ( .A(x[467]), .B(y[467]), .Z(n1672) );
  NAND U2577 ( .A(n1673), .B(n1672), .Z(n5212) );
  ANDN U2578 ( .B(n1674), .A(n5212), .Z(n1677) );
  NANDN U2579 ( .A(y[468]), .B(x[468]), .Z(n1676) );
  NANDN U2580 ( .A(y[469]), .B(x[469]), .Z(n1675) );
  AND U2581 ( .A(n1676), .B(n1675), .Z(n5214) );
  NANDN U2582 ( .A(n1677), .B(n5214), .Z(n1678) );
  NANDN U2583 ( .A(n5216), .B(n1678), .Z(n1681) );
  NANDN U2584 ( .A(y[470]), .B(x[470]), .Z(n1680) );
  NANDN U2585 ( .A(y[471]), .B(x[471]), .Z(n1679) );
  AND U2586 ( .A(n1680), .B(n1679), .Z(n5217) );
  NAND U2587 ( .A(n1681), .B(n5217), .Z(n1682) );
  NANDN U2588 ( .A(n5220), .B(n1682), .Z(n1685) );
  NANDN U2589 ( .A(y[472]), .B(x[472]), .Z(n1684) );
  NANDN U2590 ( .A(y[473]), .B(x[473]), .Z(n1683) );
  AND U2591 ( .A(n1684), .B(n1683), .Z(n5221) );
  NAND U2592 ( .A(n1685), .B(n5221), .Z(n1688) );
  NANDN U2593 ( .A(x[474]), .B(y[474]), .Z(n1687) );
  NANDN U2594 ( .A(x[473]), .B(y[473]), .Z(n1686) );
  NAND U2595 ( .A(n1687), .B(n1686), .Z(n5224) );
  ANDN U2596 ( .B(n1688), .A(n5224), .Z(n1691) );
  NANDN U2597 ( .A(y[474]), .B(x[474]), .Z(n1690) );
  NANDN U2598 ( .A(y[475]), .B(x[475]), .Z(n1689) );
  AND U2599 ( .A(n1690), .B(n1689), .Z(n5226) );
  NANDN U2600 ( .A(n1691), .B(n5226), .Z(n1692) );
  NANDN U2601 ( .A(n5228), .B(n1692), .Z(n1695) );
  NANDN U2602 ( .A(y[476]), .B(x[476]), .Z(n1694) );
  NANDN U2603 ( .A(y[477]), .B(x[477]), .Z(n1693) );
  AND U2604 ( .A(n1694), .B(n1693), .Z(n5229) );
  NAND U2605 ( .A(n1695), .B(n5229), .Z(n1696) );
  NANDN U2606 ( .A(n5232), .B(n1696), .Z(n1699) );
  NANDN U2607 ( .A(y[478]), .B(x[478]), .Z(n1698) );
  NANDN U2608 ( .A(y[479]), .B(x[479]), .Z(n1697) );
  AND U2609 ( .A(n1698), .B(n1697), .Z(n5233) );
  NAND U2610 ( .A(n1699), .B(n5233), .Z(n1702) );
  NANDN U2611 ( .A(x[480]), .B(y[480]), .Z(n1701) );
  NANDN U2612 ( .A(x[479]), .B(y[479]), .Z(n1700) );
  NAND U2613 ( .A(n1701), .B(n1700), .Z(n5236) );
  ANDN U2614 ( .B(n1702), .A(n5236), .Z(n1705) );
  NANDN U2615 ( .A(y[480]), .B(x[480]), .Z(n1704) );
  NANDN U2616 ( .A(y[481]), .B(x[481]), .Z(n1703) );
  AND U2617 ( .A(n1704), .B(n1703), .Z(n5238) );
  NANDN U2618 ( .A(n1705), .B(n5238), .Z(n1706) );
  NANDN U2619 ( .A(n5240), .B(n1706), .Z(n1709) );
  NANDN U2620 ( .A(y[482]), .B(x[482]), .Z(n1708) );
  NANDN U2621 ( .A(y[483]), .B(x[483]), .Z(n1707) );
  AND U2622 ( .A(n1708), .B(n1707), .Z(n5241) );
  NAND U2623 ( .A(n1709), .B(n5241), .Z(n1710) );
  NANDN U2624 ( .A(n5244), .B(n1710), .Z(n1713) );
  NANDN U2625 ( .A(y[484]), .B(x[484]), .Z(n1712) );
  NANDN U2626 ( .A(y[485]), .B(x[485]), .Z(n1711) );
  AND U2627 ( .A(n1712), .B(n1711), .Z(n5245) );
  NAND U2628 ( .A(n1713), .B(n5245), .Z(n1716) );
  NANDN U2629 ( .A(x[486]), .B(y[486]), .Z(n1715) );
  NANDN U2630 ( .A(x[485]), .B(y[485]), .Z(n1714) );
  NAND U2631 ( .A(n1715), .B(n1714), .Z(n5248) );
  ANDN U2632 ( .B(n1716), .A(n5248), .Z(n1719) );
  NANDN U2633 ( .A(y[486]), .B(x[486]), .Z(n1718) );
  NANDN U2634 ( .A(y[487]), .B(x[487]), .Z(n1717) );
  AND U2635 ( .A(n1718), .B(n1717), .Z(n5250) );
  NANDN U2636 ( .A(n1719), .B(n5250), .Z(n1720) );
  NANDN U2637 ( .A(n5252), .B(n1720), .Z(n1723) );
  NANDN U2638 ( .A(y[488]), .B(x[488]), .Z(n1722) );
  NANDN U2639 ( .A(y[489]), .B(x[489]), .Z(n1721) );
  AND U2640 ( .A(n1722), .B(n1721), .Z(n5253) );
  NAND U2641 ( .A(n1723), .B(n5253), .Z(n1724) );
  NANDN U2642 ( .A(n5256), .B(n1724), .Z(n1727) );
  NANDN U2643 ( .A(y[490]), .B(x[490]), .Z(n1726) );
  NANDN U2644 ( .A(y[491]), .B(x[491]), .Z(n1725) );
  AND U2645 ( .A(n1726), .B(n1725), .Z(n5257) );
  NAND U2646 ( .A(n1727), .B(n5257), .Z(n1730) );
  NANDN U2647 ( .A(x[492]), .B(y[492]), .Z(n1729) );
  NANDN U2648 ( .A(x[491]), .B(y[491]), .Z(n1728) );
  NAND U2649 ( .A(n1729), .B(n1728), .Z(n5260) );
  ANDN U2650 ( .B(n1730), .A(n5260), .Z(n1733) );
  NANDN U2651 ( .A(y[492]), .B(x[492]), .Z(n1732) );
  NANDN U2652 ( .A(y[493]), .B(x[493]), .Z(n1731) );
  AND U2653 ( .A(n1732), .B(n1731), .Z(n5262) );
  NANDN U2654 ( .A(n1733), .B(n5262), .Z(n1734) );
  NANDN U2655 ( .A(n5264), .B(n1734), .Z(n1737) );
  NANDN U2656 ( .A(y[494]), .B(x[494]), .Z(n1736) );
  NANDN U2657 ( .A(y[495]), .B(x[495]), .Z(n1735) );
  AND U2658 ( .A(n1736), .B(n1735), .Z(n5265) );
  NAND U2659 ( .A(n1737), .B(n5265), .Z(n1738) );
  NANDN U2660 ( .A(n5268), .B(n1738), .Z(n1741) );
  NANDN U2661 ( .A(y[496]), .B(x[496]), .Z(n1740) );
  NANDN U2662 ( .A(y[497]), .B(x[497]), .Z(n1739) );
  AND U2663 ( .A(n1740), .B(n1739), .Z(n5269) );
  NAND U2664 ( .A(n1741), .B(n5269), .Z(n1744) );
  NANDN U2665 ( .A(x[498]), .B(y[498]), .Z(n1743) );
  NANDN U2666 ( .A(x[497]), .B(y[497]), .Z(n1742) );
  NAND U2667 ( .A(n1743), .B(n1742), .Z(n5272) );
  ANDN U2668 ( .B(n1744), .A(n5272), .Z(n1747) );
  NANDN U2669 ( .A(y[498]), .B(x[498]), .Z(n1746) );
  NANDN U2670 ( .A(y[499]), .B(x[499]), .Z(n1745) );
  AND U2671 ( .A(n1746), .B(n1745), .Z(n5274) );
  NANDN U2672 ( .A(n1747), .B(n5274), .Z(n1748) );
  NANDN U2673 ( .A(n5276), .B(n1748), .Z(n1751) );
  NANDN U2674 ( .A(y[500]), .B(x[500]), .Z(n1750) );
  NANDN U2675 ( .A(y[501]), .B(x[501]), .Z(n1749) );
  AND U2676 ( .A(n1750), .B(n1749), .Z(n5277) );
  NAND U2677 ( .A(n1751), .B(n5277), .Z(n1752) );
  NANDN U2678 ( .A(n5280), .B(n1752), .Z(n1755) );
  NANDN U2679 ( .A(y[502]), .B(x[502]), .Z(n1754) );
  NANDN U2680 ( .A(y[503]), .B(x[503]), .Z(n1753) );
  AND U2681 ( .A(n1754), .B(n1753), .Z(n5281) );
  NAND U2682 ( .A(n1755), .B(n5281), .Z(n1756) );
  AND U2683 ( .A(n5283), .B(n1756), .Z(n1759) );
  NANDN U2684 ( .A(y[504]), .B(x[504]), .Z(n1757) );
  ANDN U2685 ( .B(x[505]), .A(y[505]), .Z(n3697) );
  ANDN U2686 ( .B(n1757), .A(n3697), .Z(n3693) );
  NANDN U2687 ( .A(n3693), .B(n1758), .Z(n5286) );
  NANDN U2688 ( .A(n1759), .B(n5286), .Z(n1760) );
  NANDN U2689 ( .A(x[506]), .B(y[506]), .Z(n5287) );
  NAND U2690 ( .A(n1760), .B(n5287), .Z(n1763) );
  NANDN U2691 ( .A(y[506]), .B(x[506]), .Z(n1762) );
  NANDN U2692 ( .A(y[507]), .B(x[507]), .Z(n1761) );
  AND U2693 ( .A(n1762), .B(n1761), .Z(n5289) );
  NAND U2694 ( .A(n1763), .B(n5289), .Z(n1764) );
  NANDN U2695 ( .A(n5292), .B(n1764), .Z(n1767) );
  NANDN U2696 ( .A(y[508]), .B(x[508]), .Z(n1766) );
  NANDN U2697 ( .A(y[509]), .B(x[509]), .Z(n1765) );
  AND U2698 ( .A(n1766), .B(n1765), .Z(n5293) );
  NAND U2699 ( .A(n1767), .B(n5293), .Z(n1770) );
  NANDN U2700 ( .A(x[510]), .B(y[510]), .Z(n1769) );
  NANDN U2701 ( .A(x[509]), .B(y[509]), .Z(n1768) );
  NAND U2702 ( .A(n1769), .B(n1768), .Z(n5296) );
  ANDN U2703 ( .B(n1770), .A(n5296), .Z(n1773) );
  NANDN U2704 ( .A(y[510]), .B(x[510]), .Z(n1772) );
  NANDN U2705 ( .A(y[511]), .B(x[511]), .Z(n1771) );
  AND U2706 ( .A(n1772), .B(n1771), .Z(n5298) );
  NANDN U2707 ( .A(n1773), .B(n5298), .Z(n1774) );
  NANDN U2708 ( .A(n5300), .B(n1774), .Z(n1777) );
  NANDN U2709 ( .A(y[512]), .B(x[512]), .Z(n1776) );
  NANDN U2710 ( .A(y[513]), .B(x[513]), .Z(n1775) );
  AND U2711 ( .A(n1776), .B(n1775), .Z(n5301) );
  NAND U2712 ( .A(n1777), .B(n5301), .Z(n1778) );
  NANDN U2713 ( .A(n5304), .B(n1778), .Z(n1781) );
  NANDN U2714 ( .A(y[514]), .B(x[514]), .Z(n1780) );
  NANDN U2715 ( .A(y[515]), .B(x[515]), .Z(n1779) );
  AND U2716 ( .A(n1780), .B(n1779), .Z(n5305) );
  NAND U2717 ( .A(n1781), .B(n5305), .Z(n1784) );
  NANDN U2718 ( .A(x[516]), .B(y[516]), .Z(n1783) );
  NANDN U2719 ( .A(x[515]), .B(y[515]), .Z(n1782) );
  NAND U2720 ( .A(n1783), .B(n1782), .Z(n5308) );
  ANDN U2721 ( .B(n1784), .A(n5308), .Z(n1787) );
  NANDN U2722 ( .A(y[516]), .B(x[516]), .Z(n1786) );
  NANDN U2723 ( .A(y[517]), .B(x[517]), .Z(n1785) );
  AND U2724 ( .A(n1786), .B(n1785), .Z(n5310) );
  NANDN U2725 ( .A(n1787), .B(n5310), .Z(n1788) );
  NANDN U2726 ( .A(n5312), .B(n1788), .Z(n1791) );
  NANDN U2727 ( .A(y[518]), .B(x[518]), .Z(n1790) );
  NANDN U2728 ( .A(y[519]), .B(x[519]), .Z(n1789) );
  AND U2729 ( .A(n1790), .B(n1789), .Z(n5313) );
  NAND U2730 ( .A(n1791), .B(n5313), .Z(n1792) );
  NANDN U2731 ( .A(n5316), .B(n1792), .Z(n1795) );
  NANDN U2732 ( .A(y[520]), .B(x[520]), .Z(n1794) );
  NANDN U2733 ( .A(y[521]), .B(x[521]), .Z(n1793) );
  AND U2734 ( .A(n1794), .B(n1793), .Z(n5317) );
  NAND U2735 ( .A(n1795), .B(n5317), .Z(n1798) );
  NANDN U2736 ( .A(x[522]), .B(y[522]), .Z(n1797) );
  NANDN U2737 ( .A(x[521]), .B(y[521]), .Z(n1796) );
  NAND U2738 ( .A(n1797), .B(n1796), .Z(n5320) );
  ANDN U2739 ( .B(n1798), .A(n5320), .Z(n1801) );
  NANDN U2740 ( .A(y[522]), .B(x[522]), .Z(n1800) );
  NANDN U2741 ( .A(y[523]), .B(x[523]), .Z(n1799) );
  AND U2742 ( .A(n1800), .B(n1799), .Z(n5322) );
  NANDN U2743 ( .A(n1801), .B(n5322), .Z(n1802) );
  NANDN U2744 ( .A(n5324), .B(n1802), .Z(n1805) );
  NANDN U2745 ( .A(y[524]), .B(x[524]), .Z(n1804) );
  NANDN U2746 ( .A(y[525]), .B(x[525]), .Z(n1803) );
  AND U2747 ( .A(n1804), .B(n1803), .Z(n5325) );
  NAND U2748 ( .A(n1805), .B(n5325), .Z(n1806) );
  NANDN U2749 ( .A(n5328), .B(n1806), .Z(n1809) );
  NANDN U2750 ( .A(y[526]), .B(x[526]), .Z(n1808) );
  NANDN U2751 ( .A(y[527]), .B(x[527]), .Z(n1807) );
  AND U2752 ( .A(n1808), .B(n1807), .Z(n5329) );
  NAND U2753 ( .A(n1809), .B(n5329), .Z(n1812) );
  NANDN U2754 ( .A(x[528]), .B(y[528]), .Z(n1811) );
  NANDN U2755 ( .A(x[527]), .B(y[527]), .Z(n1810) );
  NAND U2756 ( .A(n1811), .B(n1810), .Z(n5332) );
  ANDN U2757 ( .B(n1812), .A(n5332), .Z(n1815) );
  NANDN U2758 ( .A(y[528]), .B(x[528]), .Z(n1814) );
  NANDN U2759 ( .A(y[529]), .B(x[529]), .Z(n1813) );
  AND U2760 ( .A(n1814), .B(n1813), .Z(n5334) );
  NANDN U2761 ( .A(n1815), .B(n5334), .Z(n1816) );
  NANDN U2762 ( .A(n5336), .B(n1816), .Z(n1819) );
  NANDN U2763 ( .A(y[530]), .B(x[530]), .Z(n1818) );
  NANDN U2764 ( .A(y[531]), .B(x[531]), .Z(n1817) );
  AND U2765 ( .A(n1818), .B(n1817), .Z(n5337) );
  NAND U2766 ( .A(n1819), .B(n5337), .Z(n1820) );
  NANDN U2767 ( .A(n3726), .B(n1820), .Z(n1821) );
  NANDN U2768 ( .A(n3728), .B(n1821), .Z(n1822) );
  AND U2769 ( .A(n5347), .B(n1822), .Z(n1825) );
  NANDN U2770 ( .A(y[534]), .B(x[534]), .Z(n1824) );
  NANDN U2771 ( .A(y[535]), .B(x[535]), .Z(n1823) );
  AND U2772 ( .A(n1824), .B(n1823), .Z(n5349) );
  NANDN U2773 ( .A(n1825), .B(n5349), .Z(n1826) );
  NANDN U2774 ( .A(n5352), .B(n1826), .Z(n1829) );
  NANDN U2775 ( .A(y[536]), .B(x[536]), .Z(n1828) );
  NANDN U2776 ( .A(y[537]), .B(x[537]), .Z(n1827) );
  AND U2777 ( .A(n1828), .B(n1827), .Z(n5353) );
  NAND U2778 ( .A(n1829), .B(n5353), .Z(n1830) );
  NANDN U2779 ( .A(n5356), .B(n1830), .Z(n1833) );
  NANDN U2780 ( .A(y[538]), .B(x[538]), .Z(n1832) );
  NANDN U2781 ( .A(y[539]), .B(x[539]), .Z(n1831) );
  AND U2782 ( .A(n1832), .B(n1831), .Z(n5358) );
  NAND U2783 ( .A(n1833), .B(n5358), .Z(n1836) );
  NANDN U2784 ( .A(x[540]), .B(y[540]), .Z(n1835) );
  NANDN U2785 ( .A(x[539]), .B(y[539]), .Z(n1834) );
  NAND U2786 ( .A(n1835), .B(n1834), .Z(n5360) );
  ANDN U2787 ( .B(n1836), .A(n5360), .Z(n1839) );
  NANDN U2788 ( .A(y[540]), .B(x[540]), .Z(n1838) );
  NANDN U2789 ( .A(y[541]), .B(x[541]), .Z(n1837) );
  AND U2790 ( .A(n1838), .B(n1837), .Z(n5361) );
  NANDN U2791 ( .A(n1839), .B(n5361), .Z(n1840) );
  NANDN U2792 ( .A(n5364), .B(n1840), .Z(n1843) );
  NANDN U2793 ( .A(y[542]), .B(x[542]), .Z(n1842) );
  NANDN U2794 ( .A(y[543]), .B(x[543]), .Z(n1841) );
  AND U2795 ( .A(n1842), .B(n1841), .Z(n5365) );
  NAND U2796 ( .A(n1843), .B(n5365), .Z(n1844) );
  NANDN U2797 ( .A(n5368), .B(n1844), .Z(n1847) );
  NANDN U2798 ( .A(y[544]), .B(x[544]), .Z(n1846) );
  NANDN U2799 ( .A(y[545]), .B(x[545]), .Z(n1845) );
  AND U2800 ( .A(n1846), .B(n1845), .Z(n5370) );
  NAND U2801 ( .A(n1847), .B(n5370), .Z(n1850) );
  NANDN U2802 ( .A(x[546]), .B(y[546]), .Z(n1849) );
  NANDN U2803 ( .A(x[545]), .B(y[545]), .Z(n1848) );
  NAND U2804 ( .A(n1849), .B(n1848), .Z(n5372) );
  ANDN U2805 ( .B(n1850), .A(n5372), .Z(n1853) );
  NANDN U2806 ( .A(y[546]), .B(x[546]), .Z(n1852) );
  NANDN U2807 ( .A(y[547]), .B(x[547]), .Z(n1851) );
  AND U2808 ( .A(n1852), .B(n1851), .Z(n5373) );
  NANDN U2809 ( .A(n1853), .B(n5373), .Z(n1854) );
  NANDN U2810 ( .A(n5376), .B(n1854), .Z(n1857) );
  NANDN U2811 ( .A(y[548]), .B(x[548]), .Z(n1856) );
  NANDN U2812 ( .A(y[549]), .B(x[549]), .Z(n1855) );
  AND U2813 ( .A(n1856), .B(n1855), .Z(n5377) );
  NAND U2814 ( .A(n1857), .B(n5377), .Z(n1858) );
  NANDN U2815 ( .A(n5380), .B(n1858), .Z(n1861) );
  NANDN U2816 ( .A(y[550]), .B(x[550]), .Z(n1860) );
  NANDN U2817 ( .A(y[551]), .B(x[551]), .Z(n1859) );
  AND U2818 ( .A(n1860), .B(n1859), .Z(n5382) );
  NAND U2819 ( .A(n1861), .B(n5382), .Z(n1864) );
  NANDN U2820 ( .A(x[552]), .B(y[552]), .Z(n1863) );
  NANDN U2821 ( .A(x[551]), .B(y[551]), .Z(n1862) );
  NAND U2822 ( .A(n1863), .B(n1862), .Z(n5384) );
  ANDN U2823 ( .B(n1864), .A(n5384), .Z(n1867) );
  NANDN U2824 ( .A(y[552]), .B(x[552]), .Z(n1866) );
  NANDN U2825 ( .A(y[553]), .B(x[553]), .Z(n1865) );
  AND U2826 ( .A(n1866), .B(n1865), .Z(n5386) );
  NANDN U2827 ( .A(n1867), .B(n5386), .Z(n1868) );
  NANDN U2828 ( .A(n5388), .B(n1868), .Z(n1871) );
  NANDN U2829 ( .A(y[555]), .B(x[555]), .Z(n1870) );
  NANDN U2830 ( .A(y[554]), .B(x[554]), .Z(n1869) );
  AND U2831 ( .A(n1870), .B(n1869), .Z(n5389) );
  NAND U2832 ( .A(n1871), .B(n5389), .Z(n1872) );
  NANDN U2833 ( .A(n3752), .B(n1872), .Z(n1873) );
  NANDN U2834 ( .A(n3754), .B(n1873), .Z(n1874) );
  AND U2835 ( .A(n5399), .B(n1874), .Z(n1877) );
  NANDN U2836 ( .A(y[558]), .B(x[558]), .Z(n1876) );
  NANDN U2837 ( .A(y[559]), .B(x[559]), .Z(n1875) );
  AND U2838 ( .A(n1876), .B(n1875), .Z(n5401) );
  NANDN U2839 ( .A(n1877), .B(n5401), .Z(n1878) );
  NANDN U2840 ( .A(n5404), .B(n1878), .Z(n1881) );
  NANDN U2841 ( .A(y[560]), .B(x[560]), .Z(n1880) );
  NANDN U2842 ( .A(y[561]), .B(x[561]), .Z(n1879) );
  AND U2843 ( .A(n1880), .B(n1879), .Z(n5405) );
  NAND U2844 ( .A(n1881), .B(n5405), .Z(n1882) );
  NANDN U2845 ( .A(n5408), .B(n1882), .Z(n1885) );
  NANDN U2846 ( .A(y[562]), .B(x[562]), .Z(n1884) );
  NANDN U2847 ( .A(y[563]), .B(x[563]), .Z(n1883) );
  AND U2848 ( .A(n1884), .B(n1883), .Z(n5410) );
  NAND U2849 ( .A(n1885), .B(n5410), .Z(n1890) );
  NANDN U2850 ( .A(x[564]), .B(y[564]), .Z(n1887) );
  NANDN U2851 ( .A(x[563]), .B(y[563]), .Z(n1886) );
  AND U2852 ( .A(n1887), .B(n1886), .Z(n1889) );
  NANDN U2853 ( .A(x[565]), .B(y[565]), .Z(n1888) );
  NAND U2854 ( .A(n1889), .B(n1888), .Z(n5412) );
  ANDN U2855 ( .B(n1890), .A(n5412), .Z(n1899) );
  NANDN U2856 ( .A(y[567]), .B(x[567]), .Z(n1892) );
  NANDN U2857 ( .A(y[566]), .B(x[566]), .Z(n1891) );
  AND U2858 ( .A(n1892), .B(n1891), .Z(n1898) );
  NANDN U2859 ( .A(y[564]), .B(x[564]), .Z(n1893) );
  NANDN U2860 ( .A(x[565]), .B(n1893), .Z(n1896) );
  XNOR U2861 ( .A(n1893), .B(x[565]), .Z(n1894) );
  NAND U2862 ( .A(n1894), .B(y[565]), .Z(n1895) );
  NAND U2863 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2864 ( .A(n1898), .B(n1897), .Z(n5413) );
  NANDN U2865 ( .A(n1899), .B(n5413), .Z(n1900) );
  NANDN U2866 ( .A(n5416), .B(n1900), .Z(n1901) );
  NAND U2867 ( .A(n1901), .B(n5417), .Z(n1902) );
  NANDN U2868 ( .A(x[570]), .B(y[570]), .Z(n5419) );
  NAND U2869 ( .A(n1902), .B(n5419), .Z(n1905) );
  NANDN U2870 ( .A(y[570]), .B(x[570]), .Z(n1904) );
  NANDN U2871 ( .A(y[571]), .B(x[571]), .Z(n1903) );
  AND U2872 ( .A(n1904), .B(n1903), .Z(n5422) );
  NAND U2873 ( .A(n1905), .B(n5422), .Z(n1908) );
  NANDN U2874 ( .A(x[572]), .B(y[572]), .Z(n1907) );
  NANDN U2875 ( .A(x[571]), .B(y[571]), .Z(n1906) );
  NAND U2876 ( .A(n1907), .B(n1906), .Z(n5424) );
  ANDN U2877 ( .B(n1908), .A(n5424), .Z(n1911) );
  NANDN U2878 ( .A(y[572]), .B(x[572]), .Z(n1910) );
  NANDN U2879 ( .A(y[573]), .B(x[573]), .Z(n1909) );
  AND U2880 ( .A(n1910), .B(n1909), .Z(n5425) );
  NANDN U2881 ( .A(n1911), .B(n5425), .Z(n1912) );
  NANDN U2882 ( .A(n5428), .B(n1912), .Z(n1915) );
  NANDN U2883 ( .A(y[574]), .B(x[574]), .Z(n1914) );
  NANDN U2884 ( .A(y[575]), .B(x[575]), .Z(n1913) );
  AND U2885 ( .A(n1914), .B(n1913), .Z(n5429) );
  NAND U2886 ( .A(n1915), .B(n5429), .Z(n1916) );
  NANDN U2887 ( .A(n5432), .B(n1916), .Z(n1919) );
  NANDN U2888 ( .A(y[576]), .B(x[576]), .Z(n1918) );
  NANDN U2889 ( .A(y[577]), .B(x[577]), .Z(n1917) );
  AND U2890 ( .A(n1918), .B(n1917), .Z(n5434) );
  NAND U2891 ( .A(n1919), .B(n5434), .Z(n1922) );
  NANDN U2892 ( .A(x[578]), .B(y[578]), .Z(n1921) );
  NANDN U2893 ( .A(x[577]), .B(y[577]), .Z(n1920) );
  NAND U2894 ( .A(n1921), .B(n1920), .Z(n5436) );
  ANDN U2895 ( .B(n1922), .A(n5436), .Z(n1925) );
  NANDN U2896 ( .A(y[578]), .B(x[578]), .Z(n1924) );
  NANDN U2897 ( .A(y[579]), .B(x[579]), .Z(n1923) );
  AND U2898 ( .A(n1924), .B(n1923), .Z(n5437) );
  NANDN U2899 ( .A(n1925), .B(n5437), .Z(n1926) );
  NANDN U2900 ( .A(n5440), .B(n1926), .Z(n1929) );
  NANDN U2901 ( .A(y[580]), .B(x[580]), .Z(n1928) );
  NANDN U2902 ( .A(y[581]), .B(x[581]), .Z(n1927) );
  AND U2903 ( .A(n1928), .B(n1927), .Z(n5441) );
  NAND U2904 ( .A(n1929), .B(n5441), .Z(n1931) );
  NANDN U2905 ( .A(x[582]), .B(y[582]), .Z(n1930) );
  ANDN U2906 ( .B(y[581]), .A(x[581]), .Z(n3777) );
  ANDN U2907 ( .B(n1930), .A(n3777), .Z(n5443) );
  NAND U2908 ( .A(n1931), .B(n5443), .Z(n1932) );
  NANDN U2909 ( .A(n5445), .B(n1932), .Z(n1935) );
  NANDN U2910 ( .A(x[584]), .B(y[584]), .Z(n1934) );
  NANDN U2911 ( .A(x[583]), .B(y[583]), .Z(n1933) );
  NAND U2912 ( .A(n1934), .B(n1933), .Z(n5448) );
  ANDN U2913 ( .B(n1935), .A(n5448), .Z(n1938) );
  NANDN U2914 ( .A(y[584]), .B(x[584]), .Z(n1937) );
  NANDN U2915 ( .A(y[585]), .B(x[585]), .Z(n1936) );
  AND U2916 ( .A(n1937), .B(n1936), .Z(n5450) );
  NANDN U2917 ( .A(n1938), .B(n5450), .Z(n1939) );
  NANDN U2918 ( .A(n5452), .B(n1939), .Z(n1942) );
  NANDN U2919 ( .A(y[586]), .B(x[586]), .Z(n1941) );
  NANDN U2920 ( .A(y[587]), .B(x[587]), .Z(n1940) );
  AND U2921 ( .A(n1941), .B(n1940), .Z(n5453) );
  NAND U2922 ( .A(n1942), .B(n5453), .Z(n1943) );
  NANDN U2923 ( .A(n3788), .B(n1943), .Z(n1944) );
  NANDN U2924 ( .A(n3790), .B(n1944), .Z(n1945) );
  AND U2925 ( .A(n5463), .B(n1945), .Z(n1948) );
  NANDN U2926 ( .A(y[590]), .B(x[590]), .Z(n1947) );
  NANDN U2927 ( .A(y[591]), .B(x[591]), .Z(n1946) );
  AND U2928 ( .A(n1947), .B(n1946), .Z(n5465) );
  NANDN U2929 ( .A(n1948), .B(n5465), .Z(n1949) );
  NANDN U2930 ( .A(n5468), .B(n1949), .Z(n1952) );
  NANDN U2931 ( .A(y[592]), .B(x[592]), .Z(n1951) );
  NANDN U2932 ( .A(y[593]), .B(x[593]), .Z(n1950) );
  AND U2933 ( .A(n1951), .B(n1950), .Z(n5469) );
  NAND U2934 ( .A(n1952), .B(n5469), .Z(n1953) );
  NANDN U2935 ( .A(n5472), .B(n1953), .Z(n1956) );
  NANDN U2936 ( .A(y[594]), .B(x[594]), .Z(n1955) );
  NANDN U2937 ( .A(y[595]), .B(x[595]), .Z(n1954) );
  AND U2938 ( .A(n1955), .B(n1954), .Z(n5473) );
  NAND U2939 ( .A(n1956), .B(n5473), .Z(n1959) );
  NANDN U2940 ( .A(x[596]), .B(y[596]), .Z(n1958) );
  NANDN U2941 ( .A(x[595]), .B(y[595]), .Z(n1957) );
  NAND U2942 ( .A(n1958), .B(n1957), .Z(n5476) );
  ANDN U2943 ( .B(n1959), .A(n5476), .Z(n1962) );
  NANDN U2944 ( .A(y[596]), .B(x[596]), .Z(n1961) );
  NANDN U2945 ( .A(y[597]), .B(x[597]), .Z(n1960) );
  AND U2946 ( .A(n1961), .B(n1960), .Z(n5477) );
  NANDN U2947 ( .A(n1962), .B(n5477), .Z(n1963) );
  NANDN U2948 ( .A(n5479), .B(n1963), .Z(n1966) );
  NANDN U2949 ( .A(y[598]), .B(x[598]), .Z(n1965) );
  NANDN U2950 ( .A(y[599]), .B(x[599]), .Z(n1964) );
  AND U2951 ( .A(n1965), .B(n1964), .Z(n5481) );
  NAND U2952 ( .A(n1966), .B(n5481), .Z(n1967) );
  NANDN U2953 ( .A(n5484), .B(n1967), .Z(n1970) );
  NANDN U2954 ( .A(y[600]), .B(x[600]), .Z(n1969) );
  NANDN U2955 ( .A(y[601]), .B(x[601]), .Z(n1968) );
  AND U2956 ( .A(n1969), .B(n1968), .Z(n5485) );
  NAND U2957 ( .A(n1970), .B(n5485), .Z(n1973) );
  NANDN U2958 ( .A(x[602]), .B(y[602]), .Z(n1972) );
  NANDN U2959 ( .A(x[601]), .B(y[601]), .Z(n1971) );
  NAND U2960 ( .A(n1972), .B(n1971), .Z(n5488) );
  ANDN U2961 ( .B(n1973), .A(n5488), .Z(n1976) );
  NANDN U2962 ( .A(y[603]), .B(x[603]), .Z(n1975) );
  NANDN U2963 ( .A(y[602]), .B(x[602]), .Z(n1974) );
  AND U2964 ( .A(n1975), .B(n1974), .Z(n5489) );
  NANDN U2965 ( .A(n1976), .B(n5489), .Z(n1977) );
  AND U2966 ( .A(n1978), .B(n1977), .Z(n1979) );
  OR U2967 ( .A(n5494), .B(n1979), .Z(n1980) );
  AND U2968 ( .A(n1981), .B(n1980), .Z(n1983) );
  NANDN U2969 ( .A(y[606]), .B(x[606]), .Z(n1982) );
  NANDN U2970 ( .A(y[607]), .B(x[607]), .Z(n2939) );
  AND U2971 ( .A(n1982), .B(n2939), .Z(n5497) );
  NANDN U2972 ( .A(n1983), .B(n5497), .Z(n1984) );
  NANDN U2973 ( .A(n2942), .B(n1984), .Z(n1987) );
  NANDN U2974 ( .A(y[608]), .B(x[608]), .Z(n1986) );
  NANDN U2975 ( .A(y[609]), .B(x[609]), .Z(n1985) );
  AND U2976 ( .A(n1986), .B(n1985), .Z(n5501) );
  NAND U2977 ( .A(n1987), .B(n5501), .Z(n1988) );
  NANDN U2978 ( .A(n5503), .B(n1988), .Z(n1991) );
  NANDN U2979 ( .A(y[611]), .B(x[611]), .Z(n1990) );
  NANDN U2980 ( .A(y[610]), .B(x[610]), .Z(n1989) );
  AND U2981 ( .A(n1990), .B(n1989), .Z(n5505) );
  NAND U2982 ( .A(n1991), .B(n5505), .Z(n1992) );
  AND U2983 ( .A(n2936), .B(n1992), .Z(n1993) );
  NANDN U2984 ( .A(x[611]), .B(y[611]), .Z(n5507) );
  NAND U2985 ( .A(n1993), .B(n5507), .Z(n1995) );
  NANDN U2986 ( .A(y[612]), .B(x[612]), .Z(n1994) );
  NANDN U2987 ( .A(y[613]), .B(x[613]), .Z(n2935) );
  AND U2988 ( .A(n1994), .B(n2935), .Z(n5509) );
  NAND U2989 ( .A(n1995), .B(n5509), .Z(n1998) );
  NANDN U2990 ( .A(x[614]), .B(y[614]), .Z(n1997) );
  NANDN U2991 ( .A(x[613]), .B(y[613]), .Z(n1996) );
  NAND U2992 ( .A(n1997), .B(n1996), .Z(n2938) );
  ANDN U2993 ( .B(n1998), .A(n2938), .Z(n2001) );
  NANDN U2994 ( .A(y[614]), .B(x[614]), .Z(n2000) );
  NANDN U2995 ( .A(y[615]), .B(x[615]), .Z(n1999) );
  AND U2996 ( .A(n2000), .B(n1999), .Z(n5513) );
  NANDN U2997 ( .A(n2001), .B(n5513), .Z(n2002) );
  NANDN U2998 ( .A(n5515), .B(n2002), .Z(n2003) );
  NANDN U2999 ( .A(n5518), .B(n2003), .Z(n2004) );
  NANDN U3000 ( .A(x[618]), .B(y[618]), .Z(n5519) );
  NAND U3001 ( .A(n2004), .B(n5519), .Z(n2007) );
  NANDN U3002 ( .A(y[618]), .B(x[618]), .Z(n2006) );
  NANDN U3003 ( .A(y[619]), .B(x[619]), .Z(n2005) );
  AND U3004 ( .A(n2006), .B(n2005), .Z(n5521) );
  NAND U3005 ( .A(n2007), .B(n5521), .Z(n2010) );
  NANDN U3006 ( .A(x[620]), .B(y[620]), .Z(n2009) );
  NANDN U3007 ( .A(x[619]), .B(y[619]), .Z(n2008) );
  NAND U3008 ( .A(n2009), .B(n2008), .Z(n5524) );
  ANDN U3009 ( .B(n2010), .A(n5524), .Z(n2013) );
  NANDN U3010 ( .A(y[620]), .B(x[620]), .Z(n2012) );
  NANDN U3011 ( .A(y[621]), .B(x[621]), .Z(n2011) );
  AND U3012 ( .A(n2012), .B(n2011), .Z(n5525) );
  NANDN U3013 ( .A(n2013), .B(n5525), .Z(n2014) );
  NANDN U3014 ( .A(n5527), .B(n2014), .Z(n2017) );
  NANDN U3015 ( .A(y[623]), .B(x[623]), .Z(n2016) );
  NANDN U3016 ( .A(y[622]), .B(x[622]), .Z(n2015) );
  AND U3017 ( .A(n2016), .B(n2015), .Z(n5529) );
  NAND U3018 ( .A(n2017), .B(n5529), .Z(n2018) );
  NANDN U3019 ( .A(x[623]), .B(y[623]), .Z(n5531) );
  NAND U3020 ( .A(n2018), .B(n5531), .Z(n2020) );
  ANDN U3021 ( .B(y[624]), .A(x[624]), .Z(n2019) );
  OR U3022 ( .A(n2020), .B(n2019), .Z(n2022) );
  NANDN U3023 ( .A(y[624]), .B(x[624]), .Z(n2021) );
  NANDN U3024 ( .A(y[625]), .B(x[625]), .Z(n2929) );
  AND U3025 ( .A(n2021), .B(n2929), .Z(n5533) );
  NAND U3026 ( .A(n2022), .B(n5533), .Z(n2023) );
  NANDN U3027 ( .A(x[625]), .B(y[625]), .Z(n2928) );
  NAND U3028 ( .A(n2023), .B(n2928), .Z(n2024) );
  NANDN U3029 ( .A(x[626]), .B(y[626]), .Z(n2932) );
  NANDN U3030 ( .A(n2024), .B(n2932), .Z(n2027) );
  NANDN U3031 ( .A(y[626]), .B(x[626]), .Z(n2026) );
  NANDN U3032 ( .A(y[627]), .B(x[627]), .Z(n2025) );
  AND U3033 ( .A(n2026), .B(n2025), .Z(n5537) );
  NAND U3034 ( .A(n2027), .B(n5537), .Z(n2029) );
  NANDN U3035 ( .A(x[628]), .B(y[628]), .Z(n2028) );
  ANDN U3036 ( .B(y[627]), .A(x[627]), .Z(n5539) );
  ANDN U3037 ( .B(n2028), .A(n5539), .Z(n3834) );
  NAND U3038 ( .A(n2029), .B(n3834), .Z(n2030) );
  NANDN U3039 ( .A(n3836), .B(n2030), .Z(n2033) );
  NANDN U3040 ( .A(x[630]), .B(y[630]), .Z(n2032) );
  NANDN U3041 ( .A(x[629]), .B(y[629]), .Z(n2031) );
  AND U3042 ( .A(n2032), .B(n2031), .Z(n5545) );
  NAND U3043 ( .A(n2033), .B(n5545), .Z(n2034) );
  AND U3044 ( .A(n5547), .B(n2034), .Z(n2037) );
  NANDN U3045 ( .A(x[632]), .B(y[632]), .Z(n2036) );
  NANDN U3046 ( .A(x[631]), .B(y[631]), .Z(n2035) );
  AND U3047 ( .A(n2036), .B(n2035), .Z(n5550) );
  NANDN U3048 ( .A(n2037), .B(n5550), .Z(n2040) );
  NANDN U3049 ( .A(y[632]), .B(x[632]), .Z(n2039) );
  NANDN U3050 ( .A(y[633]), .B(x[633]), .Z(n2038) );
  AND U3051 ( .A(n2039), .B(n2038), .Z(n5551) );
  NAND U3052 ( .A(n2040), .B(n5551), .Z(n2043) );
  NANDN U3053 ( .A(x[634]), .B(y[634]), .Z(n2042) );
  NANDN U3054 ( .A(x[633]), .B(y[633]), .Z(n2041) );
  AND U3055 ( .A(n2042), .B(n2041), .Z(n5553) );
  NAND U3056 ( .A(n2043), .B(n5553), .Z(n2046) );
  NANDN U3057 ( .A(y[634]), .B(x[634]), .Z(n2045) );
  NANDN U3058 ( .A(y[635]), .B(x[635]), .Z(n2044) );
  AND U3059 ( .A(n2045), .B(n2044), .Z(n5555) );
  NAND U3060 ( .A(n2046), .B(n5555), .Z(n2049) );
  NANDN U3061 ( .A(x[636]), .B(y[636]), .Z(n2048) );
  NANDN U3062 ( .A(x[635]), .B(y[635]), .Z(n2047) );
  AND U3063 ( .A(n2048), .B(n2047), .Z(n5557) );
  NAND U3064 ( .A(n2049), .B(n5557), .Z(n2050) );
  AND U3065 ( .A(n5559), .B(n2050), .Z(n2053) );
  NANDN U3066 ( .A(x[638]), .B(y[638]), .Z(n2052) );
  NANDN U3067 ( .A(x[637]), .B(y[637]), .Z(n2051) );
  AND U3068 ( .A(n2052), .B(n2051), .Z(n5562) );
  NANDN U3069 ( .A(n2053), .B(n5562), .Z(n2056) );
  NANDN U3070 ( .A(y[638]), .B(x[638]), .Z(n2055) );
  NANDN U3071 ( .A(y[639]), .B(x[639]), .Z(n2054) );
  AND U3072 ( .A(n2055), .B(n2054), .Z(n5563) );
  NAND U3073 ( .A(n2056), .B(n5563), .Z(n2059) );
  NANDN U3074 ( .A(x[640]), .B(y[640]), .Z(n2058) );
  NANDN U3075 ( .A(x[639]), .B(y[639]), .Z(n2057) );
  AND U3076 ( .A(n2058), .B(n2057), .Z(n5565) );
  NAND U3077 ( .A(n2059), .B(n5565), .Z(n2062) );
  NANDN U3078 ( .A(y[640]), .B(x[640]), .Z(n2061) );
  NANDN U3079 ( .A(y[641]), .B(x[641]), .Z(n2060) );
  AND U3080 ( .A(n2061), .B(n2060), .Z(n5567) );
  NAND U3081 ( .A(n2062), .B(n5567), .Z(n2065) );
  NANDN U3082 ( .A(x[642]), .B(y[642]), .Z(n2064) );
  NANDN U3083 ( .A(x[641]), .B(y[641]), .Z(n2063) );
  AND U3084 ( .A(n2064), .B(n2063), .Z(n5569) );
  NAND U3085 ( .A(n2065), .B(n5569), .Z(n2066) );
  AND U3086 ( .A(n5571), .B(n2066), .Z(n2068) );
  ANDN U3087 ( .B(y[644]), .A(x[644]), .Z(n2925) );
  NANDN U3088 ( .A(x[645]), .B(y[645]), .Z(n2069) );
  NANDN U3089 ( .A(x[643]), .B(y[643]), .Z(n2067) );
  NAND U3090 ( .A(n2069), .B(n2067), .Z(n3852) );
  NOR U3091 ( .A(n2925), .B(n3852), .Z(n5574) );
  NANDN U3092 ( .A(n2068), .B(n5574), .Z(n2072) );
  ANDN U3093 ( .B(n2069), .A(y[644]), .Z(n2070) );
  NAND U3094 ( .A(n2070), .B(x[644]), .Z(n2071) );
  ANDN U3095 ( .B(x[645]), .A(y[645]), .Z(n2926) );
  ANDN U3096 ( .B(n2071), .A(n2926), .Z(n5575) );
  NAND U3097 ( .A(n2072), .B(n5575), .Z(n2073) );
  NANDN U3098 ( .A(x[646]), .B(y[646]), .Z(n5577) );
  NAND U3099 ( .A(n2073), .B(n5577), .Z(n2076) );
  NANDN U3100 ( .A(y[646]), .B(x[646]), .Z(n2075) );
  NANDN U3101 ( .A(y[647]), .B(x[647]), .Z(n2074) );
  AND U3102 ( .A(n2075), .B(n2074), .Z(n5579) );
  NAND U3103 ( .A(n2076), .B(n5579), .Z(n2079) );
  NANDN U3104 ( .A(x[648]), .B(y[648]), .Z(n2078) );
  NANDN U3105 ( .A(x[647]), .B(y[647]), .Z(n2077) );
  AND U3106 ( .A(n2078), .B(n2077), .Z(n5581) );
  NAND U3107 ( .A(n2079), .B(n5581), .Z(n2080) );
  AND U3108 ( .A(n5583), .B(n2080), .Z(n2083) );
  NANDN U3109 ( .A(x[650]), .B(y[650]), .Z(n2082) );
  NANDN U3110 ( .A(x[649]), .B(y[649]), .Z(n2081) );
  AND U3111 ( .A(n2082), .B(n2081), .Z(n5586) );
  NANDN U3112 ( .A(n2083), .B(n5586), .Z(n2086) );
  NANDN U3113 ( .A(y[650]), .B(x[650]), .Z(n2085) );
  NANDN U3114 ( .A(y[651]), .B(x[651]), .Z(n2084) );
  AND U3115 ( .A(n2085), .B(n2084), .Z(n5587) );
  NAND U3116 ( .A(n2086), .B(n5587), .Z(n2089) );
  NANDN U3117 ( .A(x[652]), .B(y[652]), .Z(n2088) );
  NANDN U3118 ( .A(x[651]), .B(y[651]), .Z(n2087) );
  AND U3119 ( .A(n2088), .B(n2087), .Z(n5589) );
  NAND U3120 ( .A(n2089), .B(n5589), .Z(n2092) );
  NANDN U3121 ( .A(y[652]), .B(x[652]), .Z(n2091) );
  NANDN U3122 ( .A(y[653]), .B(x[653]), .Z(n2090) );
  AND U3123 ( .A(n2091), .B(n2090), .Z(n5591) );
  NAND U3124 ( .A(n2092), .B(n5591), .Z(n2095) );
  NANDN U3125 ( .A(x[654]), .B(y[654]), .Z(n2094) );
  NANDN U3126 ( .A(x[653]), .B(y[653]), .Z(n2093) );
  AND U3127 ( .A(n2094), .B(n2093), .Z(n5593) );
  NAND U3128 ( .A(n2095), .B(n5593), .Z(n2096) );
  AND U3129 ( .A(n5595), .B(n2096), .Z(n2099) );
  NANDN U3130 ( .A(x[656]), .B(y[656]), .Z(n2098) );
  NANDN U3131 ( .A(x[655]), .B(y[655]), .Z(n2097) );
  AND U3132 ( .A(n2098), .B(n2097), .Z(n5598) );
  NANDN U3133 ( .A(n2099), .B(n5598), .Z(n2102) );
  NANDN U3134 ( .A(y[656]), .B(x[656]), .Z(n2101) );
  NANDN U3135 ( .A(y[657]), .B(x[657]), .Z(n2100) );
  AND U3136 ( .A(n2101), .B(n2100), .Z(n5599) );
  NAND U3137 ( .A(n2102), .B(n5599), .Z(n2105) );
  NANDN U3138 ( .A(x[658]), .B(y[658]), .Z(n2104) );
  NANDN U3139 ( .A(x[657]), .B(y[657]), .Z(n2103) );
  AND U3140 ( .A(n2104), .B(n2103), .Z(n5601) );
  NAND U3141 ( .A(n2105), .B(n5601), .Z(n2108) );
  NANDN U3142 ( .A(y[658]), .B(x[658]), .Z(n2107) );
  NANDN U3143 ( .A(y[659]), .B(x[659]), .Z(n2106) );
  AND U3144 ( .A(n2107), .B(n2106), .Z(n5603) );
  NAND U3145 ( .A(n2108), .B(n5603), .Z(n2111) );
  NANDN U3146 ( .A(x[660]), .B(y[660]), .Z(n2110) );
  NANDN U3147 ( .A(x[659]), .B(y[659]), .Z(n2109) );
  AND U3148 ( .A(n2110), .B(n2109), .Z(n5605) );
  NAND U3149 ( .A(n2111), .B(n5605), .Z(n2112) );
  AND U3150 ( .A(n5607), .B(n2112), .Z(n2115) );
  NANDN U3151 ( .A(x[662]), .B(y[662]), .Z(n2114) );
  NANDN U3152 ( .A(x[661]), .B(y[661]), .Z(n2113) );
  AND U3153 ( .A(n2114), .B(n2113), .Z(n5610) );
  NANDN U3154 ( .A(n2115), .B(n5610), .Z(n2118) );
  NANDN U3155 ( .A(y[662]), .B(x[662]), .Z(n2117) );
  NANDN U3156 ( .A(y[663]), .B(x[663]), .Z(n2116) );
  AND U3157 ( .A(n2117), .B(n2116), .Z(n5611) );
  NAND U3158 ( .A(n2118), .B(n5611), .Z(n2121) );
  NANDN U3159 ( .A(x[664]), .B(y[664]), .Z(n2120) );
  NANDN U3160 ( .A(x[663]), .B(y[663]), .Z(n2119) );
  AND U3161 ( .A(n2120), .B(n2119), .Z(n5613) );
  NAND U3162 ( .A(n2121), .B(n5613), .Z(n2124) );
  NANDN U3163 ( .A(y[664]), .B(x[664]), .Z(n2123) );
  NANDN U3164 ( .A(y[665]), .B(x[665]), .Z(n2122) );
  AND U3165 ( .A(n2123), .B(n2122), .Z(n5615) );
  NAND U3166 ( .A(n2124), .B(n5615), .Z(n2127) );
  NANDN U3167 ( .A(x[666]), .B(y[666]), .Z(n2126) );
  NANDN U3168 ( .A(x[665]), .B(y[665]), .Z(n2125) );
  AND U3169 ( .A(n2126), .B(n2125), .Z(n5617) );
  NAND U3170 ( .A(n2127), .B(n5617), .Z(n2128) );
  AND U3171 ( .A(n5619), .B(n2128), .Z(n2131) );
  NANDN U3172 ( .A(x[668]), .B(y[668]), .Z(n2130) );
  NANDN U3173 ( .A(x[667]), .B(y[667]), .Z(n2129) );
  AND U3174 ( .A(n2130), .B(n2129), .Z(n5622) );
  NANDN U3175 ( .A(n2131), .B(n5622), .Z(n2134) );
  NANDN U3176 ( .A(y[668]), .B(x[668]), .Z(n2133) );
  NANDN U3177 ( .A(y[669]), .B(x[669]), .Z(n2132) );
  AND U3178 ( .A(n2133), .B(n2132), .Z(n5623) );
  NAND U3179 ( .A(n2134), .B(n5623), .Z(n2137) );
  NANDN U3180 ( .A(x[670]), .B(y[670]), .Z(n2136) );
  NANDN U3181 ( .A(x[669]), .B(y[669]), .Z(n2135) );
  AND U3182 ( .A(n2136), .B(n2135), .Z(n5625) );
  NAND U3183 ( .A(n2137), .B(n5625), .Z(n2140) );
  NANDN U3184 ( .A(y[670]), .B(x[670]), .Z(n2139) );
  NANDN U3185 ( .A(y[671]), .B(x[671]), .Z(n2138) );
  AND U3186 ( .A(n2139), .B(n2138), .Z(n5627) );
  NAND U3187 ( .A(n2140), .B(n5627), .Z(n2143) );
  NANDN U3188 ( .A(x[672]), .B(y[672]), .Z(n2142) );
  NANDN U3189 ( .A(x[671]), .B(y[671]), .Z(n2141) );
  AND U3190 ( .A(n2142), .B(n2141), .Z(n5629) );
  NAND U3191 ( .A(n2143), .B(n5629), .Z(n2144) );
  AND U3192 ( .A(n5631), .B(n2144), .Z(n2147) );
  NANDN U3193 ( .A(x[674]), .B(y[674]), .Z(n2146) );
  NANDN U3194 ( .A(x[673]), .B(y[673]), .Z(n2145) );
  AND U3195 ( .A(n2146), .B(n2145), .Z(n5634) );
  NANDN U3196 ( .A(n2147), .B(n5634), .Z(n2150) );
  NANDN U3197 ( .A(y[674]), .B(x[674]), .Z(n2149) );
  NANDN U3198 ( .A(y[675]), .B(x[675]), .Z(n2148) );
  AND U3199 ( .A(n2149), .B(n2148), .Z(n5635) );
  NAND U3200 ( .A(n2150), .B(n5635), .Z(n2152) );
  ANDN U3201 ( .B(y[675]), .A(x[675]), .Z(n3887) );
  NOR U3202 ( .A(n3887), .B(n3891), .Z(n5637) );
  NAND U3203 ( .A(n2152), .B(n5637), .Z(n2153) );
  NANDN U3204 ( .A(n5640), .B(n2153), .Z(n2154) );
  NANDN U3205 ( .A(x[678]), .B(y[678]), .Z(n5641) );
  NAND U3206 ( .A(n2154), .B(n5641), .Z(n2155) );
  AND U3207 ( .A(n5643), .B(n2155), .Z(n2158) );
  NANDN U3208 ( .A(x[680]), .B(y[680]), .Z(n2157) );
  NANDN U3209 ( .A(x[679]), .B(y[679]), .Z(n2156) );
  AND U3210 ( .A(n2157), .B(n2156), .Z(n5645) );
  NANDN U3211 ( .A(n2158), .B(n5645), .Z(n2161) );
  NANDN U3212 ( .A(y[680]), .B(x[680]), .Z(n2160) );
  NANDN U3213 ( .A(y[681]), .B(x[681]), .Z(n2159) );
  AND U3214 ( .A(n2160), .B(n2159), .Z(n5647) );
  NAND U3215 ( .A(n2161), .B(n5647), .Z(n2164) );
  NANDN U3216 ( .A(x[682]), .B(y[682]), .Z(n2163) );
  NANDN U3217 ( .A(x[681]), .B(y[681]), .Z(n2162) );
  AND U3218 ( .A(n2163), .B(n2162), .Z(n5649) );
  NAND U3219 ( .A(n2164), .B(n5649), .Z(n2167) );
  NANDN U3220 ( .A(y[682]), .B(x[682]), .Z(n2166) );
  NANDN U3221 ( .A(y[683]), .B(x[683]), .Z(n2165) );
  AND U3222 ( .A(n2166), .B(n2165), .Z(n5652) );
  NAND U3223 ( .A(n2167), .B(n5652), .Z(n2170) );
  NANDN U3224 ( .A(x[684]), .B(y[684]), .Z(n2169) );
  NANDN U3225 ( .A(x[683]), .B(y[683]), .Z(n2168) );
  AND U3226 ( .A(n2169), .B(n2168), .Z(n5653) );
  NAND U3227 ( .A(n2170), .B(n5653), .Z(n2171) );
  AND U3228 ( .A(n5655), .B(n2171), .Z(n2174) );
  NANDN U3229 ( .A(x[686]), .B(y[686]), .Z(n2173) );
  NANDN U3230 ( .A(x[685]), .B(y[685]), .Z(n2172) );
  AND U3231 ( .A(n2173), .B(n2172), .Z(n5657) );
  NANDN U3232 ( .A(n2174), .B(n5657), .Z(n2177) );
  NANDN U3233 ( .A(y[686]), .B(x[686]), .Z(n2176) );
  NANDN U3234 ( .A(y[687]), .B(x[687]), .Z(n2175) );
  AND U3235 ( .A(n2176), .B(n2175), .Z(n5659) );
  NAND U3236 ( .A(n2177), .B(n5659), .Z(n2180) );
  NANDN U3237 ( .A(x[688]), .B(y[688]), .Z(n2179) );
  NANDN U3238 ( .A(x[687]), .B(y[687]), .Z(n2178) );
  AND U3239 ( .A(n2179), .B(n2178), .Z(n5661) );
  NAND U3240 ( .A(n2180), .B(n5661), .Z(n2183) );
  NANDN U3241 ( .A(y[688]), .B(x[688]), .Z(n2182) );
  NANDN U3242 ( .A(y[689]), .B(x[689]), .Z(n2181) );
  AND U3243 ( .A(n2182), .B(n2181), .Z(n5664) );
  NAND U3244 ( .A(n2183), .B(n5664), .Z(n2186) );
  NANDN U3245 ( .A(x[690]), .B(y[690]), .Z(n2185) );
  NANDN U3246 ( .A(x[689]), .B(y[689]), .Z(n2184) );
  AND U3247 ( .A(n2185), .B(n2184), .Z(n5665) );
  NAND U3248 ( .A(n2186), .B(n5665), .Z(n2187) );
  AND U3249 ( .A(n5667), .B(n2187), .Z(n2190) );
  NANDN U3250 ( .A(x[692]), .B(y[692]), .Z(n2189) );
  NANDN U3251 ( .A(x[691]), .B(y[691]), .Z(n2188) );
  AND U3252 ( .A(n2189), .B(n2188), .Z(n5669) );
  NANDN U3253 ( .A(n2190), .B(n5669), .Z(n2193) );
  NANDN U3254 ( .A(y[692]), .B(x[692]), .Z(n2192) );
  NANDN U3255 ( .A(y[693]), .B(x[693]), .Z(n2191) );
  AND U3256 ( .A(n2192), .B(n2191), .Z(n5671) );
  NAND U3257 ( .A(n2193), .B(n5671), .Z(n2196) );
  NANDN U3258 ( .A(x[694]), .B(y[694]), .Z(n2195) );
  NANDN U3259 ( .A(x[693]), .B(y[693]), .Z(n2194) );
  AND U3260 ( .A(n2195), .B(n2194), .Z(n5673) );
  NAND U3261 ( .A(n2196), .B(n5673), .Z(n2199) );
  NANDN U3262 ( .A(y[694]), .B(x[694]), .Z(n2198) );
  NANDN U3263 ( .A(y[695]), .B(x[695]), .Z(n2197) );
  AND U3264 ( .A(n2198), .B(n2197), .Z(n5676) );
  NAND U3265 ( .A(n2199), .B(n5676), .Z(n2201) );
  ANDN U3266 ( .B(y[695]), .A(x[695]), .Z(n3912) );
  NANDN U3267 ( .A(x[696]), .B(y[696]), .Z(n2200) );
  NANDN U3268 ( .A(x[697]), .B(y[697]), .Z(n2204) );
  NAND U3269 ( .A(n2200), .B(n2204), .Z(n3917) );
  NOR U3270 ( .A(n3912), .B(n3917), .Z(n5677) );
  NAND U3271 ( .A(n2201), .B(n5677), .Z(n2205) );
  NANDN U3272 ( .A(y[697]), .B(x[697]), .Z(n3918) );
  NANDN U3273 ( .A(y[696]), .B(x[696]), .Z(n2202) );
  AND U3274 ( .A(n3918), .B(n2202), .Z(n2203) );
  ANDN U3275 ( .B(n2204), .A(n2203), .Z(n5680) );
  ANDN U3276 ( .B(n2205), .A(n5680), .Z(n2206) );
  NANDN U3277 ( .A(x[698]), .B(y[698]), .Z(n5681) );
  NANDN U3278 ( .A(n2206), .B(n5681), .Z(n2209) );
  NANDN U3279 ( .A(y[698]), .B(x[698]), .Z(n2208) );
  NANDN U3280 ( .A(y[699]), .B(x[699]), .Z(n2207) );
  AND U3281 ( .A(n2208), .B(n2207), .Z(n5683) );
  NAND U3282 ( .A(n2209), .B(n5683), .Z(n2212) );
  NANDN U3283 ( .A(x[700]), .B(y[700]), .Z(n2211) );
  NANDN U3284 ( .A(x[699]), .B(y[699]), .Z(n2210) );
  AND U3285 ( .A(n2211), .B(n2210), .Z(n5685) );
  NAND U3286 ( .A(n2212), .B(n5685), .Z(n2215) );
  NANDN U3287 ( .A(y[700]), .B(x[700]), .Z(n2214) );
  NANDN U3288 ( .A(y[701]), .B(x[701]), .Z(n2213) );
  AND U3289 ( .A(n2214), .B(n2213), .Z(n5688) );
  NAND U3290 ( .A(n2215), .B(n5688), .Z(n2218) );
  NANDN U3291 ( .A(x[702]), .B(y[702]), .Z(n2217) );
  NANDN U3292 ( .A(x[701]), .B(y[701]), .Z(n2216) );
  AND U3293 ( .A(n2217), .B(n2216), .Z(n5689) );
  NAND U3294 ( .A(n2218), .B(n5689), .Z(n2219) );
  AND U3295 ( .A(n5691), .B(n2219), .Z(n2222) );
  NANDN U3296 ( .A(x[704]), .B(y[704]), .Z(n2221) );
  NANDN U3297 ( .A(x[703]), .B(y[703]), .Z(n2220) );
  AND U3298 ( .A(n2221), .B(n2220), .Z(n5693) );
  NANDN U3299 ( .A(n2222), .B(n5693), .Z(n2225) );
  NANDN U3300 ( .A(y[704]), .B(x[704]), .Z(n2224) );
  NANDN U3301 ( .A(y[705]), .B(x[705]), .Z(n2223) );
  AND U3302 ( .A(n2224), .B(n2223), .Z(n5695) );
  NAND U3303 ( .A(n2225), .B(n5695), .Z(n2228) );
  NANDN U3304 ( .A(x[706]), .B(y[706]), .Z(n2227) );
  NANDN U3305 ( .A(x[705]), .B(y[705]), .Z(n2226) );
  AND U3306 ( .A(n2227), .B(n2226), .Z(n5697) );
  NAND U3307 ( .A(n2228), .B(n5697), .Z(n2231) );
  NANDN U3308 ( .A(y[706]), .B(x[706]), .Z(n2230) );
  NANDN U3309 ( .A(y[707]), .B(x[707]), .Z(n2229) );
  AND U3310 ( .A(n2230), .B(n2229), .Z(n5700) );
  NAND U3311 ( .A(n2231), .B(n5700), .Z(n2236) );
  NANDN U3312 ( .A(x[708]), .B(y[708]), .Z(n2233) );
  NANDN U3313 ( .A(x[707]), .B(y[707]), .Z(n2232) );
  AND U3314 ( .A(n2233), .B(n2232), .Z(n2235) );
  NANDN U3315 ( .A(x[709]), .B(y[709]), .Z(n2234) );
  AND U3316 ( .A(n2235), .B(n2234), .Z(n5701) );
  NAND U3317 ( .A(n2236), .B(n5701), .Z(n2245) );
  NANDN U3318 ( .A(y[711]), .B(x[711]), .Z(n2238) );
  NANDN U3319 ( .A(y[710]), .B(x[710]), .Z(n2237) );
  AND U3320 ( .A(n2238), .B(n2237), .Z(n2244) );
  NANDN U3321 ( .A(y[708]), .B(x[708]), .Z(n2239) );
  NANDN U3322 ( .A(x[709]), .B(n2239), .Z(n2242) );
  XNOR U3323 ( .A(n2239), .B(x[709]), .Z(n2240) );
  NAND U3324 ( .A(n2240), .B(y[709]), .Z(n2241) );
  NAND U3325 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U3326 ( .A(n2244), .B(n2243), .Z(n5704) );
  ANDN U3327 ( .B(n2245), .A(n5704), .Z(n2246) );
  OR U3328 ( .A(n5706), .B(n2246), .Z(n2249) );
  NANDN U3329 ( .A(y[712]), .B(x[712]), .Z(n2248) );
  NANDN U3330 ( .A(y[713]), .B(x[713]), .Z(n2247) );
  AND U3331 ( .A(n2248), .B(n2247), .Z(n5707) );
  NAND U3332 ( .A(n2249), .B(n5707), .Z(n2252) );
  NANDN U3333 ( .A(x[714]), .B(y[714]), .Z(n2251) );
  NANDN U3334 ( .A(x[713]), .B(y[713]), .Z(n2250) );
  NAND U3335 ( .A(n2251), .B(n2250), .Z(n5710) );
  ANDN U3336 ( .B(n2252), .A(n5710), .Z(n2255) );
  NANDN U3337 ( .A(y[714]), .B(x[714]), .Z(n2254) );
  NANDN U3338 ( .A(y[715]), .B(x[715]), .Z(n2253) );
  AND U3339 ( .A(n2254), .B(n2253), .Z(n5712) );
  NANDN U3340 ( .A(n2255), .B(n5712), .Z(n2256) );
  NANDN U3341 ( .A(n5714), .B(n2256), .Z(n2259) );
  NANDN U3342 ( .A(y[716]), .B(x[716]), .Z(n2258) );
  NANDN U3343 ( .A(y[717]), .B(x[717]), .Z(n2257) );
  AND U3344 ( .A(n2258), .B(n2257), .Z(n5716) );
  NAND U3345 ( .A(n2259), .B(n5716), .Z(n2260) );
  NANDN U3346 ( .A(n5718), .B(n2260), .Z(n2263) );
  NANDN U3347 ( .A(y[718]), .B(x[718]), .Z(n2262) );
  NANDN U3348 ( .A(y[719]), .B(x[719]), .Z(n2261) );
  AND U3349 ( .A(n2262), .B(n2261), .Z(n5719) );
  NAND U3350 ( .A(n2263), .B(n5719), .Z(n2265) );
  ANDN U3351 ( .B(y[719]), .A(x[719]), .Z(n5722) );
  OR U3352 ( .A(n5726), .B(n5722), .Z(n3940) );
  ANDN U3353 ( .B(n2265), .A(n3940), .Z(n2266) );
  OR U3354 ( .A(n3943), .B(n2266), .Z(n2267) );
  NANDN U3355 ( .A(x[722]), .B(y[722]), .Z(n5729) );
  NAND U3356 ( .A(n2267), .B(n5729), .Z(n2270) );
  NANDN U3357 ( .A(y[722]), .B(x[722]), .Z(n2269) );
  NANDN U3358 ( .A(y[723]), .B(x[723]), .Z(n2268) );
  AND U3359 ( .A(n2269), .B(n2268), .Z(n5731) );
  NAND U3360 ( .A(n2270), .B(n5731), .Z(n2271) );
  NANDN U3361 ( .A(n5733), .B(n2271), .Z(n2274) );
  NANDN U3362 ( .A(y[724]), .B(x[724]), .Z(n2273) );
  NANDN U3363 ( .A(y[725]), .B(x[725]), .Z(n2272) );
  AND U3364 ( .A(n2273), .B(n2272), .Z(n5735) );
  NAND U3365 ( .A(n2274), .B(n5735), .Z(n2279) );
  NANDN U3366 ( .A(x[726]), .B(y[726]), .Z(n2276) );
  NANDN U3367 ( .A(x[725]), .B(y[725]), .Z(n2275) );
  AND U3368 ( .A(n2276), .B(n2275), .Z(n2278) );
  NANDN U3369 ( .A(x[727]), .B(y[727]), .Z(n2277) );
  NAND U3370 ( .A(n2278), .B(n2277), .Z(n5738) );
  ANDN U3371 ( .B(n2279), .A(n5738), .Z(n2280) );
  OR U3372 ( .A(n5740), .B(n2280), .Z(n2281) );
  NANDN U3373 ( .A(n5742), .B(n2281), .Z(n2282) );
  NAND U3374 ( .A(n2282), .B(n5743), .Z(n2283) );
  NANDN U3375 ( .A(x[732]), .B(y[732]), .Z(n5746) );
  NAND U3376 ( .A(n2283), .B(n5746), .Z(n2286) );
  NANDN U3377 ( .A(y[732]), .B(x[732]), .Z(n2285) );
  NANDN U3378 ( .A(y[733]), .B(x[733]), .Z(n2284) );
  AND U3379 ( .A(n2285), .B(n2284), .Z(n5747) );
  NAND U3380 ( .A(n2286), .B(n5747), .Z(n2289) );
  NANDN U3381 ( .A(x[734]), .B(y[734]), .Z(n2288) );
  NANDN U3382 ( .A(x[733]), .B(y[733]), .Z(n2287) );
  NAND U3383 ( .A(n2288), .B(n2287), .Z(n5750) );
  ANDN U3384 ( .B(n2289), .A(n5750), .Z(n2292) );
  NANDN U3385 ( .A(y[734]), .B(x[734]), .Z(n2291) );
  NANDN U3386 ( .A(y[735]), .B(x[735]), .Z(n2290) );
  AND U3387 ( .A(n2291), .B(n2290), .Z(n5751) );
  NANDN U3388 ( .A(n2292), .B(n5751), .Z(n2293) );
  NANDN U3389 ( .A(n5754), .B(n2293), .Z(n2296) );
  NANDN U3390 ( .A(y[736]), .B(x[736]), .Z(n2295) );
  NANDN U3391 ( .A(y[737]), .B(x[737]), .Z(n2294) );
  AND U3392 ( .A(n2295), .B(n2294), .Z(n5755) );
  NAND U3393 ( .A(n2296), .B(n5755), .Z(n2297) );
  NANDN U3394 ( .A(n5757), .B(n2297), .Z(n2300) );
  NANDN U3395 ( .A(y[738]), .B(x[738]), .Z(n2299) );
  NANDN U3396 ( .A(y[739]), .B(x[739]), .Z(n2298) );
  AND U3397 ( .A(n2299), .B(n2298), .Z(n5759) );
  NAND U3398 ( .A(n2300), .B(n5759), .Z(n2303) );
  NANDN U3399 ( .A(x[740]), .B(y[740]), .Z(n2302) );
  NANDN U3400 ( .A(x[739]), .B(y[739]), .Z(n2301) );
  NAND U3401 ( .A(n2302), .B(n2301), .Z(n5762) );
  ANDN U3402 ( .B(n2303), .A(n5762), .Z(n2306) );
  NANDN U3403 ( .A(y[740]), .B(x[740]), .Z(n2305) );
  NANDN U3404 ( .A(y[741]), .B(x[741]), .Z(n2304) );
  AND U3405 ( .A(n2305), .B(n2304), .Z(n5763) );
  NANDN U3406 ( .A(n2306), .B(n5763), .Z(n2307) );
  NANDN U3407 ( .A(n5766), .B(n2307), .Z(n2310) );
  NANDN U3408 ( .A(y[742]), .B(x[742]), .Z(n2309) );
  NANDN U3409 ( .A(y[743]), .B(x[743]), .Z(n2308) );
  AND U3410 ( .A(n2309), .B(n2308), .Z(n5767) );
  NAND U3411 ( .A(n2310), .B(n5767), .Z(n2311) );
  NANDN U3412 ( .A(n5769), .B(n2311), .Z(n2314) );
  NANDN U3413 ( .A(y[744]), .B(x[744]), .Z(n2313) );
  NANDN U3414 ( .A(y[745]), .B(x[745]), .Z(n2312) );
  AND U3415 ( .A(n2313), .B(n2312), .Z(n5771) );
  NAND U3416 ( .A(n2314), .B(n5771), .Z(n2316) );
  ANDN U3417 ( .B(y[745]), .A(x[745]), .Z(n5774) );
  OR U3418 ( .A(n5779), .B(n5774), .Z(n3966) );
  ANDN U3419 ( .B(n2316), .A(n3966), .Z(n2317) );
  OR U3420 ( .A(n3969), .B(n2317), .Z(n2318) );
  NANDN U3421 ( .A(x[748]), .B(y[748]), .Z(n5778) );
  NAND U3422 ( .A(n2318), .B(n5778), .Z(n2321) );
  NANDN U3423 ( .A(y[748]), .B(x[748]), .Z(n2320) );
  NANDN U3424 ( .A(y[749]), .B(x[749]), .Z(n2319) );
  AND U3425 ( .A(n2320), .B(n2319), .Z(n5783) );
  NAND U3426 ( .A(n2321), .B(n5783), .Z(n2322) );
  NANDN U3427 ( .A(n5786), .B(n2322), .Z(n2325) );
  NANDN U3428 ( .A(y[750]), .B(x[750]), .Z(n2324) );
  NANDN U3429 ( .A(y[751]), .B(x[751]), .Z(n2323) );
  AND U3430 ( .A(n2324), .B(n2323), .Z(n5787) );
  NAND U3431 ( .A(n2325), .B(n5787), .Z(n2328) );
  NANDN U3432 ( .A(x[752]), .B(y[752]), .Z(n2327) );
  NANDN U3433 ( .A(x[751]), .B(y[751]), .Z(n2326) );
  NAND U3434 ( .A(n2327), .B(n2326), .Z(n5790) );
  ANDN U3435 ( .B(n2328), .A(n5790), .Z(n2331) );
  NANDN U3436 ( .A(y[752]), .B(x[752]), .Z(n2330) );
  NANDN U3437 ( .A(y[753]), .B(x[753]), .Z(n2329) );
  AND U3438 ( .A(n2330), .B(n2329), .Z(n5791) );
  NANDN U3439 ( .A(n2331), .B(n5791), .Z(n2332) );
  NANDN U3440 ( .A(n3977), .B(n2332), .Z(n2333) );
  NANDN U3441 ( .A(n3979), .B(n2333), .Z(n2334) );
  NANDN U3442 ( .A(x[756]), .B(y[756]), .Z(n5801) );
  NAND U3443 ( .A(n2334), .B(n5801), .Z(n2337) );
  NANDN U3444 ( .A(y[757]), .B(x[757]), .Z(n2336) );
  NANDN U3445 ( .A(y[756]), .B(x[756]), .Z(n2335) );
  AND U3446 ( .A(n2336), .B(n2335), .Z(n5803) );
  NAND U3447 ( .A(n2337), .B(n5803), .Z(n2339) );
  ANDN U3448 ( .B(y[757]), .A(x[757]), .Z(n5805) );
  OR U3449 ( .A(n5810), .B(n5805), .Z(n3982) );
  ANDN U3450 ( .B(n2339), .A(n3982), .Z(n2340) );
  OR U3451 ( .A(n3985), .B(n2340), .Z(n2341) );
  NANDN U3452 ( .A(x[760]), .B(y[760]), .Z(n5813) );
  NAND U3453 ( .A(n2341), .B(n5813), .Z(n2344) );
  NANDN U3454 ( .A(y[760]), .B(x[760]), .Z(n2343) );
  NANDN U3455 ( .A(y[761]), .B(x[761]), .Z(n2342) );
  AND U3456 ( .A(n2343), .B(n2342), .Z(n5815) );
  NAND U3457 ( .A(n2344), .B(n5815), .Z(n2345) );
  NANDN U3458 ( .A(n5817), .B(n2345), .Z(n2348) );
  NANDN U3459 ( .A(y[762]), .B(x[762]), .Z(n2347) );
  NANDN U3460 ( .A(y[763]), .B(x[763]), .Z(n2346) );
  AND U3461 ( .A(n2347), .B(n2346), .Z(n5819) );
  NAND U3462 ( .A(n2348), .B(n5819), .Z(n2351) );
  NANDN U3463 ( .A(x[764]), .B(y[764]), .Z(n2350) );
  NANDN U3464 ( .A(x[763]), .B(y[763]), .Z(n2349) );
  NAND U3465 ( .A(n2350), .B(n2349), .Z(n5822) );
  ANDN U3466 ( .B(n2351), .A(n5822), .Z(n2354) );
  NANDN U3467 ( .A(y[764]), .B(x[764]), .Z(n2353) );
  NANDN U3468 ( .A(y[765]), .B(x[765]), .Z(n2352) );
  AND U3469 ( .A(n2353), .B(n2352), .Z(n5823) );
  NANDN U3470 ( .A(n2354), .B(n5823), .Z(n2355) );
  NANDN U3471 ( .A(n5826), .B(n2355), .Z(n2358) );
  NANDN U3472 ( .A(y[766]), .B(x[766]), .Z(n2357) );
  NANDN U3473 ( .A(y[767]), .B(x[767]), .Z(n2356) );
  AND U3474 ( .A(n2357), .B(n2356), .Z(n5827) );
  NAND U3475 ( .A(n2358), .B(n5827), .Z(n2359) );
  NANDN U3476 ( .A(n5829), .B(n2359), .Z(n2362) );
  NANDN U3477 ( .A(y[768]), .B(x[768]), .Z(n2361) );
  NANDN U3478 ( .A(y[769]), .B(x[769]), .Z(n2360) );
  AND U3479 ( .A(n2361), .B(n2360), .Z(n5831) );
  NAND U3480 ( .A(n2362), .B(n5831), .Z(n2367) );
  NANDN U3481 ( .A(x[770]), .B(y[770]), .Z(n2364) );
  NANDN U3482 ( .A(x[769]), .B(y[769]), .Z(n2363) );
  AND U3483 ( .A(n2364), .B(n2363), .Z(n2366) );
  NANDN U3484 ( .A(x[771]), .B(y[771]), .Z(n2365) );
  NAND U3485 ( .A(n2366), .B(n2365), .Z(n5834) );
  ANDN U3486 ( .B(n2367), .A(n5834), .Z(n2368) );
  NANDN U3487 ( .A(n2368), .B(n5835), .Z(n2370) );
  NAND U3488 ( .A(n2370), .B(n5839), .Z(n2371) );
  NANDN U3489 ( .A(n4000), .B(n2371), .Z(n2372) );
  NANDN U3490 ( .A(x[774]), .B(y[774]), .Z(n5843) );
  NAND U3491 ( .A(n2372), .B(n5843), .Z(n2375) );
  NANDN U3492 ( .A(y[774]), .B(x[774]), .Z(n2374) );
  NANDN U3493 ( .A(y[775]), .B(x[775]), .Z(n2373) );
  AND U3494 ( .A(n2374), .B(n2373), .Z(n5845) );
  NAND U3495 ( .A(n2375), .B(n5845), .Z(n2378) );
  NANDN U3496 ( .A(x[776]), .B(y[776]), .Z(n2377) );
  NANDN U3497 ( .A(x[775]), .B(y[775]), .Z(n2376) );
  NAND U3498 ( .A(n2377), .B(n2376), .Z(n5847) );
  ANDN U3499 ( .B(n2378), .A(n5847), .Z(n2381) );
  NANDN U3500 ( .A(y[776]), .B(x[776]), .Z(n2380) );
  NANDN U3501 ( .A(y[777]), .B(x[777]), .Z(n2379) );
  AND U3502 ( .A(n2380), .B(n2379), .Z(n5849) );
  NANDN U3503 ( .A(n2381), .B(n5849), .Z(n2382) );
  NANDN U3504 ( .A(n5852), .B(n2382), .Z(n2385) );
  NANDN U3505 ( .A(y[778]), .B(x[778]), .Z(n2384) );
  NANDN U3506 ( .A(y[779]), .B(x[779]), .Z(n2383) );
  AND U3507 ( .A(n2384), .B(n2383), .Z(n5853) );
  NAND U3508 ( .A(n2385), .B(n5853), .Z(n2386) );
  NANDN U3509 ( .A(n5856), .B(n2386), .Z(n2387) );
  NAND U3510 ( .A(n2387), .B(n5859), .Z(n2388) );
  AND U3511 ( .A(n5861), .B(n2388), .Z(n2389) );
  OR U3512 ( .A(n4011), .B(n2389), .Z(n2390) );
  NANDN U3513 ( .A(x[784]), .B(y[784]), .Z(n5865) );
  NAND U3514 ( .A(n2390), .B(n5865), .Z(n2393) );
  NANDN U3515 ( .A(y[784]), .B(x[784]), .Z(n2392) );
  NANDN U3516 ( .A(y[785]), .B(x[785]), .Z(n2391) );
  AND U3517 ( .A(n2392), .B(n2391), .Z(n5867) );
  NAND U3518 ( .A(n2393), .B(n5867), .Z(n2394) );
  NANDN U3519 ( .A(n5870), .B(n2394), .Z(n2397) );
  NANDN U3520 ( .A(y[786]), .B(x[786]), .Z(n2396) );
  NANDN U3521 ( .A(y[787]), .B(x[787]), .Z(n2395) );
  AND U3522 ( .A(n2396), .B(n2395), .Z(n5872) );
  NAND U3523 ( .A(n2397), .B(n5872), .Z(n2400) );
  NANDN U3524 ( .A(x[788]), .B(y[788]), .Z(n2399) );
  NANDN U3525 ( .A(x[787]), .B(y[787]), .Z(n2398) );
  NAND U3526 ( .A(n2399), .B(n2398), .Z(n5874) );
  ANDN U3527 ( .B(n2400), .A(n5874), .Z(n2403) );
  NANDN U3528 ( .A(y[788]), .B(x[788]), .Z(n2402) );
  NANDN U3529 ( .A(y[789]), .B(x[789]), .Z(n2401) );
  AND U3530 ( .A(n2402), .B(n2401), .Z(n5875) );
  NANDN U3531 ( .A(n2403), .B(n5875), .Z(n2404) );
  NANDN U3532 ( .A(n5878), .B(n2404), .Z(n2407) );
  NANDN U3533 ( .A(y[790]), .B(x[790]), .Z(n2406) );
  NANDN U3534 ( .A(y[791]), .B(x[791]), .Z(n2405) );
  AND U3535 ( .A(n2406), .B(n2405), .Z(n5879) );
  NAND U3536 ( .A(n2407), .B(n5879), .Z(n2408) );
  NANDN U3537 ( .A(n5882), .B(n2408), .Z(n2411) );
  NANDN U3538 ( .A(y[792]), .B(x[792]), .Z(n2410) );
  NANDN U3539 ( .A(y[793]), .B(x[793]), .Z(n2409) );
  AND U3540 ( .A(n2410), .B(n2409), .Z(n5884) );
  NAND U3541 ( .A(n2411), .B(n5884), .Z(n2414) );
  NANDN U3542 ( .A(x[794]), .B(y[794]), .Z(n2413) );
  NANDN U3543 ( .A(x[793]), .B(y[793]), .Z(n2412) );
  NAND U3544 ( .A(n2413), .B(n2412), .Z(n5886) );
  ANDN U3545 ( .B(n2414), .A(n5886), .Z(n2417) );
  NANDN U3546 ( .A(y[794]), .B(x[794]), .Z(n2416) );
  NANDN U3547 ( .A(y[795]), .B(x[795]), .Z(n2415) );
  AND U3548 ( .A(n2416), .B(n2415), .Z(n5887) );
  NANDN U3549 ( .A(n2417), .B(n5887), .Z(n2418) );
  NANDN U3550 ( .A(n5890), .B(n2418), .Z(n2421) );
  NANDN U3551 ( .A(y[796]), .B(x[796]), .Z(n2420) );
  NANDN U3552 ( .A(y[797]), .B(x[797]), .Z(n2419) );
  AND U3553 ( .A(n2420), .B(n2419), .Z(n5891) );
  NAND U3554 ( .A(n2421), .B(n5891), .Z(n2422) );
  NANDN U3555 ( .A(n5894), .B(n2422), .Z(n2425) );
  NANDN U3556 ( .A(y[798]), .B(x[798]), .Z(n2424) );
  NANDN U3557 ( .A(y[799]), .B(x[799]), .Z(n2423) );
  AND U3558 ( .A(n2424), .B(n2423), .Z(n5896) );
  NAND U3559 ( .A(n2425), .B(n5896), .Z(n2428) );
  NANDN U3560 ( .A(x[800]), .B(y[800]), .Z(n2427) );
  NANDN U3561 ( .A(x[799]), .B(y[799]), .Z(n2426) );
  NAND U3562 ( .A(n2427), .B(n2426), .Z(n5898) );
  ANDN U3563 ( .B(n2428), .A(n5898), .Z(n2431) );
  NANDN U3564 ( .A(y[800]), .B(x[800]), .Z(n2430) );
  NANDN U3565 ( .A(y[801]), .B(x[801]), .Z(n2429) );
  AND U3566 ( .A(n2430), .B(n2429), .Z(n5899) );
  NANDN U3567 ( .A(n2431), .B(n5899), .Z(n2432) );
  ANDN U3568 ( .B(y[801]), .A(x[801]), .Z(n4031) );
  NANDN U3569 ( .A(x[803]), .B(y[803]), .Z(n2434) );
  NOR U3570 ( .A(n4031), .B(n4035), .Z(n5901) );
  NAND U3571 ( .A(n2432), .B(n5901), .Z(n2435) );
  ANDN U3572 ( .B(x[803]), .A(y[803]), .Z(n4036) );
  NANDN U3573 ( .A(y[802]), .B(x[802]), .Z(n2433) );
  NANDN U3574 ( .A(n4036), .B(n2433), .Z(n4033) );
  NAND U3575 ( .A(n2434), .B(n4033), .Z(n5903) );
  NAND U3576 ( .A(n2435), .B(n5903), .Z(n2436) );
  NANDN U3577 ( .A(x[804]), .B(y[804]), .Z(n5905) );
  NAND U3578 ( .A(n2436), .B(n5905), .Z(n2439) );
  NANDN U3579 ( .A(y[804]), .B(x[804]), .Z(n2438) );
  NANDN U3580 ( .A(y[805]), .B(x[805]), .Z(n2437) );
  AND U3581 ( .A(n2438), .B(n2437), .Z(n5908) );
  NAND U3582 ( .A(n2439), .B(n5908), .Z(n2441) );
  ANDN U3583 ( .B(y[805]), .A(x[805]), .Z(n5910) );
  OR U3584 ( .A(n5916), .B(n5910), .Z(n4041) );
  ANDN U3585 ( .B(n2441), .A(n4041), .Z(n2442) );
  OR U3586 ( .A(n4043), .B(n2442), .Z(n2444) );
  NAND U3587 ( .A(n2444), .B(n5913), .Z(n2445) );
  NANDN U3588 ( .A(n5920), .B(n2445), .Z(n2446) );
  NANDN U3589 ( .A(x[810]), .B(y[810]), .Z(n5921) );
  NAND U3590 ( .A(n2446), .B(n5921), .Z(n2449) );
  NANDN U3591 ( .A(y[810]), .B(x[810]), .Z(n2448) );
  NANDN U3592 ( .A(y[811]), .B(x[811]), .Z(n2447) );
  AND U3593 ( .A(n2448), .B(n2447), .Z(n5923) );
  NAND U3594 ( .A(n2449), .B(n5923), .Z(n2452) );
  NANDN U3595 ( .A(x[812]), .B(y[812]), .Z(n2451) );
  NANDN U3596 ( .A(x[811]), .B(y[811]), .Z(n2450) );
  AND U3597 ( .A(n2451), .B(n2450), .Z(n5926) );
  NAND U3598 ( .A(n2452), .B(n5926), .Z(n2455) );
  NANDN U3599 ( .A(y[812]), .B(x[812]), .Z(n2454) );
  NANDN U3600 ( .A(y[813]), .B(x[813]), .Z(n2453) );
  AND U3601 ( .A(n2454), .B(n2453), .Z(n5927) );
  NAND U3602 ( .A(n2455), .B(n5927), .Z(n2458) );
  NANDN U3603 ( .A(x[814]), .B(y[814]), .Z(n2457) );
  NANDN U3604 ( .A(x[813]), .B(y[813]), .Z(n2456) );
  AND U3605 ( .A(n2457), .B(n2456), .Z(n5929) );
  NAND U3606 ( .A(n2458), .B(n5929), .Z(n2459) );
  AND U3607 ( .A(n5931), .B(n2459), .Z(n2462) );
  NANDN U3608 ( .A(x[816]), .B(y[816]), .Z(n2461) );
  NANDN U3609 ( .A(x[815]), .B(y[815]), .Z(n2460) );
  AND U3610 ( .A(n2461), .B(n2460), .Z(n5933) );
  NANDN U3611 ( .A(n2462), .B(n5933), .Z(n2465) );
  NANDN U3612 ( .A(y[816]), .B(x[816]), .Z(n2464) );
  NANDN U3613 ( .A(y[817]), .B(x[817]), .Z(n2463) );
  AND U3614 ( .A(n2464), .B(n2463), .Z(n5935) );
  NAND U3615 ( .A(n2465), .B(n5935), .Z(n2468) );
  NANDN U3616 ( .A(x[818]), .B(y[818]), .Z(n2467) );
  NANDN U3617 ( .A(x[817]), .B(y[817]), .Z(n2466) );
  AND U3618 ( .A(n2467), .B(n2466), .Z(n5938) );
  NAND U3619 ( .A(n2468), .B(n5938), .Z(n2471) );
  NANDN U3620 ( .A(y[818]), .B(x[818]), .Z(n2470) );
  NANDN U3621 ( .A(y[819]), .B(x[819]), .Z(n2469) );
  AND U3622 ( .A(n2470), .B(n2469), .Z(n5939) );
  NAND U3623 ( .A(n2471), .B(n5939), .Z(n2474) );
  NANDN U3624 ( .A(x[820]), .B(y[820]), .Z(n2473) );
  NANDN U3625 ( .A(x[819]), .B(y[819]), .Z(n2472) );
  AND U3626 ( .A(n2473), .B(n2472), .Z(n5941) );
  NAND U3627 ( .A(n2474), .B(n5941), .Z(n2475) );
  AND U3628 ( .A(n5943), .B(n2475), .Z(n2478) );
  NANDN U3629 ( .A(x[822]), .B(y[822]), .Z(n2477) );
  NANDN U3630 ( .A(x[821]), .B(y[821]), .Z(n2476) );
  AND U3631 ( .A(n2477), .B(n2476), .Z(n5945) );
  NANDN U3632 ( .A(n2478), .B(n5945), .Z(n2481) );
  NANDN U3633 ( .A(y[822]), .B(x[822]), .Z(n2480) );
  NANDN U3634 ( .A(y[823]), .B(x[823]), .Z(n2479) );
  AND U3635 ( .A(n2480), .B(n2479), .Z(n5947) );
  NAND U3636 ( .A(n2481), .B(n5947), .Z(n2484) );
  NANDN U3637 ( .A(x[824]), .B(y[824]), .Z(n2483) );
  NANDN U3638 ( .A(x[823]), .B(y[823]), .Z(n2482) );
  AND U3639 ( .A(n2483), .B(n2482), .Z(n5950) );
  NAND U3640 ( .A(n2484), .B(n5950), .Z(n2487) );
  NANDN U3641 ( .A(y[824]), .B(x[824]), .Z(n2486) );
  NANDN U3642 ( .A(y[825]), .B(x[825]), .Z(n2485) );
  AND U3643 ( .A(n2486), .B(n2485), .Z(n5951) );
  NAND U3644 ( .A(n2487), .B(n5951), .Z(n2490) );
  NANDN U3645 ( .A(x[826]), .B(y[826]), .Z(n2489) );
  NANDN U3646 ( .A(x[825]), .B(y[825]), .Z(n2488) );
  AND U3647 ( .A(n2489), .B(n2488), .Z(n5953) );
  NAND U3648 ( .A(n2490), .B(n5953), .Z(n2491) );
  AND U3649 ( .A(n5955), .B(n2491), .Z(n2494) );
  NANDN U3650 ( .A(x[828]), .B(y[828]), .Z(n2493) );
  NANDN U3651 ( .A(x[827]), .B(y[827]), .Z(n2492) );
  AND U3652 ( .A(n2493), .B(n2492), .Z(n5957) );
  NANDN U3653 ( .A(n2494), .B(n5957), .Z(n2497) );
  NANDN U3654 ( .A(y[828]), .B(x[828]), .Z(n2496) );
  NANDN U3655 ( .A(y[829]), .B(x[829]), .Z(n2495) );
  AND U3656 ( .A(n2496), .B(n2495), .Z(n5959) );
  NAND U3657 ( .A(n2497), .B(n5959), .Z(n2500) );
  NANDN U3658 ( .A(x[830]), .B(y[830]), .Z(n2499) );
  NANDN U3659 ( .A(x[829]), .B(y[829]), .Z(n2498) );
  AND U3660 ( .A(n2499), .B(n2498), .Z(n5962) );
  NAND U3661 ( .A(n2500), .B(n5962), .Z(n2503) );
  NANDN U3662 ( .A(y[830]), .B(x[830]), .Z(n2502) );
  NANDN U3663 ( .A(y[831]), .B(x[831]), .Z(n2501) );
  AND U3664 ( .A(n2502), .B(n2501), .Z(n5963) );
  NAND U3665 ( .A(n2503), .B(n5963), .Z(n2506) );
  NANDN U3666 ( .A(x[832]), .B(y[832]), .Z(n2505) );
  NANDN U3667 ( .A(x[831]), .B(y[831]), .Z(n2504) );
  AND U3668 ( .A(n2505), .B(n2504), .Z(n5965) );
  NAND U3669 ( .A(n2506), .B(n5965), .Z(n2507) );
  AND U3670 ( .A(n5967), .B(n2507), .Z(n2510) );
  NANDN U3671 ( .A(x[834]), .B(y[834]), .Z(n2509) );
  NANDN U3672 ( .A(x[833]), .B(y[833]), .Z(n2508) );
  AND U3673 ( .A(n2509), .B(n2508), .Z(n5969) );
  NANDN U3674 ( .A(n2510), .B(n5969), .Z(n2513) );
  NANDN U3675 ( .A(y[834]), .B(x[834]), .Z(n2512) );
  NANDN U3676 ( .A(y[835]), .B(x[835]), .Z(n2511) );
  AND U3677 ( .A(n2512), .B(n2511), .Z(n5971) );
  NAND U3678 ( .A(n2513), .B(n5971), .Z(n2516) );
  NANDN U3679 ( .A(x[836]), .B(y[836]), .Z(n2515) );
  NANDN U3680 ( .A(x[835]), .B(y[835]), .Z(n2514) );
  AND U3681 ( .A(n2515), .B(n2514), .Z(n5974) );
  NAND U3682 ( .A(n2516), .B(n5974), .Z(n2519) );
  NANDN U3683 ( .A(y[836]), .B(x[836]), .Z(n2518) );
  NANDN U3684 ( .A(y[837]), .B(x[837]), .Z(n2517) );
  AND U3685 ( .A(n2518), .B(n2517), .Z(n5975) );
  NAND U3686 ( .A(n2519), .B(n5975), .Z(n2522) );
  NANDN U3687 ( .A(x[838]), .B(y[838]), .Z(n2521) );
  NANDN U3688 ( .A(x[837]), .B(y[837]), .Z(n2520) );
  AND U3689 ( .A(n2521), .B(n2520), .Z(n5977) );
  NAND U3690 ( .A(n2522), .B(n5977), .Z(n2523) );
  AND U3691 ( .A(n5979), .B(n2523), .Z(n2526) );
  NANDN U3692 ( .A(x[840]), .B(y[840]), .Z(n2525) );
  NANDN U3693 ( .A(x[839]), .B(y[839]), .Z(n2524) );
  AND U3694 ( .A(n2525), .B(n2524), .Z(n5981) );
  NANDN U3695 ( .A(n2526), .B(n5981), .Z(n2529) );
  NANDN U3696 ( .A(y[840]), .B(x[840]), .Z(n2528) );
  NANDN U3697 ( .A(y[841]), .B(x[841]), .Z(n2527) );
  AND U3698 ( .A(n2528), .B(n2527), .Z(n5983) );
  NAND U3699 ( .A(n2529), .B(n5983), .Z(n2532) );
  NANDN U3700 ( .A(x[842]), .B(y[842]), .Z(n2531) );
  NANDN U3701 ( .A(x[841]), .B(y[841]), .Z(n2530) );
  AND U3702 ( .A(n2531), .B(n2530), .Z(n5986) );
  NAND U3703 ( .A(n2532), .B(n5986), .Z(n2535) );
  NANDN U3704 ( .A(y[842]), .B(x[842]), .Z(n2534) );
  NANDN U3705 ( .A(y[843]), .B(x[843]), .Z(n2533) );
  AND U3706 ( .A(n2534), .B(n2533), .Z(n5987) );
  NAND U3707 ( .A(n2535), .B(n5987), .Z(n2538) );
  NANDN U3708 ( .A(x[844]), .B(y[844]), .Z(n2537) );
  NANDN U3709 ( .A(x[843]), .B(y[843]), .Z(n2536) );
  AND U3710 ( .A(n2537), .B(n2536), .Z(n5989) );
  NAND U3711 ( .A(n2538), .B(n5989), .Z(n2539) );
  AND U3712 ( .A(n5991), .B(n2539), .Z(n2542) );
  NANDN U3713 ( .A(x[846]), .B(y[846]), .Z(n2541) );
  NANDN U3714 ( .A(x[845]), .B(y[845]), .Z(n2540) );
  AND U3715 ( .A(n2541), .B(n2540), .Z(n5993) );
  NANDN U3716 ( .A(n2542), .B(n5993), .Z(n2545) );
  NANDN U3717 ( .A(y[846]), .B(x[846]), .Z(n2544) );
  NANDN U3718 ( .A(y[847]), .B(x[847]), .Z(n2543) );
  AND U3719 ( .A(n2544), .B(n2543), .Z(n5995) );
  NAND U3720 ( .A(n2545), .B(n5995), .Z(n2548) );
  NANDN U3721 ( .A(x[847]), .B(y[847]), .Z(n2547) );
  NANDN U3722 ( .A(x[848]), .B(y[848]), .Z(n2546) );
  AND U3723 ( .A(n2547), .B(n2546), .Z(n5998) );
  NAND U3724 ( .A(n2548), .B(n5998), .Z(n2549) );
  NANDN U3725 ( .A(y[848]), .B(x[848]), .Z(n5999) );
  NAND U3726 ( .A(n2549), .B(n5999), .Z(n2550) );
  NANDN U3727 ( .A(x[849]), .B(y[849]), .Z(n6001) );
  NAND U3728 ( .A(n2550), .B(n6001), .Z(n2552) );
  NANDN U3729 ( .A(y[849]), .B(x[849]), .Z(n4089) );
  IV U3730 ( .A(x[850]), .Z(n2924) );
  IV U3731 ( .A(y[850]), .Z(n2923) );
  NANDN U3732 ( .A(n2924), .B(n2923), .Z(n2551) );
  NAND U3733 ( .A(n4089), .B(n2551), .Z(n6004) );
  ANDN U3734 ( .B(n2552), .A(n6004), .Z(n2554) );
  NANDN U3735 ( .A(x[850]), .B(y[850]), .Z(n2553) );
  ANDN U3736 ( .B(y[851]), .A(x[851]), .Z(n2921) );
  ANDN U3737 ( .B(n2553), .A(n2921), .Z(n6005) );
  NANDN U3738 ( .A(n2554), .B(n6005), .Z(n2555) );
  NANDN U3739 ( .A(y[851]), .B(x[851]), .Z(n6007) );
  NAND U3740 ( .A(n2555), .B(n6007), .Z(n2556) );
  NANDN U3741 ( .A(x[852]), .B(y[852]), .Z(n6010) );
  NAND U3742 ( .A(n2556), .B(n6010), .Z(n2559) );
  NANDN U3743 ( .A(y[852]), .B(x[852]), .Z(n2558) );
  NANDN U3744 ( .A(y[853]), .B(x[853]), .Z(n2557) );
  AND U3745 ( .A(n2558), .B(n2557), .Z(n6011) );
  NAND U3746 ( .A(n2559), .B(n6011), .Z(n2562) );
  NANDN U3747 ( .A(x[854]), .B(y[854]), .Z(n2561) );
  NANDN U3748 ( .A(x[853]), .B(y[853]), .Z(n2560) );
  AND U3749 ( .A(n2561), .B(n2560), .Z(n6013) );
  NAND U3750 ( .A(n2562), .B(n6013), .Z(n2563) );
  AND U3751 ( .A(n6015), .B(n2563), .Z(n2566) );
  NANDN U3752 ( .A(x[856]), .B(y[856]), .Z(n2565) );
  NANDN U3753 ( .A(x[855]), .B(y[855]), .Z(n2564) );
  AND U3754 ( .A(n2565), .B(n2564), .Z(n6017) );
  NANDN U3755 ( .A(n2566), .B(n6017), .Z(n2569) );
  NANDN U3756 ( .A(y[856]), .B(x[856]), .Z(n2568) );
  NANDN U3757 ( .A(y[857]), .B(x[857]), .Z(n2567) );
  AND U3758 ( .A(n2568), .B(n2567), .Z(n6019) );
  NAND U3759 ( .A(n2569), .B(n6019), .Z(n2570) );
  NANDN U3760 ( .A(x[857]), .B(y[857]), .Z(n6023) );
  NAND U3761 ( .A(n2570), .B(n6023), .Z(n2571) );
  NANDN U3762 ( .A(n6026), .B(n2571), .Z(n2575) );
  ANDN U3763 ( .B(y[860]), .A(x[860]), .Z(n4362) );
  ANDN U3764 ( .B(y[859]), .A(x[859]), .Z(n6027) );
  NOR U3765 ( .A(n4362), .B(n6027), .Z(n2574) );
  NANDN U3766 ( .A(x[858]), .B(y[858]), .Z(n6022) );
  NANDN U3767 ( .A(n6022), .B(n2572), .Z(n2573) );
  AND U3768 ( .A(n2574), .B(n2573), .Z(n4105) );
  NAND U3769 ( .A(n2575), .B(n4105), .Z(n2576) );
  AND U3770 ( .A(n6029), .B(n2576), .Z(n2577) );
  NANDN U3771 ( .A(x[861]), .B(y[861]), .Z(n4363) );
  NANDN U3772 ( .A(n2577), .B(n4363), .Z(n2578) );
  NANDN U3773 ( .A(n6034), .B(n2578), .Z(n2579) );
  NANDN U3774 ( .A(n6036), .B(n2579), .Z(n2580) );
  NANDN U3775 ( .A(y[863]), .B(x[863]), .Z(n6037) );
  NAND U3776 ( .A(n2580), .B(n6037), .Z(n2581) );
  NANDN U3777 ( .A(x[864]), .B(y[864]), .Z(n6039) );
  NAND U3778 ( .A(n2581), .B(n6039), .Z(n2584) );
  NANDN U3779 ( .A(y[865]), .B(x[865]), .Z(n2583) );
  NANDN U3780 ( .A(y[864]), .B(x[864]), .Z(n2582) );
  NAND U3781 ( .A(n2583), .B(n2582), .Z(n6042) );
  ANDN U3782 ( .B(n2584), .A(n6042), .Z(n2587) );
  NANDN U3783 ( .A(x[865]), .B(y[865]), .Z(n2586) );
  NANDN U3784 ( .A(x[866]), .B(y[866]), .Z(n2585) );
  AND U3785 ( .A(n2586), .B(n2585), .Z(n6044) );
  NANDN U3786 ( .A(n2587), .B(n6044), .Z(n2588) );
  NANDN U3787 ( .A(n6046), .B(n2588), .Z(n2591) );
  NANDN U3788 ( .A(x[867]), .B(y[867]), .Z(n2590) );
  NANDN U3789 ( .A(x[868]), .B(y[868]), .Z(n2589) );
  AND U3790 ( .A(n2590), .B(n2589), .Z(n6047) );
  NAND U3791 ( .A(n2591), .B(n6047), .Z(n2592) );
  NANDN U3792 ( .A(n6050), .B(n2592), .Z(n2593) );
  NANDN U3793 ( .A(x[869]), .B(y[869]), .Z(n6053) );
  NAND U3794 ( .A(n2593), .B(n6053), .Z(n2594) );
  AND U3795 ( .A(n6055), .B(n2594), .Z(n2595) );
  OR U3796 ( .A(n4128), .B(n2595), .Z(n2596) );
  NANDN U3797 ( .A(y[872]), .B(x[872]), .Z(n6061) );
  NAND U3798 ( .A(n2596), .B(n6061), .Z(n2597) );
  AND U3799 ( .A(n6059), .B(n2597), .Z(n2598) );
  NANDN U3800 ( .A(n6064), .B(n2598), .Z(n2599) );
  NANDN U3801 ( .A(n6066), .B(n2599), .Z(n2600) );
  AND U3802 ( .A(n6068), .B(n2600), .Z(n2603) );
  NANDN U3803 ( .A(y[877]), .B(x[877]), .Z(n2602) );
  NANDN U3804 ( .A(y[876]), .B(x[876]), .Z(n2601) );
  AND U3805 ( .A(n2602), .B(n2601), .Z(n6069) );
  NANDN U3806 ( .A(n2603), .B(n6069), .Z(n2606) );
  NANDN U3807 ( .A(x[877]), .B(y[877]), .Z(n2605) );
  NANDN U3808 ( .A(x[878]), .B(y[878]), .Z(n2604) );
  AND U3809 ( .A(n2605), .B(n2604), .Z(n6071) );
  NAND U3810 ( .A(n2606), .B(n6071), .Z(n2609) );
  NANDN U3811 ( .A(y[879]), .B(x[879]), .Z(n2608) );
  NANDN U3812 ( .A(y[878]), .B(x[878]), .Z(n2607) );
  AND U3813 ( .A(n2608), .B(n2607), .Z(n6073) );
  NAND U3814 ( .A(n2609), .B(n6073), .Z(n2612) );
  NANDN U3815 ( .A(x[879]), .B(y[879]), .Z(n2611) );
  NANDN U3816 ( .A(x[880]), .B(y[880]), .Z(n2610) );
  AND U3817 ( .A(n2611), .B(n2610), .Z(n6075) );
  NAND U3818 ( .A(n2612), .B(n6075), .Z(n2615) );
  NANDN U3819 ( .A(y[881]), .B(x[881]), .Z(n2614) );
  NANDN U3820 ( .A(y[880]), .B(x[880]), .Z(n2613) );
  AND U3821 ( .A(n2614), .B(n2613), .Z(n6077) );
  NAND U3822 ( .A(n2615), .B(n6077), .Z(n2616) );
  AND U3823 ( .A(n6081), .B(n2616), .Z(n2618) );
  NANDN U3824 ( .A(n2618), .B(n6083), .Z(n2619) );
  NANDN U3825 ( .A(n4149), .B(n2619), .Z(n2620) );
  NANDN U3826 ( .A(y[884]), .B(x[884]), .Z(n6087) );
  NAND U3827 ( .A(n2620), .B(n6087), .Z(n2621) );
  NANDN U3828 ( .A(n6090), .B(n2621), .Z(n2622) );
  NANDN U3829 ( .A(n6092), .B(n2622), .Z(n2623) );
  AND U3830 ( .A(n6093), .B(n2623), .Z(n2624) );
  NANDN U3831 ( .A(y[887]), .B(x[887]), .Z(n6095) );
  NANDN U3832 ( .A(n2624), .B(n6095), .Z(n2625) );
  NANDN U3833 ( .A(x[888]), .B(y[888]), .Z(n6098) );
  NAND U3834 ( .A(n2625), .B(n6098), .Z(n2628) );
  NANDN U3835 ( .A(y[889]), .B(x[889]), .Z(n2627) );
  NANDN U3836 ( .A(y[888]), .B(x[888]), .Z(n2626) );
  AND U3837 ( .A(n2627), .B(n2626), .Z(n6099) );
  NAND U3838 ( .A(n2628), .B(n6099), .Z(n2631) );
  NANDN U3839 ( .A(x[889]), .B(y[889]), .Z(n2630) );
  NANDN U3840 ( .A(x[890]), .B(y[890]), .Z(n2629) );
  AND U3841 ( .A(n2630), .B(n2629), .Z(n6101) );
  NAND U3842 ( .A(n2631), .B(n6101), .Z(n2634) );
  NANDN U3843 ( .A(y[891]), .B(x[891]), .Z(n2633) );
  NANDN U3844 ( .A(y[890]), .B(x[890]), .Z(n2632) );
  AND U3845 ( .A(n2633), .B(n2632), .Z(n6103) );
  NAND U3846 ( .A(n2634), .B(n6103), .Z(n2635) );
  AND U3847 ( .A(n6105), .B(n2635), .Z(n2636) );
  OR U3848 ( .A(n6108), .B(n2636), .Z(n2637) );
  NANDN U3849 ( .A(x[893]), .B(y[893]), .Z(n6109) );
  NAND U3850 ( .A(n2637), .B(n6109), .Z(n2638) );
  AND U3851 ( .A(n6111), .B(n2638), .Z(n2641) );
  NANDN U3852 ( .A(x[894]), .B(y[894]), .Z(n2640) );
  NANDN U3853 ( .A(x[895]), .B(y[895]), .Z(n2639) );
  AND U3854 ( .A(n2640), .B(n2639), .Z(n6113) );
  NANDN U3855 ( .A(n2641), .B(n6113), .Z(n2642) );
  NANDN U3856 ( .A(n6115), .B(n2642), .Z(n2645) );
  NANDN U3857 ( .A(x[896]), .B(y[896]), .Z(n2644) );
  NANDN U3858 ( .A(x[897]), .B(y[897]), .Z(n2643) );
  AND U3859 ( .A(n2644), .B(n2643), .Z(n6117) );
  NAND U3860 ( .A(n2645), .B(n6117), .Z(n2646) );
  NANDN U3861 ( .A(n6120), .B(n2646), .Z(n2649) );
  NANDN U3862 ( .A(x[899]), .B(y[899]), .Z(n2648) );
  NANDN U3863 ( .A(x[898]), .B(y[898]), .Z(n2647) );
  AND U3864 ( .A(n2648), .B(n2647), .Z(n6121) );
  NAND U3865 ( .A(n2649), .B(n6121), .Z(n2650) );
  AND U3866 ( .A(n6123), .B(n2650), .Z(n2651) );
  NANDN U3867 ( .A(x[900]), .B(y[900]), .Z(n6125) );
  NANDN U3868 ( .A(n2651), .B(n6125), .Z(n2652) );
  NANDN U3869 ( .A(n6127), .B(n2652), .Z(n2655) );
  NANDN U3870 ( .A(x[901]), .B(y[901]), .Z(n2654) );
  NANDN U3871 ( .A(x[902]), .B(y[902]), .Z(n2653) );
  AND U3872 ( .A(n2654), .B(n2653), .Z(n6129) );
  NAND U3873 ( .A(n2655), .B(n6129), .Z(n2656) );
  NANDN U3874 ( .A(n6132), .B(n2656), .Z(n2659) );
  NANDN U3875 ( .A(x[903]), .B(y[903]), .Z(n2658) );
  NANDN U3876 ( .A(x[904]), .B(y[904]), .Z(n2657) );
  AND U3877 ( .A(n2658), .B(n2657), .Z(n6133) );
  NAND U3878 ( .A(n2659), .B(n6133), .Z(n2662) );
  NANDN U3879 ( .A(y[905]), .B(x[905]), .Z(n2661) );
  NANDN U3880 ( .A(y[904]), .B(x[904]), .Z(n2660) );
  NAND U3881 ( .A(n2661), .B(n2660), .Z(n6136) );
  ANDN U3882 ( .B(n2662), .A(n6136), .Z(n2663) );
  NANDN U3883 ( .A(x[905]), .B(y[905]), .Z(n6138) );
  NANDN U3884 ( .A(n2663), .B(n6138), .Z(n2664) );
  NANDN U3885 ( .A(n6142), .B(n2664), .Z(n2670) );
  ANDN U3886 ( .B(y[906]), .A(x[906]), .Z(n6140) );
  ANDN U3887 ( .B(y[907]), .A(x[907]), .Z(n6143) );
  OR U3888 ( .A(n6140), .B(n6143), .Z(n2665) );
  NANDN U3889 ( .A(n2666), .B(n2665), .Z(n2669) );
  NANDN U3890 ( .A(x[909]), .B(y[909]), .Z(n2668) );
  NANDN U3891 ( .A(x[908]), .B(y[908]), .Z(n2667) );
  NAND U3892 ( .A(n2668), .B(n2667), .Z(n6147) );
  ANDN U3893 ( .B(n2669), .A(n6147), .Z(n4183) );
  NAND U3894 ( .A(n2670), .B(n4183), .Z(n2673) );
  NANDN U3895 ( .A(y[909]), .B(x[909]), .Z(n2672) );
  NANDN U3896 ( .A(y[910]), .B(x[910]), .Z(n2671) );
  AND U3897 ( .A(n2672), .B(n2671), .Z(n6149) );
  NAND U3898 ( .A(n2673), .B(n6149), .Z(n2676) );
  NANDN U3899 ( .A(x[910]), .B(y[910]), .Z(n2675) );
  NANDN U3900 ( .A(x[911]), .B(y[911]), .Z(n2674) );
  AND U3901 ( .A(n2675), .B(n2674), .Z(n6151) );
  NAND U3902 ( .A(n2676), .B(n6151), .Z(n2677) );
  AND U3903 ( .A(n6153), .B(n2677), .Z(n2678) );
  NANDN U3904 ( .A(x[912]), .B(y[912]), .Z(n6155) );
  NANDN U3905 ( .A(n2678), .B(n6155), .Z(n2681) );
  NANDN U3906 ( .A(y[912]), .B(x[912]), .Z(n2680) );
  NANDN U3907 ( .A(y[913]), .B(x[913]), .Z(n2679) );
  AND U3908 ( .A(n2680), .B(n2679), .Z(n6158) );
  NAND U3909 ( .A(n2681), .B(n6158), .Z(n2684) );
  NANDN U3910 ( .A(x[914]), .B(y[914]), .Z(n2683) );
  NANDN U3911 ( .A(x[913]), .B(y[913]), .Z(n2682) );
  AND U3912 ( .A(n2683), .B(n2682), .Z(n6159) );
  NAND U3913 ( .A(n2684), .B(n6159), .Z(n2687) );
  NANDN U3914 ( .A(y[914]), .B(x[914]), .Z(n2686) );
  NANDN U3915 ( .A(y[915]), .B(x[915]), .Z(n2685) );
  AND U3916 ( .A(n2686), .B(n2685), .Z(n6161) );
  NAND U3917 ( .A(n2687), .B(n6161), .Z(n2690) );
  NANDN U3918 ( .A(x[916]), .B(y[916]), .Z(n2689) );
  NANDN U3919 ( .A(x[915]), .B(y[915]), .Z(n2688) );
  AND U3920 ( .A(n2689), .B(n2688), .Z(n6163) );
  NAND U3921 ( .A(n2690), .B(n6163), .Z(n2691) );
  AND U3922 ( .A(n6165), .B(n2691), .Z(n2692) );
  NANDN U3923 ( .A(x[917]), .B(y[917]), .Z(n6168) );
  NANDN U3924 ( .A(n2692), .B(n6168), .Z(n2693) );
  NANDN U3925 ( .A(y[918]), .B(x[918]), .Z(n6172) );
  NAND U3926 ( .A(n2693), .B(n6172), .Z(n2694) );
  NANDN U3927 ( .A(x[919]), .B(y[919]), .Z(n6176) );
  ANDN U3928 ( .B(y[918]), .A(x[918]), .Z(n6170) );
  ANDN U3929 ( .B(n6176), .A(n6170), .Z(n4196) );
  NAND U3930 ( .A(n2694), .B(n4196), .Z(n2695) );
  NANDN U3931 ( .A(n4199), .B(n2695), .Z(n2698) );
  NANDN U3932 ( .A(x[921]), .B(y[921]), .Z(n2697) );
  NANDN U3933 ( .A(x[920]), .B(y[920]), .Z(n2696) );
  AND U3934 ( .A(n2697), .B(n2696), .Z(n6179) );
  NAND U3935 ( .A(n2698), .B(n6179), .Z(n2701) );
  NANDN U3936 ( .A(y[922]), .B(x[922]), .Z(n2700) );
  NANDN U3937 ( .A(y[921]), .B(x[921]), .Z(n2699) );
  NAND U3938 ( .A(n2700), .B(n2699), .Z(n6182) );
  ANDN U3939 ( .B(n2701), .A(n6182), .Z(n2702) );
  OR U3940 ( .A(n6184), .B(n2702), .Z(n2703) );
  NANDN U3941 ( .A(y[923]), .B(x[923]), .Z(n6185) );
  NAND U3942 ( .A(n2703), .B(n6185), .Z(n2704) );
  NANDN U3943 ( .A(x[924]), .B(y[924]), .Z(n6187) );
  NAND U3944 ( .A(n2704), .B(n6187), .Z(n2705) );
  NANDN U3945 ( .A(n6189), .B(n2705), .Z(n2708) );
  NANDN U3946 ( .A(x[925]), .B(y[925]), .Z(n2707) );
  NANDN U3947 ( .A(x[926]), .B(y[926]), .Z(n2706) );
  AND U3948 ( .A(n2707), .B(n2706), .Z(n6191) );
  NAND U3949 ( .A(n2708), .B(n6191), .Z(n2711) );
  NANDN U3950 ( .A(y[927]), .B(x[927]), .Z(n2710) );
  NANDN U3951 ( .A(y[926]), .B(x[926]), .Z(n2709) );
  NAND U3952 ( .A(n2710), .B(n2709), .Z(n6194) );
  ANDN U3953 ( .B(n2711), .A(n6194), .Z(n2714) );
  NANDN U3954 ( .A(x[927]), .B(y[927]), .Z(n2713) );
  NANDN U3955 ( .A(x[928]), .B(y[928]), .Z(n2712) );
  AND U3956 ( .A(n2713), .B(n2712), .Z(n6195) );
  NANDN U3957 ( .A(n2714), .B(n6195), .Z(n2717) );
  NANDN U3958 ( .A(y[929]), .B(x[929]), .Z(n2716) );
  NANDN U3959 ( .A(y[928]), .B(x[928]), .Z(n2715) );
  AND U3960 ( .A(n2716), .B(n2715), .Z(n6197) );
  NAND U3961 ( .A(n2717), .B(n6197), .Z(n2718) );
  AND U3962 ( .A(n6201), .B(n2718), .Z(n2721) );
  NANDN U3963 ( .A(y[930]), .B(x[930]), .Z(n2720) );
  ANDN U3964 ( .B(n2720), .A(n2719), .Z(n6204) );
  NANDN U3965 ( .A(n2721), .B(n6204), .Z(n2722) );
  NANDN U3966 ( .A(n4217), .B(n2722), .Z(n2723) );
  NANDN U3967 ( .A(y[932]), .B(x[932]), .Z(n2915) );
  NAND U3968 ( .A(n2723), .B(n2915), .Z(n2724) );
  NAND U3969 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U3970 ( .A(n2914), .B(n2726), .Z(n2727) );
  NANDN U3971 ( .A(y[934]), .B(x[934]), .Z(n6213) );
  NAND U3972 ( .A(n2727), .B(n6213), .Z(n2728) );
  NANDN U3973 ( .A(x[934]), .B(y[934]), .Z(n4220) );
  ANDN U3974 ( .B(y[935]), .A(x[935]), .Z(n4224) );
  ANDN U3975 ( .B(n4220), .A(n4224), .Z(n6215) );
  NAND U3976 ( .A(n2728), .B(n6215), .Z(n2729) );
  NANDN U3977 ( .A(y[935]), .B(x[935]), .Z(n6218) );
  NAND U3978 ( .A(n2729), .B(n6218), .Z(n2730) );
  AND U3979 ( .A(n6219), .B(n2730), .Z(n2733) );
  NANDN U3980 ( .A(y[936]), .B(x[936]), .Z(n2732) );
  NANDN U3981 ( .A(y[937]), .B(x[937]), .Z(n2731) );
  AND U3982 ( .A(n2732), .B(n2731), .Z(n6221) );
  NANDN U3983 ( .A(n2733), .B(n6221), .Z(n2734) );
  NANDN U3984 ( .A(n6224), .B(n2734), .Z(n2737) );
  NANDN U3985 ( .A(y[938]), .B(x[938]), .Z(n2736) );
  NANDN U3986 ( .A(y[939]), .B(x[939]), .Z(n2735) );
  AND U3987 ( .A(n2736), .B(n2735), .Z(n6225) );
  NAND U3988 ( .A(n2737), .B(n6225), .Z(n2738) );
  NANDN U3989 ( .A(n6228), .B(n2738), .Z(n2741) );
  NANDN U3990 ( .A(y[940]), .B(x[940]), .Z(n2740) );
  NANDN U3991 ( .A(y[941]), .B(x[941]), .Z(n2739) );
  AND U3992 ( .A(n2740), .B(n2739), .Z(n6230) );
  NAND U3993 ( .A(n2741), .B(n6230), .Z(n2742) );
  AND U3994 ( .A(n6232), .B(n2742), .Z(n2745) );
  NANDN U3995 ( .A(y[942]), .B(x[942]), .Z(n2744) );
  ANDN U3996 ( .B(n2744), .A(n2743), .Z(n6236) );
  NANDN U3997 ( .A(n2745), .B(n6236), .Z(n2746) );
  NANDN U3998 ( .A(n4234), .B(n2746), .Z(n2747) );
  NANDN U3999 ( .A(y[944]), .B(x[944]), .Z(n6239) );
  NAND U4000 ( .A(n2747), .B(n6239), .Z(n2748) );
  NANDN U4001 ( .A(x[945]), .B(y[945]), .Z(n6241) );
  NAND U4002 ( .A(n2748), .B(n6241), .Z(n2749) );
  NANDN U4003 ( .A(n6244), .B(n2749), .Z(n2751) );
  ANDN U4004 ( .B(y[947]), .A(x[947]), .Z(n2910) );
  NANDN U4005 ( .A(x[946]), .B(y[946]), .Z(n2750) );
  NANDN U4006 ( .A(n2910), .B(n2750), .Z(n6246) );
  ANDN U4007 ( .B(n2751), .A(n6246), .Z(n2752) );
  NANDN U4008 ( .A(y[947]), .B(x[947]), .Z(n6248) );
  NANDN U4009 ( .A(n2752), .B(n6248), .Z(n2753) );
  NANDN U4010 ( .A(x[948]), .B(y[948]), .Z(n6249) );
  NAND U4011 ( .A(n2753), .B(n6249), .Z(n2756) );
  NANDN U4012 ( .A(y[949]), .B(x[949]), .Z(n2755) );
  NANDN U4013 ( .A(y[948]), .B(x[948]), .Z(n2754) );
  AND U4014 ( .A(n2755), .B(n2754), .Z(n6251) );
  NAND U4015 ( .A(n2756), .B(n6251), .Z(n2759) );
  NANDN U4016 ( .A(x[949]), .B(y[949]), .Z(n2758) );
  NANDN U4017 ( .A(x[950]), .B(y[950]), .Z(n2757) );
  AND U4018 ( .A(n2758), .B(n2757), .Z(n6253) );
  NAND U4019 ( .A(n2759), .B(n6253), .Z(n2762) );
  NANDN U4020 ( .A(y[951]), .B(x[951]), .Z(n2761) );
  NANDN U4021 ( .A(y[950]), .B(x[950]), .Z(n2760) );
  AND U4022 ( .A(n2761), .B(n2760), .Z(n6255) );
  NAND U4023 ( .A(n2762), .B(n6255), .Z(n2763) );
  AND U4024 ( .A(n6257), .B(n2763), .Z(n2766) );
  NANDN U4025 ( .A(y[952]), .B(x[952]), .Z(n2765) );
  NANDN U4026 ( .A(y[953]), .B(x[953]), .Z(n2764) );
  AND U4027 ( .A(n2765), .B(n2764), .Z(n6260) );
  NANDN U4028 ( .A(n2766), .B(n6260), .Z(n2767) );
  NANDN U4029 ( .A(x[953]), .B(y[953]), .Z(n6261) );
  NAND U4030 ( .A(n2767), .B(n6261), .Z(n2768) );
  NANDN U4031 ( .A(y[954]), .B(x[954]), .Z(n6263) );
  NAND U4032 ( .A(n2768), .B(n6263), .Z(n2771) );
  NANDN U4033 ( .A(x[954]), .B(y[954]), .Z(n2770) );
  NANDN U4034 ( .A(x[955]), .B(y[955]), .Z(n2769) );
  AND U4035 ( .A(n2770), .B(n2769), .Z(n6265) );
  NAND U4036 ( .A(n2771), .B(n6265), .Z(n2774) );
  NANDN U4037 ( .A(y[956]), .B(x[956]), .Z(n2773) );
  NANDN U4038 ( .A(y[955]), .B(x[955]), .Z(n2772) );
  AND U4039 ( .A(n2773), .B(n2772), .Z(n6267) );
  NAND U4040 ( .A(n2774), .B(n6267), .Z(n2775) );
  AND U4041 ( .A(n6269), .B(n2775), .Z(n2778) );
  NANDN U4042 ( .A(y[958]), .B(x[958]), .Z(n2777) );
  NANDN U4043 ( .A(y[957]), .B(x[957]), .Z(n2776) );
  AND U4044 ( .A(n2777), .B(n2776), .Z(n6272) );
  NANDN U4045 ( .A(n2778), .B(n6272), .Z(n2781) );
  NANDN U4046 ( .A(x[959]), .B(y[959]), .Z(n2780) );
  NANDN U4047 ( .A(x[958]), .B(y[958]), .Z(n2779) );
  AND U4048 ( .A(n2780), .B(n2779), .Z(n6273) );
  NAND U4049 ( .A(n2781), .B(n6273), .Z(n2782) );
  NANDN U4050 ( .A(y[959]), .B(x[959]), .Z(n6275) );
  NAND U4051 ( .A(n2782), .B(n6275), .Z(n2783) );
  NANDN U4052 ( .A(x[960]), .B(y[960]), .Z(n6277) );
  NAND U4053 ( .A(n2783), .B(n6277), .Z(n2786) );
  NANDN U4054 ( .A(y[961]), .B(x[961]), .Z(n2785) );
  NANDN U4055 ( .A(y[960]), .B(x[960]), .Z(n2784) );
  AND U4056 ( .A(n2785), .B(n2784), .Z(n6279) );
  NAND U4057 ( .A(n2786), .B(n6279), .Z(n2787) );
  AND U4058 ( .A(n6281), .B(n2787), .Z(n2790) );
  NANDN U4059 ( .A(y[963]), .B(x[963]), .Z(n2789) );
  NANDN U4060 ( .A(y[962]), .B(x[962]), .Z(n2788) );
  AND U4061 ( .A(n2789), .B(n2788), .Z(n6284) );
  NANDN U4062 ( .A(n2790), .B(n6284), .Z(n2793) );
  NANDN U4063 ( .A(x[963]), .B(y[963]), .Z(n2792) );
  NANDN U4064 ( .A(x[964]), .B(y[964]), .Z(n2791) );
  AND U4065 ( .A(n2792), .B(n2791), .Z(n6285) );
  NAND U4066 ( .A(n2793), .B(n6285), .Z(n2796) );
  NANDN U4067 ( .A(y[964]), .B(x[964]), .Z(n2795) );
  NANDN U4068 ( .A(y[965]), .B(x[965]), .Z(n2794) );
  AND U4069 ( .A(n2795), .B(n2794), .Z(n6287) );
  NAND U4070 ( .A(n2796), .B(n6287), .Z(n2797) );
  NANDN U4071 ( .A(x[965]), .B(y[965]), .Z(n6289) );
  NAND U4072 ( .A(n2797), .B(n6289), .Z(n2798) );
  NANDN U4073 ( .A(y[966]), .B(x[966]), .Z(n6291) );
  NAND U4074 ( .A(n2798), .B(n6291), .Z(n2799) );
  AND U4075 ( .A(n6293), .B(n2799), .Z(n2802) );
  NANDN U4076 ( .A(y[968]), .B(x[968]), .Z(n2801) );
  NANDN U4077 ( .A(y[967]), .B(x[967]), .Z(n2800) );
  AND U4078 ( .A(n2801), .B(n2800), .Z(n6296) );
  NANDN U4079 ( .A(n2802), .B(n6296), .Z(n2805) );
  NANDN U4080 ( .A(x[968]), .B(y[968]), .Z(n2804) );
  NANDN U4081 ( .A(x[969]), .B(y[969]), .Z(n2803) );
  AND U4082 ( .A(n2804), .B(n2803), .Z(n6297) );
  NAND U4083 ( .A(n2805), .B(n6297), .Z(n2808) );
  NANDN U4084 ( .A(y[970]), .B(x[970]), .Z(n2807) );
  NANDN U4085 ( .A(y[969]), .B(x[969]), .Z(n2806) );
  AND U4086 ( .A(n2807), .B(n2806), .Z(n6299) );
  NAND U4087 ( .A(n2808), .B(n6299), .Z(n2811) );
  NANDN U4088 ( .A(x[971]), .B(y[971]), .Z(n2810) );
  NANDN U4089 ( .A(x[970]), .B(y[970]), .Z(n2809) );
  AND U4090 ( .A(n2810), .B(n2809), .Z(n6301) );
  NAND U4091 ( .A(n2811), .B(n6301), .Z(n2812) );
  NANDN U4092 ( .A(y[971]), .B(x[971]), .Z(n6303) );
  NAND U4093 ( .A(n2812), .B(n6303), .Z(n2813) );
  AND U4094 ( .A(n6305), .B(n2813), .Z(n2816) );
  NANDN U4095 ( .A(y[973]), .B(x[973]), .Z(n2815) );
  NANDN U4096 ( .A(y[972]), .B(x[972]), .Z(n2814) );
  AND U4097 ( .A(n2815), .B(n2814), .Z(n6308) );
  NANDN U4098 ( .A(n2816), .B(n6308), .Z(n2819) );
  NANDN U4099 ( .A(x[973]), .B(y[973]), .Z(n2818) );
  NANDN U4100 ( .A(x[974]), .B(y[974]), .Z(n2817) );
  AND U4101 ( .A(n2818), .B(n2817), .Z(n6309) );
  NAND U4102 ( .A(n2819), .B(n6309), .Z(n2822) );
  NANDN U4103 ( .A(y[975]), .B(x[975]), .Z(n2821) );
  NANDN U4104 ( .A(y[974]), .B(x[974]), .Z(n2820) );
  AND U4105 ( .A(n2821), .B(n2820), .Z(n6311) );
  NAND U4106 ( .A(n2822), .B(n6311), .Z(n2825) );
  NANDN U4107 ( .A(x[975]), .B(y[975]), .Z(n2824) );
  NANDN U4108 ( .A(x[976]), .B(y[976]), .Z(n2823) );
  AND U4109 ( .A(n2824), .B(n2823), .Z(n6313) );
  NAND U4110 ( .A(n2825), .B(n6313), .Z(n2828) );
  NANDN U4111 ( .A(y[977]), .B(x[977]), .Z(n2827) );
  NANDN U4112 ( .A(y[976]), .B(x[976]), .Z(n2826) );
  AND U4113 ( .A(n2827), .B(n2826), .Z(n6315) );
  NAND U4114 ( .A(n2828), .B(n6315), .Z(n2829) );
  AND U4115 ( .A(n6318), .B(n2829), .Z(n2832) );
  NANDN U4116 ( .A(y[978]), .B(x[978]), .Z(n2831) );
  ANDN U4117 ( .B(n2831), .A(n2830), .Z(n6321) );
  NANDN U4118 ( .A(n2832), .B(n6321), .Z(n2833) );
  NANDN U4119 ( .A(n4284), .B(n2833), .Z(n2834) );
  NANDN U4120 ( .A(y[980]), .B(x[980]), .Z(n6326) );
  NAND U4121 ( .A(n2834), .B(n6326), .Z(n2835) );
  NANDN U4122 ( .A(n6328), .B(n2835), .Z(n2836) );
  NANDN U4123 ( .A(n6330), .B(n2836), .Z(n2837) );
  AND U4124 ( .A(n6331), .B(n2837), .Z(n2838) );
  NANDN U4125 ( .A(y[983]), .B(x[983]), .Z(n6334) );
  NANDN U4126 ( .A(n2838), .B(n6334), .Z(n2839) );
  NANDN U4127 ( .A(x[984]), .B(y[984]), .Z(n6335) );
  NAND U4128 ( .A(n2839), .B(n6335), .Z(n2842) );
  NANDN U4129 ( .A(y[984]), .B(x[984]), .Z(n2841) );
  NANDN U4130 ( .A(y[985]), .B(x[985]), .Z(n2840) );
  AND U4131 ( .A(n2841), .B(n2840), .Z(n6338) );
  NAND U4132 ( .A(n2842), .B(n6338), .Z(n2843) );
  NANDN U4133 ( .A(n6340), .B(n2843), .Z(n2846) );
  NANDN U4134 ( .A(y[986]), .B(x[986]), .Z(n2845) );
  NANDN U4135 ( .A(y[987]), .B(x[987]), .Z(n2844) );
  AND U4136 ( .A(n2845), .B(n2844), .Z(n6341) );
  NAND U4137 ( .A(n2846), .B(n6341), .Z(n2849) );
  NANDN U4138 ( .A(x[988]), .B(y[988]), .Z(n2848) );
  NANDN U4139 ( .A(x[987]), .B(y[987]), .Z(n2847) );
  NAND U4140 ( .A(n2848), .B(n2847), .Z(n6344) );
  ANDN U4141 ( .B(n2849), .A(n6344), .Z(n2852) );
  NANDN U4142 ( .A(y[988]), .B(x[988]), .Z(n2851) );
  NANDN U4143 ( .A(y[989]), .B(x[989]), .Z(n2850) );
  AND U4144 ( .A(n2851), .B(n2850), .Z(n6345) );
  NANDN U4145 ( .A(n2852), .B(n6345), .Z(n2853) );
  NANDN U4146 ( .A(n4360), .B(n2853), .Z(n2854) );
  NANDN U4147 ( .A(y[990]), .B(x[990]), .Z(n4358) );
  NAND U4148 ( .A(n2854), .B(n4358), .Z(n2855) );
  NAND U4149 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U4150 ( .A(n2907), .B(n2857), .Z(n2858) );
  OR U4151 ( .A(n4310), .B(n2858), .Z(n2860) );
  NANDN U4152 ( .A(y[994]), .B(x[994]), .Z(n2859) );
  ANDN U4153 ( .B(x[993]), .A(y[993]), .Z(n2909) );
  ANDN U4154 ( .B(n2859), .A(n2909), .Z(n6353) );
  NAND U4155 ( .A(n2860), .B(n6353), .Z(n2861) );
  NANDN U4156 ( .A(n6358), .B(n2861), .Z(n2862) );
  NANDN U4157 ( .A(y[995]), .B(x[995]), .Z(n6359) );
  NAND U4158 ( .A(n2862), .B(n6359), .Z(n2863) );
  NANDN U4159 ( .A(x[996]), .B(y[996]), .Z(n6361) );
  NAND U4160 ( .A(n2863), .B(n6361), .Z(n2866) );
  NANDN U4161 ( .A(y[997]), .B(x[997]), .Z(n2865) );
  NANDN U4162 ( .A(y[996]), .B(x[996]), .Z(n2864) );
  NAND U4163 ( .A(n2865), .B(n2864), .Z(n6364) );
  ANDN U4164 ( .B(n2866), .A(n6364), .Z(n2869) );
  NANDN U4165 ( .A(x[997]), .B(y[997]), .Z(n2868) );
  NANDN U4166 ( .A(x[998]), .B(y[998]), .Z(n2867) );
  AND U4167 ( .A(n2868), .B(n2867), .Z(n6366) );
  NANDN U4168 ( .A(n2869), .B(n6366), .Z(n2870) );
  NANDN U4169 ( .A(n6368), .B(n2870), .Z(n2873) );
  NANDN U4170 ( .A(x[999]), .B(y[999]), .Z(n2872) );
  NANDN U4171 ( .A(x[1000]), .B(y[1000]), .Z(n2871) );
  AND U4172 ( .A(n2872), .B(n2871), .Z(n6369) );
  NAND U4173 ( .A(n2873), .B(n6369), .Z(n2874) );
  NANDN U4174 ( .A(x[1001]), .B(y[1001]), .Z(n6375) );
  NANDN U4175 ( .A(n2874), .B(n6375), .Z(n2875) );
  NANDN U4176 ( .A(y[1002]), .B(x[1002]), .Z(n4356) );
  NAND U4177 ( .A(n2875), .B(n4356), .Z(n2876) );
  NANDN U4178 ( .A(n4331), .B(n2876), .Z(n2877) );
  NANDN U4179 ( .A(y[1003]), .B(x[1003]), .Z(n4357) );
  NAND U4180 ( .A(n2877), .B(n4357), .Z(n2878) );
  NANDN U4181 ( .A(n2879), .B(n2878), .Z(n2880) );
  NANDN U4182 ( .A(y[1006]), .B(x[1006]), .Z(n4340) );
  IV U4183 ( .A(n4340), .Z(n6387) );
  ANDN U4184 ( .B(n2880), .A(n6387), .Z(n2881) );
  NANDN U4185 ( .A(y[1005]), .B(x[1005]), .Z(n4334) );
  NAND U4186 ( .A(n2881), .B(n4334), .Z(n2882) );
  AND U4187 ( .A(n6393), .B(n2882), .Z(n2884) );
  NANDN U4188 ( .A(x[1007]), .B(y[1007]), .Z(n2883) );
  ANDN U4189 ( .B(y[1006]), .A(x[1006]), .Z(n4337) );
  ANDN U4190 ( .B(n2883), .A(n4337), .Z(n6389) );
  NAND U4191 ( .A(n2884), .B(n6389), .Z(n2887) );
  NANDN U4192 ( .A(y[1008]), .B(x[1008]), .Z(n2886) );
  NANDN U4193 ( .A(y[1009]), .B(x[1009]), .Z(n2885) );
  AND U4194 ( .A(n2886), .B(n2885), .Z(n6395) );
  NAND U4195 ( .A(n2887), .B(n6395), .Z(n2890) );
  NANDN U4196 ( .A(x[1010]), .B(y[1010]), .Z(n2889) );
  NANDN U4197 ( .A(x[1009]), .B(y[1009]), .Z(n2888) );
  AND U4198 ( .A(n2889), .B(n2888), .Z(n6398) );
  NAND U4199 ( .A(n2890), .B(n6398), .Z(n2891) );
  AND U4200 ( .A(n6399), .B(n2891), .Z(n2897) );
  NANDN U4201 ( .A(x[1014]), .B(y[1014]), .Z(n2893) );
  NANDN U4202 ( .A(x[1013]), .B(y[1013]), .Z(n2892) );
  AND U4203 ( .A(n2893), .B(n2892), .Z(n6405) );
  NANDN U4204 ( .A(x[1012]), .B(y[1012]), .Z(n2895) );
  NANDN U4205 ( .A(x[1011]), .B(y[1011]), .Z(n2894) );
  NAND U4206 ( .A(n2895), .B(n2894), .Z(n6402) );
  ANDN U4207 ( .B(n6405), .A(n6402), .Z(n2896) );
  NANDN U4208 ( .A(n2897), .B(n2896), .Z(n2900) );
  NAND U4209 ( .A(n2899), .B(n2898), .Z(n6408) );
  ANDN U4210 ( .B(n2900), .A(n6408), .Z(n2901) );
  ANDN U4211 ( .B(n2902), .A(n2901), .Z(n4354) );
  NANDN U4212 ( .A(y[1012]), .B(x[1012]), .Z(n2904) );
  NANDN U4213 ( .A(y[1013]), .B(x[1013]), .Z(n2903) );
  NAND U4214 ( .A(n2904), .B(n2903), .Z(n6404) );
  NANDN U4215 ( .A(y[1001]), .B(x[1001]), .Z(n2906) );
  NANDN U4216 ( .A(y[1000]), .B(x[1000]), .Z(n2905) );
  NAND U4217 ( .A(n2906), .B(n2905), .Z(n6372) );
  XNOR U4218 ( .A(y[994]), .B(x[994]), .Z(n4316) );
  ANDN U4219 ( .B(n2908), .A(n2907), .Z(n6355) );
  NOR U4220 ( .A(n6355), .B(n2909), .Z(n4314) );
  ANDN U4221 ( .B(n6249), .A(n2910), .Z(n4245) );
  NANDN U4222 ( .A(y[946]), .B(x[946]), .Z(n2911) );
  AND U4223 ( .A(n6248), .B(n2911), .Z(n4243) );
  XNOR U4224 ( .A(n2913), .B(n2912), .Z(n4241) );
  NAND U4225 ( .A(n2915), .B(n2914), .Z(n6210) );
  NAND U4226 ( .A(n2916), .B(n6095), .Z(n2917) );
  AND U4227 ( .A(n2918), .B(n2917), .Z(n4160) );
  AND U4228 ( .A(n6061), .B(n2919), .Z(n4130) );
  XOR U4229 ( .A(x[862]), .B(n2920), .Z(n4112) );
  ANDN U4230 ( .B(n6010), .A(n2921), .Z(n4097) );
  NANDN U4231 ( .A(y[850]), .B(x[850]), .Z(n2922) );
  AND U4232 ( .A(n6007), .B(n2922), .Z(n4095) );
  XNOR U4233 ( .A(n2924), .B(n2923), .Z(n4093) );
  NANDN U4234 ( .A(n2926), .B(n2925), .Z(n3856) );
  NANDN U4235 ( .A(x[624]), .B(y[624]), .Z(n2927) );
  AND U4236 ( .A(n2928), .B(n2927), .Z(n2930) );
  NANDN U4237 ( .A(n2930), .B(n2929), .Z(n2931) );
  NAND U4238 ( .A(n2932), .B(n2931), .Z(n5536) );
  NANDN U4239 ( .A(n2934), .B(n2933), .Z(n3823) );
  NANDN U4240 ( .A(n2936), .B(n2935), .Z(n2937) );
  NANDN U4241 ( .A(n2938), .B(n2937), .Z(n5512) );
  NANDN U4242 ( .A(n2940), .B(n2939), .Z(n2941) );
  NANDN U4243 ( .A(n2942), .B(n2941), .Z(n5500) );
  NAND U4244 ( .A(n2944), .B(n2943), .Z(n2946) );
  NAND U4245 ( .A(n2946), .B(n2945), .Z(n5496) );
  NANDN U4246 ( .A(y[582]), .B(x[582]), .Z(n2947) );
  AND U4247 ( .A(n2948), .B(n2947), .Z(n3782) );
  XNOR U4248 ( .A(n2950), .B(n2949), .Z(n3780) );
  NANDN U4249 ( .A(n2952), .B(n2951), .Z(n2953) );
  NANDN U4250 ( .A(n2954), .B(n2953), .Z(n5048) );
  NANDN U4251 ( .A(n2956), .B(n2955), .Z(n2957) );
  NANDN U4252 ( .A(n2958), .B(n2957), .Z(n4707) );
  NANDN U4253 ( .A(n2960), .B(n2959), .Z(n2961) );
  NANDN U4254 ( .A(n2962), .B(n2961), .Z(n4623) );
  NANDN U4255 ( .A(n2964), .B(n2963), .Z(n2965) );
  NANDN U4256 ( .A(n2966), .B(n2965), .Z(n4584) );
  NANDN U4257 ( .A(n2968), .B(n2967), .Z(n2969) );
  NANDN U4258 ( .A(n2970), .B(n2969), .Z(n4498) );
  NAND U4259 ( .A(n2972), .B(n2971), .Z(n2973) );
  NANDN U4260 ( .A(n2974), .B(n2973), .Z(n4462) );
  NANDN U4261 ( .A(x[20]), .B(y[20]), .Z(n3044) );
  ANDN U4262 ( .B(n2976), .A(n2975), .Z(n3038) );
  ANDN U4263 ( .B(n2978), .A(n2977), .Z(n3032) );
  NANDN U4264 ( .A(n2980), .B(n2979), .Z(n3010) );
  ANDN U4265 ( .B(n2982), .A(n2981), .Z(n2994) );
  ANDN U4266 ( .B(x[0]), .A(y[0]), .Z(n2984) );
  ANDN U4267 ( .B(x[1]), .A(y[1]), .Z(n2983) );
  OR U4268 ( .A(n2984), .B(n2983), .Z(n2988) );
  AND U4269 ( .A(n2986), .B(n2985), .Z(n2987) );
  NAND U4270 ( .A(n2988), .B(n2987), .Z(n2989) );
  NANDN U4271 ( .A(n2990), .B(n2989), .Z(n2991) );
  OR U4272 ( .A(n2992), .B(n2991), .Z(n2993) );
  AND U4273 ( .A(n2994), .B(n2993), .Z(n2996) );
  NOR U4274 ( .A(n2996), .B(n2995), .Z(n2997) );
  NANDN U4275 ( .A(n2998), .B(n2997), .Z(n3000) );
  ANDN U4276 ( .B(n3000), .A(n2999), .Z(n3002) );
  NAND U4277 ( .A(n3002), .B(n3001), .Z(n3006) );
  NANDN U4278 ( .A(y[6]), .B(x[6]), .Z(n3004) );
  ANDN U4279 ( .B(n3004), .A(n3003), .Z(n3005) );
  NAND U4280 ( .A(n3006), .B(n3005), .Z(n3008) );
  ANDN U4281 ( .B(n3008), .A(n3007), .Z(n3009) );
  NAND U4282 ( .A(n3010), .B(n3009), .Z(n3011) );
  NANDN U4283 ( .A(n3012), .B(n3011), .Z(n3013) );
  NANDN U4284 ( .A(n3014), .B(n3013), .Z(n3015) );
  NANDN U4285 ( .A(n3016), .B(n3015), .Z(n3018) );
  ANDN U4286 ( .B(n3018), .A(n3017), .Z(n3020) );
  NOR U4287 ( .A(n3020), .B(n3019), .Z(n3021) );
  NANDN U4288 ( .A(n3022), .B(n3021), .Z(n3024) );
  ANDN U4289 ( .B(n3024), .A(n3023), .Z(n3025) );
  NANDN U4290 ( .A(n3026), .B(n3025), .Z(n3028) );
  ANDN U4291 ( .B(n3028), .A(n3027), .Z(n3029) );
  NANDN U4292 ( .A(n3030), .B(n3029), .Z(n3031) );
  NAND U4293 ( .A(n3032), .B(n3031), .Z(n3033) );
  NANDN U4294 ( .A(n3034), .B(n3033), .Z(n3035) );
  OR U4295 ( .A(n3036), .B(n3035), .Z(n3037) );
  AND U4296 ( .A(n3038), .B(n3037), .Z(n3040) );
  NOR U4297 ( .A(n3040), .B(n3039), .Z(n3041) );
  NANDN U4298 ( .A(n3042), .B(n3041), .Z(n3043) );
  AND U4299 ( .A(n3044), .B(n3043), .Z(n3045) );
  NANDN U4300 ( .A(n3046), .B(n3045), .Z(n3050) );
  NANDN U4301 ( .A(y[20]), .B(x[20]), .Z(n3047) );
  AND U4302 ( .A(n3048), .B(n3047), .Z(n3049) );
  NAND U4303 ( .A(n3050), .B(n3049), .Z(n3052) );
  ANDN U4304 ( .B(n3052), .A(n3051), .Z(n3053) );
  OR U4305 ( .A(n3054), .B(n3053), .Z(n3055) );
  NANDN U4306 ( .A(n3056), .B(n3055), .Z(n3057) );
  NANDN U4307 ( .A(n3058), .B(n3057), .Z(n3059) );
  NANDN U4308 ( .A(n3060), .B(n3059), .Z(n3061) );
  NANDN U4309 ( .A(n3062), .B(n3061), .Z(n3064) );
  ANDN U4310 ( .B(n3064), .A(n3063), .Z(n3065) );
  OR U4311 ( .A(n3066), .B(n3065), .Z(n3067) );
  NANDN U4312 ( .A(n3068), .B(n3067), .Z(n3069) );
  NANDN U4313 ( .A(n3070), .B(n3069), .Z(n3071) );
  NANDN U4314 ( .A(n3072), .B(n3071), .Z(n3073) );
  NANDN U4315 ( .A(n3074), .B(n3073), .Z(n3076) );
  ANDN U4316 ( .B(n3076), .A(n3075), .Z(n3077) );
  OR U4317 ( .A(n3078), .B(n3077), .Z(n3080) );
  NAND U4318 ( .A(n3080), .B(n3079), .Z(n3084) );
  OR U4319 ( .A(n3084), .B(y[36]), .Z(n3082) );
  ANDN U4320 ( .B(n3082), .A(n3081), .Z(n3087) );
  XNOR U4321 ( .A(n3084), .B(n3083), .Z(n3085) );
  NAND U4322 ( .A(x[36]), .B(n3085), .Z(n3086) );
  NAND U4323 ( .A(n3087), .B(n3086), .Z(n3088) );
  NANDN U4324 ( .A(n3089), .B(n3088), .Z(n3090) );
  NANDN U4325 ( .A(n3091), .B(n3090), .Z(n3093) );
  ANDN U4326 ( .B(n3093), .A(n3092), .Z(n3094) );
  OR U4327 ( .A(n3095), .B(n3094), .Z(n3096) );
  NANDN U4328 ( .A(n3097), .B(n3096), .Z(n3098) );
  NANDN U4329 ( .A(n3099), .B(n3098), .Z(n3100) );
  NANDN U4330 ( .A(n3101), .B(n3100), .Z(n3102) );
  NANDN U4331 ( .A(n3103), .B(n3102), .Z(n3105) );
  ANDN U4332 ( .B(n3105), .A(n3104), .Z(n3106) );
  OR U4333 ( .A(n3107), .B(n3106), .Z(n3108) );
  NANDN U4334 ( .A(n3109), .B(n3108), .Z(n3110) );
  NANDN U4335 ( .A(n3111), .B(n3110), .Z(n3112) );
  NANDN U4336 ( .A(n3113), .B(n3112), .Z(n3114) );
  NANDN U4337 ( .A(n3115), .B(n3114), .Z(n3117) );
  ANDN U4338 ( .B(n3117), .A(n3116), .Z(n3118) );
  OR U4339 ( .A(n3119), .B(n3118), .Z(n3120) );
  NANDN U4340 ( .A(n3121), .B(n3120), .Z(n3122) );
  NANDN U4341 ( .A(n3123), .B(n3122), .Z(n3124) );
  NANDN U4342 ( .A(n3125), .B(n3124), .Z(n3126) );
  NANDN U4343 ( .A(n3127), .B(n3126), .Z(n3129) );
  ANDN U4344 ( .B(n3129), .A(n3128), .Z(n3130) );
  OR U4345 ( .A(n3131), .B(n3130), .Z(n3132) );
  NANDN U4346 ( .A(n3133), .B(n3132), .Z(n3134) );
  NANDN U4347 ( .A(n3135), .B(n3134), .Z(n3136) );
  NANDN U4348 ( .A(n3137), .B(n3136), .Z(n3138) );
  NANDN U4349 ( .A(n3139), .B(n3138), .Z(n3141) );
  ANDN U4350 ( .B(n3141), .A(n3140), .Z(n3142) );
  OR U4351 ( .A(n3143), .B(n3142), .Z(n3144) );
  NANDN U4352 ( .A(n3145), .B(n3144), .Z(n3146) );
  NANDN U4353 ( .A(n3147), .B(n3146), .Z(n3149) );
  AND U4354 ( .A(n3149), .B(n3148), .Z(n4378) );
  NAND U4355 ( .A(n4378), .B(n4379), .Z(n3150) );
  NANDN U4356 ( .A(n3151), .B(n3150), .Z(n3152) );
  AND U4357 ( .A(n4383), .B(n3152), .Z(n3153) );
  NANDN U4358 ( .A(n3153), .B(n4385), .Z(n3154) );
  NANDN U4359 ( .A(n4387), .B(n3154), .Z(n3155) );
  NAND U4360 ( .A(n3155), .B(n4389), .Z(n3156) );
  NANDN U4361 ( .A(n4392), .B(n3156), .Z(n3157) );
  NAND U4362 ( .A(n3157), .B(n4393), .Z(n3158) );
  ANDN U4363 ( .B(n3158), .A(n4396), .Z(n3159) );
  NANDN U4364 ( .A(n3159), .B(n4397), .Z(n3160) );
  NANDN U4365 ( .A(n4399), .B(n3160), .Z(n3161) );
  NAND U4366 ( .A(n3161), .B(n4401), .Z(n3162) );
  NANDN U4367 ( .A(n4404), .B(n3162), .Z(n3163) );
  NAND U4368 ( .A(n3163), .B(n4405), .Z(n3164) );
  ANDN U4369 ( .B(n3164), .A(n4408), .Z(n3165) );
  NANDN U4370 ( .A(n3165), .B(n4409), .Z(n3166) );
  NANDN U4371 ( .A(n4411), .B(n3166), .Z(n3167) );
  NAND U4372 ( .A(n3167), .B(n4413), .Z(n3168) );
  NANDN U4373 ( .A(n3169), .B(n3168), .Z(n3170) );
  NANDN U4374 ( .A(n3171), .B(n3170), .Z(n3172) );
  AND U4375 ( .A(n4423), .B(n3172), .Z(n3173) );
  NANDN U4376 ( .A(n3173), .B(n4425), .Z(n3174) );
  NANDN U4377 ( .A(n4427), .B(n3174), .Z(n3175) );
  NAND U4378 ( .A(n3175), .B(n4429), .Z(n3176) );
  NANDN U4379 ( .A(n4432), .B(n3176), .Z(n3177) );
  NAND U4380 ( .A(n3177), .B(n4433), .Z(n3178) );
  ANDN U4381 ( .B(n3178), .A(n4436), .Z(n3179) );
  NANDN U4382 ( .A(n3179), .B(n4437), .Z(n3180) );
  NANDN U4383 ( .A(n4439), .B(n3180), .Z(n3181) );
  NAND U4384 ( .A(n3181), .B(n4441), .Z(n3182) );
  NANDN U4385 ( .A(n4444), .B(n3182), .Z(n3183) );
  NAND U4386 ( .A(n3183), .B(n4445), .Z(n3185) );
  ANDN U4387 ( .B(n3185), .A(n3184), .Z(n3187) );
  OR U4388 ( .A(n3187), .B(n3186), .Z(n3188) );
  NANDN U4389 ( .A(n4458), .B(n3188), .Z(n3189) );
  NAND U4390 ( .A(n3189), .B(n4459), .Z(n3190) );
  NANDN U4391 ( .A(n4462), .B(n3190), .Z(n3191) );
  NAND U4392 ( .A(n3191), .B(n4463), .Z(n3192) );
  ANDN U4393 ( .B(n3192), .A(n4465), .Z(n3193) );
  NANDN U4394 ( .A(n3193), .B(n4467), .Z(n3194) );
  NANDN U4395 ( .A(n4470), .B(n3194), .Z(n3195) );
  NAND U4396 ( .A(n3195), .B(n4471), .Z(n3196) );
  NANDN U4397 ( .A(n3197), .B(n3196), .Z(n3198) );
  NANDN U4398 ( .A(n3199), .B(n3198), .Z(n3200) );
  AND U4399 ( .A(n4481), .B(n3200), .Z(n3201) );
  NANDN U4400 ( .A(n3201), .B(n4483), .Z(n3202) );
  NANDN U4401 ( .A(n4486), .B(n3202), .Z(n3203) );
  NAND U4402 ( .A(n3203), .B(n4487), .Z(n3204) );
  NANDN U4403 ( .A(n4490), .B(n3204), .Z(n3205) );
  NAND U4404 ( .A(n3205), .B(n4492), .Z(n3206) );
  AND U4405 ( .A(n4493), .B(n3206), .Z(n3207) );
  OR U4406 ( .A(n3207), .B(n4496), .Z(n3208) );
  NANDN U4407 ( .A(n4498), .B(n3208), .Z(n3209) );
  NAND U4408 ( .A(n3209), .B(n4499), .Z(n3210) );
  NANDN U4409 ( .A(n3211), .B(n3210), .Z(n3212) );
  NANDN U4410 ( .A(n3213), .B(n3212), .Z(n3214) );
  AND U4411 ( .A(n4509), .B(n3214), .Z(n3215) );
  NANDN U4412 ( .A(n3215), .B(n4511), .Z(n3216) );
  AND U4413 ( .A(n3217), .B(n3216), .Z(n3219) );
  ANDN U4414 ( .B(x[128]), .A(y[128]), .Z(n3218) );
  OR U4415 ( .A(n3219), .B(n3218), .Z(n3220) );
  NANDN U4416 ( .A(n3221), .B(n3220), .Z(n3223) );
  NAND U4417 ( .A(n3223), .B(n3222), .Z(n3224) );
  NAND U4418 ( .A(n3224), .B(n4517), .Z(n3225) );
  NAND U4419 ( .A(n3225), .B(n4519), .Z(n3226) );
  ANDN U4420 ( .B(n3226), .A(n4522), .Z(n3227) );
  NANDN U4421 ( .A(n3227), .B(n4523), .Z(n3228) );
  NANDN U4422 ( .A(n3229), .B(n3228), .Z(n3230) );
  NANDN U4423 ( .A(n3231), .B(n3230), .Z(n3232) );
  NANDN U4424 ( .A(n4532), .B(n3232), .Z(n3233) );
  NAND U4425 ( .A(n3233), .B(n4533), .Z(n3234) );
  ANDN U4426 ( .B(n3234), .A(n4535), .Z(n3235) );
  NANDN U4427 ( .A(n3235), .B(n4537), .Z(n3236) );
  AND U4428 ( .A(n3237), .B(n3236), .Z(n3239) );
  ANDN U4429 ( .B(x[140]), .A(y[140]), .Z(n3238) );
  OR U4430 ( .A(n3239), .B(n3238), .Z(n3240) );
  NANDN U4431 ( .A(n3241), .B(n3240), .Z(n3243) );
  NAND U4432 ( .A(n3243), .B(n3242), .Z(n3244) );
  NAND U4433 ( .A(n3244), .B(n4545), .Z(n3245) );
  NANDN U4434 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U4435 ( .A(n3247), .B(n4549), .Z(n3248) );
  NAND U4436 ( .A(n3248), .B(n4551), .Z(n3249) );
  NAND U4437 ( .A(n3249), .B(n4554), .Z(n3250) );
  AND U4438 ( .A(n4555), .B(n3250), .Z(n3251) );
  NANDN U4439 ( .A(n3251), .B(n4557), .Z(n3252) );
  NAND U4440 ( .A(n3252), .B(n4559), .Z(n3253) );
  NAND U4441 ( .A(n3253), .B(n4561), .Z(n3254) );
  NAND U4442 ( .A(n3254), .B(n4563), .Z(n3255) );
  NANDN U4443 ( .A(n3256), .B(n3255), .Z(n3258) );
  ANDN U4444 ( .B(n3258), .A(n3257), .Z(n3259) );
  NANDN U4445 ( .A(n3259), .B(n4571), .Z(n3260) );
  NANDN U4446 ( .A(n4574), .B(n3260), .Z(n3261) );
  NAND U4447 ( .A(n3261), .B(n4576), .Z(n3262) );
  NAND U4448 ( .A(n3262), .B(n4577), .Z(n3263) );
  NAND U4449 ( .A(n3263), .B(n4579), .Z(n3264) );
  AND U4450 ( .A(n4581), .B(n3264), .Z(n3265) );
  OR U4451 ( .A(n4584), .B(n3265), .Z(n3266) );
  NAND U4452 ( .A(n3266), .B(n4585), .Z(n3268) );
  NAND U4453 ( .A(n3268), .B(n3267), .Z(n3269) );
  NAND U4454 ( .A(n3270), .B(n3269), .Z(n3271) );
  NANDN U4455 ( .A(n3272), .B(n3271), .Z(n3274) );
  ANDN U4456 ( .B(n3274), .A(n3273), .Z(n3275) );
  NANDN U4457 ( .A(n3275), .B(n4591), .Z(n3276) );
  NAND U4458 ( .A(n3276), .B(n4593), .Z(n3277) );
  NANDN U4459 ( .A(n3278), .B(n3277), .Z(n3280) );
  NAND U4460 ( .A(n3280), .B(n3279), .Z(n3281) );
  NANDN U4461 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U4462 ( .A(n4608), .B(n3283), .Z(n3284) );
  NANDN U4463 ( .A(n3284), .B(n4610), .Z(n3285) );
  NAND U4464 ( .A(n3285), .B(n4613), .Z(n3286) );
  NAND U4465 ( .A(n3286), .B(n4614), .Z(n3287) );
  NAND U4466 ( .A(n3287), .B(n4616), .Z(n3288) );
  NAND U4467 ( .A(n3288), .B(n4618), .Z(n3289) );
  ANDN U4468 ( .B(n3289), .A(n4621), .Z(n3290) );
  OR U4469 ( .A(n4623), .B(n3290), .Z(n3291) );
  NAND U4470 ( .A(n3291), .B(n4625), .Z(n3293) );
  NAND U4471 ( .A(n3293), .B(n3292), .Z(n3294) );
  NAND U4472 ( .A(n3295), .B(n3294), .Z(n3296) );
  NANDN U4473 ( .A(n3297), .B(n3296), .Z(n3299) );
  ANDN U4474 ( .B(n3299), .A(n3298), .Z(n3300) );
  NANDN U4475 ( .A(n3300), .B(n4630), .Z(n3301) );
  NAND U4476 ( .A(n3301), .B(n4632), .Z(n3302) );
  NAND U4477 ( .A(n3302), .B(n4634), .Z(n3303) );
  NAND U4478 ( .A(n3303), .B(n4637), .Z(n3304) );
  NAND U4479 ( .A(n3304), .B(n4638), .Z(n3305) );
  AND U4480 ( .A(n4640), .B(n3305), .Z(n3306) );
  NANDN U4481 ( .A(n3306), .B(n4642), .Z(n3307) );
  NAND U4482 ( .A(n3307), .B(n4644), .Z(n3308) );
  NAND U4483 ( .A(n3308), .B(n4646), .Z(n3309) );
  NAND U4484 ( .A(n3309), .B(n4649), .Z(n3310) );
  NAND U4485 ( .A(n3310), .B(n4650), .Z(n3311) );
  AND U4486 ( .A(n4652), .B(n3311), .Z(n3312) );
  NANDN U4487 ( .A(n3312), .B(n4654), .Z(n3313) );
  NAND U4488 ( .A(n3313), .B(n4656), .Z(n3314) );
  NAND U4489 ( .A(n3314), .B(n4658), .Z(n3315) );
  NAND U4490 ( .A(n3315), .B(n4661), .Z(n3316) );
  NAND U4491 ( .A(n3316), .B(n4662), .Z(n3317) );
  AND U4492 ( .A(n4664), .B(n3317), .Z(n3318) );
  NANDN U4493 ( .A(n3318), .B(n4666), .Z(n3319) );
  NAND U4494 ( .A(n3319), .B(n4668), .Z(n3321) );
  NAND U4495 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U4496 ( .A(n3323), .B(n3322), .Z(n3324) );
  NANDN U4497 ( .A(n3325), .B(n3324), .Z(n3327) );
  ANDN U4498 ( .B(n3327), .A(n3326), .Z(n3328) );
  NANDN U4499 ( .A(n3328), .B(n4674), .Z(n3329) );
  NAND U4500 ( .A(n3329), .B(n4676), .Z(n3330) );
  NAND U4501 ( .A(n3330), .B(n4678), .Z(n3331) );
  NAND U4502 ( .A(n3331), .B(n4680), .Z(n3332) );
  NAND U4503 ( .A(n3332), .B(n4682), .Z(n3333) );
  AND U4504 ( .A(n4685), .B(n3333), .Z(n3334) );
  NANDN U4505 ( .A(n3334), .B(n4686), .Z(n3335) );
  NAND U4506 ( .A(n3335), .B(n4688), .Z(n3336) );
  NAND U4507 ( .A(n3336), .B(n4690), .Z(n3337) );
  NAND U4508 ( .A(n3337), .B(n4692), .Z(n3338) );
  NAND U4509 ( .A(n3338), .B(n4694), .Z(n3339) );
  AND U4510 ( .A(n4697), .B(n3339), .Z(n3340) );
  NANDN U4511 ( .A(n3340), .B(n4698), .Z(n3341) );
  NAND U4512 ( .A(n3341), .B(n4700), .Z(n3342) );
  NAND U4513 ( .A(n3342), .B(n4702), .Z(n3343) );
  NANDN U4514 ( .A(n4705), .B(n3343), .Z(n3344) );
  NANDN U4515 ( .A(n4707), .B(n3344), .Z(n3345) );
  ANDN U4516 ( .B(n3345), .A(n4708), .Z(n3346) );
  NANDN U4517 ( .A(n3346), .B(n4710), .Z(n3347) );
  NANDN U4518 ( .A(n4713), .B(n3347), .Z(n3348) );
  NAND U4519 ( .A(n3348), .B(n4714), .Z(n3349) );
  NANDN U4520 ( .A(n4717), .B(n3349), .Z(n3350) );
  NAND U4521 ( .A(n3350), .B(n4718), .Z(n3351) );
  ANDN U4522 ( .B(n3351), .A(n4720), .Z(n3352) );
  NANDN U4523 ( .A(n3352), .B(n4722), .Z(n3353) );
  NANDN U4524 ( .A(n4724), .B(n3353), .Z(n3354) );
  NAND U4525 ( .A(n3354), .B(n4726), .Z(n3355) );
  NANDN U4526 ( .A(n4729), .B(n3355), .Z(n3356) );
  NANDN U4527 ( .A(n3357), .B(n3356), .Z(n3359) );
  ANDN U4528 ( .B(n3359), .A(n3358), .Z(n3360) );
  NANDN U4529 ( .A(n3360), .B(n4738), .Z(n3361) );
  NANDN U4530 ( .A(n4741), .B(n3361), .Z(n3362) );
  NAND U4531 ( .A(n3362), .B(n4742), .Z(n3363) );
  NANDN U4532 ( .A(n4745), .B(n3363), .Z(n3364) );
  NAND U4533 ( .A(n3364), .B(n4746), .Z(n3365) );
  ANDN U4534 ( .B(n3365), .A(n4748), .Z(n3366) );
  NANDN U4535 ( .A(n3366), .B(n4750), .Z(n3367) );
  ANDN U4536 ( .B(n3367), .A(n4753), .Z(n3368) );
  NANDN U4537 ( .A(n3368), .B(n4754), .Z(n3369) );
  NANDN U4538 ( .A(n4757), .B(n3369), .Z(n3371) );
  NAND U4539 ( .A(n3371), .B(n3370), .Z(n3372) );
  NAND U4540 ( .A(n3373), .B(n3372), .Z(n3374) );
  NANDN U4541 ( .A(n3375), .B(n3374), .Z(n3377) );
  ANDN U4542 ( .B(n3377), .A(n3376), .Z(n3378) );
  NANDN U4543 ( .A(n3378), .B(n4762), .Z(n3379) );
  NANDN U4544 ( .A(n4765), .B(n3379), .Z(n3380) );
  NAND U4545 ( .A(n3380), .B(n4766), .Z(n3381) );
  NANDN U4546 ( .A(n4769), .B(n3381), .Z(n3382) );
  NAND U4547 ( .A(n3382), .B(n4770), .Z(n3383) );
  ANDN U4548 ( .B(n3383), .A(n4772), .Z(n3384) );
  NANDN U4549 ( .A(n3384), .B(n4774), .Z(n3385) );
  NANDN U4550 ( .A(n4777), .B(n3385), .Z(n3386) );
  NAND U4551 ( .A(n3386), .B(n4778), .Z(n3387) );
  NANDN U4552 ( .A(n4781), .B(n3387), .Z(n3388) );
  NAND U4553 ( .A(n3388), .B(n4782), .Z(n3389) );
  ANDN U4554 ( .B(n3389), .A(n4784), .Z(n3390) );
  NANDN U4555 ( .A(n3390), .B(n4786), .Z(n3391) );
  NANDN U4556 ( .A(n4789), .B(n3391), .Z(n3392) );
  NAND U4557 ( .A(n3392), .B(n4790), .Z(n3393) );
  NANDN U4558 ( .A(n4793), .B(n3393), .Z(n3394) );
  NAND U4559 ( .A(n3394), .B(n4794), .Z(n3395) );
  ANDN U4560 ( .B(n3395), .A(n4796), .Z(n3396) );
  NANDN U4561 ( .A(n3396), .B(n4798), .Z(n3397) );
  NANDN U4562 ( .A(n4800), .B(n3397), .Z(n3398) );
  NAND U4563 ( .A(n3398), .B(n4802), .Z(n3399) );
  NANDN U4564 ( .A(n4805), .B(n3399), .Z(n3400) );
  NANDN U4565 ( .A(n3401), .B(n3400), .Z(n3403) );
  ANDN U4566 ( .B(n3403), .A(n3402), .Z(n3404) );
  NANDN U4567 ( .A(n3404), .B(n4814), .Z(n3405) );
  NANDN U4568 ( .A(n4817), .B(n3405), .Z(n3406) );
  NAND U4569 ( .A(n3406), .B(n4818), .Z(n3407) );
  NANDN U4570 ( .A(n4821), .B(n3407), .Z(n3408) );
  NAND U4571 ( .A(n3408), .B(n4822), .Z(n3409) );
  ANDN U4572 ( .B(n3409), .A(n4825), .Z(n3410) );
  OR U4573 ( .A(n3411), .B(n3410), .Z(n3412) );
  NANDN U4574 ( .A(n3413), .B(n3412), .Z(n3414) );
  NAND U4575 ( .A(n3414), .B(n4831), .Z(n3415) );
  NANDN U4576 ( .A(n4835), .B(n3415), .Z(n3416) );
  NAND U4577 ( .A(n3416), .B(n4836), .Z(n3417) );
  ANDN U4578 ( .B(n3417), .A(n4839), .Z(n3418) );
  NANDN U4579 ( .A(n3418), .B(n4840), .Z(n3419) );
  NANDN U4580 ( .A(n4841), .B(n3419), .Z(n3420) );
  NAND U4581 ( .A(n3420), .B(n4842), .Z(n3421) );
  NANDN U4582 ( .A(n4843), .B(n3421), .Z(n3422) );
  NAND U4583 ( .A(n3422), .B(n4844), .Z(n3423) );
  ANDN U4584 ( .B(n3423), .A(n4845), .Z(n3424) );
  OR U4585 ( .A(n3425), .B(n3424), .Z(n3426) );
  NANDN U4586 ( .A(n3427), .B(n3426), .Z(n3428) );
  NAND U4587 ( .A(n3428), .B(n4849), .Z(n3429) );
  NANDN U4588 ( .A(n4850), .B(n3429), .Z(n3430) );
  NAND U4589 ( .A(n3430), .B(n4851), .Z(n3431) );
  ANDN U4590 ( .B(n3431), .A(n4852), .Z(n3432) );
  NANDN U4591 ( .A(n3432), .B(n4853), .Z(n3433) );
  NANDN U4592 ( .A(n4854), .B(n3433), .Z(n3435) );
  NAND U4593 ( .A(n3435), .B(n3434), .Z(n3436) );
  NANDN U4594 ( .A(n3437), .B(n3436), .Z(n3438) );
  NANDN U4595 ( .A(n3439), .B(n3438), .Z(n3440) );
  ANDN U4596 ( .B(n3440), .A(n4866), .Z(n3441) );
  NANDN U4597 ( .A(n3441), .B(n4867), .Z(n3442) );
  NANDN U4598 ( .A(n4870), .B(n3442), .Z(n3443) );
  NAND U4599 ( .A(n3443), .B(n4871), .Z(n3444) );
  NANDN U4600 ( .A(n4874), .B(n3444), .Z(n3446) );
  NAND U4601 ( .A(n3446), .B(n3445), .Z(n3447) );
  AND U4602 ( .A(n3448), .B(n3447), .Z(n3449) );
  ANDN U4603 ( .B(n4879), .A(n3449), .Z(n3453) );
  NANDN U4604 ( .A(n3451), .B(n3450), .Z(n3452) );
  NAND U4605 ( .A(n3453), .B(n3452), .Z(n3454) );
  NANDN U4606 ( .A(n4882), .B(n3454), .Z(n3455) );
  NAND U4607 ( .A(n3455), .B(n4883), .Z(n3456) );
  ANDN U4608 ( .B(n3456), .A(n4886), .Z(n3457) );
  NANDN U4609 ( .A(n3457), .B(n4888), .Z(n3458) );
  ANDN U4610 ( .B(n3458), .A(n4890), .Z(n3459) );
  NANDN U4611 ( .A(n3459), .B(n4891), .Z(n3460) );
  NANDN U4612 ( .A(n4894), .B(n3460), .Z(n3462) );
  NAND U4613 ( .A(n3462), .B(n3461), .Z(n3463) );
  NAND U4614 ( .A(n3464), .B(n3463), .Z(n3465) );
  NANDN U4615 ( .A(n3466), .B(n3465), .Z(n3468) );
  ANDN U4616 ( .B(n3468), .A(n3467), .Z(n3469) );
  NANDN U4617 ( .A(n3469), .B(n4900), .Z(n3470) );
  NANDN U4618 ( .A(n4902), .B(n3470), .Z(n3471) );
  NAND U4619 ( .A(n3471), .B(n4903), .Z(n3472) );
  NANDN U4620 ( .A(n4906), .B(n3472), .Z(n3473) );
  NAND U4621 ( .A(n3473), .B(n4907), .Z(n3474) );
  ANDN U4622 ( .B(n3474), .A(n4910), .Z(n3475) );
  NANDN U4623 ( .A(n3475), .B(n4912), .Z(n3476) );
  NANDN U4624 ( .A(n4914), .B(n3476), .Z(n3477) );
  NAND U4625 ( .A(n3477), .B(n4915), .Z(n3478) );
  NANDN U4626 ( .A(n4918), .B(n3478), .Z(n3479) );
  NAND U4627 ( .A(n3479), .B(n4919), .Z(n3480) );
  ANDN U4628 ( .B(n3480), .A(n4922), .Z(n3481) );
  NANDN U4629 ( .A(n3481), .B(n4924), .Z(n3482) );
  NANDN U4630 ( .A(n4926), .B(n3482), .Z(n3484) );
  NAND U4631 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U4632 ( .A(n3486), .B(n3485), .Z(n3487) );
  NANDN U4633 ( .A(n3488), .B(n3487), .Z(n3490) );
  ANDN U4634 ( .B(n3490), .A(n3489), .Z(n3491) );
  NANDN U4635 ( .A(n3491), .B(n4931), .Z(n3492) );
  NANDN U4636 ( .A(n4934), .B(n3492), .Z(n3493) );
  NAND U4637 ( .A(n3493), .B(n4936), .Z(n3494) );
  NANDN U4638 ( .A(n4938), .B(n3494), .Z(n3495) );
  NAND U4639 ( .A(n3495), .B(n4939), .Z(n3496) );
  ANDN U4640 ( .B(n3496), .A(n4942), .Z(n3497) );
  NANDN U4641 ( .A(n3497), .B(n4943), .Z(n3498) );
  NANDN U4642 ( .A(n4946), .B(n3498), .Z(n3499) );
  NAND U4643 ( .A(n3499), .B(n4948), .Z(n3500) );
  NANDN U4644 ( .A(n4950), .B(n3500), .Z(n3501) );
  NAND U4645 ( .A(n3501), .B(n4951), .Z(n3502) );
  ANDN U4646 ( .B(n3502), .A(n4954), .Z(n3503) );
  NANDN U4647 ( .A(n3503), .B(n4955), .Z(n3504) );
  NANDN U4648 ( .A(n4958), .B(n3504), .Z(n3505) );
  NAND U4649 ( .A(n3505), .B(n4960), .Z(n3506) );
  NANDN U4650 ( .A(n4962), .B(n3506), .Z(n3507) );
  NAND U4651 ( .A(n3507), .B(n4963), .Z(n3508) );
  ANDN U4652 ( .B(n3508), .A(n4966), .Z(n3509) );
  OR U4653 ( .A(n3510), .B(n3509), .Z(n3511) );
  NANDN U4654 ( .A(n3512), .B(n3511), .Z(n3513) );
  NAND U4655 ( .A(n3513), .B(n4975), .Z(n3514) );
  NANDN U4656 ( .A(n4978), .B(n3514), .Z(n3515) );
  NAND U4657 ( .A(n3515), .B(n4980), .Z(n3516) );
  ANDN U4658 ( .B(n3516), .A(n4982), .Z(n3517) );
  NANDN U4659 ( .A(n3517), .B(n4983), .Z(n3518) );
  NANDN U4660 ( .A(n4986), .B(n3518), .Z(n3519) );
  NANDN U4661 ( .A(n3520), .B(n3519), .Z(n3521) );
  NANDN U4662 ( .A(n3522), .B(n3521), .Z(n3523) );
  NAND U4663 ( .A(n3523), .B(n4995), .Z(n3524) );
  ANDN U4664 ( .B(n3524), .A(n4998), .Z(n3525) );
  NANDN U4665 ( .A(n3525), .B(n5000), .Z(n3526) );
  NANDN U4666 ( .A(n5001), .B(n3526), .Z(n3527) );
  NANDN U4667 ( .A(n5005), .B(n3527), .Z(n3528) );
  NANDN U4668 ( .A(n3529), .B(n3528), .Z(n3530) );
  NANDN U4669 ( .A(n3531), .B(n3530), .Z(n3533) );
  ANDN U4670 ( .B(n3533), .A(n3532), .Z(n3534) );
  NANDN U4671 ( .A(n3534), .B(n5015), .Z(n3535) );
  NANDN U4672 ( .A(n5018), .B(n3535), .Z(n3536) );
  NAND U4673 ( .A(n3536), .B(n5019), .Z(n3537) );
  NANDN U4674 ( .A(n5022), .B(n3537), .Z(n3538) );
  NAND U4675 ( .A(n3538), .B(n5023), .Z(n3539) );
  ANDN U4676 ( .B(n3539), .A(n5025), .Z(n3540) );
  NANDN U4677 ( .A(n3540), .B(n5027), .Z(n3541) );
  NANDN U4678 ( .A(n5030), .B(n3541), .Z(n3542) );
  NAND U4679 ( .A(n3542), .B(n5031), .Z(n3543) );
  NANDN U4680 ( .A(n5034), .B(n3543), .Z(n3544) );
  NAND U4681 ( .A(n3544), .B(n5035), .Z(n3545) );
  ANDN U4682 ( .B(n3545), .A(n5037), .Z(n3546) );
  ANDN U4683 ( .B(n5039), .A(n3546), .Z(n3548) );
  NAND U4684 ( .A(n3548), .B(n3547), .Z(n3549) );
  ANDN U4685 ( .B(n3549), .A(n5042), .Z(n3551) );
  NANDN U4686 ( .A(n3551), .B(n3550), .Z(n3552) );
  NANDN U4687 ( .A(n5046), .B(n3552), .Z(n3553) );
  NANDN U4688 ( .A(n5048), .B(n3553), .Z(n3554) );
  NAND U4689 ( .A(n3554), .B(n5050), .Z(n3555) );
  NAND U4690 ( .A(n3555), .B(n5051), .Z(n3556) );
  AND U4691 ( .A(n5053), .B(n3556), .Z(n3557) );
  NANDN U4692 ( .A(n3557), .B(n5056), .Z(n3558) );
  NAND U4693 ( .A(n3558), .B(n5057), .Z(n3559) );
  NAND U4694 ( .A(n3559), .B(n5059), .Z(n3560) );
  NAND U4695 ( .A(n3560), .B(n5061), .Z(n3561) );
  NAND U4696 ( .A(n3561), .B(n5063), .Z(n3562) );
  AND U4697 ( .A(n5065), .B(n3562), .Z(n3563) );
  NANDN U4698 ( .A(n3563), .B(n5068), .Z(n3564) );
  NAND U4699 ( .A(n3564), .B(n5069), .Z(n3565) );
  NAND U4700 ( .A(n3565), .B(n5071), .Z(n3566) );
  NAND U4701 ( .A(n3566), .B(n5073), .Z(n3567) );
  NAND U4702 ( .A(n3567), .B(n5075), .Z(n3568) );
  AND U4703 ( .A(n5077), .B(n3568), .Z(n3569) );
  NANDN U4704 ( .A(n3569), .B(n5080), .Z(n3570) );
  AND U4705 ( .A(n5081), .B(n3570), .Z(n3571) );
  NANDN U4706 ( .A(n3571), .B(n5083), .Z(n3572) );
  NAND U4707 ( .A(n3572), .B(n5085), .Z(n3574) );
  NAND U4708 ( .A(n3574), .B(n3573), .Z(n3575) );
  NAND U4709 ( .A(n3576), .B(n3575), .Z(n3577) );
  NANDN U4710 ( .A(n3578), .B(n3577), .Z(n3580) );
  ANDN U4711 ( .B(n3580), .A(n3579), .Z(n3581) );
  NANDN U4712 ( .A(n3581), .B(n5092), .Z(n3582) );
  NAND U4713 ( .A(n3582), .B(n5093), .Z(n3583) );
  NAND U4714 ( .A(n3583), .B(n5095), .Z(n3584) );
  NAND U4715 ( .A(n3584), .B(n5097), .Z(n3585) );
  NAND U4716 ( .A(n3585), .B(n5099), .Z(n3586) );
  AND U4717 ( .A(n5101), .B(n3586), .Z(n3587) );
  NANDN U4718 ( .A(n3587), .B(n5104), .Z(n3588) );
  NAND U4719 ( .A(n3588), .B(n5105), .Z(n3589) );
  NAND U4720 ( .A(n3589), .B(n5107), .Z(n3590) );
  NAND U4721 ( .A(n3590), .B(n5109), .Z(n3591) );
  NAND U4722 ( .A(n3591), .B(n5111), .Z(n3592) );
  AND U4723 ( .A(n5113), .B(n3592), .Z(n3593) );
  NANDN U4724 ( .A(n3593), .B(n5116), .Z(n3594) );
  NAND U4725 ( .A(n3594), .B(n5117), .Z(n3595) );
  NAND U4726 ( .A(n3595), .B(n5119), .Z(n3596) );
  NAND U4727 ( .A(n3596), .B(n5121), .Z(n3597) );
  NAND U4728 ( .A(n3597), .B(n5123), .Z(n3598) );
  AND U4729 ( .A(n5125), .B(n3598), .Z(n3599) );
  NANDN U4730 ( .A(n3599), .B(n5128), .Z(n3600) );
  NAND U4731 ( .A(n3600), .B(n5129), .Z(n3601) );
  NAND U4732 ( .A(n3601), .B(n5131), .Z(n3602) );
  NAND U4733 ( .A(n3602), .B(n5133), .Z(n3603) );
  NAND U4734 ( .A(n3603), .B(n5135), .Z(n3604) );
  AND U4735 ( .A(n5137), .B(n3604), .Z(n3605) );
  NANDN U4736 ( .A(n3605), .B(n5140), .Z(n3606) );
  NAND U4737 ( .A(n3606), .B(n5141), .Z(n3607) );
  NAND U4738 ( .A(n3607), .B(n5143), .Z(n3608) );
  NAND U4739 ( .A(n3608), .B(n5145), .Z(n3609) );
  NAND U4740 ( .A(n3609), .B(n5147), .Z(n3610) );
  AND U4741 ( .A(n5149), .B(n3610), .Z(n3611) );
  NANDN U4742 ( .A(n3611), .B(n5152), .Z(n3612) );
  NAND U4743 ( .A(n3612), .B(n5153), .Z(n3613) );
  NAND U4744 ( .A(n3613), .B(n5155), .Z(n3614) );
  NAND U4745 ( .A(n3614), .B(n5157), .Z(n3615) );
  NAND U4746 ( .A(n3615), .B(n5159), .Z(n3616) );
  AND U4747 ( .A(n5161), .B(n3616), .Z(n3617) );
  NANDN U4748 ( .A(n3617), .B(n5164), .Z(n3618) );
  AND U4749 ( .A(n5165), .B(n3618), .Z(n3619) );
  NANDN U4750 ( .A(n3619), .B(n5167), .Z(n3620) );
  NAND U4751 ( .A(n3620), .B(n5169), .Z(n3622) );
  NAND U4752 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U4753 ( .A(n3624), .B(n3623), .Z(n3625) );
  NANDN U4754 ( .A(n3626), .B(n3625), .Z(n3628) );
  ANDN U4755 ( .B(n3628), .A(n3627), .Z(n3629) );
  NANDN U4756 ( .A(n3629), .B(n5176), .Z(n3630) );
  NAND U4757 ( .A(n3630), .B(n5177), .Z(n3631) );
  ANDN U4758 ( .B(n3631), .A(n5180), .Z(n3632) );
  NANDN U4759 ( .A(n3632), .B(n5181), .Z(n3633) );
  NANDN U4760 ( .A(n5184), .B(n3633), .Z(n3634) );
  NAND U4761 ( .A(n3634), .B(n5185), .Z(n3636) );
  NANDN U4762 ( .A(n3636), .B(n3635), .Z(n3637) );
  NANDN U4763 ( .A(n5187), .B(n3637), .Z(n3638) );
  NANDN U4764 ( .A(n3639), .B(n3638), .Z(n3641) );
  ANDN U4765 ( .B(x[458]), .A(y[458]), .Z(n3640) );
  OR U4766 ( .A(n3641), .B(n3640), .Z(n3642) );
  NANDN U4767 ( .A(n5192), .B(n3642), .Z(n3644) );
  NAND U4768 ( .A(n3644), .B(n3643), .Z(n3645) );
  OR U4769 ( .A(n3646), .B(n3645), .Z(n3647) );
  NANDN U4770 ( .A(n3648), .B(n3647), .Z(n3649) );
  NANDN U4771 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND U4772 ( .A(n3651), .B(n5203), .Z(n3652) );
  NAND U4773 ( .A(n3652), .B(n5205), .Z(n3653) );
  ANDN U4774 ( .B(n3653), .A(n5208), .Z(n3654) );
  NANDN U4775 ( .A(n3654), .B(n5209), .Z(n3655) );
  NANDN U4776 ( .A(n5212), .B(n3655), .Z(n3656) );
  NAND U4777 ( .A(n3656), .B(n5214), .Z(n3657) );
  NANDN U4778 ( .A(n5216), .B(n3657), .Z(n3658) );
  NAND U4779 ( .A(n3658), .B(n5217), .Z(n3659) );
  ANDN U4780 ( .B(n3659), .A(n5220), .Z(n3660) );
  NANDN U4781 ( .A(n3660), .B(n5221), .Z(n3661) );
  NANDN U4782 ( .A(n5224), .B(n3661), .Z(n3662) );
  NAND U4783 ( .A(n3662), .B(n5226), .Z(n3663) );
  NANDN U4784 ( .A(n5228), .B(n3663), .Z(n3664) );
  NAND U4785 ( .A(n3664), .B(n5229), .Z(n3665) );
  ANDN U4786 ( .B(n3665), .A(n5232), .Z(n3666) );
  NANDN U4787 ( .A(n3666), .B(n5233), .Z(n3667) );
  NANDN U4788 ( .A(n5236), .B(n3667), .Z(n3668) );
  NAND U4789 ( .A(n3668), .B(n5238), .Z(n3669) );
  NANDN U4790 ( .A(n5240), .B(n3669), .Z(n3670) );
  NAND U4791 ( .A(n3670), .B(n5241), .Z(n3671) );
  ANDN U4792 ( .B(n3671), .A(n5244), .Z(n3672) );
  NANDN U4793 ( .A(n3672), .B(n5245), .Z(n3673) );
  NANDN U4794 ( .A(n5248), .B(n3673), .Z(n3674) );
  NAND U4795 ( .A(n3674), .B(n5250), .Z(n3675) );
  NANDN U4796 ( .A(n5252), .B(n3675), .Z(n3676) );
  NAND U4797 ( .A(n3676), .B(n5253), .Z(n3677) );
  ANDN U4798 ( .B(n3677), .A(n5256), .Z(n3678) );
  NANDN U4799 ( .A(n3678), .B(n5257), .Z(n3679) );
  NANDN U4800 ( .A(n5260), .B(n3679), .Z(n3680) );
  NAND U4801 ( .A(n3680), .B(n5262), .Z(n3681) );
  NANDN U4802 ( .A(n5264), .B(n3681), .Z(n3682) );
  NAND U4803 ( .A(n3682), .B(n5265), .Z(n3683) );
  ANDN U4804 ( .B(n3683), .A(n5268), .Z(n3684) );
  NANDN U4805 ( .A(n3684), .B(n5269), .Z(n3685) );
  NANDN U4806 ( .A(n5272), .B(n3685), .Z(n3686) );
  NAND U4807 ( .A(n3686), .B(n5274), .Z(n3687) );
  NANDN U4808 ( .A(n5276), .B(n3687), .Z(n3688) );
  NAND U4809 ( .A(n3688), .B(n5277), .Z(n3689) );
  ANDN U4810 ( .B(n3689), .A(n5280), .Z(n3690) );
  NANDN U4811 ( .A(n3690), .B(n5281), .Z(n3691) );
  NANDN U4812 ( .A(n3692), .B(n3691), .Z(n3694) );
  NAND U4813 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U4814 ( .A(n5287), .B(n3695), .Z(n3699) );
  NANDN U4815 ( .A(n3697), .B(n3696), .Z(n3698) );
  AND U4816 ( .A(n3699), .B(n3698), .Z(n3700) );
  NANDN U4817 ( .A(n3700), .B(n5289), .Z(n3701) );
  NANDN U4818 ( .A(n5292), .B(n3701), .Z(n3702) );
  NAND U4819 ( .A(n3702), .B(n5293), .Z(n3703) );
  NANDN U4820 ( .A(n5296), .B(n3703), .Z(n3704) );
  NAND U4821 ( .A(n3704), .B(n5298), .Z(n3705) );
  ANDN U4822 ( .B(n3705), .A(n5300), .Z(n3706) );
  NANDN U4823 ( .A(n3706), .B(n5301), .Z(n3707) );
  NANDN U4824 ( .A(n5304), .B(n3707), .Z(n3708) );
  NAND U4825 ( .A(n3708), .B(n5305), .Z(n3709) );
  NANDN U4826 ( .A(n5308), .B(n3709), .Z(n3710) );
  NAND U4827 ( .A(n3710), .B(n5310), .Z(n3711) );
  ANDN U4828 ( .B(n3711), .A(n5312), .Z(n3712) );
  NANDN U4829 ( .A(n3712), .B(n5313), .Z(n3713) );
  NANDN U4830 ( .A(n5316), .B(n3713), .Z(n3714) );
  NAND U4831 ( .A(n3714), .B(n5317), .Z(n3715) );
  NANDN U4832 ( .A(n5320), .B(n3715), .Z(n3716) );
  NAND U4833 ( .A(n3716), .B(n5322), .Z(n3717) );
  ANDN U4834 ( .B(n3717), .A(n5324), .Z(n3718) );
  NANDN U4835 ( .A(n3718), .B(n5325), .Z(n3719) );
  NANDN U4836 ( .A(n5328), .B(n3719), .Z(n3720) );
  NAND U4837 ( .A(n3720), .B(n5329), .Z(n3721) );
  NANDN U4838 ( .A(n5332), .B(n3721), .Z(n3722) );
  NAND U4839 ( .A(n3722), .B(n5334), .Z(n3723) );
  ANDN U4840 ( .B(n3723), .A(n5336), .Z(n3724) );
  NANDN U4841 ( .A(n3724), .B(n5337), .Z(n3725) );
  NANDN U4842 ( .A(n3726), .B(n3725), .Z(n3727) );
  NANDN U4843 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U4844 ( .A(n3729), .B(n5347), .Z(n3730) );
  NAND U4845 ( .A(n3730), .B(n5349), .Z(n3731) );
  ANDN U4846 ( .B(n3731), .A(n5352), .Z(n3732) );
  NANDN U4847 ( .A(n3732), .B(n5353), .Z(n3733) );
  NANDN U4848 ( .A(n5356), .B(n3733), .Z(n3734) );
  NAND U4849 ( .A(n3734), .B(n5358), .Z(n3735) );
  NANDN U4850 ( .A(n5360), .B(n3735), .Z(n3736) );
  NAND U4851 ( .A(n3736), .B(n5361), .Z(n3737) );
  ANDN U4852 ( .B(n3737), .A(n5364), .Z(n3738) );
  NANDN U4853 ( .A(n3738), .B(n5365), .Z(n3739) );
  NANDN U4854 ( .A(n5368), .B(n3739), .Z(n3740) );
  NAND U4855 ( .A(n3740), .B(n5370), .Z(n3741) );
  NANDN U4856 ( .A(n5372), .B(n3741), .Z(n3742) );
  NAND U4857 ( .A(n3742), .B(n5373), .Z(n3743) );
  ANDN U4858 ( .B(n3743), .A(n5376), .Z(n3744) );
  NANDN U4859 ( .A(n3744), .B(n5377), .Z(n3745) );
  NANDN U4860 ( .A(n5380), .B(n3745), .Z(n3746) );
  NAND U4861 ( .A(n3746), .B(n5382), .Z(n3747) );
  NANDN U4862 ( .A(n5384), .B(n3747), .Z(n3748) );
  NAND U4863 ( .A(n3748), .B(n5386), .Z(n3749) );
  ANDN U4864 ( .B(n3749), .A(n5388), .Z(n3750) );
  NANDN U4865 ( .A(n3750), .B(n5389), .Z(n3751) );
  NANDN U4866 ( .A(n3752), .B(n3751), .Z(n3753) );
  NANDN U4867 ( .A(n3754), .B(n3753), .Z(n3755) );
  NAND U4868 ( .A(n3755), .B(n5399), .Z(n3756) );
  NAND U4869 ( .A(n3756), .B(n5401), .Z(n3757) );
  ANDN U4870 ( .B(n3757), .A(n5404), .Z(n3758) );
  NANDN U4871 ( .A(n3758), .B(n5405), .Z(n3759) );
  NANDN U4872 ( .A(n5408), .B(n3759), .Z(n3760) );
  NAND U4873 ( .A(n3760), .B(n5410), .Z(n3761) );
  NANDN U4874 ( .A(n5412), .B(n3761), .Z(n3762) );
  NAND U4875 ( .A(n3762), .B(n5413), .Z(n3763) );
  ANDN U4876 ( .B(n3763), .A(n5416), .Z(n3764) );
  NANDN U4877 ( .A(n3764), .B(n5417), .Z(n3765) );
  NAND U4878 ( .A(n3765), .B(n5419), .Z(n3766) );
  NAND U4879 ( .A(n3766), .B(n5422), .Z(n3767) );
  NANDN U4880 ( .A(n5424), .B(n3767), .Z(n3768) );
  NAND U4881 ( .A(n3768), .B(n5425), .Z(n3769) );
  ANDN U4882 ( .B(n3769), .A(n5428), .Z(n3770) );
  NANDN U4883 ( .A(n3770), .B(n5429), .Z(n3771) );
  NANDN U4884 ( .A(n5432), .B(n3771), .Z(n3772) );
  NAND U4885 ( .A(n3772), .B(n5434), .Z(n3773) );
  NANDN U4886 ( .A(n5436), .B(n3773), .Z(n3774) );
  NAND U4887 ( .A(n3774), .B(n5437), .Z(n3775) );
  ANDN U4888 ( .B(n3775), .A(n5440), .Z(n3776) );
  NANDN U4889 ( .A(n3776), .B(n5441), .Z(n3778) );
  ANDN U4890 ( .B(n3778), .A(n3777), .Z(n3779) );
  NAND U4891 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4892 ( .A(n3782), .B(n3781), .Z(n3783) );
  NANDN U4893 ( .A(n5448), .B(n3783), .Z(n3784) );
  NAND U4894 ( .A(n3784), .B(n5450), .Z(n3785) );
  ANDN U4895 ( .B(n3785), .A(n5452), .Z(n3786) );
  NANDN U4896 ( .A(n3786), .B(n5453), .Z(n3787) );
  NANDN U4897 ( .A(n3788), .B(n3787), .Z(n3789) );
  NANDN U4898 ( .A(n3790), .B(n3789), .Z(n3791) );
  NAND U4899 ( .A(n3791), .B(n5463), .Z(n3792) );
  NAND U4900 ( .A(n3792), .B(n5465), .Z(n3793) );
  ANDN U4901 ( .B(n3793), .A(n5468), .Z(n3794) );
  NANDN U4902 ( .A(n3794), .B(n5469), .Z(n3795) );
  NANDN U4903 ( .A(n5472), .B(n3795), .Z(n3796) );
  NAND U4904 ( .A(n3796), .B(n5473), .Z(n3797) );
  NANDN U4905 ( .A(n5476), .B(n3797), .Z(n3798) );
  NAND U4906 ( .A(n3798), .B(n5477), .Z(n3799) );
  ANDN U4907 ( .B(n3799), .A(n5479), .Z(n3800) );
  NANDN U4908 ( .A(n3800), .B(n5481), .Z(n3801) );
  NANDN U4909 ( .A(n5484), .B(n3801), .Z(n3802) );
  NAND U4910 ( .A(n3802), .B(n5485), .Z(n3803) );
  NANDN U4911 ( .A(n5488), .B(n3803), .Z(n3804) );
  NAND U4912 ( .A(n3804), .B(n5489), .Z(n3805) );
  AND U4913 ( .A(n5492), .B(n3805), .Z(n3806) );
  OR U4914 ( .A(n5494), .B(n3806), .Z(n3807) );
  NANDN U4915 ( .A(n5496), .B(n3807), .Z(n3808) );
  NAND U4916 ( .A(n3808), .B(n5497), .Z(n3809) );
  NANDN U4917 ( .A(n5500), .B(n3809), .Z(n3810) );
  NAND U4918 ( .A(n3810), .B(n5501), .Z(n3811) );
  ANDN U4919 ( .B(n3811), .A(n5503), .Z(n3812) );
  NANDN U4920 ( .A(n3812), .B(n5505), .Z(n3813) );
  AND U4921 ( .A(n5507), .B(n3813), .Z(n3814) );
  NANDN U4922 ( .A(n3814), .B(n5509), .Z(n3815) );
  NANDN U4923 ( .A(n5512), .B(n3815), .Z(n3816) );
  NAND U4924 ( .A(n3816), .B(n5513), .Z(n3818) );
  NAND U4925 ( .A(n3818), .B(n3817), .Z(n3820) );
  NAND U4926 ( .A(n3820), .B(n3819), .Z(n3821) );
  AND U4927 ( .A(n5519), .B(n3821), .Z(n3822) );
  NAND U4928 ( .A(n3823), .B(n3822), .Z(n3824) );
  NAND U4929 ( .A(n3824), .B(n5521), .Z(n3825) );
  NANDN U4930 ( .A(n5524), .B(n3825), .Z(n3826) );
  NAND U4931 ( .A(n3826), .B(n5525), .Z(n3827) );
  ANDN U4932 ( .B(n3827), .A(n5527), .Z(n3828) );
  NANDN U4933 ( .A(n3828), .B(n5529), .Z(n3829) );
  NAND U4934 ( .A(n3829), .B(n5531), .Z(n3830) );
  NAND U4935 ( .A(n3830), .B(n5533), .Z(n3831) );
  NANDN U4936 ( .A(n5536), .B(n3831), .Z(n3832) );
  NAND U4937 ( .A(n3832), .B(n5537), .Z(n3833) );
  AND U4938 ( .A(n3834), .B(n3833), .Z(n3835) );
  OR U4939 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4940 ( .A(n3837), .B(n5545), .Z(n3838) );
  NAND U4941 ( .A(n3838), .B(n5547), .Z(n3839) );
  NAND U4942 ( .A(n3839), .B(n5550), .Z(n3840) );
  NAND U4943 ( .A(n3840), .B(n5551), .Z(n3841) );
  AND U4944 ( .A(n5553), .B(n3841), .Z(n3842) );
  NANDN U4945 ( .A(n3842), .B(n5555), .Z(n3843) );
  NAND U4946 ( .A(n3843), .B(n5557), .Z(n3844) );
  NAND U4947 ( .A(n3844), .B(n5559), .Z(n3845) );
  NAND U4948 ( .A(n3845), .B(n5562), .Z(n3846) );
  NAND U4949 ( .A(n3846), .B(n5563), .Z(n3847) );
  AND U4950 ( .A(n5565), .B(n3847), .Z(n3848) );
  NANDN U4951 ( .A(n3848), .B(n5567), .Z(n3849) );
  NAND U4952 ( .A(n3849), .B(n5569), .Z(n3850) );
  NAND U4953 ( .A(n3850), .B(n5571), .Z(n3851) );
  NANDN U4954 ( .A(n3852), .B(n3851), .Z(n3853) );
  NAND U4955 ( .A(n3853), .B(n5575), .Z(n3854) );
  AND U4956 ( .A(n5577), .B(n3854), .Z(n3855) );
  NAND U4957 ( .A(n3856), .B(n3855), .Z(n3857) );
  NAND U4958 ( .A(n3857), .B(n5579), .Z(n3858) );
  NAND U4959 ( .A(n3858), .B(n5581), .Z(n3859) );
  NAND U4960 ( .A(n3859), .B(n5583), .Z(n3860) );
  AND U4961 ( .A(n5586), .B(n3860), .Z(n3861) );
  NANDN U4962 ( .A(n3861), .B(n5587), .Z(n3862) );
  NAND U4963 ( .A(n3862), .B(n5589), .Z(n3863) );
  NAND U4964 ( .A(n3863), .B(n5591), .Z(n3864) );
  NAND U4965 ( .A(n3864), .B(n5593), .Z(n3865) );
  NAND U4966 ( .A(n3865), .B(n5595), .Z(n3866) );
  AND U4967 ( .A(n5598), .B(n3866), .Z(n3867) );
  NANDN U4968 ( .A(n3867), .B(n5599), .Z(n3868) );
  NAND U4969 ( .A(n3868), .B(n5601), .Z(n3869) );
  NAND U4970 ( .A(n3869), .B(n5603), .Z(n3870) );
  NAND U4971 ( .A(n3870), .B(n5605), .Z(n3871) );
  NAND U4972 ( .A(n3871), .B(n5607), .Z(n3872) );
  AND U4973 ( .A(n5610), .B(n3872), .Z(n3873) );
  NANDN U4974 ( .A(n3873), .B(n5611), .Z(n3874) );
  NAND U4975 ( .A(n3874), .B(n5613), .Z(n3875) );
  NAND U4976 ( .A(n3875), .B(n5615), .Z(n3876) );
  NAND U4977 ( .A(n3876), .B(n5617), .Z(n3877) );
  NAND U4978 ( .A(n3877), .B(n5619), .Z(n3878) );
  AND U4979 ( .A(n5622), .B(n3878), .Z(n3879) );
  NANDN U4980 ( .A(n3879), .B(n5623), .Z(n3880) );
  NAND U4981 ( .A(n3880), .B(n5625), .Z(n3881) );
  NAND U4982 ( .A(n3881), .B(n5627), .Z(n3882) );
  NAND U4983 ( .A(n3882), .B(n5629), .Z(n3883) );
  NAND U4984 ( .A(n3883), .B(n5631), .Z(n3884) );
  AND U4985 ( .A(n5634), .B(n3884), .Z(n3885) );
  NANDN U4986 ( .A(n3885), .B(n5635), .Z(n3886) );
  NANDN U4987 ( .A(n3887), .B(n3886), .Z(n3889) );
  NAND U4988 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U4989 ( .A(n5641), .B(n3890), .Z(n3894) );
  NANDN U4990 ( .A(n3892), .B(n3891), .Z(n3893) );
  AND U4991 ( .A(n3894), .B(n3893), .Z(n3895) );
  NANDN U4992 ( .A(n3895), .B(n5643), .Z(n3896) );
  NAND U4993 ( .A(n3896), .B(n5645), .Z(n3897) );
  NAND U4994 ( .A(n3897), .B(n5647), .Z(n3898) );
  NAND U4995 ( .A(n3898), .B(n5649), .Z(n3899) );
  NAND U4996 ( .A(n3899), .B(n5652), .Z(n3900) );
  AND U4997 ( .A(n5653), .B(n3900), .Z(n3901) );
  NANDN U4998 ( .A(n3901), .B(n5655), .Z(n3902) );
  NAND U4999 ( .A(n3902), .B(n5657), .Z(n3903) );
  NAND U5000 ( .A(n3903), .B(n5659), .Z(n3904) );
  NAND U5001 ( .A(n3904), .B(n5661), .Z(n3905) );
  NAND U5002 ( .A(n3905), .B(n5664), .Z(n3906) );
  AND U5003 ( .A(n5665), .B(n3906), .Z(n3907) );
  NANDN U5004 ( .A(n3907), .B(n5667), .Z(n3908) );
  NAND U5005 ( .A(n3908), .B(n5669), .Z(n3909) );
  NAND U5006 ( .A(n3909), .B(n5671), .Z(n3910) );
  NAND U5007 ( .A(n3910), .B(n5673), .Z(n3911) );
  NAND U5008 ( .A(n3911), .B(n5676), .Z(n3913) );
  ANDN U5009 ( .B(n3913), .A(n3912), .Z(n3915) );
  ANDN U5010 ( .B(x[696]), .A(y[696]), .Z(n3914) );
  OR U5011 ( .A(n3915), .B(n3914), .Z(n3916) );
  NANDN U5012 ( .A(n3917), .B(n3916), .Z(n3919) );
  NAND U5013 ( .A(n3919), .B(n3918), .Z(n3920) );
  NAND U5014 ( .A(n3920), .B(n5681), .Z(n3921) );
  NAND U5015 ( .A(n3921), .B(n5683), .Z(n3922) );
  AND U5016 ( .A(n5685), .B(n3922), .Z(n3923) );
  NANDN U5017 ( .A(n3923), .B(n5688), .Z(n3924) );
  NAND U5018 ( .A(n3924), .B(n5689), .Z(n3925) );
  NAND U5019 ( .A(n3925), .B(n5691), .Z(n3926) );
  NAND U5020 ( .A(n3926), .B(n5693), .Z(n3927) );
  NAND U5021 ( .A(n3927), .B(n5695), .Z(n3928) );
  AND U5022 ( .A(n5697), .B(n3928), .Z(n3929) );
  NANDN U5023 ( .A(n3929), .B(n5700), .Z(n3930) );
  NAND U5024 ( .A(n3930), .B(n5701), .Z(n3931) );
  NANDN U5025 ( .A(n5704), .B(n3931), .Z(n3932) );
  NANDN U5026 ( .A(n5706), .B(n3932), .Z(n3933) );
  NAND U5027 ( .A(n3933), .B(n5707), .Z(n3934) );
  ANDN U5028 ( .B(n3934), .A(n5710), .Z(n3935) );
  NANDN U5029 ( .A(n3935), .B(n5712), .Z(n3936) );
  NANDN U5030 ( .A(n5714), .B(n3936), .Z(n3937) );
  NAND U5031 ( .A(n3937), .B(n5716), .Z(n3938) );
  NANDN U5032 ( .A(n5718), .B(n3938), .Z(n3939) );
  NAND U5033 ( .A(n3939), .B(n5719), .Z(n3941) );
  ANDN U5034 ( .B(n3941), .A(n3940), .Z(n3942) );
  OR U5035 ( .A(n3943), .B(n3942), .Z(n3944) );
  NAND U5036 ( .A(n3944), .B(n5729), .Z(n3945) );
  NAND U5037 ( .A(n3945), .B(n5731), .Z(n3946) );
  NANDN U5038 ( .A(n5733), .B(n3946), .Z(n3947) );
  NAND U5039 ( .A(n3947), .B(n5735), .Z(n3948) );
  ANDN U5040 ( .B(n3948), .A(n5738), .Z(n3949) );
  OR U5041 ( .A(n5740), .B(n3949), .Z(n3950) );
  NANDN U5042 ( .A(n5742), .B(n3950), .Z(n3951) );
  NAND U5043 ( .A(n3951), .B(n5743), .Z(n3952) );
  NAND U5044 ( .A(n3952), .B(n5746), .Z(n3953) );
  NAND U5045 ( .A(n3953), .B(n5747), .Z(n3954) );
  ANDN U5046 ( .B(n3954), .A(n5750), .Z(n3955) );
  NANDN U5047 ( .A(n3955), .B(n5751), .Z(n3956) );
  NANDN U5048 ( .A(n5754), .B(n3956), .Z(n3957) );
  NAND U5049 ( .A(n3957), .B(n5755), .Z(n3958) );
  NANDN U5050 ( .A(n5757), .B(n3958), .Z(n3959) );
  NAND U5051 ( .A(n3959), .B(n5759), .Z(n3960) );
  ANDN U5052 ( .B(n3960), .A(n5762), .Z(n3961) );
  NANDN U5053 ( .A(n3961), .B(n5763), .Z(n3962) );
  NANDN U5054 ( .A(n5766), .B(n3962), .Z(n3963) );
  NAND U5055 ( .A(n3963), .B(n5767), .Z(n3964) );
  NANDN U5056 ( .A(n5769), .B(n3964), .Z(n3965) );
  NAND U5057 ( .A(n3965), .B(n5771), .Z(n3967) );
  ANDN U5058 ( .B(n3967), .A(n3966), .Z(n3968) );
  OR U5059 ( .A(n3969), .B(n3968), .Z(n3970) );
  NAND U5060 ( .A(n3970), .B(n5778), .Z(n3971) );
  NAND U5061 ( .A(n3971), .B(n5783), .Z(n3972) );
  NANDN U5062 ( .A(n5786), .B(n3972), .Z(n3973) );
  NAND U5063 ( .A(n3973), .B(n5787), .Z(n3974) );
  ANDN U5064 ( .B(n3974), .A(n5790), .Z(n3975) );
  NANDN U5065 ( .A(n3975), .B(n5791), .Z(n3976) );
  NANDN U5066 ( .A(n3977), .B(n3976), .Z(n3978) );
  NANDN U5067 ( .A(n3979), .B(n3978), .Z(n3980) );
  NAND U5068 ( .A(n3980), .B(n5801), .Z(n3981) );
  NAND U5069 ( .A(n3981), .B(n5803), .Z(n3983) );
  ANDN U5070 ( .B(n3983), .A(n3982), .Z(n3984) );
  OR U5071 ( .A(n3985), .B(n3984), .Z(n3986) );
  NAND U5072 ( .A(n3986), .B(n5813), .Z(n3987) );
  NAND U5073 ( .A(n3987), .B(n5815), .Z(n3988) );
  NANDN U5074 ( .A(n5817), .B(n3988), .Z(n3989) );
  NAND U5075 ( .A(n3989), .B(n5819), .Z(n3990) );
  ANDN U5076 ( .B(n3990), .A(n5822), .Z(n3991) );
  NANDN U5077 ( .A(n3991), .B(n5823), .Z(n3992) );
  NANDN U5078 ( .A(n5826), .B(n3992), .Z(n3993) );
  NAND U5079 ( .A(n3993), .B(n5827), .Z(n3994) );
  NANDN U5080 ( .A(n5829), .B(n3994), .Z(n3995) );
  NAND U5081 ( .A(n3995), .B(n5831), .Z(n3996) );
  ANDN U5082 ( .B(n3996), .A(n5834), .Z(n3997) );
  NANDN U5083 ( .A(n3997), .B(n5835), .Z(n3998) );
  NAND U5084 ( .A(n3998), .B(n5839), .Z(n3999) );
  NANDN U5085 ( .A(n4000), .B(n3999), .Z(n4001) );
  NAND U5086 ( .A(n4001), .B(n5843), .Z(n4002) );
  NAND U5087 ( .A(n4002), .B(n5845), .Z(n4003) );
  ANDN U5088 ( .B(n4003), .A(n5847), .Z(n4004) );
  NANDN U5089 ( .A(n4004), .B(n5849), .Z(n4005) );
  NANDN U5090 ( .A(n5852), .B(n4005), .Z(n4006) );
  NAND U5091 ( .A(n4006), .B(n5853), .Z(n4007) );
  NANDN U5092 ( .A(n5856), .B(n4007), .Z(n4008) );
  NAND U5093 ( .A(n4008), .B(n5859), .Z(n4009) );
  AND U5094 ( .A(n5861), .B(n4009), .Z(n4010) );
  OR U5095 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U5096 ( .A(n4012), .B(n5865), .Z(n4013) );
  NAND U5097 ( .A(n4013), .B(n5867), .Z(n4014) );
  NANDN U5098 ( .A(n5870), .B(n4014), .Z(n4015) );
  NAND U5099 ( .A(n4015), .B(n5872), .Z(n4016) );
  ANDN U5100 ( .B(n4016), .A(n5874), .Z(n4017) );
  NANDN U5101 ( .A(n4017), .B(n5875), .Z(n4018) );
  NANDN U5102 ( .A(n5878), .B(n4018), .Z(n4019) );
  NAND U5103 ( .A(n4019), .B(n5879), .Z(n4020) );
  NANDN U5104 ( .A(n5882), .B(n4020), .Z(n4021) );
  NAND U5105 ( .A(n4021), .B(n5884), .Z(n4022) );
  ANDN U5106 ( .B(n4022), .A(n5886), .Z(n4023) );
  NANDN U5107 ( .A(n4023), .B(n5887), .Z(n4024) );
  NANDN U5108 ( .A(n5890), .B(n4024), .Z(n4025) );
  NAND U5109 ( .A(n4025), .B(n5891), .Z(n4026) );
  NANDN U5110 ( .A(n5894), .B(n4026), .Z(n4027) );
  NAND U5111 ( .A(n4027), .B(n5896), .Z(n4028) );
  ANDN U5112 ( .B(n4028), .A(n5898), .Z(n4029) );
  NANDN U5113 ( .A(n4029), .B(n5899), .Z(n4030) );
  NANDN U5114 ( .A(n4031), .B(n4030), .Z(n4032) );
  NANDN U5115 ( .A(n4033), .B(n4032), .Z(n4034) );
  AND U5116 ( .A(n5905), .B(n4034), .Z(n4038) );
  NANDN U5117 ( .A(n4036), .B(n4035), .Z(n4037) );
  AND U5118 ( .A(n4038), .B(n4037), .Z(n4039) );
  NANDN U5119 ( .A(n4039), .B(n5908), .Z(n4040) );
  NANDN U5120 ( .A(n4041), .B(n4040), .Z(n4042) );
  NANDN U5121 ( .A(n4043), .B(n4042), .Z(n4045) );
  ANDN U5122 ( .B(x[808]), .A(y[808]), .Z(n4044) );
  OR U5123 ( .A(n4045), .B(n4044), .Z(n4046) );
  NAND U5124 ( .A(n4046), .B(n5913), .Z(n4048) );
  NAND U5125 ( .A(n4048), .B(n4047), .Z(n4049) );
  NAND U5126 ( .A(n4049), .B(n5921), .Z(n4050) );
  NAND U5127 ( .A(n4050), .B(n5923), .Z(n4051) );
  AND U5128 ( .A(n5926), .B(n4051), .Z(n4052) );
  NANDN U5129 ( .A(n4052), .B(n5927), .Z(n4053) );
  NAND U5130 ( .A(n4053), .B(n5929), .Z(n4054) );
  NAND U5131 ( .A(n4054), .B(n5931), .Z(n4055) );
  NAND U5132 ( .A(n4055), .B(n5933), .Z(n4056) );
  NAND U5133 ( .A(n4056), .B(n5935), .Z(n4057) );
  AND U5134 ( .A(n5938), .B(n4057), .Z(n4058) );
  NANDN U5135 ( .A(n4058), .B(n5939), .Z(n4059) );
  NAND U5136 ( .A(n4059), .B(n5941), .Z(n4060) );
  NAND U5137 ( .A(n4060), .B(n5943), .Z(n4061) );
  NAND U5138 ( .A(n4061), .B(n5945), .Z(n4062) );
  NAND U5139 ( .A(n4062), .B(n5947), .Z(n4063) );
  AND U5140 ( .A(n5950), .B(n4063), .Z(n4064) );
  NANDN U5141 ( .A(n4064), .B(n5951), .Z(n4065) );
  NAND U5142 ( .A(n4065), .B(n5953), .Z(n4066) );
  NAND U5143 ( .A(n4066), .B(n5955), .Z(n4067) );
  NAND U5144 ( .A(n4067), .B(n5957), .Z(n4068) );
  NAND U5145 ( .A(n4068), .B(n5959), .Z(n4069) );
  AND U5146 ( .A(n5962), .B(n4069), .Z(n4070) );
  NANDN U5147 ( .A(n4070), .B(n5963), .Z(n4071) );
  NAND U5148 ( .A(n4071), .B(n5965), .Z(n4072) );
  NAND U5149 ( .A(n4072), .B(n5967), .Z(n4073) );
  NAND U5150 ( .A(n4073), .B(n5969), .Z(n4074) );
  NAND U5151 ( .A(n4074), .B(n5971), .Z(n4075) );
  AND U5152 ( .A(n5974), .B(n4075), .Z(n4076) );
  NANDN U5153 ( .A(n4076), .B(n5975), .Z(n4077) );
  NAND U5154 ( .A(n4077), .B(n5977), .Z(n4078) );
  NAND U5155 ( .A(n4078), .B(n5979), .Z(n4079) );
  NAND U5156 ( .A(n4079), .B(n5981), .Z(n4080) );
  NAND U5157 ( .A(n4080), .B(n5983), .Z(n4081) );
  AND U5158 ( .A(n5986), .B(n4081), .Z(n4082) );
  NANDN U5159 ( .A(n4082), .B(n5987), .Z(n4083) );
  NAND U5160 ( .A(n4083), .B(n5989), .Z(n4084) );
  NAND U5161 ( .A(n4084), .B(n5991), .Z(n4085) );
  NAND U5162 ( .A(n4085), .B(n5993), .Z(n4086) );
  NAND U5163 ( .A(n4086), .B(n5995), .Z(n4087) );
  AND U5164 ( .A(n5998), .B(n4087), .Z(n4088) );
  ANDN U5165 ( .B(n5999), .A(n4088), .Z(n4090) );
  NAND U5166 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U5167 ( .A(n6001), .B(n4091), .Z(n4092) );
  NAND U5168 ( .A(n4093), .B(n4092), .Z(n4094) );
  NAND U5169 ( .A(n4095), .B(n4094), .Z(n4096) );
  NAND U5170 ( .A(n4097), .B(n4096), .Z(n4098) );
  NAND U5171 ( .A(n4098), .B(n6011), .Z(n4099) );
  NAND U5172 ( .A(n4099), .B(n6013), .Z(n4100) );
  NAND U5173 ( .A(n4100), .B(n6015), .Z(n4101) );
  AND U5174 ( .A(n6017), .B(n4101), .Z(n4102) );
  NANDN U5175 ( .A(n4102), .B(n6019), .Z(n4103) );
  NAND U5176 ( .A(n4103), .B(n6023), .Z(n4104) );
  NANDN U5177 ( .A(n6026), .B(n4104), .Z(n4106) );
  NAND U5178 ( .A(n4106), .B(n4105), .Z(n4107) );
  AND U5179 ( .A(n4108), .B(n4107), .Z(n4109) );
  NAND U5180 ( .A(n4109), .B(n6029), .Z(n4110) );
  NAND U5181 ( .A(n4110), .B(n4363), .Z(n4111) );
  NAND U5182 ( .A(n4112), .B(n4111), .Z(n4113) );
  NAND U5183 ( .A(n4114), .B(n4113), .Z(n4115) );
  NAND U5184 ( .A(n4115), .B(n6037), .Z(n4116) );
  AND U5185 ( .A(n4117), .B(n4116), .Z(n4118) );
  NAND U5186 ( .A(n4118), .B(n6039), .Z(n4119) );
  NANDN U5187 ( .A(n6042), .B(n4119), .Z(n4120) );
  NAND U5188 ( .A(n4120), .B(n6044), .Z(n4121) );
  ANDN U5189 ( .B(n4121), .A(n6046), .Z(n4122) );
  NANDN U5190 ( .A(n4122), .B(n6047), .Z(n4123) );
  NANDN U5191 ( .A(n6050), .B(n4123), .Z(n4124) );
  NAND U5192 ( .A(n4124), .B(n6053), .Z(n4125) );
  NAND U5193 ( .A(n4125), .B(n6055), .Z(n4126) );
  AND U5194 ( .A(n6059), .B(n4126), .Z(n4127) );
  NANDN U5195 ( .A(n4128), .B(n4127), .Z(n4129) );
  NAND U5196 ( .A(n4130), .B(n4129), .Z(n4131) );
  NANDN U5197 ( .A(n6064), .B(n4131), .Z(n4139) );
  NANDN U5198 ( .A(n4133), .B(n4132), .Z(n4137) );
  XOR U5199 ( .A(x[875]), .B(n4133), .Z(n4134) );
  NANDN U5200 ( .A(n4135), .B(n4134), .Z(n4136) );
  NAND U5201 ( .A(n4137), .B(n4136), .Z(n4138) );
  AND U5202 ( .A(n4139), .B(n4138), .Z(n4140) );
  NANDN U5203 ( .A(n4140), .B(n6068), .Z(n4141) );
  NAND U5204 ( .A(n4141), .B(n6069), .Z(n4142) );
  NAND U5205 ( .A(n4142), .B(n6071), .Z(n4143) );
  NAND U5206 ( .A(n4143), .B(n6073), .Z(n4144) );
  NAND U5207 ( .A(n4144), .B(n6075), .Z(n4145) );
  AND U5208 ( .A(n6077), .B(n4145), .Z(n4146) );
  NANDN U5209 ( .A(n4146), .B(n6081), .Z(n4147) );
  NAND U5210 ( .A(n4147), .B(n6083), .Z(n4148) );
  NANDN U5211 ( .A(n4149), .B(n4148), .Z(n4151) );
  NANDN U5212 ( .A(n4151), .B(n4150), .Z(n4152) );
  NAND U5213 ( .A(n4152), .B(n6087), .Z(n4154) );
  OR U5214 ( .A(n4154), .B(n4153), .Z(n4157) );
  XNOR U5215 ( .A(n4154), .B(y[885]), .Z(n4155) );
  NANDN U5216 ( .A(x[885]), .B(n4155), .Z(n4156) );
  NAND U5217 ( .A(n4157), .B(n4156), .Z(n4158) );
  NANDN U5218 ( .A(n4158), .B(n6093), .Z(n4159) );
  NANDN U5219 ( .A(n4160), .B(n4159), .Z(n4161) );
  NAND U5220 ( .A(n4161), .B(n6098), .Z(n4162) );
  NAND U5221 ( .A(n4162), .B(n6099), .Z(n4163) );
  NAND U5222 ( .A(n4163), .B(n6101), .Z(n4164) );
  AND U5223 ( .A(n6103), .B(n4164), .Z(n4165) );
  NANDN U5224 ( .A(n4165), .B(n6105), .Z(n4166) );
  NANDN U5225 ( .A(n6108), .B(n4166), .Z(n4167) );
  NAND U5226 ( .A(n4167), .B(n6109), .Z(n4168) );
  NAND U5227 ( .A(n4168), .B(n6111), .Z(n4169) );
  NAND U5228 ( .A(n4169), .B(n6113), .Z(n4170) );
  ANDN U5229 ( .B(n4170), .A(n6115), .Z(n4171) );
  NANDN U5230 ( .A(n4171), .B(n6117), .Z(n4172) );
  NANDN U5231 ( .A(n6120), .B(n4172), .Z(n4173) );
  NAND U5232 ( .A(n4173), .B(n6121), .Z(n4174) );
  NAND U5233 ( .A(n4174), .B(n6123), .Z(n4175) );
  NAND U5234 ( .A(n4175), .B(n6125), .Z(n4176) );
  ANDN U5235 ( .B(n4176), .A(n6127), .Z(n4177) );
  NANDN U5236 ( .A(n4177), .B(n6129), .Z(n4178) );
  NANDN U5237 ( .A(n6132), .B(n4178), .Z(n4179) );
  NAND U5238 ( .A(n4179), .B(n6133), .Z(n4180) );
  NANDN U5239 ( .A(n6136), .B(n4180), .Z(n4181) );
  NAND U5240 ( .A(n4181), .B(n6138), .Z(n4182) );
  ANDN U5241 ( .B(n4182), .A(n6142), .Z(n4184) );
  NANDN U5242 ( .A(n4184), .B(n4183), .Z(n4185) );
  NAND U5243 ( .A(n4185), .B(n6149), .Z(n4186) );
  AND U5244 ( .A(n6151), .B(n4186), .Z(n4187) );
  NANDN U5245 ( .A(n4187), .B(n6153), .Z(n4188) );
  NAND U5246 ( .A(n4188), .B(n6155), .Z(n4189) );
  NAND U5247 ( .A(n4189), .B(n6158), .Z(n4190) );
  NAND U5248 ( .A(n4190), .B(n6159), .Z(n4191) );
  NAND U5249 ( .A(n4191), .B(n6161), .Z(n4192) );
  AND U5250 ( .A(n6163), .B(n4192), .Z(n4193) );
  NANDN U5251 ( .A(n4193), .B(n6165), .Z(n4194) );
  AND U5252 ( .A(n6168), .B(n4194), .Z(n4195) );
  NANDN U5253 ( .A(n4195), .B(n6172), .Z(n4197) );
  NAND U5254 ( .A(n4197), .B(n4196), .Z(n4198) );
  NANDN U5255 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U5256 ( .A(n4200), .B(n6179), .Z(n4201) );
  NANDN U5257 ( .A(n6182), .B(n4201), .Z(n4203) );
  NAND U5258 ( .A(n4203), .B(n4202), .Z(n4204) );
  NAND U5259 ( .A(n4204), .B(n6185), .Z(n4205) );
  AND U5260 ( .A(n4206), .B(n4205), .Z(n4207) );
  NAND U5261 ( .A(n4207), .B(n6187), .Z(n4208) );
  NANDN U5262 ( .A(n6189), .B(n4208), .Z(n4209) );
  NAND U5263 ( .A(n4209), .B(n6191), .Z(n4210) );
  ANDN U5264 ( .B(n4210), .A(n6194), .Z(n4211) );
  NANDN U5265 ( .A(n4211), .B(n6195), .Z(n4212) );
  NAND U5266 ( .A(n4212), .B(n6197), .Z(n4213) );
  NAND U5267 ( .A(n4213), .B(n6201), .Z(n4214) );
  NAND U5268 ( .A(n4214), .B(n6204), .Z(n4215) );
  AND U5269 ( .A(n6207), .B(n4215), .Z(n4216) );
  NANDN U5270 ( .A(n4217), .B(n4216), .Z(n4218) );
  NANDN U5271 ( .A(n6210), .B(n4218), .Z(n4219) );
  AND U5272 ( .A(n6211), .B(n4219), .Z(n4221) );
  NAND U5273 ( .A(n4221), .B(n4220), .Z(n4222) );
  AND U5274 ( .A(n6218), .B(n4222), .Z(n4223) );
  NAND U5275 ( .A(n4223), .B(n6213), .Z(n4225) );
  ANDN U5276 ( .B(n4225), .A(n4224), .Z(n4226) );
  NAND U5277 ( .A(n4226), .B(n6219), .Z(n4227) );
  NAND U5278 ( .A(n4227), .B(n6221), .Z(n4228) );
  ANDN U5279 ( .B(n4228), .A(n6224), .Z(n4229) );
  NANDN U5280 ( .A(n4229), .B(n6225), .Z(n4230) );
  NANDN U5281 ( .A(n6228), .B(n4230), .Z(n4231) );
  NAND U5282 ( .A(n4231), .B(n6230), .Z(n4232) );
  NAND U5283 ( .A(n4232), .B(n6232), .Z(n4233) );
  NAND U5284 ( .A(n4233), .B(n6236), .Z(n4235) );
  ANDN U5285 ( .B(n4235), .A(n4234), .Z(n4236) );
  ANDN U5286 ( .B(n6239), .A(n4236), .Z(n4238) );
  NAND U5287 ( .A(n4238), .B(n4237), .Z(n4239) );
  AND U5288 ( .A(n6241), .B(n4239), .Z(n4240) );
  NAND U5289 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND U5290 ( .A(n4243), .B(n4242), .Z(n4244) );
  NAND U5291 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U5292 ( .A(n6251), .B(n4246), .Z(n4247) );
  NANDN U5293 ( .A(n4247), .B(n6253), .Z(n4248) );
  NAND U5294 ( .A(n4248), .B(n6255), .Z(n4249) );
  NAND U5295 ( .A(n4249), .B(n6257), .Z(n4250) );
  NAND U5296 ( .A(n4250), .B(n6260), .Z(n4251) );
  NAND U5297 ( .A(n4251), .B(n6261), .Z(n4252) );
  AND U5298 ( .A(n6263), .B(n4252), .Z(n4253) );
  NANDN U5299 ( .A(n4253), .B(n6265), .Z(n4254) );
  NAND U5300 ( .A(n4254), .B(n6267), .Z(n4255) );
  NAND U5301 ( .A(n4255), .B(n6269), .Z(n4256) );
  NAND U5302 ( .A(n4256), .B(n6272), .Z(n4257) );
  NAND U5303 ( .A(n4257), .B(n6273), .Z(n4258) );
  AND U5304 ( .A(n6275), .B(n4258), .Z(n4259) );
  NANDN U5305 ( .A(n4259), .B(n6277), .Z(n4260) );
  NAND U5306 ( .A(n4260), .B(n6279), .Z(n4261) );
  NAND U5307 ( .A(n4261), .B(n6281), .Z(n4262) );
  NAND U5308 ( .A(n4262), .B(n6284), .Z(n4263) );
  NAND U5309 ( .A(n4263), .B(n6285), .Z(n4264) );
  AND U5310 ( .A(n6287), .B(n4264), .Z(n4265) );
  NANDN U5311 ( .A(n4265), .B(n6289), .Z(n4266) );
  NAND U5312 ( .A(n4266), .B(n6291), .Z(n4267) );
  NAND U5313 ( .A(n4267), .B(n6293), .Z(n4268) );
  NAND U5314 ( .A(n4268), .B(n6296), .Z(n4269) );
  NAND U5315 ( .A(n4269), .B(n6297), .Z(n4270) );
  AND U5316 ( .A(n6299), .B(n4270), .Z(n4271) );
  NANDN U5317 ( .A(n4271), .B(n6301), .Z(n4272) );
  NAND U5318 ( .A(n4272), .B(n6303), .Z(n4273) );
  NAND U5319 ( .A(n4273), .B(n6305), .Z(n4274) );
  NAND U5320 ( .A(n4274), .B(n6308), .Z(n4275) );
  NAND U5321 ( .A(n4275), .B(n6309), .Z(n4276) );
  AND U5322 ( .A(n6311), .B(n4276), .Z(n4277) );
  NANDN U5323 ( .A(n4277), .B(n6313), .Z(n4278) );
  NAND U5324 ( .A(n4278), .B(n6315), .Z(n4279) );
  NAND U5325 ( .A(n4279), .B(n6318), .Z(n4280) );
  NAND U5326 ( .A(n4280), .B(n6321), .Z(n4281) );
  AND U5327 ( .A(n4282), .B(n4281), .Z(n4283) );
  NANDN U5328 ( .A(n4284), .B(n4283), .Z(n4285) );
  AND U5329 ( .A(n4285), .B(n6326), .Z(n4286) );
  OR U5330 ( .A(n4286), .B(y[981]), .Z(n4289) );
  XOR U5331 ( .A(y[981]), .B(n4286), .Z(n4287) );
  NAND U5332 ( .A(n4287), .B(x[981]), .Z(n4288) );
  NAND U5333 ( .A(n4289), .B(n4288), .Z(n4291) );
  ANDN U5334 ( .B(n4291), .A(n4290), .Z(n4292) );
  ANDN U5335 ( .B(n6334), .A(n4292), .Z(n4294) );
  NAND U5336 ( .A(n4294), .B(n4293), .Z(n4296) );
  ANDN U5337 ( .B(n4296), .A(n4295), .Z(n4297) );
  NAND U5338 ( .A(n4297), .B(n6335), .Z(n4298) );
  NAND U5339 ( .A(n4298), .B(n6338), .Z(n4299) );
  ANDN U5340 ( .B(n4299), .A(n6340), .Z(n4300) );
  NANDN U5341 ( .A(n4300), .B(n6341), .Z(n4301) );
  NANDN U5342 ( .A(n6344), .B(n4301), .Z(n4302) );
  NAND U5343 ( .A(n4302), .B(n6345), .Z(n4304) );
  AND U5344 ( .A(n4304), .B(n4303), .Z(n4305) );
  OR U5345 ( .A(n4305), .B(x[990]), .Z(n4308) );
  XOR U5346 ( .A(x[990]), .B(n4305), .Z(n4306) );
  NAND U5347 ( .A(n4306), .B(y[990]), .Z(n4307) );
  NAND U5348 ( .A(n4308), .B(n4307), .Z(n4309) );
  ANDN U5349 ( .B(x[991]), .A(y[991]), .Z(n4359) );
  ANDN U5350 ( .B(n4309), .A(n4359), .Z(n4312) );
  NOR U5351 ( .A(n4311), .B(n4310), .Z(n6351) );
  NANDN U5352 ( .A(n4312), .B(n6351), .Z(n4313) );
  AND U5353 ( .A(n4314), .B(n4313), .Z(n4315) );
  NAND U5354 ( .A(n4316), .B(n4315), .Z(n4317) );
  NAND U5355 ( .A(n4318), .B(n4317), .Z(n4319) );
  AND U5356 ( .A(n6359), .B(n4319), .Z(n4320) );
  ANDN U5357 ( .B(n6361), .A(n4320), .Z(n4322) );
  NAND U5358 ( .A(n4322), .B(n4321), .Z(n4323) );
  ANDN U5359 ( .B(n4323), .A(n6364), .Z(n4324) );
  NANDN U5360 ( .A(n4324), .B(n6366), .Z(n4325) );
  ANDN U5361 ( .B(n4325), .A(n6368), .Z(n4326) );
  NANDN U5362 ( .A(n4326), .B(n6369), .Z(n4327) );
  NANDN U5363 ( .A(n6372), .B(n4327), .Z(n4328) );
  NAND U5364 ( .A(n4328), .B(n6375), .Z(n4329) );
  NAND U5365 ( .A(n4329), .B(n4356), .Z(n4330) );
  NANDN U5366 ( .A(n4331), .B(n4330), .Z(n4332) );
  AND U5367 ( .A(n4357), .B(n4332), .Z(n4333) );
  NANDN U5368 ( .A(n4333), .B(n6381), .Z(n4336) );
  NANDN U5369 ( .A(y[1004]), .B(x[1004]), .Z(n4335) );
  NAND U5370 ( .A(n4335), .B(n4334), .Z(n6384) );
  ANDN U5371 ( .B(n4336), .A(n6384), .Z(n4338) );
  NOR U5372 ( .A(n4338), .B(n4337), .Z(n4339) );
  NAND U5373 ( .A(n4339), .B(n6386), .Z(n4341) );
  AND U5374 ( .A(n4341), .B(n4340), .Z(n4342) );
  OR U5375 ( .A(n4342), .B(y[1007]), .Z(n4345) );
  XOR U5376 ( .A(y[1007]), .B(n4342), .Z(n4343) );
  NAND U5377 ( .A(n4343), .B(x[1007]), .Z(n4344) );
  NAND U5378 ( .A(n4345), .B(n4344), .Z(n4346) );
  AND U5379 ( .A(n6393), .B(n4346), .Z(n4347) );
  NANDN U5380 ( .A(n4347), .B(n6395), .Z(n4348) );
  NAND U5381 ( .A(n4348), .B(n6398), .Z(n4349) );
  NAND U5382 ( .A(n4349), .B(n6399), .Z(n4350) );
  NANDN U5383 ( .A(n6402), .B(n4350), .Z(n4351) );
  NANDN U5384 ( .A(n6404), .B(n4351), .Z(n4352) );
  AND U5385 ( .A(n6405), .B(n4352), .Z(n4353) );
  ANDN U5386 ( .B(n4354), .A(n4353), .Z(n4355) );
  NANDN U5387 ( .A(ebreg), .B(n4355), .Z(n5) );
  OR U5388 ( .A(n4355), .B(ebreg), .Z(n6428) );
  ANDN U5389 ( .B(x[1007]), .A(y[1007]), .Z(n6392) );
  NAND U5390 ( .A(n4357), .B(n4356), .Z(n6378) );
  NANDN U5391 ( .A(n4359), .B(n4358), .Z(n6350) );
  ANDN U5392 ( .B(n4361), .A(n4360), .Z(n6348) );
  XNOR U5393 ( .A(y[919]), .B(x[919]), .Z(n6174) );
  ANDN U5394 ( .B(n4363), .A(n4362), .Z(n6032) );
  ANDN U5395 ( .B(x[758]), .A(y[758]), .Z(n5808) );
  ANDN U5396 ( .B(n4365), .A(n4364), .Z(n5544) );
  XNOR U5397 ( .A(x[628]), .B(y[628]), .Z(n5542) );
  ANDN U5398 ( .B(n4367), .A(n4366), .Z(n5014) );
  XOR U5399 ( .A(n4368), .B(x[368]), .Z(n5012) );
  XNOR U5400 ( .A(x[295]), .B(y[295]), .Z(n4860) );
  NAND U5401 ( .A(n4371), .B(n4370), .Z(n4833) );
  XOR U5402 ( .A(n4372), .B(y[166]), .Z(n4598) );
  ANDN U5403 ( .B(n4374), .A(n4373), .Z(n4570) );
  XNOR U5404 ( .A(x[152]), .B(y[152]), .Z(n4568) );
  ANDN U5405 ( .B(n4376), .A(n4375), .Z(n4530) );
  XNOR U5406 ( .A(x[134]), .B(y[134]), .Z(n4528) );
  ANDN U5407 ( .B(x[124]), .A(y[124]), .Z(n4504) );
  ANDN U5408 ( .B(x[100]), .A(y[100]), .Z(n4450) );
  ANDN U5409 ( .B(x[86]), .A(y[86]), .Z(n4418) );
  ANDN U5410 ( .B(x[68]), .A(y[68]), .Z(n4377) );
  OR U5411 ( .A(n4378), .B(n4377), .Z(n4380) );
  NAND U5412 ( .A(n4380), .B(n4379), .Z(n4381) );
  NANDN U5413 ( .A(n4382), .B(n4381), .Z(n4384) );
  NAND U5414 ( .A(n4384), .B(n4383), .Z(n4386) );
  NAND U5415 ( .A(n4386), .B(n4385), .Z(n4388) );
  ANDN U5416 ( .B(n4388), .A(n4387), .Z(n4390) );
  NANDN U5417 ( .A(n4390), .B(n4389), .Z(n4391) );
  NANDN U5418 ( .A(n4392), .B(n4391), .Z(n4394) );
  NAND U5419 ( .A(n4394), .B(n4393), .Z(n4395) );
  NANDN U5420 ( .A(n4396), .B(n4395), .Z(n4398) );
  NAND U5421 ( .A(n4398), .B(n4397), .Z(n4400) );
  ANDN U5422 ( .B(n4400), .A(n4399), .Z(n4402) );
  NANDN U5423 ( .A(n4402), .B(n4401), .Z(n4403) );
  NANDN U5424 ( .A(n4404), .B(n4403), .Z(n4406) );
  NAND U5425 ( .A(n4406), .B(n4405), .Z(n4407) );
  NANDN U5426 ( .A(n4408), .B(n4407), .Z(n4410) );
  NAND U5427 ( .A(n4410), .B(n4409), .Z(n4412) );
  ANDN U5428 ( .B(n4412), .A(n4411), .Z(n4414) );
  NANDN U5429 ( .A(n4414), .B(n4413), .Z(n4416) );
  ANDN U5430 ( .B(n4416), .A(n4415), .Z(n4417) );
  OR U5431 ( .A(n4418), .B(n4417), .Z(n4419) );
  NANDN U5432 ( .A(n4420), .B(n4419), .Z(n4421) );
  NANDN U5433 ( .A(n4422), .B(n4421), .Z(n4424) );
  NAND U5434 ( .A(n4424), .B(n4423), .Z(n4426) );
  NAND U5435 ( .A(n4426), .B(n4425), .Z(n4428) );
  ANDN U5436 ( .B(n4428), .A(n4427), .Z(n4430) );
  NANDN U5437 ( .A(n4430), .B(n4429), .Z(n4431) );
  NANDN U5438 ( .A(n4432), .B(n4431), .Z(n4434) );
  NAND U5439 ( .A(n4434), .B(n4433), .Z(n4435) );
  NANDN U5440 ( .A(n4436), .B(n4435), .Z(n4438) );
  NAND U5441 ( .A(n4438), .B(n4437), .Z(n4440) );
  ANDN U5442 ( .B(n4440), .A(n4439), .Z(n4442) );
  NANDN U5443 ( .A(n4442), .B(n4441), .Z(n4443) );
  NANDN U5444 ( .A(n4444), .B(n4443), .Z(n4446) );
  NAND U5445 ( .A(n4446), .B(n4445), .Z(n4448) );
  ANDN U5446 ( .B(n4448), .A(n4447), .Z(n4449) );
  OR U5447 ( .A(n4450), .B(n4449), .Z(n4451) );
  NANDN U5448 ( .A(n4452), .B(n4451), .Z(n4453) );
  NANDN U5449 ( .A(n4454), .B(n4453), .Z(n4456) );
  OR U5450 ( .A(n4456), .B(n4455), .Z(n4457) );
  NANDN U5451 ( .A(n4458), .B(n4457), .Z(n4460) );
  NAND U5452 ( .A(n4460), .B(n4459), .Z(n4461) );
  NANDN U5453 ( .A(n4462), .B(n4461), .Z(n4464) );
  NAND U5454 ( .A(n4464), .B(n4463), .Z(n4466) );
  ANDN U5455 ( .B(n4466), .A(n4465), .Z(n4468) );
  NANDN U5456 ( .A(n4468), .B(n4467), .Z(n4469) );
  NANDN U5457 ( .A(n4470), .B(n4469), .Z(n4472) );
  NAND U5458 ( .A(n4472), .B(n4471), .Z(n4473) );
  NANDN U5459 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U5460 ( .A(n4476), .B(n4475), .Z(n4477) );
  NANDN U5461 ( .A(n4478), .B(n4477), .Z(n4480) );
  ANDN U5462 ( .B(n4480), .A(n4479), .Z(n4482) );
  NANDN U5463 ( .A(n4482), .B(n4481), .Z(n4484) );
  NAND U5464 ( .A(n4484), .B(n4483), .Z(n4485) );
  NANDN U5465 ( .A(n4486), .B(n4485), .Z(n4488) );
  NAND U5466 ( .A(n4488), .B(n4487), .Z(n4489) );
  NANDN U5467 ( .A(n4490), .B(n4489), .Z(n4491) );
  AND U5468 ( .A(n4492), .B(n4491), .Z(n4494) );
  NANDN U5469 ( .A(n4494), .B(n4493), .Z(n4495) );
  NANDN U5470 ( .A(n4496), .B(n4495), .Z(n4497) );
  NANDN U5471 ( .A(n4498), .B(n4497), .Z(n4500) );
  NAND U5472 ( .A(n4500), .B(n4499), .Z(n4502) );
  ANDN U5473 ( .B(n4502), .A(n4501), .Z(n4503) );
  OR U5474 ( .A(n4504), .B(n4503), .Z(n4505) );
  NANDN U5475 ( .A(n4506), .B(n4505), .Z(n4507) );
  NANDN U5476 ( .A(n4508), .B(n4507), .Z(n4510) );
  NAND U5477 ( .A(n4510), .B(n4509), .Z(n4512) );
  NAND U5478 ( .A(n4512), .B(n4511), .Z(n4514) );
  ANDN U5479 ( .B(n4514), .A(n4513), .Z(n4515) );
  OR U5480 ( .A(n4516), .B(n4515), .Z(n4518) );
  NAND U5481 ( .A(n4518), .B(n4517), .Z(n4520) );
  NAND U5482 ( .A(n4520), .B(n4519), .Z(n4521) );
  NANDN U5483 ( .A(n4522), .B(n4521), .Z(n4524) );
  NAND U5484 ( .A(n4524), .B(n4523), .Z(n4526) );
  ANDN U5485 ( .B(n4526), .A(n4525), .Z(n4527) );
  NAND U5486 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U5487 ( .A(n4530), .B(n4529), .Z(n4531) );
  NANDN U5488 ( .A(n4532), .B(n4531), .Z(n4534) );
  NAND U5489 ( .A(n4534), .B(n4533), .Z(n4536) );
  ANDN U5490 ( .B(n4536), .A(n4535), .Z(n4538) );
  NANDN U5491 ( .A(n4538), .B(n4537), .Z(n4539) );
  NANDN U5492 ( .A(n4540), .B(n4539), .Z(n4541) );
  NANDN U5493 ( .A(n4542), .B(n4541), .Z(n4543) );
  OR U5494 ( .A(n4544), .B(n4543), .Z(n4546) );
  NAND U5495 ( .A(n4546), .B(n4545), .Z(n4547) );
  NANDN U5496 ( .A(n4548), .B(n4547), .Z(n4550) );
  NAND U5497 ( .A(n4550), .B(n4549), .Z(n4552) );
  NAND U5498 ( .A(n4552), .B(n4551), .Z(n4553) );
  AND U5499 ( .A(n4554), .B(n4553), .Z(n4556) );
  NANDN U5500 ( .A(n4556), .B(n4555), .Z(n4558) );
  NAND U5501 ( .A(n4558), .B(n4557), .Z(n4560) );
  NAND U5502 ( .A(n4560), .B(n4559), .Z(n4562) );
  NAND U5503 ( .A(n4562), .B(n4561), .Z(n4564) );
  NAND U5504 ( .A(n4564), .B(n4563), .Z(n4566) );
  ANDN U5505 ( .B(n4566), .A(n4565), .Z(n4567) );
  NAND U5506 ( .A(n4568), .B(n4567), .Z(n4569) );
  NAND U5507 ( .A(n4570), .B(n4569), .Z(n4572) );
  NAND U5508 ( .A(n4572), .B(n4571), .Z(n4573) );
  NANDN U5509 ( .A(n4574), .B(n4573), .Z(n4575) );
  AND U5510 ( .A(n4576), .B(n4575), .Z(n4578) );
  NANDN U5511 ( .A(n4578), .B(n4577), .Z(n4580) );
  NAND U5512 ( .A(n4580), .B(n4579), .Z(n4582) );
  NAND U5513 ( .A(n4582), .B(n4581), .Z(n4583) );
  NANDN U5514 ( .A(n4584), .B(n4583), .Z(n4586) );
  NAND U5515 ( .A(n4586), .B(n4585), .Z(n4588) );
  ANDN U5516 ( .B(n4588), .A(n4587), .Z(n4589) );
  OR U5517 ( .A(n4590), .B(n4589), .Z(n4592) );
  NAND U5518 ( .A(n4592), .B(n4591), .Z(n4594) );
  NAND U5519 ( .A(n4594), .B(n4593), .Z(n4595) );
  NANDN U5520 ( .A(n4596), .B(n4595), .Z(n4597) );
  NAND U5521 ( .A(n4598), .B(n4597), .Z(n4599) );
  AND U5522 ( .A(n4600), .B(n4599), .Z(n4603) );
  OR U5523 ( .A(n4603), .B(x[167]), .Z(n4602) );
  ANDN U5524 ( .B(n4602), .A(n4601), .Z(n4607) );
  XNOR U5525 ( .A(n4604), .B(n4603), .Z(n4605) );
  NAND U5526 ( .A(y[167]), .B(n4605), .Z(n4606) );
  NAND U5527 ( .A(n4607), .B(n4606), .Z(n4609) );
  NAND U5528 ( .A(n4609), .B(n4608), .Z(n4611) );
  NAND U5529 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5530 ( .A(n4613), .B(n4612), .Z(n4615) );
  NANDN U5531 ( .A(n4615), .B(n4614), .Z(n4617) );
  NAND U5532 ( .A(n4617), .B(n4616), .Z(n4619) );
  NAND U5533 ( .A(n4619), .B(n4618), .Z(n4620) );
  NANDN U5534 ( .A(n4621), .B(n4620), .Z(n4622) );
  NANDN U5535 ( .A(n4623), .B(n4622), .Z(n4624) );
  AND U5536 ( .A(n4625), .B(n4624), .Z(n4626) );
  OR U5537 ( .A(n4627), .B(n4626), .Z(n4628) );
  NANDN U5538 ( .A(n4629), .B(n4628), .Z(n4631) );
  NAND U5539 ( .A(n4631), .B(n4630), .Z(n4633) );
  NAND U5540 ( .A(n4633), .B(n4632), .Z(n4635) );
  NAND U5541 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U5542 ( .A(n4637), .B(n4636), .Z(n4639) );
  NANDN U5543 ( .A(n4639), .B(n4638), .Z(n4641) );
  NAND U5544 ( .A(n4641), .B(n4640), .Z(n4643) );
  NAND U5545 ( .A(n4643), .B(n4642), .Z(n4645) );
  NAND U5546 ( .A(n4645), .B(n4644), .Z(n4647) );
  NAND U5547 ( .A(n4647), .B(n4646), .Z(n4648) );
  AND U5548 ( .A(n4649), .B(n4648), .Z(n4651) );
  NANDN U5549 ( .A(n4651), .B(n4650), .Z(n4653) );
  NAND U5550 ( .A(n4653), .B(n4652), .Z(n4655) );
  NAND U5551 ( .A(n4655), .B(n4654), .Z(n4657) );
  NAND U5552 ( .A(n4657), .B(n4656), .Z(n4659) );
  NAND U5553 ( .A(n4659), .B(n4658), .Z(n4660) );
  AND U5554 ( .A(n4661), .B(n4660), .Z(n4663) );
  NANDN U5555 ( .A(n4663), .B(n4662), .Z(n4665) );
  NAND U5556 ( .A(n4665), .B(n4664), .Z(n4667) );
  NAND U5557 ( .A(n4667), .B(n4666), .Z(n4669) );
  NAND U5558 ( .A(n4669), .B(n4668), .Z(n4670) );
  NANDN U5559 ( .A(n4671), .B(n4670), .Z(n4672) );
  AND U5560 ( .A(n4673), .B(n4672), .Z(n4675) );
  NANDN U5561 ( .A(n4675), .B(n4674), .Z(n4677) );
  NAND U5562 ( .A(n4677), .B(n4676), .Z(n4679) );
  NAND U5563 ( .A(n4679), .B(n4678), .Z(n4681) );
  NAND U5564 ( .A(n4681), .B(n4680), .Z(n4683) );
  NAND U5565 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U5566 ( .A(n4685), .B(n4684), .Z(n4687) );
  NANDN U5567 ( .A(n4687), .B(n4686), .Z(n4689) );
  NAND U5568 ( .A(n4689), .B(n4688), .Z(n4691) );
  NAND U5569 ( .A(n4691), .B(n4690), .Z(n4693) );
  NAND U5570 ( .A(n4693), .B(n4692), .Z(n4695) );
  NAND U5571 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U5572 ( .A(n4697), .B(n4696), .Z(n4699) );
  NANDN U5573 ( .A(n4699), .B(n4698), .Z(n4701) );
  NAND U5574 ( .A(n4701), .B(n4700), .Z(n4703) );
  NAND U5575 ( .A(n4703), .B(n4702), .Z(n4704) );
  NANDN U5576 ( .A(n4705), .B(n4704), .Z(n4706) );
  NANDN U5577 ( .A(n4707), .B(n4706), .Z(n4709) );
  ANDN U5578 ( .B(n4709), .A(n4708), .Z(n4711) );
  NANDN U5579 ( .A(n4711), .B(n4710), .Z(n4712) );
  NANDN U5580 ( .A(n4713), .B(n4712), .Z(n4715) );
  NAND U5581 ( .A(n4715), .B(n4714), .Z(n4716) );
  NANDN U5582 ( .A(n4717), .B(n4716), .Z(n4719) );
  NAND U5583 ( .A(n4719), .B(n4718), .Z(n4721) );
  ANDN U5584 ( .B(n4721), .A(n4720), .Z(n4723) );
  NANDN U5585 ( .A(n4723), .B(n4722), .Z(n4725) );
  ANDN U5586 ( .B(n4725), .A(n4724), .Z(n4727) );
  NANDN U5587 ( .A(n4727), .B(n4726), .Z(n4728) );
  NANDN U5588 ( .A(n4729), .B(n4728), .Z(n4730) );
  NANDN U5589 ( .A(n4731), .B(n4730), .Z(n4733) );
  NAND U5590 ( .A(n4733), .B(n4732), .Z(n4734) );
  NANDN U5591 ( .A(n4735), .B(n4734), .Z(n4737) );
  ANDN U5592 ( .B(n4737), .A(n4736), .Z(n4739) );
  NANDN U5593 ( .A(n4739), .B(n4738), .Z(n4740) );
  NANDN U5594 ( .A(n4741), .B(n4740), .Z(n4743) );
  NAND U5595 ( .A(n4743), .B(n4742), .Z(n4744) );
  NANDN U5596 ( .A(n4745), .B(n4744), .Z(n4747) );
  NAND U5597 ( .A(n4747), .B(n4746), .Z(n4749) );
  ANDN U5598 ( .B(n4749), .A(n4748), .Z(n4751) );
  NANDN U5599 ( .A(n4751), .B(n4750), .Z(n4752) );
  NANDN U5600 ( .A(n4753), .B(n4752), .Z(n4755) );
  NAND U5601 ( .A(n4755), .B(n4754), .Z(n4756) );
  NANDN U5602 ( .A(n4757), .B(n4756), .Z(n4758) );
  NANDN U5603 ( .A(n4759), .B(n4758), .Z(n4761) );
  ANDN U5604 ( .B(n4761), .A(n4760), .Z(n4763) );
  NANDN U5605 ( .A(n4763), .B(n4762), .Z(n4764) );
  NANDN U5606 ( .A(n4765), .B(n4764), .Z(n4767) );
  NAND U5607 ( .A(n4767), .B(n4766), .Z(n4768) );
  NANDN U5608 ( .A(n4769), .B(n4768), .Z(n4771) );
  NAND U5609 ( .A(n4771), .B(n4770), .Z(n4773) );
  ANDN U5610 ( .B(n4773), .A(n4772), .Z(n4775) );
  NANDN U5611 ( .A(n4775), .B(n4774), .Z(n4776) );
  NANDN U5612 ( .A(n4777), .B(n4776), .Z(n4779) );
  NAND U5613 ( .A(n4779), .B(n4778), .Z(n4780) );
  NANDN U5614 ( .A(n4781), .B(n4780), .Z(n4783) );
  NAND U5615 ( .A(n4783), .B(n4782), .Z(n4785) );
  ANDN U5616 ( .B(n4785), .A(n4784), .Z(n4787) );
  NANDN U5617 ( .A(n4787), .B(n4786), .Z(n4788) );
  NANDN U5618 ( .A(n4789), .B(n4788), .Z(n4791) );
  NAND U5619 ( .A(n4791), .B(n4790), .Z(n4792) );
  NANDN U5620 ( .A(n4793), .B(n4792), .Z(n4795) );
  NAND U5621 ( .A(n4795), .B(n4794), .Z(n4797) );
  ANDN U5622 ( .B(n4797), .A(n4796), .Z(n4799) );
  NANDN U5623 ( .A(n4799), .B(n4798), .Z(n4801) );
  ANDN U5624 ( .B(n4801), .A(n4800), .Z(n4803) );
  NANDN U5625 ( .A(n4803), .B(n4802), .Z(n4804) );
  NANDN U5626 ( .A(n4805), .B(n4804), .Z(n4806) );
  NANDN U5627 ( .A(n4807), .B(n4806), .Z(n4809) );
  NAND U5628 ( .A(n4809), .B(n4808), .Z(n4810) );
  NANDN U5629 ( .A(n4811), .B(n4810), .Z(n4813) );
  ANDN U5630 ( .B(n4813), .A(n4812), .Z(n4815) );
  NANDN U5631 ( .A(n4815), .B(n4814), .Z(n4816) );
  NANDN U5632 ( .A(n4817), .B(n4816), .Z(n4819) );
  NAND U5633 ( .A(n4819), .B(n4818), .Z(n4820) );
  NANDN U5634 ( .A(n4821), .B(n4820), .Z(n4823) );
  NAND U5635 ( .A(n4823), .B(n4822), .Z(n4824) );
  NANDN U5636 ( .A(n4825), .B(n4824), .Z(n4826) );
  NANDN U5637 ( .A(n4827), .B(n4826), .Z(n4828) );
  NANDN U5638 ( .A(n4829), .B(n4828), .Z(n4830) );
  AND U5639 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U5640 ( .A(n4833), .B(n4832), .Z(n4834) );
  NANDN U5641 ( .A(n4835), .B(n4834), .Z(n4837) );
  NAND U5642 ( .A(n4837), .B(n4836), .Z(n4838) );
  NANDN U5643 ( .A(n4855), .B(x[294]), .Z(n4858) );
  XNOR U5644 ( .A(n4855), .B(x[294]), .Z(n4856) );
  NANDN U5645 ( .A(y[294]), .B(n4856), .Z(n4857) );
  NAND U5646 ( .A(n4858), .B(n4857), .Z(n4859) );
  NAND U5647 ( .A(n4860), .B(n4859), .Z(n4861) );
  NAND U5648 ( .A(n4862), .B(n4861), .Z(n4864) );
  ANDN U5649 ( .B(n4864), .A(n4863), .Z(n4865) );
  OR U5650 ( .A(n4866), .B(n4865), .Z(n4868) );
  NAND U5651 ( .A(n4868), .B(n4867), .Z(n4869) );
  NANDN U5652 ( .A(n4870), .B(n4869), .Z(n4872) );
  NAND U5653 ( .A(n4872), .B(n4871), .Z(n4873) );
  NANDN U5654 ( .A(n4874), .B(n4873), .Z(n4876) );
  ANDN U5655 ( .B(n4876), .A(n4875), .Z(n4877) );
  OR U5656 ( .A(n4878), .B(n4877), .Z(n4880) );
  NAND U5657 ( .A(n4880), .B(n4879), .Z(n4881) );
  NANDN U5658 ( .A(n4882), .B(n4881), .Z(n4884) );
  NAND U5659 ( .A(n4884), .B(n4883), .Z(n4885) );
  NANDN U5660 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5661 ( .A(n4888), .B(n4887), .Z(n4889) );
  OR U5662 ( .A(n4890), .B(n4889), .Z(n4892) );
  NAND U5663 ( .A(n4892), .B(n4891), .Z(n4893) );
  NANDN U5664 ( .A(n4894), .B(n4893), .Z(n4895) );
  NANDN U5665 ( .A(n4896), .B(n4895), .Z(n4897) );
  NANDN U5666 ( .A(n4898), .B(n4897), .Z(n4899) );
  AND U5667 ( .A(n4900), .B(n4899), .Z(n4901) );
  OR U5668 ( .A(n4902), .B(n4901), .Z(n4904) );
  NAND U5669 ( .A(n4904), .B(n4903), .Z(n4905) );
  NANDN U5670 ( .A(n4906), .B(n4905), .Z(n4908) );
  NAND U5671 ( .A(n4908), .B(n4907), .Z(n4909) );
  NANDN U5672 ( .A(n4910), .B(n4909), .Z(n4911) );
  AND U5673 ( .A(n4912), .B(n4911), .Z(n4913) );
  OR U5674 ( .A(n4914), .B(n4913), .Z(n4916) );
  NAND U5675 ( .A(n4916), .B(n4915), .Z(n4917) );
  NANDN U5676 ( .A(n4918), .B(n4917), .Z(n4920) );
  NAND U5677 ( .A(n4920), .B(n4919), .Z(n4921) );
  NANDN U5678 ( .A(n4922), .B(n4921), .Z(n4923) );
  AND U5679 ( .A(n4924), .B(n4923), .Z(n4925) );
  OR U5680 ( .A(n4926), .B(n4925), .Z(n4927) );
  NANDN U5681 ( .A(n4928), .B(n4927), .Z(n4929) );
  NANDN U5682 ( .A(n4930), .B(n4929), .Z(n4932) );
  NAND U5683 ( .A(n4932), .B(n4931), .Z(n4933) );
  NANDN U5684 ( .A(n4934), .B(n4933), .Z(n4935) );
  AND U5685 ( .A(n4936), .B(n4935), .Z(n4937) );
  OR U5686 ( .A(n4938), .B(n4937), .Z(n4940) );
  NAND U5687 ( .A(n4940), .B(n4939), .Z(n4941) );
  NANDN U5688 ( .A(n4942), .B(n4941), .Z(n4944) );
  NAND U5689 ( .A(n4944), .B(n4943), .Z(n4945) );
  NANDN U5690 ( .A(n4946), .B(n4945), .Z(n4947) );
  AND U5691 ( .A(n4948), .B(n4947), .Z(n4949) );
  OR U5692 ( .A(n4950), .B(n4949), .Z(n4952) );
  NAND U5693 ( .A(n4952), .B(n4951), .Z(n4953) );
  NANDN U5694 ( .A(n4954), .B(n4953), .Z(n4956) );
  NAND U5695 ( .A(n4956), .B(n4955), .Z(n4957) );
  NANDN U5696 ( .A(n4958), .B(n4957), .Z(n4959) );
  AND U5697 ( .A(n4960), .B(n4959), .Z(n4961) );
  OR U5698 ( .A(n4962), .B(n4961), .Z(n4964) );
  NAND U5699 ( .A(n4964), .B(n4963), .Z(n4965) );
  NANDN U5700 ( .A(n4966), .B(n4965), .Z(n4967) );
  NANDN U5701 ( .A(n4968), .B(n4967), .Z(n4970) );
  NAND U5702 ( .A(n4970), .B(n4969), .Z(n4971) );
  NANDN U5703 ( .A(n4972), .B(n4971), .Z(n4974) );
  ANDN U5704 ( .B(n4974), .A(n4973), .Z(n4976) );
  NANDN U5705 ( .A(n4976), .B(n4975), .Z(n4977) );
  NANDN U5706 ( .A(n4978), .B(n4977), .Z(n4979) );
  AND U5707 ( .A(n4980), .B(n4979), .Z(n4981) );
  OR U5708 ( .A(n4982), .B(n4981), .Z(n4984) );
  NAND U5709 ( .A(n4984), .B(n4983), .Z(n4985) );
  NANDN U5710 ( .A(n4986), .B(n4985), .Z(n4987) );
  NANDN U5711 ( .A(n4988), .B(n4987), .Z(n4990) );
  NAND U5712 ( .A(n4990), .B(n4989), .Z(n4991) );
  NANDN U5713 ( .A(n4992), .B(n4991), .Z(n4994) );
  ANDN U5714 ( .B(n4994), .A(n4993), .Z(n4996) );
  NANDN U5715 ( .A(n4996), .B(n4995), .Z(n4997) );
  NANDN U5716 ( .A(n4998), .B(n4997), .Z(n4999) );
  AND U5717 ( .A(n5000), .B(n4999), .Z(n5004) );
  NOR U5718 ( .A(n5002), .B(n5001), .Z(n5003) );
  NANDN U5719 ( .A(n5004), .B(n5003), .Z(n5006) );
  ANDN U5720 ( .B(n5006), .A(n5005), .Z(n5008) );
  OR U5721 ( .A(n5008), .B(n5007), .Z(n5010) );
  ANDN U5722 ( .B(n5010), .A(n5009), .Z(n5011) );
  NAND U5723 ( .A(n5012), .B(n5011), .Z(n5013) );
  AND U5724 ( .A(n5014), .B(n5013), .Z(n5016) );
  NANDN U5725 ( .A(n5016), .B(n5015), .Z(n5017) );
  NANDN U5726 ( .A(n5018), .B(n5017), .Z(n5020) );
  NAND U5727 ( .A(n5020), .B(n5019), .Z(n5021) );
  NANDN U5728 ( .A(n5022), .B(n5021), .Z(n5024) );
  NAND U5729 ( .A(n5024), .B(n5023), .Z(n5026) );
  ANDN U5730 ( .B(n5026), .A(n5025), .Z(n5028) );
  NANDN U5731 ( .A(n5028), .B(n5027), .Z(n5029) );
  NANDN U5732 ( .A(n5030), .B(n5029), .Z(n5032) );
  NAND U5733 ( .A(n5032), .B(n5031), .Z(n5033) );
  NANDN U5734 ( .A(n5034), .B(n5033), .Z(n5036) );
  NAND U5735 ( .A(n5036), .B(n5035), .Z(n5038) );
  ANDN U5736 ( .B(n5038), .A(n5037), .Z(n5040) );
  NANDN U5737 ( .A(n5040), .B(n5039), .Z(n5041) );
  NANDN U5738 ( .A(n5042), .B(n5041), .Z(n5043) );
  NANDN U5739 ( .A(n5044), .B(n5043), .Z(n5045) );
  NANDN U5740 ( .A(n5046), .B(n5045), .Z(n5047) );
  NANDN U5741 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U5742 ( .A(n5050), .B(n5049), .Z(n5052) );
  NANDN U5743 ( .A(n5052), .B(n5051), .Z(n5054) );
  NAND U5744 ( .A(n5054), .B(n5053), .Z(n5055) );
  AND U5745 ( .A(n5056), .B(n5055), .Z(n5058) );
  NANDN U5746 ( .A(n5058), .B(n5057), .Z(n5060) );
  NAND U5747 ( .A(n5060), .B(n5059), .Z(n5062) );
  NAND U5748 ( .A(n5062), .B(n5061), .Z(n5064) );
  NAND U5749 ( .A(n5064), .B(n5063), .Z(n5066) );
  NAND U5750 ( .A(n5066), .B(n5065), .Z(n5067) );
  AND U5751 ( .A(n5068), .B(n5067), .Z(n5070) );
  NANDN U5752 ( .A(n5070), .B(n5069), .Z(n5072) );
  NAND U5753 ( .A(n5072), .B(n5071), .Z(n5074) );
  NAND U5754 ( .A(n5074), .B(n5073), .Z(n5076) );
  NAND U5755 ( .A(n5076), .B(n5075), .Z(n5078) );
  NAND U5756 ( .A(n5078), .B(n5077), .Z(n5079) );
  AND U5757 ( .A(n5080), .B(n5079), .Z(n5082) );
  NANDN U5758 ( .A(n5082), .B(n5081), .Z(n5084) );
  NAND U5759 ( .A(n5084), .B(n5083), .Z(n5086) );
  NAND U5760 ( .A(n5086), .B(n5085), .Z(n5087) );
  NANDN U5761 ( .A(n5088), .B(n5087), .Z(n5089) );
  NANDN U5762 ( .A(n5090), .B(n5089), .Z(n5091) );
  AND U5763 ( .A(n5092), .B(n5091), .Z(n5094) );
  NANDN U5764 ( .A(n5094), .B(n5093), .Z(n5096) );
  NAND U5765 ( .A(n5096), .B(n5095), .Z(n5098) );
  NAND U5766 ( .A(n5098), .B(n5097), .Z(n5100) );
  NAND U5767 ( .A(n5100), .B(n5099), .Z(n5102) );
  NAND U5768 ( .A(n5102), .B(n5101), .Z(n5103) );
  AND U5769 ( .A(n5104), .B(n5103), .Z(n5106) );
  NANDN U5770 ( .A(n5106), .B(n5105), .Z(n5108) );
  NAND U5771 ( .A(n5108), .B(n5107), .Z(n5110) );
  NAND U5772 ( .A(n5110), .B(n5109), .Z(n5112) );
  NAND U5773 ( .A(n5112), .B(n5111), .Z(n5114) );
  NAND U5774 ( .A(n5114), .B(n5113), .Z(n5115) );
  AND U5775 ( .A(n5116), .B(n5115), .Z(n5118) );
  NANDN U5776 ( .A(n5118), .B(n5117), .Z(n5120) );
  NAND U5777 ( .A(n5120), .B(n5119), .Z(n5122) );
  NAND U5778 ( .A(n5122), .B(n5121), .Z(n5124) );
  NAND U5779 ( .A(n5124), .B(n5123), .Z(n5126) );
  NAND U5780 ( .A(n5126), .B(n5125), .Z(n5127) );
  AND U5781 ( .A(n5128), .B(n5127), .Z(n5130) );
  NANDN U5782 ( .A(n5130), .B(n5129), .Z(n5132) );
  NAND U5783 ( .A(n5132), .B(n5131), .Z(n5134) );
  NAND U5784 ( .A(n5134), .B(n5133), .Z(n5136) );
  NAND U5785 ( .A(n5136), .B(n5135), .Z(n5138) );
  NAND U5786 ( .A(n5138), .B(n5137), .Z(n5139) );
  AND U5787 ( .A(n5140), .B(n5139), .Z(n5142) );
  NANDN U5788 ( .A(n5142), .B(n5141), .Z(n5144) );
  NAND U5789 ( .A(n5144), .B(n5143), .Z(n5146) );
  NAND U5790 ( .A(n5146), .B(n5145), .Z(n5148) );
  NAND U5791 ( .A(n5148), .B(n5147), .Z(n5150) );
  NAND U5792 ( .A(n5150), .B(n5149), .Z(n5151) );
  AND U5793 ( .A(n5152), .B(n5151), .Z(n5154) );
  NANDN U5794 ( .A(n5154), .B(n5153), .Z(n5156) );
  NAND U5795 ( .A(n5156), .B(n5155), .Z(n5158) );
  NAND U5796 ( .A(n5158), .B(n5157), .Z(n5160) );
  NAND U5797 ( .A(n5160), .B(n5159), .Z(n5162) );
  NAND U5798 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U5799 ( .A(n5164), .B(n5163), .Z(n5166) );
  NANDN U5800 ( .A(n5166), .B(n5165), .Z(n5168) );
  NAND U5801 ( .A(n5168), .B(n5167), .Z(n5170) );
  NAND U5802 ( .A(n5170), .B(n5169), .Z(n5171) );
  NANDN U5803 ( .A(n5172), .B(n5171), .Z(n5173) );
  NANDN U5804 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U5805 ( .A(n5176), .B(n5175), .Z(n5178) );
  NANDN U5806 ( .A(n5178), .B(n5177), .Z(n5179) );
  NANDN U5807 ( .A(n5180), .B(n5179), .Z(n5182) );
  NAND U5808 ( .A(n5182), .B(n5181), .Z(n5183) );
  NANDN U5809 ( .A(n5184), .B(n5183), .Z(n5186) );
  NAND U5810 ( .A(n5186), .B(n5185), .Z(n5188) );
  ANDN U5811 ( .B(n5188), .A(n5187), .Z(n5189) );
  OR U5812 ( .A(n5190), .B(n5189), .Z(n5191) );
  NANDN U5813 ( .A(n5192), .B(n5191), .Z(n5193) );
  NANDN U5814 ( .A(n5194), .B(n5193), .Z(n5195) );
  NANDN U5815 ( .A(n5196), .B(n5195), .Z(n5198) );
  NAND U5816 ( .A(n5198), .B(n5197), .Z(n5199) );
  NANDN U5817 ( .A(n5200), .B(n5199), .Z(n5202) );
  ANDN U5818 ( .B(n5202), .A(n5201), .Z(n5204) );
  NANDN U5819 ( .A(n5204), .B(n5203), .Z(n5206) );
  NAND U5820 ( .A(n5206), .B(n5205), .Z(n5207) );
  NANDN U5821 ( .A(n5208), .B(n5207), .Z(n5210) );
  NAND U5822 ( .A(n5210), .B(n5209), .Z(n5211) );
  NANDN U5823 ( .A(n5212), .B(n5211), .Z(n5213) );
  AND U5824 ( .A(n5214), .B(n5213), .Z(n5215) );
  OR U5825 ( .A(n5216), .B(n5215), .Z(n5218) );
  NAND U5826 ( .A(n5218), .B(n5217), .Z(n5219) );
  NANDN U5827 ( .A(n5220), .B(n5219), .Z(n5222) );
  NAND U5828 ( .A(n5222), .B(n5221), .Z(n5223) );
  NANDN U5829 ( .A(n5224), .B(n5223), .Z(n5225) );
  AND U5830 ( .A(n5226), .B(n5225), .Z(n5227) );
  OR U5831 ( .A(n5228), .B(n5227), .Z(n5230) );
  NAND U5832 ( .A(n5230), .B(n5229), .Z(n5231) );
  NANDN U5833 ( .A(n5232), .B(n5231), .Z(n5234) );
  NAND U5834 ( .A(n5234), .B(n5233), .Z(n5235) );
  NANDN U5835 ( .A(n5236), .B(n5235), .Z(n5237) );
  AND U5836 ( .A(n5238), .B(n5237), .Z(n5239) );
  OR U5837 ( .A(n5240), .B(n5239), .Z(n5242) );
  NAND U5838 ( .A(n5242), .B(n5241), .Z(n5243) );
  NANDN U5839 ( .A(n5244), .B(n5243), .Z(n5246) );
  NAND U5840 ( .A(n5246), .B(n5245), .Z(n5247) );
  NANDN U5841 ( .A(n5248), .B(n5247), .Z(n5249) );
  AND U5842 ( .A(n5250), .B(n5249), .Z(n5251) );
  OR U5843 ( .A(n5252), .B(n5251), .Z(n5254) );
  NAND U5844 ( .A(n5254), .B(n5253), .Z(n5255) );
  NANDN U5845 ( .A(n5256), .B(n5255), .Z(n5258) );
  NAND U5846 ( .A(n5258), .B(n5257), .Z(n5259) );
  NANDN U5847 ( .A(n5260), .B(n5259), .Z(n5261) );
  AND U5848 ( .A(n5262), .B(n5261), .Z(n5263) );
  OR U5849 ( .A(n5264), .B(n5263), .Z(n5266) );
  NAND U5850 ( .A(n5266), .B(n5265), .Z(n5267) );
  NANDN U5851 ( .A(n5268), .B(n5267), .Z(n5270) );
  NAND U5852 ( .A(n5270), .B(n5269), .Z(n5271) );
  NANDN U5853 ( .A(n5272), .B(n5271), .Z(n5273) );
  AND U5854 ( .A(n5274), .B(n5273), .Z(n5275) );
  OR U5855 ( .A(n5276), .B(n5275), .Z(n5278) );
  NAND U5856 ( .A(n5278), .B(n5277), .Z(n5279) );
  NANDN U5857 ( .A(n5280), .B(n5279), .Z(n5282) );
  NAND U5858 ( .A(n5282), .B(n5281), .Z(n5284) );
  NAND U5859 ( .A(n5284), .B(n5283), .Z(n5285) );
  AND U5860 ( .A(n5286), .B(n5285), .Z(n5288) );
  NANDN U5861 ( .A(n5288), .B(n5287), .Z(n5290) );
  NAND U5862 ( .A(n5290), .B(n5289), .Z(n5291) );
  NANDN U5863 ( .A(n5292), .B(n5291), .Z(n5294) );
  NAND U5864 ( .A(n5294), .B(n5293), .Z(n5295) );
  NANDN U5865 ( .A(n5296), .B(n5295), .Z(n5297) );
  AND U5866 ( .A(n5298), .B(n5297), .Z(n5299) );
  OR U5867 ( .A(n5300), .B(n5299), .Z(n5302) );
  NAND U5868 ( .A(n5302), .B(n5301), .Z(n5303) );
  NANDN U5869 ( .A(n5304), .B(n5303), .Z(n5306) );
  NAND U5870 ( .A(n5306), .B(n5305), .Z(n5307) );
  NANDN U5871 ( .A(n5308), .B(n5307), .Z(n5309) );
  AND U5872 ( .A(n5310), .B(n5309), .Z(n5311) );
  OR U5873 ( .A(n5312), .B(n5311), .Z(n5314) );
  NAND U5874 ( .A(n5314), .B(n5313), .Z(n5315) );
  NANDN U5875 ( .A(n5316), .B(n5315), .Z(n5318) );
  NAND U5876 ( .A(n5318), .B(n5317), .Z(n5319) );
  NANDN U5877 ( .A(n5320), .B(n5319), .Z(n5321) );
  AND U5878 ( .A(n5322), .B(n5321), .Z(n5323) );
  OR U5879 ( .A(n5324), .B(n5323), .Z(n5326) );
  NAND U5880 ( .A(n5326), .B(n5325), .Z(n5327) );
  NANDN U5881 ( .A(n5328), .B(n5327), .Z(n5330) );
  NAND U5882 ( .A(n5330), .B(n5329), .Z(n5331) );
  NANDN U5883 ( .A(n5332), .B(n5331), .Z(n5333) );
  AND U5884 ( .A(n5334), .B(n5333), .Z(n5335) );
  OR U5885 ( .A(n5336), .B(n5335), .Z(n5338) );
  NAND U5886 ( .A(n5338), .B(n5337), .Z(n5339) );
  NANDN U5887 ( .A(n5340), .B(n5339), .Z(n5342) );
  NAND U5888 ( .A(n5342), .B(n5341), .Z(n5343) );
  NANDN U5889 ( .A(n5344), .B(n5343), .Z(n5346) );
  ANDN U5890 ( .B(n5346), .A(n5345), .Z(n5348) );
  NANDN U5891 ( .A(n5348), .B(n5347), .Z(n5350) );
  NAND U5892 ( .A(n5350), .B(n5349), .Z(n5351) );
  NANDN U5893 ( .A(n5352), .B(n5351), .Z(n5354) );
  NAND U5894 ( .A(n5354), .B(n5353), .Z(n5355) );
  NANDN U5895 ( .A(n5356), .B(n5355), .Z(n5357) );
  AND U5896 ( .A(n5358), .B(n5357), .Z(n5359) );
  OR U5897 ( .A(n5360), .B(n5359), .Z(n5362) );
  NAND U5898 ( .A(n5362), .B(n5361), .Z(n5363) );
  NANDN U5899 ( .A(n5364), .B(n5363), .Z(n5366) );
  NAND U5900 ( .A(n5366), .B(n5365), .Z(n5367) );
  NANDN U5901 ( .A(n5368), .B(n5367), .Z(n5369) );
  AND U5902 ( .A(n5370), .B(n5369), .Z(n5371) );
  OR U5903 ( .A(n5372), .B(n5371), .Z(n5374) );
  NAND U5904 ( .A(n5374), .B(n5373), .Z(n5375) );
  NANDN U5905 ( .A(n5376), .B(n5375), .Z(n5378) );
  NAND U5906 ( .A(n5378), .B(n5377), .Z(n5379) );
  NANDN U5907 ( .A(n5380), .B(n5379), .Z(n5381) );
  AND U5908 ( .A(n5382), .B(n5381), .Z(n5383) );
  OR U5909 ( .A(n5384), .B(n5383), .Z(n5385) );
  AND U5910 ( .A(n5386), .B(n5385), .Z(n5387) );
  OR U5911 ( .A(n5388), .B(n5387), .Z(n5390) );
  NAND U5912 ( .A(n5390), .B(n5389), .Z(n5391) );
  NANDN U5913 ( .A(n5392), .B(n5391), .Z(n5394) );
  NAND U5914 ( .A(n5394), .B(n5393), .Z(n5395) );
  NANDN U5915 ( .A(n5396), .B(n5395), .Z(n5398) );
  ANDN U5916 ( .B(n5398), .A(n5397), .Z(n5400) );
  NANDN U5917 ( .A(n5400), .B(n5399), .Z(n5402) );
  NAND U5918 ( .A(n5402), .B(n5401), .Z(n5403) );
  NANDN U5919 ( .A(n5404), .B(n5403), .Z(n5406) );
  NAND U5920 ( .A(n5406), .B(n5405), .Z(n5407) );
  NANDN U5921 ( .A(n5408), .B(n5407), .Z(n5409) );
  AND U5922 ( .A(n5410), .B(n5409), .Z(n5411) );
  OR U5923 ( .A(n5412), .B(n5411), .Z(n5414) );
  NAND U5924 ( .A(n5414), .B(n5413), .Z(n5415) );
  NANDN U5925 ( .A(n5416), .B(n5415), .Z(n5418) );
  NAND U5926 ( .A(n5418), .B(n5417), .Z(n5420) );
  NAND U5927 ( .A(n5420), .B(n5419), .Z(n5421) );
  AND U5928 ( .A(n5422), .B(n5421), .Z(n5423) );
  OR U5929 ( .A(n5424), .B(n5423), .Z(n5426) );
  NAND U5930 ( .A(n5426), .B(n5425), .Z(n5427) );
  NANDN U5931 ( .A(n5428), .B(n5427), .Z(n5430) );
  NAND U5932 ( .A(n5430), .B(n5429), .Z(n5431) );
  NANDN U5933 ( .A(n5432), .B(n5431), .Z(n5433) );
  AND U5934 ( .A(n5434), .B(n5433), .Z(n5435) );
  OR U5935 ( .A(n5436), .B(n5435), .Z(n5438) );
  NAND U5936 ( .A(n5438), .B(n5437), .Z(n5439) );
  NANDN U5937 ( .A(n5440), .B(n5439), .Z(n5442) );
  NAND U5938 ( .A(n5442), .B(n5441), .Z(n5444) );
  NAND U5939 ( .A(n5444), .B(n5443), .Z(n5446) );
  ANDN U5940 ( .B(n5446), .A(n5445), .Z(n5447) );
  OR U5941 ( .A(n5448), .B(n5447), .Z(n5449) );
  AND U5942 ( .A(n5450), .B(n5449), .Z(n5451) );
  OR U5943 ( .A(n5452), .B(n5451), .Z(n5454) );
  NAND U5944 ( .A(n5454), .B(n5453), .Z(n5455) );
  NANDN U5945 ( .A(n5456), .B(n5455), .Z(n5458) );
  NAND U5946 ( .A(n5458), .B(n5457), .Z(n5459) );
  NANDN U5947 ( .A(n5460), .B(n5459), .Z(n5462) );
  ANDN U5948 ( .B(n5462), .A(n5461), .Z(n5464) );
  NANDN U5949 ( .A(n5464), .B(n5463), .Z(n5466) );
  NAND U5950 ( .A(n5466), .B(n5465), .Z(n5467) );
  NANDN U5951 ( .A(n5468), .B(n5467), .Z(n5470) );
  NAND U5952 ( .A(n5470), .B(n5469), .Z(n5471) );
  NANDN U5953 ( .A(n5472), .B(n5471), .Z(n5474) );
  NAND U5954 ( .A(n5474), .B(n5473), .Z(n5475) );
  NANDN U5955 ( .A(n5476), .B(n5475), .Z(n5478) );
  NAND U5956 ( .A(n5478), .B(n5477), .Z(n5480) );
  ANDN U5957 ( .B(n5480), .A(n5479), .Z(n5482) );
  NANDN U5958 ( .A(n5482), .B(n5481), .Z(n5483) );
  NANDN U5959 ( .A(n5484), .B(n5483), .Z(n5486) );
  NAND U5960 ( .A(n5486), .B(n5485), .Z(n5487) );
  NANDN U5961 ( .A(n5488), .B(n5487), .Z(n5490) );
  NAND U5962 ( .A(n5490), .B(n5489), .Z(n5491) );
  AND U5963 ( .A(n5492), .B(n5491), .Z(n5493) );
  OR U5964 ( .A(n5494), .B(n5493), .Z(n5495) );
  NANDN U5965 ( .A(n5496), .B(n5495), .Z(n5498) );
  NAND U5966 ( .A(n5498), .B(n5497), .Z(n5499) );
  NANDN U5967 ( .A(n5500), .B(n5499), .Z(n5502) );
  NAND U5968 ( .A(n5502), .B(n5501), .Z(n5504) );
  ANDN U5969 ( .B(n5504), .A(n5503), .Z(n5506) );
  NANDN U5970 ( .A(n5506), .B(n5505), .Z(n5508) );
  NAND U5971 ( .A(n5508), .B(n5507), .Z(n5510) );
  NAND U5972 ( .A(n5510), .B(n5509), .Z(n5511) );
  NANDN U5973 ( .A(n5512), .B(n5511), .Z(n5514) );
  NAND U5974 ( .A(n5514), .B(n5513), .Z(n5516) );
  ANDN U5975 ( .B(n5516), .A(n5515), .Z(n5517) );
  OR U5976 ( .A(n5518), .B(n5517), .Z(n5520) );
  NAND U5977 ( .A(n5520), .B(n5519), .Z(n5522) );
  NAND U5978 ( .A(n5522), .B(n5521), .Z(n5523) );
  NANDN U5979 ( .A(n5524), .B(n5523), .Z(n5526) );
  NAND U5980 ( .A(n5526), .B(n5525), .Z(n5528) );
  ANDN U5981 ( .B(n5528), .A(n5527), .Z(n5530) );
  NANDN U5982 ( .A(n5530), .B(n5529), .Z(n5532) );
  NAND U5983 ( .A(n5532), .B(n5531), .Z(n5534) );
  NAND U5984 ( .A(n5534), .B(n5533), .Z(n5535) );
  NANDN U5985 ( .A(n5536), .B(n5535), .Z(n5538) );
  NAND U5986 ( .A(n5538), .B(n5537), .Z(n5540) );
  ANDN U5987 ( .B(n5540), .A(n5539), .Z(n5541) );
  NAND U5988 ( .A(n5542), .B(n5541), .Z(n5543) );
  NAND U5989 ( .A(n5544), .B(n5543), .Z(n5546) );
  NAND U5990 ( .A(n5546), .B(n5545), .Z(n5548) );
  NAND U5991 ( .A(n5548), .B(n5547), .Z(n5549) );
  AND U5992 ( .A(n5550), .B(n5549), .Z(n5552) );
  NANDN U5993 ( .A(n5552), .B(n5551), .Z(n5554) );
  NAND U5994 ( .A(n5554), .B(n5553), .Z(n5556) );
  NAND U5995 ( .A(n5556), .B(n5555), .Z(n5558) );
  NAND U5996 ( .A(n5558), .B(n5557), .Z(n5560) );
  NAND U5997 ( .A(n5560), .B(n5559), .Z(n5561) );
  AND U5998 ( .A(n5562), .B(n5561), .Z(n5564) );
  NANDN U5999 ( .A(n5564), .B(n5563), .Z(n5566) );
  NAND U6000 ( .A(n5566), .B(n5565), .Z(n5568) );
  NAND U6001 ( .A(n5568), .B(n5567), .Z(n5570) );
  NAND U6002 ( .A(n5570), .B(n5569), .Z(n5572) );
  NAND U6003 ( .A(n5572), .B(n5571), .Z(n5573) );
  AND U6004 ( .A(n5574), .B(n5573), .Z(n5576) );
  NANDN U6005 ( .A(n5576), .B(n5575), .Z(n5578) );
  NAND U6006 ( .A(n5578), .B(n5577), .Z(n5580) );
  NAND U6007 ( .A(n5580), .B(n5579), .Z(n5582) );
  NAND U6008 ( .A(n5582), .B(n5581), .Z(n5584) );
  NAND U6009 ( .A(n5584), .B(n5583), .Z(n5585) );
  AND U6010 ( .A(n5586), .B(n5585), .Z(n5588) );
  NANDN U6011 ( .A(n5588), .B(n5587), .Z(n5590) );
  NAND U6012 ( .A(n5590), .B(n5589), .Z(n5592) );
  NAND U6013 ( .A(n5592), .B(n5591), .Z(n5594) );
  NAND U6014 ( .A(n5594), .B(n5593), .Z(n5596) );
  NAND U6015 ( .A(n5596), .B(n5595), .Z(n5597) );
  AND U6016 ( .A(n5598), .B(n5597), .Z(n5600) );
  NANDN U6017 ( .A(n5600), .B(n5599), .Z(n5602) );
  NAND U6018 ( .A(n5602), .B(n5601), .Z(n5604) );
  NAND U6019 ( .A(n5604), .B(n5603), .Z(n5606) );
  NAND U6020 ( .A(n5606), .B(n5605), .Z(n5608) );
  NAND U6021 ( .A(n5608), .B(n5607), .Z(n5609) );
  AND U6022 ( .A(n5610), .B(n5609), .Z(n5612) );
  NANDN U6023 ( .A(n5612), .B(n5611), .Z(n5614) );
  NAND U6024 ( .A(n5614), .B(n5613), .Z(n5616) );
  NAND U6025 ( .A(n5616), .B(n5615), .Z(n5618) );
  NAND U6026 ( .A(n5618), .B(n5617), .Z(n5620) );
  NAND U6027 ( .A(n5620), .B(n5619), .Z(n5621) );
  AND U6028 ( .A(n5622), .B(n5621), .Z(n5624) );
  NANDN U6029 ( .A(n5624), .B(n5623), .Z(n5626) );
  NAND U6030 ( .A(n5626), .B(n5625), .Z(n5628) );
  NAND U6031 ( .A(n5628), .B(n5627), .Z(n5630) );
  NAND U6032 ( .A(n5630), .B(n5629), .Z(n5632) );
  NAND U6033 ( .A(n5632), .B(n5631), .Z(n5633) );
  AND U6034 ( .A(n5634), .B(n5633), .Z(n5636) );
  NANDN U6035 ( .A(n5636), .B(n5635), .Z(n5638) );
  NAND U6036 ( .A(n5638), .B(n5637), .Z(n5639) );
  NANDN U6037 ( .A(n5640), .B(n5639), .Z(n5642) );
  NAND U6038 ( .A(n5642), .B(n5641), .Z(n5644) );
  NAND U6039 ( .A(n5644), .B(n5643), .Z(n5646) );
  NAND U6040 ( .A(n5646), .B(n5645), .Z(n5648) );
  NAND U6041 ( .A(n5648), .B(n5647), .Z(n5650) );
  NAND U6042 ( .A(n5650), .B(n5649), .Z(n5651) );
  AND U6043 ( .A(n5652), .B(n5651), .Z(n5654) );
  NANDN U6044 ( .A(n5654), .B(n5653), .Z(n5656) );
  NAND U6045 ( .A(n5656), .B(n5655), .Z(n5658) );
  NAND U6046 ( .A(n5658), .B(n5657), .Z(n5660) );
  NAND U6047 ( .A(n5660), .B(n5659), .Z(n5662) );
  NAND U6048 ( .A(n5662), .B(n5661), .Z(n5663) );
  AND U6049 ( .A(n5664), .B(n5663), .Z(n5666) );
  NANDN U6050 ( .A(n5666), .B(n5665), .Z(n5668) );
  NAND U6051 ( .A(n5668), .B(n5667), .Z(n5670) );
  NAND U6052 ( .A(n5670), .B(n5669), .Z(n5672) );
  NAND U6053 ( .A(n5672), .B(n5671), .Z(n5674) );
  NAND U6054 ( .A(n5674), .B(n5673), .Z(n5675) );
  AND U6055 ( .A(n5676), .B(n5675), .Z(n5678) );
  NANDN U6056 ( .A(n5678), .B(n5677), .Z(n5679) );
  NANDN U6057 ( .A(n5680), .B(n5679), .Z(n5682) );
  NAND U6058 ( .A(n5682), .B(n5681), .Z(n5684) );
  NAND U6059 ( .A(n5684), .B(n5683), .Z(n5686) );
  NAND U6060 ( .A(n5686), .B(n5685), .Z(n5687) );
  AND U6061 ( .A(n5688), .B(n5687), .Z(n5690) );
  NANDN U6062 ( .A(n5690), .B(n5689), .Z(n5692) );
  NAND U6063 ( .A(n5692), .B(n5691), .Z(n5694) );
  NAND U6064 ( .A(n5694), .B(n5693), .Z(n5696) );
  NAND U6065 ( .A(n5696), .B(n5695), .Z(n5698) );
  NAND U6066 ( .A(n5698), .B(n5697), .Z(n5699) );
  AND U6067 ( .A(n5700), .B(n5699), .Z(n5702) );
  NANDN U6068 ( .A(n5702), .B(n5701), .Z(n5703) );
  NANDN U6069 ( .A(n5704), .B(n5703), .Z(n5705) );
  NANDN U6070 ( .A(n5706), .B(n5705), .Z(n5708) );
  NAND U6071 ( .A(n5708), .B(n5707), .Z(n5709) );
  NANDN U6072 ( .A(n5710), .B(n5709), .Z(n5711) );
  AND U6073 ( .A(n5712), .B(n5711), .Z(n5713) );
  OR U6074 ( .A(n5714), .B(n5713), .Z(n5715) );
  AND U6075 ( .A(n5716), .B(n5715), .Z(n5717) );
  OR U6076 ( .A(n5718), .B(n5717), .Z(n5720) );
  NAND U6077 ( .A(n5720), .B(n5719), .Z(n5721) );
  NANDN U6078 ( .A(n5722), .B(n5721), .Z(n5723) );
  NAND U6079 ( .A(n5724), .B(n5723), .Z(n5725) );
  NANDN U6080 ( .A(n5726), .B(n5725), .Z(n5728) );
  ANDN U6081 ( .B(n5728), .A(n5727), .Z(n5730) );
  NANDN U6082 ( .A(n5730), .B(n5729), .Z(n5732) );
  NAND U6083 ( .A(n5732), .B(n5731), .Z(n5734) );
  ANDN U6084 ( .B(n5734), .A(n5733), .Z(n5736) );
  NANDN U6085 ( .A(n5736), .B(n5735), .Z(n5737) );
  NANDN U6086 ( .A(n5738), .B(n5737), .Z(n5739) );
  NANDN U6087 ( .A(n5740), .B(n5739), .Z(n5741) );
  NANDN U6088 ( .A(n5742), .B(n5741), .Z(n5744) );
  NAND U6089 ( .A(n5744), .B(n5743), .Z(n5745) );
  AND U6090 ( .A(n5746), .B(n5745), .Z(n5748) );
  NANDN U6091 ( .A(n5748), .B(n5747), .Z(n5749) );
  NANDN U6092 ( .A(n5750), .B(n5749), .Z(n5752) );
  NAND U6093 ( .A(n5752), .B(n5751), .Z(n5753) );
  NANDN U6094 ( .A(n5754), .B(n5753), .Z(n5756) );
  NAND U6095 ( .A(n5756), .B(n5755), .Z(n5758) );
  ANDN U6096 ( .B(n5758), .A(n5757), .Z(n5760) );
  NANDN U6097 ( .A(n5760), .B(n5759), .Z(n5761) );
  NANDN U6098 ( .A(n5762), .B(n5761), .Z(n5764) );
  NAND U6099 ( .A(n5764), .B(n5763), .Z(n5765) );
  NANDN U6100 ( .A(n5766), .B(n5765), .Z(n5768) );
  NAND U6101 ( .A(n5768), .B(n5767), .Z(n5770) );
  ANDN U6102 ( .B(n5770), .A(n5769), .Z(n5772) );
  NANDN U6103 ( .A(n5772), .B(n5771), .Z(n5773) );
  NANDN U6104 ( .A(n5774), .B(n5773), .Z(n5775) );
  NANDN U6105 ( .A(n5776), .B(n5775), .Z(n5777) );
  AND U6106 ( .A(n5778), .B(n5777), .Z(n5782) );
  NANDN U6107 ( .A(n5780), .B(n5779), .Z(n5781) );
  AND U6108 ( .A(n5782), .B(n5781), .Z(n5784) );
  NANDN U6109 ( .A(n5784), .B(n5783), .Z(n5785) );
  NANDN U6110 ( .A(n5786), .B(n5785), .Z(n5788) );
  NAND U6111 ( .A(n5788), .B(n5787), .Z(n5789) );
  NANDN U6112 ( .A(n5790), .B(n5789), .Z(n5792) );
  NAND U6113 ( .A(n5792), .B(n5791), .Z(n5794) );
  ANDN U6114 ( .B(n5794), .A(n5793), .Z(n5796) );
  ANDN U6115 ( .B(x[754]), .A(y[754]), .Z(n5795) );
  OR U6116 ( .A(n5796), .B(n5795), .Z(n5797) );
  NANDN U6117 ( .A(n5798), .B(n5797), .Z(n5799) );
  NANDN U6118 ( .A(n5800), .B(n5799), .Z(n5802) );
  NAND U6119 ( .A(n5802), .B(n5801), .Z(n5804) );
  NAND U6120 ( .A(n5804), .B(n5803), .Z(n5806) );
  ANDN U6121 ( .B(n5806), .A(n5805), .Z(n5807) );
  OR U6122 ( .A(n5808), .B(n5807), .Z(n5809) );
  NANDN U6123 ( .A(n5810), .B(n5809), .Z(n5811) );
  NANDN U6124 ( .A(n5812), .B(n5811), .Z(n5814) );
  NAND U6125 ( .A(n5814), .B(n5813), .Z(n5816) );
  NAND U6126 ( .A(n5816), .B(n5815), .Z(n5818) );
  ANDN U6127 ( .B(n5818), .A(n5817), .Z(n5820) );
  NANDN U6128 ( .A(n5820), .B(n5819), .Z(n5821) );
  NANDN U6129 ( .A(n5822), .B(n5821), .Z(n5824) );
  NAND U6130 ( .A(n5824), .B(n5823), .Z(n5825) );
  NANDN U6131 ( .A(n5826), .B(n5825), .Z(n5828) );
  NAND U6132 ( .A(n5828), .B(n5827), .Z(n5830) );
  ANDN U6133 ( .B(n5830), .A(n5829), .Z(n5832) );
  NANDN U6134 ( .A(n5832), .B(n5831), .Z(n5833) );
  NANDN U6135 ( .A(n5834), .B(n5833), .Z(n5836) );
  NAND U6136 ( .A(n5836), .B(n5835), .Z(n5838) );
  ANDN U6137 ( .B(x[772]), .A(y[772]), .Z(n5837) );
  OR U6138 ( .A(n5838), .B(n5837), .Z(n5840) );
  NAND U6139 ( .A(n5840), .B(n5839), .Z(n5841) );
  NANDN U6140 ( .A(n5842), .B(n5841), .Z(n5844) );
  NAND U6141 ( .A(n5844), .B(n5843), .Z(n5846) );
  NAND U6142 ( .A(n5846), .B(n5845), .Z(n5848) );
  ANDN U6143 ( .B(n5848), .A(n5847), .Z(n5850) );
  NANDN U6144 ( .A(n5850), .B(n5849), .Z(n5851) );
  NANDN U6145 ( .A(n5852), .B(n5851), .Z(n5854) );
  NAND U6146 ( .A(n5854), .B(n5853), .Z(n5855) );
  NANDN U6147 ( .A(n5856), .B(n5855), .Z(n5858) );
  ANDN U6148 ( .B(n5858), .A(n5857), .Z(n5860) );
  NAND U6149 ( .A(n5860), .B(n5859), .Z(n5862) );
  NAND U6150 ( .A(n5862), .B(n5861), .Z(n5864) );
  NAND U6151 ( .A(n5864), .B(n5863), .Z(n5866) );
  NAND U6152 ( .A(n5866), .B(n5865), .Z(n5868) );
  NAND U6153 ( .A(n5868), .B(n5867), .Z(n5869) );
  NANDN U6154 ( .A(n5870), .B(n5869), .Z(n5871) );
  AND U6155 ( .A(n5872), .B(n5871), .Z(n5873) );
  OR U6156 ( .A(n5874), .B(n5873), .Z(n5876) );
  NAND U6157 ( .A(n5876), .B(n5875), .Z(n5877) );
  NANDN U6158 ( .A(n5878), .B(n5877), .Z(n5880) );
  NAND U6159 ( .A(n5880), .B(n5879), .Z(n5881) );
  NANDN U6160 ( .A(n5882), .B(n5881), .Z(n5883) );
  AND U6161 ( .A(n5884), .B(n5883), .Z(n5885) );
  OR U6162 ( .A(n5886), .B(n5885), .Z(n5888) );
  NAND U6163 ( .A(n5888), .B(n5887), .Z(n5889) );
  NANDN U6164 ( .A(n5890), .B(n5889), .Z(n5892) );
  NAND U6165 ( .A(n5892), .B(n5891), .Z(n5893) );
  NANDN U6166 ( .A(n5894), .B(n5893), .Z(n5895) );
  AND U6167 ( .A(n5896), .B(n5895), .Z(n5897) );
  OR U6168 ( .A(n5898), .B(n5897), .Z(n5900) );
  NAND U6169 ( .A(n5900), .B(n5899), .Z(n5902) );
  NAND U6170 ( .A(n5902), .B(n5901), .Z(n5904) );
  NAND U6171 ( .A(n5904), .B(n5903), .Z(n5906) );
  NAND U6172 ( .A(n5906), .B(n5905), .Z(n5907) );
  AND U6173 ( .A(n5908), .B(n5907), .Z(n5909) );
  OR U6174 ( .A(n5910), .B(n5909), .Z(n5911) );
  NANDN U6175 ( .A(n5912), .B(n5911), .Z(n5914) );
  NAND U6176 ( .A(n5914), .B(n5913), .Z(n5918) );
  NAND U6177 ( .A(n5916), .B(n5915), .Z(n5917) );
  NANDN U6178 ( .A(n5918), .B(n5917), .Z(n5919) );
  NANDN U6179 ( .A(n5920), .B(n5919), .Z(n5922) );
  NAND U6180 ( .A(n5922), .B(n5921), .Z(n5924) );
  NAND U6181 ( .A(n5924), .B(n5923), .Z(n5925) );
  AND U6182 ( .A(n5926), .B(n5925), .Z(n5928) );
  NANDN U6183 ( .A(n5928), .B(n5927), .Z(n5930) );
  NAND U6184 ( .A(n5930), .B(n5929), .Z(n5932) );
  NAND U6185 ( .A(n5932), .B(n5931), .Z(n5934) );
  NAND U6186 ( .A(n5934), .B(n5933), .Z(n5936) );
  NAND U6187 ( .A(n5936), .B(n5935), .Z(n5937) );
  AND U6188 ( .A(n5938), .B(n5937), .Z(n5940) );
  NANDN U6189 ( .A(n5940), .B(n5939), .Z(n5942) );
  NAND U6190 ( .A(n5942), .B(n5941), .Z(n5944) );
  NAND U6191 ( .A(n5944), .B(n5943), .Z(n5946) );
  NAND U6192 ( .A(n5946), .B(n5945), .Z(n5948) );
  NAND U6193 ( .A(n5948), .B(n5947), .Z(n5949) );
  AND U6194 ( .A(n5950), .B(n5949), .Z(n5952) );
  NANDN U6195 ( .A(n5952), .B(n5951), .Z(n5954) );
  NAND U6196 ( .A(n5954), .B(n5953), .Z(n5956) );
  NAND U6197 ( .A(n5956), .B(n5955), .Z(n5958) );
  NAND U6198 ( .A(n5958), .B(n5957), .Z(n5960) );
  NAND U6199 ( .A(n5960), .B(n5959), .Z(n5961) );
  AND U6200 ( .A(n5962), .B(n5961), .Z(n5964) );
  NANDN U6201 ( .A(n5964), .B(n5963), .Z(n5966) );
  NAND U6202 ( .A(n5966), .B(n5965), .Z(n5968) );
  NAND U6203 ( .A(n5968), .B(n5967), .Z(n5970) );
  NAND U6204 ( .A(n5970), .B(n5969), .Z(n5972) );
  NAND U6205 ( .A(n5972), .B(n5971), .Z(n5973) );
  AND U6206 ( .A(n5974), .B(n5973), .Z(n5976) );
  NANDN U6207 ( .A(n5976), .B(n5975), .Z(n5978) );
  NAND U6208 ( .A(n5978), .B(n5977), .Z(n5980) );
  NAND U6209 ( .A(n5980), .B(n5979), .Z(n5982) );
  NAND U6210 ( .A(n5982), .B(n5981), .Z(n5984) );
  NAND U6211 ( .A(n5984), .B(n5983), .Z(n5985) );
  AND U6212 ( .A(n5986), .B(n5985), .Z(n5988) );
  NANDN U6213 ( .A(n5988), .B(n5987), .Z(n5990) );
  NAND U6214 ( .A(n5990), .B(n5989), .Z(n5992) );
  NAND U6215 ( .A(n5992), .B(n5991), .Z(n5994) );
  NAND U6216 ( .A(n5994), .B(n5993), .Z(n5996) );
  NAND U6217 ( .A(n5996), .B(n5995), .Z(n5997) );
  AND U6218 ( .A(n5998), .B(n5997), .Z(n6000) );
  NANDN U6219 ( .A(n6000), .B(n5999), .Z(n6002) );
  NAND U6220 ( .A(n6002), .B(n6001), .Z(n6003) );
  NANDN U6221 ( .A(n6004), .B(n6003), .Z(n6006) );
  NAND U6222 ( .A(n6006), .B(n6005), .Z(n6008) );
  NAND U6223 ( .A(n6008), .B(n6007), .Z(n6009) );
  AND U6224 ( .A(n6010), .B(n6009), .Z(n6012) );
  NANDN U6225 ( .A(n6012), .B(n6011), .Z(n6014) );
  NAND U6226 ( .A(n6014), .B(n6013), .Z(n6016) );
  NAND U6227 ( .A(n6016), .B(n6015), .Z(n6018) );
  NAND U6228 ( .A(n6018), .B(n6017), .Z(n6020) );
  NAND U6229 ( .A(n6020), .B(n6019), .Z(n6021) );
  AND U6230 ( .A(n6022), .B(n6021), .Z(n6024) );
  NAND U6231 ( .A(n6024), .B(n6023), .Z(n6025) );
  NANDN U6232 ( .A(n6026), .B(n6025), .Z(n6028) );
  ANDN U6233 ( .B(n6028), .A(n6027), .Z(n6030) );
  NANDN U6234 ( .A(n6030), .B(n6029), .Z(n6031) );
  AND U6235 ( .A(n6032), .B(n6031), .Z(n6033) );
  OR U6236 ( .A(n6034), .B(n6033), .Z(n6035) );
  NANDN U6237 ( .A(n6036), .B(n6035), .Z(n6038) );
  NAND U6238 ( .A(n6038), .B(n6037), .Z(n6040) );
  NAND U6239 ( .A(n6040), .B(n6039), .Z(n6041) );
  NANDN U6240 ( .A(n6042), .B(n6041), .Z(n6043) );
  AND U6241 ( .A(n6044), .B(n6043), .Z(n6045) );
  OR U6242 ( .A(n6046), .B(n6045), .Z(n6048) );
  NAND U6243 ( .A(n6048), .B(n6047), .Z(n6049) );
  NANDN U6244 ( .A(n6050), .B(n6049), .Z(n6052) );
  ANDN U6245 ( .B(n6052), .A(n6051), .Z(n6054) );
  NAND U6246 ( .A(n6054), .B(n6053), .Z(n6056) );
  NAND U6247 ( .A(n6056), .B(n6055), .Z(n6058) );
  AND U6248 ( .A(n6058), .B(n6057), .Z(n6060) );
  NAND U6249 ( .A(n6060), .B(n6059), .Z(n6062) );
  NAND U6250 ( .A(n6062), .B(n6061), .Z(n6063) );
  NANDN U6251 ( .A(n6064), .B(n6063), .Z(n6065) );
  NANDN U6252 ( .A(n6066), .B(n6065), .Z(n6067) );
  AND U6253 ( .A(n6068), .B(n6067), .Z(n6070) );
  NANDN U6254 ( .A(n6070), .B(n6069), .Z(n6072) );
  NAND U6255 ( .A(n6072), .B(n6071), .Z(n6074) );
  NAND U6256 ( .A(n6074), .B(n6073), .Z(n6076) );
  NAND U6257 ( .A(n6076), .B(n6075), .Z(n6078) );
  NAND U6258 ( .A(n6078), .B(n6077), .Z(n6079) );
  AND U6259 ( .A(n6080), .B(n6079), .Z(n6082) );
  NAND U6260 ( .A(n6082), .B(n6081), .Z(n6084) );
  NAND U6261 ( .A(n6084), .B(n6083), .Z(n6086) );
  ANDN U6262 ( .B(n6086), .A(n6085), .Z(n6088) );
  NANDN U6263 ( .A(n6088), .B(n6087), .Z(n6089) );
  NANDN U6264 ( .A(n6090), .B(n6089), .Z(n6091) );
  NANDN U6265 ( .A(n6092), .B(n6091), .Z(n6094) );
  NAND U6266 ( .A(n6094), .B(n6093), .Z(n6096) );
  NAND U6267 ( .A(n6096), .B(n6095), .Z(n6097) );
  AND U6268 ( .A(n6098), .B(n6097), .Z(n6100) );
  NANDN U6269 ( .A(n6100), .B(n6099), .Z(n6102) );
  NAND U6270 ( .A(n6102), .B(n6101), .Z(n6104) );
  NAND U6271 ( .A(n6104), .B(n6103), .Z(n6106) );
  NAND U6272 ( .A(n6106), .B(n6105), .Z(n6107) );
  NANDN U6273 ( .A(n6108), .B(n6107), .Z(n6110) );
  NAND U6274 ( .A(n6110), .B(n6109), .Z(n6112) );
  NAND U6275 ( .A(n6112), .B(n6111), .Z(n6114) );
  NAND U6276 ( .A(n6114), .B(n6113), .Z(n6116) );
  ANDN U6277 ( .B(n6116), .A(n6115), .Z(n6118) );
  NANDN U6278 ( .A(n6118), .B(n6117), .Z(n6119) );
  NANDN U6279 ( .A(n6120), .B(n6119), .Z(n6122) );
  NAND U6280 ( .A(n6122), .B(n6121), .Z(n6124) );
  NAND U6281 ( .A(n6124), .B(n6123), .Z(n6126) );
  NAND U6282 ( .A(n6126), .B(n6125), .Z(n6128) );
  ANDN U6283 ( .B(n6128), .A(n6127), .Z(n6130) );
  NANDN U6284 ( .A(n6130), .B(n6129), .Z(n6131) );
  NANDN U6285 ( .A(n6132), .B(n6131), .Z(n6134) );
  NAND U6286 ( .A(n6134), .B(n6133), .Z(n6135) );
  NANDN U6287 ( .A(n6136), .B(n6135), .Z(n6137) );
  AND U6288 ( .A(n6138), .B(n6137), .Z(n6139) );
  NANDN U6289 ( .A(n6140), .B(n6139), .Z(n6141) );
  NANDN U6290 ( .A(n6142), .B(n6141), .Z(n6146) );
  NAND U6291 ( .A(n6144), .B(n6143), .Z(n6145) );
  NAND U6292 ( .A(n6146), .B(n6145), .Z(n6148) );
  OR U6293 ( .A(n6148), .B(n6147), .Z(n6150) );
  NAND U6294 ( .A(n6150), .B(n6149), .Z(n6152) );
  NAND U6295 ( .A(n6152), .B(n6151), .Z(n6154) );
  NAND U6296 ( .A(n6154), .B(n6153), .Z(n6156) );
  NAND U6297 ( .A(n6156), .B(n6155), .Z(n6157) );
  AND U6298 ( .A(n6158), .B(n6157), .Z(n6160) );
  NANDN U6299 ( .A(n6160), .B(n6159), .Z(n6162) );
  NAND U6300 ( .A(n6162), .B(n6161), .Z(n6164) );
  NAND U6301 ( .A(n6164), .B(n6163), .Z(n6166) );
  NAND U6302 ( .A(n6166), .B(n6165), .Z(n6167) );
  AND U6303 ( .A(n6168), .B(n6167), .Z(n6169) );
  NANDN U6304 ( .A(n6170), .B(n6169), .Z(n6171) );
  AND U6305 ( .A(n6172), .B(n6171), .Z(n6173) );
  NAND U6306 ( .A(n6174), .B(n6173), .Z(n6175) );
  NAND U6307 ( .A(n6176), .B(n6175), .Z(n6178) );
  ANDN U6308 ( .B(n6178), .A(n6177), .Z(n6180) );
  NANDN U6309 ( .A(n6180), .B(n6179), .Z(n6181) );
  NANDN U6310 ( .A(n6182), .B(n6181), .Z(n6183) );
  NANDN U6311 ( .A(n6184), .B(n6183), .Z(n6186) );
  NAND U6312 ( .A(n6186), .B(n6185), .Z(n6188) );
  NAND U6313 ( .A(n6188), .B(n6187), .Z(n6190) );
  ANDN U6314 ( .B(n6190), .A(n6189), .Z(n6192) );
  NANDN U6315 ( .A(n6192), .B(n6191), .Z(n6193) );
  NANDN U6316 ( .A(n6194), .B(n6193), .Z(n6196) );
  NAND U6317 ( .A(n6196), .B(n6195), .Z(n6198) );
  NAND U6318 ( .A(n6198), .B(n6197), .Z(n6200) );
  ANDN U6319 ( .B(n6200), .A(n6199), .Z(n6202) );
  NAND U6320 ( .A(n6202), .B(n6201), .Z(n6206) );
  NANDN U6321 ( .A(n6204), .B(n6203), .Z(n6205) );
  AND U6322 ( .A(n6206), .B(n6205), .Z(n6208) );
  NANDN U6323 ( .A(n6208), .B(n6207), .Z(n6209) );
  NANDN U6324 ( .A(n6210), .B(n6209), .Z(n6212) );
  NAND U6325 ( .A(n6212), .B(n6211), .Z(n6214) );
  NAND U6326 ( .A(n6214), .B(n6213), .Z(n6216) );
  NAND U6327 ( .A(n6216), .B(n6215), .Z(n6217) );
  AND U6328 ( .A(n6218), .B(n6217), .Z(n6220) );
  NANDN U6329 ( .A(n6220), .B(n6219), .Z(n6222) );
  NAND U6330 ( .A(n6222), .B(n6221), .Z(n6223) );
  NANDN U6331 ( .A(n6224), .B(n6223), .Z(n6226) );
  NAND U6332 ( .A(n6226), .B(n6225), .Z(n6227) );
  NANDN U6333 ( .A(n6228), .B(n6227), .Z(n6229) );
  AND U6334 ( .A(n6230), .B(n6229), .Z(n6234) );
  ANDN U6335 ( .B(n6232), .A(n6231), .Z(n6233) );
  NANDN U6336 ( .A(n6234), .B(n6233), .Z(n6235) );
  AND U6337 ( .A(n6236), .B(n6235), .Z(n6237) );
  OR U6338 ( .A(n6238), .B(n6237), .Z(n6240) );
  NAND U6339 ( .A(n6240), .B(n6239), .Z(n6242) );
  NAND U6340 ( .A(n6242), .B(n6241), .Z(n6243) );
  NANDN U6341 ( .A(n6244), .B(n6243), .Z(n6245) );
  NANDN U6342 ( .A(n6246), .B(n6245), .Z(n6247) );
  AND U6343 ( .A(n6248), .B(n6247), .Z(n6250) );
  NANDN U6344 ( .A(n6250), .B(n6249), .Z(n6252) );
  NAND U6345 ( .A(n6252), .B(n6251), .Z(n6254) );
  NAND U6346 ( .A(n6254), .B(n6253), .Z(n6256) );
  NAND U6347 ( .A(n6256), .B(n6255), .Z(n6258) );
  NAND U6348 ( .A(n6258), .B(n6257), .Z(n6259) );
  AND U6349 ( .A(n6260), .B(n6259), .Z(n6262) );
  NANDN U6350 ( .A(n6262), .B(n6261), .Z(n6264) );
  NAND U6351 ( .A(n6264), .B(n6263), .Z(n6266) );
  NAND U6352 ( .A(n6266), .B(n6265), .Z(n6268) );
  NAND U6353 ( .A(n6268), .B(n6267), .Z(n6270) );
  NAND U6354 ( .A(n6270), .B(n6269), .Z(n6271) );
  AND U6355 ( .A(n6272), .B(n6271), .Z(n6274) );
  NANDN U6356 ( .A(n6274), .B(n6273), .Z(n6276) );
  NAND U6357 ( .A(n6276), .B(n6275), .Z(n6278) );
  NAND U6358 ( .A(n6278), .B(n6277), .Z(n6280) );
  NAND U6359 ( .A(n6280), .B(n6279), .Z(n6282) );
  NAND U6360 ( .A(n6282), .B(n6281), .Z(n6283) );
  AND U6361 ( .A(n6284), .B(n6283), .Z(n6286) );
  NANDN U6362 ( .A(n6286), .B(n6285), .Z(n6288) );
  NAND U6363 ( .A(n6288), .B(n6287), .Z(n6290) );
  NAND U6364 ( .A(n6290), .B(n6289), .Z(n6292) );
  NAND U6365 ( .A(n6292), .B(n6291), .Z(n6294) );
  NAND U6366 ( .A(n6294), .B(n6293), .Z(n6295) );
  AND U6367 ( .A(n6296), .B(n6295), .Z(n6298) );
  NANDN U6368 ( .A(n6298), .B(n6297), .Z(n6300) );
  NAND U6369 ( .A(n6300), .B(n6299), .Z(n6302) );
  NAND U6370 ( .A(n6302), .B(n6301), .Z(n6304) );
  NAND U6371 ( .A(n6304), .B(n6303), .Z(n6306) );
  NAND U6372 ( .A(n6306), .B(n6305), .Z(n6307) );
  AND U6373 ( .A(n6308), .B(n6307), .Z(n6310) );
  NANDN U6374 ( .A(n6310), .B(n6309), .Z(n6312) );
  NAND U6375 ( .A(n6312), .B(n6311), .Z(n6314) );
  NAND U6376 ( .A(n6314), .B(n6313), .Z(n6316) );
  NAND U6377 ( .A(n6316), .B(n6315), .Z(n6317) );
  AND U6378 ( .A(n6318), .B(n6317), .Z(n6319) );
  NANDN U6379 ( .A(n6320), .B(n6319), .Z(n6322) );
  NAND U6380 ( .A(n6322), .B(n6321), .Z(n6323) );
  NANDN U6381 ( .A(n6324), .B(n6323), .Z(n6325) );
  AND U6382 ( .A(n6326), .B(n6325), .Z(n6327) );
  OR U6383 ( .A(n6328), .B(n6327), .Z(n6329) );
  NANDN U6384 ( .A(n6330), .B(n6329), .Z(n6332) );
  NAND U6385 ( .A(n6332), .B(n6331), .Z(n6333) );
  NAND U6386 ( .A(n6334), .B(n6333), .Z(n6336) );
  NAND U6387 ( .A(n6336), .B(n6335), .Z(n6337) );
  AND U6388 ( .A(n6338), .B(n6337), .Z(n6339) );
  OR U6389 ( .A(n6340), .B(n6339), .Z(n6342) );
  NAND U6390 ( .A(n6342), .B(n6341), .Z(n6343) );
  NANDN U6391 ( .A(n6344), .B(n6343), .Z(n6346) );
  NAND U6392 ( .A(n6346), .B(n6345), .Z(n6347) );
  AND U6393 ( .A(n6348), .B(n6347), .Z(n6349) );
  OR U6394 ( .A(n6350), .B(n6349), .Z(n6352) );
  NAND U6395 ( .A(n6352), .B(n6351), .Z(n6354) );
  NAND U6396 ( .A(n6354), .B(n6353), .Z(n6356) );
  OR U6397 ( .A(n6356), .B(n6355), .Z(n6357) );
  NANDN U6398 ( .A(n6358), .B(n6357), .Z(n6360) );
  NAND U6399 ( .A(n6360), .B(n6359), .Z(n6362) );
  NAND U6400 ( .A(n6362), .B(n6361), .Z(n6363) );
  NANDN U6401 ( .A(n6364), .B(n6363), .Z(n6365) );
  AND U6402 ( .A(n6366), .B(n6365), .Z(n6367) );
  OR U6403 ( .A(n6368), .B(n6367), .Z(n6370) );
  NAND U6404 ( .A(n6370), .B(n6369), .Z(n6371) );
  NANDN U6405 ( .A(n6372), .B(n6371), .Z(n6374) );
  ANDN U6406 ( .B(n6374), .A(n6373), .Z(n6376) );
  NAND U6407 ( .A(n6376), .B(n6375), .Z(n6377) );
  NANDN U6408 ( .A(n6378), .B(n6377), .Z(n6380) );
  ANDN U6409 ( .B(n6380), .A(n6379), .Z(n6382) );
  NAND U6410 ( .A(n6382), .B(n6381), .Z(n6383) );
  NANDN U6411 ( .A(n6384), .B(n6383), .Z(n6385) );
  AND U6412 ( .A(n6386), .B(n6385), .Z(n6388) );
  OR U6413 ( .A(n6388), .B(n6387), .Z(n6390) );
  NAND U6414 ( .A(n6390), .B(n6389), .Z(n6391) );
  NANDN U6415 ( .A(n6392), .B(n6391), .Z(n6394) );
  NAND U6416 ( .A(n6394), .B(n6393), .Z(n6396) );
  NAND U6417 ( .A(n6396), .B(n6395), .Z(n6397) );
  AND U6418 ( .A(n6398), .B(n6397), .Z(n6400) );
  NANDN U6419 ( .A(n6400), .B(n6399), .Z(n6401) );
  NANDN U6420 ( .A(n6402), .B(n6401), .Z(n6403) );
  NANDN U6421 ( .A(n6404), .B(n6403), .Z(n6406) );
  NAND U6422 ( .A(n6406), .B(n6405), .Z(n6407) );
  NANDN U6423 ( .A(n6408), .B(n6407), .Z(n6410) );
  ANDN U6424 ( .B(n6410), .A(n6409), .Z(n6411) );
  OR U6425 ( .A(n6412), .B(n6411), .Z(n6413) );
  NANDN U6426 ( .A(n6414), .B(n6413), .Z(n6415) );
  NANDN U6427 ( .A(n6416), .B(n6415), .Z(n6417) );
  NANDN U6428 ( .A(n6418), .B(n6417), .Z(n6419) );
  NANDN U6429 ( .A(n6420), .B(n6419), .Z(n6422) );
  ANDN U6430 ( .B(n6422), .A(n6421), .Z(n6423) );
  OR U6431 ( .A(n6424), .B(n6423), .Z(n6425) );
  AND U6432 ( .A(n6426), .B(n6425), .Z(n6427) );
  NANDN U6433 ( .A(n6428), .B(n6427), .Z(n6430) );
  NAND U6434 ( .A(n6428), .B(g), .Z(n6429) );
  NAND U6435 ( .A(n6430), .B(n6429), .Z(n4) );
endmodule

