
module mult_N256_CC256 ( clk, rst, a, b, c );
  input [255:0] a;
  input [0:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530;
  wire   [511:0] sreg;

  DFF \sreg_reg[510]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[510]) );
  DFF \sreg_reg[509]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[509]) );
  DFF \sreg_reg[508]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[508]) );
  DFF \sreg_reg[507]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U4 ( .A(sreg[258]), .B(n771), .Z(n1) );
  NANDN U5 ( .A(n772), .B(n1), .Z(n2) );
  NAND U6 ( .A(sreg[258]), .B(n771), .Z(n3) );
  AND U7 ( .A(n2), .B(n3), .Z(n775) );
  XOR U8 ( .A(sreg[261]), .B(n780), .Z(n4) );
  NANDN U9 ( .A(n781), .B(n4), .Z(n5) );
  NAND U10 ( .A(sreg[261]), .B(n780), .Z(n6) );
  AND U11 ( .A(n5), .B(n6), .Z(n784) );
  XOR U12 ( .A(sreg[264]), .B(n789), .Z(n7) );
  NANDN U13 ( .A(n790), .B(n7), .Z(n8) );
  NAND U14 ( .A(sreg[264]), .B(n789), .Z(n9) );
  AND U15 ( .A(n8), .B(n9), .Z(n793) );
  XOR U16 ( .A(sreg[267]), .B(n798), .Z(n10) );
  NANDN U17 ( .A(n799), .B(n10), .Z(n11) );
  NAND U18 ( .A(sreg[267]), .B(n798), .Z(n12) );
  AND U19 ( .A(n11), .B(n12), .Z(n802) );
  XOR U20 ( .A(sreg[270]), .B(n807), .Z(n13) );
  NANDN U21 ( .A(n808), .B(n13), .Z(n14) );
  NAND U22 ( .A(sreg[270]), .B(n807), .Z(n15) );
  AND U23 ( .A(n14), .B(n15), .Z(n811) );
  XOR U24 ( .A(sreg[273]), .B(n816), .Z(n16) );
  NANDN U25 ( .A(n817), .B(n16), .Z(n17) );
  NAND U26 ( .A(sreg[273]), .B(n816), .Z(n18) );
  AND U27 ( .A(n17), .B(n18), .Z(n820) );
  XOR U28 ( .A(sreg[276]), .B(n825), .Z(n19) );
  NANDN U29 ( .A(n826), .B(n19), .Z(n20) );
  NAND U30 ( .A(sreg[276]), .B(n825), .Z(n21) );
  AND U31 ( .A(n20), .B(n21), .Z(n829) );
  XOR U32 ( .A(sreg[279]), .B(n834), .Z(n22) );
  NANDN U33 ( .A(n835), .B(n22), .Z(n23) );
  NAND U34 ( .A(sreg[279]), .B(n834), .Z(n24) );
  AND U35 ( .A(n23), .B(n24), .Z(n838) );
  XOR U36 ( .A(sreg[282]), .B(n843), .Z(n25) );
  NANDN U37 ( .A(n844), .B(n25), .Z(n26) );
  NAND U38 ( .A(sreg[282]), .B(n843), .Z(n27) );
  AND U39 ( .A(n26), .B(n27), .Z(n847) );
  XOR U40 ( .A(sreg[285]), .B(n852), .Z(n28) );
  NANDN U41 ( .A(n853), .B(n28), .Z(n29) );
  NAND U42 ( .A(sreg[285]), .B(n852), .Z(n30) );
  AND U43 ( .A(n29), .B(n30), .Z(n856) );
  XOR U44 ( .A(sreg[288]), .B(n861), .Z(n31) );
  NANDN U45 ( .A(n862), .B(n31), .Z(n32) );
  NAND U46 ( .A(sreg[288]), .B(n861), .Z(n33) );
  AND U47 ( .A(n32), .B(n33), .Z(n865) );
  XOR U48 ( .A(sreg[291]), .B(n870), .Z(n34) );
  NANDN U49 ( .A(n871), .B(n34), .Z(n35) );
  NAND U50 ( .A(sreg[291]), .B(n870), .Z(n36) );
  AND U51 ( .A(n35), .B(n36), .Z(n874) );
  XOR U52 ( .A(sreg[294]), .B(n879), .Z(n37) );
  NANDN U53 ( .A(n880), .B(n37), .Z(n38) );
  NAND U54 ( .A(sreg[294]), .B(n879), .Z(n39) );
  AND U55 ( .A(n38), .B(n39), .Z(n883) );
  XOR U56 ( .A(sreg[297]), .B(n888), .Z(n40) );
  NANDN U57 ( .A(n889), .B(n40), .Z(n41) );
  NAND U58 ( .A(sreg[297]), .B(n888), .Z(n42) );
  AND U59 ( .A(n41), .B(n42), .Z(n892) );
  XOR U60 ( .A(sreg[300]), .B(n897), .Z(n43) );
  NANDN U61 ( .A(n898), .B(n43), .Z(n44) );
  NAND U62 ( .A(sreg[300]), .B(n897), .Z(n45) );
  AND U63 ( .A(n44), .B(n45), .Z(n901) );
  XOR U64 ( .A(sreg[303]), .B(n906), .Z(n46) );
  NANDN U65 ( .A(n907), .B(n46), .Z(n47) );
  NAND U66 ( .A(sreg[303]), .B(n906), .Z(n48) );
  AND U67 ( .A(n47), .B(n48), .Z(n910) );
  XOR U68 ( .A(sreg[306]), .B(n915), .Z(n49) );
  NANDN U69 ( .A(n916), .B(n49), .Z(n50) );
  NAND U70 ( .A(sreg[306]), .B(n915), .Z(n51) );
  AND U71 ( .A(n50), .B(n51), .Z(n919) );
  XOR U72 ( .A(sreg[309]), .B(n924), .Z(n52) );
  NANDN U73 ( .A(n925), .B(n52), .Z(n53) );
  NAND U74 ( .A(sreg[309]), .B(n924), .Z(n54) );
  AND U75 ( .A(n53), .B(n54), .Z(n928) );
  XOR U76 ( .A(sreg[312]), .B(n933), .Z(n55) );
  NANDN U77 ( .A(n934), .B(n55), .Z(n56) );
  NAND U78 ( .A(sreg[312]), .B(n933), .Z(n57) );
  AND U79 ( .A(n56), .B(n57), .Z(n937) );
  XOR U80 ( .A(sreg[315]), .B(n942), .Z(n58) );
  NANDN U81 ( .A(n943), .B(n58), .Z(n59) );
  NAND U82 ( .A(sreg[315]), .B(n942), .Z(n60) );
  AND U83 ( .A(n59), .B(n60), .Z(n946) );
  XOR U84 ( .A(sreg[318]), .B(n951), .Z(n61) );
  NANDN U85 ( .A(n952), .B(n61), .Z(n62) );
  NAND U86 ( .A(sreg[318]), .B(n951), .Z(n63) );
  AND U87 ( .A(n62), .B(n63), .Z(n955) );
  XOR U88 ( .A(sreg[321]), .B(n960), .Z(n64) );
  NANDN U89 ( .A(n961), .B(n64), .Z(n65) );
  NAND U90 ( .A(sreg[321]), .B(n960), .Z(n66) );
  AND U91 ( .A(n65), .B(n66), .Z(n964) );
  XOR U92 ( .A(sreg[324]), .B(n969), .Z(n67) );
  NANDN U93 ( .A(n970), .B(n67), .Z(n68) );
  NAND U94 ( .A(sreg[324]), .B(n969), .Z(n69) );
  AND U95 ( .A(n68), .B(n69), .Z(n973) );
  XOR U96 ( .A(sreg[327]), .B(n978), .Z(n70) );
  NANDN U97 ( .A(n979), .B(n70), .Z(n71) );
  NAND U98 ( .A(sreg[327]), .B(n978), .Z(n72) );
  AND U99 ( .A(n71), .B(n72), .Z(n982) );
  XOR U100 ( .A(sreg[330]), .B(n987), .Z(n73) );
  NANDN U101 ( .A(n988), .B(n73), .Z(n74) );
  NAND U102 ( .A(sreg[330]), .B(n987), .Z(n75) );
  AND U103 ( .A(n74), .B(n75), .Z(n991) );
  XOR U104 ( .A(sreg[333]), .B(n996), .Z(n76) );
  NANDN U105 ( .A(n997), .B(n76), .Z(n77) );
  NAND U106 ( .A(sreg[333]), .B(n996), .Z(n78) );
  AND U107 ( .A(n77), .B(n78), .Z(n1000) );
  XOR U108 ( .A(sreg[336]), .B(n1005), .Z(n79) );
  NANDN U109 ( .A(n1006), .B(n79), .Z(n80) );
  NAND U110 ( .A(sreg[336]), .B(n1005), .Z(n81) );
  AND U111 ( .A(n80), .B(n81), .Z(n1009) );
  XOR U112 ( .A(sreg[339]), .B(n1014), .Z(n82) );
  NANDN U113 ( .A(n1015), .B(n82), .Z(n83) );
  NAND U114 ( .A(sreg[339]), .B(n1014), .Z(n84) );
  AND U115 ( .A(n83), .B(n84), .Z(n1018) );
  XOR U116 ( .A(sreg[342]), .B(n1023), .Z(n85) );
  NANDN U117 ( .A(n1024), .B(n85), .Z(n86) );
  NAND U118 ( .A(sreg[342]), .B(n1023), .Z(n87) );
  AND U119 ( .A(n86), .B(n87), .Z(n1027) );
  XOR U120 ( .A(sreg[345]), .B(n1032), .Z(n88) );
  NANDN U121 ( .A(n1033), .B(n88), .Z(n89) );
  NAND U122 ( .A(sreg[345]), .B(n1032), .Z(n90) );
  AND U123 ( .A(n89), .B(n90), .Z(n1036) );
  XOR U124 ( .A(sreg[348]), .B(n1041), .Z(n91) );
  NANDN U125 ( .A(n1042), .B(n91), .Z(n92) );
  NAND U126 ( .A(sreg[348]), .B(n1041), .Z(n93) );
  AND U127 ( .A(n92), .B(n93), .Z(n1045) );
  XOR U128 ( .A(sreg[351]), .B(n1050), .Z(n94) );
  NANDN U129 ( .A(n1051), .B(n94), .Z(n95) );
  NAND U130 ( .A(sreg[351]), .B(n1050), .Z(n96) );
  AND U131 ( .A(n95), .B(n96), .Z(n1054) );
  XOR U132 ( .A(sreg[354]), .B(n1059), .Z(n97) );
  NANDN U133 ( .A(n1060), .B(n97), .Z(n98) );
  NAND U134 ( .A(sreg[354]), .B(n1059), .Z(n99) );
  AND U135 ( .A(n98), .B(n99), .Z(n1063) );
  XOR U136 ( .A(sreg[357]), .B(n1068), .Z(n100) );
  NANDN U137 ( .A(n1069), .B(n100), .Z(n101) );
  NAND U138 ( .A(sreg[357]), .B(n1068), .Z(n102) );
  AND U139 ( .A(n101), .B(n102), .Z(n1072) );
  XOR U140 ( .A(sreg[360]), .B(n1077), .Z(n103) );
  NANDN U141 ( .A(n1078), .B(n103), .Z(n104) );
  NAND U142 ( .A(sreg[360]), .B(n1077), .Z(n105) );
  AND U143 ( .A(n104), .B(n105), .Z(n1081) );
  XOR U144 ( .A(sreg[363]), .B(n1086), .Z(n106) );
  NANDN U145 ( .A(n1087), .B(n106), .Z(n107) );
  NAND U146 ( .A(sreg[363]), .B(n1086), .Z(n108) );
  AND U147 ( .A(n107), .B(n108), .Z(n1090) );
  XOR U148 ( .A(sreg[366]), .B(n1095), .Z(n109) );
  NANDN U149 ( .A(n1096), .B(n109), .Z(n110) );
  NAND U150 ( .A(sreg[366]), .B(n1095), .Z(n111) );
  AND U151 ( .A(n110), .B(n111), .Z(n1099) );
  XOR U152 ( .A(sreg[369]), .B(n1104), .Z(n112) );
  NANDN U153 ( .A(n1105), .B(n112), .Z(n113) );
  NAND U154 ( .A(sreg[369]), .B(n1104), .Z(n114) );
  AND U155 ( .A(n113), .B(n114), .Z(n1108) );
  XOR U156 ( .A(sreg[372]), .B(n1113), .Z(n115) );
  NANDN U157 ( .A(n1114), .B(n115), .Z(n116) );
  NAND U158 ( .A(sreg[372]), .B(n1113), .Z(n117) );
  AND U159 ( .A(n116), .B(n117), .Z(n1117) );
  XOR U160 ( .A(sreg[375]), .B(n1122), .Z(n118) );
  NANDN U161 ( .A(n1123), .B(n118), .Z(n119) );
  NAND U162 ( .A(sreg[375]), .B(n1122), .Z(n120) );
  AND U163 ( .A(n119), .B(n120), .Z(n1126) );
  XOR U164 ( .A(sreg[378]), .B(n1131), .Z(n121) );
  NANDN U165 ( .A(n1132), .B(n121), .Z(n122) );
  NAND U166 ( .A(sreg[378]), .B(n1131), .Z(n123) );
  AND U167 ( .A(n122), .B(n123), .Z(n1135) );
  XOR U168 ( .A(sreg[381]), .B(n1140), .Z(n124) );
  NANDN U169 ( .A(n1141), .B(n124), .Z(n125) );
  NAND U170 ( .A(sreg[381]), .B(n1140), .Z(n126) );
  AND U171 ( .A(n125), .B(n126), .Z(n1144) );
  XOR U172 ( .A(sreg[384]), .B(n1149), .Z(n127) );
  NANDN U173 ( .A(n1150), .B(n127), .Z(n128) );
  NAND U174 ( .A(sreg[384]), .B(n1149), .Z(n129) );
  AND U175 ( .A(n128), .B(n129), .Z(n1153) );
  XOR U176 ( .A(sreg[387]), .B(n1158), .Z(n130) );
  NANDN U177 ( .A(n1159), .B(n130), .Z(n131) );
  NAND U178 ( .A(sreg[387]), .B(n1158), .Z(n132) );
  AND U179 ( .A(n131), .B(n132), .Z(n1162) );
  XOR U180 ( .A(sreg[390]), .B(n1167), .Z(n133) );
  NANDN U181 ( .A(n1168), .B(n133), .Z(n134) );
  NAND U182 ( .A(sreg[390]), .B(n1167), .Z(n135) );
  AND U183 ( .A(n134), .B(n135), .Z(n1171) );
  XOR U184 ( .A(sreg[393]), .B(n1176), .Z(n136) );
  NANDN U185 ( .A(n1177), .B(n136), .Z(n137) );
  NAND U186 ( .A(sreg[393]), .B(n1176), .Z(n138) );
  AND U187 ( .A(n137), .B(n138), .Z(n1180) );
  XOR U188 ( .A(sreg[396]), .B(n1185), .Z(n139) );
  NANDN U189 ( .A(n1186), .B(n139), .Z(n140) );
  NAND U190 ( .A(sreg[396]), .B(n1185), .Z(n141) );
  AND U191 ( .A(n140), .B(n141), .Z(n1189) );
  XOR U192 ( .A(sreg[399]), .B(n1194), .Z(n142) );
  NANDN U193 ( .A(n1195), .B(n142), .Z(n143) );
  NAND U194 ( .A(sreg[399]), .B(n1194), .Z(n144) );
  AND U195 ( .A(n143), .B(n144), .Z(n1198) );
  XOR U196 ( .A(sreg[402]), .B(n1203), .Z(n145) );
  NANDN U197 ( .A(n1204), .B(n145), .Z(n146) );
  NAND U198 ( .A(sreg[402]), .B(n1203), .Z(n147) );
  AND U199 ( .A(n146), .B(n147), .Z(n1207) );
  XOR U200 ( .A(sreg[405]), .B(n1212), .Z(n148) );
  NANDN U201 ( .A(n1213), .B(n148), .Z(n149) );
  NAND U202 ( .A(sreg[405]), .B(n1212), .Z(n150) );
  AND U203 ( .A(n149), .B(n150), .Z(n1216) );
  XOR U204 ( .A(sreg[408]), .B(n1221), .Z(n151) );
  NANDN U205 ( .A(n1222), .B(n151), .Z(n152) );
  NAND U206 ( .A(sreg[408]), .B(n1221), .Z(n153) );
  AND U207 ( .A(n152), .B(n153), .Z(n1225) );
  XOR U208 ( .A(sreg[411]), .B(n1230), .Z(n154) );
  NANDN U209 ( .A(n1231), .B(n154), .Z(n155) );
  NAND U210 ( .A(sreg[411]), .B(n1230), .Z(n156) );
  AND U211 ( .A(n155), .B(n156), .Z(n1234) );
  XOR U212 ( .A(sreg[414]), .B(n1239), .Z(n157) );
  NANDN U213 ( .A(n1240), .B(n157), .Z(n158) );
  NAND U214 ( .A(sreg[414]), .B(n1239), .Z(n159) );
  AND U215 ( .A(n158), .B(n159), .Z(n1243) );
  XOR U216 ( .A(sreg[417]), .B(n1248), .Z(n160) );
  NANDN U217 ( .A(n1249), .B(n160), .Z(n161) );
  NAND U218 ( .A(sreg[417]), .B(n1248), .Z(n162) );
  AND U219 ( .A(n161), .B(n162), .Z(n1252) );
  XOR U220 ( .A(sreg[420]), .B(n1257), .Z(n163) );
  NANDN U221 ( .A(n1258), .B(n163), .Z(n164) );
  NAND U222 ( .A(sreg[420]), .B(n1257), .Z(n165) );
  AND U223 ( .A(n164), .B(n165), .Z(n1261) );
  XOR U224 ( .A(sreg[423]), .B(n1266), .Z(n166) );
  NANDN U225 ( .A(n1267), .B(n166), .Z(n167) );
  NAND U226 ( .A(sreg[423]), .B(n1266), .Z(n168) );
  AND U227 ( .A(n167), .B(n168), .Z(n1270) );
  XOR U228 ( .A(sreg[426]), .B(n1275), .Z(n169) );
  NANDN U229 ( .A(n1276), .B(n169), .Z(n170) );
  NAND U230 ( .A(sreg[426]), .B(n1275), .Z(n171) );
  AND U231 ( .A(n170), .B(n171), .Z(n1279) );
  XOR U232 ( .A(sreg[429]), .B(n1284), .Z(n172) );
  NANDN U233 ( .A(n1285), .B(n172), .Z(n173) );
  NAND U234 ( .A(sreg[429]), .B(n1284), .Z(n174) );
  AND U235 ( .A(n173), .B(n174), .Z(n1288) );
  XOR U236 ( .A(sreg[432]), .B(n1293), .Z(n175) );
  NANDN U237 ( .A(n1294), .B(n175), .Z(n176) );
  NAND U238 ( .A(sreg[432]), .B(n1293), .Z(n177) );
  AND U239 ( .A(n176), .B(n177), .Z(n1297) );
  XOR U240 ( .A(sreg[435]), .B(n1302), .Z(n178) );
  NANDN U241 ( .A(n1303), .B(n178), .Z(n179) );
  NAND U242 ( .A(sreg[435]), .B(n1302), .Z(n180) );
  AND U243 ( .A(n179), .B(n180), .Z(n1306) );
  XOR U244 ( .A(sreg[438]), .B(n1311), .Z(n181) );
  NANDN U245 ( .A(n1312), .B(n181), .Z(n182) );
  NAND U246 ( .A(sreg[438]), .B(n1311), .Z(n183) );
  AND U247 ( .A(n182), .B(n183), .Z(n1315) );
  XOR U248 ( .A(sreg[441]), .B(n1320), .Z(n184) );
  NANDN U249 ( .A(n1321), .B(n184), .Z(n185) );
  NAND U250 ( .A(sreg[441]), .B(n1320), .Z(n186) );
  AND U251 ( .A(n185), .B(n186), .Z(n1324) );
  XOR U252 ( .A(sreg[444]), .B(n1329), .Z(n187) );
  NANDN U253 ( .A(n1330), .B(n187), .Z(n188) );
  NAND U254 ( .A(sreg[444]), .B(n1329), .Z(n189) );
  AND U255 ( .A(n188), .B(n189), .Z(n1333) );
  XOR U256 ( .A(sreg[447]), .B(n1338), .Z(n190) );
  NANDN U257 ( .A(n1339), .B(n190), .Z(n191) );
  NAND U258 ( .A(sreg[447]), .B(n1338), .Z(n192) );
  AND U259 ( .A(n191), .B(n192), .Z(n1342) );
  XOR U260 ( .A(sreg[450]), .B(n1347), .Z(n193) );
  NANDN U261 ( .A(n1348), .B(n193), .Z(n194) );
  NAND U262 ( .A(sreg[450]), .B(n1347), .Z(n195) );
  AND U263 ( .A(n194), .B(n195), .Z(n1351) );
  XOR U264 ( .A(sreg[453]), .B(n1356), .Z(n196) );
  NANDN U265 ( .A(n1357), .B(n196), .Z(n197) );
  NAND U266 ( .A(sreg[453]), .B(n1356), .Z(n198) );
  AND U267 ( .A(n197), .B(n198), .Z(n1360) );
  XOR U268 ( .A(sreg[456]), .B(n1365), .Z(n199) );
  NANDN U269 ( .A(n1366), .B(n199), .Z(n200) );
  NAND U270 ( .A(sreg[456]), .B(n1365), .Z(n201) );
  AND U271 ( .A(n200), .B(n201), .Z(n1369) );
  XOR U272 ( .A(sreg[459]), .B(n1374), .Z(n202) );
  NANDN U273 ( .A(n1375), .B(n202), .Z(n203) );
  NAND U274 ( .A(sreg[459]), .B(n1374), .Z(n204) );
  AND U275 ( .A(n203), .B(n204), .Z(n1378) );
  XOR U276 ( .A(sreg[462]), .B(n1383), .Z(n205) );
  NANDN U277 ( .A(n1384), .B(n205), .Z(n206) );
  NAND U278 ( .A(sreg[462]), .B(n1383), .Z(n207) );
  AND U279 ( .A(n206), .B(n207), .Z(n1387) );
  XOR U280 ( .A(sreg[465]), .B(n1392), .Z(n208) );
  NANDN U281 ( .A(n1393), .B(n208), .Z(n209) );
  NAND U282 ( .A(sreg[465]), .B(n1392), .Z(n210) );
  AND U283 ( .A(n209), .B(n210), .Z(n1396) );
  XOR U284 ( .A(sreg[468]), .B(n1401), .Z(n211) );
  NANDN U285 ( .A(n1402), .B(n211), .Z(n212) );
  NAND U286 ( .A(sreg[468]), .B(n1401), .Z(n213) );
  AND U287 ( .A(n212), .B(n213), .Z(n1405) );
  XOR U288 ( .A(sreg[471]), .B(n1410), .Z(n214) );
  NANDN U289 ( .A(n1411), .B(n214), .Z(n215) );
  NAND U290 ( .A(sreg[471]), .B(n1410), .Z(n216) );
  AND U291 ( .A(n215), .B(n216), .Z(n1414) );
  XOR U292 ( .A(sreg[474]), .B(n1419), .Z(n217) );
  NANDN U293 ( .A(n1420), .B(n217), .Z(n218) );
  NAND U294 ( .A(sreg[474]), .B(n1419), .Z(n219) );
  AND U295 ( .A(n218), .B(n219), .Z(n1423) );
  XOR U296 ( .A(sreg[477]), .B(n1428), .Z(n220) );
  NANDN U297 ( .A(n1429), .B(n220), .Z(n221) );
  NAND U298 ( .A(sreg[477]), .B(n1428), .Z(n222) );
  AND U299 ( .A(n221), .B(n222), .Z(n1432) );
  XOR U300 ( .A(sreg[480]), .B(n1437), .Z(n223) );
  NANDN U301 ( .A(n1438), .B(n223), .Z(n224) );
  NAND U302 ( .A(sreg[480]), .B(n1437), .Z(n225) );
  AND U303 ( .A(n224), .B(n225), .Z(n1441) );
  XOR U304 ( .A(sreg[483]), .B(n1446), .Z(n226) );
  NANDN U305 ( .A(n1447), .B(n226), .Z(n227) );
  NAND U306 ( .A(sreg[483]), .B(n1446), .Z(n228) );
  AND U307 ( .A(n227), .B(n228), .Z(n1450) );
  XOR U308 ( .A(sreg[486]), .B(n1455), .Z(n229) );
  NANDN U309 ( .A(n1456), .B(n229), .Z(n230) );
  NAND U310 ( .A(sreg[486]), .B(n1455), .Z(n231) );
  AND U311 ( .A(n230), .B(n231), .Z(n1459) );
  XOR U312 ( .A(sreg[489]), .B(n1464), .Z(n232) );
  NANDN U313 ( .A(n1465), .B(n232), .Z(n233) );
  NAND U314 ( .A(sreg[489]), .B(n1464), .Z(n234) );
  AND U315 ( .A(n233), .B(n234), .Z(n1468) );
  XOR U316 ( .A(sreg[492]), .B(n1473), .Z(n235) );
  NANDN U317 ( .A(n1474), .B(n235), .Z(n236) );
  NAND U318 ( .A(sreg[492]), .B(n1473), .Z(n237) );
  AND U319 ( .A(n236), .B(n237), .Z(n1477) );
  XOR U320 ( .A(sreg[495]), .B(n1482), .Z(n238) );
  NANDN U321 ( .A(n1483), .B(n238), .Z(n239) );
  NAND U322 ( .A(sreg[495]), .B(n1482), .Z(n240) );
  AND U323 ( .A(n239), .B(n240), .Z(n1486) );
  XOR U324 ( .A(sreg[498]), .B(n1491), .Z(n241) );
  NANDN U325 ( .A(n1492), .B(n241), .Z(n242) );
  NAND U326 ( .A(sreg[498]), .B(n1491), .Z(n243) );
  AND U327 ( .A(n242), .B(n243), .Z(n1495) );
  XOR U328 ( .A(sreg[501]), .B(n1500), .Z(n244) );
  NANDN U329 ( .A(n1501), .B(n244), .Z(n245) );
  NAND U330 ( .A(sreg[501]), .B(n1500), .Z(n246) );
  AND U331 ( .A(n245), .B(n246), .Z(n1504) );
  XOR U332 ( .A(sreg[504]), .B(n1509), .Z(n247) );
  NANDN U333 ( .A(n1510), .B(n247), .Z(n248) );
  NAND U334 ( .A(sreg[504]), .B(n1509), .Z(n249) );
  AND U335 ( .A(n248), .B(n249), .Z(n1513) );
  XOR U336 ( .A(sreg[507]), .B(n1518), .Z(n250) );
  NANDN U337 ( .A(n1519), .B(n250), .Z(n251) );
  NAND U338 ( .A(sreg[507]), .B(n1518), .Z(n252) );
  AND U339 ( .A(n251), .B(n252), .Z(n1522) );
  XOR U340 ( .A(n765), .B(sreg[256]), .Z(n253) );
  NANDN U341 ( .A(n766), .B(n253), .Z(n254) );
  NAND U342 ( .A(n765), .B(sreg[256]), .Z(n255) );
  AND U343 ( .A(n254), .B(n255), .Z(n769) );
  XOR U344 ( .A(sreg[259]), .B(n774), .Z(n256) );
  NANDN U345 ( .A(n775), .B(n256), .Z(n257) );
  NAND U346 ( .A(sreg[259]), .B(n774), .Z(n258) );
  AND U347 ( .A(n257), .B(n258), .Z(n778) );
  XOR U348 ( .A(sreg[262]), .B(n783), .Z(n259) );
  NANDN U349 ( .A(n784), .B(n259), .Z(n260) );
  NAND U350 ( .A(sreg[262]), .B(n783), .Z(n261) );
  AND U351 ( .A(n260), .B(n261), .Z(n787) );
  XOR U352 ( .A(sreg[265]), .B(n792), .Z(n262) );
  NANDN U353 ( .A(n793), .B(n262), .Z(n263) );
  NAND U354 ( .A(sreg[265]), .B(n792), .Z(n264) );
  AND U355 ( .A(n263), .B(n264), .Z(n796) );
  XOR U356 ( .A(sreg[268]), .B(n801), .Z(n265) );
  NANDN U357 ( .A(n802), .B(n265), .Z(n266) );
  NAND U358 ( .A(sreg[268]), .B(n801), .Z(n267) );
  AND U359 ( .A(n266), .B(n267), .Z(n805) );
  XOR U360 ( .A(sreg[271]), .B(n810), .Z(n268) );
  NANDN U361 ( .A(n811), .B(n268), .Z(n269) );
  NAND U362 ( .A(sreg[271]), .B(n810), .Z(n270) );
  AND U363 ( .A(n269), .B(n270), .Z(n814) );
  XOR U364 ( .A(sreg[274]), .B(n819), .Z(n271) );
  NANDN U365 ( .A(n820), .B(n271), .Z(n272) );
  NAND U366 ( .A(sreg[274]), .B(n819), .Z(n273) );
  AND U367 ( .A(n272), .B(n273), .Z(n823) );
  XOR U368 ( .A(sreg[277]), .B(n828), .Z(n274) );
  NANDN U369 ( .A(n829), .B(n274), .Z(n275) );
  NAND U370 ( .A(sreg[277]), .B(n828), .Z(n276) );
  AND U371 ( .A(n275), .B(n276), .Z(n832) );
  XOR U372 ( .A(sreg[280]), .B(n837), .Z(n277) );
  NANDN U373 ( .A(n838), .B(n277), .Z(n278) );
  NAND U374 ( .A(sreg[280]), .B(n837), .Z(n279) );
  AND U375 ( .A(n278), .B(n279), .Z(n841) );
  XOR U376 ( .A(sreg[283]), .B(n846), .Z(n280) );
  NANDN U377 ( .A(n847), .B(n280), .Z(n281) );
  NAND U378 ( .A(sreg[283]), .B(n846), .Z(n282) );
  AND U379 ( .A(n281), .B(n282), .Z(n850) );
  XOR U380 ( .A(sreg[286]), .B(n855), .Z(n283) );
  NANDN U381 ( .A(n856), .B(n283), .Z(n284) );
  NAND U382 ( .A(sreg[286]), .B(n855), .Z(n285) );
  AND U383 ( .A(n284), .B(n285), .Z(n859) );
  XOR U384 ( .A(sreg[289]), .B(n864), .Z(n286) );
  NANDN U385 ( .A(n865), .B(n286), .Z(n287) );
  NAND U386 ( .A(sreg[289]), .B(n864), .Z(n288) );
  AND U387 ( .A(n287), .B(n288), .Z(n868) );
  XOR U388 ( .A(sreg[292]), .B(n873), .Z(n289) );
  NANDN U389 ( .A(n874), .B(n289), .Z(n290) );
  NAND U390 ( .A(sreg[292]), .B(n873), .Z(n291) );
  AND U391 ( .A(n290), .B(n291), .Z(n877) );
  XOR U392 ( .A(sreg[295]), .B(n882), .Z(n292) );
  NANDN U393 ( .A(n883), .B(n292), .Z(n293) );
  NAND U394 ( .A(sreg[295]), .B(n882), .Z(n294) );
  AND U395 ( .A(n293), .B(n294), .Z(n886) );
  XOR U396 ( .A(sreg[298]), .B(n891), .Z(n295) );
  NANDN U397 ( .A(n892), .B(n295), .Z(n296) );
  NAND U398 ( .A(sreg[298]), .B(n891), .Z(n297) );
  AND U399 ( .A(n296), .B(n297), .Z(n895) );
  XOR U400 ( .A(sreg[301]), .B(n900), .Z(n298) );
  NANDN U401 ( .A(n901), .B(n298), .Z(n299) );
  NAND U402 ( .A(sreg[301]), .B(n900), .Z(n300) );
  AND U403 ( .A(n299), .B(n300), .Z(n904) );
  XOR U404 ( .A(sreg[304]), .B(n909), .Z(n301) );
  NANDN U405 ( .A(n910), .B(n301), .Z(n302) );
  NAND U406 ( .A(sreg[304]), .B(n909), .Z(n303) );
  AND U407 ( .A(n302), .B(n303), .Z(n913) );
  XOR U408 ( .A(sreg[307]), .B(n918), .Z(n304) );
  NANDN U409 ( .A(n919), .B(n304), .Z(n305) );
  NAND U410 ( .A(sreg[307]), .B(n918), .Z(n306) );
  AND U411 ( .A(n305), .B(n306), .Z(n922) );
  XOR U412 ( .A(sreg[310]), .B(n927), .Z(n307) );
  NANDN U413 ( .A(n928), .B(n307), .Z(n308) );
  NAND U414 ( .A(sreg[310]), .B(n927), .Z(n309) );
  AND U415 ( .A(n308), .B(n309), .Z(n931) );
  XOR U416 ( .A(sreg[313]), .B(n936), .Z(n310) );
  NANDN U417 ( .A(n937), .B(n310), .Z(n311) );
  NAND U418 ( .A(sreg[313]), .B(n936), .Z(n312) );
  AND U419 ( .A(n311), .B(n312), .Z(n940) );
  XOR U420 ( .A(sreg[316]), .B(n945), .Z(n313) );
  NANDN U421 ( .A(n946), .B(n313), .Z(n314) );
  NAND U422 ( .A(sreg[316]), .B(n945), .Z(n315) );
  AND U423 ( .A(n314), .B(n315), .Z(n949) );
  XOR U424 ( .A(sreg[319]), .B(n954), .Z(n316) );
  NANDN U425 ( .A(n955), .B(n316), .Z(n317) );
  NAND U426 ( .A(sreg[319]), .B(n954), .Z(n318) );
  AND U427 ( .A(n317), .B(n318), .Z(n958) );
  XOR U428 ( .A(sreg[322]), .B(n963), .Z(n319) );
  NANDN U429 ( .A(n964), .B(n319), .Z(n320) );
  NAND U430 ( .A(sreg[322]), .B(n963), .Z(n321) );
  AND U431 ( .A(n320), .B(n321), .Z(n967) );
  XOR U432 ( .A(sreg[325]), .B(n972), .Z(n322) );
  NANDN U433 ( .A(n973), .B(n322), .Z(n323) );
  NAND U434 ( .A(sreg[325]), .B(n972), .Z(n324) );
  AND U435 ( .A(n323), .B(n324), .Z(n976) );
  XOR U436 ( .A(sreg[328]), .B(n981), .Z(n325) );
  NANDN U437 ( .A(n982), .B(n325), .Z(n326) );
  NAND U438 ( .A(sreg[328]), .B(n981), .Z(n327) );
  AND U439 ( .A(n326), .B(n327), .Z(n985) );
  XOR U440 ( .A(sreg[331]), .B(n990), .Z(n328) );
  NANDN U441 ( .A(n991), .B(n328), .Z(n329) );
  NAND U442 ( .A(sreg[331]), .B(n990), .Z(n330) );
  AND U443 ( .A(n329), .B(n330), .Z(n994) );
  XOR U444 ( .A(sreg[334]), .B(n999), .Z(n331) );
  NANDN U445 ( .A(n1000), .B(n331), .Z(n332) );
  NAND U446 ( .A(sreg[334]), .B(n999), .Z(n333) );
  AND U447 ( .A(n332), .B(n333), .Z(n1003) );
  XOR U448 ( .A(sreg[337]), .B(n1008), .Z(n334) );
  NANDN U449 ( .A(n1009), .B(n334), .Z(n335) );
  NAND U450 ( .A(sreg[337]), .B(n1008), .Z(n336) );
  AND U451 ( .A(n335), .B(n336), .Z(n1012) );
  XOR U452 ( .A(sreg[340]), .B(n1017), .Z(n337) );
  NANDN U453 ( .A(n1018), .B(n337), .Z(n338) );
  NAND U454 ( .A(sreg[340]), .B(n1017), .Z(n339) );
  AND U455 ( .A(n338), .B(n339), .Z(n1021) );
  XOR U456 ( .A(sreg[343]), .B(n1026), .Z(n340) );
  NANDN U457 ( .A(n1027), .B(n340), .Z(n341) );
  NAND U458 ( .A(sreg[343]), .B(n1026), .Z(n342) );
  AND U459 ( .A(n341), .B(n342), .Z(n1030) );
  XOR U460 ( .A(sreg[346]), .B(n1035), .Z(n343) );
  NANDN U461 ( .A(n1036), .B(n343), .Z(n344) );
  NAND U462 ( .A(sreg[346]), .B(n1035), .Z(n345) );
  AND U463 ( .A(n344), .B(n345), .Z(n1039) );
  XOR U464 ( .A(sreg[349]), .B(n1044), .Z(n346) );
  NANDN U465 ( .A(n1045), .B(n346), .Z(n347) );
  NAND U466 ( .A(sreg[349]), .B(n1044), .Z(n348) );
  AND U467 ( .A(n347), .B(n348), .Z(n1048) );
  XOR U468 ( .A(sreg[352]), .B(n1053), .Z(n349) );
  NANDN U469 ( .A(n1054), .B(n349), .Z(n350) );
  NAND U470 ( .A(sreg[352]), .B(n1053), .Z(n351) );
  AND U471 ( .A(n350), .B(n351), .Z(n1057) );
  XOR U472 ( .A(sreg[355]), .B(n1062), .Z(n352) );
  NANDN U473 ( .A(n1063), .B(n352), .Z(n353) );
  NAND U474 ( .A(sreg[355]), .B(n1062), .Z(n354) );
  AND U475 ( .A(n353), .B(n354), .Z(n1066) );
  XOR U476 ( .A(sreg[358]), .B(n1071), .Z(n355) );
  NANDN U477 ( .A(n1072), .B(n355), .Z(n356) );
  NAND U478 ( .A(sreg[358]), .B(n1071), .Z(n357) );
  AND U479 ( .A(n356), .B(n357), .Z(n1075) );
  XOR U480 ( .A(sreg[361]), .B(n1080), .Z(n358) );
  NANDN U481 ( .A(n1081), .B(n358), .Z(n359) );
  NAND U482 ( .A(sreg[361]), .B(n1080), .Z(n360) );
  AND U483 ( .A(n359), .B(n360), .Z(n1084) );
  XOR U484 ( .A(sreg[364]), .B(n1089), .Z(n361) );
  NANDN U485 ( .A(n1090), .B(n361), .Z(n362) );
  NAND U486 ( .A(sreg[364]), .B(n1089), .Z(n363) );
  AND U487 ( .A(n362), .B(n363), .Z(n1093) );
  XOR U488 ( .A(sreg[367]), .B(n1098), .Z(n364) );
  NANDN U489 ( .A(n1099), .B(n364), .Z(n365) );
  NAND U490 ( .A(sreg[367]), .B(n1098), .Z(n366) );
  AND U491 ( .A(n365), .B(n366), .Z(n1102) );
  XOR U492 ( .A(sreg[370]), .B(n1107), .Z(n367) );
  NANDN U493 ( .A(n1108), .B(n367), .Z(n368) );
  NAND U494 ( .A(sreg[370]), .B(n1107), .Z(n369) );
  AND U495 ( .A(n368), .B(n369), .Z(n1111) );
  XOR U496 ( .A(sreg[373]), .B(n1116), .Z(n370) );
  NANDN U497 ( .A(n1117), .B(n370), .Z(n371) );
  NAND U498 ( .A(sreg[373]), .B(n1116), .Z(n372) );
  AND U499 ( .A(n371), .B(n372), .Z(n1120) );
  XOR U500 ( .A(sreg[376]), .B(n1125), .Z(n373) );
  NANDN U501 ( .A(n1126), .B(n373), .Z(n374) );
  NAND U502 ( .A(sreg[376]), .B(n1125), .Z(n375) );
  AND U503 ( .A(n374), .B(n375), .Z(n1129) );
  XOR U504 ( .A(sreg[379]), .B(n1134), .Z(n376) );
  NANDN U505 ( .A(n1135), .B(n376), .Z(n377) );
  NAND U506 ( .A(sreg[379]), .B(n1134), .Z(n378) );
  AND U507 ( .A(n377), .B(n378), .Z(n1138) );
  XOR U508 ( .A(sreg[382]), .B(n1143), .Z(n379) );
  NANDN U509 ( .A(n1144), .B(n379), .Z(n380) );
  NAND U510 ( .A(sreg[382]), .B(n1143), .Z(n381) );
  AND U511 ( .A(n380), .B(n381), .Z(n1147) );
  XOR U512 ( .A(sreg[385]), .B(n1152), .Z(n382) );
  NANDN U513 ( .A(n1153), .B(n382), .Z(n383) );
  NAND U514 ( .A(sreg[385]), .B(n1152), .Z(n384) );
  AND U515 ( .A(n383), .B(n384), .Z(n1156) );
  XOR U516 ( .A(sreg[388]), .B(n1161), .Z(n385) );
  NANDN U517 ( .A(n1162), .B(n385), .Z(n386) );
  NAND U518 ( .A(sreg[388]), .B(n1161), .Z(n387) );
  AND U519 ( .A(n386), .B(n387), .Z(n1165) );
  XOR U520 ( .A(sreg[391]), .B(n1170), .Z(n388) );
  NANDN U521 ( .A(n1171), .B(n388), .Z(n389) );
  NAND U522 ( .A(sreg[391]), .B(n1170), .Z(n390) );
  AND U523 ( .A(n389), .B(n390), .Z(n1174) );
  XOR U524 ( .A(sreg[394]), .B(n1179), .Z(n391) );
  NANDN U525 ( .A(n1180), .B(n391), .Z(n392) );
  NAND U526 ( .A(sreg[394]), .B(n1179), .Z(n393) );
  AND U527 ( .A(n392), .B(n393), .Z(n1183) );
  XOR U528 ( .A(sreg[397]), .B(n1188), .Z(n394) );
  NANDN U529 ( .A(n1189), .B(n394), .Z(n395) );
  NAND U530 ( .A(sreg[397]), .B(n1188), .Z(n396) );
  AND U531 ( .A(n395), .B(n396), .Z(n1192) );
  XOR U532 ( .A(sreg[400]), .B(n1197), .Z(n397) );
  NANDN U533 ( .A(n1198), .B(n397), .Z(n398) );
  NAND U534 ( .A(sreg[400]), .B(n1197), .Z(n399) );
  AND U535 ( .A(n398), .B(n399), .Z(n1201) );
  XOR U536 ( .A(sreg[403]), .B(n1206), .Z(n400) );
  NANDN U537 ( .A(n1207), .B(n400), .Z(n401) );
  NAND U538 ( .A(sreg[403]), .B(n1206), .Z(n402) );
  AND U539 ( .A(n401), .B(n402), .Z(n1210) );
  XOR U540 ( .A(sreg[406]), .B(n1215), .Z(n403) );
  NANDN U541 ( .A(n1216), .B(n403), .Z(n404) );
  NAND U542 ( .A(sreg[406]), .B(n1215), .Z(n405) );
  AND U543 ( .A(n404), .B(n405), .Z(n1219) );
  XOR U544 ( .A(sreg[409]), .B(n1224), .Z(n406) );
  NANDN U545 ( .A(n1225), .B(n406), .Z(n407) );
  NAND U546 ( .A(sreg[409]), .B(n1224), .Z(n408) );
  AND U547 ( .A(n407), .B(n408), .Z(n1228) );
  XOR U548 ( .A(sreg[412]), .B(n1233), .Z(n409) );
  NANDN U549 ( .A(n1234), .B(n409), .Z(n410) );
  NAND U550 ( .A(sreg[412]), .B(n1233), .Z(n411) );
  AND U551 ( .A(n410), .B(n411), .Z(n1237) );
  XOR U552 ( .A(sreg[415]), .B(n1242), .Z(n412) );
  NANDN U553 ( .A(n1243), .B(n412), .Z(n413) );
  NAND U554 ( .A(sreg[415]), .B(n1242), .Z(n414) );
  AND U555 ( .A(n413), .B(n414), .Z(n1246) );
  XOR U556 ( .A(sreg[418]), .B(n1251), .Z(n415) );
  NANDN U557 ( .A(n1252), .B(n415), .Z(n416) );
  NAND U558 ( .A(sreg[418]), .B(n1251), .Z(n417) );
  AND U559 ( .A(n416), .B(n417), .Z(n1255) );
  XOR U560 ( .A(sreg[421]), .B(n1260), .Z(n418) );
  NANDN U561 ( .A(n1261), .B(n418), .Z(n419) );
  NAND U562 ( .A(sreg[421]), .B(n1260), .Z(n420) );
  AND U563 ( .A(n419), .B(n420), .Z(n1264) );
  XOR U564 ( .A(sreg[424]), .B(n1269), .Z(n421) );
  NANDN U565 ( .A(n1270), .B(n421), .Z(n422) );
  NAND U566 ( .A(sreg[424]), .B(n1269), .Z(n423) );
  AND U567 ( .A(n422), .B(n423), .Z(n1273) );
  XOR U568 ( .A(sreg[427]), .B(n1278), .Z(n424) );
  NANDN U569 ( .A(n1279), .B(n424), .Z(n425) );
  NAND U570 ( .A(sreg[427]), .B(n1278), .Z(n426) );
  AND U571 ( .A(n425), .B(n426), .Z(n1282) );
  XOR U572 ( .A(sreg[430]), .B(n1287), .Z(n427) );
  NANDN U573 ( .A(n1288), .B(n427), .Z(n428) );
  NAND U574 ( .A(sreg[430]), .B(n1287), .Z(n429) );
  AND U575 ( .A(n428), .B(n429), .Z(n1291) );
  XOR U576 ( .A(sreg[433]), .B(n1296), .Z(n430) );
  NANDN U577 ( .A(n1297), .B(n430), .Z(n431) );
  NAND U578 ( .A(sreg[433]), .B(n1296), .Z(n432) );
  AND U579 ( .A(n431), .B(n432), .Z(n1300) );
  XOR U580 ( .A(sreg[436]), .B(n1305), .Z(n433) );
  NANDN U581 ( .A(n1306), .B(n433), .Z(n434) );
  NAND U582 ( .A(sreg[436]), .B(n1305), .Z(n435) );
  AND U583 ( .A(n434), .B(n435), .Z(n1309) );
  XOR U584 ( .A(sreg[439]), .B(n1314), .Z(n436) );
  NANDN U585 ( .A(n1315), .B(n436), .Z(n437) );
  NAND U586 ( .A(sreg[439]), .B(n1314), .Z(n438) );
  AND U587 ( .A(n437), .B(n438), .Z(n1318) );
  XOR U588 ( .A(sreg[442]), .B(n1323), .Z(n439) );
  NANDN U589 ( .A(n1324), .B(n439), .Z(n440) );
  NAND U590 ( .A(sreg[442]), .B(n1323), .Z(n441) );
  AND U591 ( .A(n440), .B(n441), .Z(n1327) );
  XOR U592 ( .A(sreg[445]), .B(n1332), .Z(n442) );
  NANDN U593 ( .A(n1333), .B(n442), .Z(n443) );
  NAND U594 ( .A(sreg[445]), .B(n1332), .Z(n444) );
  AND U595 ( .A(n443), .B(n444), .Z(n1336) );
  XOR U596 ( .A(sreg[448]), .B(n1341), .Z(n445) );
  NANDN U597 ( .A(n1342), .B(n445), .Z(n446) );
  NAND U598 ( .A(sreg[448]), .B(n1341), .Z(n447) );
  AND U599 ( .A(n446), .B(n447), .Z(n1345) );
  XOR U600 ( .A(sreg[451]), .B(n1350), .Z(n448) );
  NANDN U601 ( .A(n1351), .B(n448), .Z(n449) );
  NAND U602 ( .A(sreg[451]), .B(n1350), .Z(n450) );
  AND U603 ( .A(n449), .B(n450), .Z(n1354) );
  XOR U604 ( .A(sreg[454]), .B(n1359), .Z(n451) );
  NANDN U605 ( .A(n1360), .B(n451), .Z(n452) );
  NAND U606 ( .A(sreg[454]), .B(n1359), .Z(n453) );
  AND U607 ( .A(n452), .B(n453), .Z(n1363) );
  XOR U608 ( .A(sreg[457]), .B(n1368), .Z(n454) );
  NANDN U609 ( .A(n1369), .B(n454), .Z(n455) );
  NAND U610 ( .A(sreg[457]), .B(n1368), .Z(n456) );
  AND U611 ( .A(n455), .B(n456), .Z(n1372) );
  XOR U612 ( .A(sreg[460]), .B(n1377), .Z(n457) );
  NANDN U613 ( .A(n1378), .B(n457), .Z(n458) );
  NAND U614 ( .A(sreg[460]), .B(n1377), .Z(n459) );
  AND U615 ( .A(n458), .B(n459), .Z(n1381) );
  XOR U616 ( .A(sreg[463]), .B(n1386), .Z(n460) );
  NANDN U617 ( .A(n1387), .B(n460), .Z(n461) );
  NAND U618 ( .A(sreg[463]), .B(n1386), .Z(n462) );
  AND U619 ( .A(n461), .B(n462), .Z(n1390) );
  XOR U620 ( .A(sreg[466]), .B(n1395), .Z(n463) );
  NANDN U621 ( .A(n1396), .B(n463), .Z(n464) );
  NAND U622 ( .A(sreg[466]), .B(n1395), .Z(n465) );
  AND U623 ( .A(n464), .B(n465), .Z(n1399) );
  XOR U624 ( .A(sreg[469]), .B(n1404), .Z(n466) );
  NANDN U625 ( .A(n1405), .B(n466), .Z(n467) );
  NAND U626 ( .A(sreg[469]), .B(n1404), .Z(n468) );
  AND U627 ( .A(n467), .B(n468), .Z(n1408) );
  XOR U628 ( .A(sreg[472]), .B(n1413), .Z(n469) );
  NANDN U629 ( .A(n1414), .B(n469), .Z(n470) );
  NAND U630 ( .A(sreg[472]), .B(n1413), .Z(n471) );
  AND U631 ( .A(n470), .B(n471), .Z(n1417) );
  XOR U632 ( .A(sreg[475]), .B(n1422), .Z(n472) );
  NANDN U633 ( .A(n1423), .B(n472), .Z(n473) );
  NAND U634 ( .A(sreg[475]), .B(n1422), .Z(n474) );
  AND U635 ( .A(n473), .B(n474), .Z(n1426) );
  XOR U636 ( .A(sreg[478]), .B(n1431), .Z(n475) );
  NANDN U637 ( .A(n1432), .B(n475), .Z(n476) );
  NAND U638 ( .A(sreg[478]), .B(n1431), .Z(n477) );
  AND U639 ( .A(n476), .B(n477), .Z(n1435) );
  XOR U640 ( .A(sreg[481]), .B(n1440), .Z(n478) );
  NANDN U641 ( .A(n1441), .B(n478), .Z(n479) );
  NAND U642 ( .A(sreg[481]), .B(n1440), .Z(n480) );
  AND U643 ( .A(n479), .B(n480), .Z(n1444) );
  XOR U644 ( .A(sreg[484]), .B(n1449), .Z(n481) );
  NANDN U645 ( .A(n1450), .B(n481), .Z(n482) );
  NAND U646 ( .A(sreg[484]), .B(n1449), .Z(n483) );
  AND U647 ( .A(n482), .B(n483), .Z(n1453) );
  XOR U648 ( .A(sreg[487]), .B(n1458), .Z(n484) );
  NANDN U649 ( .A(n1459), .B(n484), .Z(n485) );
  NAND U650 ( .A(sreg[487]), .B(n1458), .Z(n486) );
  AND U651 ( .A(n485), .B(n486), .Z(n1462) );
  XOR U652 ( .A(sreg[490]), .B(n1467), .Z(n487) );
  NANDN U653 ( .A(n1468), .B(n487), .Z(n488) );
  NAND U654 ( .A(sreg[490]), .B(n1467), .Z(n489) );
  AND U655 ( .A(n488), .B(n489), .Z(n1471) );
  XOR U656 ( .A(sreg[493]), .B(n1476), .Z(n490) );
  NANDN U657 ( .A(n1477), .B(n490), .Z(n491) );
  NAND U658 ( .A(sreg[493]), .B(n1476), .Z(n492) );
  AND U659 ( .A(n491), .B(n492), .Z(n1480) );
  XOR U660 ( .A(sreg[496]), .B(n1485), .Z(n493) );
  NANDN U661 ( .A(n1486), .B(n493), .Z(n494) );
  NAND U662 ( .A(sreg[496]), .B(n1485), .Z(n495) );
  AND U663 ( .A(n494), .B(n495), .Z(n1489) );
  XOR U664 ( .A(sreg[499]), .B(n1494), .Z(n496) );
  NANDN U665 ( .A(n1495), .B(n496), .Z(n497) );
  NAND U666 ( .A(sreg[499]), .B(n1494), .Z(n498) );
  AND U667 ( .A(n497), .B(n498), .Z(n1498) );
  XOR U668 ( .A(sreg[502]), .B(n1503), .Z(n499) );
  NANDN U669 ( .A(n1504), .B(n499), .Z(n500) );
  NAND U670 ( .A(sreg[502]), .B(n1503), .Z(n501) );
  AND U671 ( .A(n500), .B(n501), .Z(n1507) );
  XOR U672 ( .A(sreg[505]), .B(n1512), .Z(n502) );
  NANDN U673 ( .A(n1513), .B(n502), .Z(n503) );
  NAND U674 ( .A(sreg[505]), .B(n1512), .Z(n504) );
  AND U675 ( .A(n503), .B(n504), .Z(n1516) );
  XOR U676 ( .A(sreg[508]), .B(n1521), .Z(n505) );
  NANDN U677 ( .A(n1522), .B(n505), .Z(n506) );
  NAND U678 ( .A(sreg[508]), .B(n1521), .Z(n507) );
  AND U679 ( .A(n506), .B(n507), .Z(n1525) );
  XOR U680 ( .A(sreg[257]), .B(n768), .Z(n508) );
  NANDN U681 ( .A(n769), .B(n508), .Z(n509) );
  NAND U682 ( .A(sreg[257]), .B(n768), .Z(n510) );
  AND U683 ( .A(n509), .B(n510), .Z(n772) );
  XOR U684 ( .A(sreg[260]), .B(n777), .Z(n511) );
  NANDN U685 ( .A(n778), .B(n511), .Z(n512) );
  NAND U686 ( .A(sreg[260]), .B(n777), .Z(n513) );
  AND U687 ( .A(n512), .B(n513), .Z(n781) );
  XOR U688 ( .A(sreg[263]), .B(n786), .Z(n514) );
  NANDN U689 ( .A(n787), .B(n514), .Z(n515) );
  NAND U690 ( .A(sreg[263]), .B(n786), .Z(n516) );
  AND U691 ( .A(n515), .B(n516), .Z(n790) );
  XOR U692 ( .A(sreg[266]), .B(n795), .Z(n517) );
  NANDN U693 ( .A(n796), .B(n517), .Z(n518) );
  NAND U694 ( .A(sreg[266]), .B(n795), .Z(n519) );
  AND U695 ( .A(n518), .B(n519), .Z(n799) );
  XOR U696 ( .A(sreg[269]), .B(n804), .Z(n520) );
  NANDN U697 ( .A(n805), .B(n520), .Z(n521) );
  NAND U698 ( .A(sreg[269]), .B(n804), .Z(n522) );
  AND U699 ( .A(n521), .B(n522), .Z(n808) );
  XOR U700 ( .A(sreg[272]), .B(n813), .Z(n523) );
  NANDN U701 ( .A(n814), .B(n523), .Z(n524) );
  NAND U702 ( .A(sreg[272]), .B(n813), .Z(n525) );
  AND U703 ( .A(n524), .B(n525), .Z(n817) );
  XOR U704 ( .A(sreg[275]), .B(n822), .Z(n526) );
  NANDN U705 ( .A(n823), .B(n526), .Z(n527) );
  NAND U706 ( .A(sreg[275]), .B(n822), .Z(n528) );
  AND U707 ( .A(n527), .B(n528), .Z(n826) );
  XOR U708 ( .A(sreg[278]), .B(n831), .Z(n529) );
  NANDN U709 ( .A(n832), .B(n529), .Z(n530) );
  NAND U710 ( .A(sreg[278]), .B(n831), .Z(n531) );
  AND U711 ( .A(n530), .B(n531), .Z(n835) );
  XOR U712 ( .A(sreg[281]), .B(n840), .Z(n532) );
  NANDN U713 ( .A(n841), .B(n532), .Z(n533) );
  NAND U714 ( .A(sreg[281]), .B(n840), .Z(n534) );
  AND U715 ( .A(n533), .B(n534), .Z(n844) );
  XOR U716 ( .A(sreg[284]), .B(n849), .Z(n535) );
  NANDN U717 ( .A(n850), .B(n535), .Z(n536) );
  NAND U718 ( .A(sreg[284]), .B(n849), .Z(n537) );
  AND U719 ( .A(n536), .B(n537), .Z(n853) );
  XOR U720 ( .A(sreg[287]), .B(n858), .Z(n538) );
  NANDN U721 ( .A(n859), .B(n538), .Z(n539) );
  NAND U722 ( .A(sreg[287]), .B(n858), .Z(n540) );
  AND U723 ( .A(n539), .B(n540), .Z(n862) );
  XOR U724 ( .A(sreg[290]), .B(n867), .Z(n541) );
  NANDN U725 ( .A(n868), .B(n541), .Z(n542) );
  NAND U726 ( .A(sreg[290]), .B(n867), .Z(n543) );
  AND U727 ( .A(n542), .B(n543), .Z(n871) );
  XOR U728 ( .A(sreg[293]), .B(n876), .Z(n544) );
  NANDN U729 ( .A(n877), .B(n544), .Z(n545) );
  NAND U730 ( .A(sreg[293]), .B(n876), .Z(n546) );
  AND U731 ( .A(n545), .B(n546), .Z(n880) );
  XOR U732 ( .A(sreg[296]), .B(n885), .Z(n547) );
  NANDN U733 ( .A(n886), .B(n547), .Z(n548) );
  NAND U734 ( .A(sreg[296]), .B(n885), .Z(n549) );
  AND U735 ( .A(n548), .B(n549), .Z(n889) );
  XOR U736 ( .A(sreg[299]), .B(n894), .Z(n550) );
  NANDN U737 ( .A(n895), .B(n550), .Z(n551) );
  NAND U738 ( .A(sreg[299]), .B(n894), .Z(n552) );
  AND U739 ( .A(n551), .B(n552), .Z(n898) );
  XOR U740 ( .A(sreg[302]), .B(n903), .Z(n553) );
  NANDN U741 ( .A(n904), .B(n553), .Z(n554) );
  NAND U742 ( .A(sreg[302]), .B(n903), .Z(n555) );
  AND U743 ( .A(n554), .B(n555), .Z(n907) );
  XOR U744 ( .A(sreg[305]), .B(n912), .Z(n556) );
  NANDN U745 ( .A(n913), .B(n556), .Z(n557) );
  NAND U746 ( .A(sreg[305]), .B(n912), .Z(n558) );
  AND U747 ( .A(n557), .B(n558), .Z(n916) );
  XOR U748 ( .A(sreg[308]), .B(n921), .Z(n559) );
  NANDN U749 ( .A(n922), .B(n559), .Z(n560) );
  NAND U750 ( .A(sreg[308]), .B(n921), .Z(n561) );
  AND U751 ( .A(n560), .B(n561), .Z(n925) );
  XOR U752 ( .A(sreg[311]), .B(n930), .Z(n562) );
  NANDN U753 ( .A(n931), .B(n562), .Z(n563) );
  NAND U754 ( .A(sreg[311]), .B(n930), .Z(n564) );
  AND U755 ( .A(n563), .B(n564), .Z(n934) );
  XOR U756 ( .A(sreg[314]), .B(n939), .Z(n565) );
  NANDN U757 ( .A(n940), .B(n565), .Z(n566) );
  NAND U758 ( .A(sreg[314]), .B(n939), .Z(n567) );
  AND U759 ( .A(n566), .B(n567), .Z(n943) );
  XOR U760 ( .A(sreg[317]), .B(n948), .Z(n568) );
  NANDN U761 ( .A(n949), .B(n568), .Z(n569) );
  NAND U762 ( .A(sreg[317]), .B(n948), .Z(n570) );
  AND U763 ( .A(n569), .B(n570), .Z(n952) );
  XOR U764 ( .A(sreg[320]), .B(n957), .Z(n571) );
  NANDN U765 ( .A(n958), .B(n571), .Z(n572) );
  NAND U766 ( .A(sreg[320]), .B(n957), .Z(n573) );
  AND U767 ( .A(n572), .B(n573), .Z(n961) );
  XOR U768 ( .A(sreg[323]), .B(n966), .Z(n574) );
  NANDN U769 ( .A(n967), .B(n574), .Z(n575) );
  NAND U770 ( .A(sreg[323]), .B(n966), .Z(n576) );
  AND U771 ( .A(n575), .B(n576), .Z(n970) );
  XOR U772 ( .A(sreg[326]), .B(n975), .Z(n577) );
  NANDN U773 ( .A(n976), .B(n577), .Z(n578) );
  NAND U774 ( .A(sreg[326]), .B(n975), .Z(n579) );
  AND U775 ( .A(n578), .B(n579), .Z(n979) );
  XOR U776 ( .A(sreg[329]), .B(n984), .Z(n580) );
  NANDN U777 ( .A(n985), .B(n580), .Z(n581) );
  NAND U778 ( .A(sreg[329]), .B(n984), .Z(n582) );
  AND U779 ( .A(n581), .B(n582), .Z(n988) );
  XOR U780 ( .A(sreg[332]), .B(n993), .Z(n583) );
  NANDN U781 ( .A(n994), .B(n583), .Z(n584) );
  NAND U782 ( .A(sreg[332]), .B(n993), .Z(n585) );
  AND U783 ( .A(n584), .B(n585), .Z(n997) );
  XOR U784 ( .A(sreg[335]), .B(n1002), .Z(n586) );
  NANDN U785 ( .A(n1003), .B(n586), .Z(n587) );
  NAND U786 ( .A(sreg[335]), .B(n1002), .Z(n588) );
  AND U787 ( .A(n587), .B(n588), .Z(n1006) );
  XOR U788 ( .A(sreg[338]), .B(n1011), .Z(n589) );
  NANDN U789 ( .A(n1012), .B(n589), .Z(n590) );
  NAND U790 ( .A(sreg[338]), .B(n1011), .Z(n591) );
  AND U791 ( .A(n590), .B(n591), .Z(n1015) );
  XOR U792 ( .A(sreg[341]), .B(n1020), .Z(n592) );
  NANDN U793 ( .A(n1021), .B(n592), .Z(n593) );
  NAND U794 ( .A(sreg[341]), .B(n1020), .Z(n594) );
  AND U795 ( .A(n593), .B(n594), .Z(n1024) );
  XOR U796 ( .A(sreg[344]), .B(n1029), .Z(n595) );
  NANDN U797 ( .A(n1030), .B(n595), .Z(n596) );
  NAND U798 ( .A(sreg[344]), .B(n1029), .Z(n597) );
  AND U799 ( .A(n596), .B(n597), .Z(n1033) );
  XOR U800 ( .A(sreg[347]), .B(n1038), .Z(n598) );
  NANDN U801 ( .A(n1039), .B(n598), .Z(n599) );
  NAND U802 ( .A(sreg[347]), .B(n1038), .Z(n600) );
  AND U803 ( .A(n599), .B(n600), .Z(n1042) );
  XOR U804 ( .A(sreg[350]), .B(n1047), .Z(n601) );
  NANDN U805 ( .A(n1048), .B(n601), .Z(n602) );
  NAND U806 ( .A(sreg[350]), .B(n1047), .Z(n603) );
  AND U807 ( .A(n602), .B(n603), .Z(n1051) );
  XOR U808 ( .A(sreg[353]), .B(n1056), .Z(n604) );
  NANDN U809 ( .A(n1057), .B(n604), .Z(n605) );
  NAND U810 ( .A(sreg[353]), .B(n1056), .Z(n606) );
  AND U811 ( .A(n605), .B(n606), .Z(n1060) );
  XOR U812 ( .A(sreg[356]), .B(n1065), .Z(n607) );
  NANDN U813 ( .A(n1066), .B(n607), .Z(n608) );
  NAND U814 ( .A(sreg[356]), .B(n1065), .Z(n609) );
  AND U815 ( .A(n608), .B(n609), .Z(n1069) );
  XOR U816 ( .A(sreg[359]), .B(n1074), .Z(n610) );
  NANDN U817 ( .A(n1075), .B(n610), .Z(n611) );
  NAND U818 ( .A(sreg[359]), .B(n1074), .Z(n612) );
  AND U819 ( .A(n611), .B(n612), .Z(n1078) );
  XOR U820 ( .A(sreg[362]), .B(n1083), .Z(n613) );
  NANDN U821 ( .A(n1084), .B(n613), .Z(n614) );
  NAND U822 ( .A(sreg[362]), .B(n1083), .Z(n615) );
  AND U823 ( .A(n614), .B(n615), .Z(n1087) );
  XOR U824 ( .A(sreg[365]), .B(n1092), .Z(n616) );
  NANDN U825 ( .A(n1093), .B(n616), .Z(n617) );
  NAND U826 ( .A(sreg[365]), .B(n1092), .Z(n618) );
  AND U827 ( .A(n617), .B(n618), .Z(n1096) );
  XOR U828 ( .A(sreg[368]), .B(n1101), .Z(n619) );
  NANDN U829 ( .A(n1102), .B(n619), .Z(n620) );
  NAND U830 ( .A(sreg[368]), .B(n1101), .Z(n621) );
  AND U831 ( .A(n620), .B(n621), .Z(n1105) );
  XOR U832 ( .A(sreg[371]), .B(n1110), .Z(n622) );
  NANDN U833 ( .A(n1111), .B(n622), .Z(n623) );
  NAND U834 ( .A(sreg[371]), .B(n1110), .Z(n624) );
  AND U835 ( .A(n623), .B(n624), .Z(n1114) );
  XOR U836 ( .A(sreg[374]), .B(n1119), .Z(n625) );
  NANDN U837 ( .A(n1120), .B(n625), .Z(n626) );
  NAND U838 ( .A(sreg[374]), .B(n1119), .Z(n627) );
  AND U839 ( .A(n626), .B(n627), .Z(n1123) );
  XOR U840 ( .A(sreg[377]), .B(n1128), .Z(n628) );
  NANDN U841 ( .A(n1129), .B(n628), .Z(n629) );
  NAND U842 ( .A(sreg[377]), .B(n1128), .Z(n630) );
  AND U843 ( .A(n629), .B(n630), .Z(n1132) );
  XOR U844 ( .A(sreg[380]), .B(n1137), .Z(n631) );
  NANDN U845 ( .A(n1138), .B(n631), .Z(n632) );
  NAND U846 ( .A(sreg[380]), .B(n1137), .Z(n633) );
  AND U847 ( .A(n632), .B(n633), .Z(n1141) );
  XOR U848 ( .A(sreg[383]), .B(n1146), .Z(n634) );
  NANDN U849 ( .A(n1147), .B(n634), .Z(n635) );
  NAND U850 ( .A(sreg[383]), .B(n1146), .Z(n636) );
  AND U851 ( .A(n635), .B(n636), .Z(n1150) );
  XOR U852 ( .A(sreg[386]), .B(n1155), .Z(n637) );
  NANDN U853 ( .A(n1156), .B(n637), .Z(n638) );
  NAND U854 ( .A(sreg[386]), .B(n1155), .Z(n639) );
  AND U855 ( .A(n638), .B(n639), .Z(n1159) );
  XOR U856 ( .A(sreg[389]), .B(n1164), .Z(n640) );
  NANDN U857 ( .A(n1165), .B(n640), .Z(n641) );
  NAND U858 ( .A(sreg[389]), .B(n1164), .Z(n642) );
  AND U859 ( .A(n641), .B(n642), .Z(n1168) );
  XOR U860 ( .A(sreg[392]), .B(n1173), .Z(n643) );
  NANDN U861 ( .A(n1174), .B(n643), .Z(n644) );
  NAND U862 ( .A(sreg[392]), .B(n1173), .Z(n645) );
  AND U863 ( .A(n644), .B(n645), .Z(n1177) );
  XOR U864 ( .A(sreg[395]), .B(n1182), .Z(n646) );
  NANDN U865 ( .A(n1183), .B(n646), .Z(n647) );
  NAND U866 ( .A(sreg[395]), .B(n1182), .Z(n648) );
  AND U867 ( .A(n647), .B(n648), .Z(n1186) );
  XOR U868 ( .A(sreg[398]), .B(n1191), .Z(n649) );
  NANDN U869 ( .A(n1192), .B(n649), .Z(n650) );
  NAND U870 ( .A(sreg[398]), .B(n1191), .Z(n651) );
  AND U871 ( .A(n650), .B(n651), .Z(n1195) );
  XOR U872 ( .A(sreg[401]), .B(n1200), .Z(n652) );
  NANDN U873 ( .A(n1201), .B(n652), .Z(n653) );
  NAND U874 ( .A(sreg[401]), .B(n1200), .Z(n654) );
  AND U875 ( .A(n653), .B(n654), .Z(n1204) );
  XOR U876 ( .A(sreg[404]), .B(n1209), .Z(n655) );
  NANDN U877 ( .A(n1210), .B(n655), .Z(n656) );
  NAND U878 ( .A(sreg[404]), .B(n1209), .Z(n657) );
  AND U879 ( .A(n656), .B(n657), .Z(n1213) );
  XOR U880 ( .A(sreg[407]), .B(n1218), .Z(n658) );
  NANDN U881 ( .A(n1219), .B(n658), .Z(n659) );
  NAND U882 ( .A(sreg[407]), .B(n1218), .Z(n660) );
  AND U883 ( .A(n659), .B(n660), .Z(n1222) );
  XOR U884 ( .A(sreg[410]), .B(n1227), .Z(n661) );
  NANDN U885 ( .A(n1228), .B(n661), .Z(n662) );
  NAND U886 ( .A(sreg[410]), .B(n1227), .Z(n663) );
  AND U887 ( .A(n662), .B(n663), .Z(n1231) );
  XOR U888 ( .A(sreg[413]), .B(n1236), .Z(n664) );
  NANDN U889 ( .A(n1237), .B(n664), .Z(n665) );
  NAND U890 ( .A(sreg[413]), .B(n1236), .Z(n666) );
  AND U891 ( .A(n665), .B(n666), .Z(n1240) );
  XOR U892 ( .A(sreg[416]), .B(n1245), .Z(n667) );
  NANDN U893 ( .A(n1246), .B(n667), .Z(n668) );
  NAND U894 ( .A(sreg[416]), .B(n1245), .Z(n669) );
  AND U895 ( .A(n668), .B(n669), .Z(n1249) );
  XOR U896 ( .A(sreg[419]), .B(n1254), .Z(n670) );
  NANDN U897 ( .A(n1255), .B(n670), .Z(n671) );
  NAND U898 ( .A(sreg[419]), .B(n1254), .Z(n672) );
  AND U899 ( .A(n671), .B(n672), .Z(n1258) );
  XOR U900 ( .A(sreg[422]), .B(n1263), .Z(n673) );
  NANDN U901 ( .A(n1264), .B(n673), .Z(n674) );
  NAND U902 ( .A(sreg[422]), .B(n1263), .Z(n675) );
  AND U903 ( .A(n674), .B(n675), .Z(n1267) );
  XOR U904 ( .A(sreg[425]), .B(n1272), .Z(n676) );
  NANDN U905 ( .A(n1273), .B(n676), .Z(n677) );
  NAND U906 ( .A(sreg[425]), .B(n1272), .Z(n678) );
  AND U907 ( .A(n677), .B(n678), .Z(n1276) );
  XOR U908 ( .A(sreg[428]), .B(n1281), .Z(n679) );
  NANDN U909 ( .A(n1282), .B(n679), .Z(n680) );
  NAND U910 ( .A(sreg[428]), .B(n1281), .Z(n681) );
  AND U911 ( .A(n680), .B(n681), .Z(n1285) );
  XOR U912 ( .A(sreg[431]), .B(n1290), .Z(n682) );
  NANDN U913 ( .A(n1291), .B(n682), .Z(n683) );
  NAND U914 ( .A(sreg[431]), .B(n1290), .Z(n684) );
  AND U915 ( .A(n683), .B(n684), .Z(n1294) );
  XOR U916 ( .A(sreg[434]), .B(n1299), .Z(n685) );
  NANDN U917 ( .A(n1300), .B(n685), .Z(n686) );
  NAND U918 ( .A(sreg[434]), .B(n1299), .Z(n687) );
  AND U919 ( .A(n686), .B(n687), .Z(n1303) );
  XOR U920 ( .A(sreg[437]), .B(n1308), .Z(n688) );
  NANDN U921 ( .A(n1309), .B(n688), .Z(n689) );
  NAND U922 ( .A(sreg[437]), .B(n1308), .Z(n690) );
  AND U923 ( .A(n689), .B(n690), .Z(n1312) );
  XOR U924 ( .A(sreg[440]), .B(n1317), .Z(n691) );
  NANDN U925 ( .A(n1318), .B(n691), .Z(n692) );
  NAND U926 ( .A(sreg[440]), .B(n1317), .Z(n693) );
  AND U927 ( .A(n692), .B(n693), .Z(n1321) );
  XOR U928 ( .A(sreg[443]), .B(n1326), .Z(n694) );
  NANDN U929 ( .A(n1327), .B(n694), .Z(n695) );
  NAND U930 ( .A(sreg[443]), .B(n1326), .Z(n696) );
  AND U931 ( .A(n695), .B(n696), .Z(n1330) );
  XOR U932 ( .A(sreg[446]), .B(n1335), .Z(n697) );
  NANDN U933 ( .A(n1336), .B(n697), .Z(n698) );
  NAND U934 ( .A(sreg[446]), .B(n1335), .Z(n699) );
  AND U935 ( .A(n698), .B(n699), .Z(n1339) );
  XOR U936 ( .A(sreg[449]), .B(n1344), .Z(n700) );
  NANDN U937 ( .A(n1345), .B(n700), .Z(n701) );
  NAND U938 ( .A(sreg[449]), .B(n1344), .Z(n702) );
  AND U939 ( .A(n701), .B(n702), .Z(n1348) );
  XOR U940 ( .A(sreg[452]), .B(n1353), .Z(n703) );
  NANDN U941 ( .A(n1354), .B(n703), .Z(n704) );
  NAND U942 ( .A(sreg[452]), .B(n1353), .Z(n705) );
  AND U943 ( .A(n704), .B(n705), .Z(n1357) );
  XOR U944 ( .A(sreg[455]), .B(n1362), .Z(n706) );
  NANDN U945 ( .A(n1363), .B(n706), .Z(n707) );
  NAND U946 ( .A(sreg[455]), .B(n1362), .Z(n708) );
  AND U947 ( .A(n707), .B(n708), .Z(n1366) );
  XOR U948 ( .A(sreg[458]), .B(n1371), .Z(n709) );
  NANDN U949 ( .A(n1372), .B(n709), .Z(n710) );
  NAND U950 ( .A(sreg[458]), .B(n1371), .Z(n711) );
  AND U951 ( .A(n710), .B(n711), .Z(n1375) );
  XOR U952 ( .A(sreg[461]), .B(n1380), .Z(n712) );
  NANDN U953 ( .A(n1381), .B(n712), .Z(n713) );
  NAND U954 ( .A(sreg[461]), .B(n1380), .Z(n714) );
  AND U955 ( .A(n713), .B(n714), .Z(n1384) );
  XOR U956 ( .A(sreg[464]), .B(n1389), .Z(n715) );
  NANDN U957 ( .A(n1390), .B(n715), .Z(n716) );
  NAND U958 ( .A(sreg[464]), .B(n1389), .Z(n717) );
  AND U959 ( .A(n716), .B(n717), .Z(n1393) );
  XOR U960 ( .A(sreg[467]), .B(n1398), .Z(n718) );
  NANDN U961 ( .A(n1399), .B(n718), .Z(n719) );
  NAND U962 ( .A(sreg[467]), .B(n1398), .Z(n720) );
  AND U963 ( .A(n719), .B(n720), .Z(n1402) );
  XOR U964 ( .A(sreg[470]), .B(n1407), .Z(n721) );
  NANDN U965 ( .A(n1408), .B(n721), .Z(n722) );
  NAND U966 ( .A(sreg[470]), .B(n1407), .Z(n723) );
  AND U967 ( .A(n722), .B(n723), .Z(n1411) );
  XOR U968 ( .A(sreg[473]), .B(n1416), .Z(n724) );
  NANDN U969 ( .A(n1417), .B(n724), .Z(n725) );
  NAND U970 ( .A(sreg[473]), .B(n1416), .Z(n726) );
  AND U971 ( .A(n725), .B(n726), .Z(n1420) );
  XOR U972 ( .A(sreg[476]), .B(n1425), .Z(n727) );
  NANDN U973 ( .A(n1426), .B(n727), .Z(n728) );
  NAND U974 ( .A(sreg[476]), .B(n1425), .Z(n729) );
  AND U975 ( .A(n728), .B(n729), .Z(n1429) );
  XOR U976 ( .A(sreg[479]), .B(n1434), .Z(n730) );
  NANDN U977 ( .A(n1435), .B(n730), .Z(n731) );
  NAND U978 ( .A(sreg[479]), .B(n1434), .Z(n732) );
  AND U979 ( .A(n731), .B(n732), .Z(n1438) );
  XOR U980 ( .A(sreg[482]), .B(n1443), .Z(n733) );
  NANDN U981 ( .A(n1444), .B(n733), .Z(n734) );
  NAND U982 ( .A(sreg[482]), .B(n1443), .Z(n735) );
  AND U983 ( .A(n734), .B(n735), .Z(n1447) );
  XOR U984 ( .A(sreg[485]), .B(n1452), .Z(n736) );
  NANDN U985 ( .A(n1453), .B(n736), .Z(n737) );
  NAND U986 ( .A(sreg[485]), .B(n1452), .Z(n738) );
  AND U987 ( .A(n737), .B(n738), .Z(n1456) );
  XOR U988 ( .A(sreg[488]), .B(n1461), .Z(n739) );
  NANDN U989 ( .A(n1462), .B(n739), .Z(n740) );
  NAND U990 ( .A(sreg[488]), .B(n1461), .Z(n741) );
  AND U991 ( .A(n740), .B(n741), .Z(n1465) );
  XOR U992 ( .A(sreg[491]), .B(n1470), .Z(n742) );
  NANDN U993 ( .A(n1471), .B(n742), .Z(n743) );
  NAND U994 ( .A(sreg[491]), .B(n1470), .Z(n744) );
  AND U995 ( .A(n743), .B(n744), .Z(n1474) );
  XOR U996 ( .A(sreg[494]), .B(n1479), .Z(n745) );
  NANDN U997 ( .A(n1480), .B(n745), .Z(n746) );
  NAND U998 ( .A(sreg[494]), .B(n1479), .Z(n747) );
  AND U999 ( .A(n746), .B(n747), .Z(n1483) );
  XOR U1000 ( .A(sreg[497]), .B(n1488), .Z(n748) );
  NANDN U1001 ( .A(n1489), .B(n748), .Z(n749) );
  NAND U1002 ( .A(sreg[497]), .B(n1488), .Z(n750) );
  AND U1003 ( .A(n749), .B(n750), .Z(n1492) );
  XOR U1004 ( .A(sreg[500]), .B(n1497), .Z(n751) );
  NANDN U1005 ( .A(n1498), .B(n751), .Z(n752) );
  NAND U1006 ( .A(sreg[500]), .B(n1497), .Z(n753) );
  AND U1007 ( .A(n752), .B(n753), .Z(n1501) );
  XOR U1008 ( .A(sreg[503]), .B(n1506), .Z(n754) );
  NANDN U1009 ( .A(n1507), .B(n754), .Z(n755) );
  NAND U1010 ( .A(sreg[503]), .B(n1506), .Z(n756) );
  AND U1011 ( .A(n755), .B(n756), .Z(n1510) );
  XOR U1012 ( .A(sreg[506]), .B(n1515), .Z(n757) );
  NANDN U1013 ( .A(n1516), .B(n757), .Z(n758) );
  NAND U1014 ( .A(sreg[506]), .B(n1515), .Z(n759) );
  AND U1015 ( .A(n758), .B(n759), .Z(n1519) );
  XOR U1016 ( .A(sreg[509]), .B(n1524), .Z(n760) );
  NANDN U1017 ( .A(n1525), .B(n760), .Z(n761) );
  NAND U1018 ( .A(sreg[509]), .B(n1524), .Z(n762) );
  AND U1019 ( .A(n761), .B(n762), .Z(n1528) );
  AND U1020 ( .A(b[0]), .B(a[0]), .Z(n763) );
  XOR U1021 ( .A(n763), .B(sreg[255]), .Z(c[255]) );
  NAND U1022 ( .A(b[0]), .B(a[1]), .Z(n766) );
  AND U1023 ( .A(n763), .B(sreg[255]), .Z(n765) );
  XOR U1024 ( .A(sreg[256]), .B(n765), .Z(n764) );
  XNOR U1025 ( .A(n766), .B(n764), .Z(c[256]) );
  AND U1026 ( .A(b[0]), .B(a[2]), .Z(n768) );
  XNOR U1027 ( .A(n769), .B(sreg[257]), .Z(n767) );
  XOR U1028 ( .A(n768), .B(n767), .Z(c[257]) );
  AND U1029 ( .A(b[0]), .B(a[3]), .Z(n771) );
  XNOR U1030 ( .A(n772), .B(sreg[258]), .Z(n770) );
  XOR U1031 ( .A(n771), .B(n770), .Z(c[258]) );
  AND U1032 ( .A(b[0]), .B(a[4]), .Z(n774) );
  XNOR U1033 ( .A(n775), .B(sreg[259]), .Z(n773) );
  XOR U1034 ( .A(n774), .B(n773), .Z(c[259]) );
  AND U1035 ( .A(b[0]), .B(a[5]), .Z(n777) );
  XNOR U1036 ( .A(n778), .B(sreg[260]), .Z(n776) );
  XOR U1037 ( .A(n777), .B(n776), .Z(c[260]) );
  AND U1038 ( .A(b[0]), .B(a[6]), .Z(n780) );
  XNOR U1039 ( .A(n781), .B(sreg[261]), .Z(n779) );
  XOR U1040 ( .A(n780), .B(n779), .Z(c[261]) );
  AND U1041 ( .A(b[0]), .B(a[7]), .Z(n783) );
  XNOR U1042 ( .A(n784), .B(sreg[262]), .Z(n782) );
  XOR U1043 ( .A(n783), .B(n782), .Z(c[262]) );
  AND U1044 ( .A(b[0]), .B(a[8]), .Z(n786) );
  XNOR U1045 ( .A(n787), .B(sreg[263]), .Z(n785) );
  XOR U1046 ( .A(n786), .B(n785), .Z(c[263]) );
  AND U1047 ( .A(b[0]), .B(a[9]), .Z(n789) );
  XNOR U1048 ( .A(n790), .B(sreg[264]), .Z(n788) );
  XOR U1049 ( .A(n789), .B(n788), .Z(c[264]) );
  AND U1050 ( .A(b[0]), .B(a[10]), .Z(n792) );
  XNOR U1051 ( .A(n793), .B(sreg[265]), .Z(n791) );
  XOR U1052 ( .A(n792), .B(n791), .Z(c[265]) );
  AND U1053 ( .A(b[0]), .B(a[11]), .Z(n795) );
  XNOR U1054 ( .A(n796), .B(sreg[266]), .Z(n794) );
  XOR U1055 ( .A(n795), .B(n794), .Z(c[266]) );
  AND U1056 ( .A(b[0]), .B(a[12]), .Z(n798) );
  XNOR U1057 ( .A(n799), .B(sreg[267]), .Z(n797) );
  XOR U1058 ( .A(n798), .B(n797), .Z(c[267]) );
  AND U1059 ( .A(b[0]), .B(a[13]), .Z(n801) );
  XNOR U1060 ( .A(n802), .B(sreg[268]), .Z(n800) );
  XOR U1061 ( .A(n801), .B(n800), .Z(c[268]) );
  AND U1062 ( .A(b[0]), .B(a[14]), .Z(n804) );
  XNOR U1063 ( .A(n805), .B(sreg[269]), .Z(n803) );
  XOR U1064 ( .A(n804), .B(n803), .Z(c[269]) );
  AND U1065 ( .A(b[0]), .B(a[15]), .Z(n807) );
  XNOR U1066 ( .A(n808), .B(sreg[270]), .Z(n806) );
  XOR U1067 ( .A(n807), .B(n806), .Z(c[270]) );
  AND U1068 ( .A(b[0]), .B(a[16]), .Z(n810) );
  XNOR U1069 ( .A(n811), .B(sreg[271]), .Z(n809) );
  XOR U1070 ( .A(n810), .B(n809), .Z(c[271]) );
  AND U1071 ( .A(b[0]), .B(a[17]), .Z(n813) );
  XNOR U1072 ( .A(n814), .B(sreg[272]), .Z(n812) );
  XOR U1073 ( .A(n813), .B(n812), .Z(c[272]) );
  AND U1074 ( .A(b[0]), .B(a[18]), .Z(n816) );
  XNOR U1075 ( .A(n817), .B(sreg[273]), .Z(n815) );
  XOR U1076 ( .A(n816), .B(n815), .Z(c[273]) );
  AND U1077 ( .A(b[0]), .B(a[19]), .Z(n819) );
  XNOR U1078 ( .A(n820), .B(sreg[274]), .Z(n818) );
  XOR U1079 ( .A(n819), .B(n818), .Z(c[274]) );
  AND U1080 ( .A(b[0]), .B(a[20]), .Z(n822) );
  XNOR U1081 ( .A(n823), .B(sreg[275]), .Z(n821) );
  XOR U1082 ( .A(n822), .B(n821), .Z(c[275]) );
  AND U1083 ( .A(b[0]), .B(a[21]), .Z(n825) );
  XNOR U1084 ( .A(n826), .B(sreg[276]), .Z(n824) );
  XOR U1085 ( .A(n825), .B(n824), .Z(c[276]) );
  AND U1086 ( .A(b[0]), .B(a[22]), .Z(n828) );
  XNOR U1087 ( .A(n829), .B(sreg[277]), .Z(n827) );
  XOR U1088 ( .A(n828), .B(n827), .Z(c[277]) );
  AND U1089 ( .A(b[0]), .B(a[23]), .Z(n831) );
  XNOR U1090 ( .A(n832), .B(sreg[278]), .Z(n830) );
  XOR U1091 ( .A(n831), .B(n830), .Z(c[278]) );
  AND U1092 ( .A(b[0]), .B(a[24]), .Z(n834) );
  XNOR U1093 ( .A(n835), .B(sreg[279]), .Z(n833) );
  XOR U1094 ( .A(n834), .B(n833), .Z(c[279]) );
  AND U1095 ( .A(b[0]), .B(a[25]), .Z(n837) );
  XNOR U1096 ( .A(n838), .B(sreg[280]), .Z(n836) );
  XOR U1097 ( .A(n837), .B(n836), .Z(c[280]) );
  AND U1098 ( .A(b[0]), .B(a[26]), .Z(n840) );
  XNOR U1099 ( .A(n841), .B(sreg[281]), .Z(n839) );
  XOR U1100 ( .A(n840), .B(n839), .Z(c[281]) );
  AND U1101 ( .A(b[0]), .B(a[27]), .Z(n843) );
  XNOR U1102 ( .A(n844), .B(sreg[282]), .Z(n842) );
  XOR U1103 ( .A(n843), .B(n842), .Z(c[282]) );
  AND U1104 ( .A(b[0]), .B(a[28]), .Z(n846) );
  XNOR U1105 ( .A(n847), .B(sreg[283]), .Z(n845) );
  XOR U1106 ( .A(n846), .B(n845), .Z(c[283]) );
  AND U1107 ( .A(b[0]), .B(a[29]), .Z(n849) );
  XNOR U1108 ( .A(n850), .B(sreg[284]), .Z(n848) );
  XOR U1109 ( .A(n849), .B(n848), .Z(c[284]) );
  AND U1110 ( .A(b[0]), .B(a[30]), .Z(n852) );
  XNOR U1111 ( .A(n853), .B(sreg[285]), .Z(n851) );
  XOR U1112 ( .A(n852), .B(n851), .Z(c[285]) );
  AND U1113 ( .A(b[0]), .B(a[31]), .Z(n855) );
  XNOR U1114 ( .A(n856), .B(sreg[286]), .Z(n854) );
  XOR U1115 ( .A(n855), .B(n854), .Z(c[286]) );
  AND U1116 ( .A(b[0]), .B(a[32]), .Z(n858) );
  XNOR U1117 ( .A(n859), .B(sreg[287]), .Z(n857) );
  XOR U1118 ( .A(n858), .B(n857), .Z(c[287]) );
  AND U1119 ( .A(b[0]), .B(a[33]), .Z(n861) );
  XNOR U1120 ( .A(n862), .B(sreg[288]), .Z(n860) );
  XOR U1121 ( .A(n861), .B(n860), .Z(c[288]) );
  AND U1122 ( .A(b[0]), .B(a[34]), .Z(n864) );
  XNOR U1123 ( .A(n865), .B(sreg[289]), .Z(n863) );
  XOR U1124 ( .A(n864), .B(n863), .Z(c[289]) );
  AND U1125 ( .A(b[0]), .B(a[35]), .Z(n867) );
  XNOR U1126 ( .A(n868), .B(sreg[290]), .Z(n866) );
  XOR U1127 ( .A(n867), .B(n866), .Z(c[290]) );
  AND U1128 ( .A(b[0]), .B(a[36]), .Z(n870) );
  XNOR U1129 ( .A(n871), .B(sreg[291]), .Z(n869) );
  XOR U1130 ( .A(n870), .B(n869), .Z(c[291]) );
  AND U1131 ( .A(b[0]), .B(a[37]), .Z(n873) );
  XNOR U1132 ( .A(n874), .B(sreg[292]), .Z(n872) );
  XOR U1133 ( .A(n873), .B(n872), .Z(c[292]) );
  AND U1134 ( .A(b[0]), .B(a[38]), .Z(n876) );
  XNOR U1135 ( .A(n877), .B(sreg[293]), .Z(n875) );
  XOR U1136 ( .A(n876), .B(n875), .Z(c[293]) );
  AND U1137 ( .A(b[0]), .B(a[39]), .Z(n879) );
  XNOR U1138 ( .A(n880), .B(sreg[294]), .Z(n878) );
  XOR U1139 ( .A(n879), .B(n878), .Z(c[294]) );
  AND U1140 ( .A(b[0]), .B(a[40]), .Z(n882) );
  XNOR U1141 ( .A(n883), .B(sreg[295]), .Z(n881) );
  XOR U1142 ( .A(n882), .B(n881), .Z(c[295]) );
  AND U1143 ( .A(b[0]), .B(a[41]), .Z(n885) );
  XNOR U1144 ( .A(n886), .B(sreg[296]), .Z(n884) );
  XOR U1145 ( .A(n885), .B(n884), .Z(c[296]) );
  AND U1146 ( .A(b[0]), .B(a[42]), .Z(n888) );
  XNOR U1147 ( .A(n889), .B(sreg[297]), .Z(n887) );
  XOR U1148 ( .A(n888), .B(n887), .Z(c[297]) );
  AND U1149 ( .A(b[0]), .B(a[43]), .Z(n891) );
  XNOR U1150 ( .A(n892), .B(sreg[298]), .Z(n890) );
  XOR U1151 ( .A(n891), .B(n890), .Z(c[298]) );
  AND U1152 ( .A(b[0]), .B(a[44]), .Z(n894) );
  XNOR U1153 ( .A(n895), .B(sreg[299]), .Z(n893) );
  XOR U1154 ( .A(n894), .B(n893), .Z(c[299]) );
  AND U1155 ( .A(b[0]), .B(a[45]), .Z(n897) );
  XNOR U1156 ( .A(n898), .B(sreg[300]), .Z(n896) );
  XOR U1157 ( .A(n897), .B(n896), .Z(c[300]) );
  AND U1158 ( .A(b[0]), .B(a[46]), .Z(n900) );
  XNOR U1159 ( .A(n901), .B(sreg[301]), .Z(n899) );
  XOR U1160 ( .A(n900), .B(n899), .Z(c[301]) );
  AND U1161 ( .A(b[0]), .B(a[47]), .Z(n903) );
  XNOR U1162 ( .A(n904), .B(sreg[302]), .Z(n902) );
  XOR U1163 ( .A(n903), .B(n902), .Z(c[302]) );
  AND U1164 ( .A(b[0]), .B(a[48]), .Z(n906) );
  XNOR U1165 ( .A(n907), .B(sreg[303]), .Z(n905) );
  XOR U1166 ( .A(n906), .B(n905), .Z(c[303]) );
  AND U1167 ( .A(b[0]), .B(a[49]), .Z(n909) );
  XNOR U1168 ( .A(n910), .B(sreg[304]), .Z(n908) );
  XOR U1169 ( .A(n909), .B(n908), .Z(c[304]) );
  AND U1170 ( .A(b[0]), .B(a[50]), .Z(n912) );
  XNOR U1171 ( .A(n913), .B(sreg[305]), .Z(n911) );
  XOR U1172 ( .A(n912), .B(n911), .Z(c[305]) );
  AND U1173 ( .A(b[0]), .B(a[51]), .Z(n915) );
  XNOR U1174 ( .A(n916), .B(sreg[306]), .Z(n914) );
  XOR U1175 ( .A(n915), .B(n914), .Z(c[306]) );
  AND U1176 ( .A(b[0]), .B(a[52]), .Z(n918) );
  XNOR U1177 ( .A(n919), .B(sreg[307]), .Z(n917) );
  XOR U1178 ( .A(n918), .B(n917), .Z(c[307]) );
  AND U1179 ( .A(b[0]), .B(a[53]), .Z(n921) );
  XNOR U1180 ( .A(n922), .B(sreg[308]), .Z(n920) );
  XOR U1181 ( .A(n921), .B(n920), .Z(c[308]) );
  AND U1182 ( .A(b[0]), .B(a[54]), .Z(n924) );
  XNOR U1183 ( .A(n925), .B(sreg[309]), .Z(n923) );
  XOR U1184 ( .A(n924), .B(n923), .Z(c[309]) );
  AND U1185 ( .A(b[0]), .B(a[55]), .Z(n927) );
  XNOR U1186 ( .A(n928), .B(sreg[310]), .Z(n926) );
  XOR U1187 ( .A(n927), .B(n926), .Z(c[310]) );
  AND U1188 ( .A(b[0]), .B(a[56]), .Z(n930) );
  XNOR U1189 ( .A(n931), .B(sreg[311]), .Z(n929) );
  XOR U1190 ( .A(n930), .B(n929), .Z(c[311]) );
  AND U1191 ( .A(b[0]), .B(a[57]), .Z(n933) );
  XNOR U1192 ( .A(n934), .B(sreg[312]), .Z(n932) );
  XOR U1193 ( .A(n933), .B(n932), .Z(c[312]) );
  AND U1194 ( .A(b[0]), .B(a[58]), .Z(n936) );
  XNOR U1195 ( .A(n937), .B(sreg[313]), .Z(n935) );
  XOR U1196 ( .A(n936), .B(n935), .Z(c[313]) );
  AND U1197 ( .A(b[0]), .B(a[59]), .Z(n939) );
  XNOR U1198 ( .A(n940), .B(sreg[314]), .Z(n938) );
  XOR U1199 ( .A(n939), .B(n938), .Z(c[314]) );
  AND U1200 ( .A(b[0]), .B(a[60]), .Z(n942) );
  XNOR U1201 ( .A(n943), .B(sreg[315]), .Z(n941) );
  XOR U1202 ( .A(n942), .B(n941), .Z(c[315]) );
  AND U1203 ( .A(b[0]), .B(a[61]), .Z(n945) );
  XNOR U1204 ( .A(n946), .B(sreg[316]), .Z(n944) );
  XOR U1205 ( .A(n945), .B(n944), .Z(c[316]) );
  AND U1206 ( .A(b[0]), .B(a[62]), .Z(n948) );
  XNOR U1207 ( .A(n949), .B(sreg[317]), .Z(n947) );
  XOR U1208 ( .A(n948), .B(n947), .Z(c[317]) );
  AND U1209 ( .A(b[0]), .B(a[63]), .Z(n951) );
  XNOR U1210 ( .A(n952), .B(sreg[318]), .Z(n950) );
  XOR U1211 ( .A(n951), .B(n950), .Z(c[318]) );
  AND U1212 ( .A(b[0]), .B(a[64]), .Z(n954) );
  XNOR U1213 ( .A(n955), .B(sreg[319]), .Z(n953) );
  XOR U1214 ( .A(n954), .B(n953), .Z(c[319]) );
  AND U1215 ( .A(b[0]), .B(a[65]), .Z(n957) );
  XNOR U1216 ( .A(n958), .B(sreg[320]), .Z(n956) );
  XOR U1217 ( .A(n957), .B(n956), .Z(c[320]) );
  AND U1218 ( .A(b[0]), .B(a[66]), .Z(n960) );
  XNOR U1219 ( .A(n961), .B(sreg[321]), .Z(n959) );
  XOR U1220 ( .A(n960), .B(n959), .Z(c[321]) );
  AND U1221 ( .A(b[0]), .B(a[67]), .Z(n963) );
  XNOR U1222 ( .A(n964), .B(sreg[322]), .Z(n962) );
  XOR U1223 ( .A(n963), .B(n962), .Z(c[322]) );
  AND U1224 ( .A(b[0]), .B(a[68]), .Z(n966) );
  XNOR U1225 ( .A(n967), .B(sreg[323]), .Z(n965) );
  XOR U1226 ( .A(n966), .B(n965), .Z(c[323]) );
  AND U1227 ( .A(b[0]), .B(a[69]), .Z(n969) );
  XNOR U1228 ( .A(n970), .B(sreg[324]), .Z(n968) );
  XOR U1229 ( .A(n969), .B(n968), .Z(c[324]) );
  AND U1230 ( .A(b[0]), .B(a[70]), .Z(n972) );
  XNOR U1231 ( .A(n973), .B(sreg[325]), .Z(n971) );
  XOR U1232 ( .A(n972), .B(n971), .Z(c[325]) );
  AND U1233 ( .A(b[0]), .B(a[71]), .Z(n975) );
  XNOR U1234 ( .A(n976), .B(sreg[326]), .Z(n974) );
  XOR U1235 ( .A(n975), .B(n974), .Z(c[326]) );
  AND U1236 ( .A(b[0]), .B(a[72]), .Z(n978) );
  XNOR U1237 ( .A(n979), .B(sreg[327]), .Z(n977) );
  XOR U1238 ( .A(n978), .B(n977), .Z(c[327]) );
  AND U1239 ( .A(b[0]), .B(a[73]), .Z(n981) );
  XNOR U1240 ( .A(n982), .B(sreg[328]), .Z(n980) );
  XOR U1241 ( .A(n981), .B(n980), .Z(c[328]) );
  AND U1242 ( .A(b[0]), .B(a[74]), .Z(n984) );
  XNOR U1243 ( .A(n985), .B(sreg[329]), .Z(n983) );
  XOR U1244 ( .A(n984), .B(n983), .Z(c[329]) );
  AND U1245 ( .A(b[0]), .B(a[75]), .Z(n987) );
  XNOR U1246 ( .A(n988), .B(sreg[330]), .Z(n986) );
  XOR U1247 ( .A(n987), .B(n986), .Z(c[330]) );
  AND U1248 ( .A(b[0]), .B(a[76]), .Z(n990) );
  XNOR U1249 ( .A(n991), .B(sreg[331]), .Z(n989) );
  XOR U1250 ( .A(n990), .B(n989), .Z(c[331]) );
  AND U1251 ( .A(b[0]), .B(a[77]), .Z(n993) );
  XNOR U1252 ( .A(n994), .B(sreg[332]), .Z(n992) );
  XOR U1253 ( .A(n993), .B(n992), .Z(c[332]) );
  AND U1254 ( .A(b[0]), .B(a[78]), .Z(n996) );
  XNOR U1255 ( .A(n997), .B(sreg[333]), .Z(n995) );
  XOR U1256 ( .A(n996), .B(n995), .Z(c[333]) );
  AND U1257 ( .A(b[0]), .B(a[79]), .Z(n999) );
  XNOR U1258 ( .A(n1000), .B(sreg[334]), .Z(n998) );
  XOR U1259 ( .A(n999), .B(n998), .Z(c[334]) );
  AND U1260 ( .A(b[0]), .B(a[80]), .Z(n1002) );
  XNOR U1261 ( .A(n1003), .B(sreg[335]), .Z(n1001) );
  XOR U1262 ( .A(n1002), .B(n1001), .Z(c[335]) );
  AND U1263 ( .A(b[0]), .B(a[81]), .Z(n1005) );
  XNOR U1264 ( .A(n1006), .B(sreg[336]), .Z(n1004) );
  XOR U1265 ( .A(n1005), .B(n1004), .Z(c[336]) );
  AND U1266 ( .A(b[0]), .B(a[82]), .Z(n1008) );
  XNOR U1267 ( .A(n1009), .B(sreg[337]), .Z(n1007) );
  XOR U1268 ( .A(n1008), .B(n1007), .Z(c[337]) );
  AND U1269 ( .A(b[0]), .B(a[83]), .Z(n1011) );
  XNOR U1270 ( .A(n1012), .B(sreg[338]), .Z(n1010) );
  XOR U1271 ( .A(n1011), .B(n1010), .Z(c[338]) );
  AND U1272 ( .A(b[0]), .B(a[84]), .Z(n1014) );
  XNOR U1273 ( .A(n1015), .B(sreg[339]), .Z(n1013) );
  XOR U1274 ( .A(n1014), .B(n1013), .Z(c[339]) );
  AND U1275 ( .A(b[0]), .B(a[85]), .Z(n1017) );
  XNOR U1276 ( .A(n1018), .B(sreg[340]), .Z(n1016) );
  XOR U1277 ( .A(n1017), .B(n1016), .Z(c[340]) );
  AND U1278 ( .A(b[0]), .B(a[86]), .Z(n1020) );
  XNOR U1279 ( .A(n1021), .B(sreg[341]), .Z(n1019) );
  XOR U1280 ( .A(n1020), .B(n1019), .Z(c[341]) );
  AND U1281 ( .A(b[0]), .B(a[87]), .Z(n1023) );
  XNOR U1282 ( .A(n1024), .B(sreg[342]), .Z(n1022) );
  XOR U1283 ( .A(n1023), .B(n1022), .Z(c[342]) );
  AND U1284 ( .A(b[0]), .B(a[88]), .Z(n1026) );
  XNOR U1285 ( .A(n1027), .B(sreg[343]), .Z(n1025) );
  XOR U1286 ( .A(n1026), .B(n1025), .Z(c[343]) );
  AND U1287 ( .A(b[0]), .B(a[89]), .Z(n1029) );
  XNOR U1288 ( .A(n1030), .B(sreg[344]), .Z(n1028) );
  XOR U1289 ( .A(n1029), .B(n1028), .Z(c[344]) );
  AND U1290 ( .A(b[0]), .B(a[90]), .Z(n1032) );
  XNOR U1291 ( .A(n1033), .B(sreg[345]), .Z(n1031) );
  XOR U1292 ( .A(n1032), .B(n1031), .Z(c[345]) );
  AND U1293 ( .A(b[0]), .B(a[91]), .Z(n1035) );
  XNOR U1294 ( .A(n1036), .B(sreg[346]), .Z(n1034) );
  XOR U1295 ( .A(n1035), .B(n1034), .Z(c[346]) );
  AND U1296 ( .A(b[0]), .B(a[92]), .Z(n1038) );
  XNOR U1297 ( .A(n1039), .B(sreg[347]), .Z(n1037) );
  XOR U1298 ( .A(n1038), .B(n1037), .Z(c[347]) );
  AND U1299 ( .A(b[0]), .B(a[93]), .Z(n1041) );
  XNOR U1300 ( .A(n1042), .B(sreg[348]), .Z(n1040) );
  XOR U1301 ( .A(n1041), .B(n1040), .Z(c[348]) );
  AND U1302 ( .A(b[0]), .B(a[94]), .Z(n1044) );
  XNOR U1303 ( .A(n1045), .B(sreg[349]), .Z(n1043) );
  XOR U1304 ( .A(n1044), .B(n1043), .Z(c[349]) );
  AND U1305 ( .A(b[0]), .B(a[95]), .Z(n1047) );
  XNOR U1306 ( .A(n1048), .B(sreg[350]), .Z(n1046) );
  XOR U1307 ( .A(n1047), .B(n1046), .Z(c[350]) );
  AND U1308 ( .A(b[0]), .B(a[96]), .Z(n1050) );
  XNOR U1309 ( .A(n1051), .B(sreg[351]), .Z(n1049) );
  XOR U1310 ( .A(n1050), .B(n1049), .Z(c[351]) );
  AND U1311 ( .A(b[0]), .B(a[97]), .Z(n1053) );
  XNOR U1312 ( .A(n1054), .B(sreg[352]), .Z(n1052) );
  XOR U1313 ( .A(n1053), .B(n1052), .Z(c[352]) );
  AND U1314 ( .A(b[0]), .B(a[98]), .Z(n1056) );
  XNOR U1315 ( .A(n1057), .B(sreg[353]), .Z(n1055) );
  XOR U1316 ( .A(n1056), .B(n1055), .Z(c[353]) );
  AND U1317 ( .A(b[0]), .B(a[99]), .Z(n1059) );
  XNOR U1318 ( .A(n1060), .B(sreg[354]), .Z(n1058) );
  XOR U1319 ( .A(n1059), .B(n1058), .Z(c[354]) );
  AND U1320 ( .A(b[0]), .B(a[100]), .Z(n1062) );
  XNOR U1321 ( .A(n1063), .B(sreg[355]), .Z(n1061) );
  XOR U1322 ( .A(n1062), .B(n1061), .Z(c[355]) );
  AND U1323 ( .A(b[0]), .B(a[101]), .Z(n1065) );
  XNOR U1324 ( .A(n1066), .B(sreg[356]), .Z(n1064) );
  XOR U1325 ( .A(n1065), .B(n1064), .Z(c[356]) );
  AND U1326 ( .A(b[0]), .B(a[102]), .Z(n1068) );
  XNOR U1327 ( .A(n1069), .B(sreg[357]), .Z(n1067) );
  XOR U1328 ( .A(n1068), .B(n1067), .Z(c[357]) );
  AND U1329 ( .A(b[0]), .B(a[103]), .Z(n1071) );
  XNOR U1330 ( .A(n1072), .B(sreg[358]), .Z(n1070) );
  XOR U1331 ( .A(n1071), .B(n1070), .Z(c[358]) );
  AND U1332 ( .A(b[0]), .B(a[104]), .Z(n1074) );
  XNOR U1333 ( .A(n1075), .B(sreg[359]), .Z(n1073) );
  XOR U1334 ( .A(n1074), .B(n1073), .Z(c[359]) );
  AND U1335 ( .A(b[0]), .B(a[105]), .Z(n1077) );
  XNOR U1336 ( .A(n1078), .B(sreg[360]), .Z(n1076) );
  XOR U1337 ( .A(n1077), .B(n1076), .Z(c[360]) );
  AND U1338 ( .A(b[0]), .B(a[106]), .Z(n1080) );
  XNOR U1339 ( .A(n1081), .B(sreg[361]), .Z(n1079) );
  XOR U1340 ( .A(n1080), .B(n1079), .Z(c[361]) );
  AND U1341 ( .A(b[0]), .B(a[107]), .Z(n1083) );
  XNOR U1342 ( .A(n1084), .B(sreg[362]), .Z(n1082) );
  XOR U1343 ( .A(n1083), .B(n1082), .Z(c[362]) );
  AND U1344 ( .A(b[0]), .B(a[108]), .Z(n1086) );
  XNOR U1345 ( .A(n1087), .B(sreg[363]), .Z(n1085) );
  XOR U1346 ( .A(n1086), .B(n1085), .Z(c[363]) );
  AND U1347 ( .A(b[0]), .B(a[109]), .Z(n1089) );
  XNOR U1348 ( .A(n1090), .B(sreg[364]), .Z(n1088) );
  XOR U1349 ( .A(n1089), .B(n1088), .Z(c[364]) );
  AND U1350 ( .A(b[0]), .B(a[110]), .Z(n1092) );
  XNOR U1351 ( .A(n1093), .B(sreg[365]), .Z(n1091) );
  XOR U1352 ( .A(n1092), .B(n1091), .Z(c[365]) );
  AND U1353 ( .A(b[0]), .B(a[111]), .Z(n1095) );
  XNOR U1354 ( .A(n1096), .B(sreg[366]), .Z(n1094) );
  XOR U1355 ( .A(n1095), .B(n1094), .Z(c[366]) );
  AND U1356 ( .A(b[0]), .B(a[112]), .Z(n1098) );
  XNOR U1357 ( .A(n1099), .B(sreg[367]), .Z(n1097) );
  XOR U1358 ( .A(n1098), .B(n1097), .Z(c[367]) );
  AND U1359 ( .A(b[0]), .B(a[113]), .Z(n1101) );
  XNOR U1360 ( .A(n1102), .B(sreg[368]), .Z(n1100) );
  XOR U1361 ( .A(n1101), .B(n1100), .Z(c[368]) );
  AND U1362 ( .A(b[0]), .B(a[114]), .Z(n1104) );
  XNOR U1363 ( .A(n1105), .B(sreg[369]), .Z(n1103) );
  XOR U1364 ( .A(n1104), .B(n1103), .Z(c[369]) );
  AND U1365 ( .A(b[0]), .B(a[115]), .Z(n1107) );
  XNOR U1366 ( .A(n1108), .B(sreg[370]), .Z(n1106) );
  XOR U1367 ( .A(n1107), .B(n1106), .Z(c[370]) );
  AND U1368 ( .A(b[0]), .B(a[116]), .Z(n1110) );
  XNOR U1369 ( .A(n1111), .B(sreg[371]), .Z(n1109) );
  XOR U1370 ( .A(n1110), .B(n1109), .Z(c[371]) );
  AND U1371 ( .A(b[0]), .B(a[117]), .Z(n1113) );
  XNOR U1372 ( .A(n1114), .B(sreg[372]), .Z(n1112) );
  XOR U1373 ( .A(n1113), .B(n1112), .Z(c[372]) );
  AND U1374 ( .A(b[0]), .B(a[118]), .Z(n1116) );
  XNOR U1375 ( .A(n1117), .B(sreg[373]), .Z(n1115) );
  XOR U1376 ( .A(n1116), .B(n1115), .Z(c[373]) );
  AND U1377 ( .A(b[0]), .B(a[119]), .Z(n1119) );
  XNOR U1378 ( .A(n1120), .B(sreg[374]), .Z(n1118) );
  XOR U1379 ( .A(n1119), .B(n1118), .Z(c[374]) );
  AND U1380 ( .A(b[0]), .B(a[120]), .Z(n1122) );
  XNOR U1381 ( .A(n1123), .B(sreg[375]), .Z(n1121) );
  XOR U1382 ( .A(n1122), .B(n1121), .Z(c[375]) );
  AND U1383 ( .A(b[0]), .B(a[121]), .Z(n1125) );
  XNOR U1384 ( .A(n1126), .B(sreg[376]), .Z(n1124) );
  XOR U1385 ( .A(n1125), .B(n1124), .Z(c[376]) );
  AND U1386 ( .A(b[0]), .B(a[122]), .Z(n1128) );
  XNOR U1387 ( .A(n1129), .B(sreg[377]), .Z(n1127) );
  XOR U1388 ( .A(n1128), .B(n1127), .Z(c[377]) );
  AND U1389 ( .A(b[0]), .B(a[123]), .Z(n1131) );
  XNOR U1390 ( .A(n1132), .B(sreg[378]), .Z(n1130) );
  XOR U1391 ( .A(n1131), .B(n1130), .Z(c[378]) );
  AND U1392 ( .A(b[0]), .B(a[124]), .Z(n1134) );
  XNOR U1393 ( .A(n1135), .B(sreg[379]), .Z(n1133) );
  XOR U1394 ( .A(n1134), .B(n1133), .Z(c[379]) );
  AND U1395 ( .A(b[0]), .B(a[125]), .Z(n1137) );
  XNOR U1396 ( .A(n1138), .B(sreg[380]), .Z(n1136) );
  XOR U1397 ( .A(n1137), .B(n1136), .Z(c[380]) );
  AND U1398 ( .A(b[0]), .B(a[126]), .Z(n1140) );
  XNOR U1399 ( .A(n1141), .B(sreg[381]), .Z(n1139) );
  XOR U1400 ( .A(n1140), .B(n1139), .Z(c[381]) );
  AND U1401 ( .A(b[0]), .B(a[127]), .Z(n1143) );
  XNOR U1402 ( .A(n1144), .B(sreg[382]), .Z(n1142) );
  XOR U1403 ( .A(n1143), .B(n1142), .Z(c[382]) );
  AND U1404 ( .A(b[0]), .B(a[128]), .Z(n1146) );
  XNOR U1405 ( .A(n1147), .B(sreg[383]), .Z(n1145) );
  XOR U1406 ( .A(n1146), .B(n1145), .Z(c[383]) );
  AND U1407 ( .A(b[0]), .B(a[129]), .Z(n1149) );
  XNOR U1408 ( .A(n1150), .B(sreg[384]), .Z(n1148) );
  XOR U1409 ( .A(n1149), .B(n1148), .Z(c[384]) );
  AND U1410 ( .A(b[0]), .B(a[130]), .Z(n1152) );
  XNOR U1411 ( .A(n1153), .B(sreg[385]), .Z(n1151) );
  XOR U1412 ( .A(n1152), .B(n1151), .Z(c[385]) );
  AND U1413 ( .A(b[0]), .B(a[131]), .Z(n1155) );
  XNOR U1414 ( .A(n1156), .B(sreg[386]), .Z(n1154) );
  XOR U1415 ( .A(n1155), .B(n1154), .Z(c[386]) );
  AND U1416 ( .A(b[0]), .B(a[132]), .Z(n1158) );
  XNOR U1417 ( .A(n1159), .B(sreg[387]), .Z(n1157) );
  XOR U1418 ( .A(n1158), .B(n1157), .Z(c[387]) );
  AND U1419 ( .A(b[0]), .B(a[133]), .Z(n1161) );
  XNOR U1420 ( .A(n1162), .B(sreg[388]), .Z(n1160) );
  XOR U1421 ( .A(n1161), .B(n1160), .Z(c[388]) );
  AND U1422 ( .A(b[0]), .B(a[134]), .Z(n1164) );
  XNOR U1423 ( .A(n1165), .B(sreg[389]), .Z(n1163) );
  XOR U1424 ( .A(n1164), .B(n1163), .Z(c[389]) );
  AND U1425 ( .A(b[0]), .B(a[135]), .Z(n1167) );
  XNOR U1426 ( .A(n1168), .B(sreg[390]), .Z(n1166) );
  XOR U1427 ( .A(n1167), .B(n1166), .Z(c[390]) );
  AND U1428 ( .A(b[0]), .B(a[136]), .Z(n1170) );
  XNOR U1429 ( .A(n1171), .B(sreg[391]), .Z(n1169) );
  XOR U1430 ( .A(n1170), .B(n1169), .Z(c[391]) );
  AND U1431 ( .A(b[0]), .B(a[137]), .Z(n1173) );
  XNOR U1432 ( .A(n1174), .B(sreg[392]), .Z(n1172) );
  XOR U1433 ( .A(n1173), .B(n1172), .Z(c[392]) );
  AND U1434 ( .A(b[0]), .B(a[138]), .Z(n1176) );
  XNOR U1435 ( .A(n1177), .B(sreg[393]), .Z(n1175) );
  XOR U1436 ( .A(n1176), .B(n1175), .Z(c[393]) );
  AND U1437 ( .A(b[0]), .B(a[139]), .Z(n1179) );
  XNOR U1438 ( .A(n1180), .B(sreg[394]), .Z(n1178) );
  XOR U1439 ( .A(n1179), .B(n1178), .Z(c[394]) );
  AND U1440 ( .A(b[0]), .B(a[140]), .Z(n1182) );
  XNOR U1441 ( .A(n1183), .B(sreg[395]), .Z(n1181) );
  XOR U1442 ( .A(n1182), .B(n1181), .Z(c[395]) );
  AND U1443 ( .A(b[0]), .B(a[141]), .Z(n1185) );
  XNOR U1444 ( .A(n1186), .B(sreg[396]), .Z(n1184) );
  XOR U1445 ( .A(n1185), .B(n1184), .Z(c[396]) );
  AND U1446 ( .A(b[0]), .B(a[142]), .Z(n1188) );
  XNOR U1447 ( .A(n1189), .B(sreg[397]), .Z(n1187) );
  XOR U1448 ( .A(n1188), .B(n1187), .Z(c[397]) );
  AND U1449 ( .A(b[0]), .B(a[143]), .Z(n1191) );
  XNOR U1450 ( .A(n1192), .B(sreg[398]), .Z(n1190) );
  XOR U1451 ( .A(n1191), .B(n1190), .Z(c[398]) );
  AND U1452 ( .A(b[0]), .B(a[144]), .Z(n1194) );
  XNOR U1453 ( .A(n1195), .B(sreg[399]), .Z(n1193) );
  XOR U1454 ( .A(n1194), .B(n1193), .Z(c[399]) );
  AND U1455 ( .A(b[0]), .B(a[145]), .Z(n1197) );
  XNOR U1456 ( .A(n1198), .B(sreg[400]), .Z(n1196) );
  XOR U1457 ( .A(n1197), .B(n1196), .Z(c[400]) );
  AND U1458 ( .A(b[0]), .B(a[146]), .Z(n1200) );
  XNOR U1459 ( .A(n1201), .B(sreg[401]), .Z(n1199) );
  XOR U1460 ( .A(n1200), .B(n1199), .Z(c[401]) );
  AND U1461 ( .A(b[0]), .B(a[147]), .Z(n1203) );
  XNOR U1462 ( .A(n1204), .B(sreg[402]), .Z(n1202) );
  XOR U1463 ( .A(n1203), .B(n1202), .Z(c[402]) );
  AND U1464 ( .A(b[0]), .B(a[148]), .Z(n1206) );
  XNOR U1465 ( .A(n1207), .B(sreg[403]), .Z(n1205) );
  XOR U1466 ( .A(n1206), .B(n1205), .Z(c[403]) );
  AND U1467 ( .A(b[0]), .B(a[149]), .Z(n1209) );
  XNOR U1468 ( .A(n1210), .B(sreg[404]), .Z(n1208) );
  XOR U1469 ( .A(n1209), .B(n1208), .Z(c[404]) );
  AND U1470 ( .A(b[0]), .B(a[150]), .Z(n1212) );
  XNOR U1471 ( .A(n1213), .B(sreg[405]), .Z(n1211) );
  XOR U1472 ( .A(n1212), .B(n1211), .Z(c[405]) );
  AND U1473 ( .A(b[0]), .B(a[151]), .Z(n1215) );
  XNOR U1474 ( .A(n1216), .B(sreg[406]), .Z(n1214) );
  XOR U1475 ( .A(n1215), .B(n1214), .Z(c[406]) );
  AND U1476 ( .A(b[0]), .B(a[152]), .Z(n1218) );
  XNOR U1477 ( .A(n1219), .B(sreg[407]), .Z(n1217) );
  XOR U1478 ( .A(n1218), .B(n1217), .Z(c[407]) );
  AND U1479 ( .A(b[0]), .B(a[153]), .Z(n1221) );
  XNOR U1480 ( .A(n1222), .B(sreg[408]), .Z(n1220) );
  XOR U1481 ( .A(n1221), .B(n1220), .Z(c[408]) );
  AND U1482 ( .A(b[0]), .B(a[154]), .Z(n1224) );
  XNOR U1483 ( .A(n1225), .B(sreg[409]), .Z(n1223) );
  XOR U1484 ( .A(n1224), .B(n1223), .Z(c[409]) );
  AND U1485 ( .A(b[0]), .B(a[155]), .Z(n1227) );
  XNOR U1486 ( .A(n1228), .B(sreg[410]), .Z(n1226) );
  XOR U1487 ( .A(n1227), .B(n1226), .Z(c[410]) );
  AND U1488 ( .A(b[0]), .B(a[156]), .Z(n1230) );
  XNOR U1489 ( .A(n1231), .B(sreg[411]), .Z(n1229) );
  XOR U1490 ( .A(n1230), .B(n1229), .Z(c[411]) );
  AND U1491 ( .A(b[0]), .B(a[157]), .Z(n1233) );
  XNOR U1492 ( .A(n1234), .B(sreg[412]), .Z(n1232) );
  XOR U1493 ( .A(n1233), .B(n1232), .Z(c[412]) );
  AND U1494 ( .A(b[0]), .B(a[158]), .Z(n1236) );
  XNOR U1495 ( .A(n1237), .B(sreg[413]), .Z(n1235) );
  XOR U1496 ( .A(n1236), .B(n1235), .Z(c[413]) );
  AND U1497 ( .A(b[0]), .B(a[159]), .Z(n1239) );
  XNOR U1498 ( .A(n1240), .B(sreg[414]), .Z(n1238) );
  XOR U1499 ( .A(n1239), .B(n1238), .Z(c[414]) );
  AND U1500 ( .A(b[0]), .B(a[160]), .Z(n1242) );
  XNOR U1501 ( .A(n1243), .B(sreg[415]), .Z(n1241) );
  XOR U1502 ( .A(n1242), .B(n1241), .Z(c[415]) );
  AND U1503 ( .A(b[0]), .B(a[161]), .Z(n1245) );
  XNOR U1504 ( .A(n1246), .B(sreg[416]), .Z(n1244) );
  XOR U1505 ( .A(n1245), .B(n1244), .Z(c[416]) );
  AND U1506 ( .A(b[0]), .B(a[162]), .Z(n1248) );
  XNOR U1507 ( .A(n1249), .B(sreg[417]), .Z(n1247) );
  XOR U1508 ( .A(n1248), .B(n1247), .Z(c[417]) );
  AND U1509 ( .A(b[0]), .B(a[163]), .Z(n1251) );
  XNOR U1510 ( .A(n1252), .B(sreg[418]), .Z(n1250) );
  XOR U1511 ( .A(n1251), .B(n1250), .Z(c[418]) );
  AND U1512 ( .A(b[0]), .B(a[164]), .Z(n1254) );
  XNOR U1513 ( .A(n1255), .B(sreg[419]), .Z(n1253) );
  XOR U1514 ( .A(n1254), .B(n1253), .Z(c[419]) );
  AND U1515 ( .A(b[0]), .B(a[165]), .Z(n1257) );
  XNOR U1516 ( .A(n1258), .B(sreg[420]), .Z(n1256) );
  XOR U1517 ( .A(n1257), .B(n1256), .Z(c[420]) );
  AND U1518 ( .A(b[0]), .B(a[166]), .Z(n1260) );
  XNOR U1519 ( .A(n1261), .B(sreg[421]), .Z(n1259) );
  XOR U1520 ( .A(n1260), .B(n1259), .Z(c[421]) );
  AND U1521 ( .A(b[0]), .B(a[167]), .Z(n1263) );
  XNOR U1522 ( .A(n1264), .B(sreg[422]), .Z(n1262) );
  XOR U1523 ( .A(n1263), .B(n1262), .Z(c[422]) );
  AND U1524 ( .A(b[0]), .B(a[168]), .Z(n1266) );
  XNOR U1525 ( .A(n1267), .B(sreg[423]), .Z(n1265) );
  XOR U1526 ( .A(n1266), .B(n1265), .Z(c[423]) );
  AND U1527 ( .A(b[0]), .B(a[169]), .Z(n1269) );
  XNOR U1528 ( .A(n1270), .B(sreg[424]), .Z(n1268) );
  XOR U1529 ( .A(n1269), .B(n1268), .Z(c[424]) );
  AND U1530 ( .A(b[0]), .B(a[170]), .Z(n1272) );
  XNOR U1531 ( .A(n1273), .B(sreg[425]), .Z(n1271) );
  XOR U1532 ( .A(n1272), .B(n1271), .Z(c[425]) );
  AND U1533 ( .A(b[0]), .B(a[171]), .Z(n1275) );
  XNOR U1534 ( .A(n1276), .B(sreg[426]), .Z(n1274) );
  XOR U1535 ( .A(n1275), .B(n1274), .Z(c[426]) );
  AND U1536 ( .A(b[0]), .B(a[172]), .Z(n1278) );
  XNOR U1537 ( .A(n1279), .B(sreg[427]), .Z(n1277) );
  XOR U1538 ( .A(n1278), .B(n1277), .Z(c[427]) );
  AND U1539 ( .A(b[0]), .B(a[173]), .Z(n1281) );
  XNOR U1540 ( .A(n1282), .B(sreg[428]), .Z(n1280) );
  XOR U1541 ( .A(n1281), .B(n1280), .Z(c[428]) );
  AND U1542 ( .A(b[0]), .B(a[174]), .Z(n1284) );
  XNOR U1543 ( .A(n1285), .B(sreg[429]), .Z(n1283) );
  XOR U1544 ( .A(n1284), .B(n1283), .Z(c[429]) );
  AND U1545 ( .A(b[0]), .B(a[175]), .Z(n1287) );
  XNOR U1546 ( .A(n1288), .B(sreg[430]), .Z(n1286) );
  XOR U1547 ( .A(n1287), .B(n1286), .Z(c[430]) );
  AND U1548 ( .A(b[0]), .B(a[176]), .Z(n1290) );
  XNOR U1549 ( .A(n1291), .B(sreg[431]), .Z(n1289) );
  XOR U1550 ( .A(n1290), .B(n1289), .Z(c[431]) );
  AND U1551 ( .A(b[0]), .B(a[177]), .Z(n1293) );
  XNOR U1552 ( .A(n1294), .B(sreg[432]), .Z(n1292) );
  XOR U1553 ( .A(n1293), .B(n1292), .Z(c[432]) );
  AND U1554 ( .A(b[0]), .B(a[178]), .Z(n1296) );
  XNOR U1555 ( .A(n1297), .B(sreg[433]), .Z(n1295) );
  XOR U1556 ( .A(n1296), .B(n1295), .Z(c[433]) );
  AND U1557 ( .A(b[0]), .B(a[179]), .Z(n1299) );
  XNOR U1558 ( .A(n1300), .B(sreg[434]), .Z(n1298) );
  XOR U1559 ( .A(n1299), .B(n1298), .Z(c[434]) );
  AND U1560 ( .A(b[0]), .B(a[180]), .Z(n1302) );
  XNOR U1561 ( .A(n1303), .B(sreg[435]), .Z(n1301) );
  XOR U1562 ( .A(n1302), .B(n1301), .Z(c[435]) );
  AND U1563 ( .A(b[0]), .B(a[181]), .Z(n1305) );
  XNOR U1564 ( .A(n1306), .B(sreg[436]), .Z(n1304) );
  XOR U1565 ( .A(n1305), .B(n1304), .Z(c[436]) );
  AND U1566 ( .A(b[0]), .B(a[182]), .Z(n1308) );
  XNOR U1567 ( .A(n1309), .B(sreg[437]), .Z(n1307) );
  XOR U1568 ( .A(n1308), .B(n1307), .Z(c[437]) );
  AND U1569 ( .A(b[0]), .B(a[183]), .Z(n1311) );
  XNOR U1570 ( .A(n1312), .B(sreg[438]), .Z(n1310) );
  XOR U1571 ( .A(n1311), .B(n1310), .Z(c[438]) );
  AND U1572 ( .A(b[0]), .B(a[184]), .Z(n1314) );
  XNOR U1573 ( .A(n1315), .B(sreg[439]), .Z(n1313) );
  XOR U1574 ( .A(n1314), .B(n1313), .Z(c[439]) );
  AND U1575 ( .A(b[0]), .B(a[185]), .Z(n1317) );
  XNOR U1576 ( .A(n1318), .B(sreg[440]), .Z(n1316) );
  XOR U1577 ( .A(n1317), .B(n1316), .Z(c[440]) );
  AND U1578 ( .A(b[0]), .B(a[186]), .Z(n1320) );
  XNOR U1579 ( .A(n1321), .B(sreg[441]), .Z(n1319) );
  XOR U1580 ( .A(n1320), .B(n1319), .Z(c[441]) );
  AND U1581 ( .A(b[0]), .B(a[187]), .Z(n1323) );
  XNOR U1582 ( .A(n1324), .B(sreg[442]), .Z(n1322) );
  XOR U1583 ( .A(n1323), .B(n1322), .Z(c[442]) );
  AND U1584 ( .A(b[0]), .B(a[188]), .Z(n1326) );
  XNOR U1585 ( .A(n1327), .B(sreg[443]), .Z(n1325) );
  XOR U1586 ( .A(n1326), .B(n1325), .Z(c[443]) );
  AND U1587 ( .A(b[0]), .B(a[189]), .Z(n1329) );
  XNOR U1588 ( .A(n1330), .B(sreg[444]), .Z(n1328) );
  XOR U1589 ( .A(n1329), .B(n1328), .Z(c[444]) );
  AND U1590 ( .A(b[0]), .B(a[190]), .Z(n1332) );
  XNOR U1591 ( .A(n1333), .B(sreg[445]), .Z(n1331) );
  XOR U1592 ( .A(n1332), .B(n1331), .Z(c[445]) );
  AND U1593 ( .A(b[0]), .B(a[191]), .Z(n1335) );
  XNOR U1594 ( .A(n1336), .B(sreg[446]), .Z(n1334) );
  XOR U1595 ( .A(n1335), .B(n1334), .Z(c[446]) );
  AND U1596 ( .A(b[0]), .B(a[192]), .Z(n1338) );
  XNOR U1597 ( .A(n1339), .B(sreg[447]), .Z(n1337) );
  XOR U1598 ( .A(n1338), .B(n1337), .Z(c[447]) );
  AND U1599 ( .A(b[0]), .B(a[193]), .Z(n1341) );
  XNOR U1600 ( .A(n1342), .B(sreg[448]), .Z(n1340) );
  XOR U1601 ( .A(n1341), .B(n1340), .Z(c[448]) );
  AND U1602 ( .A(b[0]), .B(a[194]), .Z(n1344) );
  XNOR U1603 ( .A(n1345), .B(sreg[449]), .Z(n1343) );
  XOR U1604 ( .A(n1344), .B(n1343), .Z(c[449]) );
  AND U1605 ( .A(b[0]), .B(a[195]), .Z(n1347) );
  XNOR U1606 ( .A(n1348), .B(sreg[450]), .Z(n1346) );
  XOR U1607 ( .A(n1347), .B(n1346), .Z(c[450]) );
  AND U1608 ( .A(b[0]), .B(a[196]), .Z(n1350) );
  XNOR U1609 ( .A(n1351), .B(sreg[451]), .Z(n1349) );
  XOR U1610 ( .A(n1350), .B(n1349), .Z(c[451]) );
  AND U1611 ( .A(b[0]), .B(a[197]), .Z(n1353) );
  XNOR U1612 ( .A(n1354), .B(sreg[452]), .Z(n1352) );
  XOR U1613 ( .A(n1353), .B(n1352), .Z(c[452]) );
  AND U1614 ( .A(b[0]), .B(a[198]), .Z(n1356) );
  XNOR U1615 ( .A(n1357), .B(sreg[453]), .Z(n1355) );
  XOR U1616 ( .A(n1356), .B(n1355), .Z(c[453]) );
  AND U1617 ( .A(b[0]), .B(a[199]), .Z(n1359) );
  XNOR U1618 ( .A(n1360), .B(sreg[454]), .Z(n1358) );
  XOR U1619 ( .A(n1359), .B(n1358), .Z(c[454]) );
  AND U1620 ( .A(b[0]), .B(a[200]), .Z(n1362) );
  XNOR U1621 ( .A(n1363), .B(sreg[455]), .Z(n1361) );
  XOR U1622 ( .A(n1362), .B(n1361), .Z(c[455]) );
  AND U1623 ( .A(b[0]), .B(a[201]), .Z(n1365) );
  XNOR U1624 ( .A(n1366), .B(sreg[456]), .Z(n1364) );
  XOR U1625 ( .A(n1365), .B(n1364), .Z(c[456]) );
  AND U1626 ( .A(b[0]), .B(a[202]), .Z(n1368) );
  XNOR U1627 ( .A(n1369), .B(sreg[457]), .Z(n1367) );
  XOR U1628 ( .A(n1368), .B(n1367), .Z(c[457]) );
  AND U1629 ( .A(b[0]), .B(a[203]), .Z(n1371) );
  XNOR U1630 ( .A(n1372), .B(sreg[458]), .Z(n1370) );
  XOR U1631 ( .A(n1371), .B(n1370), .Z(c[458]) );
  AND U1632 ( .A(b[0]), .B(a[204]), .Z(n1374) );
  XNOR U1633 ( .A(n1375), .B(sreg[459]), .Z(n1373) );
  XOR U1634 ( .A(n1374), .B(n1373), .Z(c[459]) );
  AND U1635 ( .A(b[0]), .B(a[205]), .Z(n1377) );
  XNOR U1636 ( .A(n1378), .B(sreg[460]), .Z(n1376) );
  XOR U1637 ( .A(n1377), .B(n1376), .Z(c[460]) );
  AND U1638 ( .A(b[0]), .B(a[206]), .Z(n1380) );
  XNOR U1639 ( .A(n1381), .B(sreg[461]), .Z(n1379) );
  XOR U1640 ( .A(n1380), .B(n1379), .Z(c[461]) );
  AND U1641 ( .A(b[0]), .B(a[207]), .Z(n1383) );
  XNOR U1642 ( .A(n1384), .B(sreg[462]), .Z(n1382) );
  XOR U1643 ( .A(n1383), .B(n1382), .Z(c[462]) );
  AND U1644 ( .A(b[0]), .B(a[208]), .Z(n1386) );
  XNOR U1645 ( .A(n1387), .B(sreg[463]), .Z(n1385) );
  XOR U1646 ( .A(n1386), .B(n1385), .Z(c[463]) );
  AND U1647 ( .A(b[0]), .B(a[209]), .Z(n1389) );
  XNOR U1648 ( .A(n1390), .B(sreg[464]), .Z(n1388) );
  XOR U1649 ( .A(n1389), .B(n1388), .Z(c[464]) );
  AND U1650 ( .A(b[0]), .B(a[210]), .Z(n1392) );
  XNOR U1651 ( .A(n1393), .B(sreg[465]), .Z(n1391) );
  XOR U1652 ( .A(n1392), .B(n1391), .Z(c[465]) );
  AND U1653 ( .A(b[0]), .B(a[211]), .Z(n1395) );
  XNOR U1654 ( .A(n1396), .B(sreg[466]), .Z(n1394) );
  XOR U1655 ( .A(n1395), .B(n1394), .Z(c[466]) );
  AND U1656 ( .A(b[0]), .B(a[212]), .Z(n1398) );
  XNOR U1657 ( .A(n1399), .B(sreg[467]), .Z(n1397) );
  XOR U1658 ( .A(n1398), .B(n1397), .Z(c[467]) );
  AND U1659 ( .A(b[0]), .B(a[213]), .Z(n1401) );
  XNOR U1660 ( .A(n1402), .B(sreg[468]), .Z(n1400) );
  XOR U1661 ( .A(n1401), .B(n1400), .Z(c[468]) );
  AND U1662 ( .A(b[0]), .B(a[214]), .Z(n1404) );
  XNOR U1663 ( .A(n1405), .B(sreg[469]), .Z(n1403) );
  XOR U1664 ( .A(n1404), .B(n1403), .Z(c[469]) );
  AND U1665 ( .A(b[0]), .B(a[215]), .Z(n1407) );
  XNOR U1666 ( .A(n1408), .B(sreg[470]), .Z(n1406) );
  XOR U1667 ( .A(n1407), .B(n1406), .Z(c[470]) );
  AND U1668 ( .A(b[0]), .B(a[216]), .Z(n1410) );
  XNOR U1669 ( .A(n1411), .B(sreg[471]), .Z(n1409) );
  XOR U1670 ( .A(n1410), .B(n1409), .Z(c[471]) );
  AND U1671 ( .A(b[0]), .B(a[217]), .Z(n1413) );
  XNOR U1672 ( .A(n1414), .B(sreg[472]), .Z(n1412) );
  XOR U1673 ( .A(n1413), .B(n1412), .Z(c[472]) );
  AND U1674 ( .A(b[0]), .B(a[218]), .Z(n1416) );
  XNOR U1675 ( .A(n1417), .B(sreg[473]), .Z(n1415) );
  XOR U1676 ( .A(n1416), .B(n1415), .Z(c[473]) );
  AND U1677 ( .A(b[0]), .B(a[219]), .Z(n1419) );
  XNOR U1678 ( .A(n1420), .B(sreg[474]), .Z(n1418) );
  XOR U1679 ( .A(n1419), .B(n1418), .Z(c[474]) );
  AND U1680 ( .A(b[0]), .B(a[220]), .Z(n1422) );
  XNOR U1681 ( .A(n1423), .B(sreg[475]), .Z(n1421) );
  XOR U1682 ( .A(n1422), .B(n1421), .Z(c[475]) );
  AND U1683 ( .A(b[0]), .B(a[221]), .Z(n1425) );
  XNOR U1684 ( .A(n1426), .B(sreg[476]), .Z(n1424) );
  XOR U1685 ( .A(n1425), .B(n1424), .Z(c[476]) );
  AND U1686 ( .A(b[0]), .B(a[222]), .Z(n1428) );
  XNOR U1687 ( .A(n1429), .B(sreg[477]), .Z(n1427) );
  XOR U1688 ( .A(n1428), .B(n1427), .Z(c[477]) );
  AND U1689 ( .A(b[0]), .B(a[223]), .Z(n1431) );
  XNOR U1690 ( .A(n1432), .B(sreg[478]), .Z(n1430) );
  XOR U1691 ( .A(n1431), .B(n1430), .Z(c[478]) );
  AND U1692 ( .A(b[0]), .B(a[224]), .Z(n1434) );
  XNOR U1693 ( .A(n1435), .B(sreg[479]), .Z(n1433) );
  XOR U1694 ( .A(n1434), .B(n1433), .Z(c[479]) );
  AND U1695 ( .A(b[0]), .B(a[225]), .Z(n1437) );
  XNOR U1696 ( .A(n1438), .B(sreg[480]), .Z(n1436) );
  XOR U1697 ( .A(n1437), .B(n1436), .Z(c[480]) );
  AND U1698 ( .A(b[0]), .B(a[226]), .Z(n1440) );
  XNOR U1699 ( .A(n1441), .B(sreg[481]), .Z(n1439) );
  XOR U1700 ( .A(n1440), .B(n1439), .Z(c[481]) );
  AND U1701 ( .A(b[0]), .B(a[227]), .Z(n1443) );
  XNOR U1702 ( .A(n1444), .B(sreg[482]), .Z(n1442) );
  XOR U1703 ( .A(n1443), .B(n1442), .Z(c[482]) );
  AND U1704 ( .A(b[0]), .B(a[228]), .Z(n1446) );
  XNOR U1705 ( .A(n1447), .B(sreg[483]), .Z(n1445) );
  XOR U1706 ( .A(n1446), .B(n1445), .Z(c[483]) );
  AND U1707 ( .A(b[0]), .B(a[229]), .Z(n1449) );
  XNOR U1708 ( .A(n1450), .B(sreg[484]), .Z(n1448) );
  XOR U1709 ( .A(n1449), .B(n1448), .Z(c[484]) );
  AND U1710 ( .A(b[0]), .B(a[230]), .Z(n1452) );
  XNOR U1711 ( .A(n1453), .B(sreg[485]), .Z(n1451) );
  XOR U1712 ( .A(n1452), .B(n1451), .Z(c[485]) );
  AND U1713 ( .A(b[0]), .B(a[231]), .Z(n1455) );
  XNOR U1714 ( .A(n1456), .B(sreg[486]), .Z(n1454) );
  XOR U1715 ( .A(n1455), .B(n1454), .Z(c[486]) );
  AND U1716 ( .A(b[0]), .B(a[232]), .Z(n1458) );
  XNOR U1717 ( .A(n1459), .B(sreg[487]), .Z(n1457) );
  XOR U1718 ( .A(n1458), .B(n1457), .Z(c[487]) );
  AND U1719 ( .A(b[0]), .B(a[233]), .Z(n1461) );
  XNOR U1720 ( .A(n1462), .B(sreg[488]), .Z(n1460) );
  XOR U1721 ( .A(n1461), .B(n1460), .Z(c[488]) );
  AND U1722 ( .A(b[0]), .B(a[234]), .Z(n1464) );
  XNOR U1723 ( .A(n1465), .B(sreg[489]), .Z(n1463) );
  XOR U1724 ( .A(n1464), .B(n1463), .Z(c[489]) );
  AND U1725 ( .A(b[0]), .B(a[235]), .Z(n1467) );
  XNOR U1726 ( .A(n1468), .B(sreg[490]), .Z(n1466) );
  XOR U1727 ( .A(n1467), .B(n1466), .Z(c[490]) );
  AND U1728 ( .A(b[0]), .B(a[236]), .Z(n1470) );
  XNOR U1729 ( .A(n1471), .B(sreg[491]), .Z(n1469) );
  XOR U1730 ( .A(n1470), .B(n1469), .Z(c[491]) );
  AND U1731 ( .A(b[0]), .B(a[237]), .Z(n1473) );
  XNOR U1732 ( .A(n1474), .B(sreg[492]), .Z(n1472) );
  XOR U1733 ( .A(n1473), .B(n1472), .Z(c[492]) );
  AND U1734 ( .A(b[0]), .B(a[238]), .Z(n1476) );
  XNOR U1735 ( .A(n1477), .B(sreg[493]), .Z(n1475) );
  XOR U1736 ( .A(n1476), .B(n1475), .Z(c[493]) );
  AND U1737 ( .A(b[0]), .B(a[239]), .Z(n1479) );
  XNOR U1738 ( .A(n1480), .B(sreg[494]), .Z(n1478) );
  XOR U1739 ( .A(n1479), .B(n1478), .Z(c[494]) );
  AND U1740 ( .A(b[0]), .B(a[240]), .Z(n1482) );
  XNOR U1741 ( .A(n1483), .B(sreg[495]), .Z(n1481) );
  XOR U1742 ( .A(n1482), .B(n1481), .Z(c[495]) );
  AND U1743 ( .A(b[0]), .B(a[241]), .Z(n1485) );
  XNOR U1744 ( .A(n1486), .B(sreg[496]), .Z(n1484) );
  XOR U1745 ( .A(n1485), .B(n1484), .Z(c[496]) );
  AND U1746 ( .A(b[0]), .B(a[242]), .Z(n1488) );
  XNOR U1747 ( .A(n1489), .B(sreg[497]), .Z(n1487) );
  XOR U1748 ( .A(n1488), .B(n1487), .Z(c[497]) );
  AND U1749 ( .A(b[0]), .B(a[243]), .Z(n1491) );
  XNOR U1750 ( .A(n1492), .B(sreg[498]), .Z(n1490) );
  XOR U1751 ( .A(n1491), .B(n1490), .Z(c[498]) );
  AND U1752 ( .A(b[0]), .B(a[244]), .Z(n1494) );
  XNOR U1753 ( .A(n1495), .B(sreg[499]), .Z(n1493) );
  XOR U1754 ( .A(n1494), .B(n1493), .Z(c[499]) );
  AND U1755 ( .A(b[0]), .B(a[245]), .Z(n1497) );
  XNOR U1756 ( .A(n1498), .B(sreg[500]), .Z(n1496) );
  XOR U1757 ( .A(n1497), .B(n1496), .Z(c[500]) );
  AND U1758 ( .A(b[0]), .B(a[246]), .Z(n1500) );
  XNOR U1759 ( .A(n1501), .B(sreg[501]), .Z(n1499) );
  XOR U1760 ( .A(n1500), .B(n1499), .Z(c[501]) );
  AND U1761 ( .A(b[0]), .B(a[247]), .Z(n1503) );
  XNOR U1762 ( .A(n1504), .B(sreg[502]), .Z(n1502) );
  XOR U1763 ( .A(n1503), .B(n1502), .Z(c[502]) );
  AND U1764 ( .A(b[0]), .B(a[248]), .Z(n1506) );
  XNOR U1765 ( .A(n1507), .B(sreg[503]), .Z(n1505) );
  XOR U1766 ( .A(n1506), .B(n1505), .Z(c[503]) );
  AND U1767 ( .A(b[0]), .B(a[249]), .Z(n1509) );
  XNOR U1768 ( .A(n1510), .B(sreg[504]), .Z(n1508) );
  XOR U1769 ( .A(n1509), .B(n1508), .Z(c[504]) );
  AND U1770 ( .A(b[0]), .B(a[250]), .Z(n1512) );
  XNOR U1771 ( .A(n1513), .B(sreg[505]), .Z(n1511) );
  XOR U1772 ( .A(n1512), .B(n1511), .Z(c[505]) );
  AND U1773 ( .A(b[0]), .B(a[251]), .Z(n1515) );
  XNOR U1774 ( .A(n1516), .B(sreg[506]), .Z(n1514) );
  XOR U1775 ( .A(n1515), .B(n1514), .Z(c[506]) );
  AND U1776 ( .A(b[0]), .B(a[252]), .Z(n1518) );
  XNOR U1777 ( .A(n1519), .B(sreg[507]), .Z(n1517) );
  XOR U1778 ( .A(n1518), .B(n1517), .Z(c[507]) );
  AND U1779 ( .A(b[0]), .B(a[253]), .Z(n1521) );
  XNOR U1780 ( .A(n1522), .B(sreg[508]), .Z(n1520) );
  XOR U1781 ( .A(n1521), .B(n1520), .Z(c[508]) );
  AND U1782 ( .A(b[0]), .B(a[254]), .Z(n1524) );
  XNOR U1783 ( .A(n1525), .B(sreg[509]), .Z(n1523) );
  XOR U1784 ( .A(n1524), .B(n1523), .Z(c[509]) );
  NAND U1785 ( .A(b[0]), .B(a[255]), .Z(n1526) );
  XNOR U1786 ( .A(sreg[510]), .B(n1528), .Z(n1527) );
  XNOR U1787 ( .A(n1526), .B(n1527), .Z(c[510]) );
  NAND U1788 ( .A(n1527), .B(n1526), .Z(n1530) );
  NANDN U1789 ( .A(sreg[510]), .B(n1528), .Z(n1529) );
  AND U1790 ( .A(n1530), .B(n1529), .Z(c[511]) );
endmodule

