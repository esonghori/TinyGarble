
module modexp_1_N_N4_CC2 ( clk, rst, m, e, n, c );
  input [3:0] m;
  input [3:0] e;
  input [3:0] n;
  output [3:0] c;
  input clk, rst;
  wire   \cin[0][2] , \cin[0][1] , init, \keep_1[0] , N10, N11, N12, N13,
         \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ,
         \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ,
         \MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 , n6, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823;
  wire   [3:0] ein;
  wire   [3:0] ereg;
  assign \MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4  = m[0];

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \ereg_reg[2]  ( .D(ein[0]), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(ein[1]), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \creg_reg[0]  ( .D(N10), .CLK(clk), .RST(rst), .Q(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ) );
  DFF \creg_reg[1]  ( .D(N11), .CLK(clk), .RST(rst), .Q(\cin[0][1] ) );
  DFF \creg_reg[2]  ( .D(N12), .CLK(clk), .RST(rst), .Q(\cin[0][2] ) );
  DFF \creg_reg[3]  ( .D(N13), .CLK(clk), .RST(rst), .Q(
        \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .Q(\keep_1[0] ) );
  XOR U552 ( .A(n960), .B(n959), .Z(n356) );
  NANDN U553 ( .A(n[1]), .B(n356), .Z(n357) );
  NAND U554 ( .A(n960), .B(n959), .Z(n358) );
  AND U555 ( .A(n357), .B(n358), .Z(n964) );
  XOR U556 ( .A(n1529), .B(n1526), .Z(n359) );
  NANDN U557 ( .A(n[1]), .B(n359), .Z(n360) );
  NAND U558 ( .A(n1529), .B(n1526), .Z(n361) );
  AND U559 ( .A(n360), .B(n361), .Z(n1534) );
  NAND U560 ( .A(n1224), .B(n1225), .Z(n362) );
  XOR U561 ( .A(n1224), .B(n1225), .Z(n363) );
  NANDN U562 ( .A(n1223), .B(n363), .Z(n364) );
  NAND U563 ( .A(n362), .B(n364), .Z(n1237) );
  NAND U564 ( .A(n1634), .B(m[2]), .Z(n365) );
  XOR U565 ( .A(n1634), .B(m[2]), .Z(n366) );
  NAND U566 ( .A(n366), .B(n1633), .Z(n367) );
  NAND U567 ( .A(n365), .B(n367), .Z(n1639) );
  NAND U568 ( .A(n709), .B(n1782), .Z(n368) );
  ANDN U569 ( .B(n368), .A(n1797), .Z(n369) );
  NOR U570 ( .A(n[0]), .B(n696), .Z(n370) );
  NAND U571 ( .A(n370), .B(n714), .Z(n371) );
  XOR U572 ( .A(n370), .B(n714), .Z(n372) );
  NANDN U573 ( .A(n[1]), .B(n372), .Z(n373) );
  NAND U574 ( .A(n371), .B(n373), .Z(n374) );
  XNOR U575 ( .A(n709), .B(n[2]), .Z(n375) );
  NAND U576 ( .A(n374), .B(n375), .Z(n376) );
  NAND U577 ( .A(n369), .B(n376), .Z(n377) );
  AND U578 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n377), .Z(n712) );
  XOR U579 ( .A(n1782), .B(n963), .Z(n378) );
  NOR U580 ( .A(n[0]), .B(n956), .Z(n379) );
  NAND U581 ( .A(n379), .B(n960), .Z(n380) );
  XOR U582 ( .A(n379), .B(n960), .Z(n381) );
  NANDN U583 ( .A(n[1]), .B(n381), .Z(n382) );
  NAND U584 ( .A(n380), .B(n382), .Z(n383) );
  NAND U585 ( .A(n378), .B(n383), .Z(n384) );
  NAND U586 ( .A(n1782), .B(n963), .Z(n385) );
  AND U587 ( .A(n384), .B(n385), .Z(n970) );
  NAND U588 ( .A(n[0]), .B(n1279), .Z(n386) );
  NANDN U589 ( .A(n[1]), .B(n1275), .Z(n387) );
  XNOR U590 ( .A(n[1]), .B(n1275), .Z(n388) );
  NAND U591 ( .A(n388), .B(n386), .Z(n389) );
  NAND U592 ( .A(n387), .B(n389), .Z(n390) );
  NAND U593 ( .A(n1293), .B(n1782), .Z(n391) );
  XOR U594 ( .A(n1293), .B(n1782), .Z(n392) );
  NAND U595 ( .A(n392), .B(n390), .Z(n393) );
  NAND U596 ( .A(n391), .B(n393), .Z(n394) );
  ANDN U597 ( .B(n1270), .A(n1797), .Z(n395) );
  NAND U598 ( .A(n1272), .B(n395), .Z(n396) );
  NAND U599 ( .A(n1797), .B(n394), .Z(n397) );
  AND U600 ( .A(n396), .B(n397), .Z(n398) );
  XOR U601 ( .A(n1797), .B(n394), .Z(n399) );
  NAND U602 ( .A(n399), .B(n1292), .Z(n400) );
  AND U603 ( .A(n398), .B(n400), .Z(n1290) );
  NOR U604 ( .A(n[0]), .B(n1531), .Z(n401) );
  NAND U605 ( .A(n401), .B(n1529), .Z(n402) );
  XOR U606 ( .A(n401), .B(n1529), .Z(n403) );
  NANDN U607 ( .A(n[1]), .B(n403), .Z(n404) );
  NAND U608 ( .A(n402), .B(n404), .Z(n405) );
  XOR U609 ( .A(n1782), .B(n1533), .Z(n406) );
  NAND U610 ( .A(n406), .B(n405), .Z(n407) );
  NAND U611 ( .A(n1782), .B(n1533), .Z(n408) );
  AND U612 ( .A(n407), .B(n408), .Z(n1540) );
  XOR U613 ( .A(n1445), .B(n1384), .Z(n409) );
  NAND U614 ( .A(n1445), .B(n1384), .Z(n410) );
  NANDN U615 ( .A(n1381), .B(n409), .Z(n411) );
  NAND U616 ( .A(n410), .B(n411), .Z(n1356) );
  NAND U617 ( .A(n[1]), .B(n1693), .Z(n412) );
  XOR U618 ( .A(n[1]), .B(n1693), .Z(n413) );
  NANDN U619 ( .A(n1690), .B(n413), .Z(n414) );
  NAND U620 ( .A(n412), .B(n414), .Z(n1677) );
  ANDN U621 ( .B(n1186), .A(n[0]), .Z(n415) );
  NAND U622 ( .A(n1193), .B(n415), .Z(n416) );
  NANDN U623 ( .A(n1184), .B(n416), .Z(n417) );
  OR U624 ( .A(n1196), .B(n417), .Z(n418) );
  ANDN U625 ( .B(n418), .A(n1195), .Z(n419) );
  NANDN U626 ( .A(n[3]), .B(n1204), .Z(n420) );
  ANDN U627 ( .B(n420), .A(n1199), .Z(n421) );
  XNOR U628 ( .A(n1204), .B(n[3]), .Z(n422) );
  NAND U629 ( .A(n419), .B(n422), .Z(n423) );
  AND U630 ( .A(n421), .B(n423), .Z(n424) );
  AND U631 ( .A(n1198), .B(n424), .Z(n1202) );
  XNOR U632 ( .A(m[3]), .B(n1722), .Z(n425) );
  AND U633 ( .A(n1806), .B(n425), .Z(n426) );
  XNOR U634 ( .A(n1723), .B(n426), .Z(n1764) );
  XOR U635 ( .A(n729), .B(n728), .Z(n732) );
  NANDN U636 ( .A(n1797), .B(n971), .Z(n427) );
  NANDN U637 ( .A(n970), .B(n[3]), .Z(n428) );
  NANDN U638 ( .A(n971), .B(n428), .Z(n429) );
  AND U639 ( .A(n427), .B(n429), .Z(n430) );
  NAND U640 ( .A(n972), .B(n430), .Z(n431) );
  NANDN U641 ( .A(n[1]), .B(n980), .Z(n432) );
  XNOR U642 ( .A(n[1]), .B(n980), .Z(n433) );
  NAND U643 ( .A(n[0]), .B(n976), .Z(n434) );
  NAND U644 ( .A(n433), .B(n434), .Z(n435) );
  NAND U645 ( .A(n432), .B(n435), .Z(n436) );
  XOR U646 ( .A(n1782), .B(n436), .Z(n437) );
  NAND U647 ( .A(n437), .B(n992), .Z(n438) );
  NAND U648 ( .A(n1782), .B(n436), .Z(n439) );
  AND U649 ( .A(n438), .B(n439), .Z(n440) );
  OR U650 ( .A(n1797), .B(n1007), .Z(n441) );
  NANDN U651 ( .A(n440), .B(n441), .Z(n442) );
  AND U652 ( .A(n431), .B(n442), .Z(n1005) );
  XOR U653 ( .A(n1262), .B(n1259), .Z(n443) );
  NANDN U654 ( .A(n[1]), .B(n443), .Z(n444) );
  NAND U655 ( .A(n1262), .B(n1259), .Z(n445) );
  AND U656 ( .A(n444), .B(n445), .Z(n1265) );
  XNOR U657 ( .A(m[3]), .B(n1000), .Z(n446) );
  AND U658 ( .A(n1220), .B(n446), .Z(n447) );
  XNOR U659 ( .A(n998), .B(n447), .Z(n1051) );
  NAND U660 ( .A(n[0]), .B(n1551), .Z(n448) );
  NANDN U661 ( .A(n[1]), .B(n1545), .Z(n449) );
  XNOR U662 ( .A(n[1]), .B(n1545), .Z(n450) );
  NAND U663 ( .A(n450), .B(n448), .Z(n451) );
  NAND U664 ( .A(n449), .B(n451), .Z(n452) );
  XOR U665 ( .A(n1782), .B(n452), .Z(n453) );
  NAND U666 ( .A(n453), .B(n1556), .Z(n454) );
  NAND U667 ( .A(n1782), .B(n452), .Z(n455) );
  AND U668 ( .A(n454), .B(n455), .Z(n456) );
  NANDN U669 ( .A(n1540), .B(n[3]), .Z(n457) );
  NANDN U670 ( .A(n1797), .B(n1541), .Z(n458) );
  NANDN U671 ( .A(n1541), .B(n457), .Z(n459) );
  AND U672 ( .A(n458), .B(n459), .Z(n460) );
  NAND U673 ( .A(n1542), .B(n460), .Z(n461) );
  OR U674 ( .A(n1797), .B(n1571), .Z(n462) );
  NANDN U675 ( .A(n456), .B(n462), .Z(n463) );
  AND U676 ( .A(n461), .B(n463), .Z(n1569) );
  NOR U677 ( .A(n[0]), .B(n891), .Z(n464) );
  NANDN U678 ( .A(n829), .B(n464), .Z(n465) );
  NANDN U679 ( .A(n830), .B(n465), .Z(n466) );
  ANDN U680 ( .B(n843), .A(n844), .Z(n467) );
  OR U681 ( .A(n466), .B(n841), .Z(n468) );
  AND U682 ( .A(n467), .B(n468), .Z(n469) );
  NOR U683 ( .A(n849), .B(n839), .Z(n470) );
  ANDN U684 ( .B(n470), .A(n469), .Z(n471) );
  NANDN U685 ( .A(n848), .B(n471), .Z(n852) );
  ANDN U686 ( .B(n1320), .A(n[1]), .Z(n1322) );
  ANDN U687 ( .B(n1605), .A(n[1]), .Z(n1594) );
  XNOR U688 ( .A(m[3]), .B(n1564), .Z(n472) );
  AND U689 ( .A(n1814), .B(n472), .Z(n473) );
  XNOR U690 ( .A(n1562), .B(n473), .Z(n1601) );
  AND U691 ( .A(n[1]), .B(n1394), .Z(n1396) );
  AND U692 ( .A(n[0]), .B(n1709), .Z(n474) );
  NAND U693 ( .A(n1703), .B(n[1]), .Z(n475) );
  XOR U694 ( .A(n1703), .B(n[1]), .Z(n476) );
  NAND U695 ( .A(n476), .B(n474), .Z(n477) );
  NAND U696 ( .A(n475), .B(n477), .Z(n478) );
  XNOR U697 ( .A(n1782), .B(n1699), .Z(n479) );
  NAND U698 ( .A(n478), .B(n479), .Z(n480) );
  NAND U699 ( .A(n1697), .B(n480), .Z(n481) );
  OR U700 ( .A(n1797), .B(n1726), .Z(n482) );
  NANDN U701 ( .A(n481), .B(n482), .Z(n483) );
  ANDN U702 ( .B(n483), .A(n1698), .Z(n1704) );
  NANDN U703 ( .A(n1200), .B(n1204), .Z(n484) );
  NANDN U704 ( .A(n1797), .B(n484), .Z(n485) );
  NANDN U705 ( .A(n1198), .B(n485), .Z(n486) );
  ANDN U706 ( .B(n486), .A(n1199), .Z(n487) );
  NANDN U707 ( .A(n[3]), .B(n1244), .Z(n488) );
  AND U708 ( .A(n487), .B(n488), .Z(n489) );
  XNOR U709 ( .A(n[3]), .B(n1244), .Z(n490) );
  NANDN U710 ( .A(n[1]), .B(n1225), .Z(n491) );
  XNOR U711 ( .A(n[1]), .B(n1225), .Z(n492) );
  NAND U712 ( .A(n[0]), .B(n1212), .Z(n493) );
  NAND U713 ( .A(n492), .B(n493), .Z(n494) );
  NAND U714 ( .A(n491), .B(n494), .Z(n495) );
  XNOR U715 ( .A(n1236), .B(n1782), .Z(n496) );
  NANDN U716 ( .A(n495), .B(n496), .Z(n497) );
  NANDN U717 ( .A(n1782), .B(n1236), .Z(n498) );
  AND U718 ( .A(n497), .B(n498), .Z(n499) );
  NAND U719 ( .A(n490), .B(n499), .Z(n500) );
  AND U720 ( .A(n489), .B(n500), .Z(n1240) );
  ANDN U721 ( .B(n1746), .A(n[0]), .Z(n501) );
  NAND U722 ( .A(n1743), .B(n501), .Z(n502) );
  NANDN U723 ( .A(n1744), .B(n502), .Z(n503) );
  OR U724 ( .A(n1756), .B(n503), .Z(n504) );
  ANDN U725 ( .B(n504), .A(n1755), .Z(n505) );
  NANDN U726 ( .A(n[3]), .B(n1764), .Z(n506) );
  ANDN U727 ( .B(n506), .A(n1759), .Z(n507) );
  XNOR U728 ( .A(n1764), .B(n[3]), .Z(n508) );
  NAND U729 ( .A(n505), .B(n508), .Z(n509) );
  AND U730 ( .A(n507), .B(n509), .Z(n510) );
  NANDN U731 ( .A(n1758), .B(n510), .Z(n1762) );
  XNOR U732 ( .A(n981), .B(n980), .Z(n982) );
  AND U733 ( .A(n[0]), .B(n717), .Z(n511) );
  NAND U734 ( .A(n511), .B(n[1]), .Z(n512) );
  XOR U735 ( .A(n511), .B(n[1]), .Z(n513) );
  NANDN U736 ( .A(n726), .B(n513), .Z(n514) );
  NAND U737 ( .A(n512), .B(n514), .Z(n515) );
  NANDN U738 ( .A(n1797), .B(n744), .Z(n516) );
  NANDN U739 ( .A(n744), .B(n1782), .Z(n517) );
  NANDN U740 ( .A(n747), .B(n517), .Z(n518) );
  NAND U741 ( .A(n516), .B(n518), .Z(n519) );
  NAND U742 ( .A(n1782), .B(n747), .Z(n520) );
  NAND U743 ( .A(n515), .B(n520), .Z(n521) );
  NANDN U744 ( .A(n519), .B(n521), .Z(n743) );
  ANDN U745 ( .B(n764), .A(n[1]), .Z(n756) );
  ANDN U746 ( .B(n1033), .A(n[1]), .Z(n1024) );
  XNOR U747 ( .A(n822), .B(n823), .Z(n848) );
  NAND U748 ( .A(n1300), .B(n1299), .Z(n522) );
  XNOR U749 ( .A(n1302), .B(n522), .Z(n523) );
  NAND U750 ( .A(n1302), .B(n1301), .Z(n524) );
  NAND U751 ( .A(n523), .B(n524), .Z(n1343) );
  OR U752 ( .A(n1602), .B(n1594), .Z(n525) );
  AND U753 ( .A(n1595), .B(n525), .Z(n1606) );
  XOR U754 ( .A(n864), .B(n863), .Z(n867) );
  AND U755 ( .A(n[0]), .B(n1136), .Z(n526) );
  XOR U756 ( .A(n[1]), .B(n1145), .Z(n527) );
  NAND U757 ( .A(n527), .B(n526), .Z(n528) );
  NAND U758 ( .A(n[1]), .B(n1145), .Z(n529) );
  AND U759 ( .A(n528), .B(n529), .Z(n530) );
  XNOR U760 ( .A(n1782), .B(n1141), .Z(n531) );
  NANDN U761 ( .A(n530), .B(n531), .Z(n532) );
  AND U762 ( .A(n1140), .B(n532), .Z(n533) );
  OR U763 ( .A(n1797), .B(n1163), .Z(n534) );
  NAND U764 ( .A(n533), .B(n534), .Z(n535) );
  NANDN U765 ( .A(n1139), .B(n535), .Z(n1162) );
  NAND U766 ( .A(n941), .B(n942), .Z(n536) );
  XOR U767 ( .A(n941), .B(n942), .Z(n537) );
  NANDN U768 ( .A(n940), .B(n537), .Z(n538) );
  NAND U769 ( .A(n536), .B(n538), .Z(n944) );
  XOR U770 ( .A(n1369), .B(n1368), .Z(n1374) );
  AND U771 ( .A(n[0]), .B(n1444), .Z(n539) );
  NAND U772 ( .A(n1420), .B(n[1]), .Z(n540) );
  XOR U773 ( .A(n1420), .B(n[1]), .Z(n541) );
  NAND U774 ( .A(n541), .B(n539), .Z(n542) );
  NAND U775 ( .A(n540), .B(n542), .Z(n543) );
  XNOR U776 ( .A(n1782), .B(n1426), .Z(n544) );
  NAND U777 ( .A(n543), .B(n544), .Z(n545) );
  NAND U778 ( .A(n1424), .B(n545), .Z(n546) );
  NANDN U779 ( .A(n1797), .B(n1433), .Z(n547) );
  NANDN U780 ( .A(n546), .B(n547), .Z(n548) );
  ANDN U781 ( .B(n548), .A(n1423), .Z(n1425) );
  XNOR U782 ( .A(n[1]), .B(n1190), .Z(n549) );
  ANDN U783 ( .B(n549), .A(n1202), .Z(n550) );
  XNOR U784 ( .A(n1191), .B(n550), .Z(n1225) );
  XNOR U785 ( .A(n1657), .B(n1658), .Z(n1682) );
  OR U786 ( .A(n1703), .B(n1702), .Z(n551) );
  NAND U787 ( .A(n1707), .B(n1706), .Z(n552) );
  AND U788 ( .A(n551), .B(n552), .Z(n1718) );
  ANDN U789 ( .B(n1505), .A(n1797), .Z(n553) );
  OR U790 ( .A(n1507), .B(n1506), .Z(n554) );
  AND U791 ( .A(n553), .B(n554), .Z(n555) );
  AND U792 ( .A(n[0]), .B(n1510), .Z(n556) );
  NAND U793 ( .A(n1620), .B(n[1]), .Z(n557) );
  XOR U794 ( .A(n1620), .B(n[1]), .Z(n558) );
  NAND U795 ( .A(n558), .B(n556), .Z(n559) );
  NAND U796 ( .A(n557), .B(n559), .Z(n560) );
  XNOR U797 ( .A(n1782), .B(n1512), .Z(n561) );
  NAND U798 ( .A(n561), .B(n560), .Z(n562) );
  NANDN U799 ( .A(n1782), .B(n1512), .Z(n563) );
  NAND U800 ( .A(n562), .B(n563), .Z(n564) );
  OR U801 ( .A(n564), .B(n1521), .Z(n565) );
  ANDN U802 ( .B(n565), .A(n1498), .Z(n566) );
  XOR U803 ( .A(n564), .B(n1521), .Z(n567) );
  NAND U804 ( .A(n1797), .B(n567), .Z(n568) );
  NAND U805 ( .A(n566), .B(n568), .Z(n569) );
  XNOR U806 ( .A(n1508), .B(n555), .Z(n570) );
  NANDN U807 ( .A(n569), .B(n570), .Z(n1517) );
  AND U808 ( .A(n[0]), .B(n1775), .Z(n571) );
  XOR U809 ( .A(n[1]), .B(n1781), .Z(n572) );
  NAND U810 ( .A(n572), .B(n571), .Z(n573) );
  NAND U811 ( .A(n[1]), .B(n1781), .Z(n574) );
  AND U812 ( .A(n573), .B(n574), .Z(n575) );
  XNOR U813 ( .A(n1792), .B(n1782), .Z(n576) );
  NANDN U814 ( .A(n575), .B(n576), .Z(n577) );
  NANDN U815 ( .A(n1782), .B(n1792), .Z(n578) );
  AND U816 ( .A(n577), .B(n578), .Z(n579) );
  ANDN U817 ( .B(n1762), .A(n1797), .Z(n580) );
  NANDN U818 ( .A(n1760), .B(n1764), .Z(n581) );
  AND U819 ( .A(n580), .B(n581), .Z(n582) );
  XNOR U820 ( .A(n582), .B(n1758), .Z(n583) );
  NANDN U821 ( .A(n1759), .B(n583), .Z(n584) );
  NANDN U822 ( .A(n[3]), .B(n579), .Z(n585) );
  ANDN U823 ( .B(n585), .A(n584), .Z(n586) );
  XNOR U824 ( .A(n579), .B(n[3]), .Z(n587) );
  NAND U825 ( .A(n587), .B(n1801), .Z(n588) );
  NAND U826 ( .A(n586), .B(n588), .Z(n1796) );
  XNOR U827 ( .A(n727), .B(n726), .Z(n728) );
  XNOR U828 ( .A(n983), .B(n982), .Z(n987) );
  ANDN U829 ( .B(n[0]), .A(n786), .Z(n589) );
  XOR U830 ( .A(n[1]), .B(n790), .Z(n590) );
  NAND U831 ( .A(n590), .B(n589), .Z(n591) );
  NAND U832 ( .A(n[1]), .B(n790), .Z(n592) );
  AND U833 ( .A(n591), .B(n592), .Z(n593) );
  XNOR U834 ( .A(n[2]), .B(n809), .Z(n594) );
  NAND U835 ( .A(n594), .B(n593), .Z(n595) );
  NANDN U836 ( .A(n[2]), .B(n809), .Z(n596) );
  NAND U837 ( .A(n595), .B(n596), .Z(n597) );
  NAND U838 ( .A(n779), .B(n778), .Z(n598) );
  NANDN U839 ( .A(n825), .B(n598), .Z(n599) );
  NANDN U840 ( .A(n[3]), .B(n597), .Z(n600) );
  ANDN U841 ( .B(n600), .A(n599), .Z(n601) );
  XNOR U842 ( .A(n[3]), .B(n597), .Z(n602) );
  NAND U843 ( .A(n602), .B(n819), .Z(n603) );
  NAND U844 ( .A(n601), .B(n603), .Z(n815) );
  ANDN U845 ( .B(n[0]), .A(n1059), .Z(n604) );
  XOR U846 ( .A(n[1]), .B(n1053), .Z(n605) );
  NAND U847 ( .A(n605), .B(n604), .Z(n606) );
  NAND U848 ( .A(n[1]), .B(n1053), .Z(n607) );
  AND U849 ( .A(n606), .B(n607), .Z(n608) );
  XNOR U850 ( .A(n[2]), .B(n1072), .Z(n609) );
  NAND U851 ( .A(n609), .B(n608), .Z(n610) );
  NANDN U852 ( .A(n[2]), .B(n1072), .Z(n611) );
  NAND U853 ( .A(n610), .B(n611), .Z(n612) );
  NAND U854 ( .A(n1088), .B(n1046), .Z(n613) );
  NANDN U855 ( .A(n[3]), .B(n612), .Z(n614) );
  ANDN U856 ( .B(n614), .A(n613), .Z(n615) );
  XNOR U857 ( .A(n[3]), .B(n612), .Z(n616) );
  NAND U858 ( .A(n616), .B(n1080), .Z(n617) );
  NAND U859 ( .A(n615), .B(n617), .Z(n1078) );
  NAND U860 ( .A(n1266), .B(n1272), .Z(n618) );
  XNOR U861 ( .A(n1267), .B(n618), .Z(n1293) );
  AND U862 ( .A(n[0]), .B(n856), .Z(n619) );
  XOR U863 ( .A(n[1]), .B(n862), .Z(n620) );
  NAND U864 ( .A(n620), .B(n619), .Z(n621) );
  NAND U865 ( .A(n[1]), .B(n862), .Z(n622) );
  AND U866 ( .A(n621), .B(n622), .Z(n623) );
  XNOR U867 ( .A(n[2]), .B(n877), .Z(n624) );
  NAND U868 ( .A(n624), .B(n623), .Z(n625) );
  NANDN U869 ( .A(n[2]), .B(n877), .Z(n626) );
  NAND U870 ( .A(n625), .B(n626), .Z(n627) );
  OR U871 ( .A(n906), .B(n849), .Z(n628) );
  NANDN U872 ( .A(n[3]), .B(n627), .Z(n629) );
  ANDN U873 ( .B(n629), .A(n628), .Z(n630) );
  XNOR U874 ( .A(n[3]), .B(n627), .Z(n631) );
  NAND U875 ( .A(n631), .B(n900), .Z(n632) );
  NAND U876 ( .A(n630), .B(n632), .Z(n883) );
  NAND U877 ( .A(n[1]), .B(n1132), .Z(n633) );
  XOR U878 ( .A(n[1]), .B(n1132), .Z(n634) );
  NANDN U879 ( .A(n1128), .B(n634), .Z(n635) );
  NAND U880 ( .A(n633), .B(n635), .Z(n1123) );
  XNOR U881 ( .A(n1085), .B(n1086), .Z(n1115) );
  XNOR U882 ( .A(n1159), .B(n1158), .Z(n1168) );
  AND U883 ( .A(n[0]), .B(n1346), .Z(n636) );
  XOR U884 ( .A(n[1]), .B(n1348), .Z(n637) );
  NAND U885 ( .A(n637), .B(n636), .Z(n638) );
  NAND U886 ( .A(n[1]), .B(n1348), .Z(n639) );
  AND U887 ( .A(n638), .B(n639), .Z(n640) );
  XOR U888 ( .A(n1782), .B(n1361), .Z(n641) );
  NAND U889 ( .A(n641), .B(n640), .Z(n642) );
  NAND U890 ( .A(n1782), .B(n1361), .Z(n643) );
  AND U891 ( .A(n642), .B(n643), .Z(n644) );
  NANDN U892 ( .A(n1797), .B(n644), .Z(n645) );
  XNOR U893 ( .A(n644), .B(n1797), .Z(n646) );
  NAND U894 ( .A(n646), .B(n1371), .Z(n647) );
  NAND U895 ( .A(n645), .B(n647), .Z(n648) );
  ANDN U896 ( .B(n648), .A(n1377), .Z(n649) );
  NAND U897 ( .A(n649), .B(n1343), .Z(n1367) );
  AND U898 ( .A(n[0]), .B(n1624), .Z(n650) );
  XOR U899 ( .A(n[1]), .B(n1628), .Z(n651) );
  NAND U900 ( .A(n651), .B(n650), .Z(n652) );
  NAND U901 ( .A(n[1]), .B(n1628), .Z(n653) );
  AND U902 ( .A(n652), .B(n653), .Z(n654) );
  NAND U903 ( .A(n1644), .B(n1782), .Z(n655) );
  XOR U904 ( .A(n1644), .B(n1782), .Z(n656) );
  NAND U905 ( .A(n656), .B(n654), .Z(n657) );
  NAND U906 ( .A(n655), .B(n657), .Z(n658) );
  NAND U907 ( .A(n1654), .B(n1797), .Z(n659) );
  ANDN U908 ( .B(n659), .A(n1660), .Z(n660) );
  XOR U909 ( .A(n1654), .B(n1797), .Z(n661) );
  NAND U910 ( .A(n661), .B(n658), .Z(n662) );
  AND U911 ( .A(n660), .B(n662), .Z(n663) );
  NAND U912 ( .A(n663), .B(n1618), .Z(n1650) );
  NAND U913 ( .A(n[0]), .B(n1134), .Z(n664) );
  NANDN U914 ( .A(n[1]), .B(n942), .Z(n665) );
  XNOR U915 ( .A(n[1]), .B(n942), .Z(n666) );
  NAND U916 ( .A(n666), .B(n664), .Z(n667) );
  NAND U917 ( .A(n665), .B(n667), .Z(n668) );
  XNOR U918 ( .A(n943), .B(n1782), .Z(n669) );
  NANDN U919 ( .A(n668), .B(n669), .Z(n670) );
  NANDN U920 ( .A(n1782), .B(n943), .Z(n671) );
  AND U921 ( .A(n670), .B(n671), .Z(n672) );
  NANDN U922 ( .A(n934), .B(n938), .Z(n673) );
  NANDN U923 ( .A(n1797), .B(n673), .Z(n674) );
  NANDN U924 ( .A(n932), .B(n674), .Z(n675) );
  ANDN U925 ( .B(n675), .A(n933), .Z(n676) );
  NANDN U926 ( .A(n[3]), .B(n951), .Z(n677) );
  AND U927 ( .A(n676), .B(n677), .Z(n678) );
  XNOR U928 ( .A(n[3]), .B(n951), .Z(n679) );
  NAND U929 ( .A(n679), .B(n672), .Z(n680) );
  AND U930 ( .A(n678), .B(n680), .Z(n947) );
  NAND U931 ( .A(n1212), .B(n1211), .Z(n1224) );
  XNOR U932 ( .A(n1718), .B(n1717), .Z(n1705) );
  XNOR U933 ( .A(n1438), .B(n1439), .Z(n1461) );
  NOR U934 ( .A(n1411), .B(n1412), .Z(n681) );
  OR U935 ( .A(n1413), .B(n1414), .Z(n682) );
  NAND U936 ( .A(n681), .B(n682), .Z(n683) );
  XNOR U937 ( .A(n1415), .B(n683), .Z(n1454) );
  NOR U938 ( .A(n1694), .B(n1676), .Z(n684) );
  OR U939 ( .A(n1684), .B(n1681), .Z(n685) );
  NAND U940 ( .A(n684), .B(n685), .Z(n686) );
  XNOR U941 ( .A(n1682), .B(n686), .Z(n1733) );
  XOR U942 ( .A(n1620), .B(n1622), .Z(n687) );
  NAND U943 ( .A(n687), .B(n1619), .Z(n688) );
  NAND U944 ( .A(n1620), .B(n1622), .Z(n689) );
  AND U945 ( .A(n688), .B(n689), .Z(n1511) );
  XOR U946 ( .A(n1781), .B(n1779), .Z(n690) );
  NANDN U947 ( .A(n1780), .B(n690), .Z(n691) );
  NAND U948 ( .A(n1781), .B(n1779), .Z(n692) );
  AND U949 ( .A(n691), .B(n692), .Z(n1793) );
  NANDN U950 ( .A(\keep_1[0] ), .B(n1765), .Z(n1823) );
  NAND U951 ( .A(ereg[3]), .B(init), .Z(n694) );
  NANDN U952 ( .A(init), .B(e[3]), .Z(n693) );
  AND U953 ( .A(n694), .B(n693), .Z(n1765) );
  ANDN U954 ( .B(\keep_1[0] ), .A(n1765), .Z(n1246) );
  IV U955 ( .A(n1246), .Z(n1227) );
  IV U956 ( .A(n[2]), .Z(n1782) );
  NAND U957 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[0][1] ), .Z(n891) );
  IV U958 ( .A(n891), .Z(n913) );
  NAND U959 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), .Z(
        n696) );
  AND U960 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(\cin[0][2] ), .Z(n709) );
  IV U961 ( .A(n[3]), .Z(n1797) );
  AND U962 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(\cin[0][1] ), .Z(n714) );
  NAND U963 ( .A(n712), .B(n[0]), .Z(n695) );
  XNOR U964 ( .A(n696), .B(n695), .Z(n717) );
  AND U965 ( .A(n[0]), .B(n696), .Z(n698) );
  IV U966 ( .A(n698), .Z(n710) );
  ANDN U967 ( .B(n[1]), .A(n710), .Z(n697) );
  NANDN U968 ( .A(n697), .B(n714), .Z(n700) );
  NOR U969 ( .A(n698), .B(n[1]), .Z(n699) );
  ANDN U970 ( .B(n700), .A(n699), .Z(n701) );
  NANDN U971 ( .A(n1782), .B(n701), .Z(n703) );
  XNOR U972 ( .A(n1782), .B(n701), .Z(n707) );
  NANDN U973 ( .A(n709), .B(n707), .Z(n702) );
  NAND U974 ( .A(n703), .B(n702), .Z(n704) );
  NANDN U975 ( .A(n704), .B(n1797), .Z(n705) );
  NAND U976 ( .A(n712), .B(n705), .Z(n706) );
  NAND U977 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n706), .Z(n744) );
  NAND U978 ( .A(n712), .B(n707), .Z(n708) );
  XNOR U979 ( .A(n709), .B(n708), .Z(n747) );
  XNOR U980 ( .A(n[1]), .B(n710), .Z(n711) );
  NAND U981 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U982 ( .A(n714), .B(n713), .Z(n726) );
  NANDN U983 ( .A(n744), .B(n1797), .Z(n715) );
  AND U984 ( .A(n743), .B(n715), .Z(n725) );
  ANDN U985 ( .B(n[0]), .A(n725), .Z(n716) );
  AND U986 ( .A(n717), .B(n716), .Z(n729) );
  ANDN U987 ( .B(n[1]), .A(n725), .Z(n727) );
  XOR U988 ( .A(n717), .B(n716), .Z(n720) );
  NANDN U989 ( .A(n720), .B(\cin[0][1] ), .Z(n733) );
  NAND U990 ( .A(n733), .B(\cin[0][2] ), .Z(n718) );
  XNOR U991 ( .A(n732), .B(n718), .Z(n769) );
  NAND U992 ( .A(\cin[0][2] ), .B(\cin[0][1] ), .Z(n719) );
  XOR U993 ( .A(n720), .B(n719), .Z(n764) );
  NANDN U994 ( .A(n764), .B(n[1]), .Z(n758) );
  NAND U995 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[0][2] ), .Z(n766) );
  NOR U996 ( .A(n766), .B(n[0]), .Z(n721) );
  NAND U997 ( .A(n758), .B(n721), .Z(n722) );
  NANDN U998 ( .A(n756), .B(n722), .Z(n723) );
  OR U999 ( .A(n723), .B(n1782), .Z(n724) );
  ANDN U1000 ( .B(n724), .A(n769), .Z(n738) );
  NOR U1001 ( .A(n1782), .B(n725), .Z(n746) );
  XNOR U1002 ( .A(n747), .B(n746), .Z(n749) );
  NANDN U1003 ( .A(n727), .B(n726), .Z(n731) );
  NANDN U1004 ( .A(n729), .B(n728), .Z(n730) );
  NAND U1005 ( .A(n731), .B(n730), .Z(n748) );
  XOR U1006 ( .A(n749), .B(n748), .Z(n741) );
  OR U1007 ( .A(n741), .B(\cin[0][2] ), .Z(n737) );
  NAND U1008 ( .A(n733), .B(n732), .Z(n740) );
  NANDN U1009 ( .A(n741), .B(
        \MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), .Z(n734)
         );
  XOR U1010 ( .A(n740), .B(n734), .Z(n735) );
  NAND U1011 ( .A(\cin[0][2] ), .B(n735), .Z(n736) );
  NAND U1012 ( .A(n737), .B(n736), .Z(n784) );
  NANDN U1013 ( .A(n1797), .B(n784), .Z(n772) );
  NAND U1014 ( .A(n738), .B(n772), .Z(n739) );
  ANDN U1015 ( .B(n1797), .A(n784), .Z(n775) );
  ANDN U1016 ( .B(n739), .A(n775), .Z(n755) );
  OR U1017 ( .A(n741), .B(n740), .Z(n742) );
  AND U1018 ( .A(\cin[0][2] ), .B(n742), .Z(n779) );
  OR U1019 ( .A(n743), .B(n1797), .Z(n745) );
  ANDN U1020 ( .B(n745), .A(n744), .Z(n753) );
  ANDN U1021 ( .B(n747), .A(n746), .Z(n751) );
  AND U1022 ( .A(n749), .B(n748), .Z(n750) );
  NOR U1023 ( .A(n751), .B(n750), .Z(n752) );
  XOR U1024 ( .A(n753), .B(n752), .Z(n778) );
  OR U1025 ( .A(n779), .B(n778), .Z(n754) );
  ANDN U1026 ( .B(n755), .A(n754), .Z(n781) );
  AND U1027 ( .A(n[0]), .B(n766), .Z(n761) );
  NANDN U1028 ( .A(n756), .B(n761), .Z(n757) );
  NAND U1029 ( .A(n758), .B(n757), .Z(n767) );
  XOR U1030 ( .A(n[2]), .B(n767), .Z(n759) );
  NANDN U1031 ( .A(n781), .B(n759), .Z(n760) );
  XOR U1032 ( .A(n769), .B(n760), .Z(n809) );
  XOR U1033 ( .A(n[1]), .B(n761), .Z(n762) );
  NANDN U1034 ( .A(n781), .B(n762), .Z(n763) );
  XOR U1035 ( .A(n764), .B(n763), .Z(n790) );
  NANDN U1036 ( .A(n781), .B(n[0]), .Z(n765) );
  XOR U1037 ( .A(n766), .B(n765), .Z(n786) );
  XNOR U1038 ( .A(n1782), .B(n769), .Z(n768) );
  NAND U1039 ( .A(n768), .B(n767), .Z(n771) );
  NANDN U1040 ( .A(n1782), .B(n769), .Z(n770) );
  AND U1041 ( .A(n771), .B(n770), .Z(n780) );
  NAND U1042 ( .A(n780), .B(n772), .Z(n773) );
  ANDN U1043 ( .B(n773), .A(n781), .Z(n774) );
  NANDN U1044 ( .A(n775), .B(n774), .Z(n777) );
  XNOR U1045 ( .A(n779), .B(n778), .Z(n776) );
  XOR U1046 ( .A(n777), .B(n776), .Z(n825) );
  XOR U1047 ( .A(n780), .B(n1797), .Z(n782) );
  ANDN U1048 ( .B(n782), .A(n781), .Z(n783) );
  XNOR U1049 ( .A(n784), .B(n783), .Z(n819) );
  AND U1050 ( .A(n[0]), .B(n815), .Z(n785) );
  ANDN U1051 ( .B(n785), .A(n786), .Z(n792) );
  NAND U1052 ( .A(n[1]), .B(n815), .Z(n789) );
  XNOR U1053 ( .A(n790), .B(n789), .Z(n791) );
  XOR U1054 ( .A(n792), .B(n791), .Z(n795) );
  XOR U1055 ( .A(n786), .B(n785), .Z(n801) );
  XOR U1056 ( .A(\cin[0][2] ), .B(n801), .Z(n787) );
  NAND U1057 ( .A(\cin[0][1] ), .B(n787), .Z(n788) );
  XOR U1058 ( .A(n795), .B(n788), .Z(n834) );
  OR U1059 ( .A(n834), .B(n1782), .Z(n843) );
  ANDN U1060 ( .B(n815), .A(n1782), .Z(n810) );
  XNOR U1061 ( .A(n809), .B(n810), .Z(n812) );
  NANDN U1062 ( .A(n790), .B(n789), .Z(n794) );
  NANDN U1063 ( .A(n792), .B(n791), .Z(n793) );
  NAND U1064 ( .A(n794), .B(n793), .Z(n811) );
  XOR U1065 ( .A(n812), .B(n811), .Z(n803) );
  IV U1066 ( .A(n803), .Z(n802) );
  NANDN U1067 ( .A(n795), .B(\cin[0][2] ), .Z(n798) );
  XNOR U1068 ( .A(\cin[0][2] ), .B(n795), .Z(n796) );
  NAND U1069 ( .A(n801), .B(n796), .Z(n797) );
  NAND U1070 ( .A(n798), .B(n797), .Z(n804) );
  XOR U1071 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n804), .Z(n799) );
  NAND U1072 ( .A(\cin[0][1] ), .B(n799), .Z(n800) );
  XOR U1073 ( .A(n802), .B(n800), .Z(n854) );
  NOR U1074 ( .A(n1797), .B(n854), .Z(n844) );
  XNOR U1075 ( .A(\cin[0][1] ), .B(n801), .Z(n838) );
  NOR U1076 ( .A(n838), .B(n[1]), .Z(n830) );
  AND U1077 ( .A(n[1]), .B(n838), .Z(n829) );
  AND U1078 ( .A(n834), .B(n1782), .Z(n841) );
  AND U1079 ( .A(n854), .B(n1797), .Z(n839) );
  ANDN U1080 ( .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .A(n802), .Z(n807) );
  XOR U1081 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n803), .Z(n805) );
  AND U1082 ( .A(n805), .B(n804), .Z(n806) );
  OR U1083 ( .A(n807), .B(n806), .Z(n808) );
  AND U1084 ( .A(\cin[0][1] ), .B(n808), .Z(n823) );
  NANDN U1085 ( .A(n810), .B(n809), .Z(n814) );
  NAND U1086 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1087 ( .A(n814), .B(n813), .Z(n816) );
  NANDN U1088 ( .A(n1797), .B(n815), .Z(n818) );
  XOR U1089 ( .A(n819), .B(n818), .Z(n817) );
  XNOR U1090 ( .A(n816), .B(n817), .Z(n822) );
  NAND U1091 ( .A(n817), .B(n816), .Z(n821) );
  NAND U1092 ( .A(n819), .B(n818), .Z(n820) );
  AND U1093 ( .A(n821), .B(n820), .Z(n827) );
  ANDN U1094 ( .B(n823), .A(n822), .Z(n824) );
  XNOR U1095 ( .A(n825), .B(n824), .Z(n826) );
  XNOR U1096 ( .A(n827), .B(n826), .Z(n849) );
  NAND U1097 ( .A(n852), .B(n[0]), .Z(n828) );
  XOR U1098 ( .A(n913), .B(n828), .Z(n856) );
  ANDN U1099 ( .B(n[0]), .A(n913), .Z(n835) );
  OR U1100 ( .A(n829), .B(n835), .Z(n831) );
  ANDN U1101 ( .B(n831), .A(n830), .Z(n840) );
  XNOR U1102 ( .A(n1782), .B(n840), .Z(n832) );
  NAND U1103 ( .A(n852), .B(n832), .Z(n833) );
  XNOR U1104 ( .A(n834), .B(n833), .Z(n877) );
  XOR U1105 ( .A(n[1]), .B(n835), .Z(n836) );
  NAND U1106 ( .A(n852), .B(n836), .Z(n837) );
  XNOR U1107 ( .A(n838), .B(n837), .Z(n862) );
  ANDN U1108 ( .B(n852), .A(n839), .Z(n846) );
  NANDN U1109 ( .A(n841), .B(n840), .Z(n842) );
  AND U1110 ( .A(n843), .B(n842), .Z(n850) );
  NANDN U1111 ( .A(n844), .B(n850), .Z(n845) );
  AND U1112 ( .A(n846), .B(n845), .Z(n847) );
  XOR U1113 ( .A(n848), .B(n847), .Z(n906) );
  XOR U1114 ( .A(n1797), .B(n850), .Z(n851) );
  NAND U1115 ( .A(n852), .B(n851), .Z(n853) );
  XNOR U1116 ( .A(n854), .B(n853), .Z(n900) );
  AND U1117 ( .A(n[0]), .B(n883), .Z(n855) );
  NAND U1118 ( .A(n856), .B(n855), .Z(n863) );
  NAND U1119 ( .A(n[1]), .B(n883), .Z(n861) );
  XOR U1120 ( .A(n862), .B(n861), .Z(n864) );
  XNOR U1121 ( .A(\cin[0][2] ), .B(n867), .Z(n868) );
  XOR U1122 ( .A(n856), .B(n855), .Z(n915) );
  ANDN U1123 ( .B(\cin[0][1] ), .A(n915), .Z(n857) );
  XOR U1124 ( .A(n868), .B(n857), .Z(n858) );
  NAND U1125 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n858), .Z(n860) );
  OR U1126 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .B(
        n867), .Z(n859) );
  AND U1127 ( .A(n860), .B(n859), .Z(n927) );
  ANDN U1128 ( .B(n883), .A(n1782), .Z(n878) );
  XNOR U1129 ( .A(n877), .B(n878), .Z(n880) );
  NANDN U1130 ( .A(n862), .B(n861), .Z(n866) );
  NANDN U1131 ( .A(n864), .B(n863), .Z(n865) );
  NAND U1132 ( .A(n866), .B(n865), .Z(n879) );
  XOR U1133 ( .A(n880), .B(n879), .Z(n872) );
  IV U1134 ( .A(n872), .Z(n887) );
  ANDN U1135 ( .B(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .A(n887), .Z(n875) );
  NANDN U1136 ( .A(n867), .B(\cin[0][2] ), .Z(n871) );
  NANDN U1137 ( .A(n915), .B(\cin[0][1] ), .Z(n869) );
  NANDN U1138 ( .A(n869), .B(n868), .Z(n870) );
  AND U1139 ( .A(n871), .B(n870), .Z(n884) );
  XOR U1140 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n872), .Z(n873) );
  NANDN U1141 ( .A(n884), .B(n873), .Z(n874) );
  NANDN U1142 ( .A(n875), .B(n874), .Z(n876) );
  AND U1143 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n876), .Z(n904) );
  NANDN U1144 ( .A(n878), .B(n877), .Z(n882) );
  NAND U1145 ( .A(n880), .B(n879), .Z(n881) );
  NAND U1146 ( .A(n882), .B(n881), .Z(n897) );
  ANDN U1147 ( .B(n883), .A(n1797), .Z(n899) );
  XNOR U1148 ( .A(n900), .B(n899), .Z(n898) );
  XOR U1149 ( .A(n897), .B(n898), .Z(n903) );
  XNOR U1150 ( .A(n904), .B(n903), .Z(n932) );
  NANDN U1151 ( .A(n1782), .B(n927), .Z(n890) );
  XNOR U1152 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[0].modmult_step_/z2[3] ), 
        .B(n884), .Z(n885) );
  NAND U1153 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n885), .Z(n886) );
  XOR U1154 ( .A(n887), .B(n886), .Z(n938) );
  NANDN U1155 ( .A(n927), .B(n1797), .Z(n888) );
  NANDN U1156 ( .A(n938), .B(n888), .Z(n889) );
  NAND U1157 ( .A(n890), .B(n889), .Z(n896) );
  XNOR U1158 ( .A(n891), .B(n915), .Z(n924) );
  NANDN U1159 ( .A(n[0]), .B(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n892) );
  NAND U1160 ( .A(n924), .B(n892), .Z(n893) );
  NANDN U1161 ( .A(n[1]), .B(n893), .Z(n894) );
  NANDN U1162 ( .A(n927), .B(n1782), .Z(n931) );
  NAND U1163 ( .A(n894), .B(n931), .Z(n895) );
  NANDN U1164 ( .A(n896), .B(n895), .Z(n909) );
  NAND U1165 ( .A(n898), .B(n897), .Z(n902) );
  ANDN U1166 ( .B(n900), .A(n899), .Z(n901) );
  ANDN U1167 ( .B(n902), .A(n901), .Z(n908) );
  AND U1168 ( .A(n904), .B(n903), .Z(n905) );
  XNOR U1169 ( .A(n906), .B(n905), .Z(n907) );
  XNOR U1170 ( .A(n908), .B(n907), .Z(n933) );
  ANDN U1171 ( .B(n909), .A(n933), .Z(n910) );
  AND U1172 ( .A(n932), .B(n910), .Z(n912) );
  NAND U1173 ( .A(n1797), .B(n938), .Z(n911) );
  NAND U1174 ( .A(n912), .B(n911), .Z(n925) );
  IV U1175 ( .A(n925), .Z(n936) );
  ANDN U1176 ( .B(n[0]), .A(
        \MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n921) );
  XNOR U1177 ( .A(n915), .B(n913), .Z(n914) );
  NANDN U1178 ( .A(n921), .B(n914), .Z(n918) );
  NAND U1179 ( .A(n921), .B(n915), .Z(n916) );
  NANDN U1180 ( .A(n[1]), .B(n916), .Z(n917) );
  AND U1181 ( .A(n918), .B(n917), .Z(n928) );
  XOR U1182 ( .A(n[2]), .B(n928), .Z(n919) );
  NANDN U1183 ( .A(n936), .B(n919), .Z(n920) );
  XNOR U1184 ( .A(n927), .B(n920), .Z(n943) );
  XOR U1185 ( .A(n[1]), .B(n921), .Z(n922) );
  NANDN U1186 ( .A(n936), .B(n922), .Z(n923) );
  XOR U1187 ( .A(n924), .B(n923), .Z(n942) );
  AND U1188 ( .A(n[0]), .B(n925), .Z(n926) );
  XNOR U1189 ( .A(\MODMULT1[0].modmult_1/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n926), .Z(n1134) );
  ANDN U1190 ( .B(n927), .A(n1782), .Z(n929) );
  OR U1191 ( .A(n929), .B(n928), .Z(n930) );
  AND U1192 ( .A(n931), .B(n930), .Z(n934) );
  XNOR U1193 ( .A(n1797), .B(n934), .Z(n935) );
  NANDN U1194 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U1195 ( .A(n938), .B(n937), .Z(n951) );
  ANDN U1196 ( .B(n[1]), .A(n947), .Z(n940) );
  ANDN U1197 ( .B(n[0]), .A(n947), .Z(n1133) );
  NAND U1198 ( .A(n1134), .B(n1133), .Z(n941) );
  XOR U1199 ( .A(n942), .B(n941), .Z(n939) );
  XNOR U1200 ( .A(n940), .B(n939), .Z(n1215) );
  NAND U1201 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1215), .Z(n1107) );
  XNOR U1202 ( .A(n943), .B(n944), .Z(n974) );
  ANDN U1203 ( .B(n[2]), .A(n947), .Z(n973) );
  NAND U1204 ( .A(n974), .B(n973), .Z(n946) );
  NANDN U1205 ( .A(n944), .B(n943), .Z(n945) );
  AND U1206 ( .A(n946), .B(n945), .Z(n949) );
  OR U1207 ( .A(n947), .B(n1797), .Z(n948) );
  XNOR U1208 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1209 ( .A(n951), .B(n950), .Z(n1230) );
  NAND U1210 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1230), .Z(n956) );
  AND U1211 ( .A(m[3]), .B(n1230), .Z(n972) );
  AND U1212 ( .A(m[1]), .B(n1230), .Z(n960) );
  AND U1213 ( .A(m[2]), .B(n1230), .Z(n963) );
  XNOR U1214 ( .A(n1797), .B(n970), .Z(n952) );
  NANDN U1215 ( .A(n972), .B(n952), .Z(n954) );
  NANDN U1216 ( .A(n1797), .B(n970), .Z(n953) );
  NAND U1217 ( .A(n954), .B(n953), .Z(n968) );
  NANDN U1218 ( .A(n968), .B(n[0]), .Z(n955) );
  XNOR U1219 ( .A(n956), .B(n955), .Z(n976) );
  NAND U1220 ( .A(n[0]), .B(n956), .Z(n959) );
  XNOR U1221 ( .A(n[1]), .B(n959), .Z(n957) );
  NANDN U1222 ( .A(n968), .B(n957), .Z(n958) );
  XNOR U1223 ( .A(n960), .B(n958), .Z(n980) );
  XNOR U1224 ( .A(n1782), .B(n964), .Z(n962) );
  NANDN U1225 ( .A(n968), .B(n962), .Z(n961) );
  XOR U1226 ( .A(n963), .B(n961), .Z(n979) );
  IV U1227 ( .A(n979), .Z(n992) );
  NANDN U1228 ( .A(n963), .B(n962), .Z(n966) );
  NANDN U1229 ( .A(n1782), .B(n964), .Z(n965) );
  AND U1230 ( .A(n966), .B(n965), .Z(n971) );
  XOR U1231 ( .A(n1797), .B(n971), .Z(n967) );
  NANDN U1232 ( .A(n968), .B(n967), .Z(n969) );
  AND U1233 ( .A(n972), .B(n969), .Z(n1007) );
  ANDN U1234 ( .B(n[0]), .A(n1005), .Z(n975) );
  AND U1235 ( .A(n976), .B(n975), .Z(n983) );
  ANDN U1236 ( .B(n[1]), .A(n1005), .Z(n981) );
  IV U1237 ( .A(n987), .Z(n986) );
  XNOR U1238 ( .A(n974), .B(n973), .Z(n1220) );
  XOR U1239 ( .A(n976), .B(n975), .Z(n1015) );
  ANDN U1240 ( .B(m[1]), .A(n1015), .Z(n989) );
  XOR U1241 ( .A(m[2]), .B(n989), .Z(n977) );
  NAND U1242 ( .A(n1220), .B(n977), .Z(n978) );
  XOR U1243 ( .A(n986), .B(n978), .Z(n1029) );
  NOR U1244 ( .A(n1782), .B(n1005), .Z(n993) );
  XOR U1245 ( .A(n979), .B(n993), .Z(n995) );
  NANDN U1246 ( .A(n981), .B(n980), .Z(n985) );
  NANDN U1247 ( .A(n983), .B(n982), .Z(n984) );
  NAND U1248 ( .A(n985), .B(n984), .Z(n994) );
  XOR U1249 ( .A(n995), .B(n994), .Z(n999) );
  IV U1250 ( .A(n999), .Z(n998) );
  NANDN U1251 ( .A(n986), .B(m[2]), .Z(n991) );
  XOR U1252 ( .A(m[2]), .B(n987), .Z(n988) );
  NAND U1253 ( .A(n989), .B(n988), .Z(n990) );
  AND U1254 ( .A(n991), .B(n990), .Z(n1000) );
  AND U1255 ( .A(n1051), .B(n1797), .Z(n1036) );
  NANDN U1256 ( .A(n993), .B(n992), .Z(n997) );
  NAND U1257 ( .A(n995), .B(n994), .Z(n996) );
  AND U1258 ( .A(n997), .B(n996), .Z(n1011) );
  ANDN U1259 ( .B(m[3]), .A(n998), .Z(n1003) );
  XOR U1260 ( .A(m[3]), .B(n999), .Z(n1001) );
  ANDN U1261 ( .B(n1001), .A(n1000), .Z(n1002) );
  OR U1262 ( .A(n1003), .B(n1002), .Z(n1004) );
  AND U1263 ( .A(n1220), .B(n1004), .Z(n1013) );
  XOR U1264 ( .A(n1011), .B(n1013), .Z(n1009) );
  OR U1265 ( .A(n1005), .B(n1797), .Z(n1006) );
  AND U1266 ( .A(n1007), .B(n1006), .Z(n1010) );
  XNOR U1267 ( .A(n1013), .B(n1010), .Z(n1008) );
  NAND U1268 ( .A(n1009), .B(n1008), .Z(n1046) );
  XNOR U1269 ( .A(n1011), .B(n1010), .Z(n1012) );
  XNOR U1270 ( .A(n1013), .B(n1012), .Z(n1045) );
  ANDN U1271 ( .B(n1046), .A(n1045), .Z(n1022) );
  OR U1272 ( .A(n1029), .B(n1782), .Z(n1040) );
  NOR U1273 ( .A(n1797), .B(n1051), .Z(n1041) );
  ANDN U1274 ( .B(n1040), .A(n1041), .Z(n1020) );
  NAND U1275 ( .A(n1220), .B(m[1]), .Z(n1014) );
  XOR U1276 ( .A(n1015), .B(n1014), .Z(n1033) );
  NANDN U1277 ( .A(n1033), .B(n[1]), .Z(n1026) );
  NAND U1278 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1220), .Z(n1035) );
  NOR U1279 ( .A(n1035), .B(n[0]), .Z(n1016) );
  NAND U1280 ( .A(n1026), .B(n1016), .Z(n1017) );
  NANDN U1281 ( .A(n1024), .B(n1017), .Z(n1018) );
  AND U1282 ( .A(n1029), .B(n1782), .Z(n1038) );
  OR U1283 ( .A(n1018), .B(n1038), .Z(n1019) );
  AND U1284 ( .A(n1020), .B(n1019), .Z(n1021) );
  ANDN U1285 ( .B(n1022), .A(n1021), .Z(n1023) );
  NANDN U1286 ( .A(n1036), .B(n1023), .Z(n1049) );
  AND U1287 ( .A(n[0]), .B(n1035), .Z(n1030) );
  NANDN U1288 ( .A(n1024), .B(n1030), .Z(n1025) );
  AND U1289 ( .A(n1026), .B(n1025), .Z(n1037) );
  XOR U1290 ( .A(n1782), .B(n1037), .Z(n1027) );
  NAND U1291 ( .A(n1049), .B(n1027), .Z(n1028) );
  XNOR U1292 ( .A(n1029), .B(n1028), .Z(n1072) );
  XOR U1293 ( .A(n[1]), .B(n1030), .Z(n1031) );
  NAND U1294 ( .A(n1049), .B(n1031), .Z(n1032) );
  XOR U1295 ( .A(n1033), .B(n1032), .Z(n1053) );
  NAND U1296 ( .A(n1049), .B(n[0]), .Z(n1034) );
  XOR U1297 ( .A(n1035), .B(n1034), .Z(n1059) );
  ANDN U1298 ( .B(n1049), .A(n1036), .Z(n1043) );
  OR U1299 ( .A(n1038), .B(n1037), .Z(n1039) );
  AND U1300 ( .A(n1040), .B(n1039), .Z(n1047) );
  NANDN U1301 ( .A(n1041), .B(n1047), .Z(n1042) );
  AND U1302 ( .A(n1043), .B(n1042), .Z(n1044) );
  XNOR U1303 ( .A(n1045), .B(n1044), .Z(n1088) );
  XOR U1304 ( .A(n1797), .B(n1047), .Z(n1048) );
  NAND U1305 ( .A(n1049), .B(n1048), .Z(n1050) );
  XNOR U1306 ( .A(n1051), .B(n1050), .Z(n1080) );
  ANDN U1307 ( .B(n1078), .A(n1782), .Z(n1073) );
  XNOR U1308 ( .A(n1072), .B(n1073), .Z(n1075) );
  NAND U1309 ( .A(n[1]), .B(n1078), .Z(n1052) );
  NANDN U1310 ( .A(n1053), .B(n1052), .Z(n1055) );
  AND U1311 ( .A(n[0]), .B(n1078), .Z(n1058) );
  ANDN U1312 ( .B(n1058), .A(n1059), .Z(n1057) );
  XNOR U1313 ( .A(n1053), .B(n1052), .Z(n1056) );
  NANDN U1314 ( .A(n1057), .B(n1056), .Z(n1054) );
  NAND U1315 ( .A(n1055), .B(n1054), .Z(n1074) );
  XOR U1316 ( .A(n1075), .B(n1074), .Z(n1066) );
  IV U1317 ( .A(n1066), .Z(n1065) );
  XOR U1318 ( .A(n1057), .B(n1056), .Z(n1095) );
  NANDN U1319 ( .A(n1095), .B(m[2]), .Z(n1062) );
  XNOR U1320 ( .A(m[2]), .B(n1095), .Z(n1060) );
  XOR U1321 ( .A(n1059), .B(n1058), .Z(n1098) );
  AND U1322 ( .A(m[1]), .B(n1098), .Z(n1092) );
  NAND U1323 ( .A(n1060), .B(n1092), .Z(n1061) );
  NAND U1324 ( .A(n1062), .B(n1061), .Z(n1067) );
  XOR U1325 ( .A(m[3]), .B(n1067), .Z(n1063) );
  NAND U1326 ( .A(n1215), .B(n1063), .Z(n1064) );
  XOR U1327 ( .A(n1065), .B(n1064), .Z(n1120) );
  AND U1328 ( .A(n1120), .B(n1797), .Z(n1106) );
  ANDN U1329 ( .B(m[3]), .A(n1065), .Z(n1070) );
  XOR U1330 ( .A(m[3]), .B(n1066), .Z(n1068) );
  AND U1331 ( .A(n1068), .B(n1067), .Z(n1069) );
  OR U1332 ( .A(n1070), .B(n1069), .Z(n1071) );
  AND U1333 ( .A(n1215), .B(n1071), .Z(n1086) );
  NANDN U1334 ( .A(n1073), .B(n1072), .Z(n1077) );
  NAND U1335 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U1336 ( .A(n1077), .B(n1076), .Z(n1081) );
  NANDN U1337 ( .A(n1797), .B(n1078), .Z(n1079) );
  XOR U1338 ( .A(n1080), .B(n1079), .Z(n1082) );
  XNOR U1339 ( .A(n1081), .B(n1082), .Z(n1085) );
  NOR U1340 ( .A(n1106), .B(n1115), .Z(n1091) );
  AND U1341 ( .A(n1080), .B(n1079), .Z(n1084) );
  AND U1342 ( .A(n1082), .B(n1081), .Z(n1083) );
  NOR U1343 ( .A(n1084), .B(n1083), .Z(n1090) );
  ANDN U1344 ( .B(n1086), .A(n1085), .Z(n1087) );
  XOR U1345 ( .A(n1088), .B(n1087), .Z(n1089) );
  XNOR U1346 ( .A(n1090), .B(n1089), .Z(n1116) );
  ANDN U1347 ( .B(n1091), .A(n1116), .Z(n1104) );
  NOR U1348 ( .A(n1797), .B(n1120), .Z(n1111) );
  XOR U1349 ( .A(n1092), .B(m[2]), .Z(n1093) );
  NAND U1350 ( .A(n1215), .B(n1093), .Z(n1094) );
  XNOR U1351 ( .A(n1095), .B(n1094), .Z(n1127) );
  ANDN U1352 ( .B(n1127), .A(n1782), .Z(n1108) );
  NOR U1353 ( .A(n1111), .B(n1108), .Z(n1102) );
  OR U1354 ( .A(n[0]), .B(n1107), .Z(n1096) );
  NAND U1355 ( .A(n[1]), .B(n1096), .Z(n1099) );
  NAND U1356 ( .A(m[1]), .B(n1215), .Z(n1097) );
  XOR U1357 ( .A(n1098), .B(n1097), .Z(n1132) );
  ANDN U1358 ( .B(n1099), .A(n1132), .Z(n1100) );
  ANDN U1359 ( .B(n1782), .A(n1127), .Z(n1109) );
  OR U1360 ( .A(n1100), .B(n1109), .Z(n1101) );
  AND U1361 ( .A(n1102), .B(n1101), .Z(n1103) );
  ANDN U1362 ( .B(n1104), .A(n1103), .Z(n1130) );
  NANDN U1363 ( .A(n1130), .B(n[0]), .Z(n1105) );
  XNOR U1364 ( .A(n1107), .B(n1105), .Z(n1136) );
  IV U1365 ( .A(n1130), .Z(n1125) );
  ANDN U1366 ( .B(n1125), .A(n1106), .Z(n1113) );
  NAND U1367 ( .A(n[0]), .B(n1107), .Z(n1128) );
  OR U1368 ( .A(n1108), .B(n1123), .Z(n1110) );
  ANDN U1369 ( .B(n1110), .A(n1109), .Z(n1117) );
  OR U1370 ( .A(n1111), .B(n1117), .Z(n1112) );
  NAND U1371 ( .A(n1113), .B(n1112), .Z(n1114) );
  XNOR U1372 ( .A(n1115), .B(n1114), .Z(n1177) );
  NOR U1373 ( .A(n1177), .B(n1116), .Z(n1122) );
  XNOR U1374 ( .A(n1797), .B(n1117), .Z(n1118) );
  NANDN U1375 ( .A(n1130), .B(n1118), .Z(n1119) );
  XNOR U1376 ( .A(n1120), .B(n1119), .Z(n1163) );
  NAND U1377 ( .A(n1797), .B(n1163), .Z(n1121) );
  NAND U1378 ( .A(n1122), .B(n1121), .Z(n1139) );
  XNOR U1379 ( .A(n1782), .B(n1123), .Z(n1124) );
  NAND U1380 ( .A(n1125), .B(n1124), .Z(n1126) );
  XNOR U1381 ( .A(n1127), .B(n1126), .Z(n1141) );
  XNOR U1382 ( .A(n[1]), .B(n1128), .Z(n1129) );
  NANDN U1383 ( .A(n1130), .B(n1129), .Z(n1131) );
  XNOR U1384 ( .A(n1132), .B(n1131), .Z(n1145) );
  NANDN U1385 ( .A(n1782), .B(n1141), .Z(n1140) );
  AND U1386 ( .A(n[0]), .B(n1162), .Z(n1135) );
  AND U1387 ( .A(n1136), .B(n1135), .Z(n1147) );
  NAND U1388 ( .A(n1162), .B(n[1]), .Z(n1144) );
  XNOR U1389 ( .A(n1145), .B(n1144), .Z(n1146) );
  XOR U1390 ( .A(n1147), .B(n1146), .Z(n1150) );
  XNOR U1391 ( .A(n1134), .B(n1133), .Z(n1206) );
  XNOR U1392 ( .A(n1136), .B(n1135), .Z(n1181) );
  AND U1393 ( .A(m[1]), .B(n1181), .Z(n1152) );
  XOR U1394 ( .A(n1152), .B(m[2]), .Z(n1137) );
  NAND U1395 ( .A(n1206), .B(n1137), .Z(n1138) );
  XNOR U1396 ( .A(n1150), .B(n1138), .Z(n1189) );
  NANDN U1397 ( .A(n1140), .B(n1139), .Z(n1143) );
  NAND U1398 ( .A(n[2]), .B(n1162), .Z(n1142) );
  ANDN U1399 ( .B(n1142), .A(n1141), .Z(n1160) );
  ANDN U1400 ( .B(n1143), .A(n1160), .Z(n1158) );
  NANDN U1401 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1402 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1403 ( .A(n1149), .B(n1148), .Z(n1159) );
  IV U1404 ( .A(n1168), .Z(n1167) );
  NANDN U1405 ( .A(n1150), .B(m[2]), .Z(n1154) );
  XNOR U1406 ( .A(m[2]), .B(n1150), .Z(n1151) );
  NAND U1407 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1408 ( .A(n1154), .B(n1153), .Z(n1169) );
  IV U1409 ( .A(n1169), .Z(n1155) );
  XOR U1410 ( .A(m[3]), .B(n1155), .Z(n1156) );
  NAND U1411 ( .A(n1206), .B(n1156), .Z(n1157) );
  XOR U1412 ( .A(n1167), .B(n1157), .Z(n1204) );
  NANDN U1413 ( .A(n1159), .B(n1158), .Z(n1161) );
  ANDN U1414 ( .B(n1161), .A(n1160), .Z(n1175) );
  AND U1415 ( .A(n1162), .B(n[3]), .Z(n1164) );
  XNOR U1416 ( .A(n1163), .B(n1164), .Z(n1174) );
  NANDN U1417 ( .A(n1175), .B(n1174), .Z(n1166) );
  NANDN U1418 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1419 ( .A(n1166), .B(n1165), .Z(n1179) );
  ANDN U1420 ( .B(m[3]), .A(n1167), .Z(n1172) );
  XOR U1421 ( .A(m[3]), .B(n1168), .Z(n1170) );
  ANDN U1422 ( .B(n1170), .A(n1169), .Z(n1171) );
  OR U1423 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U1424 ( .A(n1206), .B(n1173), .Z(n1183) );
  XNOR U1425 ( .A(n1175), .B(n1174), .Z(n1182) );
  AND U1426 ( .A(n1183), .B(n1182), .Z(n1176) );
  XNOR U1427 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1428 ( .A(n1179), .B(n1178), .Z(n1199) );
  NAND U1429 ( .A(n1206), .B(m[1]), .Z(n1180) );
  XOR U1430 ( .A(n1181), .B(n1180), .Z(n1191) );
  NOR U1431 ( .A(n1191), .B(n[1]), .Z(n1184) );
  NAND U1432 ( .A(n[1]), .B(n1191), .Z(n1186) );
  AND U1433 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1206), .Z(n1193) );
  ANDN U1434 ( .B(n1782), .A(n1189), .Z(n1196) );
  ANDN U1435 ( .B(n1189), .A(n1782), .Z(n1195) );
  XNOR U1436 ( .A(n1183), .B(n1182), .Z(n1198) );
  NANDN U1437 ( .A(n1193), .B(n[0]), .Z(n1190) );
  OR U1438 ( .A(n1184), .B(n1190), .Z(n1185) );
  AND U1439 ( .A(n1186), .B(n1185), .Z(n1194) );
  XOR U1440 ( .A(n1782), .B(n1194), .Z(n1187) );
  NANDN U1441 ( .A(n1202), .B(n1187), .Z(n1188) );
  XNOR U1442 ( .A(n1189), .B(n1188), .Z(n1236) );
  NANDN U1443 ( .A(n1202), .B(n[0]), .Z(n1192) );
  XOR U1444 ( .A(n1193), .B(n1192), .Z(n1212) );
  NANDN U1445 ( .A(n1195), .B(n1194), .Z(n1197) );
  ANDN U1446 ( .B(n1197), .A(n1196), .Z(n1200) );
  XNOR U1447 ( .A(n1797), .B(n1200), .Z(n1201) );
  NANDN U1448 ( .A(n1202), .B(n1201), .Z(n1203) );
  XNOR U1449 ( .A(n1204), .B(n1203), .Z(n1244) );
  ANDN U1450 ( .B(n[0]), .A(n1240), .Z(n1211) );
  XNOR U1451 ( .A(n1211), .B(n1212), .Z(n1205) );
  NANDN U1452 ( .A(n1227), .B(n1205), .Z(n1210) );
  ANDN U1453 ( .B(\keep_1[0] ), .A(n1246), .Z(n1231) );
  NAND U1454 ( .A(n1231), .B(n1206), .Z(n1208) );
  NANDN U1455 ( .A(\keep_1[0] ), .B(
        \MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1207)
         );
  NAND U1456 ( .A(n1208), .B(n1207), .Z(n1209) );
  ANDN U1457 ( .B(n1210), .A(n1209), .Z(n1468) );
  IV U1458 ( .A(n1468), .Z(n1483) );
  ANDN U1459 ( .B(n[1]), .A(n1240), .Z(n1223) );
  XOR U1460 ( .A(n1224), .B(n1223), .Z(n1213) );
  XNOR U1461 ( .A(n1213), .B(n1225), .Z(n1214) );
  NANDN U1462 ( .A(n1227), .B(n1214), .Z(n1219) );
  NAND U1463 ( .A(n1231), .B(n1215), .Z(n1217) );
  NANDN U1464 ( .A(\keep_1[0] ), .B(m[1]), .Z(n1216) );
  NAND U1465 ( .A(n1217), .B(n1216), .Z(n1218) );
  ANDN U1466 ( .B(n1219), .A(n1218), .Z(n1464) );
  IV U1467 ( .A(n1464), .Z(n1344) );
  NAND U1468 ( .A(n1231), .B(n1220), .Z(n1222) );
  NANDN U1469 ( .A(\keep_1[0] ), .B(m[2]), .Z(n1221) );
  NAND U1470 ( .A(n1222), .B(n1221), .Z(n1229) );
  NOR U1471 ( .A(n1782), .B(n1240), .Z(n1235) );
  XNOR U1472 ( .A(n1236), .B(n1237), .Z(n1234) );
  XNOR U1473 ( .A(n1235), .B(n1234), .Z(n1226) );
  NANDN U1474 ( .A(n1227), .B(n1226), .Z(n1228) );
  NANDN U1475 ( .A(n1229), .B(n1228), .Z(n1445) );
  AND U1476 ( .A(n1445), .B(n1483), .Z(n1317) );
  NAND U1477 ( .A(n1231), .B(n1230), .Z(n1233) );
  NANDN U1478 ( .A(\keep_1[0] ), .B(m[3]), .Z(n1232) );
  AND U1479 ( .A(n1233), .B(n1232), .Z(n1248) );
  NAND U1480 ( .A(n1235), .B(n1234), .Z(n1239) );
  NANDN U1481 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1482 ( .A(n1239), .B(n1238), .Z(n1242) );
  OR U1483 ( .A(n1240), .B(n1797), .Z(n1241) );
  XNOR U1484 ( .A(n1242), .B(n1241), .Z(n1243) );
  XNOR U1485 ( .A(n1244), .B(n1243), .Z(n1245) );
  NAND U1486 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U1487 ( .A(n1248), .B(n1247), .Z(n1440) );
  IV U1488 ( .A(n1440), .Z(n1457) );
  AND U1489 ( .A(n1445), .B(n1457), .Z(n1267) );
  NAND U1490 ( .A(n1267), .B(n1782), .Z(n1250) );
  AND U1491 ( .A(n1457), .B(n1797), .Z(n1249) );
  ANDN U1492 ( .B(n1250), .A(n1249), .Z(n1258) );
  ANDN U1493 ( .B(n1457), .A(n1464), .Z(n1262) );
  NANDN U1494 ( .A(n1262), .B(n[1]), .Z(n1254) );
  NANDN U1495 ( .A(n[1]), .B(n1262), .Z(n1252) );
  NANDN U1496 ( .A(n1468), .B(n1457), .Z(n1264) );
  OR U1497 ( .A(n1264), .B(n[0]), .Z(n1251) );
  NAND U1498 ( .A(n1252), .B(n1251), .Z(n1253) );
  NAND U1499 ( .A(n1254), .B(n1253), .Z(n1256) );
  XNOR U1500 ( .A(n1267), .B(n[2]), .Z(n1255) );
  NANDN U1501 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U1502 ( .A(n1258), .B(n1257), .Z(n1272) );
  NAND U1503 ( .A(n[0]), .B(n1264), .Z(n1259) );
  XNOR U1504 ( .A(n1265), .B(n1782), .Z(n1266) );
  XNOR U1505 ( .A(n[1]), .B(n1259), .Z(n1260) );
  NAND U1506 ( .A(n1272), .B(n1260), .Z(n1261) );
  XNOR U1507 ( .A(n1262), .B(n1261), .Z(n1275) );
  NAND U1508 ( .A(n1272), .B(n[0]), .Z(n1263) );
  XNOR U1509 ( .A(n1264), .B(n1263), .Z(n1279) );
  NANDN U1510 ( .A(n1782), .B(n1265), .Z(n1269) );
  NANDN U1511 ( .A(n1267), .B(n1266), .Z(n1268) );
  NAND U1512 ( .A(n1269), .B(n1268), .Z(n1270) );
  XNOR U1513 ( .A(n1270), .B(n1797), .Z(n1271) );
  NAND U1514 ( .A(n1272), .B(n1271), .Z(n1273) );
  ANDN U1515 ( .B(n1273), .A(n1440), .Z(n1292) );
  NOR U1516 ( .A(n1782), .B(n1290), .Z(n1294) );
  XNOR U1517 ( .A(n1293), .B(n1294), .Z(n1296) );
  ANDN U1518 ( .B(n[1]), .A(n1290), .Z(n1274) );
  NANDN U1519 ( .A(n1274), .B(n1275), .Z(n1277) );
  ANDN U1520 ( .B(n[0]), .A(n1290), .Z(n1278) );
  AND U1521 ( .A(n1279), .B(n1278), .Z(n1281) );
  XNOR U1522 ( .A(n1275), .B(n1274), .Z(n1280) );
  NANDN U1523 ( .A(n1281), .B(n1280), .Z(n1276) );
  NAND U1524 ( .A(n1277), .B(n1276), .Z(n1295) );
  XOR U1525 ( .A(n1296), .B(n1295), .Z(n1288) );
  XOR U1526 ( .A(n1279), .B(n1278), .Z(n1307) );
  NANDN U1527 ( .A(n1307), .B(n1344), .Z(n1303) );
  XOR U1528 ( .A(n1281), .B(n1280), .Z(n1305) );
  AND U1529 ( .A(n1303), .B(n1305), .Z(n1286) );
  IV U1530 ( .A(n1286), .Z(n1282) );
  XNOR U1531 ( .A(n1282), .B(n1440), .Z(n1283) );
  NAND U1532 ( .A(n1445), .B(n1283), .Z(n1284) );
  XOR U1533 ( .A(n1288), .B(n1284), .Z(n1334) );
  ANDN U1534 ( .B(n1797), .A(n1334), .Z(n1335) );
  XOR U1535 ( .A(n1457), .B(n1288), .Z(n1285) );
  NANDN U1536 ( .A(n1286), .B(n1285), .Z(n1287) );
  NANDN U1537 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U1538 ( .A(n1289), .B(n1445), .Z(n1302) );
  OR U1539 ( .A(n1290), .B(n1797), .Z(n1291) );
  NAND U1540 ( .A(n1292), .B(n1291), .Z(n1299) );
  NANDN U1541 ( .A(n1294), .B(n1293), .Z(n1298) );
  NAND U1542 ( .A(n1296), .B(n1295), .Z(n1297) );
  AND U1543 ( .A(n1298), .B(n1297), .Z(n1300) );
  XOR U1544 ( .A(n1300), .B(n1299), .Z(n1301) );
  XNOR U1545 ( .A(n1302), .B(n1301), .Z(n1342) );
  ANDN U1546 ( .B(n1343), .A(n1342), .Z(n1314) );
  ANDN U1547 ( .B(n1334), .A(n1797), .Z(n1338) );
  NAND U1548 ( .A(n1445), .B(n1303), .Z(n1304) );
  XOR U1549 ( .A(n1305), .B(n1304), .Z(n1327) );
  NOR U1550 ( .A(n1782), .B(n1327), .Z(n1329) );
  NOR U1551 ( .A(n1338), .B(n1329), .Z(n1312) );
  NANDN U1552 ( .A(n1464), .B(n1445), .Z(n1306) );
  XOR U1553 ( .A(n1307), .B(n1306), .Z(n1320) );
  NANDN U1554 ( .A(n1320), .B(n[1]), .Z(n1324) );
  ANDN U1555 ( .B(n1317), .A(n[0]), .Z(n1308) );
  NAND U1556 ( .A(n1324), .B(n1308), .Z(n1309) );
  NANDN U1557 ( .A(n1322), .B(n1309), .Z(n1310) );
  AND U1558 ( .A(n1327), .B(n1782), .Z(n1330) );
  OR U1559 ( .A(n1310), .B(n1330), .Z(n1311) );
  AND U1560 ( .A(n1312), .B(n1311), .Z(n1313) );
  ANDN U1561 ( .B(n1314), .A(n1313), .Z(n1315) );
  NANDN U1562 ( .A(n1335), .B(n1315), .Z(n1336) );
  NAND U1563 ( .A(n1336), .B(n[0]), .Z(n1316) );
  XOR U1564 ( .A(n1317), .B(n1316), .Z(n1346) );
  ANDN U1565 ( .B(n[0]), .A(n1317), .Z(n1321) );
  XOR U1566 ( .A(n[1]), .B(n1321), .Z(n1318) );
  NAND U1567 ( .A(n1336), .B(n1318), .Z(n1319) );
  XOR U1568 ( .A(n1320), .B(n1319), .Z(n1348) );
  NANDN U1569 ( .A(n1322), .B(n1321), .Z(n1323) );
  AND U1570 ( .A(n1324), .B(n1323), .Z(n1328) );
  XOR U1571 ( .A(n1782), .B(n1328), .Z(n1325) );
  AND U1572 ( .A(n1336), .B(n1325), .Z(n1326) );
  XOR U1573 ( .A(n1327), .B(n1326), .Z(n1361) );
  NANDN U1574 ( .A(n1329), .B(n1328), .Z(n1331) );
  ANDN U1575 ( .B(n1331), .A(n1330), .Z(n1337) );
  XNOR U1576 ( .A(n1797), .B(n1337), .Z(n1332) );
  NAND U1577 ( .A(n1336), .B(n1332), .Z(n1333) );
  XNOR U1578 ( .A(n1334), .B(n1333), .Z(n1371) );
  ANDN U1579 ( .B(n1336), .A(n1335), .Z(n1340) );
  OR U1580 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U1581 ( .A(n1340), .B(n1339), .Z(n1341) );
  XOR U1582 ( .A(n1342), .B(n1341), .Z(n1377) );
  AND U1583 ( .A(n[0]), .B(n1367), .Z(n1345) );
  XOR U1584 ( .A(n1346), .B(n1345), .Z(n1381) );
  XOR U1585 ( .A(n1344), .B(n1381), .Z(n1394) );
  NOR U1586 ( .A(n1464), .B(n1468), .Z(n1403) );
  ANDN U1587 ( .B(n[0]), .A(n1403), .Z(n1395) );
  XOR U1588 ( .A(n[1]), .B(n1395), .Z(n1392) );
  ANDN U1589 ( .B(n1367), .A(n1782), .Z(n1362) );
  XNOR U1590 ( .A(n1361), .B(n1362), .Z(n1364) );
  NAND U1591 ( .A(n[1]), .B(n1367), .Z(n1347) );
  NANDN U1592 ( .A(n1348), .B(n1347), .Z(n1350) );
  NAND U1593 ( .A(n1346), .B(n1345), .Z(n1352) );
  XNOR U1594 ( .A(n1348), .B(n1347), .Z(n1351) );
  NAND U1595 ( .A(n1352), .B(n1351), .Z(n1349) );
  NAND U1596 ( .A(n1350), .B(n1349), .Z(n1363) );
  XOR U1597 ( .A(n1364), .B(n1363), .Z(n1355) );
  XOR U1598 ( .A(n1352), .B(n1351), .Z(n1384) );
  XNOR U1599 ( .A(n1356), .B(n1440), .Z(n1353) );
  NANDN U1600 ( .A(n1464), .B(n1353), .Z(n1354) );
  XOR U1601 ( .A(n1355), .B(n1354), .Z(n1410) );
  ANDN U1602 ( .B(n1797), .A(n1410), .Z(n1412) );
  ANDN U1603 ( .B(n1355), .A(n1440), .Z(n1359) );
  XOR U1604 ( .A(n1457), .B(n1355), .Z(n1357) );
  AND U1605 ( .A(n1357), .B(n1356), .Z(n1358) );
  OR U1606 ( .A(n1359), .B(n1358), .Z(n1360) );
  ANDN U1607 ( .B(n1360), .A(n1464), .Z(n1375) );
  NANDN U1608 ( .A(n1362), .B(n1361), .Z(n1366) );
  NAND U1609 ( .A(n1364), .B(n1363), .Z(n1365) );
  NAND U1610 ( .A(n1366), .B(n1365), .Z(n1368) );
  ANDN U1611 ( .B(n1367), .A(n1797), .Z(n1370) );
  XNOR U1612 ( .A(n1371), .B(n1370), .Z(n1369) );
  XNOR U1613 ( .A(n1375), .B(n1374), .Z(n1415) );
  NOR U1614 ( .A(n1412), .B(n1415), .Z(n1380) );
  NANDN U1615 ( .A(n1369), .B(n1368), .Z(n1373) );
  OR U1616 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U1617 ( .A(n1373), .B(n1372), .Z(n1379) );
  ANDN U1618 ( .B(n1375), .A(n1374), .Z(n1376) );
  XNOR U1619 ( .A(n1377), .B(n1376), .Z(n1378) );
  XNOR U1620 ( .A(n1379), .B(n1378), .Z(n1416) );
  ANDN U1621 ( .B(n1380), .A(n1416), .Z(n1391) );
  ANDN U1622 ( .B(n1410), .A(n1797), .Z(n1414) );
  XNOR U1623 ( .A(n1381), .B(n1445), .Z(n1382) );
  NANDN U1624 ( .A(n1464), .B(n1382), .Z(n1383) );
  XOR U1625 ( .A(n1384), .B(n1383), .Z(n1401) );
  ANDN U1626 ( .B(n1401), .A(n1782), .Z(n1405) );
  NOR U1627 ( .A(n1414), .B(n1405), .Z(n1389) );
  NOR U1628 ( .A(n1394), .B(n[1]), .Z(n1397) );
  IV U1629 ( .A(n1403), .Z(n1484) );
  NOR U1630 ( .A(n1484), .B(n[0]), .Z(n1385) );
  NANDN U1631 ( .A(n1396), .B(n1385), .Z(n1386) );
  NANDN U1632 ( .A(n1397), .B(n1386), .Z(n1387) );
  ANDN U1633 ( .B(n1782), .A(n1401), .Z(n1406) );
  OR U1634 ( .A(n1387), .B(n1406), .Z(n1388) );
  AND U1635 ( .A(n1389), .B(n1388), .Z(n1390) );
  ANDN U1636 ( .B(n1391), .A(n1390), .Z(n1411) );
  ANDN U1637 ( .B(n1392), .A(n1411), .Z(n1393) );
  XOR U1638 ( .A(n1394), .B(n1393), .Z(n1420) );
  OR U1639 ( .A(n1396), .B(n1395), .Z(n1398) );
  ANDN U1640 ( .B(n1398), .A(n1397), .Z(n1404) );
  XNOR U1641 ( .A(n1782), .B(n1404), .Z(n1399) );
  NANDN U1642 ( .A(n1411), .B(n1399), .Z(n1400) );
  XNOR U1643 ( .A(n1401), .B(n1400), .Z(n1426) );
  NANDN U1644 ( .A(n1411), .B(n[0]), .Z(n1402) );
  XOR U1645 ( .A(n1403), .B(n1402), .Z(n1444) );
  NANDN U1646 ( .A(n1782), .B(n1426), .Z(n1424) );
  OR U1647 ( .A(n1405), .B(n1404), .Z(n1407) );
  ANDN U1648 ( .B(n1407), .A(n1406), .Z(n1413) );
  XNOR U1649 ( .A(n1797), .B(n1413), .Z(n1408) );
  NANDN U1650 ( .A(n1411), .B(n1408), .Z(n1409) );
  XNOR U1651 ( .A(n1410), .B(n1409), .Z(n1433) );
  NOR U1652 ( .A(n1454), .B(n1416), .Z(n1418) );
  NANDN U1653 ( .A(n1433), .B(n1797), .Z(n1417) );
  NAND U1654 ( .A(n1418), .B(n1417), .Z(n1423) );
  NANDN U1655 ( .A(n1425), .B(n[1]), .Z(n1419) );
  NANDN U1656 ( .A(n1420), .B(n1419), .Z(n1422) );
  XOR U1657 ( .A(n1420), .B(n1419), .Z(n1441) );
  ANDN U1658 ( .B(n[0]), .A(n1425), .Z(n1443) );
  NAND U1659 ( .A(n1444), .B(n1443), .Z(n1442) );
  NANDN U1660 ( .A(n1441), .B(n1442), .Z(n1421) );
  AND U1661 ( .A(n1422), .B(n1421), .Z(n1438) );
  NANDN U1662 ( .A(n1424), .B(n1423), .Z(n1428) );
  IV U1663 ( .A(n1425), .Z(n1431) );
  NAND U1664 ( .A(n1431), .B(n[2]), .Z(n1427) );
  ANDN U1665 ( .B(n1427), .A(n1426), .Z(n1429) );
  ANDN U1666 ( .B(n1428), .A(n1429), .Z(n1439) );
  NANDN U1667 ( .A(n1438), .B(n1439), .Z(n1430) );
  ANDN U1668 ( .B(n1430), .A(n1429), .Z(n1436) );
  NANDN U1669 ( .A(n1797), .B(n1431), .Z(n1432) );
  XNOR U1670 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1671 ( .A(n1436), .B(n1437), .Z(n1435) );
  NANDN U1672 ( .A(n1433), .B(n1432), .Z(n1434) );
  AND U1673 ( .A(n1435), .B(n1434), .Z(n1456) );
  XNOR U1674 ( .A(n1437), .B(n1436), .Z(n1479) );
  ANDN U1675 ( .B(n1461), .A(n1440), .Z(n1451) );
  XOR U1676 ( .A(n1457), .B(n1461), .Z(n1449) );
  XOR U1677 ( .A(n1442), .B(n1441), .Z(n1469) );
  NANDN U1678 ( .A(n1469), .B(n1445), .Z(n1448) );
  XOR U1679 ( .A(n1444), .B(n1443), .Z(n1487) );
  IV U1680 ( .A(n1487), .Z(n1485) );
  NANDN U1681 ( .A(n1464), .B(n1485), .Z(n1446) );
  XOR U1682 ( .A(n1445), .B(n1469), .Z(n1466) );
  OR U1683 ( .A(n1446), .B(n1466), .Z(n1447) );
  AND U1684 ( .A(n1448), .B(n1447), .Z(n1458) );
  ANDN U1685 ( .B(n1449), .A(n1458), .Z(n1450) );
  OR U1686 ( .A(n1451), .B(n1450), .Z(n1452) );
  ANDN U1687 ( .B(n1452), .A(n1468), .Z(n1478) );
  AND U1688 ( .A(n1479), .B(n1478), .Z(n1453) );
  XNOR U1689 ( .A(n1454), .B(n1453), .Z(n1455) );
  XNOR U1690 ( .A(n1456), .B(n1455), .Z(n1498) );
  XNOR U1691 ( .A(n1458), .B(n1457), .Z(n1459) );
  NANDN U1692 ( .A(n1468), .B(n1459), .Z(n1460) );
  XOR U1693 ( .A(n1461), .B(n1460), .Z(n1507) );
  XOR U1694 ( .A(n1484), .B(n1485), .Z(n1497) );
  NANDN U1695 ( .A(n[0]), .B(n1483), .Z(n1462) );
  NAND U1696 ( .A(n1497), .B(n1462), .Z(n1463) );
  NANDN U1697 ( .A(n[1]), .B(n1463), .Z(n1472) );
  ANDN U1698 ( .B(n1485), .A(n1464), .Z(n1465) );
  XNOR U1699 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1700 ( .A(n1483), .B(n1467), .Z(n1471) );
  NANDN U1701 ( .A(n1469), .B(n1468), .Z(n1470) );
  AND U1702 ( .A(n1471), .B(n1470), .Z(n1493) );
  NANDN U1703 ( .A(n1493), .B(n1782), .Z(n1502) );
  NAND U1704 ( .A(n1472), .B(n1502), .Z(n1473) );
  NANDN U1705 ( .A(n1782), .B(n1493), .Z(n1499) );
  NAND U1706 ( .A(n1473), .B(n1499), .Z(n1474) );
  NAND U1707 ( .A(n1507), .B(n1474), .Z(n1477) );
  XOR U1708 ( .A(n1507), .B(n1474), .Z(n1475) );
  NANDN U1709 ( .A(n1797), .B(n1475), .Z(n1476) );
  NAND U1710 ( .A(n1477), .B(n1476), .Z(n1480) );
  XOR U1711 ( .A(n1479), .B(n1478), .Z(n1508) );
  ANDN U1712 ( .B(n1480), .A(n1508), .Z(n1481) );
  NANDN U1713 ( .A(n1498), .B(n1481), .Z(n1505) );
  NAND U1714 ( .A(n1505), .B(n[0]), .Z(n1482) );
  XOR U1715 ( .A(n1483), .B(n1482), .Z(n1510) );
  ANDN U1716 ( .B(n[0]), .A(n1483), .Z(n1494) );
  XNOR U1717 ( .A(n1485), .B(n1484), .Z(n1486) );
  NANDN U1718 ( .A(n1494), .B(n1486), .Z(n1490) );
  NAND U1719 ( .A(n1487), .B(n1494), .Z(n1488) );
  NANDN U1720 ( .A(n[1]), .B(n1488), .Z(n1489) );
  NAND U1721 ( .A(n1490), .B(n1489), .Z(n1500) );
  XOR U1722 ( .A(n1782), .B(n1500), .Z(n1491) );
  NAND U1723 ( .A(n1505), .B(n1491), .Z(n1492) );
  XNOR U1724 ( .A(n1493), .B(n1492), .Z(n1512) );
  XOR U1725 ( .A(n[1]), .B(n1494), .Z(n1495) );
  AND U1726 ( .A(n1505), .B(n1495), .Z(n1496) );
  XOR U1727 ( .A(n1497), .B(n1496), .Z(n1620) );
  NAND U1728 ( .A(n1500), .B(n1499), .Z(n1501) );
  AND U1729 ( .A(n1502), .B(n1501), .Z(n1506) );
  XNOR U1730 ( .A(n1797), .B(n1506), .Z(n1503) );
  NAND U1731 ( .A(n1505), .B(n1503), .Z(n1504) );
  XNOR U1732 ( .A(n1507), .B(n1504), .Z(n1521) );
  AND U1733 ( .A(n[0]), .B(n1517), .Z(n1509) );
  XNOR U1734 ( .A(n1510), .B(n1509), .Z(n1806) );
  AND U1735 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1806), .Z(n1743) );
  AND U1736 ( .A(n1510), .B(n1509), .Z(n1619) );
  AND U1737 ( .A(n[1]), .B(n1517), .Z(n1622) );
  XNOR U1738 ( .A(n1512), .B(n1511), .Z(n1514) );
  ANDN U1739 ( .B(n1517), .A(n1782), .Z(n1513) );
  XNOR U1740 ( .A(n1514), .B(n1513), .Z(n1814) );
  NAND U1741 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1814), .Z(n1593) );
  ANDN U1742 ( .B(n1512), .A(n1511), .Z(n1516) );
  AND U1743 ( .A(n1514), .B(n1513), .Z(n1515) );
  NOR U1744 ( .A(n1516), .B(n1515), .Z(n1519) );
  ANDN U1745 ( .B(n1517), .A(n1797), .Z(n1518) );
  XNOR U1746 ( .A(n1519), .B(n1518), .Z(n1520) );
  XNOR U1747 ( .A(n1521), .B(n1520), .Z(n1818) );
  AND U1748 ( .A(m[2]), .B(n1818), .Z(n1533) );
  AND U1749 ( .A(m[3]), .B(n1818), .Z(n1542) );
  AND U1750 ( .A(m[1]), .B(n1818), .Z(n1529) );
  NAND U1751 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1818), .Z(n1531) );
  XNOR U1752 ( .A(n1797), .B(n1540), .Z(n1522) );
  NANDN U1753 ( .A(n1542), .B(n1522), .Z(n1524) );
  NANDN U1754 ( .A(n1797), .B(n1540), .Z(n1523) );
  NAND U1755 ( .A(n1524), .B(n1523), .Z(n1538) );
  NAND U1756 ( .A(n[0]), .B(n1531), .Z(n1526) );
  XNOR U1757 ( .A(n1782), .B(n1534), .Z(n1532) );
  NANDN U1758 ( .A(n1538), .B(n1532), .Z(n1525) );
  XOR U1759 ( .A(n1533), .B(n1525), .Z(n1543) );
  XNOR U1760 ( .A(n[1]), .B(n1526), .Z(n1527) );
  NANDN U1761 ( .A(n1538), .B(n1527), .Z(n1528) );
  XNOR U1762 ( .A(n1529), .B(n1528), .Z(n1545) );
  NANDN U1763 ( .A(n1538), .B(n[0]), .Z(n1530) );
  XNOR U1764 ( .A(n1531), .B(n1530), .Z(n1551) );
  IV U1765 ( .A(n1543), .Z(n1556) );
  NANDN U1766 ( .A(n1533), .B(n1532), .Z(n1536) );
  NANDN U1767 ( .A(n1782), .B(n1534), .Z(n1535) );
  AND U1768 ( .A(n1536), .B(n1535), .Z(n1541) );
  XOR U1769 ( .A(n1797), .B(n1541), .Z(n1537) );
  NANDN U1770 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1771 ( .A(n1542), .B(n1539), .Z(n1571) );
  NOR U1772 ( .A(n1782), .B(n1569), .Z(n1557) );
  XOR U1773 ( .A(n1543), .B(n1557), .Z(n1559) );
  ANDN U1774 ( .B(n[1]), .A(n1569), .Z(n1544) );
  NANDN U1775 ( .A(n1544), .B(n1545), .Z(n1547) );
  ANDN U1776 ( .B(n[0]), .A(n1569), .Z(n1550) );
  AND U1777 ( .A(n1551), .B(n1550), .Z(n1549) );
  XNOR U1778 ( .A(n1545), .B(n1544), .Z(n1548) );
  NANDN U1779 ( .A(n1549), .B(n1548), .Z(n1546) );
  NAND U1780 ( .A(n1547), .B(n1546), .Z(n1558) );
  XOR U1781 ( .A(n1559), .B(n1558), .Z(n1563) );
  IV U1782 ( .A(n1563), .Z(n1562) );
  XNOR U1783 ( .A(n1549), .B(n1548), .Z(n1552) );
  IV U1784 ( .A(n1552), .Z(n1581) );
  NANDN U1785 ( .A(n1581), .B(m[2]), .Z(n1555) );
  XOR U1786 ( .A(n1551), .B(n1550), .Z(n1583) );
  ANDN U1787 ( .B(m[1]), .A(n1583), .Z(n1578) );
  XOR U1788 ( .A(m[2]), .B(n1552), .Z(n1553) );
  NAND U1789 ( .A(n1578), .B(n1553), .Z(n1554) );
  AND U1790 ( .A(n1555), .B(n1554), .Z(n1564) );
  AND U1791 ( .A(n1601), .B(n1797), .Z(n1610) );
  NANDN U1792 ( .A(n1557), .B(n1556), .Z(n1561) );
  NAND U1793 ( .A(n1559), .B(n1558), .Z(n1560) );
  AND U1794 ( .A(n1561), .B(n1560), .Z(n1575) );
  ANDN U1795 ( .B(m[3]), .A(n1562), .Z(n1567) );
  XOR U1796 ( .A(m[3]), .B(n1563), .Z(n1565) );
  ANDN U1797 ( .B(n1565), .A(n1564), .Z(n1566) );
  OR U1798 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1799 ( .A(n1814), .B(n1568), .Z(n1577) );
  XOR U1800 ( .A(n1575), .B(n1577), .Z(n1573) );
  OR U1801 ( .A(n1569), .B(n1797), .Z(n1570) );
  AND U1802 ( .A(n1571), .B(n1570), .Z(n1574) );
  XNOR U1803 ( .A(n1577), .B(n1574), .Z(n1572) );
  NAND U1804 ( .A(n1573), .B(n1572), .Z(n1618) );
  XNOR U1805 ( .A(n1575), .B(n1574), .Z(n1576) );
  XNOR U1806 ( .A(n1577), .B(n1576), .Z(n1617) );
  ANDN U1807 ( .B(n1618), .A(n1617), .Z(n1590) );
  XOR U1808 ( .A(m[2]), .B(n1578), .Z(n1579) );
  NAND U1809 ( .A(n1814), .B(n1579), .Z(n1580) );
  XOR U1810 ( .A(n1581), .B(n1580), .Z(n1609) );
  OR U1811 ( .A(n1609), .B(n1782), .Z(n1598) );
  NOR U1812 ( .A(n1797), .B(n1601), .Z(n1613) );
  ANDN U1813 ( .B(n1598), .A(n1613), .Z(n1588) );
  NAND U1814 ( .A(n1814), .B(m[1]), .Z(n1582) );
  XOR U1815 ( .A(n1583), .B(n1582), .Z(n1605) );
  NANDN U1816 ( .A(n1605), .B(n[1]), .Z(n1595) );
  NOR U1817 ( .A(n1593), .B(n[0]), .Z(n1584) );
  NAND U1818 ( .A(n1595), .B(n1584), .Z(n1585) );
  NANDN U1819 ( .A(n1594), .B(n1585), .Z(n1586) );
  AND U1820 ( .A(n1609), .B(n1782), .Z(n1596) );
  OR U1821 ( .A(n1586), .B(n1596), .Z(n1587) );
  AND U1822 ( .A(n1588), .B(n1587), .Z(n1589) );
  ANDN U1823 ( .B(n1590), .A(n1589), .Z(n1591) );
  NANDN U1824 ( .A(n1610), .B(n1591), .Z(n1611) );
  NAND U1825 ( .A(n1611), .B(n[0]), .Z(n1592) );
  XNOR U1826 ( .A(n1593), .B(n1592), .Z(n1624) );
  NAND U1827 ( .A(n[0]), .B(n1593), .Z(n1602) );
  OR U1828 ( .A(n1596), .B(n1606), .Z(n1597) );
  AND U1829 ( .A(n1598), .B(n1597), .Z(n1612) );
  XOR U1830 ( .A(n1797), .B(n1612), .Z(n1599) );
  AND U1831 ( .A(n1611), .B(n1599), .Z(n1600) );
  XOR U1832 ( .A(n1601), .B(n1600), .Z(n1654) );
  XNOR U1833 ( .A(n[1]), .B(n1602), .Z(n1603) );
  NAND U1834 ( .A(n1611), .B(n1603), .Z(n1604) );
  XOR U1835 ( .A(n1605), .B(n1604), .Z(n1628) );
  XOR U1836 ( .A(n1782), .B(n1606), .Z(n1607) );
  AND U1837 ( .A(n1611), .B(n1607), .Z(n1608) );
  XOR U1838 ( .A(n1609), .B(n1608), .Z(n1644) );
  ANDN U1839 ( .B(n1611), .A(n1610), .Z(n1615) );
  NANDN U1840 ( .A(n1613), .B(n1612), .Z(n1614) );
  AND U1841 ( .A(n1615), .B(n1614), .Z(n1616) );
  XOR U1842 ( .A(n1617), .B(n1616), .Z(n1660) );
  AND U1843 ( .A(n[0]), .B(n1650), .Z(n1623) );
  NAND U1844 ( .A(n1624), .B(n1623), .Z(n1630) );
  NAND U1845 ( .A(n[1]), .B(n1650), .Z(n1627) );
  XNOR U1846 ( .A(n1628), .B(n1627), .Z(n1629) );
  XOR U1847 ( .A(n1630), .B(n1629), .Z(n1633) );
  XOR U1848 ( .A(n1620), .B(n1619), .Z(n1621) );
  XNOR U1849 ( .A(n1622), .B(n1621), .Z(n1809) );
  XNOR U1850 ( .A(n1624), .B(n1623), .Z(n1666) );
  AND U1851 ( .A(m[1]), .B(n1666), .Z(n1634) );
  XOR U1852 ( .A(n1634), .B(m[2]), .Z(n1625) );
  NAND U1853 ( .A(n1809), .B(n1625), .Z(n1626) );
  XOR U1854 ( .A(n1633), .B(n1626), .Z(n1675) );
  ANDN U1855 ( .B(n1650), .A(n1782), .Z(n1645) );
  XNOR U1856 ( .A(n1644), .B(n1645), .Z(n1647) );
  NANDN U1857 ( .A(n1628), .B(n1627), .Z(n1632) );
  NAND U1858 ( .A(n1630), .B(n1629), .Z(n1631) );
  NAND U1859 ( .A(n1632), .B(n1631), .Z(n1646) );
  XOR U1860 ( .A(n1647), .B(n1646), .Z(n1638) );
  IV U1861 ( .A(n1638), .Z(n1637) );
  XOR U1862 ( .A(m[3]), .B(n1639), .Z(n1635) );
  NAND U1863 ( .A(n1809), .B(n1635), .Z(n1636) );
  XOR U1864 ( .A(n1637), .B(n1636), .Z(n1687) );
  AND U1865 ( .A(n1687), .B(n1797), .Z(n1676) );
  ANDN U1866 ( .B(m[3]), .A(n1637), .Z(n1642) );
  XOR U1867 ( .A(m[3]), .B(n1638), .Z(n1640) );
  AND U1868 ( .A(n1640), .B(n1639), .Z(n1641) );
  OR U1869 ( .A(n1642), .B(n1641), .Z(n1643) );
  AND U1870 ( .A(n1809), .B(n1643), .Z(n1658) );
  NANDN U1871 ( .A(n1645), .B(n1644), .Z(n1649) );
  NAND U1872 ( .A(n1647), .B(n1646), .Z(n1648) );
  NAND U1873 ( .A(n1649), .B(n1648), .Z(n1651) );
  NANDN U1874 ( .A(n1797), .B(n1650), .Z(n1653) );
  XOR U1875 ( .A(n1654), .B(n1653), .Z(n1652) );
  XNOR U1876 ( .A(n1651), .B(n1652), .Z(n1657) );
  NOR U1877 ( .A(n1676), .B(n1682), .Z(n1663) );
  NAND U1878 ( .A(n1652), .B(n1651), .Z(n1656) );
  NAND U1879 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U1880 ( .A(n1656), .B(n1655), .Z(n1662) );
  ANDN U1881 ( .B(n1658), .A(n1657), .Z(n1659) );
  XNOR U1882 ( .A(n1660), .B(n1659), .Z(n1661) );
  XNOR U1883 ( .A(n1662), .B(n1661), .Z(n1683) );
  ANDN U1884 ( .B(n1663), .A(n1683), .Z(n1672) );
  NOR U1885 ( .A(n1797), .B(n1687), .Z(n1681) );
  ANDN U1886 ( .B(n1675), .A(n1782), .Z(n1678) );
  NOR U1887 ( .A(n1681), .B(n1678), .Z(n1670) );
  NAND U1888 ( .A(\MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1809), .Z(n1696) );
  OR U1889 ( .A(n[0]), .B(n1696), .Z(n1664) );
  NAND U1890 ( .A(n[1]), .B(n1664), .Z(n1667) );
  NAND U1891 ( .A(n1809), .B(m[1]), .Z(n1665) );
  XOR U1892 ( .A(n1666), .B(n1665), .Z(n1693) );
  ANDN U1893 ( .B(n1667), .A(n1693), .Z(n1668) );
  ANDN U1894 ( .B(n1782), .A(n1675), .Z(n1679) );
  OR U1895 ( .A(n1668), .B(n1679), .Z(n1669) );
  AND U1896 ( .A(n1670), .B(n1669), .Z(n1671) );
  ANDN U1897 ( .B(n1672), .A(n1671), .Z(n1694) );
  NAND U1898 ( .A(n[0]), .B(n1696), .Z(n1690) );
  XNOR U1899 ( .A(n1782), .B(n1677), .Z(n1673) );
  NANDN U1900 ( .A(n1694), .B(n1673), .Z(n1674) );
  XNOR U1901 ( .A(n1675), .B(n1674), .Z(n1699) );
  NANDN U1902 ( .A(n1782), .B(n1699), .Z(n1697) );
  OR U1903 ( .A(n1678), .B(n1677), .Z(n1680) );
  ANDN U1904 ( .B(n1680), .A(n1679), .Z(n1684) );
  NOR U1905 ( .A(n1733), .B(n1683), .Z(n1689) );
  XNOR U1906 ( .A(n1797), .B(n1684), .Z(n1685) );
  NANDN U1907 ( .A(n1694), .B(n1685), .Z(n1686) );
  XNOR U1908 ( .A(n1687), .B(n1686), .Z(n1726) );
  NAND U1909 ( .A(n1797), .B(n1726), .Z(n1688) );
  NAND U1910 ( .A(n1689), .B(n1688), .Z(n1698) );
  NANDN U1911 ( .A(n1697), .B(n1698), .Z(n1701) );
  XNOR U1912 ( .A(n[1]), .B(n1690), .Z(n1691) );
  NANDN U1913 ( .A(n1694), .B(n1691), .Z(n1692) );
  XNOR U1914 ( .A(n1693), .B(n1692), .Z(n1703) );
  NANDN U1915 ( .A(n1694), .B(n[0]), .Z(n1695) );
  XNOR U1916 ( .A(n1696), .B(n1695), .Z(n1709) );
  IV U1917 ( .A(n1704), .Z(n1721) );
  NAND U1918 ( .A(n1721), .B(n[2]), .Z(n1700) );
  ANDN U1919 ( .B(n1700), .A(n1699), .Z(n1719) );
  ANDN U1920 ( .B(n1701), .A(n1719), .Z(n1717) );
  ANDN U1921 ( .B(n[1]), .A(n1704), .Z(n1702) );
  XOR U1922 ( .A(n1703), .B(n1702), .Z(n1706) );
  ANDN U1923 ( .B(n[0]), .A(n1704), .Z(n1708) );
  NAND U1924 ( .A(n1709), .B(n1708), .Z(n1707) );
  IV U1925 ( .A(n1705), .Z(n1723) );
  ANDN U1926 ( .B(m[3]), .A(n1723), .Z(n1715) );
  XOR U1927 ( .A(m[3]), .B(n1705), .Z(n1713) );
  XNOR U1928 ( .A(n1707), .B(n1706), .Z(n1741) );
  NANDN U1929 ( .A(n1741), .B(m[2]), .Z(n1712) );
  XNOR U1930 ( .A(n1709), .B(n1708), .Z(n1737) );
  AND U1931 ( .A(m[1]), .B(n1737), .Z(n1738) );
  XNOR U1932 ( .A(m[2]), .B(n1741), .Z(n1710) );
  NAND U1933 ( .A(n1738), .B(n1710), .Z(n1711) );
  AND U1934 ( .A(n1712), .B(n1711), .Z(n1722) );
  ANDN U1935 ( .B(n1713), .A(n1722), .Z(n1714) );
  OR U1936 ( .A(n1715), .B(n1714), .Z(n1716) );
  AND U1937 ( .A(n1806), .B(n1716), .Z(n1731) );
  NANDN U1938 ( .A(n1718), .B(n1717), .Z(n1720) );
  ANDN U1939 ( .B(n1720), .A(n1719), .Z(n1725) );
  AND U1940 ( .A(n1721), .B(n[3]), .Z(n1727) );
  XNOR U1941 ( .A(n1726), .B(n1727), .Z(n1724) );
  XNOR U1942 ( .A(n1725), .B(n1724), .Z(n1730) );
  XOR U1943 ( .A(n1731), .B(n1730), .Z(n1758) );
  NANDN U1944 ( .A(n1725), .B(n1724), .Z(n1729) );
  NANDN U1945 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U1946 ( .A(n1729), .B(n1728), .Z(n1735) );
  AND U1947 ( .A(n1731), .B(n1730), .Z(n1732) );
  XNOR U1948 ( .A(n1733), .B(n1732), .Z(n1734) );
  XNOR U1949 ( .A(n1735), .B(n1734), .Z(n1759) );
  NAND U1950 ( .A(n1806), .B(m[1]), .Z(n1736) );
  XOR U1951 ( .A(n1737), .B(n1736), .Z(n1753) );
  NOR U1952 ( .A(n1753), .B(n[1]), .Z(n1744) );
  NAND U1953 ( .A(n[1]), .B(n1753), .Z(n1746) );
  XOR U1954 ( .A(n1738), .B(m[2]), .Z(n1739) );
  NAND U1955 ( .A(n1806), .B(n1739), .Z(n1740) );
  XNOR U1956 ( .A(n1741), .B(n1740), .Z(n1749) );
  NOR U1957 ( .A(n[2]), .B(n1749), .Z(n1756) );
  ANDN U1958 ( .B(n1749), .A(n1782), .Z(n1755) );
  NAND U1959 ( .A(n1762), .B(n[0]), .Z(n1742) );
  XOR U1960 ( .A(n1743), .B(n1742), .Z(n1775) );
  ANDN U1961 ( .B(n[0]), .A(n1743), .Z(n1750) );
  NANDN U1962 ( .A(n1744), .B(n1750), .Z(n1745) );
  AND U1963 ( .A(n1746), .B(n1745), .Z(n1754) );
  XOR U1964 ( .A(n1782), .B(n1754), .Z(n1747) );
  NAND U1965 ( .A(n1762), .B(n1747), .Z(n1748) );
  XNOR U1966 ( .A(n1749), .B(n1748), .Z(n1792) );
  XOR U1967 ( .A(n[1]), .B(n1750), .Z(n1751) );
  NAND U1968 ( .A(n1762), .B(n1751), .Z(n1752) );
  XNOR U1969 ( .A(n1753), .B(n1752), .Z(n1781) );
  NANDN U1970 ( .A(n1755), .B(n1754), .Z(n1757) );
  ANDN U1971 ( .B(n1757), .A(n1756), .Z(n1760) );
  XNOR U1972 ( .A(n1797), .B(n1760), .Z(n1761) );
  NAND U1973 ( .A(n1762), .B(n1761), .Z(n1763) );
  XNOR U1974 ( .A(n1764), .B(n1763), .Z(n1801) );
  AND U1975 ( .A(n[0]), .B(n1796), .Z(n1774) );
  XOR U1976 ( .A(n1775), .B(n1774), .Z(n1805) );
  NANDN U1977 ( .A(ereg[2]), .B(init), .Z(n1767) );
  OR U1978 ( .A(init), .B(e[2]), .Z(n1766) );
  AND U1979 ( .A(n1767), .B(n1766), .Z(n1822) );
  IV U1980 ( .A(n1822), .Z(n1815) );
  ANDN U1981 ( .B(n1823), .A(n1815), .Z(n1802) );
  NANDN U1982 ( .A(n1805), .B(n1802), .Z(n1769) );
  NANDN U1983 ( .A(n1823), .B(
        \MODMULT2[1].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1768)
         );
  NAND U1984 ( .A(n1769), .B(n1768), .Z(n1771) );
  NANDN U1985 ( .A(n1822), .B(n1823), .Z(n1787) );
  NANDN U1986 ( .A(n1787), .B(n1806), .Z(n1770) );
  NANDN U1987 ( .A(n1771), .B(n1770), .Z(N10) );
  NANDN U1988 ( .A(n1787), .B(n1809), .Z(n1773) );
  NANDN U1989 ( .A(n1823), .B(m[1]), .Z(n1772) );
  AND U1990 ( .A(n1773), .B(n1772), .Z(n1778) );
  AND U1991 ( .A(n[1]), .B(n1796), .Z(n1779) );
  NAND U1992 ( .A(n1775), .B(n1774), .Z(n1780) );
  XOR U1993 ( .A(n1781), .B(n1780), .Z(n1776) );
  XOR U1994 ( .A(n1779), .B(n1776), .Z(n1810) );
  NAND U1995 ( .A(n1802), .B(n1810), .Z(n1777) );
  NAND U1996 ( .A(n1778), .B(n1777), .Z(N11) );
  XNOR U1997 ( .A(n1792), .B(n1793), .Z(n1791) );
  ANDN U1998 ( .B(n1796), .A(n1782), .Z(n1790) );
  XOR U1999 ( .A(n1791), .B(n1790), .Z(n1813) );
  NANDN U2000 ( .A(n1813), .B(n1802), .Z(n1784) );
  NANDN U2001 ( .A(n1823), .B(m[2]), .Z(n1783) );
  NAND U2002 ( .A(n1784), .B(n1783), .Z(n1786) );
  NANDN U2003 ( .A(n1787), .B(n1814), .Z(n1785) );
  NANDN U2004 ( .A(n1786), .B(n1785), .Z(N12) );
  NANDN U2005 ( .A(n1787), .B(n1818), .Z(n1789) );
  NANDN U2006 ( .A(n1823), .B(m[3]), .Z(n1788) );
  AND U2007 ( .A(n1789), .B(n1788), .Z(n1804) );
  NAND U2008 ( .A(n1791), .B(n1790), .Z(n1795) );
  NANDN U2009 ( .A(n1793), .B(n1792), .Z(n1794) );
  AND U2010 ( .A(n1795), .B(n1794), .Z(n1799) );
  NANDN U2011 ( .A(n1797), .B(n1796), .Z(n1798) );
  XNOR U2012 ( .A(n1799), .B(n1798), .Z(n1800) );
  XNOR U2013 ( .A(n1801), .B(n1800), .Z(n1819) );
  NAND U2014 ( .A(n1802), .B(n1819), .Z(n1803) );
  NAND U2015 ( .A(n1804), .B(n1803), .Z(N13) );
  OR U2016 ( .A(n1805), .B(n1815), .Z(n1808) );
  NAND U2017 ( .A(n1815), .B(n1806), .Z(n1807) );
  NAND U2018 ( .A(n1808), .B(n1807), .Z(c[0]) );
  NANDN U2019 ( .A(n1822), .B(n1809), .Z(n1812) );
  NAND U2020 ( .A(n1822), .B(n1810), .Z(n1811) );
  NAND U2021 ( .A(n1812), .B(n1811), .Z(c[1]) );
  OR U2022 ( .A(n1813), .B(n1815), .Z(n1817) );
  NAND U2023 ( .A(n1815), .B(n1814), .Z(n1816) );
  NAND U2024 ( .A(n1817), .B(n1816), .Z(c[2]) );
  NANDN U2025 ( .A(n1822), .B(n1818), .Z(n1821) );
  NAND U2026 ( .A(n1822), .B(n1819), .Z(n1820) );
  NAND U2027 ( .A(n1821), .B(n1820), .Z(c[3]) );
  ANDN U2028 ( .B(e[0]), .A(init), .Z(ein[0]) );
  ANDN U2029 ( .B(e[1]), .A(init), .Z(ein[1]) );
  OR U2030 ( .A(n1823), .B(n1822), .Z(n6) );
endmodule

