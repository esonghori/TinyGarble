
module SubBytes_0 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U2967 ( .A(n3911), .B(n3519), .Z(n3521) );
  AND U2968 ( .A(n3543), .B(n3528), .Z(n1966) );
  NAND U2969 ( .A(n3514), .B(n1966), .Z(n1967) );
  NANDN U2970 ( .A(n3528), .B(n3543), .Z(n1968) );
  XNOR U2971 ( .A(x[96]), .B(n1968), .Z(n1969) );
  NANDN U2972 ( .A(n3514), .B(n1969), .Z(n1970) );
  NAND U2973 ( .A(n1967), .B(n1970), .Z(n1971) );
  XNOR U2974 ( .A(n3469), .B(n3472), .Z(n1972) );
  XNOR U2975 ( .A(n1971), .B(n1972), .Z(n3497) );
  XNOR U2976 ( .A(n2823), .B(n2821), .Z(n1973) );
  NANDN U2977 ( .A(n2826), .B(n1973), .Z(n1974) );
  NAND U2978 ( .A(n2826), .B(n2822), .Z(n1975) );
  NANDN U2979 ( .A(n2825), .B(n1975), .Z(n1976) );
  NAND U2980 ( .A(n1974), .B(n1976), .Z(n2881) );
  XNOR U2981 ( .A(n2938), .B(n2936), .Z(n1977) );
  NANDN U2982 ( .A(n2941), .B(n1977), .Z(n1978) );
  NAND U2983 ( .A(n2941), .B(n2937), .Z(n1979) );
  NANDN U2984 ( .A(n2940), .B(n1979), .Z(n1980) );
  NAND U2985 ( .A(n1978), .B(n1980), .Z(n2996) );
  XNOR U2986 ( .A(n3398), .B(n3396), .Z(n1981) );
  NANDN U2987 ( .A(n3401), .B(n1981), .Z(n1982) );
  NAND U2988 ( .A(n3401), .B(n3397), .Z(n1983) );
  NANDN U2989 ( .A(n3400), .B(n1983), .Z(n1984) );
  NAND U2990 ( .A(n1982), .B(n1984), .Z(n3456) );
  AND U2991 ( .A(n2297), .B(n2296), .Z(n1985) );
  XNOR U2992 ( .A(n2295), .B(n1985), .Z(n2309) );
  XNOR U2993 ( .A(n2708), .B(n2706), .Z(n1986) );
  NANDN U2994 ( .A(n2711), .B(n1986), .Z(n1987) );
  NAND U2995 ( .A(n2711), .B(n2707), .Z(n1988) );
  NANDN U2996 ( .A(n2710), .B(n1988), .Z(n1989) );
  NAND U2997 ( .A(n1987), .B(n1989), .Z(n2766) );
  XNOR U2998 ( .A(n2478), .B(n2476), .Z(n1990) );
  NANDN U2999 ( .A(n2481), .B(n1990), .Z(n1991) );
  NAND U3000 ( .A(n2481), .B(n2477), .Z(n1992) );
  NANDN U3001 ( .A(n2480), .B(n1992), .Z(n1993) );
  NAND U3002 ( .A(n1991), .B(n1993), .Z(n2536) );
  XNOR U3003 ( .A(n3168), .B(n3166), .Z(n1994) );
  NANDN U3004 ( .A(n3171), .B(n1994), .Z(n1995) );
  NAND U3005 ( .A(n3171), .B(n3167), .Z(n1996) );
  NANDN U3006 ( .A(n3170), .B(n1996), .Z(n1997) );
  NAND U3007 ( .A(n1995), .B(n1997), .Z(n3226) );
  XNOR U3008 ( .A(n3727), .B(n3725), .Z(n1998) );
  NANDN U3009 ( .A(n3730), .B(n1998), .Z(n1999) );
  NAND U3010 ( .A(n3730), .B(n3726), .Z(n2000) );
  NANDN U3011 ( .A(n3729), .B(n2000), .Z(n2001) );
  NAND U3012 ( .A(n1999), .B(n2001), .Z(n3785) );
  XNOR U3013 ( .A(n2593), .B(n2591), .Z(n2002) );
  NANDN U3014 ( .A(n2596), .B(n2002), .Z(n2003) );
  NAND U3015 ( .A(n2596), .B(n2592), .Z(n2004) );
  NANDN U3016 ( .A(n2595), .B(n2004), .Z(n2005) );
  NAND U3017 ( .A(n2003), .B(n2005), .Z(n2651) );
  XNOR U3018 ( .A(n3842), .B(n3840), .Z(n2006) );
  NANDN U3019 ( .A(n3845), .B(n2006), .Z(n2007) );
  NAND U3020 ( .A(n3845), .B(n3841), .Z(n2008) );
  NANDN U3021 ( .A(n3844), .B(n2008), .Z(n2009) );
  NAND U3022 ( .A(n2007), .B(n2009), .Z(n3900) );
  XNOR U3023 ( .A(n3283), .B(n3281), .Z(n2010) );
  NANDN U3024 ( .A(n3286), .B(n2010), .Z(n2011) );
  NAND U3025 ( .A(n3286), .B(n3282), .Z(n2012) );
  NANDN U3026 ( .A(n3285), .B(n2012), .Z(n2013) );
  NAND U3027 ( .A(n2011), .B(n2013), .Z(n3341) );
  XNOR U3028 ( .A(n2135), .B(n2133), .Z(n2014) );
  NANDN U3029 ( .A(n2138), .B(n2014), .Z(n2015) );
  NAND U3030 ( .A(n2138), .B(n2134), .Z(n2016) );
  NANDN U3031 ( .A(n2137), .B(n2016), .Z(n2017) );
  NAND U3032 ( .A(n2015), .B(n2017), .Z(n2193) );
  XNOR U3033 ( .A(n3612), .B(n3610), .Z(n2018) );
  NANDN U3034 ( .A(n3615), .B(n2018), .Z(n2019) );
  NAND U3035 ( .A(n3615), .B(n3611), .Z(n2020) );
  NANDN U3036 ( .A(n3614), .B(n2020), .Z(n2021) );
  NAND U3037 ( .A(n2019), .B(n2021), .Z(n3670) );
  XNOR U3038 ( .A(n2363), .B(n2361), .Z(n2022) );
  NANDN U3039 ( .A(n2366), .B(n2022), .Z(n2023) );
  NAND U3040 ( .A(n2366), .B(n2362), .Z(n2024) );
  NANDN U3041 ( .A(n2365), .B(n2024), .Z(n2025) );
  NAND U3042 ( .A(n2023), .B(n2025), .Z(n2421) );
  XNOR U3043 ( .A(n3053), .B(n3051), .Z(n2026) );
  NANDN U3044 ( .A(n3056), .B(n2026), .Z(n2027) );
  NAND U3045 ( .A(n3056), .B(n3052), .Z(n2028) );
  NANDN U3046 ( .A(n3055), .B(n2028), .Z(n2029) );
  NAND U3047 ( .A(n2027), .B(n2029), .Z(n3111) );
  XOR U3048 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3049 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3050 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3051 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3052 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3053 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3054 ( .A(n2522), .B(n2536), .Z(n2499) );
  ANDN U3055 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3056 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3057 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3058 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3059 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3060 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3061 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3062 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3063 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3064 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U3065 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3066 ( .A(n2407), .B(n2421), .Z(n2384) );
  NANDN U3067 ( .A(n2825), .B(n2826), .Z(n2032) );
  AND U3068 ( .A(n2825), .B(n2823), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n2824), .Z(n2034) );
  NANDN U3070 ( .A(n2826), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n2840) );
  NANDN U3072 ( .A(n2595), .B(n2596), .Z(n2036) );
  AND U3073 ( .A(n2595), .B(n2593), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n2594), .Z(n2038) );
  NANDN U3075 ( .A(n2596), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n2610) );
  NANDN U3077 ( .A(n2940), .B(n2941), .Z(n2040) );
  AND U3078 ( .A(n2940), .B(n2938), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n2939), .Z(n2042) );
  NANDN U3080 ( .A(n2941), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n2955) );
  NANDN U3082 ( .A(n3844), .B(n3845), .Z(n2044) );
  AND U3083 ( .A(n3844), .B(n3842), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n3843), .Z(n2046) );
  NANDN U3085 ( .A(n3845), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n3859) );
  NANDN U3087 ( .A(n2480), .B(n2481), .Z(n2048) );
  AND U3088 ( .A(n2480), .B(n2478), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n2479), .Z(n2050) );
  NANDN U3090 ( .A(n2481), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n2495) );
  NANDN U3092 ( .A(n2710), .B(n2711), .Z(n2052) );
  AND U3093 ( .A(n2710), .B(n2708), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n2709), .Z(n2054) );
  NANDN U3095 ( .A(n2711), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n2725) );
  NANDN U3097 ( .A(n3400), .B(n3401), .Z(n2056) );
  AND U3098 ( .A(n3400), .B(n3398), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n3399), .Z(n2058) );
  NANDN U3100 ( .A(n3401), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n3415) );
  XOR U3102 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3103 ( .A(n3285), .B(n3286), .Z(n2060) );
  AND U3104 ( .A(n3285), .B(n3283), .Z(n2061) );
  XNOR U3105 ( .A(n2061), .B(n3284), .Z(n2062) );
  NANDN U3106 ( .A(n3286), .B(n2062), .Z(n2063) );
  NAND U3107 ( .A(n2060), .B(n2063), .Z(n3300) );
  NANDN U3108 ( .A(n3170), .B(n3171), .Z(n2064) );
  AND U3109 ( .A(n3170), .B(n3168), .Z(n2065) );
  XNOR U3110 ( .A(n2065), .B(n3169), .Z(n2066) );
  NANDN U3111 ( .A(n3171), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2064), .B(n2067), .Z(n3185) );
  NANDN U3113 ( .A(n3729), .B(n3730), .Z(n2068) );
  AND U3114 ( .A(n3729), .B(n3727), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n3728), .Z(n2070) );
  NANDN U3116 ( .A(n3730), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n3744) );
  NANDN U3118 ( .A(n2137), .B(n2138), .Z(n2072) );
  AND U3119 ( .A(n2137), .B(n2135), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n2136), .Z(n2074) );
  NANDN U3121 ( .A(n2138), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n2152) );
  NANDN U3123 ( .A(n3614), .B(n3615), .Z(n2076) );
  AND U3124 ( .A(n3614), .B(n3612), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3613), .Z(n2078) );
  NANDN U3126 ( .A(n3615), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3629) );
  NANDN U3128 ( .A(n3055), .B(n3056), .Z(n2080) );
  AND U3129 ( .A(n3055), .B(n3053), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n3054), .Z(n2082) );
  NANDN U3131 ( .A(n3056), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n3070) );
  NANDN U3133 ( .A(n2365), .B(n2366), .Z(n2084) );
  AND U3134 ( .A(n2365), .B(n2363), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n2364), .Z(n2086) );
  NANDN U3136 ( .A(n2366), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n2380) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_1 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  XOR U2962 ( .A(n3544), .B(n3555), .Z(n3542) );
  AND U2963 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2964 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2965 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2966 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2967 ( .A(n3911), .B(n3519), .Z(n3521) );
  XNOR U2968 ( .A(n2593), .B(n2591), .Z(n1966) );
  NANDN U2969 ( .A(n2596), .B(n1966), .Z(n1967) );
  NAND U2970 ( .A(n2596), .B(n2592), .Z(n1968) );
  NANDN U2971 ( .A(n2595), .B(n1968), .Z(n1969) );
  NAND U2972 ( .A(n1967), .B(n1969), .Z(n2651) );
  XNOR U2973 ( .A(n3168), .B(n3166), .Z(n1970) );
  NANDN U2974 ( .A(n3171), .B(n1970), .Z(n1971) );
  NAND U2975 ( .A(n3171), .B(n3167), .Z(n1972) );
  NANDN U2976 ( .A(n3170), .B(n1972), .Z(n1973) );
  NAND U2977 ( .A(n1971), .B(n1973), .Z(n3226) );
  XNOR U2978 ( .A(n3727), .B(n3725), .Z(n1974) );
  NANDN U2979 ( .A(n3730), .B(n1974), .Z(n1975) );
  NAND U2980 ( .A(n3730), .B(n3726), .Z(n1976) );
  NANDN U2981 ( .A(n3729), .B(n1976), .Z(n1977) );
  NAND U2982 ( .A(n1975), .B(n1977), .Z(n3785) );
  XNOR U2983 ( .A(n2478), .B(n2476), .Z(n1978) );
  NANDN U2984 ( .A(n2481), .B(n1978), .Z(n1979) );
  NAND U2985 ( .A(n2481), .B(n2477), .Z(n1980) );
  NANDN U2986 ( .A(n2480), .B(n1980), .Z(n1981) );
  NAND U2987 ( .A(n1979), .B(n1981), .Z(n2536) );
  XNOR U2988 ( .A(n3053), .B(n3051), .Z(n1982) );
  NANDN U2989 ( .A(n3056), .B(n1982), .Z(n1983) );
  NAND U2990 ( .A(n3056), .B(n3052), .Z(n1984) );
  NANDN U2991 ( .A(n3055), .B(n1984), .Z(n1985) );
  NAND U2992 ( .A(n1983), .B(n1985), .Z(n3111) );
  XNOR U2993 ( .A(n3612), .B(n3610), .Z(n1986) );
  NANDN U2994 ( .A(n3615), .B(n1986), .Z(n1987) );
  NAND U2995 ( .A(n3615), .B(n3611), .Z(n1988) );
  NANDN U2996 ( .A(n3614), .B(n1988), .Z(n1989) );
  NAND U2997 ( .A(n1987), .B(n1989), .Z(n3670) );
  XNOR U2998 ( .A(n2363), .B(n2361), .Z(n1990) );
  NANDN U2999 ( .A(n2366), .B(n1990), .Z(n1991) );
  NAND U3000 ( .A(n2366), .B(n2362), .Z(n1992) );
  NANDN U3001 ( .A(n2365), .B(n1992), .Z(n1993) );
  NAND U3002 ( .A(n1991), .B(n1993), .Z(n2421) );
  XNOR U3003 ( .A(n2938), .B(n2936), .Z(n1994) );
  NANDN U3004 ( .A(n2941), .B(n1994), .Z(n1995) );
  NAND U3005 ( .A(n2941), .B(n2937), .Z(n1996) );
  NANDN U3006 ( .A(n2940), .B(n1996), .Z(n1997) );
  NAND U3007 ( .A(n1995), .B(n1997), .Z(n2996) );
  AND U3008 ( .A(n3543), .B(n3528), .Z(n1998) );
  NAND U3009 ( .A(n3514), .B(n1998), .Z(n1999) );
  NANDN U3010 ( .A(n3528), .B(n3543), .Z(n2000) );
  XNOR U3011 ( .A(x[96]), .B(n2000), .Z(n2001) );
  NANDN U3012 ( .A(n3514), .B(n2001), .Z(n2002) );
  NAND U3013 ( .A(n1999), .B(n2002), .Z(n2003) );
  XNOR U3014 ( .A(n3469), .B(n3472), .Z(n2004) );
  XNOR U3015 ( .A(n2003), .B(n2004), .Z(n3497) );
  AND U3016 ( .A(n2297), .B(n2296), .Z(n2005) );
  XNOR U3017 ( .A(n2295), .B(n2005), .Z(n2309) );
  XNOR U3018 ( .A(n2823), .B(n2821), .Z(n2006) );
  NANDN U3019 ( .A(n2826), .B(n2006), .Z(n2007) );
  NAND U3020 ( .A(n2826), .B(n2822), .Z(n2008) );
  NANDN U3021 ( .A(n2825), .B(n2008), .Z(n2009) );
  NAND U3022 ( .A(n2007), .B(n2009), .Z(n2881) );
  XNOR U3023 ( .A(n3398), .B(n3396), .Z(n2010) );
  NANDN U3024 ( .A(n3401), .B(n2010), .Z(n2011) );
  NAND U3025 ( .A(n3401), .B(n3397), .Z(n2012) );
  NANDN U3026 ( .A(n3400), .B(n2012), .Z(n2013) );
  NAND U3027 ( .A(n2011), .B(n2013), .Z(n3456) );
  XNOR U3028 ( .A(n2135), .B(n2133), .Z(n2014) );
  NANDN U3029 ( .A(n2138), .B(n2014), .Z(n2015) );
  NAND U3030 ( .A(n2138), .B(n2134), .Z(n2016) );
  NANDN U3031 ( .A(n2137), .B(n2016), .Z(n2017) );
  NAND U3032 ( .A(n2015), .B(n2017), .Z(n2193) );
  XNOR U3033 ( .A(n2708), .B(n2706), .Z(n2018) );
  NANDN U3034 ( .A(n2711), .B(n2018), .Z(n2019) );
  NAND U3035 ( .A(n2711), .B(n2707), .Z(n2020) );
  NANDN U3036 ( .A(n2710), .B(n2020), .Z(n2021) );
  NAND U3037 ( .A(n2019), .B(n2021), .Z(n2766) );
  XNOR U3038 ( .A(n3283), .B(n3281), .Z(n2022) );
  NANDN U3039 ( .A(n3286), .B(n2022), .Z(n2023) );
  NAND U3040 ( .A(n3286), .B(n3282), .Z(n2024) );
  NANDN U3041 ( .A(n3285), .B(n2024), .Z(n2025) );
  NAND U3042 ( .A(n2023), .B(n2025), .Z(n3341) );
  XNOR U3043 ( .A(n3842), .B(n3840), .Z(n2026) );
  NANDN U3044 ( .A(n3845), .B(n2026), .Z(n2027) );
  NAND U3045 ( .A(n3845), .B(n3841), .Z(n2028) );
  NANDN U3046 ( .A(n3844), .B(n2028), .Z(n2029) );
  NAND U3047 ( .A(n2027), .B(n2029), .Z(n3900) );
  XOR U3048 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3049 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3050 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3051 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3052 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3053 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3054 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3055 ( .A(n2982), .B(n2996), .Z(n2959) );
  ANDN U3056 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3057 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3058 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3059 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3060 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3061 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3062 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3063 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3064 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3065 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U3066 ( .A(n3470), .B(n3471), .Z(n3546) );
  NANDN U3067 ( .A(n2595), .B(n2596), .Z(n2032) );
  AND U3068 ( .A(n2595), .B(n2593), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n2594), .Z(n2034) );
  NANDN U3070 ( .A(n2596), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n2610) );
  NANDN U3072 ( .A(n3170), .B(n3171), .Z(n2036) );
  AND U3073 ( .A(n3170), .B(n3168), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n3169), .Z(n2038) );
  NANDN U3075 ( .A(n3171), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n3185) );
  NANDN U3077 ( .A(n3729), .B(n3730), .Z(n2040) );
  AND U3078 ( .A(n3729), .B(n3727), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n3728), .Z(n2042) );
  NANDN U3080 ( .A(n3730), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n3744) );
  NANDN U3082 ( .A(n2480), .B(n2481), .Z(n2044) );
  AND U3083 ( .A(n2480), .B(n2478), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n2479), .Z(n2046) );
  NANDN U3085 ( .A(n2481), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n2495) );
  NANDN U3087 ( .A(n3055), .B(n3056), .Z(n2048) );
  AND U3088 ( .A(n3055), .B(n3053), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n3054), .Z(n2050) );
  NANDN U3090 ( .A(n3056), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n3070) );
  NANDN U3092 ( .A(n3614), .B(n3615), .Z(n2052) );
  AND U3093 ( .A(n3614), .B(n3612), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n3613), .Z(n2054) );
  NANDN U3095 ( .A(n3615), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n3629) );
  NANDN U3097 ( .A(n2365), .B(n2366), .Z(n2056) );
  AND U3098 ( .A(n2365), .B(n2363), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n2364), .Z(n2058) );
  NANDN U3100 ( .A(n2366), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n2380) );
  NANDN U3102 ( .A(n2940), .B(n2941), .Z(n2060) );
  AND U3103 ( .A(n2940), .B(n2938), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n2939), .Z(n2062) );
  NANDN U3105 ( .A(n2941), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n2955) );
  XOR U3107 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3108 ( .A(n2825), .B(n2826), .Z(n2064) );
  AND U3109 ( .A(n2825), .B(n2823), .Z(n2065) );
  XNOR U3110 ( .A(n2065), .B(n2824), .Z(n2066) );
  NANDN U3111 ( .A(n2826), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2064), .B(n2067), .Z(n2840) );
  NANDN U3113 ( .A(n3400), .B(n3401), .Z(n2068) );
  AND U3114 ( .A(n3400), .B(n3398), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n3399), .Z(n2070) );
  NANDN U3116 ( .A(n3401), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n3415) );
  NANDN U3118 ( .A(n2137), .B(n2138), .Z(n2072) );
  AND U3119 ( .A(n2137), .B(n2135), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n2136), .Z(n2074) );
  NANDN U3121 ( .A(n2138), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n2152) );
  NANDN U3123 ( .A(n2710), .B(n2711), .Z(n2076) );
  AND U3124 ( .A(n2710), .B(n2708), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n2709), .Z(n2078) );
  NANDN U3126 ( .A(n2711), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n2725) );
  NANDN U3128 ( .A(n3285), .B(n3286), .Z(n2080) );
  AND U3129 ( .A(n3285), .B(n3283), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n3284), .Z(n2082) );
  NANDN U3131 ( .A(n3286), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n3300) );
  NANDN U3133 ( .A(n3844), .B(n3845), .Z(n2084) );
  AND U3134 ( .A(n3844), .B(n3842), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3843), .Z(n2086) );
  NANDN U3136 ( .A(n3845), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3859) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_2 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3544), .B(n3555), .Z(n3542) );
  XNOR U2967 ( .A(n2708), .B(n2706), .Z(n1966) );
  NANDN U2968 ( .A(n2711), .B(n1966), .Z(n1967) );
  NAND U2969 ( .A(n2711), .B(n2707), .Z(n1968) );
  NANDN U2970 ( .A(n2710), .B(n1968), .Z(n1969) );
  NAND U2971 ( .A(n1967), .B(n1969), .Z(n2766) );
  XNOR U2972 ( .A(n2938), .B(n2936), .Z(n1970) );
  NANDN U2973 ( .A(n2941), .B(n1970), .Z(n1971) );
  NAND U2974 ( .A(n2941), .B(n2937), .Z(n1972) );
  NANDN U2975 ( .A(n2940), .B(n1972), .Z(n1973) );
  NAND U2976 ( .A(n1971), .B(n1973), .Z(n2996) );
  XOR U2977 ( .A(n3911), .B(n3519), .Z(n3521) );
  AND U2978 ( .A(n3543), .B(n3528), .Z(n1974) );
  NAND U2979 ( .A(n3514), .B(n1974), .Z(n1975) );
  NANDN U2980 ( .A(n3528), .B(n3543), .Z(n1976) );
  XNOR U2981 ( .A(x[96]), .B(n1976), .Z(n1977) );
  NANDN U2982 ( .A(n3514), .B(n1977), .Z(n1978) );
  NAND U2983 ( .A(n1975), .B(n1978), .Z(n1979) );
  XNOR U2984 ( .A(n3469), .B(n3472), .Z(n1980) );
  XNOR U2985 ( .A(n1979), .B(n1980), .Z(n3497) );
  XNOR U2986 ( .A(n2823), .B(n2821), .Z(n1981) );
  NANDN U2987 ( .A(n2826), .B(n1981), .Z(n1982) );
  NAND U2988 ( .A(n2826), .B(n2822), .Z(n1983) );
  NANDN U2989 ( .A(n2825), .B(n1983), .Z(n1984) );
  NAND U2990 ( .A(n1982), .B(n1984), .Z(n2881) );
  XNOR U2991 ( .A(n2478), .B(n2476), .Z(n1985) );
  NANDN U2992 ( .A(n2481), .B(n1985), .Z(n1986) );
  NAND U2993 ( .A(n2481), .B(n2477), .Z(n1987) );
  NANDN U2994 ( .A(n2480), .B(n1987), .Z(n1988) );
  NAND U2995 ( .A(n1986), .B(n1988), .Z(n2536) );
  XNOR U2996 ( .A(n3612), .B(n3610), .Z(n1989) );
  NANDN U2997 ( .A(n3615), .B(n1989), .Z(n1990) );
  NAND U2998 ( .A(n3615), .B(n3611), .Z(n1991) );
  NANDN U2999 ( .A(n3614), .B(n1991), .Z(n1992) );
  NAND U3000 ( .A(n1990), .B(n1992), .Z(n3670) );
  XNOR U3001 ( .A(n2363), .B(n2361), .Z(n1993) );
  NANDN U3002 ( .A(n2366), .B(n1993), .Z(n1994) );
  NAND U3003 ( .A(n2366), .B(n2362), .Z(n1995) );
  NANDN U3004 ( .A(n2365), .B(n1995), .Z(n1996) );
  NAND U3005 ( .A(n1994), .B(n1996), .Z(n2421) );
  XNOR U3006 ( .A(n3053), .B(n3051), .Z(n1997) );
  NANDN U3007 ( .A(n3056), .B(n1997), .Z(n1998) );
  NAND U3008 ( .A(n3056), .B(n3052), .Z(n1999) );
  NANDN U3009 ( .A(n3055), .B(n1999), .Z(n2000) );
  NAND U3010 ( .A(n1998), .B(n2000), .Z(n3111) );
  AND U3011 ( .A(n2297), .B(n2296), .Z(n2001) );
  XNOR U3012 ( .A(n2295), .B(n2001), .Z(n2309) );
  XNOR U3013 ( .A(n3398), .B(n3396), .Z(n2002) );
  NANDN U3014 ( .A(n3401), .B(n2002), .Z(n2003) );
  NAND U3015 ( .A(n3401), .B(n3397), .Z(n2004) );
  NANDN U3016 ( .A(n3400), .B(n2004), .Z(n2005) );
  NAND U3017 ( .A(n2003), .B(n2005), .Z(n3456) );
  XNOR U3018 ( .A(n3842), .B(n3840), .Z(n2006) );
  NANDN U3019 ( .A(n3845), .B(n2006), .Z(n2007) );
  NAND U3020 ( .A(n3845), .B(n3841), .Z(n2008) );
  NANDN U3021 ( .A(n3844), .B(n2008), .Z(n2009) );
  NAND U3022 ( .A(n2007), .B(n2009), .Z(n3900) );
  XNOR U3023 ( .A(n2135), .B(n2133), .Z(n2010) );
  NANDN U3024 ( .A(n2138), .B(n2010), .Z(n2011) );
  NAND U3025 ( .A(n2138), .B(n2134), .Z(n2012) );
  NANDN U3026 ( .A(n2137), .B(n2012), .Z(n2013) );
  NAND U3027 ( .A(n2011), .B(n2013), .Z(n2193) );
  XNOR U3028 ( .A(n3283), .B(n3281), .Z(n2014) );
  NANDN U3029 ( .A(n3286), .B(n2014), .Z(n2015) );
  NAND U3030 ( .A(n3286), .B(n3282), .Z(n2016) );
  NANDN U3031 ( .A(n3285), .B(n2016), .Z(n2017) );
  NAND U3032 ( .A(n2015), .B(n2017), .Z(n3341) );
  XNOR U3033 ( .A(n2593), .B(n2591), .Z(n2018) );
  NANDN U3034 ( .A(n2596), .B(n2018), .Z(n2019) );
  NAND U3035 ( .A(n2596), .B(n2592), .Z(n2020) );
  NANDN U3036 ( .A(n2595), .B(n2020), .Z(n2021) );
  NAND U3037 ( .A(n2019), .B(n2021), .Z(n2651) );
  XNOR U3038 ( .A(n3168), .B(n3166), .Z(n2022) );
  NANDN U3039 ( .A(n3171), .B(n2022), .Z(n2023) );
  NAND U3040 ( .A(n3171), .B(n3167), .Z(n2024) );
  NANDN U3041 ( .A(n3170), .B(n2024), .Z(n2025) );
  NAND U3042 ( .A(n2023), .B(n2025), .Z(n3226) );
  XNOR U3043 ( .A(n3727), .B(n3725), .Z(n2026) );
  NANDN U3044 ( .A(n3730), .B(n2026), .Z(n2027) );
  NAND U3045 ( .A(n3730), .B(n3726), .Z(n2028) );
  NANDN U3046 ( .A(n3729), .B(n2028), .Z(n2029) );
  NAND U3047 ( .A(n2027), .B(n2029), .Z(n3785) );
  XOR U3048 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3049 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3050 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3051 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3052 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3053 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3054 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3055 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3056 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3057 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3058 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3059 ( .A(n2407), .B(n2421), .Z(n2384) );
  ANDN U3060 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3061 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3062 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3063 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3064 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3065 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U3066 ( .A(n3470), .B(n3471), .Z(n3546) );
  NANDN U3067 ( .A(n2710), .B(n2711), .Z(n2032) );
  AND U3068 ( .A(n2710), .B(n2708), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n2709), .Z(n2034) );
  NANDN U3070 ( .A(n2711), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n2725) );
  NANDN U3072 ( .A(n3285), .B(n3286), .Z(n2036) );
  AND U3073 ( .A(n3285), .B(n3283), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n3284), .Z(n2038) );
  NANDN U3075 ( .A(n3286), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n3300) );
  NANDN U3077 ( .A(n2940), .B(n2941), .Z(n2040) );
  AND U3078 ( .A(n2940), .B(n2938), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n2939), .Z(n2042) );
  NANDN U3080 ( .A(n2941), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n2955) );
  NANDN U3082 ( .A(n3844), .B(n3845), .Z(n2044) );
  AND U3083 ( .A(n3844), .B(n3842), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n3843), .Z(n2046) );
  NANDN U3085 ( .A(n3845), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n3859) );
  NANDN U3087 ( .A(n2595), .B(n2596), .Z(n2048) );
  AND U3088 ( .A(n2595), .B(n2593), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n2594), .Z(n2050) );
  NANDN U3090 ( .A(n2596), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n2610) );
  NANDN U3092 ( .A(n3170), .B(n3171), .Z(n2052) );
  AND U3093 ( .A(n3170), .B(n3168), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n3169), .Z(n2054) );
  NANDN U3095 ( .A(n3171), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n3185) );
  NANDN U3097 ( .A(n2825), .B(n2826), .Z(n2056) );
  AND U3098 ( .A(n2825), .B(n2823), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n2824), .Z(n2058) );
  NANDN U3100 ( .A(n2826), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n2840) );
  NANDN U3102 ( .A(n3400), .B(n3401), .Z(n2060) );
  AND U3103 ( .A(n3400), .B(n3398), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n3399), .Z(n2062) );
  NANDN U3105 ( .A(n3401), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n3415) );
  NANDN U3107 ( .A(n2480), .B(n2481), .Z(n2064) );
  AND U3108 ( .A(n2480), .B(n2478), .Z(n2065) );
  XNOR U3109 ( .A(n2065), .B(n2479), .Z(n2066) );
  NANDN U3110 ( .A(n2481), .B(n2066), .Z(n2067) );
  NAND U3111 ( .A(n2064), .B(n2067), .Z(n2495) );
  NANDN U3112 ( .A(n3614), .B(n3615), .Z(n2068) );
  AND U3113 ( .A(n3614), .B(n3612), .Z(n2069) );
  XNOR U3114 ( .A(n2069), .B(n3613), .Z(n2070) );
  NANDN U3115 ( .A(n3615), .B(n2070), .Z(n2071) );
  NAND U3116 ( .A(n2068), .B(n2071), .Z(n3629) );
  NANDN U3117 ( .A(n3055), .B(n3056), .Z(n2072) );
  AND U3118 ( .A(n3055), .B(n3053), .Z(n2073) );
  XNOR U3119 ( .A(n2073), .B(n3054), .Z(n2074) );
  NANDN U3120 ( .A(n3056), .B(n2074), .Z(n2075) );
  NAND U3121 ( .A(n2072), .B(n2075), .Z(n3070) );
  NANDN U3122 ( .A(n2365), .B(n2366), .Z(n2076) );
  AND U3123 ( .A(n2365), .B(n2363), .Z(n2077) );
  XNOR U3124 ( .A(n2077), .B(n2364), .Z(n2078) );
  NANDN U3125 ( .A(n2366), .B(n2078), .Z(n2079) );
  NAND U3126 ( .A(n2076), .B(n2079), .Z(n2380) );
  XOR U3127 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3128 ( .A(n2137), .B(n2138), .Z(n2080) );
  AND U3129 ( .A(n2137), .B(n2135), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2136), .Z(n2082) );
  NANDN U3131 ( .A(n2138), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2152) );
  NANDN U3133 ( .A(n3729), .B(n3730), .Z(n2084) );
  AND U3134 ( .A(n3729), .B(n3727), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3728), .Z(n2086) );
  NANDN U3136 ( .A(n3730), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3744) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_3 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U2967 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U2968 ( .A(n3911), .B(n3519), .Z(n3521) );
  XNOR U2969 ( .A(n2363), .B(n2361), .Z(n1966) );
  NANDN U2970 ( .A(n2366), .B(n1966), .Z(n1967) );
  NAND U2971 ( .A(n2366), .B(n2362), .Z(n1968) );
  NANDN U2972 ( .A(n2365), .B(n1968), .Z(n1969) );
  NAND U2973 ( .A(n1967), .B(n1969), .Z(n2421) );
  XNOR U2974 ( .A(n3053), .B(n3051), .Z(n1970) );
  NANDN U2975 ( .A(n3056), .B(n1970), .Z(n1971) );
  NAND U2976 ( .A(n3056), .B(n3052), .Z(n1972) );
  NANDN U2977 ( .A(n3055), .B(n1972), .Z(n1973) );
  NAND U2978 ( .A(n1971), .B(n1973), .Z(n3111) );
  XNOR U2979 ( .A(n3612), .B(n3610), .Z(n1974) );
  NANDN U2980 ( .A(n3615), .B(n1974), .Z(n1975) );
  NAND U2981 ( .A(n3615), .B(n3611), .Z(n1976) );
  NANDN U2982 ( .A(n3614), .B(n1976), .Z(n1977) );
  NAND U2983 ( .A(n1975), .B(n1977), .Z(n3670) );
  XNOR U2984 ( .A(n2938), .B(n2936), .Z(n1978) );
  NANDN U2985 ( .A(n2941), .B(n1978), .Z(n1979) );
  NAND U2986 ( .A(n2941), .B(n2937), .Z(n1980) );
  NANDN U2987 ( .A(n2940), .B(n1980), .Z(n1981) );
  NAND U2988 ( .A(n1979), .B(n1981), .Z(n2996) );
  AND U2989 ( .A(n3543), .B(n3528), .Z(n1982) );
  NAND U2990 ( .A(n3514), .B(n1982), .Z(n1983) );
  NANDN U2991 ( .A(n3528), .B(n3543), .Z(n1984) );
  XNOR U2992 ( .A(x[96]), .B(n1984), .Z(n1985) );
  NANDN U2993 ( .A(n3514), .B(n1985), .Z(n1986) );
  NAND U2994 ( .A(n1983), .B(n1986), .Z(n1987) );
  XNOR U2995 ( .A(n3469), .B(n3472), .Z(n1988) );
  XNOR U2996 ( .A(n1987), .B(n1988), .Z(n3497) );
  XNOR U2997 ( .A(n2823), .B(n2821), .Z(n1989) );
  NANDN U2998 ( .A(n2826), .B(n1989), .Z(n1990) );
  NAND U2999 ( .A(n2826), .B(n2822), .Z(n1991) );
  NANDN U3000 ( .A(n2825), .B(n1991), .Z(n1992) );
  NAND U3001 ( .A(n1990), .B(n1992), .Z(n2881) );
  XNOR U3002 ( .A(n3283), .B(n3281), .Z(n1993) );
  NANDN U3003 ( .A(n3286), .B(n1993), .Z(n1994) );
  NAND U3004 ( .A(n3286), .B(n3282), .Z(n1995) );
  NANDN U3005 ( .A(n3285), .B(n1995), .Z(n1996) );
  NAND U3006 ( .A(n1994), .B(n1996), .Z(n3341) );
  XNOR U3007 ( .A(n2135), .B(n2133), .Z(n1997) );
  NANDN U3008 ( .A(n2138), .B(n1997), .Z(n1998) );
  NAND U3009 ( .A(n2138), .B(n2134), .Z(n1999) );
  NANDN U3010 ( .A(n2137), .B(n1999), .Z(n2000) );
  NAND U3011 ( .A(n1998), .B(n2000), .Z(n2193) );
  XNOR U3012 ( .A(n3398), .B(n3396), .Z(n2001) );
  NANDN U3013 ( .A(n3401), .B(n2001), .Z(n2002) );
  NAND U3014 ( .A(n3401), .B(n3397), .Z(n2003) );
  NANDN U3015 ( .A(n3400), .B(n2003), .Z(n2004) );
  NAND U3016 ( .A(n2002), .B(n2004), .Z(n3456) );
  AND U3017 ( .A(n2297), .B(n2296), .Z(n2005) );
  XNOR U3018 ( .A(n2295), .B(n2005), .Z(n2309) );
  XNOR U3019 ( .A(n2478), .B(n2476), .Z(n2006) );
  NANDN U3020 ( .A(n2481), .B(n2006), .Z(n2007) );
  NAND U3021 ( .A(n2481), .B(n2477), .Z(n2008) );
  NANDN U3022 ( .A(n2480), .B(n2008), .Z(n2009) );
  NAND U3023 ( .A(n2007), .B(n2009), .Z(n2536) );
  XNOR U3024 ( .A(n2708), .B(n2706), .Z(n2010) );
  NANDN U3025 ( .A(n2711), .B(n2010), .Z(n2011) );
  NAND U3026 ( .A(n2711), .B(n2707), .Z(n2012) );
  NANDN U3027 ( .A(n2710), .B(n2012), .Z(n2013) );
  NAND U3028 ( .A(n2011), .B(n2013), .Z(n2766) );
  XNOR U3029 ( .A(n3842), .B(n3840), .Z(n2014) );
  NANDN U3030 ( .A(n3845), .B(n2014), .Z(n2015) );
  NAND U3031 ( .A(n3845), .B(n3841), .Z(n2016) );
  NANDN U3032 ( .A(n3844), .B(n2016), .Z(n2017) );
  NAND U3033 ( .A(n2015), .B(n2017), .Z(n3900) );
  NANDN U3034 ( .A(n3170), .B(n3171), .Z(n2018) );
  AND U3035 ( .A(n3170), .B(n3168), .Z(n2019) );
  XNOR U3036 ( .A(n2019), .B(n3169), .Z(n2020) );
  NANDN U3037 ( .A(n3171), .B(n2020), .Z(n2021) );
  NAND U3038 ( .A(n2018), .B(n2021), .Z(n3185) );
  XNOR U3039 ( .A(n3727), .B(n3725), .Z(n2022) );
  NANDN U3040 ( .A(n3730), .B(n2022), .Z(n2023) );
  NAND U3041 ( .A(n3730), .B(n3726), .Z(n2024) );
  NANDN U3042 ( .A(n3729), .B(n2024), .Z(n2025) );
  NAND U3043 ( .A(n2023), .B(n2025), .Z(n3785) );
  XNOR U3044 ( .A(n2593), .B(n2591), .Z(n2026) );
  NANDN U3045 ( .A(n2596), .B(n2026), .Z(n2027) );
  NAND U3046 ( .A(n2596), .B(n2592), .Z(n2028) );
  NANDN U3047 ( .A(n2595), .B(n2028), .Z(n2029) );
  NAND U3048 ( .A(n2027), .B(n2029), .Z(n2651) );
  ANDN U3049 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3050 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3051 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3052 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3053 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3054 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3055 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3056 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3057 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3058 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3059 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3060 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3061 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3062 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3063 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3064 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U3065 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3066 ( .A(n3771), .B(n3785), .Z(n3748) );
  NANDN U3067 ( .A(n3055), .B(n3056), .Z(n2032) );
  AND U3068 ( .A(n3055), .B(n3053), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n3054), .Z(n2034) );
  NANDN U3070 ( .A(n3056), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n3070) );
  NANDN U3072 ( .A(n2365), .B(n2366), .Z(n2036) );
  AND U3073 ( .A(n2365), .B(n2363), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n2364), .Z(n2038) );
  NANDN U3075 ( .A(n2366), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n2380) );
  NANDN U3077 ( .A(n2940), .B(n2941), .Z(n2040) );
  AND U3078 ( .A(n2940), .B(n2938), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n2939), .Z(n2042) );
  NANDN U3080 ( .A(n2941), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n2955) );
  NANDN U3082 ( .A(n2825), .B(n2826), .Z(n2044) );
  AND U3083 ( .A(n2825), .B(n2823), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n2824), .Z(n2046) );
  NANDN U3085 ( .A(n2826), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n2840) );
  NANDN U3087 ( .A(n2137), .B(n2138), .Z(n2048) );
  AND U3088 ( .A(n2137), .B(n2135), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n2136), .Z(n2050) );
  NANDN U3090 ( .A(n2138), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n2152) );
  NANDN U3092 ( .A(n3614), .B(n3615), .Z(n2052) );
  AND U3093 ( .A(n3614), .B(n3612), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n3613), .Z(n2054) );
  NANDN U3095 ( .A(n3615), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n3629) );
  NANDN U3097 ( .A(n3844), .B(n3845), .Z(n2056) );
  AND U3098 ( .A(n3844), .B(n3842), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n3843), .Z(n2058) );
  NANDN U3100 ( .A(n3845), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n3859) );
  NANDN U3102 ( .A(n3285), .B(n3286), .Z(n2060) );
  AND U3103 ( .A(n3285), .B(n3283), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n3284), .Z(n2062) );
  NANDN U3105 ( .A(n3286), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n3300) );
  NANDN U3107 ( .A(n3400), .B(n3401), .Z(n2064) );
  AND U3108 ( .A(n3400), .B(n3398), .Z(n2065) );
  XNOR U3109 ( .A(n2065), .B(n3399), .Z(n2066) );
  NANDN U3110 ( .A(n3401), .B(n2066), .Z(n2067) );
  NAND U3111 ( .A(n2064), .B(n2067), .Z(n3415) );
  XOR U3112 ( .A(n2283), .B(n2293), .Z(n3960) );
  XNOR U3113 ( .A(n3168), .B(n3166), .Z(n2068) );
  NANDN U3114 ( .A(n3171), .B(n2068), .Z(n2069) );
  NAND U3115 ( .A(n3171), .B(n3167), .Z(n2070) );
  NANDN U3116 ( .A(n3170), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2069), .B(n2071), .Z(n3226) );
  NANDN U3118 ( .A(n2595), .B(n2596), .Z(n2072) );
  AND U3119 ( .A(n2595), .B(n2593), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n2594), .Z(n2074) );
  NANDN U3121 ( .A(n2596), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n2610) );
  NANDN U3123 ( .A(n2480), .B(n2481), .Z(n2076) );
  AND U3124 ( .A(n2480), .B(n2478), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n2479), .Z(n2078) );
  NANDN U3126 ( .A(n2481), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n2495) );
  NANDN U3128 ( .A(n2710), .B(n2711), .Z(n2080) );
  AND U3129 ( .A(n2710), .B(n2708), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2709), .Z(n2082) );
  NANDN U3131 ( .A(n2711), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2725) );
  NANDN U3133 ( .A(n3729), .B(n3730), .Z(n2084) );
  AND U3134 ( .A(n3729), .B(n3727), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3728), .Z(n2086) );
  NANDN U3136 ( .A(n3730), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3744) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_4 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3912), .B(n3520), .Z(n3530) );
  AND U2967 ( .A(n2297), .B(n2296), .Z(n1966) );
  XNOR U2968 ( .A(n2295), .B(n1966), .Z(n2309) );
  XOR U2969 ( .A(n3911), .B(n3519), .Z(n3521) );
  XNOR U2970 ( .A(n3398), .B(n3396), .Z(n1967) );
  NANDN U2971 ( .A(n3401), .B(n1967), .Z(n1968) );
  NAND U2972 ( .A(n3401), .B(n3397), .Z(n1969) );
  NANDN U2973 ( .A(n3400), .B(n1969), .Z(n1970) );
  NAND U2974 ( .A(n1968), .B(n1970), .Z(n3456) );
  AND U2975 ( .A(n3543), .B(n3528), .Z(n1971) );
  NAND U2976 ( .A(n3514), .B(n1971), .Z(n1972) );
  NANDN U2977 ( .A(n3528), .B(n3543), .Z(n1973) );
  XNOR U2978 ( .A(x[96]), .B(n1973), .Z(n1974) );
  NANDN U2979 ( .A(n3514), .B(n1974), .Z(n1975) );
  NAND U2980 ( .A(n1972), .B(n1975), .Z(n1976) );
  XNOR U2981 ( .A(n3469), .B(n3472), .Z(n1977) );
  XNOR U2982 ( .A(n1976), .B(n1977), .Z(n3497) );
  XNOR U2983 ( .A(n2823), .B(n2821), .Z(n1978) );
  NANDN U2984 ( .A(n2826), .B(n1978), .Z(n1979) );
  NAND U2985 ( .A(n2826), .B(n2822), .Z(n1980) );
  NANDN U2986 ( .A(n2825), .B(n1980), .Z(n1981) );
  NAND U2987 ( .A(n1979), .B(n1981), .Z(n2881) );
  XOR U2988 ( .A(n3886), .B(n3900), .Z(n3863) );
  XNOR U2989 ( .A(n3283), .B(n3281), .Z(n1982) );
  NANDN U2990 ( .A(n3286), .B(n1982), .Z(n1983) );
  NAND U2991 ( .A(n3286), .B(n3282), .Z(n1984) );
  NANDN U2992 ( .A(n3285), .B(n1984), .Z(n1985) );
  NAND U2993 ( .A(n1983), .B(n1985), .Z(n3341) );
  XNOR U2994 ( .A(n2135), .B(n2133), .Z(n1986) );
  NANDN U2995 ( .A(n2138), .B(n1986), .Z(n1987) );
  NAND U2996 ( .A(n2138), .B(n2134), .Z(n1988) );
  NANDN U2997 ( .A(n2137), .B(n1988), .Z(n1989) );
  NAND U2998 ( .A(n1987), .B(n1989), .Z(n2193) );
  XNOR U2999 ( .A(n2938), .B(n2936), .Z(n1990) );
  NANDN U3000 ( .A(n2941), .B(n1990), .Z(n1991) );
  NAND U3001 ( .A(n2941), .B(n2937), .Z(n1992) );
  NANDN U3002 ( .A(n2940), .B(n1992), .Z(n1993) );
  NAND U3003 ( .A(n1991), .B(n1993), .Z(n2996) );
  XNOR U3004 ( .A(n2478), .B(n2476), .Z(n1994) );
  NANDN U3005 ( .A(n2481), .B(n1994), .Z(n1995) );
  NAND U3006 ( .A(n2481), .B(n2477), .Z(n1996) );
  NANDN U3007 ( .A(n2480), .B(n1996), .Z(n1997) );
  NAND U3008 ( .A(n1995), .B(n1997), .Z(n2536) );
  XNOR U3009 ( .A(n3727), .B(n3725), .Z(n1998) );
  NANDN U3010 ( .A(n3730), .B(n1998), .Z(n1999) );
  NAND U3011 ( .A(n3730), .B(n3726), .Z(n2000) );
  NANDN U3012 ( .A(n3729), .B(n2000), .Z(n2001) );
  NAND U3013 ( .A(n1999), .B(n2001), .Z(n3785) );
  XNOR U3014 ( .A(n3168), .B(n3166), .Z(n2002) );
  NANDN U3015 ( .A(n3171), .B(n2002), .Z(n2003) );
  NAND U3016 ( .A(n3171), .B(n3167), .Z(n2004) );
  NANDN U3017 ( .A(n3170), .B(n2004), .Z(n2005) );
  NAND U3018 ( .A(n2003), .B(n2005), .Z(n3226) );
  XNOR U3019 ( .A(n2593), .B(n2591), .Z(n2006) );
  NANDN U3020 ( .A(n2596), .B(n2006), .Z(n2007) );
  NAND U3021 ( .A(n2596), .B(n2592), .Z(n2008) );
  NANDN U3022 ( .A(n2595), .B(n2008), .Z(n2009) );
  NAND U3023 ( .A(n2007), .B(n2009), .Z(n2651) );
  XNOR U3024 ( .A(n3612), .B(n3610), .Z(n2010) );
  NANDN U3025 ( .A(n3615), .B(n2010), .Z(n2011) );
  NAND U3026 ( .A(n3615), .B(n3611), .Z(n2012) );
  NANDN U3027 ( .A(n3614), .B(n2012), .Z(n2013) );
  NAND U3028 ( .A(n2011), .B(n2013), .Z(n3670) );
  XNOR U3029 ( .A(n2363), .B(n2361), .Z(n2014) );
  NANDN U3030 ( .A(n2366), .B(n2014), .Z(n2015) );
  NAND U3031 ( .A(n2366), .B(n2362), .Z(n2016) );
  NANDN U3032 ( .A(n2365), .B(n2016), .Z(n2017) );
  NAND U3033 ( .A(n2015), .B(n2017), .Z(n2421) );
  XNOR U3034 ( .A(n3053), .B(n3051), .Z(n2018) );
  NANDN U3035 ( .A(n3056), .B(n2018), .Z(n2019) );
  NAND U3036 ( .A(n3056), .B(n3052), .Z(n2020) );
  NANDN U3037 ( .A(n3055), .B(n2020), .Z(n2021) );
  NAND U3038 ( .A(n2019), .B(n2021), .Z(n3111) );
  XNOR U3039 ( .A(n2708), .B(n2706), .Z(n2022) );
  NANDN U3040 ( .A(n2711), .B(n2022), .Z(n2023) );
  NAND U3041 ( .A(n2711), .B(n2707), .Z(n2024) );
  NANDN U3042 ( .A(n2710), .B(n2024), .Z(n2025) );
  NAND U3043 ( .A(n2023), .B(n2025), .Z(n2766) );
  NANDN U3044 ( .A(n3844), .B(n3845), .Z(n2026) );
  AND U3045 ( .A(n3844), .B(n3842), .Z(n2027) );
  XNOR U3046 ( .A(n2027), .B(n3843), .Z(n2028) );
  NANDN U3047 ( .A(n3845), .B(n2028), .Z(n2029) );
  NAND U3048 ( .A(n2026), .B(n2029), .Z(n3859) );
  XOR U3049 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3050 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3051 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3052 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3053 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3054 ( .A(n3327), .B(n3341), .Z(n3304) );
  ANDN U3055 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3056 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3057 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3058 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3059 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3060 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3061 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3062 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3063 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3064 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3065 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U3066 ( .A(n2752), .B(n2766), .Z(n2729) );
  NANDN U3067 ( .A(n3170), .B(n3171), .Z(n2032) );
  AND U3068 ( .A(n3170), .B(n3168), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n3169), .Z(n2034) );
  NANDN U3070 ( .A(n3171), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n3185) );
  XOR U3072 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3073 ( .A(n3400), .B(n3401), .Z(n2036) );
  AND U3074 ( .A(n3400), .B(n3398), .Z(n2037) );
  XNOR U3075 ( .A(n2037), .B(n3399), .Z(n2038) );
  NANDN U3076 ( .A(n3401), .B(n2038), .Z(n2039) );
  NAND U3077 ( .A(n2036), .B(n2039), .Z(n3415) );
  NANDN U3078 ( .A(n2825), .B(n2826), .Z(n2040) );
  AND U3079 ( .A(n2825), .B(n2823), .Z(n2041) );
  XNOR U3080 ( .A(n2041), .B(n2824), .Z(n2042) );
  NANDN U3081 ( .A(n2826), .B(n2042), .Z(n2043) );
  NAND U3082 ( .A(n2040), .B(n2043), .Z(n2840) );
  NANDN U3083 ( .A(n3285), .B(n3286), .Z(n2044) );
  AND U3084 ( .A(n3285), .B(n3283), .Z(n2045) );
  XNOR U3085 ( .A(n2045), .B(n3284), .Z(n2046) );
  NANDN U3086 ( .A(n3286), .B(n2046), .Z(n2047) );
  NAND U3087 ( .A(n2044), .B(n2047), .Z(n3300) );
  NANDN U3088 ( .A(n2137), .B(n2138), .Z(n2048) );
  AND U3089 ( .A(n2137), .B(n2135), .Z(n2049) );
  XNOR U3090 ( .A(n2049), .B(n2136), .Z(n2050) );
  NANDN U3091 ( .A(n2138), .B(n2050), .Z(n2051) );
  NAND U3092 ( .A(n2048), .B(n2051), .Z(n2152) );
  XNOR U3093 ( .A(n3842), .B(n3840), .Z(n2052) );
  NANDN U3094 ( .A(n3845), .B(n2052), .Z(n2053) );
  NAND U3095 ( .A(n3845), .B(n3841), .Z(n2054) );
  NANDN U3096 ( .A(n3844), .B(n2054), .Z(n2055) );
  NAND U3097 ( .A(n2053), .B(n2055), .Z(n3900) );
  NANDN U3098 ( .A(n2940), .B(n2941), .Z(n2056) );
  AND U3099 ( .A(n2940), .B(n2938), .Z(n2057) );
  XNOR U3100 ( .A(n2057), .B(n2939), .Z(n2058) );
  NANDN U3101 ( .A(n2941), .B(n2058), .Z(n2059) );
  NAND U3102 ( .A(n2056), .B(n2059), .Z(n2955) );
  NANDN U3103 ( .A(n2480), .B(n2481), .Z(n2060) );
  AND U3104 ( .A(n2480), .B(n2478), .Z(n2061) );
  XNOR U3105 ( .A(n2061), .B(n2479), .Z(n2062) );
  NANDN U3106 ( .A(n2481), .B(n2062), .Z(n2063) );
  NAND U3107 ( .A(n2060), .B(n2063), .Z(n2495) );
  NANDN U3108 ( .A(n2595), .B(n2596), .Z(n2064) );
  AND U3109 ( .A(n2595), .B(n2593), .Z(n2065) );
  XNOR U3110 ( .A(n2065), .B(n2594), .Z(n2066) );
  NANDN U3111 ( .A(n2596), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2064), .B(n2067), .Z(n2610) );
  NANDN U3113 ( .A(n3729), .B(n3730), .Z(n2068) );
  AND U3114 ( .A(n3729), .B(n3727), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n3728), .Z(n2070) );
  NANDN U3116 ( .A(n3730), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n3744) );
  NANDN U3118 ( .A(n3614), .B(n3615), .Z(n2072) );
  AND U3119 ( .A(n3614), .B(n3612), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n3613), .Z(n2074) );
  NANDN U3121 ( .A(n3615), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n3629) );
  NANDN U3123 ( .A(n3055), .B(n3056), .Z(n2076) );
  AND U3124 ( .A(n3055), .B(n3053), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3054), .Z(n2078) );
  NANDN U3126 ( .A(n3056), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3070) );
  NANDN U3128 ( .A(n2365), .B(n2366), .Z(n2080) );
  AND U3129 ( .A(n2365), .B(n2363), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2364), .Z(n2082) );
  NANDN U3131 ( .A(n2366), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2380) );
  NANDN U3133 ( .A(n2710), .B(n2711), .Z(n2084) );
  AND U3134 ( .A(n2710), .B(n2708), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n2709), .Z(n2086) );
  NANDN U3136 ( .A(n2711), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n2725) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_5 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U2967 ( .A(n3911), .B(n3519), .Z(n3521) );
  AND U2968 ( .A(n3543), .B(n3528), .Z(n1966) );
  NAND U2969 ( .A(n3514), .B(n1966), .Z(n1967) );
  NANDN U2970 ( .A(n3528), .B(n3543), .Z(n1968) );
  XNOR U2971 ( .A(x[96]), .B(n1968), .Z(n1969) );
  NANDN U2972 ( .A(n3514), .B(n1969), .Z(n1970) );
  NAND U2973 ( .A(n1967), .B(n1970), .Z(n1971) );
  XNOR U2974 ( .A(n3469), .B(n3472), .Z(n1972) );
  XNOR U2975 ( .A(n1971), .B(n1972), .Z(n3497) );
  XNOR U2976 ( .A(n2823), .B(n2821), .Z(n1973) );
  NANDN U2977 ( .A(n2826), .B(n1973), .Z(n1974) );
  NAND U2978 ( .A(n2826), .B(n2822), .Z(n1975) );
  NANDN U2979 ( .A(n2825), .B(n1975), .Z(n1976) );
  NAND U2980 ( .A(n1974), .B(n1976), .Z(n2881) );
  XNOR U2981 ( .A(n2938), .B(n2936), .Z(n1977) );
  NANDN U2982 ( .A(n2941), .B(n1977), .Z(n1978) );
  NAND U2983 ( .A(n2941), .B(n2937), .Z(n1979) );
  NANDN U2984 ( .A(n2940), .B(n1979), .Z(n1980) );
  NAND U2985 ( .A(n1978), .B(n1980), .Z(n2996) );
  XNOR U2986 ( .A(n2708), .B(n2706), .Z(n1981) );
  NANDN U2987 ( .A(n2711), .B(n1981), .Z(n1982) );
  NAND U2988 ( .A(n2711), .B(n2707), .Z(n1983) );
  NANDN U2989 ( .A(n2710), .B(n1983), .Z(n1984) );
  NAND U2990 ( .A(n1982), .B(n1984), .Z(n2766) );
  XNOR U2991 ( .A(n3398), .B(n3396), .Z(n1985) );
  NANDN U2992 ( .A(n3401), .B(n1985), .Z(n1986) );
  NAND U2993 ( .A(n3401), .B(n3397), .Z(n1987) );
  NANDN U2994 ( .A(n3400), .B(n1987), .Z(n1988) );
  NAND U2995 ( .A(n1986), .B(n1988), .Z(n3456) );
  AND U2996 ( .A(n2297), .B(n2296), .Z(n1989) );
  XNOR U2997 ( .A(n2295), .B(n1989), .Z(n2309) );
  XNOR U2998 ( .A(n2478), .B(n2476), .Z(n1990) );
  NANDN U2999 ( .A(n2481), .B(n1990), .Z(n1991) );
  NAND U3000 ( .A(n2481), .B(n2477), .Z(n1992) );
  NANDN U3001 ( .A(n2480), .B(n1992), .Z(n1993) );
  NAND U3002 ( .A(n1991), .B(n1993), .Z(n2536) );
  XNOR U3003 ( .A(n3168), .B(n3166), .Z(n1994) );
  NANDN U3004 ( .A(n3171), .B(n1994), .Z(n1995) );
  NAND U3005 ( .A(n3171), .B(n3167), .Z(n1996) );
  NANDN U3006 ( .A(n3170), .B(n1996), .Z(n1997) );
  NAND U3007 ( .A(n1995), .B(n1997), .Z(n3226) );
  XNOR U3008 ( .A(n3727), .B(n3725), .Z(n1998) );
  NANDN U3009 ( .A(n3730), .B(n1998), .Z(n1999) );
  NAND U3010 ( .A(n3730), .B(n3726), .Z(n2000) );
  NANDN U3011 ( .A(n3729), .B(n2000), .Z(n2001) );
  NAND U3012 ( .A(n1999), .B(n2001), .Z(n3785) );
  XNOR U3013 ( .A(n2593), .B(n2591), .Z(n2002) );
  NANDN U3014 ( .A(n2596), .B(n2002), .Z(n2003) );
  NAND U3015 ( .A(n2596), .B(n2592), .Z(n2004) );
  NANDN U3016 ( .A(n2595), .B(n2004), .Z(n2005) );
  NAND U3017 ( .A(n2003), .B(n2005), .Z(n2651) );
  XNOR U3018 ( .A(n3283), .B(n3281), .Z(n2006) );
  NANDN U3019 ( .A(n3286), .B(n2006), .Z(n2007) );
  NAND U3020 ( .A(n3286), .B(n3282), .Z(n2008) );
  NANDN U3021 ( .A(n3285), .B(n2008), .Z(n2009) );
  NAND U3022 ( .A(n2007), .B(n2009), .Z(n3341) );
  XNOR U3023 ( .A(n3842), .B(n3840), .Z(n2010) );
  NANDN U3024 ( .A(n3845), .B(n2010), .Z(n2011) );
  NAND U3025 ( .A(n3845), .B(n3841), .Z(n2012) );
  NANDN U3026 ( .A(n3844), .B(n2012), .Z(n2013) );
  NAND U3027 ( .A(n2011), .B(n2013), .Z(n3900) );
  XNOR U3028 ( .A(n2135), .B(n2133), .Z(n2014) );
  NANDN U3029 ( .A(n2138), .B(n2014), .Z(n2015) );
  NAND U3030 ( .A(n2138), .B(n2134), .Z(n2016) );
  NANDN U3031 ( .A(n2137), .B(n2016), .Z(n2017) );
  NAND U3032 ( .A(n2015), .B(n2017), .Z(n2193) );
  XNOR U3033 ( .A(n3612), .B(n3610), .Z(n2018) );
  NANDN U3034 ( .A(n3615), .B(n2018), .Z(n2019) );
  NAND U3035 ( .A(n3615), .B(n3611), .Z(n2020) );
  NANDN U3036 ( .A(n3614), .B(n2020), .Z(n2021) );
  NAND U3037 ( .A(n2019), .B(n2021), .Z(n3670) );
  XNOR U3038 ( .A(n2363), .B(n2361), .Z(n2022) );
  NANDN U3039 ( .A(n2366), .B(n2022), .Z(n2023) );
  NAND U3040 ( .A(n2366), .B(n2362), .Z(n2024) );
  NANDN U3041 ( .A(n2365), .B(n2024), .Z(n2025) );
  NAND U3042 ( .A(n2023), .B(n2025), .Z(n2421) );
  XNOR U3043 ( .A(n3053), .B(n3051), .Z(n2026) );
  NANDN U3044 ( .A(n3056), .B(n2026), .Z(n2027) );
  NAND U3045 ( .A(n3056), .B(n3052), .Z(n2028) );
  NANDN U3046 ( .A(n3055), .B(n2028), .Z(n2029) );
  NAND U3047 ( .A(n2027), .B(n2029), .Z(n3111) );
  XOR U3048 ( .A(n2867), .B(n2881), .Z(n2844) );
  ANDN U3049 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3050 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3051 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3052 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3053 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3054 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3055 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3056 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3057 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3058 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3059 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3060 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3061 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3062 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U3063 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3064 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3065 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3066 ( .A(n2407), .B(n2421), .Z(n2384) );
  NANDN U3067 ( .A(n2825), .B(n2826), .Z(n2032) );
  AND U3068 ( .A(n2825), .B(n2823), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n2824), .Z(n2034) );
  NANDN U3070 ( .A(n2826), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n2840) );
  NANDN U3072 ( .A(n3844), .B(n3845), .Z(n2036) );
  AND U3073 ( .A(n3844), .B(n3842), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n3843), .Z(n2038) );
  NANDN U3075 ( .A(n3845), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n3859) );
  NANDN U3077 ( .A(n2480), .B(n2481), .Z(n2040) );
  AND U3078 ( .A(n2480), .B(n2478), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n2479), .Z(n2042) );
  NANDN U3080 ( .A(n2481), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n2495) );
  NANDN U3082 ( .A(n2595), .B(n2596), .Z(n2044) );
  AND U3083 ( .A(n2595), .B(n2593), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n2594), .Z(n2046) );
  NANDN U3085 ( .A(n2596), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n2610) );
  NANDN U3087 ( .A(n2940), .B(n2941), .Z(n2048) );
  AND U3088 ( .A(n2940), .B(n2938), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n2939), .Z(n2050) );
  NANDN U3090 ( .A(n2941), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n2955) );
  NANDN U3092 ( .A(n2710), .B(n2711), .Z(n2052) );
  AND U3093 ( .A(n2710), .B(n2708), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n2709), .Z(n2054) );
  NANDN U3095 ( .A(n2711), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n2725) );
  NANDN U3097 ( .A(n3285), .B(n3286), .Z(n2056) );
  AND U3098 ( .A(n3285), .B(n3283), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n3284), .Z(n2058) );
  NANDN U3100 ( .A(n3286), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n3300) );
  NANDN U3102 ( .A(n3400), .B(n3401), .Z(n2060) );
  AND U3103 ( .A(n3400), .B(n3398), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n3399), .Z(n2062) );
  NANDN U3105 ( .A(n3401), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n3415) );
  XOR U3107 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3108 ( .A(n3170), .B(n3171), .Z(n2064) );
  AND U3109 ( .A(n3170), .B(n3168), .Z(n2065) );
  XNOR U3110 ( .A(n2065), .B(n3169), .Z(n2066) );
  NANDN U3111 ( .A(n3171), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2064), .B(n2067), .Z(n3185) );
  NANDN U3113 ( .A(n3729), .B(n3730), .Z(n2068) );
  AND U3114 ( .A(n3729), .B(n3727), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n3728), .Z(n2070) );
  NANDN U3116 ( .A(n3730), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n3744) );
  NANDN U3118 ( .A(n2137), .B(n2138), .Z(n2072) );
  AND U3119 ( .A(n2137), .B(n2135), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n2136), .Z(n2074) );
  NANDN U3121 ( .A(n2138), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n2152) );
  NANDN U3123 ( .A(n3614), .B(n3615), .Z(n2076) );
  AND U3124 ( .A(n3614), .B(n3612), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3613), .Z(n2078) );
  NANDN U3126 ( .A(n3615), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3629) );
  NANDN U3128 ( .A(n3055), .B(n3056), .Z(n2080) );
  AND U3129 ( .A(n3055), .B(n3053), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n3054), .Z(n2082) );
  NANDN U3131 ( .A(n3056), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n3070) );
  NANDN U3133 ( .A(n2365), .B(n2366), .Z(n2084) );
  AND U3134 ( .A(n2365), .B(n2363), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n2364), .Z(n2086) );
  NANDN U3136 ( .A(n2366), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n2380) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_6 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3912), .B(n3520), .Z(n3530) );
  XNOR U2967 ( .A(n2938), .B(n2936), .Z(n1966) );
  NANDN U2968 ( .A(n2941), .B(n1966), .Z(n1967) );
  NAND U2969 ( .A(n2941), .B(n2937), .Z(n1968) );
  NANDN U2970 ( .A(n2940), .B(n1968), .Z(n1969) );
  NAND U2971 ( .A(n1967), .B(n1969), .Z(n2996) );
  XNOR U2972 ( .A(n3612), .B(n3610), .Z(n1970) );
  NANDN U2973 ( .A(n3615), .B(n1970), .Z(n1971) );
  NAND U2974 ( .A(n3615), .B(n3611), .Z(n1972) );
  NANDN U2975 ( .A(n3614), .B(n1972), .Z(n1973) );
  NAND U2976 ( .A(n1971), .B(n1973), .Z(n3670) );
  XNOR U2977 ( .A(n2363), .B(n2361), .Z(n1974) );
  NANDN U2978 ( .A(n2366), .B(n1974), .Z(n1975) );
  NAND U2979 ( .A(n2366), .B(n2362), .Z(n1976) );
  NANDN U2980 ( .A(n2365), .B(n1976), .Z(n1977) );
  NAND U2981 ( .A(n1975), .B(n1977), .Z(n2421) );
  XNOR U2982 ( .A(n3053), .B(n3051), .Z(n1978) );
  NANDN U2983 ( .A(n3056), .B(n1978), .Z(n1979) );
  NAND U2984 ( .A(n3056), .B(n3052), .Z(n1980) );
  NANDN U2985 ( .A(n3055), .B(n1980), .Z(n1981) );
  NAND U2986 ( .A(n1979), .B(n1981), .Z(n3111) );
  XOR U2987 ( .A(n3911), .B(n3519), .Z(n3521) );
  AND U2988 ( .A(n3543), .B(n3528), .Z(n1982) );
  NAND U2989 ( .A(n3514), .B(n1982), .Z(n1983) );
  NANDN U2990 ( .A(n3528), .B(n3543), .Z(n1984) );
  XNOR U2991 ( .A(x[96]), .B(n1984), .Z(n1985) );
  NANDN U2992 ( .A(n3514), .B(n1985), .Z(n1986) );
  NAND U2993 ( .A(n1983), .B(n1986), .Z(n1987) );
  XNOR U2994 ( .A(n3469), .B(n3472), .Z(n1988) );
  XNOR U2995 ( .A(n1987), .B(n1988), .Z(n3497) );
  XNOR U2996 ( .A(n2823), .B(n2821), .Z(n1989) );
  NANDN U2997 ( .A(n2826), .B(n1989), .Z(n1990) );
  NAND U2998 ( .A(n2826), .B(n2822), .Z(n1991) );
  NANDN U2999 ( .A(n2825), .B(n1991), .Z(n1992) );
  NAND U3000 ( .A(n1990), .B(n1992), .Z(n2881) );
  XNOR U3001 ( .A(n3842), .B(n3840), .Z(n1993) );
  NANDN U3002 ( .A(n3845), .B(n1993), .Z(n1994) );
  NAND U3003 ( .A(n3845), .B(n3841), .Z(n1995) );
  NANDN U3004 ( .A(n3844), .B(n1995), .Z(n1996) );
  NAND U3005 ( .A(n1994), .B(n1996), .Z(n3900) );
  XNOR U3006 ( .A(n2593), .B(n2591), .Z(n1997) );
  NANDN U3007 ( .A(n2596), .B(n1997), .Z(n1998) );
  NAND U3008 ( .A(n2596), .B(n2592), .Z(n1999) );
  NANDN U3009 ( .A(n2595), .B(n1999), .Z(n2000) );
  NAND U3010 ( .A(n1998), .B(n2000), .Z(n2651) );
  XNOR U3011 ( .A(n3727), .B(n3725), .Z(n2001) );
  NANDN U3012 ( .A(n3730), .B(n2001), .Z(n2002) );
  NAND U3013 ( .A(n3730), .B(n3726), .Z(n2003) );
  NANDN U3014 ( .A(n3729), .B(n2003), .Z(n2004) );
  NAND U3015 ( .A(n2002), .B(n2004), .Z(n3785) );
  XNOR U3016 ( .A(n2708), .B(n2706), .Z(n2005) );
  NANDN U3017 ( .A(n2711), .B(n2005), .Z(n2006) );
  NAND U3018 ( .A(n2711), .B(n2707), .Z(n2007) );
  NANDN U3019 ( .A(n2710), .B(n2007), .Z(n2008) );
  NAND U3020 ( .A(n2006), .B(n2008), .Z(n2766) );
  XNOR U3021 ( .A(n3283), .B(n3281), .Z(n2009) );
  NANDN U3022 ( .A(n3286), .B(n2009), .Z(n2010) );
  NAND U3023 ( .A(n3286), .B(n3282), .Z(n2011) );
  NANDN U3024 ( .A(n3285), .B(n2011), .Z(n2012) );
  NAND U3025 ( .A(n2010), .B(n2012), .Z(n3341) );
  XNOR U3026 ( .A(n2135), .B(n2133), .Z(n2013) );
  NANDN U3027 ( .A(n2138), .B(n2013), .Z(n2014) );
  NAND U3028 ( .A(n2138), .B(n2134), .Z(n2015) );
  NANDN U3029 ( .A(n2137), .B(n2015), .Z(n2016) );
  NAND U3030 ( .A(n2014), .B(n2016), .Z(n2193) );
  XNOR U3031 ( .A(n3398), .B(n3396), .Z(n2017) );
  NANDN U3032 ( .A(n3401), .B(n2017), .Z(n2018) );
  NAND U3033 ( .A(n3401), .B(n3397), .Z(n2019) );
  NANDN U3034 ( .A(n3400), .B(n2019), .Z(n2020) );
  NAND U3035 ( .A(n2018), .B(n2020), .Z(n3456) );
  AND U3036 ( .A(n2297), .B(n2296), .Z(n2021) );
  XNOR U3037 ( .A(n2295), .B(n2021), .Z(n2309) );
  XNOR U3038 ( .A(n2478), .B(n2476), .Z(n2022) );
  NANDN U3039 ( .A(n2481), .B(n2022), .Z(n2023) );
  NAND U3040 ( .A(n2481), .B(n2477), .Z(n2024) );
  NANDN U3041 ( .A(n2480), .B(n2024), .Z(n2025) );
  NAND U3042 ( .A(n2023), .B(n2025), .Z(n2536) );
  XNOR U3043 ( .A(n3168), .B(n3166), .Z(n2026) );
  NANDN U3044 ( .A(n3171), .B(n2026), .Z(n2027) );
  NAND U3045 ( .A(n3171), .B(n3167), .Z(n2028) );
  NANDN U3046 ( .A(n3170), .B(n2028), .Z(n2029) );
  NAND U3047 ( .A(n2027), .B(n2029), .Z(n3226) );
  XOR U3048 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3049 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3050 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3051 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3052 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3053 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3054 ( .A(n2407), .B(n2421), .Z(n2384) );
  ANDN U3055 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3056 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3057 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3058 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3059 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3060 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3061 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3062 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3063 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3064 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3065 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3066 ( .A(n3544), .B(n3555), .Z(n3542) );
  NANDN U3067 ( .A(n3844), .B(n3845), .Z(n2032) );
  AND U3068 ( .A(n3844), .B(n3842), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n3843), .Z(n2034) );
  NANDN U3070 ( .A(n3845), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n3859) );
  NANDN U3072 ( .A(n2595), .B(n2596), .Z(n2036) );
  AND U3073 ( .A(n2595), .B(n2593), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n2594), .Z(n2038) );
  NANDN U3075 ( .A(n2596), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n2610) );
  NANDN U3077 ( .A(n2940), .B(n2941), .Z(n2040) );
  AND U3078 ( .A(n2940), .B(n2938), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n2939), .Z(n2042) );
  NANDN U3080 ( .A(n2941), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n2955) );
  NANDN U3082 ( .A(n2137), .B(n2138), .Z(n2044) );
  AND U3083 ( .A(n2137), .B(n2135), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n2136), .Z(n2046) );
  NANDN U3085 ( .A(n2138), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n2152) );
  NANDN U3087 ( .A(n3055), .B(n3056), .Z(n2048) );
  AND U3088 ( .A(n3055), .B(n3053), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n3054), .Z(n2050) );
  NANDN U3090 ( .A(n3056), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n3070) );
  NANDN U3092 ( .A(n3614), .B(n3615), .Z(n2052) );
  AND U3093 ( .A(n3614), .B(n3612), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n3613), .Z(n2054) );
  NANDN U3095 ( .A(n3615), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n3629) );
  NANDN U3097 ( .A(n2365), .B(n2366), .Z(n2056) );
  AND U3098 ( .A(n2365), .B(n2363), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n2364), .Z(n2058) );
  NANDN U3100 ( .A(n2366), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n2380) );
  NANDN U3102 ( .A(n2825), .B(n2826), .Z(n2060) );
  AND U3103 ( .A(n2825), .B(n2823), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n2824), .Z(n2062) );
  NANDN U3105 ( .A(n2826), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n2840) );
  NANDN U3107 ( .A(n2710), .B(n2711), .Z(n2064) );
  AND U3108 ( .A(n2710), .B(n2708), .Z(n2065) );
  XNOR U3109 ( .A(n2065), .B(n2709), .Z(n2066) );
  NANDN U3110 ( .A(n2711), .B(n2066), .Z(n2067) );
  NAND U3111 ( .A(n2064), .B(n2067), .Z(n2725) );
  NANDN U3112 ( .A(n2480), .B(n2481), .Z(n2068) );
  AND U3113 ( .A(n2480), .B(n2478), .Z(n2069) );
  XNOR U3114 ( .A(n2069), .B(n2479), .Z(n2070) );
  NANDN U3115 ( .A(n2481), .B(n2070), .Z(n2071) );
  NAND U3116 ( .A(n2068), .B(n2071), .Z(n2495) );
  NANDN U3117 ( .A(n3729), .B(n3730), .Z(n2072) );
  AND U3118 ( .A(n3729), .B(n3727), .Z(n2073) );
  XNOR U3119 ( .A(n2073), .B(n3728), .Z(n2074) );
  NANDN U3120 ( .A(n3730), .B(n2074), .Z(n2075) );
  NAND U3121 ( .A(n2072), .B(n2075), .Z(n3744) );
  NANDN U3122 ( .A(n3285), .B(n3286), .Z(n2076) );
  AND U3123 ( .A(n3285), .B(n3283), .Z(n2077) );
  XNOR U3124 ( .A(n2077), .B(n3284), .Z(n2078) );
  NANDN U3125 ( .A(n3286), .B(n2078), .Z(n2079) );
  NAND U3126 ( .A(n2076), .B(n2079), .Z(n3300) );
  NANDN U3127 ( .A(n3400), .B(n3401), .Z(n2080) );
  AND U3128 ( .A(n3400), .B(n3398), .Z(n2081) );
  XNOR U3129 ( .A(n2081), .B(n3399), .Z(n2082) );
  NANDN U3130 ( .A(n3401), .B(n2082), .Z(n2083) );
  NAND U3131 ( .A(n2080), .B(n2083), .Z(n3415) );
  XOR U3132 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3133 ( .A(n3170), .B(n3171), .Z(n2084) );
  AND U3134 ( .A(n3170), .B(n3168), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3169), .Z(n2086) );
  NANDN U3136 ( .A(n3171), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3185) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_7 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U2967 ( .A(n3212), .B(n3226), .Z(n3189) );
  XNOR U2968 ( .A(n3283), .B(n3281), .Z(n1966) );
  NANDN U2969 ( .A(n3286), .B(n1966), .Z(n1967) );
  NAND U2970 ( .A(n3286), .B(n3282), .Z(n1968) );
  NANDN U2971 ( .A(n3285), .B(n1968), .Z(n1969) );
  NAND U2972 ( .A(n1967), .B(n1969), .Z(n3341) );
  XNOR U2973 ( .A(n2135), .B(n2133), .Z(n1970) );
  NANDN U2974 ( .A(n2138), .B(n1970), .Z(n1971) );
  NAND U2975 ( .A(n2138), .B(n2134), .Z(n1972) );
  NANDN U2976 ( .A(n2137), .B(n1972), .Z(n1973) );
  NAND U2977 ( .A(n1971), .B(n1973), .Z(n2193) );
  XNOR U2978 ( .A(n2938), .B(n2936), .Z(n1974) );
  NANDN U2979 ( .A(n2941), .B(n1974), .Z(n1975) );
  NAND U2980 ( .A(n2941), .B(n2937), .Z(n1976) );
  NANDN U2981 ( .A(n2940), .B(n1976), .Z(n1977) );
  NAND U2982 ( .A(n1975), .B(n1977), .Z(n2996) );
  XNOR U2983 ( .A(n3612), .B(n3610), .Z(n1978) );
  NANDN U2984 ( .A(n3615), .B(n1978), .Z(n1979) );
  NAND U2985 ( .A(n3615), .B(n3611), .Z(n1980) );
  NANDN U2986 ( .A(n3614), .B(n1980), .Z(n1981) );
  NAND U2987 ( .A(n1979), .B(n1981), .Z(n3670) );
  XNOR U2988 ( .A(n2363), .B(n2361), .Z(n1982) );
  NANDN U2989 ( .A(n2366), .B(n1982), .Z(n1983) );
  NAND U2990 ( .A(n2366), .B(n2362), .Z(n1984) );
  NANDN U2991 ( .A(n2365), .B(n1984), .Z(n1985) );
  NAND U2992 ( .A(n1983), .B(n1985), .Z(n2421) );
  XNOR U2993 ( .A(n3053), .B(n3051), .Z(n1986) );
  NANDN U2994 ( .A(n3056), .B(n1986), .Z(n1987) );
  NAND U2995 ( .A(n3056), .B(n3052), .Z(n1988) );
  NANDN U2996 ( .A(n3055), .B(n1988), .Z(n1989) );
  NAND U2997 ( .A(n1987), .B(n1989), .Z(n3111) );
  XNOR U2998 ( .A(n2478), .B(n2476), .Z(n1990) );
  NANDN U2999 ( .A(n2481), .B(n1990), .Z(n1991) );
  NAND U3000 ( .A(n2481), .B(n2477), .Z(n1992) );
  NANDN U3001 ( .A(n2480), .B(n1992), .Z(n1993) );
  NAND U3002 ( .A(n1991), .B(n1993), .Z(n2536) );
  XNOR U3003 ( .A(n2708), .B(n2706), .Z(n1994) );
  NANDN U3004 ( .A(n2711), .B(n1994), .Z(n1995) );
  NAND U3005 ( .A(n2711), .B(n2707), .Z(n1996) );
  NANDN U3006 ( .A(n2710), .B(n1996), .Z(n1997) );
  NAND U3007 ( .A(n1995), .B(n1997), .Z(n2766) );
  XNOR U3008 ( .A(n3842), .B(n3840), .Z(n1998) );
  NANDN U3009 ( .A(n3845), .B(n1998), .Z(n1999) );
  NAND U3010 ( .A(n3845), .B(n3841), .Z(n2000) );
  NANDN U3011 ( .A(n3844), .B(n2000), .Z(n2001) );
  NAND U3012 ( .A(n1999), .B(n2001), .Z(n3900) );
  AND U3013 ( .A(n2297), .B(n2296), .Z(n2002) );
  XNOR U3014 ( .A(n2295), .B(n2002), .Z(n2309) );
  XOR U3015 ( .A(n3911), .B(n3519), .Z(n3521) );
  XNOR U3016 ( .A(n3398), .B(n3396), .Z(n2003) );
  NANDN U3017 ( .A(n3401), .B(n2003), .Z(n2004) );
  NAND U3018 ( .A(n3401), .B(n3397), .Z(n2005) );
  NANDN U3019 ( .A(n3400), .B(n2005), .Z(n2006) );
  NAND U3020 ( .A(n2004), .B(n2006), .Z(n3456) );
  AND U3021 ( .A(n3543), .B(n3528), .Z(n2007) );
  NAND U3022 ( .A(n3514), .B(n2007), .Z(n2008) );
  NANDN U3023 ( .A(n3528), .B(n3543), .Z(n2009) );
  XNOR U3024 ( .A(x[96]), .B(n2009), .Z(n2010) );
  NANDN U3025 ( .A(n3514), .B(n2010), .Z(n2011) );
  NAND U3026 ( .A(n2008), .B(n2011), .Z(n2012) );
  XNOR U3027 ( .A(n3469), .B(n3472), .Z(n2013) );
  XNOR U3028 ( .A(n2012), .B(n2013), .Z(n3497) );
  XNOR U3029 ( .A(n2823), .B(n2821), .Z(n2014) );
  NANDN U3030 ( .A(n2826), .B(n2014), .Z(n2015) );
  NAND U3031 ( .A(n2826), .B(n2822), .Z(n2016) );
  NANDN U3032 ( .A(n2825), .B(n2016), .Z(n2017) );
  NAND U3033 ( .A(n2015), .B(n2017), .Z(n2881) );
  NANDN U3034 ( .A(n3170), .B(n3171), .Z(n2018) );
  AND U3035 ( .A(n3170), .B(n3168), .Z(n2019) );
  XNOR U3036 ( .A(n2019), .B(n3169), .Z(n2020) );
  NANDN U3037 ( .A(n3171), .B(n2020), .Z(n2021) );
  NAND U3038 ( .A(n2018), .B(n2021), .Z(n3185) );
  XNOR U3039 ( .A(n3727), .B(n3725), .Z(n2022) );
  NANDN U3040 ( .A(n3730), .B(n2022), .Z(n2023) );
  NAND U3041 ( .A(n3730), .B(n3726), .Z(n2024) );
  NANDN U3042 ( .A(n3729), .B(n2024), .Z(n2025) );
  NAND U3043 ( .A(n2023), .B(n2025), .Z(n3785) );
  XNOR U3044 ( .A(n2593), .B(n2591), .Z(n2026) );
  NANDN U3045 ( .A(n2596), .B(n2026), .Z(n2027) );
  NAND U3046 ( .A(n2596), .B(n2592), .Z(n2028) );
  NANDN U3047 ( .A(n2595), .B(n2028), .Z(n2029) );
  NAND U3048 ( .A(n2027), .B(n2029), .Z(n2651) );
  XOR U3049 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3050 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3051 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3052 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3053 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3054 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3055 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3056 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3057 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3058 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3059 ( .A(n2752), .B(n2766), .Z(n2729) );
  ANDN U3060 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3061 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3062 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3063 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3064 ( .A(n3771), .B(n3785), .Z(n3748) );
  NANDN U3065 ( .A(n2137), .B(n2138), .Z(n2032) );
  AND U3066 ( .A(n2137), .B(n2135), .Z(n2033) );
  XNOR U3067 ( .A(n2033), .B(n2136), .Z(n2034) );
  NANDN U3068 ( .A(n2138), .B(n2034), .Z(n2035) );
  NAND U3069 ( .A(n2032), .B(n2035), .Z(n2152) );
  XOR U3070 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3071 ( .A(n3544), .B(n3555), .Z(n3542) );
  NANDN U3072 ( .A(n2940), .B(n2941), .Z(n2036) );
  AND U3073 ( .A(n2940), .B(n2938), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n2939), .Z(n2038) );
  NANDN U3075 ( .A(n2941), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n2955) );
  NANDN U3077 ( .A(n3285), .B(n3286), .Z(n2040) );
  AND U3078 ( .A(n3285), .B(n3283), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n3284), .Z(n2042) );
  NANDN U3080 ( .A(n3286), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n3300) );
  XNOR U3082 ( .A(n3168), .B(n3166), .Z(n2044) );
  NANDN U3083 ( .A(n3171), .B(n2044), .Z(n2045) );
  NAND U3084 ( .A(n3171), .B(n3167), .Z(n2046) );
  NANDN U3085 ( .A(n3170), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2045), .B(n2047), .Z(n3226) );
  NANDN U3087 ( .A(n3844), .B(n3845), .Z(n2048) );
  AND U3088 ( .A(n3844), .B(n3842), .Z(n2049) );
  XNOR U3089 ( .A(n2049), .B(n3843), .Z(n2050) );
  NANDN U3090 ( .A(n3845), .B(n2050), .Z(n2051) );
  NAND U3091 ( .A(n2048), .B(n2051), .Z(n3859) );
  NANDN U3092 ( .A(n3614), .B(n3615), .Z(n2052) );
  AND U3093 ( .A(n3614), .B(n3612), .Z(n2053) );
  XNOR U3094 ( .A(n2053), .B(n3613), .Z(n2054) );
  NANDN U3095 ( .A(n3615), .B(n2054), .Z(n2055) );
  NAND U3096 ( .A(n2052), .B(n2055), .Z(n3629) );
  NANDN U3097 ( .A(n3055), .B(n3056), .Z(n2056) );
  AND U3098 ( .A(n3055), .B(n3053), .Z(n2057) );
  XNOR U3099 ( .A(n2057), .B(n3054), .Z(n2058) );
  NANDN U3100 ( .A(n3056), .B(n2058), .Z(n2059) );
  NAND U3101 ( .A(n2056), .B(n2059), .Z(n3070) );
  NANDN U3102 ( .A(n2365), .B(n2366), .Z(n2060) );
  AND U3103 ( .A(n2365), .B(n2363), .Z(n2061) );
  XNOR U3104 ( .A(n2061), .B(n2364), .Z(n2062) );
  NANDN U3105 ( .A(n2366), .B(n2062), .Z(n2063) );
  NAND U3106 ( .A(n2060), .B(n2063), .Z(n2380) );
  NANDN U3107 ( .A(n2480), .B(n2481), .Z(n2064) );
  AND U3108 ( .A(n2480), .B(n2478), .Z(n2065) );
  XNOR U3109 ( .A(n2065), .B(n2479), .Z(n2066) );
  NANDN U3110 ( .A(n2481), .B(n2066), .Z(n2067) );
  NAND U3111 ( .A(n2064), .B(n2067), .Z(n2495) );
  NANDN U3112 ( .A(n2595), .B(n2596), .Z(n2068) );
  AND U3113 ( .A(n2595), .B(n2593), .Z(n2069) );
  XNOR U3114 ( .A(n2069), .B(n2594), .Z(n2070) );
  NANDN U3115 ( .A(n2596), .B(n2070), .Z(n2071) );
  NAND U3116 ( .A(n2068), .B(n2071), .Z(n2610) );
  NANDN U3117 ( .A(n2710), .B(n2711), .Z(n2072) );
  AND U3118 ( .A(n2710), .B(n2708), .Z(n2073) );
  XNOR U3119 ( .A(n2073), .B(n2709), .Z(n2074) );
  NANDN U3120 ( .A(n2711), .B(n2074), .Z(n2075) );
  NAND U3121 ( .A(n2072), .B(n2075), .Z(n2725) );
  XOR U3122 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3123 ( .A(n3400), .B(n3401), .Z(n2076) );
  AND U3124 ( .A(n3400), .B(n3398), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3399), .Z(n2078) );
  NANDN U3126 ( .A(n3401), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3415) );
  NANDN U3128 ( .A(n2825), .B(n2826), .Z(n2080) );
  AND U3129 ( .A(n2825), .B(n2823), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2824), .Z(n2082) );
  NANDN U3131 ( .A(n2826), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2840) );
  NANDN U3133 ( .A(n3729), .B(n3730), .Z(n2084) );
  AND U3134 ( .A(n3729), .B(n3727), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3728), .Z(n2086) );
  NANDN U3136 ( .A(n3730), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3744) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_8 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U2967 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U2968 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U2969 ( .A(n3911), .B(n3519), .Z(n3521) );
  XNOR U2970 ( .A(n3283), .B(n3281), .Z(n1966) );
  NANDN U2971 ( .A(n3286), .B(n1966), .Z(n1967) );
  NAND U2972 ( .A(n3286), .B(n3282), .Z(n1968) );
  NANDN U2973 ( .A(n3285), .B(n1968), .Z(n1969) );
  NAND U2974 ( .A(n1967), .B(n1969), .Z(n3341) );
  XNOR U2975 ( .A(n2135), .B(n2133), .Z(n1970) );
  NANDN U2976 ( .A(n2138), .B(n1970), .Z(n1971) );
  NAND U2977 ( .A(n2138), .B(n2134), .Z(n1972) );
  NANDN U2978 ( .A(n2137), .B(n1972), .Z(n1973) );
  NAND U2979 ( .A(n1971), .B(n1973), .Z(n2193) );
  AND U2980 ( .A(n2297), .B(n2296), .Z(n1974) );
  XNOR U2981 ( .A(n2295), .B(n1974), .Z(n2309) );
  XNOR U2982 ( .A(n2363), .B(n2361), .Z(n1975) );
  NANDN U2983 ( .A(n2366), .B(n1975), .Z(n1976) );
  NAND U2984 ( .A(n2366), .B(n2362), .Z(n1977) );
  NANDN U2985 ( .A(n2365), .B(n1977), .Z(n1978) );
  NAND U2986 ( .A(n1976), .B(n1978), .Z(n2421) );
  XNOR U2987 ( .A(n3053), .B(n3051), .Z(n1979) );
  NANDN U2988 ( .A(n3056), .B(n1979), .Z(n1980) );
  NAND U2989 ( .A(n3056), .B(n3052), .Z(n1981) );
  NANDN U2990 ( .A(n3055), .B(n1981), .Z(n1982) );
  NAND U2991 ( .A(n1980), .B(n1982), .Z(n3111) );
  XNOR U2992 ( .A(n3398), .B(n3396), .Z(n1983) );
  NANDN U2993 ( .A(n3401), .B(n1983), .Z(n1984) );
  NAND U2994 ( .A(n3401), .B(n3397), .Z(n1985) );
  NANDN U2995 ( .A(n3400), .B(n1985), .Z(n1986) );
  NAND U2996 ( .A(n1984), .B(n1986), .Z(n3456) );
  AND U2997 ( .A(n3543), .B(n3528), .Z(n1987) );
  NAND U2998 ( .A(n3514), .B(n1987), .Z(n1988) );
  NANDN U2999 ( .A(n3528), .B(n3543), .Z(n1989) );
  XNOR U3000 ( .A(x[96]), .B(n1989), .Z(n1990) );
  NANDN U3001 ( .A(n3514), .B(n1990), .Z(n1991) );
  NAND U3002 ( .A(n1988), .B(n1991), .Z(n1992) );
  XNOR U3003 ( .A(n3469), .B(n3472), .Z(n1993) );
  XNOR U3004 ( .A(n1992), .B(n1993), .Z(n3497) );
  XNOR U3005 ( .A(n2823), .B(n2821), .Z(n1994) );
  NANDN U3006 ( .A(n2826), .B(n1994), .Z(n1995) );
  NAND U3007 ( .A(n2826), .B(n2822), .Z(n1996) );
  NANDN U3008 ( .A(n2825), .B(n1996), .Z(n1997) );
  NAND U3009 ( .A(n1995), .B(n1997), .Z(n2881) );
  XNOR U3010 ( .A(n2478), .B(n2476), .Z(n1998) );
  NANDN U3011 ( .A(n2481), .B(n1998), .Z(n1999) );
  NAND U3012 ( .A(n2481), .B(n2477), .Z(n2000) );
  NANDN U3013 ( .A(n2480), .B(n2000), .Z(n2001) );
  NAND U3014 ( .A(n1999), .B(n2001), .Z(n2536) );
  XNOR U3015 ( .A(n2938), .B(n2936), .Z(n2002) );
  NANDN U3016 ( .A(n2941), .B(n2002), .Z(n2003) );
  NAND U3017 ( .A(n2941), .B(n2937), .Z(n2004) );
  NANDN U3018 ( .A(n2940), .B(n2004), .Z(n2005) );
  NAND U3019 ( .A(n2003), .B(n2005), .Z(n2996) );
  XNOR U3020 ( .A(n3612), .B(n3610), .Z(n2006) );
  NANDN U3021 ( .A(n3615), .B(n2006), .Z(n2007) );
  NAND U3022 ( .A(n3615), .B(n3611), .Z(n2008) );
  NANDN U3023 ( .A(n3614), .B(n2008), .Z(n2009) );
  NAND U3024 ( .A(n2007), .B(n2009), .Z(n3670) );
  XNOR U3025 ( .A(n2708), .B(n2706), .Z(n2010) );
  NANDN U3026 ( .A(n2711), .B(n2010), .Z(n2011) );
  NAND U3027 ( .A(n2711), .B(n2707), .Z(n2012) );
  NANDN U3028 ( .A(n2710), .B(n2012), .Z(n2013) );
  NAND U3029 ( .A(n2011), .B(n2013), .Z(n2766) );
  XNOR U3030 ( .A(n3842), .B(n3840), .Z(n2014) );
  NANDN U3031 ( .A(n3845), .B(n2014), .Z(n2015) );
  NAND U3032 ( .A(n3845), .B(n3841), .Z(n2016) );
  NANDN U3033 ( .A(n3844), .B(n2016), .Z(n2017) );
  NAND U3034 ( .A(n2015), .B(n2017), .Z(n3900) );
  NANDN U3035 ( .A(n3170), .B(n3171), .Z(n2018) );
  AND U3036 ( .A(n3170), .B(n3168), .Z(n2019) );
  XNOR U3037 ( .A(n2019), .B(n3169), .Z(n2020) );
  NANDN U3038 ( .A(n3171), .B(n2020), .Z(n2021) );
  NAND U3039 ( .A(n2018), .B(n2021), .Z(n3185) );
  NANDN U3040 ( .A(n2595), .B(n2596), .Z(n2022) );
  AND U3041 ( .A(n2595), .B(n2593), .Z(n2023) );
  XNOR U3042 ( .A(n2023), .B(n2594), .Z(n2024) );
  NANDN U3043 ( .A(n2596), .B(n2024), .Z(n2025) );
  NAND U3044 ( .A(n2022), .B(n2025), .Z(n2610) );
  XNOR U3045 ( .A(n3727), .B(n3725), .Z(n2026) );
  NANDN U3046 ( .A(n3730), .B(n2026), .Z(n2027) );
  NAND U3047 ( .A(n3730), .B(n3726), .Z(n2028) );
  NANDN U3048 ( .A(n3729), .B(n2028), .Z(n2029) );
  NAND U3049 ( .A(n2027), .B(n2029), .Z(n3785) );
  XOR U3050 ( .A(n3097), .B(n3111), .Z(n3074) );
  ANDN U3051 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3052 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3053 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3054 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3055 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3056 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3057 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3058 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3059 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3060 ( .A(n3886), .B(n3900), .Z(n3863) );
  XOR U3061 ( .A(n2522), .B(n2536), .Z(n2499) );
  XOR U3062 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3063 ( .A(n2752), .B(n2766), .Z(n2729) );
  XOR U3064 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U3065 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3066 ( .A(n3771), .B(n3785), .Z(n3748) );
  NANDN U3067 ( .A(n2825), .B(n2826), .Z(n2032) );
  AND U3068 ( .A(n2825), .B(n2823), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n2824), .Z(n2034) );
  NANDN U3070 ( .A(n2826), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n2840) );
  NANDN U3072 ( .A(n2137), .B(n2138), .Z(n2036) );
  AND U3073 ( .A(n2137), .B(n2135), .Z(n2037) );
  XNOR U3074 ( .A(n2037), .B(n2136), .Z(n2038) );
  NANDN U3075 ( .A(n2138), .B(n2038), .Z(n2039) );
  NAND U3076 ( .A(n2036), .B(n2039), .Z(n2152) );
  NANDN U3077 ( .A(n3285), .B(n3286), .Z(n2040) );
  AND U3078 ( .A(n3285), .B(n3283), .Z(n2041) );
  XNOR U3079 ( .A(n2041), .B(n3284), .Z(n2042) );
  NANDN U3080 ( .A(n3286), .B(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2040), .B(n2043), .Z(n3300) );
  NANDN U3082 ( .A(n3400), .B(n3401), .Z(n2044) );
  AND U3083 ( .A(n3400), .B(n3398), .Z(n2045) );
  XNOR U3084 ( .A(n2045), .B(n3399), .Z(n2046) );
  NANDN U3085 ( .A(n3401), .B(n2046), .Z(n2047) );
  NAND U3086 ( .A(n2044), .B(n2047), .Z(n3415) );
  XOR U3087 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3088 ( .A(n2940), .B(n2941), .Z(n2048) );
  AND U3089 ( .A(n2940), .B(n2938), .Z(n2049) );
  XNOR U3090 ( .A(n2049), .B(n2939), .Z(n2050) );
  NANDN U3091 ( .A(n2941), .B(n2050), .Z(n2051) );
  NAND U3092 ( .A(n2048), .B(n2051), .Z(n2955) );
  NANDN U3093 ( .A(n3055), .B(n3056), .Z(n2052) );
  AND U3094 ( .A(n3055), .B(n3053), .Z(n2053) );
  XNOR U3095 ( .A(n2053), .B(n3054), .Z(n2054) );
  NANDN U3096 ( .A(n3056), .B(n2054), .Z(n2055) );
  NAND U3097 ( .A(n2052), .B(n2055), .Z(n3070) );
  NANDN U3098 ( .A(n2365), .B(n2366), .Z(n2056) );
  AND U3099 ( .A(n2365), .B(n2363), .Z(n2057) );
  XNOR U3100 ( .A(n2057), .B(n2364), .Z(n2058) );
  NANDN U3101 ( .A(n2366), .B(n2058), .Z(n2059) );
  NAND U3102 ( .A(n2056), .B(n2059), .Z(n2380) );
  NANDN U3103 ( .A(n3844), .B(n3845), .Z(n2060) );
  AND U3104 ( .A(n3844), .B(n3842), .Z(n2061) );
  XNOR U3105 ( .A(n2061), .B(n3843), .Z(n2062) );
  NANDN U3106 ( .A(n3845), .B(n2062), .Z(n2063) );
  NAND U3107 ( .A(n2060), .B(n2063), .Z(n3859) );
  XNOR U3108 ( .A(n3168), .B(n3166), .Z(n2064) );
  NANDN U3109 ( .A(n3171), .B(n2064), .Z(n2065) );
  NAND U3110 ( .A(n3171), .B(n3167), .Z(n2066) );
  NANDN U3111 ( .A(n3170), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2065), .B(n2067), .Z(n3226) );
  NANDN U3113 ( .A(n2480), .B(n2481), .Z(n2068) );
  AND U3114 ( .A(n2480), .B(n2478), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n2479), .Z(n2070) );
  NANDN U3116 ( .A(n2481), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n2495) );
  XNOR U3118 ( .A(n2593), .B(n2591), .Z(n2072) );
  NANDN U3119 ( .A(n2596), .B(n2072), .Z(n2073) );
  NAND U3120 ( .A(n2596), .B(n2592), .Z(n2074) );
  NANDN U3121 ( .A(n2595), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2073), .B(n2075), .Z(n2651) );
  NANDN U3123 ( .A(n3614), .B(n3615), .Z(n2076) );
  AND U3124 ( .A(n3614), .B(n3612), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3613), .Z(n2078) );
  NANDN U3126 ( .A(n3615), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3629) );
  NANDN U3128 ( .A(n2710), .B(n2711), .Z(n2080) );
  AND U3129 ( .A(n2710), .B(n2708), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2709), .Z(n2082) );
  NANDN U3131 ( .A(n2711), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2725) );
  NANDN U3133 ( .A(n3729), .B(n3730), .Z(n2084) );
  AND U3134 ( .A(n3729), .B(n3727), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n3728), .Z(n2086) );
  NANDN U3136 ( .A(n3730), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n3744) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module SubBytes_9 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965;

  AND U2962 ( .A(n2250), .B(n2258), .Z(n1963) );
  XNOR U2963 ( .A(n2306), .B(n2266), .Z(n1964) );
  XNOR U2964 ( .A(n1963), .B(n1964), .Z(n1965) );
  XOR U2965 ( .A(n2209), .B(n1965), .Z(n2225) );
  XOR U2966 ( .A(n3912), .B(n3520), .Z(n3530) );
  XOR U2967 ( .A(n3911), .B(n3519), .Z(n3521) );
  AND U2968 ( .A(n3543), .B(n3528), .Z(n1966) );
  NAND U2969 ( .A(n3514), .B(n1966), .Z(n1967) );
  NANDN U2970 ( .A(n3528), .B(n3543), .Z(n1968) );
  XNOR U2971 ( .A(x[96]), .B(n1968), .Z(n1969) );
  NANDN U2972 ( .A(n3514), .B(n1969), .Z(n1970) );
  NAND U2973 ( .A(n1967), .B(n1970), .Z(n1971) );
  XNOR U2974 ( .A(n3469), .B(n3472), .Z(n1972) );
  XNOR U2975 ( .A(n1971), .B(n1972), .Z(n3497) );
  XNOR U2976 ( .A(n3398), .B(n3396), .Z(n1973) );
  NANDN U2977 ( .A(n3401), .B(n1973), .Z(n1974) );
  NAND U2978 ( .A(n3401), .B(n3397), .Z(n1975) );
  NANDN U2979 ( .A(n3400), .B(n1975), .Z(n1976) );
  NAND U2980 ( .A(n1974), .B(n1976), .Z(n3456) );
  AND U2981 ( .A(n2297), .B(n2296), .Z(n1977) );
  XNOR U2982 ( .A(n2295), .B(n1977), .Z(n2309) );
  XNOR U2983 ( .A(n2823), .B(n2821), .Z(n1978) );
  NANDN U2984 ( .A(n2826), .B(n1978), .Z(n1979) );
  NAND U2985 ( .A(n2826), .B(n2822), .Z(n1980) );
  NANDN U2986 ( .A(n2825), .B(n1980), .Z(n1981) );
  NAND U2987 ( .A(n1979), .B(n1981), .Z(n2881) );
  XNOR U2988 ( .A(n2938), .B(n2936), .Z(n1982) );
  NANDN U2989 ( .A(n2941), .B(n1982), .Z(n1983) );
  NAND U2990 ( .A(n2941), .B(n2937), .Z(n1984) );
  NANDN U2991 ( .A(n2940), .B(n1984), .Z(n1985) );
  NAND U2992 ( .A(n1983), .B(n1985), .Z(n2996) );
  XNOR U2993 ( .A(n2478), .B(n2476), .Z(n1986) );
  NANDN U2994 ( .A(n2481), .B(n1986), .Z(n1987) );
  NAND U2995 ( .A(n2481), .B(n2477), .Z(n1988) );
  NANDN U2996 ( .A(n2480), .B(n1988), .Z(n1989) );
  NAND U2997 ( .A(n1987), .B(n1989), .Z(n2536) );
  XOR U2998 ( .A(n3886), .B(n3900), .Z(n3863) );
  XNOR U2999 ( .A(n3283), .B(n3281), .Z(n1990) );
  NANDN U3000 ( .A(n3286), .B(n1990), .Z(n1991) );
  NAND U3001 ( .A(n3286), .B(n3282), .Z(n1992) );
  NANDN U3002 ( .A(n3285), .B(n1992), .Z(n1993) );
  NAND U3003 ( .A(n1991), .B(n1993), .Z(n3341) );
  XNOR U3004 ( .A(n2135), .B(n2133), .Z(n1994) );
  NANDN U3005 ( .A(n2138), .B(n1994), .Z(n1995) );
  NAND U3006 ( .A(n2138), .B(n2134), .Z(n1996) );
  NANDN U3007 ( .A(n2137), .B(n1996), .Z(n1997) );
  NAND U3008 ( .A(n1995), .B(n1997), .Z(n2193) );
  XNOR U3009 ( .A(n2593), .B(n2591), .Z(n1998) );
  NANDN U3010 ( .A(n2596), .B(n1998), .Z(n1999) );
  NAND U3011 ( .A(n2596), .B(n2592), .Z(n2000) );
  NANDN U3012 ( .A(n2595), .B(n2000), .Z(n2001) );
  NAND U3013 ( .A(n1999), .B(n2001), .Z(n2651) );
  XNOR U3014 ( .A(n3168), .B(n3166), .Z(n2002) );
  NANDN U3015 ( .A(n3171), .B(n2002), .Z(n2003) );
  NAND U3016 ( .A(n3171), .B(n3167), .Z(n2004) );
  NANDN U3017 ( .A(n3170), .B(n2004), .Z(n2005) );
  NAND U3018 ( .A(n2003), .B(n2005), .Z(n3226) );
  XNOR U3019 ( .A(n3727), .B(n3725), .Z(n2006) );
  NANDN U3020 ( .A(n3730), .B(n2006), .Z(n2007) );
  NAND U3021 ( .A(n3730), .B(n3726), .Z(n2008) );
  NANDN U3022 ( .A(n3729), .B(n2008), .Z(n2009) );
  NAND U3023 ( .A(n2007), .B(n2009), .Z(n3785) );
  XNOR U3024 ( .A(n3612), .B(n3610), .Z(n2010) );
  NANDN U3025 ( .A(n3615), .B(n2010), .Z(n2011) );
  NAND U3026 ( .A(n3615), .B(n3611), .Z(n2012) );
  NANDN U3027 ( .A(n3614), .B(n2012), .Z(n2013) );
  NAND U3028 ( .A(n2011), .B(n2013), .Z(n3670) );
  XNOR U3029 ( .A(n2363), .B(n2361), .Z(n2014) );
  NANDN U3030 ( .A(n2366), .B(n2014), .Z(n2015) );
  NAND U3031 ( .A(n2366), .B(n2362), .Z(n2016) );
  NANDN U3032 ( .A(n2365), .B(n2016), .Z(n2017) );
  NAND U3033 ( .A(n2015), .B(n2017), .Z(n2421) );
  XNOR U3034 ( .A(n3053), .B(n3051), .Z(n2018) );
  NANDN U3035 ( .A(n3056), .B(n2018), .Z(n2019) );
  NAND U3036 ( .A(n3056), .B(n3052), .Z(n2020) );
  NANDN U3037 ( .A(n3055), .B(n2020), .Z(n2021) );
  NAND U3038 ( .A(n2019), .B(n2021), .Z(n3111) );
  XNOR U3039 ( .A(n2708), .B(n2706), .Z(n2022) );
  NANDN U3040 ( .A(n2711), .B(n2022), .Z(n2023) );
  NAND U3041 ( .A(n2711), .B(n2707), .Z(n2024) );
  NANDN U3042 ( .A(n2710), .B(n2024), .Z(n2025) );
  NAND U3043 ( .A(n2023), .B(n2025), .Z(n2766) );
  NANDN U3044 ( .A(n3844), .B(n3845), .Z(n2026) );
  AND U3045 ( .A(n3844), .B(n3842), .Z(n2027) );
  XNOR U3046 ( .A(n2027), .B(n3843), .Z(n2028) );
  NANDN U3047 ( .A(n3845), .B(n2028), .Z(n2029) );
  NAND U3048 ( .A(n2026), .B(n2029), .Z(n3859) );
  XOR U3049 ( .A(n3656), .B(n3670), .Z(n3633) );
  XOR U3050 ( .A(n2522), .B(n2536), .Z(n2499) );
  ANDN U3051 ( .B(n2211), .A(x[9]), .Z(n2030) );
  XNOR U3052 ( .A(n2210), .B(n2225), .Z(n2031) );
  XNOR U3053 ( .A(n2030), .B(n2031), .Z(n2228) );
  XOR U3054 ( .A(n3097), .B(n3111), .Z(n3074) );
  XOR U3055 ( .A(n3442), .B(n3456), .Z(n3419) );
  XOR U3056 ( .A(n3212), .B(n3226), .Z(n3189) );
  XOR U3057 ( .A(n2867), .B(n2881), .Z(n2844) );
  XOR U3058 ( .A(n2982), .B(n2996), .Z(n2959) );
  XOR U3059 ( .A(n2637), .B(n2651), .Z(n2614) );
  XOR U3060 ( .A(n2179), .B(n2193), .Z(n2156) );
  XOR U3061 ( .A(n3327), .B(n3341), .Z(n3304) );
  XOR U3062 ( .A(n3771), .B(n3785), .Z(n3748) );
  XOR U3063 ( .A(n2407), .B(n2421), .Z(n2384) );
  XOR U3064 ( .A(n3470), .B(n3471), .Z(n3546) );
  XOR U3065 ( .A(n3544), .B(n3555), .Z(n3542) );
  XOR U3066 ( .A(n2752), .B(n2766), .Z(n2729) );
  NANDN U3067 ( .A(n3400), .B(n3401), .Z(n2032) );
  AND U3068 ( .A(n3400), .B(n3398), .Z(n2033) );
  XNOR U3069 ( .A(n2033), .B(n3399), .Z(n2034) );
  NANDN U3070 ( .A(n3401), .B(n2034), .Z(n2035) );
  NAND U3071 ( .A(n2032), .B(n2035), .Z(n3415) );
  XOR U3072 ( .A(n2283), .B(n2293), .Z(n3960) );
  NANDN U3073 ( .A(n3170), .B(n3171), .Z(n2036) );
  AND U3074 ( .A(n3170), .B(n3168), .Z(n2037) );
  XNOR U3075 ( .A(n2037), .B(n3169), .Z(n2038) );
  NANDN U3076 ( .A(n3171), .B(n2038), .Z(n2039) );
  NAND U3077 ( .A(n2036), .B(n2039), .Z(n3185) );
  NANDN U3078 ( .A(n2825), .B(n2826), .Z(n2040) );
  AND U3079 ( .A(n2825), .B(n2823), .Z(n2041) );
  XNOR U3080 ( .A(n2041), .B(n2824), .Z(n2042) );
  NANDN U3081 ( .A(n2826), .B(n2042), .Z(n2043) );
  NAND U3082 ( .A(n2040), .B(n2043), .Z(n2840) );
  NANDN U3083 ( .A(n2940), .B(n2941), .Z(n2044) );
  AND U3084 ( .A(n2940), .B(n2938), .Z(n2045) );
  XNOR U3085 ( .A(n2045), .B(n2939), .Z(n2046) );
  NANDN U3086 ( .A(n2941), .B(n2046), .Z(n2047) );
  NAND U3087 ( .A(n2044), .B(n2047), .Z(n2955) );
  NANDN U3088 ( .A(n2480), .B(n2481), .Z(n2048) );
  AND U3089 ( .A(n2480), .B(n2478), .Z(n2049) );
  XNOR U3090 ( .A(n2049), .B(n2479), .Z(n2050) );
  NANDN U3091 ( .A(n2481), .B(n2050), .Z(n2051) );
  NAND U3092 ( .A(n2048), .B(n2051), .Z(n2495) );
  NANDN U3093 ( .A(n2595), .B(n2596), .Z(n2052) );
  AND U3094 ( .A(n2595), .B(n2593), .Z(n2053) );
  XNOR U3095 ( .A(n2053), .B(n2594), .Z(n2054) );
  NANDN U3096 ( .A(n2596), .B(n2054), .Z(n2055) );
  NAND U3097 ( .A(n2052), .B(n2055), .Z(n2610) );
  XNOR U3098 ( .A(n3842), .B(n3840), .Z(n2056) );
  NANDN U3099 ( .A(n3845), .B(n2056), .Z(n2057) );
  NAND U3100 ( .A(n3845), .B(n3841), .Z(n2058) );
  NANDN U3101 ( .A(n3844), .B(n2058), .Z(n2059) );
  NAND U3102 ( .A(n2057), .B(n2059), .Z(n3900) );
  NANDN U3103 ( .A(n2137), .B(n2138), .Z(n2060) );
  AND U3104 ( .A(n2137), .B(n2135), .Z(n2061) );
  XNOR U3105 ( .A(n2061), .B(n2136), .Z(n2062) );
  NANDN U3106 ( .A(n2138), .B(n2062), .Z(n2063) );
  NAND U3107 ( .A(n2060), .B(n2063), .Z(n2152) );
  NANDN U3108 ( .A(n3285), .B(n3286), .Z(n2064) );
  AND U3109 ( .A(n3285), .B(n3283), .Z(n2065) );
  XNOR U3110 ( .A(n2065), .B(n3284), .Z(n2066) );
  NANDN U3111 ( .A(n3286), .B(n2066), .Z(n2067) );
  NAND U3112 ( .A(n2064), .B(n2067), .Z(n3300) );
  NANDN U3113 ( .A(n3729), .B(n3730), .Z(n2068) );
  AND U3114 ( .A(n3729), .B(n3727), .Z(n2069) );
  XNOR U3115 ( .A(n2069), .B(n3728), .Z(n2070) );
  NANDN U3116 ( .A(n3730), .B(n2070), .Z(n2071) );
  NAND U3117 ( .A(n2068), .B(n2071), .Z(n3744) );
  NANDN U3118 ( .A(n3055), .B(n3056), .Z(n2072) );
  AND U3119 ( .A(n3055), .B(n3053), .Z(n2073) );
  XNOR U3120 ( .A(n2073), .B(n3054), .Z(n2074) );
  NANDN U3121 ( .A(n3056), .B(n2074), .Z(n2075) );
  NAND U3122 ( .A(n2072), .B(n2075), .Z(n3070) );
  NANDN U3123 ( .A(n3614), .B(n3615), .Z(n2076) );
  AND U3124 ( .A(n3614), .B(n3612), .Z(n2077) );
  XNOR U3125 ( .A(n2077), .B(n3613), .Z(n2078) );
  NANDN U3126 ( .A(n3615), .B(n2078), .Z(n2079) );
  NAND U3127 ( .A(n2076), .B(n2079), .Z(n3629) );
  NANDN U3128 ( .A(n2365), .B(n2366), .Z(n2080) );
  AND U3129 ( .A(n2365), .B(n2363), .Z(n2081) );
  XNOR U3130 ( .A(n2081), .B(n2364), .Z(n2082) );
  NANDN U3131 ( .A(n2366), .B(n2082), .Z(n2083) );
  NAND U3132 ( .A(n2080), .B(n2083), .Z(n2380) );
  NANDN U3133 ( .A(n2710), .B(n2711), .Z(n2084) );
  AND U3134 ( .A(n2710), .B(n2708), .Z(n2085) );
  XNOR U3135 ( .A(n2085), .B(n2709), .Z(n2086) );
  NANDN U3136 ( .A(n2711), .B(n2086), .Z(n2087) );
  NAND U3137 ( .A(n2084), .B(n2087), .Z(n2725) );
  XOR U3138 ( .A(x[1]), .B(x[3]), .Z(n2091) );
  XOR U3139 ( .A(x[0]), .B(x[6]), .Z(n2089) );
  XNOR U3140 ( .A(n2091), .B(n2089), .Z(n2088) );
  XNOR U3141 ( .A(x[2]), .B(n2088), .Z(n2159) );
  IV U3142 ( .A(n2159), .Z(n2093) );
  XNOR U3143 ( .A(x[0]), .B(n2093), .Z(n2141) );
  XNOR U3144 ( .A(x[4]), .B(x[7]), .Z(n2090) );
  IV U3145 ( .A(n2090), .Z(n2154) );
  AND U3146 ( .A(n2141), .B(n2154), .Z(n2098) );
  XOR U3147 ( .A(x[7]), .B(x[2]), .Z(n2181) );
  XNOR U3148 ( .A(n2089), .B(x[5]), .Z(n2104) );
  IV U3149 ( .A(n2104), .Z(n2150) );
  XOR U3150 ( .A(n2091), .B(n2090), .Z(n2115) );
  IV U3151 ( .A(n2115), .Z(n2130) );
  XNOR U3152 ( .A(n2130), .B(x[0]), .Z(n2131) );
  XNOR U3153 ( .A(n2150), .B(n2131), .Z(n2143) );
  NAND U3154 ( .A(n2181), .B(n2143), .Z(n2092) );
  XNOR U3155 ( .A(n2098), .B(n2092), .Z(n2111) );
  XOR U3156 ( .A(x[1]), .B(x[7]), .Z(n2149) );
  XOR U3157 ( .A(n2093), .B(n2150), .Z(n2139) );
  ANDN U3158 ( .B(n2149), .A(n2139), .Z(n2100) );
  XOR U3159 ( .A(x[7]), .B(n2150), .Z(n2192) );
  IV U3160 ( .A(n2192), .Z(n2103) );
  NAND U3161 ( .A(n2093), .B(n2103), .Z(n2094) );
  XOR U3162 ( .A(n2100), .B(n2094), .Z(n2095) );
  XNOR U3163 ( .A(n2111), .B(n2095), .Z(n2135) );
  NANDN U3164 ( .A(x[1]), .B(n2104), .Z(n2102) );
  XNOR U3165 ( .A(n2130), .B(n2139), .Z(n2174) );
  XOR U3166 ( .A(x[4]), .B(x[2]), .Z(n2157) );
  AND U3167 ( .A(n2174), .B(n2157), .Z(n2097) );
  XNOR U3168 ( .A(n2159), .B(n2192), .Z(n2096) );
  XNOR U3169 ( .A(n2097), .B(n2096), .Z(n2099) );
  XOR U3170 ( .A(n2099), .B(n2098), .Z(n2119) );
  XNOR U3171 ( .A(n2100), .B(n2119), .Z(n2101) );
  XNOR U3172 ( .A(n2102), .B(n2101), .Z(n2133) );
  IV U3173 ( .A(n2133), .Z(n2136) );
  NAND U3174 ( .A(n2135), .B(n2136), .Z(n2129) );
  NANDN U3175 ( .A(n2135), .B(n2136), .Z(n2123) );
  XNOR U3176 ( .A(x[2]), .B(n2103), .Z(n2110) );
  XNOR U3177 ( .A(x[1]), .B(n2110), .Z(n2114) );
  IV U3178 ( .A(n2114), .Z(n2168) );
  XNOR U3179 ( .A(x[4]), .B(n2104), .Z(n2180) );
  OR U3180 ( .A(x[0]), .B(n2180), .Z(n2105) );
  XNOR U3181 ( .A(n2168), .B(n2105), .Z(n2106) );
  NANDN U3182 ( .A(n2115), .B(n2106), .Z(n2109) );
  ANDN U3183 ( .B(x[0]), .A(n2180), .Z(n2107) );
  NAND U3184 ( .A(n2115), .B(n2107), .Z(n2108) );
  NAND U3185 ( .A(n2109), .B(n2108), .Z(n2113) );
  XNOR U3186 ( .A(n2111), .B(n2110), .Z(n2112) );
  XOR U3187 ( .A(n2113), .B(n2112), .Z(n2137) );
  IV U3188 ( .A(n2135), .Z(n2134) );
  ANDN U3189 ( .B(n2137), .A(n2134), .Z(n2120) );
  AND U3190 ( .A(x[0]), .B(n2114), .Z(n2117) );
  NAND U3191 ( .A(n2115), .B(n2180), .Z(n2116) );
  XNOR U3192 ( .A(n2117), .B(n2116), .Z(n2118) );
  XNOR U3193 ( .A(n2119), .B(n2118), .Z(n2138) );
  XNOR U3194 ( .A(n2120), .B(n2138), .Z(n2121) );
  NAND U3195 ( .A(n2133), .B(n2121), .Z(n2122) );
  NAND U3196 ( .A(n2123), .B(n2122), .Z(n2167) );
  IV U3197 ( .A(n2167), .Z(n2142) );
  OR U3198 ( .A(n2137), .B(n2133), .Z(n2124) );
  NAND U3199 ( .A(n2134), .B(n2124), .Z(n2127) );
  XOR U3200 ( .A(n2137), .B(n2138), .Z(n2125) );
  NANDN U3201 ( .A(n2136), .B(n2125), .Z(n2126) );
  NAND U3202 ( .A(n2127), .B(n2126), .Z(n2179) );
  NANDN U3203 ( .A(n2142), .B(n2179), .Z(n2128) );
  AND U3204 ( .A(n2129), .B(n2128), .Z(n2170) );
  AND U3205 ( .A(n2170), .B(n2130), .Z(n2145) );
  OR U3206 ( .A(n2131), .B(n2142), .Z(n2132) );
  XNOR U3207 ( .A(n2145), .B(n2132), .Z(n2178) );
  XOR U3208 ( .A(n2193), .B(n2152), .Z(n2148) );
  ANDN U3209 ( .B(n2148), .A(n2139), .Z(n2160) );
  NAND U3210 ( .A(n2150), .B(n2152), .Z(n2140) );
  XNOR U3211 ( .A(n2160), .B(n2140), .Z(n2185) );
  XNOR U3212 ( .A(n2178), .B(n2185), .Z(z[2]) );
  AND U3213 ( .A(x[0]), .B(n2179), .Z(n2147) );
  AND U3214 ( .A(n2141), .B(n2156), .Z(n2177) );
  XOR U3215 ( .A(n2142), .B(n2152), .Z(n2155) );
  IV U3216 ( .A(n2155), .Z(n2182) );
  NAND U3217 ( .A(n2182), .B(n2143), .Z(n2144) );
  XNOR U3218 ( .A(n2177), .B(n2144), .Z(n2161) );
  XNOR U3219 ( .A(n2145), .B(n2161), .Z(n2146) );
  XNOR U3220 ( .A(n2147), .B(n2146), .Z(n3955) );
  AND U3221 ( .A(n2149), .B(n2148), .Z(n2194) );
  XOR U3222 ( .A(x[1]), .B(n2150), .Z(n2151) );
  NAND U3223 ( .A(n2152), .B(n2151), .Z(n2153) );
  XNOR U3224 ( .A(n2194), .B(n2153), .Z(n2165) );
  AND U3225 ( .A(n2156), .B(n2154), .Z(n2184) );
  XNOR U3226 ( .A(n2156), .B(n2155), .Z(n2175) );
  NAND U3227 ( .A(n2175), .B(n2157), .Z(n2158) );
  XNOR U3228 ( .A(n2184), .B(n2158), .Z(n2171) );
  AND U3229 ( .A(n2193), .B(n2159), .Z(n2163) );
  XNOR U3230 ( .A(n2161), .B(n2160), .Z(n2162) );
  XNOR U3231 ( .A(n2163), .B(n2162), .Z(n3943) );
  XNOR U3232 ( .A(n2171), .B(n3943), .Z(n2164) );
  XNOR U3233 ( .A(n2165), .B(n2164), .Z(n2166) );
  XNOR U3234 ( .A(n3955), .B(n2166), .Z(z[5]) );
  AND U3235 ( .A(n2168), .B(n2167), .Z(n2173) );
  XOR U3236 ( .A(n2168), .B(n2180), .Z(n2169) );
  AND U3237 ( .A(n2170), .B(n2169), .Z(n2189) );
  XNOR U3238 ( .A(n2171), .B(n2189), .Z(n2172) );
  XNOR U3239 ( .A(n2173), .B(n2172), .Z(n2200) );
  NAND U3240 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U3241 ( .A(n2177), .B(n2176), .Z(n2188) );
  XNOR U3242 ( .A(n2178), .B(n2188), .Z(n3910) );
  XNOR U3243 ( .A(n2200), .B(n3910), .Z(n2198) );
  AND U3244 ( .A(n2180), .B(n2179), .Z(n2187) );
  NAND U3245 ( .A(n2182), .B(n2181), .Z(n2183) );
  XNOR U3246 ( .A(n2184), .B(n2183), .Z(n2195) );
  XNOR U3247 ( .A(n2195), .B(n2185), .Z(n2186) );
  XNOR U3248 ( .A(n2187), .B(n2186), .Z(n2191) );
  XNOR U3249 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U3250 ( .A(n2191), .B(n2190), .Z(n2199) );
  XNOR U3251 ( .A(n2198), .B(n2199), .Z(z[1]) );
  AND U3252 ( .A(n2193), .B(n2192), .Z(n2197) );
  XNOR U3253 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U3254 ( .A(n2197), .B(n2196), .Z(n2202) );
  XNOR U3255 ( .A(n2198), .B(n2202), .Z(z[6]) );
  XOR U3256 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3257 ( .A(n2202), .B(n2201), .Z(z[3]) );
  XNOR U3258 ( .A(x[8]), .B(x[14]), .Z(n2203) );
  XNOR U3259 ( .A(x[13]), .B(n2203), .Z(n2301) );
  XNOR U3260 ( .A(n2301), .B(x[15]), .Z(n2266) );
  XNOR U3261 ( .A(x[10]), .B(n2266), .Z(n2218) );
  XOR U3262 ( .A(x[9]), .B(n2218), .Z(n2252) );
  XOR U3263 ( .A(x[11]), .B(x[9]), .Z(n2205) );
  XOR U3264 ( .A(n2203), .B(x[10]), .Z(n2204) );
  XOR U3265 ( .A(n2205), .B(n2204), .Z(n2306) );
  XNOR U3266 ( .A(x[8]), .B(n2306), .Z(n2257) );
  XOR U3267 ( .A(x[15]), .B(x[12]), .Z(n2241) );
  AND U3268 ( .A(n2257), .B(n2241), .Z(n2209) );
  XOR U3269 ( .A(x[10]), .B(x[15]), .Z(n2268) );
  XNOR U3270 ( .A(n2205), .B(n2241), .Z(n2221) );
  IV U3271 ( .A(n2221), .Z(n2261) );
  XNOR U3272 ( .A(x[8]), .B(n2261), .Z(n2264) );
  XNOR U3273 ( .A(n2301), .B(n2264), .Z(n2296) );
  NAND U3274 ( .A(n2268), .B(n2296), .Z(n2206) );
  XNOR U3275 ( .A(n2209), .B(n2206), .Z(n2220) );
  NAND U3276 ( .A(n2306), .B(n2266), .Z(n2207) );
  IV U3277 ( .A(n2301), .Z(n2211) );
  XOR U3278 ( .A(n2306), .B(n2211), .Z(n2278) );
  XOR U3279 ( .A(x[9]), .B(x[15]), .Z(n2273) );
  NAND U3280 ( .A(n2278), .B(n2273), .Z(n2210) );
  XNOR U3281 ( .A(n2207), .B(n2210), .Z(n2208) );
  XNOR U3282 ( .A(n2220), .B(n2208), .Z(n2244) );
  XOR U3283 ( .A(x[10]), .B(x[12]), .Z(n2250) );
  XNOR U3284 ( .A(n2221), .B(n2278), .Z(n2258) );
  IV U3285 ( .A(n2228), .Z(n2246) );
  NANDN U3286 ( .A(n2244), .B(n2246), .Z(n2230) );
  XNOR U3287 ( .A(x[12]), .B(n2211), .Z(n2276) );
  NOR U3288 ( .A(n2276), .B(x[8]), .Z(n2212) );
  XOR U3289 ( .A(n2212), .B(n2252), .Z(n2213) );
  NANDN U3290 ( .A(n2221), .B(n2213), .Z(n2216) );
  ANDN U3291 ( .B(x[8]), .A(n2276), .Z(n2214) );
  NAND U3292 ( .A(n2221), .B(n2214), .Z(n2215) );
  NAND U3293 ( .A(n2216), .B(n2215), .Z(n2217) );
  XNOR U3294 ( .A(n2218), .B(n2217), .Z(n2219) );
  XOR U3295 ( .A(n2220), .B(n2219), .Z(n2243) );
  IV U3296 ( .A(n2244), .Z(n2236) );
  ANDN U3297 ( .B(n2243), .A(n2236), .Z(n2226) );
  AND U3298 ( .A(n2276), .B(n2221), .Z(n2223) );
  NANDN U3299 ( .A(n2252), .B(x[8]), .Z(n2222) );
  XNOR U3300 ( .A(n2223), .B(n2222), .Z(n2224) );
  XNOR U3301 ( .A(n2225), .B(n2224), .Z(n2248) );
  XNOR U3302 ( .A(n2226), .B(n2248), .Z(n2227) );
  NAND U3303 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U3304 ( .A(n2230), .B(n2229), .Z(n2242) );
  AND U3305 ( .A(n2252), .B(n2242), .Z(n2255) );
  NANDN U3306 ( .A(n2244), .B(n2243), .Z(n2231) );
  NAND U3307 ( .A(n2246), .B(n2231), .Z(n2234) );
  IV U3308 ( .A(n2248), .Z(n2237) );
  XOR U3309 ( .A(n2243), .B(n2237), .Z(n2232) );
  NAND U3310 ( .A(n2244), .B(n2232), .Z(n2233) );
  AND U3311 ( .A(n2234), .B(n2233), .Z(n2294) );
  XNOR U3312 ( .A(n2246), .B(n2236), .Z(n2235) );
  NAND U3313 ( .A(n2237), .B(n2235), .Z(n2240) );
  NANDN U3314 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U3315 ( .A(n2243), .B(n2238), .Z(n2239) );
  NAND U3316 ( .A(n2240), .B(n2239), .Z(n2307) );
  XOR U3317 ( .A(n2294), .B(n2307), .Z(n2256) );
  NAND U3318 ( .A(n2241), .B(n2256), .Z(n2270) );
  IV U3319 ( .A(n2242), .Z(n2263) );
  NAND U3320 ( .A(n2248), .B(n2243), .Z(n2272) );
  NAND U3321 ( .A(n2244), .B(n2243), .Z(n2245) );
  XNOR U3322 ( .A(n2246), .B(n2245), .Z(n2247) );
  NANDN U3323 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U3324 ( .A(n2272), .B(n2249), .Z(n2303) );
  XOR U3325 ( .A(n2263), .B(n2303), .Z(n2267) );
  XNOR U3326 ( .A(n2256), .B(n2267), .Z(n2259) );
  NAND U3327 ( .A(n2259), .B(n2250), .Z(n2251) );
  XOR U3328 ( .A(n2270), .B(n2251), .Z(n2312) );
  XNOR U3329 ( .A(n2294), .B(n2263), .Z(n2262) );
  XOR U3330 ( .A(n2276), .B(n2252), .Z(n2253) );
  AND U3331 ( .A(n2262), .B(n2253), .Z(n2280) );
  XNOR U3332 ( .A(n2312), .B(n2280), .Z(n2254) );
  XNOR U3333 ( .A(n2255), .B(n2254), .Z(n2287) );
  AND U3334 ( .A(n2257), .B(n2256), .Z(n2295) );
  NAND U3335 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U3336 ( .A(n2295), .B(n2260), .Z(n2283) );
  AND U3337 ( .A(n2262), .B(n2261), .Z(n2298) );
  OR U3338 ( .A(n2264), .B(n2263), .Z(n2265) );
  XNOR U3339 ( .A(n2298), .B(n2265), .Z(n2293) );
  XNOR U3340 ( .A(n2287), .B(n3960), .Z(n2291) );
  ANDN U3341 ( .B(n2307), .A(n2266), .Z(n2275) );
  IV U3342 ( .A(n2267), .Z(n2297) );
  NAND U3343 ( .A(n2297), .B(n2268), .Z(n2269) );
  XNOR U3344 ( .A(n2270), .B(n2269), .Z(n2286) );
  NAND U3345 ( .A(n2307), .B(n2303), .Z(n2271) );
  AND U3346 ( .A(n2272), .B(n2271), .Z(n2277) );
  AND U3347 ( .A(n2273), .B(n2277), .Z(n2305) );
  XOR U3348 ( .A(n2286), .B(n2305), .Z(n2274) );
  XNOR U3349 ( .A(n2275), .B(n2274), .Z(n2289) );
  XNOR U3350 ( .A(n2291), .B(n2289), .Z(z[14]) );
  AND U3351 ( .A(n2276), .B(n2294), .Z(n2282) );
  AND U3352 ( .A(n2278), .B(n2277), .Z(n2308) );
  NAND U3353 ( .A(n2301), .B(n2303), .Z(n2279) );
  XNOR U3354 ( .A(n2308), .B(n2279), .Z(n2292) );
  XNOR U3355 ( .A(n2280), .B(n2292), .Z(n2281) );
  XNOR U3356 ( .A(n2282), .B(n2281), .Z(n2284) );
  XNOR U3357 ( .A(n2284), .B(n2283), .Z(n2285) );
  XNOR U3358 ( .A(n2286), .B(n2285), .Z(n2290) );
  XOR U3359 ( .A(n2287), .B(n2290), .Z(n2288) );
  XNOR U3360 ( .A(n2289), .B(n2288), .Z(z[11]) );
  XNOR U3361 ( .A(n2291), .B(n2290), .Z(z[9]) );
  XNOR U3362 ( .A(n2293), .B(n2292), .Z(z[10]) );
  AND U3363 ( .A(x[8]), .B(n2294), .Z(n2300) );
  XOR U3364 ( .A(n2309), .B(n2298), .Z(n2299) );
  XNOR U3365 ( .A(n2300), .B(n2299), .Z(n3929) );
  XOR U3366 ( .A(x[9]), .B(n2301), .Z(n2302) );
  NAND U3367 ( .A(n2303), .B(n2302), .Z(n2304) );
  XNOR U3368 ( .A(n2305), .B(n2304), .Z(n2314) );
  ANDN U3369 ( .B(n2307), .A(n2306), .Z(n2311) );
  XOR U3370 ( .A(n2309), .B(n2308), .Z(n2310) );
  XNOR U3371 ( .A(n2311), .B(n2310), .Z(n3961) );
  XNOR U3372 ( .A(n2312), .B(n3961), .Z(n2313) );
  XNOR U3373 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U3374 ( .A(n3929), .B(n2315), .Z(z[13]) );
  XOR U3375 ( .A(x[17]), .B(x[19]), .Z(n2319) );
  XOR U3376 ( .A(x[16]), .B(x[22]), .Z(n2317) );
  XNOR U3377 ( .A(n2319), .B(n2317), .Z(n2316) );
  XNOR U3378 ( .A(x[18]), .B(n2316), .Z(n2387) );
  IV U3379 ( .A(n2387), .Z(n2321) );
  XNOR U3380 ( .A(x[16]), .B(n2321), .Z(n2369) );
  XNOR U3381 ( .A(x[20]), .B(x[23]), .Z(n2318) );
  IV U3382 ( .A(n2318), .Z(n2382) );
  AND U3383 ( .A(n2369), .B(n2382), .Z(n2326) );
  XOR U3384 ( .A(x[23]), .B(x[18]), .Z(n2409) );
  XNOR U3385 ( .A(n2317), .B(x[21]), .Z(n2332) );
  IV U3386 ( .A(n2332), .Z(n2378) );
  XOR U3387 ( .A(n2319), .B(n2318), .Z(n2343) );
  IV U3388 ( .A(n2343), .Z(n2358) );
  XNOR U3389 ( .A(n2358), .B(x[16]), .Z(n2359) );
  XNOR U3390 ( .A(n2378), .B(n2359), .Z(n2371) );
  NAND U3391 ( .A(n2409), .B(n2371), .Z(n2320) );
  XNOR U3392 ( .A(n2326), .B(n2320), .Z(n2339) );
  XOR U3393 ( .A(x[17]), .B(x[23]), .Z(n2377) );
  XOR U3394 ( .A(n2321), .B(n2378), .Z(n2367) );
  ANDN U3395 ( .B(n2377), .A(n2367), .Z(n2328) );
  XOR U3396 ( .A(x[23]), .B(n2378), .Z(n2420) );
  IV U3397 ( .A(n2420), .Z(n2331) );
  NAND U3398 ( .A(n2321), .B(n2331), .Z(n2322) );
  XOR U3399 ( .A(n2328), .B(n2322), .Z(n2323) );
  XNOR U3400 ( .A(n2339), .B(n2323), .Z(n2363) );
  NANDN U3401 ( .A(x[17]), .B(n2332), .Z(n2330) );
  XNOR U3402 ( .A(n2358), .B(n2367), .Z(n2402) );
  XOR U3403 ( .A(x[20]), .B(x[18]), .Z(n2385) );
  AND U3404 ( .A(n2402), .B(n2385), .Z(n2325) );
  XNOR U3405 ( .A(n2387), .B(n2420), .Z(n2324) );
  XNOR U3406 ( .A(n2325), .B(n2324), .Z(n2327) );
  XOR U3407 ( .A(n2327), .B(n2326), .Z(n2347) );
  XNOR U3408 ( .A(n2328), .B(n2347), .Z(n2329) );
  XNOR U3409 ( .A(n2330), .B(n2329), .Z(n2361) );
  IV U3410 ( .A(n2361), .Z(n2364) );
  NAND U3411 ( .A(n2363), .B(n2364), .Z(n2357) );
  NANDN U3412 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U3413 ( .A(x[18]), .B(n2331), .Z(n2338) );
  XNOR U3414 ( .A(x[17]), .B(n2338), .Z(n2342) );
  IV U3415 ( .A(n2342), .Z(n2396) );
  XNOR U3416 ( .A(x[20]), .B(n2332), .Z(n2408) );
  OR U3417 ( .A(x[16]), .B(n2408), .Z(n2333) );
  XNOR U3418 ( .A(n2396), .B(n2333), .Z(n2334) );
  NANDN U3419 ( .A(n2343), .B(n2334), .Z(n2337) );
  ANDN U3420 ( .B(x[16]), .A(n2408), .Z(n2335) );
  NAND U3421 ( .A(n2343), .B(n2335), .Z(n2336) );
  NAND U3422 ( .A(n2337), .B(n2336), .Z(n2341) );
  XNOR U3423 ( .A(n2339), .B(n2338), .Z(n2340) );
  XOR U3424 ( .A(n2341), .B(n2340), .Z(n2365) );
  IV U3425 ( .A(n2363), .Z(n2362) );
  ANDN U3426 ( .B(n2365), .A(n2362), .Z(n2348) );
  AND U3427 ( .A(x[16]), .B(n2342), .Z(n2345) );
  NAND U3428 ( .A(n2343), .B(n2408), .Z(n2344) );
  XNOR U3429 ( .A(n2345), .B(n2344), .Z(n2346) );
  XNOR U3430 ( .A(n2347), .B(n2346), .Z(n2366) );
  XNOR U3431 ( .A(n2348), .B(n2366), .Z(n2349) );
  NAND U3432 ( .A(n2361), .B(n2349), .Z(n2350) );
  NAND U3433 ( .A(n2351), .B(n2350), .Z(n2395) );
  IV U3434 ( .A(n2395), .Z(n2370) );
  OR U3435 ( .A(n2365), .B(n2361), .Z(n2352) );
  NAND U3436 ( .A(n2362), .B(n2352), .Z(n2355) );
  XOR U3437 ( .A(n2365), .B(n2366), .Z(n2353) );
  NANDN U3438 ( .A(n2364), .B(n2353), .Z(n2354) );
  NAND U3439 ( .A(n2355), .B(n2354), .Z(n2407) );
  NANDN U3440 ( .A(n2370), .B(n2407), .Z(n2356) );
  AND U3441 ( .A(n2357), .B(n2356), .Z(n2398) );
  AND U3442 ( .A(n2398), .B(n2358), .Z(n2373) );
  OR U3443 ( .A(n2359), .B(n2370), .Z(n2360) );
  XNOR U3444 ( .A(n2373), .B(n2360), .Z(n2406) );
  XOR U3445 ( .A(n2421), .B(n2380), .Z(n2376) );
  ANDN U3446 ( .B(n2376), .A(n2367), .Z(n2388) );
  NAND U3447 ( .A(n2378), .B(n2380), .Z(n2368) );
  XNOR U3448 ( .A(n2388), .B(n2368), .Z(n2413) );
  XNOR U3449 ( .A(n2406), .B(n2413), .Z(z[18]) );
  AND U3450 ( .A(x[16]), .B(n2407), .Z(n2375) );
  AND U3451 ( .A(n2369), .B(n2384), .Z(n2405) );
  XOR U3452 ( .A(n2370), .B(n2380), .Z(n2383) );
  IV U3453 ( .A(n2383), .Z(n2410) );
  NAND U3454 ( .A(n2410), .B(n2371), .Z(n2372) );
  XNOR U3455 ( .A(n2405), .B(n2372), .Z(n2389) );
  XNOR U3456 ( .A(n2373), .B(n2389), .Z(n2374) );
  XNOR U3457 ( .A(n2375), .B(n2374), .Z(n3932) );
  AND U3458 ( .A(n2377), .B(n2376), .Z(n2422) );
  XOR U3459 ( .A(x[17]), .B(n2378), .Z(n2379) );
  NAND U3460 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U3461 ( .A(n2422), .B(n2381), .Z(n2393) );
  AND U3462 ( .A(n2384), .B(n2382), .Z(n2412) );
  XNOR U3463 ( .A(n2384), .B(n2383), .Z(n2403) );
  NAND U3464 ( .A(n2403), .B(n2385), .Z(n2386) );
  XNOR U3465 ( .A(n2412), .B(n2386), .Z(n2399) );
  AND U3466 ( .A(n2421), .B(n2387), .Z(n2391) );
  XNOR U3467 ( .A(n2389), .B(n2388), .Z(n2390) );
  XNOR U3468 ( .A(n2391), .B(n2390), .Z(n3931) );
  XNOR U3469 ( .A(n2399), .B(n3931), .Z(n2392) );
  XNOR U3470 ( .A(n2393), .B(n2392), .Z(n2394) );
  XNOR U3471 ( .A(n3932), .B(n2394), .Z(z[21]) );
  AND U3472 ( .A(n2396), .B(n2395), .Z(n2401) );
  XOR U3473 ( .A(n2396), .B(n2408), .Z(n2397) );
  AND U3474 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U3475 ( .A(n2399), .B(n2417), .Z(n2400) );
  XNOR U3476 ( .A(n2401), .B(n2400), .Z(n2428) );
  NAND U3477 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U3478 ( .A(n2405), .B(n2404), .Z(n2416) );
  XNOR U3479 ( .A(n2406), .B(n2416), .Z(n3930) );
  XNOR U3480 ( .A(n2428), .B(n3930), .Z(n2426) );
  AND U3481 ( .A(n2408), .B(n2407), .Z(n2415) );
  NAND U3482 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U3483 ( .A(n2412), .B(n2411), .Z(n2423) );
  XNOR U3484 ( .A(n2423), .B(n2413), .Z(n2414) );
  XNOR U3485 ( .A(n2415), .B(n2414), .Z(n2419) );
  XNOR U3486 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U3487 ( .A(n2419), .B(n2418), .Z(n2427) );
  XNOR U3488 ( .A(n2426), .B(n2427), .Z(z[17]) );
  AND U3489 ( .A(n2421), .B(n2420), .Z(n2425) );
  XNOR U3490 ( .A(n2423), .B(n2422), .Z(n2424) );
  XNOR U3491 ( .A(n2425), .B(n2424), .Z(n2430) );
  XNOR U3492 ( .A(n2426), .B(n2430), .Z(z[22]) );
  XOR U3493 ( .A(n2428), .B(n2427), .Z(n2429) );
  XNOR U3494 ( .A(n2430), .B(n2429), .Z(z[19]) );
  XOR U3495 ( .A(x[25]), .B(x[27]), .Z(n2434) );
  XOR U3496 ( .A(x[24]), .B(x[30]), .Z(n2432) );
  XNOR U3497 ( .A(n2434), .B(n2432), .Z(n2431) );
  XNOR U3498 ( .A(x[26]), .B(n2431), .Z(n2502) );
  IV U3499 ( .A(n2502), .Z(n2436) );
  XNOR U3500 ( .A(x[24]), .B(n2436), .Z(n2484) );
  XNOR U3501 ( .A(x[28]), .B(x[31]), .Z(n2433) );
  IV U3502 ( .A(n2433), .Z(n2497) );
  AND U3503 ( .A(n2484), .B(n2497), .Z(n2441) );
  XOR U3504 ( .A(x[31]), .B(x[26]), .Z(n2524) );
  XNOR U3505 ( .A(n2432), .B(x[29]), .Z(n2447) );
  IV U3506 ( .A(n2447), .Z(n2493) );
  XOR U3507 ( .A(n2434), .B(n2433), .Z(n2458) );
  IV U3508 ( .A(n2458), .Z(n2473) );
  XNOR U3509 ( .A(n2473), .B(x[24]), .Z(n2474) );
  XNOR U3510 ( .A(n2493), .B(n2474), .Z(n2486) );
  NAND U3511 ( .A(n2524), .B(n2486), .Z(n2435) );
  XNOR U3512 ( .A(n2441), .B(n2435), .Z(n2454) );
  XOR U3513 ( .A(x[25]), .B(x[31]), .Z(n2492) );
  XOR U3514 ( .A(n2436), .B(n2493), .Z(n2482) );
  ANDN U3515 ( .B(n2492), .A(n2482), .Z(n2443) );
  XOR U3516 ( .A(x[31]), .B(n2493), .Z(n2535) );
  IV U3517 ( .A(n2535), .Z(n2446) );
  NAND U3518 ( .A(n2436), .B(n2446), .Z(n2437) );
  XOR U3519 ( .A(n2443), .B(n2437), .Z(n2438) );
  XNOR U3520 ( .A(n2454), .B(n2438), .Z(n2478) );
  NANDN U3521 ( .A(x[25]), .B(n2447), .Z(n2445) );
  XNOR U3522 ( .A(n2473), .B(n2482), .Z(n2517) );
  XOR U3523 ( .A(x[28]), .B(x[26]), .Z(n2500) );
  AND U3524 ( .A(n2517), .B(n2500), .Z(n2440) );
  XNOR U3525 ( .A(n2502), .B(n2535), .Z(n2439) );
  XNOR U3526 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U3527 ( .A(n2442), .B(n2441), .Z(n2462) );
  XNOR U3528 ( .A(n2443), .B(n2462), .Z(n2444) );
  XNOR U3529 ( .A(n2445), .B(n2444), .Z(n2476) );
  IV U3530 ( .A(n2476), .Z(n2479) );
  NAND U3531 ( .A(n2478), .B(n2479), .Z(n2472) );
  NANDN U3532 ( .A(n2478), .B(n2479), .Z(n2466) );
  XNOR U3533 ( .A(x[26]), .B(n2446), .Z(n2453) );
  XNOR U3534 ( .A(x[25]), .B(n2453), .Z(n2457) );
  IV U3535 ( .A(n2457), .Z(n2511) );
  XNOR U3536 ( .A(x[28]), .B(n2447), .Z(n2523) );
  OR U3537 ( .A(x[24]), .B(n2523), .Z(n2448) );
  XNOR U3538 ( .A(n2511), .B(n2448), .Z(n2449) );
  NANDN U3539 ( .A(n2458), .B(n2449), .Z(n2452) );
  ANDN U3540 ( .B(x[24]), .A(n2523), .Z(n2450) );
  NAND U3541 ( .A(n2458), .B(n2450), .Z(n2451) );
  NAND U3542 ( .A(n2452), .B(n2451), .Z(n2456) );
  XNOR U3543 ( .A(n2454), .B(n2453), .Z(n2455) );
  XOR U3544 ( .A(n2456), .B(n2455), .Z(n2480) );
  IV U3545 ( .A(n2478), .Z(n2477) );
  ANDN U3546 ( .B(n2480), .A(n2477), .Z(n2463) );
  AND U3547 ( .A(x[24]), .B(n2457), .Z(n2460) );
  NAND U3548 ( .A(n2458), .B(n2523), .Z(n2459) );
  XNOR U3549 ( .A(n2460), .B(n2459), .Z(n2461) );
  XNOR U3550 ( .A(n2462), .B(n2461), .Z(n2481) );
  XNOR U3551 ( .A(n2463), .B(n2481), .Z(n2464) );
  NAND U3552 ( .A(n2476), .B(n2464), .Z(n2465) );
  NAND U3553 ( .A(n2466), .B(n2465), .Z(n2510) );
  IV U3554 ( .A(n2510), .Z(n2485) );
  OR U3555 ( .A(n2480), .B(n2476), .Z(n2467) );
  NAND U3556 ( .A(n2477), .B(n2467), .Z(n2470) );
  XOR U3557 ( .A(n2480), .B(n2481), .Z(n2468) );
  NANDN U3558 ( .A(n2479), .B(n2468), .Z(n2469) );
  NAND U3559 ( .A(n2470), .B(n2469), .Z(n2522) );
  NANDN U3560 ( .A(n2485), .B(n2522), .Z(n2471) );
  AND U3561 ( .A(n2472), .B(n2471), .Z(n2513) );
  AND U3562 ( .A(n2513), .B(n2473), .Z(n2488) );
  OR U3563 ( .A(n2474), .B(n2485), .Z(n2475) );
  XNOR U3564 ( .A(n2488), .B(n2475), .Z(n2521) );
  XOR U3565 ( .A(n2536), .B(n2495), .Z(n2491) );
  ANDN U3566 ( .B(n2491), .A(n2482), .Z(n2503) );
  NAND U3567 ( .A(n2493), .B(n2495), .Z(n2483) );
  XNOR U3568 ( .A(n2503), .B(n2483), .Z(n2528) );
  XNOR U3569 ( .A(n2521), .B(n2528), .Z(z[26]) );
  AND U3570 ( .A(x[24]), .B(n2522), .Z(n2490) );
  AND U3571 ( .A(n2484), .B(n2499), .Z(n2520) );
  XOR U3572 ( .A(n2485), .B(n2495), .Z(n2498) );
  IV U3573 ( .A(n2498), .Z(n2525) );
  NAND U3574 ( .A(n2525), .B(n2486), .Z(n2487) );
  XNOR U3575 ( .A(n2520), .B(n2487), .Z(n2504) );
  XNOR U3576 ( .A(n2488), .B(n2504), .Z(n2489) );
  XNOR U3577 ( .A(n2490), .B(n2489), .Z(n3935) );
  AND U3578 ( .A(n2492), .B(n2491), .Z(n2537) );
  XOR U3579 ( .A(x[25]), .B(n2493), .Z(n2494) );
  NAND U3580 ( .A(n2495), .B(n2494), .Z(n2496) );
  XNOR U3581 ( .A(n2537), .B(n2496), .Z(n2508) );
  AND U3582 ( .A(n2499), .B(n2497), .Z(n2527) );
  XNOR U3583 ( .A(n2499), .B(n2498), .Z(n2518) );
  NAND U3584 ( .A(n2518), .B(n2500), .Z(n2501) );
  XNOR U3585 ( .A(n2527), .B(n2501), .Z(n2514) );
  AND U3586 ( .A(n2536), .B(n2502), .Z(n2506) );
  XNOR U3587 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3588 ( .A(n2506), .B(n2505), .Z(n3934) );
  XNOR U3589 ( .A(n2514), .B(n3934), .Z(n2507) );
  XNOR U3590 ( .A(n2508), .B(n2507), .Z(n2509) );
  XNOR U3591 ( .A(n3935), .B(n2509), .Z(z[29]) );
  AND U3592 ( .A(n2511), .B(n2510), .Z(n2516) );
  XOR U3593 ( .A(n2511), .B(n2523), .Z(n2512) );
  AND U3594 ( .A(n2513), .B(n2512), .Z(n2532) );
  XNOR U3595 ( .A(n2514), .B(n2532), .Z(n2515) );
  XNOR U3596 ( .A(n2516), .B(n2515), .Z(n2543) );
  NAND U3597 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U3598 ( .A(n2520), .B(n2519), .Z(n2531) );
  XNOR U3599 ( .A(n2521), .B(n2531), .Z(n3933) );
  XNOR U3600 ( .A(n2543), .B(n3933), .Z(n2541) );
  AND U3601 ( .A(n2523), .B(n2522), .Z(n2530) );
  NAND U3602 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3603 ( .A(n2527), .B(n2526), .Z(n2538) );
  XNOR U3604 ( .A(n2538), .B(n2528), .Z(n2529) );
  XNOR U3605 ( .A(n2530), .B(n2529), .Z(n2534) );
  XNOR U3606 ( .A(n2532), .B(n2531), .Z(n2533) );
  XNOR U3607 ( .A(n2534), .B(n2533), .Z(n2542) );
  XNOR U3608 ( .A(n2541), .B(n2542), .Z(z[25]) );
  AND U3609 ( .A(n2536), .B(n2535), .Z(n2540) );
  XNOR U3610 ( .A(n2538), .B(n2537), .Z(n2539) );
  XNOR U3611 ( .A(n2540), .B(n2539), .Z(n2545) );
  XNOR U3612 ( .A(n2541), .B(n2545), .Z(z[30]) );
  XOR U3613 ( .A(n2543), .B(n2542), .Z(n2544) );
  XNOR U3614 ( .A(n2545), .B(n2544), .Z(z[27]) );
  XOR U3615 ( .A(x[33]), .B(x[35]), .Z(n2549) );
  XOR U3616 ( .A(x[32]), .B(x[38]), .Z(n2547) );
  XNOR U3617 ( .A(n2549), .B(n2547), .Z(n2546) );
  XNOR U3618 ( .A(x[34]), .B(n2546), .Z(n2617) );
  IV U3619 ( .A(n2617), .Z(n2551) );
  XNOR U3620 ( .A(x[32]), .B(n2551), .Z(n2599) );
  XNOR U3621 ( .A(x[36]), .B(x[39]), .Z(n2548) );
  IV U3622 ( .A(n2548), .Z(n2612) );
  AND U3623 ( .A(n2599), .B(n2612), .Z(n2556) );
  XOR U3624 ( .A(x[39]), .B(x[34]), .Z(n2639) );
  XNOR U3625 ( .A(n2547), .B(x[37]), .Z(n2562) );
  IV U3626 ( .A(n2562), .Z(n2608) );
  XOR U3627 ( .A(n2549), .B(n2548), .Z(n2573) );
  IV U3628 ( .A(n2573), .Z(n2588) );
  XNOR U3629 ( .A(n2588), .B(x[32]), .Z(n2589) );
  XNOR U3630 ( .A(n2608), .B(n2589), .Z(n2601) );
  NAND U3631 ( .A(n2639), .B(n2601), .Z(n2550) );
  XNOR U3632 ( .A(n2556), .B(n2550), .Z(n2569) );
  XOR U3633 ( .A(x[33]), .B(x[39]), .Z(n2607) );
  XOR U3634 ( .A(n2551), .B(n2608), .Z(n2597) );
  ANDN U3635 ( .B(n2607), .A(n2597), .Z(n2558) );
  XOR U3636 ( .A(x[39]), .B(n2608), .Z(n2650) );
  IV U3637 ( .A(n2650), .Z(n2561) );
  NAND U3638 ( .A(n2551), .B(n2561), .Z(n2552) );
  XOR U3639 ( .A(n2558), .B(n2552), .Z(n2553) );
  XNOR U3640 ( .A(n2569), .B(n2553), .Z(n2593) );
  NANDN U3641 ( .A(x[33]), .B(n2562), .Z(n2560) );
  XNOR U3642 ( .A(n2588), .B(n2597), .Z(n2632) );
  XOR U3643 ( .A(x[36]), .B(x[34]), .Z(n2615) );
  AND U3644 ( .A(n2632), .B(n2615), .Z(n2555) );
  XNOR U3645 ( .A(n2617), .B(n2650), .Z(n2554) );
  XNOR U3646 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U3647 ( .A(n2557), .B(n2556), .Z(n2577) );
  XNOR U3648 ( .A(n2558), .B(n2577), .Z(n2559) );
  XNOR U3649 ( .A(n2560), .B(n2559), .Z(n2591) );
  IV U3650 ( .A(n2591), .Z(n2594) );
  NAND U3651 ( .A(n2593), .B(n2594), .Z(n2587) );
  NANDN U3652 ( .A(n2593), .B(n2594), .Z(n2581) );
  XNOR U3653 ( .A(x[34]), .B(n2561), .Z(n2568) );
  XNOR U3654 ( .A(x[33]), .B(n2568), .Z(n2572) );
  IV U3655 ( .A(n2572), .Z(n2626) );
  XNOR U3656 ( .A(x[36]), .B(n2562), .Z(n2638) );
  OR U3657 ( .A(x[32]), .B(n2638), .Z(n2563) );
  XNOR U3658 ( .A(n2626), .B(n2563), .Z(n2564) );
  NANDN U3659 ( .A(n2573), .B(n2564), .Z(n2567) );
  ANDN U3660 ( .B(x[32]), .A(n2638), .Z(n2565) );
  NAND U3661 ( .A(n2573), .B(n2565), .Z(n2566) );
  NAND U3662 ( .A(n2567), .B(n2566), .Z(n2571) );
  XNOR U3663 ( .A(n2569), .B(n2568), .Z(n2570) );
  XOR U3664 ( .A(n2571), .B(n2570), .Z(n2595) );
  IV U3665 ( .A(n2593), .Z(n2592) );
  ANDN U3666 ( .B(n2595), .A(n2592), .Z(n2578) );
  AND U3667 ( .A(x[32]), .B(n2572), .Z(n2575) );
  NAND U3668 ( .A(n2573), .B(n2638), .Z(n2574) );
  XNOR U3669 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U3670 ( .A(n2577), .B(n2576), .Z(n2596) );
  XNOR U3671 ( .A(n2578), .B(n2596), .Z(n2579) );
  NAND U3672 ( .A(n2591), .B(n2579), .Z(n2580) );
  NAND U3673 ( .A(n2581), .B(n2580), .Z(n2625) );
  IV U3674 ( .A(n2625), .Z(n2600) );
  OR U3675 ( .A(n2595), .B(n2591), .Z(n2582) );
  NAND U3676 ( .A(n2592), .B(n2582), .Z(n2585) );
  XOR U3677 ( .A(n2595), .B(n2596), .Z(n2583) );
  NANDN U3678 ( .A(n2594), .B(n2583), .Z(n2584) );
  NAND U3679 ( .A(n2585), .B(n2584), .Z(n2637) );
  NANDN U3680 ( .A(n2600), .B(n2637), .Z(n2586) );
  AND U3681 ( .A(n2587), .B(n2586), .Z(n2628) );
  AND U3682 ( .A(n2628), .B(n2588), .Z(n2603) );
  OR U3683 ( .A(n2589), .B(n2600), .Z(n2590) );
  XNOR U3684 ( .A(n2603), .B(n2590), .Z(n2636) );
  XOR U3685 ( .A(n2651), .B(n2610), .Z(n2606) );
  ANDN U3686 ( .B(n2606), .A(n2597), .Z(n2618) );
  NAND U3687 ( .A(n2608), .B(n2610), .Z(n2598) );
  XNOR U3688 ( .A(n2618), .B(n2598), .Z(n2643) );
  XNOR U3689 ( .A(n2636), .B(n2643), .Z(z[34]) );
  AND U3690 ( .A(x[32]), .B(n2637), .Z(n2605) );
  AND U3691 ( .A(n2599), .B(n2614), .Z(n2635) );
  XOR U3692 ( .A(n2600), .B(n2610), .Z(n2613) );
  IV U3693 ( .A(n2613), .Z(n2640) );
  NAND U3694 ( .A(n2640), .B(n2601), .Z(n2602) );
  XNOR U3695 ( .A(n2635), .B(n2602), .Z(n2619) );
  XNOR U3696 ( .A(n2603), .B(n2619), .Z(n2604) );
  XNOR U3697 ( .A(n2605), .B(n2604), .Z(n3938) );
  AND U3698 ( .A(n2607), .B(n2606), .Z(n2652) );
  XOR U3699 ( .A(x[33]), .B(n2608), .Z(n2609) );
  NAND U3700 ( .A(n2610), .B(n2609), .Z(n2611) );
  XNOR U3701 ( .A(n2652), .B(n2611), .Z(n2623) );
  AND U3702 ( .A(n2614), .B(n2612), .Z(n2642) );
  XNOR U3703 ( .A(n2614), .B(n2613), .Z(n2633) );
  NAND U3704 ( .A(n2633), .B(n2615), .Z(n2616) );
  XNOR U3705 ( .A(n2642), .B(n2616), .Z(n2629) );
  AND U3706 ( .A(n2651), .B(n2617), .Z(n2621) );
  XNOR U3707 ( .A(n2619), .B(n2618), .Z(n2620) );
  XNOR U3708 ( .A(n2621), .B(n2620), .Z(n3937) );
  XNOR U3709 ( .A(n2629), .B(n3937), .Z(n2622) );
  XNOR U3710 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U3711 ( .A(n3938), .B(n2624), .Z(z[37]) );
  AND U3712 ( .A(n2626), .B(n2625), .Z(n2631) );
  XOR U3713 ( .A(n2626), .B(n2638), .Z(n2627) );
  AND U3714 ( .A(n2628), .B(n2627), .Z(n2647) );
  XNOR U3715 ( .A(n2629), .B(n2647), .Z(n2630) );
  XNOR U3716 ( .A(n2631), .B(n2630), .Z(n2658) );
  NAND U3717 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U3718 ( .A(n2635), .B(n2634), .Z(n2646) );
  XNOR U3719 ( .A(n2636), .B(n2646), .Z(n3936) );
  XNOR U3720 ( .A(n2658), .B(n3936), .Z(n2656) );
  AND U3721 ( .A(n2638), .B(n2637), .Z(n2645) );
  NAND U3722 ( .A(n2640), .B(n2639), .Z(n2641) );
  XNOR U3723 ( .A(n2642), .B(n2641), .Z(n2653) );
  XNOR U3724 ( .A(n2653), .B(n2643), .Z(n2644) );
  XNOR U3725 ( .A(n2645), .B(n2644), .Z(n2649) );
  XNOR U3726 ( .A(n2647), .B(n2646), .Z(n2648) );
  XNOR U3727 ( .A(n2649), .B(n2648), .Z(n2657) );
  XNOR U3728 ( .A(n2656), .B(n2657), .Z(z[33]) );
  AND U3729 ( .A(n2651), .B(n2650), .Z(n2655) );
  XNOR U3730 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3731 ( .A(n2655), .B(n2654), .Z(n2660) );
  XNOR U3732 ( .A(n2656), .B(n2660), .Z(z[38]) );
  XOR U3733 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U3734 ( .A(n2660), .B(n2659), .Z(z[35]) );
  XOR U3735 ( .A(x[41]), .B(x[43]), .Z(n2664) );
  XOR U3736 ( .A(x[40]), .B(x[46]), .Z(n2662) );
  XNOR U3737 ( .A(n2664), .B(n2662), .Z(n2661) );
  XNOR U3738 ( .A(x[42]), .B(n2661), .Z(n2732) );
  IV U3739 ( .A(n2732), .Z(n2666) );
  XNOR U3740 ( .A(x[40]), .B(n2666), .Z(n2714) );
  XNOR U3741 ( .A(x[44]), .B(x[47]), .Z(n2663) );
  IV U3742 ( .A(n2663), .Z(n2727) );
  AND U3743 ( .A(n2714), .B(n2727), .Z(n2671) );
  XOR U3744 ( .A(x[47]), .B(x[42]), .Z(n2754) );
  XNOR U3745 ( .A(n2662), .B(x[45]), .Z(n2677) );
  IV U3746 ( .A(n2677), .Z(n2723) );
  XOR U3747 ( .A(n2664), .B(n2663), .Z(n2688) );
  IV U3748 ( .A(n2688), .Z(n2703) );
  XNOR U3749 ( .A(n2703), .B(x[40]), .Z(n2704) );
  XNOR U3750 ( .A(n2723), .B(n2704), .Z(n2716) );
  NAND U3751 ( .A(n2754), .B(n2716), .Z(n2665) );
  XNOR U3752 ( .A(n2671), .B(n2665), .Z(n2684) );
  XOR U3753 ( .A(x[41]), .B(x[47]), .Z(n2722) );
  XOR U3754 ( .A(n2666), .B(n2723), .Z(n2712) );
  ANDN U3755 ( .B(n2722), .A(n2712), .Z(n2673) );
  XOR U3756 ( .A(x[47]), .B(n2723), .Z(n2765) );
  IV U3757 ( .A(n2765), .Z(n2676) );
  NAND U3758 ( .A(n2666), .B(n2676), .Z(n2667) );
  XOR U3759 ( .A(n2673), .B(n2667), .Z(n2668) );
  XNOR U3760 ( .A(n2684), .B(n2668), .Z(n2708) );
  NANDN U3761 ( .A(x[41]), .B(n2677), .Z(n2675) );
  XNOR U3762 ( .A(n2703), .B(n2712), .Z(n2747) );
  XOR U3763 ( .A(x[44]), .B(x[42]), .Z(n2730) );
  AND U3764 ( .A(n2747), .B(n2730), .Z(n2670) );
  XNOR U3765 ( .A(n2732), .B(n2765), .Z(n2669) );
  XNOR U3766 ( .A(n2670), .B(n2669), .Z(n2672) );
  XOR U3767 ( .A(n2672), .B(n2671), .Z(n2692) );
  XNOR U3768 ( .A(n2673), .B(n2692), .Z(n2674) );
  XNOR U3769 ( .A(n2675), .B(n2674), .Z(n2706) );
  IV U3770 ( .A(n2706), .Z(n2709) );
  NAND U3771 ( .A(n2708), .B(n2709), .Z(n2702) );
  NANDN U3772 ( .A(n2708), .B(n2709), .Z(n2696) );
  XNOR U3773 ( .A(x[42]), .B(n2676), .Z(n2683) );
  XNOR U3774 ( .A(x[41]), .B(n2683), .Z(n2687) );
  IV U3775 ( .A(n2687), .Z(n2741) );
  XNOR U3776 ( .A(x[44]), .B(n2677), .Z(n2753) );
  OR U3777 ( .A(x[40]), .B(n2753), .Z(n2678) );
  XNOR U3778 ( .A(n2741), .B(n2678), .Z(n2679) );
  NANDN U3779 ( .A(n2688), .B(n2679), .Z(n2682) );
  ANDN U3780 ( .B(x[40]), .A(n2753), .Z(n2680) );
  NAND U3781 ( .A(n2688), .B(n2680), .Z(n2681) );
  NAND U3782 ( .A(n2682), .B(n2681), .Z(n2686) );
  XNOR U3783 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3784 ( .A(n2686), .B(n2685), .Z(n2710) );
  IV U3785 ( .A(n2708), .Z(n2707) );
  ANDN U3786 ( .B(n2710), .A(n2707), .Z(n2693) );
  AND U3787 ( .A(x[40]), .B(n2687), .Z(n2690) );
  NAND U3788 ( .A(n2688), .B(n2753), .Z(n2689) );
  XNOR U3789 ( .A(n2690), .B(n2689), .Z(n2691) );
  XNOR U3790 ( .A(n2692), .B(n2691), .Z(n2711) );
  XNOR U3791 ( .A(n2693), .B(n2711), .Z(n2694) );
  NAND U3792 ( .A(n2706), .B(n2694), .Z(n2695) );
  NAND U3793 ( .A(n2696), .B(n2695), .Z(n2740) );
  IV U3794 ( .A(n2740), .Z(n2715) );
  OR U3795 ( .A(n2710), .B(n2706), .Z(n2697) );
  NAND U3796 ( .A(n2707), .B(n2697), .Z(n2700) );
  XOR U3797 ( .A(n2710), .B(n2711), .Z(n2698) );
  NANDN U3798 ( .A(n2709), .B(n2698), .Z(n2699) );
  NAND U3799 ( .A(n2700), .B(n2699), .Z(n2752) );
  NANDN U3800 ( .A(n2715), .B(n2752), .Z(n2701) );
  AND U3801 ( .A(n2702), .B(n2701), .Z(n2743) );
  AND U3802 ( .A(n2743), .B(n2703), .Z(n2718) );
  OR U3803 ( .A(n2704), .B(n2715), .Z(n2705) );
  XNOR U3804 ( .A(n2718), .B(n2705), .Z(n2751) );
  XOR U3805 ( .A(n2766), .B(n2725), .Z(n2721) );
  ANDN U3806 ( .B(n2721), .A(n2712), .Z(n2733) );
  NAND U3807 ( .A(n2723), .B(n2725), .Z(n2713) );
  XNOR U3808 ( .A(n2733), .B(n2713), .Z(n2758) );
  XNOR U3809 ( .A(n2751), .B(n2758), .Z(z[42]) );
  AND U3810 ( .A(x[40]), .B(n2752), .Z(n2720) );
  AND U3811 ( .A(n2714), .B(n2729), .Z(n2750) );
  XOR U3812 ( .A(n2715), .B(n2725), .Z(n2728) );
  IV U3813 ( .A(n2728), .Z(n2755) );
  NAND U3814 ( .A(n2755), .B(n2716), .Z(n2717) );
  XNOR U3815 ( .A(n2750), .B(n2717), .Z(n2734) );
  XNOR U3816 ( .A(n2718), .B(n2734), .Z(n2719) );
  XNOR U3817 ( .A(n2720), .B(n2719), .Z(n3941) );
  AND U3818 ( .A(n2722), .B(n2721), .Z(n2767) );
  XOR U3819 ( .A(x[41]), .B(n2723), .Z(n2724) );
  NAND U3820 ( .A(n2725), .B(n2724), .Z(n2726) );
  XNOR U3821 ( .A(n2767), .B(n2726), .Z(n2738) );
  AND U3822 ( .A(n2729), .B(n2727), .Z(n2757) );
  XNOR U3823 ( .A(n2729), .B(n2728), .Z(n2748) );
  NAND U3824 ( .A(n2748), .B(n2730), .Z(n2731) );
  XNOR U3825 ( .A(n2757), .B(n2731), .Z(n2744) );
  AND U3826 ( .A(n2766), .B(n2732), .Z(n2736) );
  XNOR U3827 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U3828 ( .A(n2736), .B(n2735), .Z(n3940) );
  XNOR U3829 ( .A(n2744), .B(n3940), .Z(n2737) );
  XNOR U3830 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U3831 ( .A(n3941), .B(n2739), .Z(z[45]) );
  AND U3832 ( .A(n2741), .B(n2740), .Z(n2746) );
  XOR U3833 ( .A(n2741), .B(n2753), .Z(n2742) );
  AND U3834 ( .A(n2743), .B(n2742), .Z(n2762) );
  XNOR U3835 ( .A(n2744), .B(n2762), .Z(n2745) );
  XNOR U3836 ( .A(n2746), .B(n2745), .Z(n2773) );
  NAND U3837 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3838 ( .A(n2750), .B(n2749), .Z(n2761) );
  XNOR U3839 ( .A(n2751), .B(n2761), .Z(n3939) );
  XNOR U3840 ( .A(n2773), .B(n3939), .Z(n2771) );
  AND U3841 ( .A(n2753), .B(n2752), .Z(n2760) );
  NAND U3842 ( .A(n2755), .B(n2754), .Z(n2756) );
  XNOR U3843 ( .A(n2757), .B(n2756), .Z(n2768) );
  XNOR U3844 ( .A(n2768), .B(n2758), .Z(n2759) );
  XNOR U3845 ( .A(n2760), .B(n2759), .Z(n2764) );
  XNOR U3846 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U3847 ( .A(n2764), .B(n2763), .Z(n2772) );
  XNOR U3848 ( .A(n2771), .B(n2772), .Z(z[41]) );
  AND U3849 ( .A(n2766), .B(n2765), .Z(n2770) );
  XNOR U3850 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U3851 ( .A(n2770), .B(n2769), .Z(n2775) );
  XNOR U3852 ( .A(n2771), .B(n2775), .Z(z[46]) );
  XOR U3853 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U3854 ( .A(n2775), .B(n2774), .Z(z[43]) );
  XOR U3855 ( .A(x[49]), .B(x[51]), .Z(n2779) );
  XOR U3856 ( .A(x[48]), .B(x[54]), .Z(n2777) );
  XNOR U3857 ( .A(n2779), .B(n2777), .Z(n2776) );
  XNOR U3858 ( .A(x[50]), .B(n2776), .Z(n2847) );
  IV U3859 ( .A(n2847), .Z(n2781) );
  XNOR U3860 ( .A(x[48]), .B(n2781), .Z(n2829) );
  XNOR U3861 ( .A(x[52]), .B(x[55]), .Z(n2778) );
  IV U3862 ( .A(n2778), .Z(n2842) );
  AND U3863 ( .A(n2829), .B(n2842), .Z(n2786) );
  XOR U3864 ( .A(x[55]), .B(x[50]), .Z(n2869) );
  XNOR U3865 ( .A(n2777), .B(x[53]), .Z(n2792) );
  IV U3866 ( .A(n2792), .Z(n2838) );
  XOR U3867 ( .A(n2779), .B(n2778), .Z(n2803) );
  IV U3868 ( .A(n2803), .Z(n2818) );
  XNOR U3869 ( .A(n2818), .B(x[48]), .Z(n2819) );
  XNOR U3870 ( .A(n2838), .B(n2819), .Z(n2831) );
  NAND U3871 ( .A(n2869), .B(n2831), .Z(n2780) );
  XNOR U3872 ( .A(n2786), .B(n2780), .Z(n2799) );
  XOR U3873 ( .A(x[49]), .B(x[55]), .Z(n2837) );
  XOR U3874 ( .A(n2781), .B(n2838), .Z(n2827) );
  ANDN U3875 ( .B(n2837), .A(n2827), .Z(n2788) );
  XOR U3876 ( .A(x[55]), .B(n2838), .Z(n2880) );
  IV U3877 ( .A(n2880), .Z(n2791) );
  NAND U3878 ( .A(n2781), .B(n2791), .Z(n2782) );
  XOR U3879 ( .A(n2788), .B(n2782), .Z(n2783) );
  XNOR U3880 ( .A(n2799), .B(n2783), .Z(n2823) );
  NANDN U3881 ( .A(x[49]), .B(n2792), .Z(n2790) );
  XNOR U3882 ( .A(n2818), .B(n2827), .Z(n2862) );
  XOR U3883 ( .A(x[52]), .B(x[50]), .Z(n2845) );
  AND U3884 ( .A(n2862), .B(n2845), .Z(n2785) );
  XNOR U3885 ( .A(n2847), .B(n2880), .Z(n2784) );
  XNOR U3886 ( .A(n2785), .B(n2784), .Z(n2787) );
  XOR U3887 ( .A(n2787), .B(n2786), .Z(n2807) );
  XNOR U3888 ( .A(n2788), .B(n2807), .Z(n2789) );
  XNOR U3889 ( .A(n2790), .B(n2789), .Z(n2821) );
  IV U3890 ( .A(n2821), .Z(n2824) );
  NAND U3891 ( .A(n2823), .B(n2824), .Z(n2817) );
  NANDN U3892 ( .A(n2823), .B(n2824), .Z(n2811) );
  XNOR U3893 ( .A(x[50]), .B(n2791), .Z(n2798) );
  XNOR U3894 ( .A(x[49]), .B(n2798), .Z(n2802) );
  IV U3895 ( .A(n2802), .Z(n2856) );
  XNOR U3896 ( .A(x[52]), .B(n2792), .Z(n2868) );
  OR U3897 ( .A(x[48]), .B(n2868), .Z(n2793) );
  XNOR U3898 ( .A(n2856), .B(n2793), .Z(n2794) );
  NANDN U3899 ( .A(n2803), .B(n2794), .Z(n2797) );
  ANDN U3900 ( .B(x[48]), .A(n2868), .Z(n2795) );
  NAND U3901 ( .A(n2803), .B(n2795), .Z(n2796) );
  NAND U3902 ( .A(n2797), .B(n2796), .Z(n2801) );
  XNOR U3903 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3904 ( .A(n2801), .B(n2800), .Z(n2825) );
  IV U3905 ( .A(n2823), .Z(n2822) );
  ANDN U3906 ( .B(n2825), .A(n2822), .Z(n2808) );
  AND U3907 ( .A(x[48]), .B(n2802), .Z(n2805) );
  NAND U3908 ( .A(n2803), .B(n2868), .Z(n2804) );
  XNOR U3909 ( .A(n2805), .B(n2804), .Z(n2806) );
  XNOR U3910 ( .A(n2807), .B(n2806), .Z(n2826) );
  XNOR U3911 ( .A(n2808), .B(n2826), .Z(n2809) );
  NAND U3912 ( .A(n2821), .B(n2809), .Z(n2810) );
  NAND U3913 ( .A(n2811), .B(n2810), .Z(n2855) );
  IV U3914 ( .A(n2855), .Z(n2830) );
  OR U3915 ( .A(n2825), .B(n2821), .Z(n2812) );
  NAND U3916 ( .A(n2822), .B(n2812), .Z(n2815) );
  XOR U3917 ( .A(n2825), .B(n2826), .Z(n2813) );
  NANDN U3918 ( .A(n2824), .B(n2813), .Z(n2814) );
  NAND U3919 ( .A(n2815), .B(n2814), .Z(n2867) );
  NANDN U3920 ( .A(n2830), .B(n2867), .Z(n2816) );
  AND U3921 ( .A(n2817), .B(n2816), .Z(n2858) );
  AND U3922 ( .A(n2858), .B(n2818), .Z(n2833) );
  OR U3923 ( .A(n2819), .B(n2830), .Z(n2820) );
  XNOR U3924 ( .A(n2833), .B(n2820), .Z(n2866) );
  XOR U3925 ( .A(n2881), .B(n2840), .Z(n2836) );
  ANDN U3926 ( .B(n2836), .A(n2827), .Z(n2848) );
  NAND U3927 ( .A(n2838), .B(n2840), .Z(n2828) );
  XNOR U3928 ( .A(n2848), .B(n2828), .Z(n2873) );
  XNOR U3929 ( .A(n2866), .B(n2873), .Z(z[50]) );
  AND U3930 ( .A(x[48]), .B(n2867), .Z(n2835) );
  AND U3931 ( .A(n2829), .B(n2844), .Z(n2865) );
  XOR U3932 ( .A(n2830), .B(n2840), .Z(n2843) );
  IV U3933 ( .A(n2843), .Z(n2870) );
  NAND U3934 ( .A(n2870), .B(n2831), .Z(n2832) );
  XNOR U3935 ( .A(n2865), .B(n2832), .Z(n2849) );
  XNOR U3936 ( .A(n2833), .B(n2849), .Z(n2834) );
  XNOR U3937 ( .A(n2835), .B(n2834), .Z(n3945) );
  AND U3938 ( .A(n2837), .B(n2836), .Z(n2882) );
  XOR U3939 ( .A(x[49]), .B(n2838), .Z(n2839) );
  NAND U3940 ( .A(n2840), .B(n2839), .Z(n2841) );
  XNOR U3941 ( .A(n2882), .B(n2841), .Z(n2853) );
  AND U3942 ( .A(n2844), .B(n2842), .Z(n2872) );
  XNOR U3943 ( .A(n2844), .B(n2843), .Z(n2863) );
  NAND U3944 ( .A(n2863), .B(n2845), .Z(n2846) );
  XNOR U3945 ( .A(n2872), .B(n2846), .Z(n2859) );
  AND U3946 ( .A(n2881), .B(n2847), .Z(n2851) );
  XNOR U3947 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U3948 ( .A(n2851), .B(n2850), .Z(n3944) );
  XNOR U3949 ( .A(n2859), .B(n3944), .Z(n2852) );
  XNOR U3950 ( .A(n2853), .B(n2852), .Z(n2854) );
  XNOR U3951 ( .A(n3945), .B(n2854), .Z(z[53]) );
  AND U3952 ( .A(n2856), .B(n2855), .Z(n2861) );
  XOR U3953 ( .A(n2856), .B(n2868), .Z(n2857) );
  AND U3954 ( .A(n2858), .B(n2857), .Z(n2877) );
  XNOR U3955 ( .A(n2859), .B(n2877), .Z(n2860) );
  XNOR U3956 ( .A(n2861), .B(n2860), .Z(n2888) );
  NAND U3957 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3958 ( .A(n2865), .B(n2864), .Z(n2876) );
  XNOR U3959 ( .A(n2866), .B(n2876), .Z(n3942) );
  XNOR U3960 ( .A(n2888), .B(n3942), .Z(n2886) );
  AND U3961 ( .A(n2868), .B(n2867), .Z(n2875) );
  NAND U3962 ( .A(n2870), .B(n2869), .Z(n2871) );
  XNOR U3963 ( .A(n2872), .B(n2871), .Z(n2883) );
  XNOR U3964 ( .A(n2883), .B(n2873), .Z(n2874) );
  XNOR U3965 ( .A(n2875), .B(n2874), .Z(n2879) );
  XNOR U3966 ( .A(n2877), .B(n2876), .Z(n2878) );
  XNOR U3967 ( .A(n2879), .B(n2878), .Z(n2887) );
  XNOR U3968 ( .A(n2886), .B(n2887), .Z(z[49]) );
  AND U3969 ( .A(n2881), .B(n2880), .Z(n2885) );
  XNOR U3970 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U3971 ( .A(n2885), .B(n2884), .Z(n2890) );
  XNOR U3972 ( .A(n2886), .B(n2890), .Z(z[54]) );
  XOR U3973 ( .A(n2888), .B(n2887), .Z(n2889) );
  XNOR U3974 ( .A(n2890), .B(n2889), .Z(z[51]) );
  XOR U3975 ( .A(x[57]), .B(x[59]), .Z(n2894) );
  XOR U3976 ( .A(x[56]), .B(x[62]), .Z(n2892) );
  XNOR U3977 ( .A(n2894), .B(n2892), .Z(n2891) );
  XNOR U3978 ( .A(x[58]), .B(n2891), .Z(n2962) );
  IV U3979 ( .A(n2962), .Z(n2896) );
  XNOR U3980 ( .A(x[56]), .B(n2896), .Z(n2944) );
  XNOR U3981 ( .A(x[60]), .B(x[63]), .Z(n2893) );
  IV U3982 ( .A(n2893), .Z(n2957) );
  AND U3983 ( .A(n2944), .B(n2957), .Z(n2901) );
  XOR U3984 ( .A(x[63]), .B(x[58]), .Z(n2984) );
  XNOR U3985 ( .A(n2892), .B(x[61]), .Z(n2907) );
  IV U3986 ( .A(n2907), .Z(n2953) );
  XOR U3987 ( .A(n2894), .B(n2893), .Z(n2918) );
  IV U3988 ( .A(n2918), .Z(n2933) );
  XNOR U3989 ( .A(n2933), .B(x[56]), .Z(n2934) );
  XNOR U3990 ( .A(n2953), .B(n2934), .Z(n2946) );
  NAND U3991 ( .A(n2984), .B(n2946), .Z(n2895) );
  XNOR U3992 ( .A(n2901), .B(n2895), .Z(n2914) );
  XOR U3993 ( .A(x[57]), .B(x[63]), .Z(n2952) );
  XOR U3994 ( .A(n2896), .B(n2953), .Z(n2942) );
  ANDN U3995 ( .B(n2952), .A(n2942), .Z(n2903) );
  XOR U3996 ( .A(x[63]), .B(n2953), .Z(n2995) );
  IV U3997 ( .A(n2995), .Z(n2906) );
  NAND U3998 ( .A(n2896), .B(n2906), .Z(n2897) );
  XOR U3999 ( .A(n2903), .B(n2897), .Z(n2898) );
  XNOR U4000 ( .A(n2914), .B(n2898), .Z(n2938) );
  NANDN U4001 ( .A(x[57]), .B(n2907), .Z(n2905) );
  XNOR U4002 ( .A(n2933), .B(n2942), .Z(n2977) );
  XOR U4003 ( .A(x[60]), .B(x[58]), .Z(n2960) );
  AND U4004 ( .A(n2977), .B(n2960), .Z(n2900) );
  XNOR U4005 ( .A(n2962), .B(n2995), .Z(n2899) );
  XNOR U4006 ( .A(n2900), .B(n2899), .Z(n2902) );
  XOR U4007 ( .A(n2902), .B(n2901), .Z(n2922) );
  XNOR U4008 ( .A(n2903), .B(n2922), .Z(n2904) );
  XNOR U4009 ( .A(n2905), .B(n2904), .Z(n2936) );
  IV U4010 ( .A(n2936), .Z(n2939) );
  NAND U4011 ( .A(n2938), .B(n2939), .Z(n2932) );
  NANDN U4012 ( .A(n2938), .B(n2939), .Z(n2926) );
  XNOR U4013 ( .A(x[58]), .B(n2906), .Z(n2913) );
  XNOR U4014 ( .A(x[57]), .B(n2913), .Z(n2917) );
  IV U4015 ( .A(n2917), .Z(n2971) );
  XNOR U4016 ( .A(x[60]), .B(n2907), .Z(n2983) );
  OR U4017 ( .A(x[56]), .B(n2983), .Z(n2908) );
  XNOR U4018 ( .A(n2971), .B(n2908), .Z(n2909) );
  NANDN U4019 ( .A(n2918), .B(n2909), .Z(n2912) );
  ANDN U4020 ( .B(x[56]), .A(n2983), .Z(n2910) );
  NAND U4021 ( .A(n2918), .B(n2910), .Z(n2911) );
  NAND U4022 ( .A(n2912), .B(n2911), .Z(n2916) );
  XNOR U4023 ( .A(n2914), .B(n2913), .Z(n2915) );
  XOR U4024 ( .A(n2916), .B(n2915), .Z(n2940) );
  IV U4025 ( .A(n2938), .Z(n2937) );
  ANDN U4026 ( .B(n2940), .A(n2937), .Z(n2923) );
  AND U4027 ( .A(x[56]), .B(n2917), .Z(n2920) );
  NAND U4028 ( .A(n2918), .B(n2983), .Z(n2919) );
  XNOR U4029 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4030 ( .A(n2922), .B(n2921), .Z(n2941) );
  XNOR U4031 ( .A(n2923), .B(n2941), .Z(n2924) );
  NAND U4032 ( .A(n2936), .B(n2924), .Z(n2925) );
  NAND U4033 ( .A(n2926), .B(n2925), .Z(n2970) );
  IV U4034 ( .A(n2970), .Z(n2945) );
  OR U4035 ( .A(n2940), .B(n2936), .Z(n2927) );
  NAND U4036 ( .A(n2937), .B(n2927), .Z(n2930) );
  XOR U4037 ( .A(n2940), .B(n2941), .Z(n2928) );
  NANDN U4038 ( .A(n2939), .B(n2928), .Z(n2929) );
  NAND U4039 ( .A(n2930), .B(n2929), .Z(n2982) );
  NANDN U4040 ( .A(n2945), .B(n2982), .Z(n2931) );
  AND U4041 ( .A(n2932), .B(n2931), .Z(n2973) );
  AND U4042 ( .A(n2973), .B(n2933), .Z(n2948) );
  OR U4043 ( .A(n2934), .B(n2945), .Z(n2935) );
  XNOR U4044 ( .A(n2948), .B(n2935), .Z(n2981) );
  XOR U4045 ( .A(n2996), .B(n2955), .Z(n2951) );
  ANDN U4046 ( .B(n2951), .A(n2942), .Z(n2963) );
  NAND U4047 ( .A(n2953), .B(n2955), .Z(n2943) );
  XNOR U4048 ( .A(n2963), .B(n2943), .Z(n2988) );
  XNOR U4049 ( .A(n2981), .B(n2988), .Z(z[58]) );
  AND U4050 ( .A(x[56]), .B(n2982), .Z(n2950) );
  AND U4051 ( .A(n2944), .B(n2959), .Z(n2980) );
  XOR U4052 ( .A(n2945), .B(n2955), .Z(n2958) );
  IV U4053 ( .A(n2958), .Z(n2985) );
  NAND U4054 ( .A(n2985), .B(n2946), .Z(n2947) );
  XNOR U4055 ( .A(n2980), .B(n2947), .Z(n2964) );
  XNOR U4056 ( .A(n2948), .B(n2964), .Z(n2949) );
  XNOR U4057 ( .A(n2950), .B(n2949), .Z(n3948) );
  AND U4058 ( .A(n2952), .B(n2951), .Z(n2997) );
  XOR U4059 ( .A(x[57]), .B(n2953), .Z(n2954) );
  NAND U4060 ( .A(n2955), .B(n2954), .Z(n2956) );
  XNOR U4061 ( .A(n2997), .B(n2956), .Z(n2968) );
  AND U4062 ( .A(n2959), .B(n2957), .Z(n2987) );
  XNOR U4063 ( .A(n2959), .B(n2958), .Z(n2978) );
  NAND U4064 ( .A(n2978), .B(n2960), .Z(n2961) );
  XNOR U4065 ( .A(n2987), .B(n2961), .Z(n2974) );
  AND U4066 ( .A(n2996), .B(n2962), .Z(n2966) );
  XNOR U4067 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U4068 ( .A(n2966), .B(n2965), .Z(n3947) );
  XNOR U4069 ( .A(n2974), .B(n3947), .Z(n2967) );
  XNOR U4070 ( .A(n2968), .B(n2967), .Z(n2969) );
  XNOR U4071 ( .A(n3948), .B(n2969), .Z(z[61]) );
  AND U4072 ( .A(n2971), .B(n2970), .Z(n2976) );
  XOR U4073 ( .A(n2971), .B(n2983), .Z(n2972) );
  AND U4074 ( .A(n2973), .B(n2972), .Z(n2992) );
  XNOR U4075 ( .A(n2974), .B(n2992), .Z(n2975) );
  XNOR U4076 ( .A(n2976), .B(n2975), .Z(n3003) );
  NAND U4077 ( .A(n2978), .B(n2977), .Z(n2979) );
  XNOR U4078 ( .A(n2980), .B(n2979), .Z(n2991) );
  XNOR U4079 ( .A(n2981), .B(n2991), .Z(n3946) );
  XNOR U4080 ( .A(n3003), .B(n3946), .Z(n3001) );
  AND U4081 ( .A(n2983), .B(n2982), .Z(n2990) );
  NAND U4082 ( .A(n2985), .B(n2984), .Z(n2986) );
  XNOR U4083 ( .A(n2987), .B(n2986), .Z(n2998) );
  XNOR U4084 ( .A(n2998), .B(n2988), .Z(n2989) );
  XNOR U4085 ( .A(n2990), .B(n2989), .Z(n2994) );
  XNOR U4086 ( .A(n2992), .B(n2991), .Z(n2993) );
  XNOR U4087 ( .A(n2994), .B(n2993), .Z(n3002) );
  XNOR U4088 ( .A(n3001), .B(n3002), .Z(z[57]) );
  AND U4089 ( .A(n2996), .B(n2995), .Z(n3000) );
  XNOR U4090 ( .A(n2998), .B(n2997), .Z(n2999) );
  XNOR U4091 ( .A(n3000), .B(n2999), .Z(n3005) );
  XNOR U4092 ( .A(n3001), .B(n3005), .Z(z[62]) );
  XOR U4093 ( .A(n3003), .B(n3002), .Z(n3004) );
  XNOR U4094 ( .A(n3005), .B(n3004), .Z(z[59]) );
  XOR U4095 ( .A(x[65]), .B(x[67]), .Z(n3009) );
  XOR U4096 ( .A(x[64]), .B(x[70]), .Z(n3007) );
  XNOR U4097 ( .A(n3009), .B(n3007), .Z(n3006) );
  XNOR U4098 ( .A(x[66]), .B(n3006), .Z(n3077) );
  IV U4099 ( .A(n3077), .Z(n3011) );
  XNOR U4100 ( .A(x[64]), .B(n3011), .Z(n3059) );
  XNOR U4101 ( .A(x[68]), .B(x[71]), .Z(n3008) );
  IV U4102 ( .A(n3008), .Z(n3072) );
  AND U4103 ( .A(n3059), .B(n3072), .Z(n3016) );
  XOR U4104 ( .A(x[71]), .B(x[66]), .Z(n3099) );
  XNOR U4105 ( .A(n3007), .B(x[69]), .Z(n3022) );
  IV U4106 ( .A(n3022), .Z(n3068) );
  XOR U4107 ( .A(n3009), .B(n3008), .Z(n3033) );
  IV U4108 ( .A(n3033), .Z(n3048) );
  XNOR U4109 ( .A(n3048), .B(x[64]), .Z(n3049) );
  XNOR U4110 ( .A(n3068), .B(n3049), .Z(n3061) );
  NAND U4111 ( .A(n3099), .B(n3061), .Z(n3010) );
  XNOR U4112 ( .A(n3016), .B(n3010), .Z(n3029) );
  XOR U4113 ( .A(x[65]), .B(x[71]), .Z(n3067) );
  XOR U4114 ( .A(n3011), .B(n3068), .Z(n3057) );
  ANDN U4115 ( .B(n3067), .A(n3057), .Z(n3018) );
  XOR U4116 ( .A(x[71]), .B(n3068), .Z(n3110) );
  IV U4117 ( .A(n3110), .Z(n3021) );
  NAND U4118 ( .A(n3011), .B(n3021), .Z(n3012) );
  XOR U4119 ( .A(n3018), .B(n3012), .Z(n3013) );
  XNOR U4120 ( .A(n3029), .B(n3013), .Z(n3053) );
  NANDN U4121 ( .A(x[65]), .B(n3022), .Z(n3020) );
  XNOR U4122 ( .A(n3048), .B(n3057), .Z(n3092) );
  XOR U4123 ( .A(x[68]), .B(x[66]), .Z(n3075) );
  AND U4124 ( .A(n3092), .B(n3075), .Z(n3015) );
  XNOR U4125 ( .A(n3077), .B(n3110), .Z(n3014) );
  XNOR U4126 ( .A(n3015), .B(n3014), .Z(n3017) );
  XOR U4127 ( .A(n3017), .B(n3016), .Z(n3037) );
  XNOR U4128 ( .A(n3018), .B(n3037), .Z(n3019) );
  XNOR U4129 ( .A(n3020), .B(n3019), .Z(n3051) );
  IV U4130 ( .A(n3051), .Z(n3054) );
  NAND U4131 ( .A(n3053), .B(n3054), .Z(n3047) );
  NANDN U4132 ( .A(n3053), .B(n3054), .Z(n3041) );
  XNOR U4133 ( .A(x[66]), .B(n3021), .Z(n3028) );
  XNOR U4134 ( .A(x[65]), .B(n3028), .Z(n3032) );
  IV U4135 ( .A(n3032), .Z(n3086) );
  XNOR U4136 ( .A(x[68]), .B(n3022), .Z(n3098) );
  OR U4137 ( .A(x[64]), .B(n3098), .Z(n3023) );
  XNOR U4138 ( .A(n3086), .B(n3023), .Z(n3024) );
  NANDN U4139 ( .A(n3033), .B(n3024), .Z(n3027) );
  ANDN U4140 ( .B(x[64]), .A(n3098), .Z(n3025) );
  NAND U4141 ( .A(n3033), .B(n3025), .Z(n3026) );
  NAND U4142 ( .A(n3027), .B(n3026), .Z(n3031) );
  XNOR U4143 ( .A(n3029), .B(n3028), .Z(n3030) );
  XOR U4144 ( .A(n3031), .B(n3030), .Z(n3055) );
  IV U4145 ( .A(n3053), .Z(n3052) );
  ANDN U4146 ( .B(n3055), .A(n3052), .Z(n3038) );
  AND U4147 ( .A(x[64]), .B(n3032), .Z(n3035) );
  NAND U4148 ( .A(n3033), .B(n3098), .Z(n3034) );
  XNOR U4149 ( .A(n3035), .B(n3034), .Z(n3036) );
  XNOR U4150 ( .A(n3037), .B(n3036), .Z(n3056) );
  XNOR U4151 ( .A(n3038), .B(n3056), .Z(n3039) );
  NAND U4152 ( .A(n3051), .B(n3039), .Z(n3040) );
  NAND U4153 ( .A(n3041), .B(n3040), .Z(n3085) );
  IV U4154 ( .A(n3085), .Z(n3060) );
  OR U4155 ( .A(n3055), .B(n3051), .Z(n3042) );
  NAND U4156 ( .A(n3052), .B(n3042), .Z(n3045) );
  XOR U4157 ( .A(n3055), .B(n3056), .Z(n3043) );
  NANDN U4158 ( .A(n3054), .B(n3043), .Z(n3044) );
  NAND U4159 ( .A(n3045), .B(n3044), .Z(n3097) );
  NANDN U4160 ( .A(n3060), .B(n3097), .Z(n3046) );
  AND U4161 ( .A(n3047), .B(n3046), .Z(n3088) );
  AND U4162 ( .A(n3088), .B(n3048), .Z(n3063) );
  OR U4163 ( .A(n3049), .B(n3060), .Z(n3050) );
  XNOR U4164 ( .A(n3063), .B(n3050), .Z(n3096) );
  XOR U4165 ( .A(n3111), .B(n3070), .Z(n3066) );
  ANDN U4166 ( .B(n3066), .A(n3057), .Z(n3078) );
  NAND U4167 ( .A(n3068), .B(n3070), .Z(n3058) );
  XNOR U4168 ( .A(n3078), .B(n3058), .Z(n3103) );
  XNOR U4169 ( .A(n3096), .B(n3103), .Z(z[66]) );
  AND U4170 ( .A(x[64]), .B(n3097), .Z(n3065) );
  AND U4171 ( .A(n3059), .B(n3074), .Z(n3095) );
  XOR U4172 ( .A(n3060), .B(n3070), .Z(n3073) );
  IV U4173 ( .A(n3073), .Z(n3100) );
  NAND U4174 ( .A(n3100), .B(n3061), .Z(n3062) );
  XNOR U4175 ( .A(n3095), .B(n3062), .Z(n3079) );
  XNOR U4176 ( .A(n3063), .B(n3079), .Z(n3064) );
  XNOR U4177 ( .A(n3065), .B(n3064), .Z(n3951) );
  AND U4178 ( .A(n3067), .B(n3066), .Z(n3112) );
  XOR U4179 ( .A(x[65]), .B(n3068), .Z(n3069) );
  NAND U4180 ( .A(n3070), .B(n3069), .Z(n3071) );
  XNOR U4181 ( .A(n3112), .B(n3071), .Z(n3083) );
  AND U4182 ( .A(n3074), .B(n3072), .Z(n3102) );
  XNOR U4183 ( .A(n3074), .B(n3073), .Z(n3093) );
  NAND U4184 ( .A(n3093), .B(n3075), .Z(n3076) );
  XNOR U4185 ( .A(n3102), .B(n3076), .Z(n3089) );
  AND U4186 ( .A(n3111), .B(n3077), .Z(n3081) );
  XNOR U4187 ( .A(n3079), .B(n3078), .Z(n3080) );
  XNOR U4188 ( .A(n3081), .B(n3080), .Z(n3950) );
  XNOR U4189 ( .A(n3089), .B(n3950), .Z(n3082) );
  XNOR U4190 ( .A(n3083), .B(n3082), .Z(n3084) );
  XNOR U4191 ( .A(n3951), .B(n3084), .Z(z[69]) );
  AND U4192 ( .A(n3086), .B(n3085), .Z(n3091) );
  XOR U4193 ( .A(n3086), .B(n3098), .Z(n3087) );
  AND U4194 ( .A(n3088), .B(n3087), .Z(n3107) );
  XNOR U4195 ( .A(n3089), .B(n3107), .Z(n3090) );
  XNOR U4196 ( .A(n3091), .B(n3090), .Z(n3118) );
  NAND U4197 ( .A(n3093), .B(n3092), .Z(n3094) );
  XNOR U4198 ( .A(n3095), .B(n3094), .Z(n3106) );
  XNOR U4199 ( .A(n3096), .B(n3106), .Z(n3949) );
  XNOR U4200 ( .A(n3118), .B(n3949), .Z(n3116) );
  AND U4201 ( .A(n3098), .B(n3097), .Z(n3105) );
  NAND U4202 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U4203 ( .A(n3102), .B(n3101), .Z(n3113) );
  XNOR U4204 ( .A(n3113), .B(n3103), .Z(n3104) );
  XNOR U4205 ( .A(n3105), .B(n3104), .Z(n3109) );
  XNOR U4206 ( .A(n3107), .B(n3106), .Z(n3108) );
  XNOR U4207 ( .A(n3109), .B(n3108), .Z(n3117) );
  XNOR U4208 ( .A(n3116), .B(n3117), .Z(z[65]) );
  AND U4209 ( .A(n3111), .B(n3110), .Z(n3115) );
  XNOR U4210 ( .A(n3113), .B(n3112), .Z(n3114) );
  XNOR U4211 ( .A(n3115), .B(n3114), .Z(n3120) );
  XNOR U4212 ( .A(n3116), .B(n3120), .Z(z[70]) );
  XOR U4213 ( .A(n3118), .B(n3117), .Z(n3119) );
  XNOR U4214 ( .A(n3120), .B(n3119), .Z(z[67]) );
  XOR U4215 ( .A(x[73]), .B(x[75]), .Z(n3124) );
  XOR U4216 ( .A(x[72]), .B(x[78]), .Z(n3122) );
  XNOR U4217 ( .A(n3124), .B(n3122), .Z(n3121) );
  XNOR U4218 ( .A(x[74]), .B(n3121), .Z(n3192) );
  IV U4219 ( .A(n3192), .Z(n3126) );
  XNOR U4220 ( .A(x[72]), .B(n3126), .Z(n3174) );
  XNOR U4221 ( .A(x[76]), .B(x[79]), .Z(n3123) );
  IV U4222 ( .A(n3123), .Z(n3187) );
  AND U4223 ( .A(n3174), .B(n3187), .Z(n3131) );
  XOR U4224 ( .A(x[79]), .B(x[74]), .Z(n3214) );
  XNOR U4225 ( .A(n3122), .B(x[77]), .Z(n3137) );
  IV U4226 ( .A(n3137), .Z(n3183) );
  XOR U4227 ( .A(n3124), .B(n3123), .Z(n3148) );
  IV U4228 ( .A(n3148), .Z(n3163) );
  XNOR U4229 ( .A(n3163), .B(x[72]), .Z(n3164) );
  XNOR U4230 ( .A(n3183), .B(n3164), .Z(n3176) );
  NAND U4231 ( .A(n3214), .B(n3176), .Z(n3125) );
  XNOR U4232 ( .A(n3131), .B(n3125), .Z(n3144) );
  XOR U4233 ( .A(x[73]), .B(x[79]), .Z(n3182) );
  XOR U4234 ( .A(n3126), .B(n3183), .Z(n3172) );
  ANDN U4235 ( .B(n3182), .A(n3172), .Z(n3133) );
  XOR U4236 ( .A(x[79]), .B(n3183), .Z(n3225) );
  IV U4237 ( .A(n3225), .Z(n3136) );
  NAND U4238 ( .A(n3126), .B(n3136), .Z(n3127) );
  XOR U4239 ( .A(n3133), .B(n3127), .Z(n3128) );
  XNOR U4240 ( .A(n3144), .B(n3128), .Z(n3168) );
  NANDN U4241 ( .A(x[73]), .B(n3137), .Z(n3135) );
  XNOR U4242 ( .A(n3163), .B(n3172), .Z(n3207) );
  XOR U4243 ( .A(x[76]), .B(x[74]), .Z(n3190) );
  AND U4244 ( .A(n3207), .B(n3190), .Z(n3130) );
  XNOR U4245 ( .A(n3192), .B(n3225), .Z(n3129) );
  XNOR U4246 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4247 ( .A(n3132), .B(n3131), .Z(n3152) );
  XNOR U4248 ( .A(n3133), .B(n3152), .Z(n3134) );
  XNOR U4249 ( .A(n3135), .B(n3134), .Z(n3166) );
  IV U4250 ( .A(n3166), .Z(n3169) );
  NAND U4251 ( .A(n3168), .B(n3169), .Z(n3162) );
  NANDN U4252 ( .A(n3168), .B(n3169), .Z(n3156) );
  XNOR U4253 ( .A(x[74]), .B(n3136), .Z(n3143) );
  XNOR U4254 ( .A(x[73]), .B(n3143), .Z(n3147) );
  IV U4255 ( .A(n3147), .Z(n3201) );
  XNOR U4256 ( .A(x[76]), .B(n3137), .Z(n3213) );
  OR U4257 ( .A(x[72]), .B(n3213), .Z(n3138) );
  XNOR U4258 ( .A(n3201), .B(n3138), .Z(n3139) );
  NANDN U4259 ( .A(n3148), .B(n3139), .Z(n3142) );
  ANDN U4260 ( .B(x[72]), .A(n3213), .Z(n3140) );
  NAND U4261 ( .A(n3148), .B(n3140), .Z(n3141) );
  NAND U4262 ( .A(n3142), .B(n3141), .Z(n3146) );
  XNOR U4263 ( .A(n3144), .B(n3143), .Z(n3145) );
  XOR U4264 ( .A(n3146), .B(n3145), .Z(n3170) );
  IV U4265 ( .A(n3168), .Z(n3167) );
  ANDN U4266 ( .B(n3170), .A(n3167), .Z(n3153) );
  AND U4267 ( .A(x[72]), .B(n3147), .Z(n3150) );
  NAND U4268 ( .A(n3148), .B(n3213), .Z(n3149) );
  XNOR U4269 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U4270 ( .A(n3152), .B(n3151), .Z(n3171) );
  XNOR U4271 ( .A(n3153), .B(n3171), .Z(n3154) );
  NAND U4272 ( .A(n3166), .B(n3154), .Z(n3155) );
  NAND U4273 ( .A(n3156), .B(n3155), .Z(n3200) );
  IV U4274 ( .A(n3200), .Z(n3175) );
  OR U4275 ( .A(n3170), .B(n3166), .Z(n3157) );
  NAND U4276 ( .A(n3167), .B(n3157), .Z(n3160) );
  XOR U4277 ( .A(n3170), .B(n3171), .Z(n3158) );
  NANDN U4278 ( .A(n3169), .B(n3158), .Z(n3159) );
  NAND U4279 ( .A(n3160), .B(n3159), .Z(n3212) );
  NANDN U4280 ( .A(n3175), .B(n3212), .Z(n3161) );
  AND U4281 ( .A(n3162), .B(n3161), .Z(n3203) );
  AND U4282 ( .A(n3203), .B(n3163), .Z(n3178) );
  OR U4283 ( .A(n3164), .B(n3175), .Z(n3165) );
  XNOR U4284 ( .A(n3178), .B(n3165), .Z(n3211) );
  XOR U4285 ( .A(n3226), .B(n3185), .Z(n3181) );
  ANDN U4286 ( .B(n3181), .A(n3172), .Z(n3193) );
  NAND U4287 ( .A(n3183), .B(n3185), .Z(n3173) );
  XNOR U4288 ( .A(n3193), .B(n3173), .Z(n3218) );
  XNOR U4289 ( .A(n3211), .B(n3218), .Z(z[74]) );
  AND U4290 ( .A(x[72]), .B(n3212), .Z(n3180) );
  AND U4291 ( .A(n3174), .B(n3189), .Z(n3210) );
  XOR U4292 ( .A(n3175), .B(n3185), .Z(n3188) );
  IV U4293 ( .A(n3188), .Z(n3215) );
  NAND U4294 ( .A(n3215), .B(n3176), .Z(n3177) );
  XNOR U4295 ( .A(n3210), .B(n3177), .Z(n3194) );
  XNOR U4296 ( .A(n3178), .B(n3194), .Z(n3179) );
  XNOR U4297 ( .A(n3180), .B(n3179), .Z(n3954) );
  AND U4298 ( .A(n3182), .B(n3181), .Z(n3227) );
  XOR U4299 ( .A(x[73]), .B(n3183), .Z(n3184) );
  NAND U4300 ( .A(n3185), .B(n3184), .Z(n3186) );
  XNOR U4301 ( .A(n3227), .B(n3186), .Z(n3198) );
  AND U4302 ( .A(n3189), .B(n3187), .Z(n3217) );
  XNOR U4303 ( .A(n3189), .B(n3188), .Z(n3208) );
  NAND U4304 ( .A(n3208), .B(n3190), .Z(n3191) );
  XNOR U4305 ( .A(n3217), .B(n3191), .Z(n3204) );
  AND U4306 ( .A(n3226), .B(n3192), .Z(n3196) );
  XNOR U4307 ( .A(n3194), .B(n3193), .Z(n3195) );
  XNOR U4308 ( .A(n3196), .B(n3195), .Z(n3953) );
  XNOR U4309 ( .A(n3204), .B(n3953), .Z(n3197) );
  XNOR U4310 ( .A(n3198), .B(n3197), .Z(n3199) );
  XNOR U4311 ( .A(n3954), .B(n3199), .Z(z[77]) );
  AND U4312 ( .A(n3201), .B(n3200), .Z(n3206) );
  XOR U4313 ( .A(n3201), .B(n3213), .Z(n3202) );
  AND U4314 ( .A(n3203), .B(n3202), .Z(n3222) );
  XNOR U4315 ( .A(n3204), .B(n3222), .Z(n3205) );
  XNOR U4316 ( .A(n3206), .B(n3205), .Z(n3233) );
  NAND U4317 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U4318 ( .A(n3210), .B(n3209), .Z(n3221) );
  XNOR U4319 ( .A(n3211), .B(n3221), .Z(n3952) );
  XNOR U4320 ( .A(n3233), .B(n3952), .Z(n3231) );
  AND U4321 ( .A(n3213), .B(n3212), .Z(n3220) );
  NAND U4322 ( .A(n3215), .B(n3214), .Z(n3216) );
  XNOR U4323 ( .A(n3217), .B(n3216), .Z(n3228) );
  XNOR U4324 ( .A(n3228), .B(n3218), .Z(n3219) );
  XNOR U4325 ( .A(n3220), .B(n3219), .Z(n3224) );
  XNOR U4326 ( .A(n3222), .B(n3221), .Z(n3223) );
  XNOR U4327 ( .A(n3224), .B(n3223), .Z(n3232) );
  XNOR U4328 ( .A(n3231), .B(n3232), .Z(z[73]) );
  AND U4329 ( .A(n3226), .B(n3225), .Z(n3230) );
  XNOR U4330 ( .A(n3228), .B(n3227), .Z(n3229) );
  XNOR U4331 ( .A(n3230), .B(n3229), .Z(n3235) );
  XNOR U4332 ( .A(n3231), .B(n3235), .Z(z[78]) );
  XOR U4333 ( .A(n3233), .B(n3232), .Z(n3234) );
  XNOR U4334 ( .A(n3235), .B(n3234), .Z(z[75]) );
  XOR U4335 ( .A(x[81]), .B(x[83]), .Z(n3239) );
  XOR U4336 ( .A(x[80]), .B(x[86]), .Z(n3237) );
  XNOR U4337 ( .A(n3239), .B(n3237), .Z(n3236) );
  XNOR U4338 ( .A(x[82]), .B(n3236), .Z(n3307) );
  IV U4339 ( .A(n3307), .Z(n3241) );
  XNOR U4340 ( .A(x[80]), .B(n3241), .Z(n3289) );
  XNOR U4341 ( .A(x[84]), .B(x[87]), .Z(n3238) );
  IV U4342 ( .A(n3238), .Z(n3302) );
  AND U4343 ( .A(n3289), .B(n3302), .Z(n3246) );
  XOR U4344 ( .A(x[87]), .B(x[82]), .Z(n3329) );
  XNOR U4345 ( .A(n3237), .B(x[85]), .Z(n3252) );
  IV U4346 ( .A(n3252), .Z(n3298) );
  XOR U4347 ( .A(n3239), .B(n3238), .Z(n3263) );
  IV U4348 ( .A(n3263), .Z(n3278) );
  XNOR U4349 ( .A(n3278), .B(x[80]), .Z(n3279) );
  XNOR U4350 ( .A(n3298), .B(n3279), .Z(n3291) );
  NAND U4351 ( .A(n3329), .B(n3291), .Z(n3240) );
  XNOR U4352 ( .A(n3246), .B(n3240), .Z(n3259) );
  XOR U4353 ( .A(x[81]), .B(x[87]), .Z(n3297) );
  XOR U4354 ( .A(n3241), .B(n3298), .Z(n3287) );
  ANDN U4355 ( .B(n3297), .A(n3287), .Z(n3248) );
  XOR U4356 ( .A(x[87]), .B(n3298), .Z(n3340) );
  IV U4357 ( .A(n3340), .Z(n3251) );
  NAND U4358 ( .A(n3241), .B(n3251), .Z(n3242) );
  XOR U4359 ( .A(n3248), .B(n3242), .Z(n3243) );
  XNOR U4360 ( .A(n3259), .B(n3243), .Z(n3283) );
  NANDN U4361 ( .A(x[81]), .B(n3252), .Z(n3250) );
  XNOR U4362 ( .A(n3278), .B(n3287), .Z(n3322) );
  XOR U4363 ( .A(x[84]), .B(x[82]), .Z(n3305) );
  AND U4364 ( .A(n3322), .B(n3305), .Z(n3245) );
  XNOR U4365 ( .A(n3307), .B(n3340), .Z(n3244) );
  XNOR U4366 ( .A(n3245), .B(n3244), .Z(n3247) );
  XOR U4367 ( .A(n3247), .B(n3246), .Z(n3267) );
  XNOR U4368 ( .A(n3248), .B(n3267), .Z(n3249) );
  XNOR U4369 ( .A(n3250), .B(n3249), .Z(n3281) );
  IV U4370 ( .A(n3281), .Z(n3284) );
  NAND U4371 ( .A(n3283), .B(n3284), .Z(n3277) );
  NANDN U4372 ( .A(n3283), .B(n3284), .Z(n3271) );
  XNOR U4373 ( .A(x[82]), .B(n3251), .Z(n3258) );
  XNOR U4374 ( .A(x[81]), .B(n3258), .Z(n3262) );
  IV U4375 ( .A(n3262), .Z(n3316) );
  XNOR U4376 ( .A(x[84]), .B(n3252), .Z(n3328) );
  OR U4377 ( .A(x[80]), .B(n3328), .Z(n3253) );
  XNOR U4378 ( .A(n3316), .B(n3253), .Z(n3254) );
  NANDN U4379 ( .A(n3263), .B(n3254), .Z(n3257) );
  ANDN U4380 ( .B(x[80]), .A(n3328), .Z(n3255) );
  NAND U4381 ( .A(n3263), .B(n3255), .Z(n3256) );
  NAND U4382 ( .A(n3257), .B(n3256), .Z(n3261) );
  XNOR U4383 ( .A(n3259), .B(n3258), .Z(n3260) );
  XOR U4384 ( .A(n3261), .B(n3260), .Z(n3285) );
  IV U4385 ( .A(n3283), .Z(n3282) );
  ANDN U4386 ( .B(n3285), .A(n3282), .Z(n3268) );
  AND U4387 ( .A(x[80]), .B(n3262), .Z(n3265) );
  NAND U4388 ( .A(n3263), .B(n3328), .Z(n3264) );
  XNOR U4389 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U4390 ( .A(n3267), .B(n3266), .Z(n3286) );
  XNOR U4391 ( .A(n3268), .B(n3286), .Z(n3269) );
  NAND U4392 ( .A(n3281), .B(n3269), .Z(n3270) );
  NAND U4393 ( .A(n3271), .B(n3270), .Z(n3315) );
  IV U4394 ( .A(n3315), .Z(n3290) );
  OR U4395 ( .A(n3285), .B(n3281), .Z(n3272) );
  NAND U4396 ( .A(n3282), .B(n3272), .Z(n3275) );
  XOR U4397 ( .A(n3285), .B(n3286), .Z(n3273) );
  NANDN U4398 ( .A(n3284), .B(n3273), .Z(n3274) );
  NAND U4399 ( .A(n3275), .B(n3274), .Z(n3327) );
  NANDN U4400 ( .A(n3290), .B(n3327), .Z(n3276) );
  AND U4401 ( .A(n3277), .B(n3276), .Z(n3318) );
  AND U4402 ( .A(n3318), .B(n3278), .Z(n3293) );
  OR U4403 ( .A(n3279), .B(n3290), .Z(n3280) );
  XNOR U4404 ( .A(n3293), .B(n3280), .Z(n3326) );
  XOR U4405 ( .A(n3341), .B(n3300), .Z(n3296) );
  ANDN U4406 ( .B(n3296), .A(n3287), .Z(n3308) );
  NAND U4407 ( .A(n3298), .B(n3300), .Z(n3288) );
  XNOR U4408 ( .A(n3308), .B(n3288), .Z(n3333) );
  XNOR U4409 ( .A(n3326), .B(n3333), .Z(z[82]) );
  AND U4410 ( .A(x[80]), .B(n3327), .Z(n3295) );
  AND U4411 ( .A(n3289), .B(n3304), .Z(n3325) );
  XOR U4412 ( .A(n3290), .B(n3300), .Z(n3303) );
  IV U4413 ( .A(n3303), .Z(n3330) );
  NAND U4414 ( .A(n3330), .B(n3291), .Z(n3292) );
  XNOR U4415 ( .A(n3325), .B(n3292), .Z(n3309) );
  XNOR U4416 ( .A(n3293), .B(n3309), .Z(n3294) );
  XNOR U4417 ( .A(n3295), .B(n3294), .Z(n3958) );
  AND U4418 ( .A(n3297), .B(n3296), .Z(n3342) );
  XOR U4419 ( .A(x[81]), .B(n3298), .Z(n3299) );
  NAND U4420 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U4421 ( .A(n3342), .B(n3301), .Z(n3313) );
  AND U4422 ( .A(n3304), .B(n3302), .Z(n3332) );
  XNOR U4423 ( .A(n3304), .B(n3303), .Z(n3323) );
  NAND U4424 ( .A(n3323), .B(n3305), .Z(n3306) );
  XNOR U4425 ( .A(n3332), .B(n3306), .Z(n3319) );
  AND U4426 ( .A(n3341), .B(n3307), .Z(n3311) );
  XNOR U4427 ( .A(n3309), .B(n3308), .Z(n3310) );
  XNOR U4428 ( .A(n3311), .B(n3310), .Z(n3957) );
  XNOR U4429 ( .A(n3319), .B(n3957), .Z(n3312) );
  XNOR U4430 ( .A(n3313), .B(n3312), .Z(n3314) );
  XNOR U4431 ( .A(n3958), .B(n3314), .Z(z[85]) );
  AND U4432 ( .A(n3316), .B(n3315), .Z(n3321) );
  XOR U4433 ( .A(n3316), .B(n3328), .Z(n3317) );
  AND U4434 ( .A(n3318), .B(n3317), .Z(n3337) );
  XNOR U4435 ( .A(n3319), .B(n3337), .Z(n3320) );
  XNOR U4436 ( .A(n3321), .B(n3320), .Z(n3348) );
  NAND U4437 ( .A(n3323), .B(n3322), .Z(n3324) );
  XNOR U4438 ( .A(n3325), .B(n3324), .Z(n3336) );
  XNOR U4439 ( .A(n3326), .B(n3336), .Z(n3956) );
  XNOR U4440 ( .A(n3348), .B(n3956), .Z(n3346) );
  AND U4441 ( .A(n3328), .B(n3327), .Z(n3335) );
  NAND U4442 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U4443 ( .A(n3332), .B(n3331), .Z(n3343) );
  XNOR U4444 ( .A(n3343), .B(n3333), .Z(n3334) );
  XNOR U4445 ( .A(n3335), .B(n3334), .Z(n3339) );
  XNOR U4446 ( .A(n3337), .B(n3336), .Z(n3338) );
  XNOR U4447 ( .A(n3339), .B(n3338), .Z(n3347) );
  XNOR U4448 ( .A(n3346), .B(n3347), .Z(z[81]) );
  AND U4449 ( .A(n3341), .B(n3340), .Z(n3345) );
  XNOR U4450 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U4451 ( .A(n3345), .B(n3344), .Z(n3350) );
  XNOR U4452 ( .A(n3346), .B(n3350), .Z(z[86]) );
  XOR U4453 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4454 ( .A(n3350), .B(n3349), .Z(z[83]) );
  XOR U4455 ( .A(x[89]), .B(x[91]), .Z(n3354) );
  XOR U4456 ( .A(x[88]), .B(x[94]), .Z(n3352) );
  XNOR U4457 ( .A(n3354), .B(n3352), .Z(n3351) );
  XNOR U4458 ( .A(x[90]), .B(n3351), .Z(n3422) );
  IV U4459 ( .A(n3422), .Z(n3356) );
  XNOR U4460 ( .A(x[88]), .B(n3356), .Z(n3404) );
  XNOR U4461 ( .A(x[92]), .B(x[95]), .Z(n3353) );
  IV U4462 ( .A(n3353), .Z(n3417) );
  AND U4463 ( .A(n3404), .B(n3417), .Z(n3361) );
  XOR U4464 ( .A(x[95]), .B(x[90]), .Z(n3444) );
  XNOR U4465 ( .A(n3352), .B(x[93]), .Z(n3367) );
  IV U4466 ( .A(n3367), .Z(n3413) );
  XOR U4467 ( .A(n3354), .B(n3353), .Z(n3378) );
  IV U4468 ( .A(n3378), .Z(n3393) );
  XNOR U4469 ( .A(n3393), .B(x[88]), .Z(n3394) );
  XNOR U4470 ( .A(n3413), .B(n3394), .Z(n3406) );
  NAND U4471 ( .A(n3444), .B(n3406), .Z(n3355) );
  XNOR U4472 ( .A(n3361), .B(n3355), .Z(n3374) );
  XOR U4473 ( .A(x[89]), .B(x[95]), .Z(n3412) );
  XOR U4474 ( .A(n3356), .B(n3413), .Z(n3402) );
  ANDN U4475 ( .B(n3412), .A(n3402), .Z(n3363) );
  XOR U4476 ( .A(x[95]), .B(n3413), .Z(n3455) );
  IV U4477 ( .A(n3455), .Z(n3366) );
  NAND U4478 ( .A(n3356), .B(n3366), .Z(n3357) );
  XOR U4479 ( .A(n3363), .B(n3357), .Z(n3358) );
  XNOR U4480 ( .A(n3374), .B(n3358), .Z(n3398) );
  NANDN U4481 ( .A(x[89]), .B(n3367), .Z(n3365) );
  XNOR U4482 ( .A(n3393), .B(n3402), .Z(n3437) );
  XOR U4483 ( .A(x[92]), .B(x[90]), .Z(n3420) );
  AND U4484 ( .A(n3437), .B(n3420), .Z(n3360) );
  XNOR U4485 ( .A(n3422), .B(n3455), .Z(n3359) );
  XNOR U4486 ( .A(n3360), .B(n3359), .Z(n3362) );
  XOR U4487 ( .A(n3362), .B(n3361), .Z(n3382) );
  XNOR U4488 ( .A(n3363), .B(n3382), .Z(n3364) );
  XNOR U4489 ( .A(n3365), .B(n3364), .Z(n3396) );
  IV U4490 ( .A(n3396), .Z(n3399) );
  NAND U4491 ( .A(n3398), .B(n3399), .Z(n3392) );
  NANDN U4492 ( .A(n3398), .B(n3399), .Z(n3386) );
  XNOR U4493 ( .A(x[90]), .B(n3366), .Z(n3373) );
  XNOR U4494 ( .A(x[89]), .B(n3373), .Z(n3377) );
  IV U4495 ( .A(n3377), .Z(n3431) );
  XNOR U4496 ( .A(x[92]), .B(n3367), .Z(n3443) );
  OR U4497 ( .A(x[88]), .B(n3443), .Z(n3368) );
  XNOR U4498 ( .A(n3431), .B(n3368), .Z(n3369) );
  NANDN U4499 ( .A(n3378), .B(n3369), .Z(n3372) );
  ANDN U4500 ( .B(x[88]), .A(n3443), .Z(n3370) );
  NAND U4501 ( .A(n3378), .B(n3370), .Z(n3371) );
  NAND U4502 ( .A(n3372), .B(n3371), .Z(n3376) );
  XNOR U4503 ( .A(n3374), .B(n3373), .Z(n3375) );
  XOR U4504 ( .A(n3376), .B(n3375), .Z(n3400) );
  IV U4505 ( .A(n3398), .Z(n3397) );
  ANDN U4506 ( .B(n3400), .A(n3397), .Z(n3383) );
  AND U4507 ( .A(x[88]), .B(n3377), .Z(n3380) );
  NAND U4508 ( .A(n3378), .B(n3443), .Z(n3379) );
  XNOR U4509 ( .A(n3380), .B(n3379), .Z(n3381) );
  XNOR U4510 ( .A(n3382), .B(n3381), .Z(n3401) );
  XNOR U4511 ( .A(n3383), .B(n3401), .Z(n3384) );
  NAND U4512 ( .A(n3396), .B(n3384), .Z(n3385) );
  NAND U4513 ( .A(n3386), .B(n3385), .Z(n3430) );
  IV U4514 ( .A(n3430), .Z(n3405) );
  OR U4515 ( .A(n3400), .B(n3396), .Z(n3387) );
  NAND U4516 ( .A(n3397), .B(n3387), .Z(n3390) );
  XOR U4517 ( .A(n3400), .B(n3401), .Z(n3388) );
  NANDN U4518 ( .A(n3399), .B(n3388), .Z(n3389) );
  NAND U4519 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U4520 ( .A(n3405), .B(n3442), .Z(n3391) );
  AND U4521 ( .A(n3392), .B(n3391), .Z(n3433) );
  AND U4522 ( .A(n3433), .B(n3393), .Z(n3408) );
  OR U4523 ( .A(n3394), .B(n3405), .Z(n3395) );
  XNOR U4524 ( .A(n3408), .B(n3395), .Z(n3441) );
  XOR U4525 ( .A(n3456), .B(n3415), .Z(n3411) );
  ANDN U4526 ( .B(n3411), .A(n3402), .Z(n3423) );
  NAND U4527 ( .A(n3413), .B(n3415), .Z(n3403) );
  XNOR U4528 ( .A(n3423), .B(n3403), .Z(n3448) );
  XNOR U4529 ( .A(n3441), .B(n3448), .Z(z[90]) );
  AND U4530 ( .A(x[88]), .B(n3442), .Z(n3410) );
  AND U4531 ( .A(n3404), .B(n3419), .Z(n3440) );
  XOR U4532 ( .A(n3405), .B(n3415), .Z(n3418) );
  IV U4533 ( .A(n3418), .Z(n3445) );
  NAND U4534 ( .A(n3445), .B(n3406), .Z(n3407) );
  XNOR U4535 ( .A(n3440), .B(n3407), .Z(n3424) );
  XNOR U4536 ( .A(n3408), .B(n3424), .Z(n3409) );
  XNOR U4537 ( .A(n3410), .B(n3409), .Z(n3963) );
  AND U4538 ( .A(n3412), .B(n3411), .Z(n3457) );
  XOR U4539 ( .A(x[89]), .B(n3413), .Z(n3414) );
  NAND U4540 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4541 ( .A(n3457), .B(n3416), .Z(n3428) );
  AND U4542 ( .A(n3419), .B(n3417), .Z(n3447) );
  XNOR U4543 ( .A(n3419), .B(n3418), .Z(n3438) );
  NAND U4544 ( .A(n3438), .B(n3420), .Z(n3421) );
  XNOR U4545 ( .A(n3447), .B(n3421), .Z(n3434) );
  AND U4546 ( .A(n3456), .B(n3422), .Z(n3426) );
  XNOR U4547 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4548 ( .A(n3426), .B(n3425), .Z(n3962) );
  XNOR U4549 ( .A(n3434), .B(n3962), .Z(n3427) );
  XNOR U4550 ( .A(n3428), .B(n3427), .Z(n3429) );
  XNOR U4551 ( .A(n3963), .B(n3429), .Z(z[93]) );
  AND U4552 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4553 ( .A(n3431), .B(n3443), .Z(n3432) );
  AND U4554 ( .A(n3433), .B(n3432), .Z(n3452) );
  XNOR U4555 ( .A(n3434), .B(n3452), .Z(n3435) );
  XNOR U4556 ( .A(n3436), .B(n3435), .Z(n3463) );
  NAND U4557 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U4558 ( .A(n3440), .B(n3439), .Z(n3451) );
  XNOR U4559 ( .A(n3441), .B(n3451), .Z(n3959) );
  XNOR U4560 ( .A(n3463), .B(n3959), .Z(n3461) );
  AND U4561 ( .A(n3443), .B(n3442), .Z(n3450) );
  NAND U4562 ( .A(n3445), .B(n3444), .Z(n3446) );
  XNOR U4563 ( .A(n3447), .B(n3446), .Z(n3458) );
  XNOR U4564 ( .A(n3458), .B(n3448), .Z(n3449) );
  XNOR U4565 ( .A(n3450), .B(n3449), .Z(n3454) );
  XNOR U4566 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U4567 ( .A(n3454), .B(n3453), .Z(n3462) );
  XNOR U4568 ( .A(n3461), .B(n3462), .Z(z[89]) );
  AND U4569 ( .A(n3456), .B(n3455), .Z(n3460) );
  XNOR U4570 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U4571 ( .A(n3460), .B(n3459), .Z(n3465) );
  XNOR U4572 ( .A(n3461), .B(n3465), .Z(z[94]) );
  XOR U4573 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4574 ( .A(n3465), .B(n3464), .Z(z[91]) );
  XNOR U4575 ( .A(x[102]), .B(x[96]), .Z(n3471) );
  XNOR U4576 ( .A(x[101]), .B(n3471), .Z(n3537) );
  IV U4577 ( .A(n3537), .Z(n3475) );
  XOR U4578 ( .A(x[103]), .B(n3475), .Z(n3468) );
  IV U4579 ( .A(n3468), .Z(n3491) );
  XOR U4580 ( .A(x[97]), .B(x[99]), .Z(n3466) );
  XNOR U4581 ( .A(x[98]), .B(n3466), .Z(n3470) );
  XNOR U4582 ( .A(x[102]), .B(n3470), .Z(n3519) );
  XOR U4583 ( .A(x[100]), .B(x[103]), .Z(n3496) );
  AND U4584 ( .A(n3519), .B(n3496), .Z(n3478) );
  XOR U4585 ( .A(n3466), .B(n3496), .Z(n3543) );
  XOR U4586 ( .A(x[96]), .B(n3543), .Z(n3554) );
  XOR U4587 ( .A(n3537), .B(n3554), .Z(n3911) );
  XOR U4588 ( .A(x[98]), .B(x[103]), .Z(n3509) );
  NAND U4589 ( .A(n3911), .B(n3509), .Z(n3467) );
  XNOR U4590 ( .A(n3478), .B(n3467), .Z(n3472) );
  XNOR U4591 ( .A(x[98]), .B(n3468), .Z(n3469) );
  XOR U4592 ( .A(x[97]), .B(n3469), .Z(n3528) );
  XNOR U4593 ( .A(x[100]), .B(n3475), .Z(n3514) );
  IV U4594 ( .A(n3497), .Z(n3498) );
  XOR U4595 ( .A(x[97]), .B(x[103]), .Z(n3511) );
  XNOR U4596 ( .A(x[101]), .B(n3470), .Z(n3524) );
  AND U4597 ( .A(n3511), .B(n3524), .Z(n3480) );
  NOR U4598 ( .A(n3491), .B(n3546), .Z(n3473) );
  XNOR U4599 ( .A(n3473), .B(n3472), .Z(n3474) );
  XNOR U4600 ( .A(n3480), .B(n3474), .Z(n3502) );
  NANDN U4601 ( .A(x[97]), .B(n3475), .Z(n3482) );
  XOR U4602 ( .A(x[98]), .B(x[100]), .Z(n3529) );
  AND U4603 ( .A(n3529), .B(n3521), .Z(n3477) );
  XNOR U4604 ( .A(n3491), .B(n3546), .Z(n3476) );
  XNOR U4605 ( .A(n3477), .B(n3476), .Z(n3479) );
  XOR U4606 ( .A(n3479), .B(n3478), .Z(n3485) );
  XNOR U4607 ( .A(n3485), .B(n3480), .Z(n3481) );
  XNOR U4608 ( .A(n3482), .B(n3481), .Z(n3506) );
  XOR U4609 ( .A(n3502), .B(n3506), .Z(n3483) );
  NAND U4610 ( .A(n3498), .B(n3483), .Z(n3490) );
  ANDN U4611 ( .B(n3514), .A(n3543), .Z(n3487) );
  ANDN U4612 ( .B(x[96]), .A(n3528), .Z(n3484) );
  XNOR U4613 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4614 ( .A(n3487), .B(n3486), .Z(n3503) );
  NANDN U4615 ( .A(n3498), .B(n3502), .Z(n3488) );
  NANDN U4616 ( .A(n3503), .B(n3488), .Z(n3489) );
  NAND U4617 ( .A(n3490), .B(n3489), .Z(n3547) );
  ANDN U4618 ( .B(n3491), .A(n3547), .Z(n3513) );
  XOR U4619 ( .A(n3497), .B(n3503), .Z(n3492) );
  NAND U4620 ( .A(n3506), .B(n3492), .Z(n3495) );
  OR U4621 ( .A(n3506), .B(n3498), .Z(n3493) );
  NANDN U4622 ( .A(n3502), .B(n3493), .Z(n3494) );
  NAND U4623 ( .A(n3495), .B(n3494), .Z(n3544) );
  XNOR U4624 ( .A(n3547), .B(n3544), .Z(n3520) );
  AND U4625 ( .A(n3496), .B(n3520), .Z(n3532) );
  NANDN U4626 ( .A(n3503), .B(n3497), .Z(n3501) );
  AND U4627 ( .A(n3502), .B(n3498), .Z(n3504) );
  XOR U4628 ( .A(n3506), .B(n3504), .Z(n3499) );
  NAND U4629 ( .A(n3503), .B(n3499), .Z(n3500) );
  NAND U4630 ( .A(n3501), .B(n3500), .Z(n3539) );
  OR U4631 ( .A(n3506), .B(n3502), .Z(n3508) );
  XOR U4632 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U4633 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U4634 ( .A(n3508), .B(n3507), .Z(n3555) );
  XOR U4635 ( .A(n3539), .B(n3555), .Z(n3912) );
  NAND U4636 ( .A(n3912), .B(n3509), .Z(n3510) );
  XNOR U4637 ( .A(n3532), .B(n3510), .Z(n3516) );
  XNOR U4638 ( .A(n3547), .B(n3539), .Z(n3523) );
  AND U4639 ( .A(n3511), .B(n3523), .Z(n3541) );
  XNOR U4640 ( .A(n3516), .B(n3541), .Z(n3512) );
  XNOR U4641 ( .A(n3513), .B(n3512), .Z(n3561) );
  AND U4642 ( .A(n3514), .B(n3544), .Z(n3518) );
  XOR U4643 ( .A(n3528), .B(n3514), .Z(n3515) );
  AND U4644 ( .A(n3542), .B(n3515), .Z(n3533) );
  XNOR U4645 ( .A(n3516), .B(n3533), .Z(n3517) );
  XNOR U4646 ( .A(n3518), .B(n3517), .Z(n3527) );
  AND U4647 ( .A(n3519), .B(n3520), .Z(n3916) );
  NAND U4648 ( .A(n3530), .B(n3521), .Z(n3522) );
  XNOR U4649 ( .A(n3916), .B(n3522), .Z(n3558) );
  AND U4650 ( .A(n3524), .B(n3523), .Z(n3549) );
  NAND U4651 ( .A(n3537), .B(n3539), .Z(n3525) );
  XNOR U4652 ( .A(n3549), .B(n3525), .Z(n3564) );
  XNOR U4653 ( .A(n3558), .B(n3564), .Z(n3526) );
  XNOR U4654 ( .A(n3527), .B(n3526), .Z(n3560) );
  AND U4655 ( .A(n3528), .B(n3555), .Z(n3535) );
  NAND U4656 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U4657 ( .A(n3532), .B(n3531), .Z(n3553) );
  XNOR U4658 ( .A(n3533), .B(n3553), .Z(n3534) );
  XNOR U4659 ( .A(n3535), .B(n3534), .Z(n3559) );
  XOR U4660 ( .A(n3560), .B(n3559), .Z(n3536) );
  XNOR U4661 ( .A(n3561), .B(n3536), .Z(z[99]) );
  XOR U4662 ( .A(x[97]), .B(n3537), .Z(n3538) );
  NAND U4663 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U4664 ( .A(n3541), .B(n3540), .Z(n3551) );
  AND U4665 ( .A(n3543), .B(n3542), .Z(n3557) );
  NAND U4666 ( .A(n3544), .B(x[96]), .Z(n3545) );
  XNOR U4667 ( .A(n3557), .B(n3545), .Z(n3915) );
  NANDN U4668 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U4669 ( .A(n3549), .B(n3548), .Z(n3913) );
  XNOR U4670 ( .A(n3915), .B(n3913), .Z(n3550) );
  XNOR U4671 ( .A(n3551), .B(n3550), .Z(n3552) );
  XNOR U4672 ( .A(n3553), .B(n3552), .Z(z[101]) );
  NAND U4673 ( .A(n3555), .B(n3554), .Z(n3556) );
  XNOR U4674 ( .A(n3557), .B(n3556), .Z(n3563) );
  XNOR U4675 ( .A(n3558), .B(n3563), .Z(n3964) );
  XNOR U4676 ( .A(n3559), .B(n3964), .Z(n3562) );
  XNOR U4677 ( .A(n3560), .B(n3562), .Z(z[97]) );
  XNOR U4678 ( .A(n3562), .B(n3561), .Z(z[102]) );
  XNOR U4679 ( .A(n3564), .B(n3563), .Z(z[98]) );
  XOR U4680 ( .A(x[105]), .B(x[107]), .Z(n3568) );
  XOR U4681 ( .A(x[104]), .B(x[110]), .Z(n3566) );
  XNOR U4682 ( .A(n3568), .B(n3566), .Z(n3565) );
  XNOR U4683 ( .A(x[106]), .B(n3565), .Z(n3636) );
  IV U4684 ( .A(n3636), .Z(n3570) );
  XNOR U4685 ( .A(x[104]), .B(n3570), .Z(n3618) );
  XNOR U4686 ( .A(x[108]), .B(x[111]), .Z(n3567) );
  IV U4687 ( .A(n3567), .Z(n3631) );
  AND U4688 ( .A(n3618), .B(n3631), .Z(n3575) );
  XOR U4689 ( .A(x[111]), .B(x[106]), .Z(n3658) );
  XNOR U4690 ( .A(n3566), .B(x[109]), .Z(n3581) );
  IV U4691 ( .A(n3581), .Z(n3627) );
  XOR U4692 ( .A(n3568), .B(n3567), .Z(n3592) );
  IV U4693 ( .A(n3592), .Z(n3607) );
  XNOR U4694 ( .A(n3607), .B(x[104]), .Z(n3608) );
  XNOR U4695 ( .A(n3627), .B(n3608), .Z(n3620) );
  NAND U4696 ( .A(n3658), .B(n3620), .Z(n3569) );
  XNOR U4697 ( .A(n3575), .B(n3569), .Z(n3588) );
  XOR U4698 ( .A(x[105]), .B(x[111]), .Z(n3626) );
  XOR U4699 ( .A(n3570), .B(n3627), .Z(n3616) );
  ANDN U4700 ( .B(n3626), .A(n3616), .Z(n3577) );
  XOR U4701 ( .A(x[111]), .B(n3627), .Z(n3669) );
  IV U4702 ( .A(n3669), .Z(n3580) );
  NAND U4703 ( .A(n3570), .B(n3580), .Z(n3571) );
  XOR U4704 ( .A(n3577), .B(n3571), .Z(n3572) );
  XNOR U4705 ( .A(n3588), .B(n3572), .Z(n3612) );
  NANDN U4706 ( .A(x[105]), .B(n3581), .Z(n3579) );
  XNOR U4707 ( .A(n3607), .B(n3616), .Z(n3651) );
  XOR U4708 ( .A(x[108]), .B(x[106]), .Z(n3634) );
  AND U4709 ( .A(n3651), .B(n3634), .Z(n3574) );
  XNOR U4710 ( .A(n3636), .B(n3669), .Z(n3573) );
  XNOR U4711 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U4712 ( .A(n3576), .B(n3575), .Z(n3596) );
  XNOR U4713 ( .A(n3577), .B(n3596), .Z(n3578) );
  XNOR U4714 ( .A(n3579), .B(n3578), .Z(n3610) );
  IV U4715 ( .A(n3610), .Z(n3613) );
  NAND U4716 ( .A(n3612), .B(n3613), .Z(n3606) );
  NANDN U4717 ( .A(n3612), .B(n3613), .Z(n3600) );
  XNOR U4718 ( .A(x[106]), .B(n3580), .Z(n3587) );
  XNOR U4719 ( .A(x[105]), .B(n3587), .Z(n3591) );
  IV U4720 ( .A(n3591), .Z(n3645) );
  XNOR U4721 ( .A(x[108]), .B(n3581), .Z(n3657) );
  OR U4722 ( .A(x[104]), .B(n3657), .Z(n3582) );
  XNOR U4723 ( .A(n3645), .B(n3582), .Z(n3583) );
  NANDN U4724 ( .A(n3592), .B(n3583), .Z(n3586) );
  ANDN U4725 ( .B(x[104]), .A(n3657), .Z(n3584) );
  NAND U4726 ( .A(n3592), .B(n3584), .Z(n3585) );
  NAND U4727 ( .A(n3586), .B(n3585), .Z(n3590) );
  XNOR U4728 ( .A(n3588), .B(n3587), .Z(n3589) );
  XOR U4729 ( .A(n3590), .B(n3589), .Z(n3614) );
  IV U4730 ( .A(n3612), .Z(n3611) );
  ANDN U4731 ( .B(n3614), .A(n3611), .Z(n3597) );
  AND U4732 ( .A(x[104]), .B(n3591), .Z(n3594) );
  NAND U4733 ( .A(n3592), .B(n3657), .Z(n3593) );
  XNOR U4734 ( .A(n3594), .B(n3593), .Z(n3595) );
  XNOR U4735 ( .A(n3596), .B(n3595), .Z(n3615) );
  XNOR U4736 ( .A(n3597), .B(n3615), .Z(n3598) );
  NAND U4737 ( .A(n3610), .B(n3598), .Z(n3599) );
  NAND U4738 ( .A(n3600), .B(n3599), .Z(n3644) );
  IV U4739 ( .A(n3644), .Z(n3619) );
  OR U4740 ( .A(n3614), .B(n3610), .Z(n3601) );
  NAND U4741 ( .A(n3611), .B(n3601), .Z(n3604) );
  XOR U4742 ( .A(n3614), .B(n3615), .Z(n3602) );
  NANDN U4743 ( .A(n3613), .B(n3602), .Z(n3603) );
  NAND U4744 ( .A(n3604), .B(n3603), .Z(n3656) );
  NANDN U4745 ( .A(n3619), .B(n3656), .Z(n3605) );
  AND U4746 ( .A(n3606), .B(n3605), .Z(n3647) );
  AND U4747 ( .A(n3647), .B(n3607), .Z(n3622) );
  OR U4748 ( .A(n3608), .B(n3619), .Z(n3609) );
  XNOR U4749 ( .A(n3622), .B(n3609), .Z(n3655) );
  XOR U4750 ( .A(n3670), .B(n3629), .Z(n3625) );
  ANDN U4751 ( .B(n3625), .A(n3616), .Z(n3637) );
  NAND U4752 ( .A(n3627), .B(n3629), .Z(n3617) );
  XNOR U4753 ( .A(n3637), .B(n3617), .Z(n3662) );
  XNOR U4754 ( .A(n3655), .B(n3662), .Z(z[106]) );
  AND U4755 ( .A(x[104]), .B(n3656), .Z(n3624) );
  AND U4756 ( .A(n3618), .B(n3633), .Z(n3654) );
  XOR U4757 ( .A(n3619), .B(n3629), .Z(n3632) );
  IV U4758 ( .A(n3632), .Z(n3659) );
  NAND U4759 ( .A(n3659), .B(n3620), .Z(n3621) );
  XNOR U4760 ( .A(n3654), .B(n3621), .Z(n3638) );
  XNOR U4761 ( .A(n3622), .B(n3638), .Z(n3623) );
  XNOR U4762 ( .A(n3624), .B(n3623), .Z(n3922) );
  AND U4763 ( .A(n3626), .B(n3625), .Z(n3671) );
  XOR U4764 ( .A(x[105]), .B(n3627), .Z(n3628) );
  NAND U4765 ( .A(n3629), .B(n3628), .Z(n3630) );
  XNOR U4766 ( .A(n3671), .B(n3630), .Z(n3642) );
  AND U4767 ( .A(n3633), .B(n3631), .Z(n3661) );
  XNOR U4768 ( .A(n3633), .B(n3632), .Z(n3652) );
  NAND U4769 ( .A(n3652), .B(n3634), .Z(n3635) );
  XNOR U4770 ( .A(n3661), .B(n3635), .Z(n3648) );
  AND U4771 ( .A(n3670), .B(n3636), .Z(n3640) );
  XNOR U4772 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U4773 ( .A(n3640), .B(n3639), .Z(n3921) );
  XNOR U4774 ( .A(n3648), .B(n3921), .Z(n3641) );
  XNOR U4775 ( .A(n3642), .B(n3641), .Z(n3643) );
  XNOR U4776 ( .A(n3922), .B(n3643), .Z(z[109]) );
  AND U4777 ( .A(n3645), .B(n3644), .Z(n3650) );
  XOR U4778 ( .A(n3645), .B(n3657), .Z(n3646) );
  AND U4779 ( .A(n3647), .B(n3646), .Z(n3666) );
  XNOR U4780 ( .A(n3648), .B(n3666), .Z(n3649) );
  XNOR U4781 ( .A(n3650), .B(n3649), .Z(n3677) );
  NAND U4782 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U4783 ( .A(n3654), .B(n3653), .Z(n3665) );
  XNOR U4784 ( .A(n3655), .B(n3665), .Z(n3920) );
  XNOR U4785 ( .A(n3677), .B(n3920), .Z(n3675) );
  AND U4786 ( .A(n3657), .B(n3656), .Z(n3664) );
  NAND U4787 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4788 ( .A(n3661), .B(n3660), .Z(n3672) );
  XNOR U4789 ( .A(n3672), .B(n3662), .Z(n3663) );
  XNOR U4790 ( .A(n3664), .B(n3663), .Z(n3668) );
  XNOR U4791 ( .A(n3666), .B(n3665), .Z(n3667) );
  XNOR U4792 ( .A(n3668), .B(n3667), .Z(n3676) );
  XNOR U4793 ( .A(n3675), .B(n3676), .Z(z[105]) );
  AND U4794 ( .A(n3670), .B(n3669), .Z(n3674) );
  XNOR U4795 ( .A(n3672), .B(n3671), .Z(n3673) );
  XNOR U4796 ( .A(n3674), .B(n3673), .Z(n3679) );
  XNOR U4797 ( .A(n3675), .B(n3679), .Z(z[110]) );
  XOR U4798 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4799 ( .A(n3679), .B(n3678), .Z(z[107]) );
  XOR U4800 ( .A(x[113]), .B(x[115]), .Z(n3683) );
  XOR U4801 ( .A(x[112]), .B(x[118]), .Z(n3681) );
  XNOR U4802 ( .A(n3683), .B(n3681), .Z(n3680) );
  XNOR U4803 ( .A(x[114]), .B(n3680), .Z(n3751) );
  IV U4804 ( .A(n3751), .Z(n3685) );
  XNOR U4805 ( .A(x[112]), .B(n3685), .Z(n3733) );
  XNOR U4806 ( .A(x[116]), .B(x[119]), .Z(n3682) );
  IV U4807 ( .A(n3682), .Z(n3746) );
  AND U4808 ( .A(n3733), .B(n3746), .Z(n3690) );
  XOR U4809 ( .A(x[119]), .B(x[114]), .Z(n3773) );
  XNOR U4810 ( .A(n3681), .B(x[117]), .Z(n3696) );
  IV U4811 ( .A(n3696), .Z(n3742) );
  XOR U4812 ( .A(n3683), .B(n3682), .Z(n3707) );
  IV U4813 ( .A(n3707), .Z(n3722) );
  XNOR U4814 ( .A(n3722), .B(x[112]), .Z(n3723) );
  XNOR U4815 ( .A(n3742), .B(n3723), .Z(n3735) );
  NAND U4816 ( .A(n3773), .B(n3735), .Z(n3684) );
  XNOR U4817 ( .A(n3690), .B(n3684), .Z(n3703) );
  XOR U4818 ( .A(x[113]), .B(x[119]), .Z(n3741) );
  XOR U4819 ( .A(n3685), .B(n3742), .Z(n3731) );
  ANDN U4820 ( .B(n3741), .A(n3731), .Z(n3692) );
  XOR U4821 ( .A(x[119]), .B(n3742), .Z(n3784) );
  IV U4822 ( .A(n3784), .Z(n3695) );
  NAND U4823 ( .A(n3685), .B(n3695), .Z(n3686) );
  XOR U4824 ( .A(n3692), .B(n3686), .Z(n3687) );
  XNOR U4825 ( .A(n3703), .B(n3687), .Z(n3727) );
  NANDN U4826 ( .A(x[113]), .B(n3696), .Z(n3694) );
  XNOR U4827 ( .A(n3722), .B(n3731), .Z(n3766) );
  XOR U4828 ( .A(x[116]), .B(x[114]), .Z(n3749) );
  AND U4829 ( .A(n3766), .B(n3749), .Z(n3689) );
  XNOR U4830 ( .A(n3751), .B(n3784), .Z(n3688) );
  XNOR U4831 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4832 ( .A(n3691), .B(n3690), .Z(n3711) );
  XNOR U4833 ( .A(n3692), .B(n3711), .Z(n3693) );
  XNOR U4834 ( .A(n3694), .B(n3693), .Z(n3725) );
  IV U4835 ( .A(n3725), .Z(n3728) );
  NAND U4836 ( .A(n3727), .B(n3728), .Z(n3721) );
  NANDN U4837 ( .A(n3727), .B(n3728), .Z(n3715) );
  XNOR U4838 ( .A(x[114]), .B(n3695), .Z(n3702) );
  XNOR U4839 ( .A(x[113]), .B(n3702), .Z(n3706) );
  IV U4840 ( .A(n3706), .Z(n3760) );
  XNOR U4841 ( .A(x[116]), .B(n3696), .Z(n3772) );
  OR U4842 ( .A(x[112]), .B(n3772), .Z(n3697) );
  XNOR U4843 ( .A(n3760), .B(n3697), .Z(n3698) );
  NANDN U4844 ( .A(n3707), .B(n3698), .Z(n3701) );
  ANDN U4845 ( .B(x[112]), .A(n3772), .Z(n3699) );
  NAND U4846 ( .A(n3707), .B(n3699), .Z(n3700) );
  NAND U4847 ( .A(n3701), .B(n3700), .Z(n3705) );
  XNOR U4848 ( .A(n3703), .B(n3702), .Z(n3704) );
  XOR U4849 ( .A(n3705), .B(n3704), .Z(n3729) );
  IV U4850 ( .A(n3727), .Z(n3726) );
  ANDN U4851 ( .B(n3729), .A(n3726), .Z(n3712) );
  AND U4852 ( .A(x[112]), .B(n3706), .Z(n3709) );
  NAND U4853 ( .A(n3707), .B(n3772), .Z(n3708) );
  XNOR U4854 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U4855 ( .A(n3711), .B(n3710), .Z(n3730) );
  XNOR U4856 ( .A(n3712), .B(n3730), .Z(n3713) );
  NAND U4857 ( .A(n3725), .B(n3713), .Z(n3714) );
  NAND U4858 ( .A(n3715), .B(n3714), .Z(n3759) );
  IV U4859 ( .A(n3759), .Z(n3734) );
  OR U4860 ( .A(n3729), .B(n3725), .Z(n3716) );
  NAND U4861 ( .A(n3726), .B(n3716), .Z(n3719) );
  XOR U4862 ( .A(n3729), .B(n3730), .Z(n3717) );
  NANDN U4863 ( .A(n3728), .B(n3717), .Z(n3718) );
  NAND U4864 ( .A(n3719), .B(n3718), .Z(n3771) );
  NANDN U4865 ( .A(n3734), .B(n3771), .Z(n3720) );
  AND U4866 ( .A(n3721), .B(n3720), .Z(n3762) );
  AND U4867 ( .A(n3762), .B(n3722), .Z(n3737) );
  OR U4868 ( .A(n3723), .B(n3734), .Z(n3724) );
  XNOR U4869 ( .A(n3737), .B(n3724), .Z(n3770) );
  XOR U4870 ( .A(n3785), .B(n3744), .Z(n3740) );
  ANDN U4871 ( .B(n3740), .A(n3731), .Z(n3752) );
  NAND U4872 ( .A(n3742), .B(n3744), .Z(n3732) );
  XNOR U4873 ( .A(n3752), .B(n3732), .Z(n3777) );
  XNOR U4874 ( .A(n3770), .B(n3777), .Z(z[114]) );
  AND U4875 ( .A(x[112]), .B(n3771), .Z(n3739) );
  AND U4876 ( .A(n3733), .B(n3748), .Z(n3769) );
  XOR U4877 ( .A(n3734), .B(n3744), .Z(n3747) );
  IV U4878 ( .A(n3747), .Z(n3774) );
  NAND U4879 ( .A(n3774), .B(n3735), .Z(n3736) );
  XNOR U4880 ( .A(n3769), .B(n3736), .Z(n3753) );
  XNOR U4881 ( .A(n3737), .B(n3753), .Z(n3738) );
  XNOR U4882 ( .A(n3739), .B(n3738), .Z(n3925) );
  AND U4883 ( .A(n3741), .B(n3740), .Z(n3786) );
  XOR U4884 ( .A(x[113]), .B(n3742), .Z(n3743) );
  NAND U4885 ( .A(n3744), .B(n3743), .Z(n3745) );
  XNOR U4886 ( .A(n3786), .B(n3745), .Z(n3757) );
  AND U4887 ( .A(n3748), .B(n3746), .Z(n3776) );
  XNOR U4888 ( .A(n3748), .B(n3747), .Z(n3767) );
  NAND U4889 ( .A(n3767), .B(n3749), .Z(n3750) );
  XNOR U4890 ( .A(n3776), .B(n3750), .Z(n3763) );
  AND U4891 ( .A(n3785), .B(n3751), .Z(n3755) );
  XNOR U4892 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U4893 ( .A(n3755), .B(n3754), .Z(n3924) );
  XNOR U4894 ( .A(n3763), .B(n3924), .Z(n3756) );
  XNOR U4895 ( .A(n3757), .B(n3756), .Z(n3758) );
  XNOR U4896 ( .A(n3925), .B(n3758), .Z(z[117]) );
  AND U4897 ( .A(n3760), .B(n3759), .Z(n3765) );
  XOR U4898 ( .A(n3760), .B(n3772), .Z(n3761) );
  AND U4899 ( .A(n3762), .B(n3761), .Z(n3781) );
  XNOR U4900 ( .A(n3763), .B(n3781), .Z(n3764) );
  XNOR U4901 ( .A(n3765), .B(n3764), .Z(n3792) );
  NAND U4902 ( .A(n3767), .B(n3766), .Z(n3768) );
  XNOR U4903 ( .A(n3769), .B(n3768), .Z(n3780) );
  XNOR U4904 ( .A(n3770), .B(n3780), .Z(n3923) );
  XNOR U4905 ( .A(n3792), .B(n3923), .Z(n3790) );
  AND U4906 ( .A(n3772), .B(n3771), .Z(n3779) );
  NAND U4907 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4908 ( .A(n3776), .B(n3775), .Z(n3787) );
  XNOR U4909 ( .A(n3787), .B(n3777), .Z(n3778) );
  XNOR U4910 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4911 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR U4912 ( .A(n3783), .B(n3782), .Z(n3791) );
  XNOR U4913 ( .A(n3790), .B(n3791), .Z(z[113]) );
  AND U4914 ( .A(n3785), .B(n3784), .Z(n3789) );
  XNOR U4915 ( .A(n3787), .B(n3786), .Z(n3788) );
  XNOR U4916 ( .A(n3789), .B(n3788), .Z(n3794) );
  XNOR U4917 ( .A(n3790), .B(n3794), .Z(z[118]) );
  XOR U4918 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U4919 ( .A(n3794), .B(n3793), .Z(z[115]) );
  XOR U4920 ( .A(x[121]), .B(x[123]), .Z(n3798) );
  XOR U4921 ( .A(x[120]), .B(x[126]), .Z(n3796) );
  XNOR U4922 ( .A(n3798), .B(n3796), .Z(n3795) );
  XNOR U4923 ( .A(x[122]), .B(n3795), .Z(n3866) );
  IV U4924 ( .A(n3866), .Z(n3800) );
  XNOR U4925 ( .A(x[120]), .B(n3800), .Z(n3848) );
  XNOR U4926 ( .A(x[124]), .B(x[127]), .Z(n3797) );
  IV U4927 ( .A(n3797), .Z(n3861) );
  AND U4928 ( .A(n3848), .B(n3861), .Z(n3805) );
  XOR U4929 ( .A(x[127]), .B(x[122]), .Z(n3888) );
  XNOR U4930 ( .A(n3796), .B(x[125]), .Z(n3811) );
  IV U4931 ( .A(n3811), .Z(n3857) );
  XOR U4932 ( .A(n3798), .B(n3797), .Z(n3822) );
  IV U4933 ( .A(n3822), .Z(n3837) );
  XNOR U4934 ( .A(n3837), .B(x[120]), .Z(n3838) );
  XNOR U4935 ( .A(n3857), .B(n3838), .Z(n3850) );
  NAND U4936 ( .A(n3888), .B(n3850), .Z(n3799) );
  XNOR U4937 ( .A(n3805), .B(n3799), .Z(n3818) );
  XOR U4938 ( .A(x[121]), .B(x[127]), .Z(n3856) );
  XOR U4939 ( .A(n3800), .B(n3857), .Z(n3846) );
  ANDN U4940 ( .B(n3856), .A(n3846), .Z(n3807) );
  XOR U4941 ( .A(x[127]), .B(n3857), .Z(n3899) );
  IV U4942 ( .A(n3899), .Z(n3810) );
  NAND U4943 ( .A(n3800), .B(n3810), .Z(n3801) );
  XOR U4944 ( .A(n3807), .B(n3801), .Z(n3802) );
  XNOR U4945 ( .A(n3818), .B(n3802), .Z(n3842) );
  NANDN U4946 ( .A(x[121]), .B(n3811), .Z(n3809) );
  XNOR U4947 ( .A(n3837), .B(n3846), .Z(n3881) );
  XOR U4948 ( .A(x[124]), .B(x[122]), .Z(n3864) );
  AND U4949 ( .A(n3881), .B(n3864), .Z(n3804) );
  XNOR U4950 ( .A(n3866), .B(n3899), .Z(n3803) );
  XNOR U4951 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U4952 ( .A(n3806), .B(n3805), .Z(n3826) );
  XNOR U4953 ( .A(n3807), .B(n3826), .Z(n3808) );
  XNOR U4954 ( .A(n3809), .B(n3808), .Z(n3840) );
  IV U4955 ( .A(n3840), .Z(n3843) );
  NAND U4956 ( .A(n3842), .B(n3843), .Z(n3836) );
  NANDN U4957 ( .A(n3842), .B(n3843), .Z(n3830) );
  XNOR U4958 ( .A(x[122]), .B(n3810), .Z(n3817) );
  XNOR U4959 ( .A(x[121]), .B(n3817), .Z(n3821) );
  IV U4960 ( .A(n3821), .Z(n3875) );
  XNOR U4961 ( .A(x[124]), .B(n3811), .Z(n3887) );
  OR U4962 ( .A(x[120]), .B(n3887), .Z(n3812) );
  XNOR U4963 ( .A(n3875), .B(n3812), .Z(n3813) );
  NANDN U4964 ( .A(n3822), .B(n3813), .Z(n3816) );
  ANDN U4965 ( .B(x[120]), .A(n3887), .Z(n3814) );
  NAND U4966 ( .A(n3822), .B(n3814), .Z(n3815) );
  NAND U4967 ( .A(n3816), .B(n3815), .Z(n3820) );
  XNOR U4968 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U4969 ( .A(n3820), .B(n3819), .Z(n3844) );
  IV U4970 ( .A(n3842), .Z(n3841) );
  ANDN U4971 ( .B(n3844), .A(n3841), .Z(n3827) );
  AND U4972 ( .A(x[120]), .B(n3821), .Z(n3824) );
  NAND U4973 ( .A(n3822), .B(n3887), .Z(n3823) );
  XNOR U4974 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U4975 ( .A(n3826), .B(n3825), .Z(n3845) );
  XNOR U4976 ( .A(n3827), .B(n3845), .Z(n3828) );
  NAND U4977 ( .A(n3840), .B(n3828), .Z(n3829) );
  NAND U4978 ( .A(n3830), .B(n3829), .Z(n3874) );
  IV U4979 ( .A(n3874), .Z(n3849) );
  OR U4980 ( .A(n3844), .B(n3840), .Z(n3831) );
  NAND U4981 ( .A(n3841), .B(n3831), .Z(n3834) );
  XOR U4982 ( .A(n3844), .B(n3845), .Z(n3832) );
  NANDN U4983 ( .A(n3843), .B(n3832), .Z(n3833) );
  NAND U4984 ( .A(n3834), .B(n3833), .Z(n3886) );
  NANDN U4985 ( .A(n3849), .B(n3886), .Z(n3835) );
  AND U4986 ( .A(n3836), .B(n3835), .Z(n3877) );
  AND U4987 ( .A(n3877), .B(n3837), .Z(n3852) );
  OR U4988 ( .A(n3838), .B(n3849), .Z(n3839) );
  XNOR U4989 ( .A(n3852), .B(n3839), .Z(n3885) );
  XOR U4990 ( .A(n3900), .B(n3859), .Z(n3855) );
  ANDN U4991 ( .B(n3855), .A(n3846), .Z(n3867) );
  NAND U4992 ( .A(n3857), .B(n3859), .Z(n3847) );
  XNOR U4993 ( .A(n3867), .B(n3847), .Z(n3892) );
  XNOR U4994 ( .A(n3885), .B(n3892), .Z(z[122]) );
  AND U4995 ( .A(x[120]), .B(n3886), .Z(n3854) );
  AND U4996 ( .A(n3848), .B(n3863), .Z(n3884) );
  XOR U4997 ( .A(n3849), .B(n3859), .Z(n3862) );
  IV U4998 ( .A(n3862), .Z(n3889) );
  NAND U4999 ( .A(n3889), .B(n3850), .Z(n3851) );
  XNOR U5000 ( .A(n3884), .B(n3851), .Z(n3868) );
  XNOR U5001 ( .A(n3852), .B(n3868), .Z(n3853) );
  XNOR U5002 ( .A(n3854), .B(n3853), .Z(n3928) );
  AND U5003 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U5004 ( .A(x[121]), .B(n3857), .Z(n3858) );
  NAND U5005 ( .A(n3859), .B(n3858), .Z(n3860) );
  XNOR U5006 ( .A(n3901), .B(n3860), .Z(n3872) );
  AND U5007 ( .A(n3863), .B(n3861), .Z(n3891) );
  XNOR U5008 ( .A(n3863), .B(n3862), .Z(n3882) );
  NAND U5009 ( .A(n3882), .B(n3864), .Z(n3865) );
  XNOR U5010 ( .A(n3891), .B(n3865), .Z(n3878) );
  AND U5011 ( .A(n3900), .B(n3866), .Z(n3870) );
  XNOR U5012 ( .A(n3868), .B(n3867), .Z(n3869) );
  XNOR U5013 ( .A(n3870), .B(n3869), .Z(n3927) );
  XNOR U5014 ( .A(n3878), .B(n3927), .Z(n3871) );
  XNOR U5015 ( .A(n3872), .B(n3871), .Z(n3873) );
  XNOR U5016 ( .A(n3928), .B(n3873), .Z(z[125]) );
  AND U5017 ( .A(n3875), .B(n3874), .Z(n3880) );
  XOR U5018 ( .A(n3875), .B(n3887), .Z(n3876) );
  AND U5019 ( .A(n3877), .B(n3876), .Z(n3896) );
  XNOR U5020 ( .A(n3878), .B(n3896), .Z(n3879) );
  XNOR U5021 ( .A(n3880), .B(n3879), .Z(n3907) );
  NAND U5022 ( .A(n3882), .B(n3881), .Z(n3883) );
  XNOR U5023 ( .A(n3884), .B(n3883), .Z(n3895) );
  XNOR U5024 ( .A(n3885), .B(n3895), .Z(n3926) );
  XNOR U5025 ( .A(n3907), .B(n3926), .Z(n3905) );
  AND U5026 ( .A(n3887), .B(n3886), .Z(n3894) );
  NAND U5027 ( .A(n3889), .B(n3888), .Z(n3890) );
  XNOR U5028 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U5029 ( .A(n3902), .B(n3892), .Z(n3893) );
  XNOR U5030 ( .A(n3894), .B(n3893), .Z(n3898) );
  XNOR U5031 ( .A(n3896), .B(n3895), .Z(n3897) );
  XNOR U5032 ( .A(n3898), .B(n3897), .Z(n3906) );
  XNOR U5033 ( .A(n3905), .B(n3906), .Z(z[121]) );
  AND U5034 ( .A(n3900), .B(n3899), .Z(n3904) );
  XNOR U5035 ( .A(n3902), .B(n3901), .Z(n3903) );
  XNOR U5036 ( .A(n3904), .B(n3903), .Z(n3909) );
  XNOR U5037 ( .A(n3905), .B(n3909), .Z(z[126]) );
  XOR U5038 ( .A(n3907), .B(n3906), .Z(n3908) );
  XNOR U5039 ( .A(n3909), .B(n3908), .Z(z[123]) );
  XOR U5040 ( .A(n3943), .B(n3910), .Z(z[0]) );
  AND U5041 ( .A(n3912), .B(n3911), .Z(n3918) );
  XNOR U5042 ( .A(n3916), .B(n3913), .Z(n3914) );
  XNOR U5043 ( .A(n3918), .B(n3914), .Z(n3965) );
  XOR U5044 ( .A(n3965), .B(z[98]), .Z(z[100]) );
  XNOR U5045 ( .A(n3916), .B(n3915), .Z(n3917) );
  XNOR U5046 ( .A(n3918), .B(n3917), .Z(n3919) );
  XOR U5047 ( .A(n3919), .B(z[97]), .Z(z[103]) );
  XOR U5048 ( .A(n3921), .B(n3920), .Z(z[104]) );
  XOR U5049 ( .A(n3921), .B(z[106]), .Z(z[108]) );
  XOR U5050 ( .A(n3922), .B(z[105]), .Z(z[111]) );
  XOR U5051 ( .A(n3924), .B(n3923), .Z(z[112]) );
  XOR U5052 ( .A(n3924), .B(z[114]), .Z(z[116]) );
  XOR U5053 ( .A(n3925), .B(z[113]), .Z(z[119]) );
  XOR U5054 ( .A(n3927), .B(n3926), .Z(z[120]) );
  XOR U5055 ( .A(n3927), .B(z[122]), .Z(z[124]) );
  XOR U5056 ( .A(n3928), .B(z[121]), .Z(z[127]) );
  XOR U5057 ( .A(n3961), .B(z[10]), .Z(z[12]) );
  XOR U5058 ( .A(n3929), .B(z[9]), .Z(z[15]) );
  XOR U5059 ( .A(n3931), .B(n3930), .Z(z[16]) );
  XOR U5060 ( .A(n3931), .B(z[18]), .Z(z[20]) );
  XOR U5061 ( .A(n3932), .B(z[17]), .Z(z[23]) );
  XOR U5062 ( .A(n3934), .B(n3933), .Z(z[24]) );
  XOR U5063 ( .A(n3934), .B(z[26]), .Z(z[28]) );
  XOR U5064 ( .A(n3935), .B(z[25]), .Z(z[31]) );
  XOR U5065 ( .A(n3937), .B(n3936), .Z(z[32]) );
  XOR U5066 ( .A(n3937), .B(z[34]), .Z(z[36]) );
  XOR U5067 ( .A(n3938), .B(z[33]), .Z(z[39]) );
  XOR U5068 ( .A(n3940), .B(n3939), .Z(z[40]) );
  XOR U5069 ( .A(n3940), .B(z[42]), .Z(z[44]) );
  XOR U5070 ( .A(n3941), .B(z[41]), .Z(z[47]) );
  XOR U5071 ( .A(n3944), .B(n3942), .Z(z[48]) );
  XOR U5072 ( .A(n3943), .B(z[2]), .Z(z[4]) );
  XOR U5073 ( .A(n3944), .B(z[50]), .Z(z[52]) );
  XOR U5074 ( .A(n3945), .B(z[49]), .Z(z[55]) );
  XOR U5075 ( .A(n3947), .B(n3946), .Z(z[56]) );
  XOR U5076 ( .A(n3947), .B(z[58]), .Z(z[60]) );
  XOR U5077 ( .A(n3948), .B(z[57]), .Z(z[63]) );
  XOR U5078 ( .A(n3950), .B(n3949), .Z(z[64]) );
  XOR U5079 ( .A(n3950), .B(z[66]), .Z(z[68]) );
  XOR U5080 ( .A(n3951), .B(z[65]), .Z(z[71]) );
  XOR U5081 ( .A(n3953), .B(n3952), .Z(z[72]) );
  XOR U5082 ( .A(n3953), .B(z[74]), .Z(z[76]) );
  XOR U5083 ( .A(n3954), .B(z[73]), .Z(z[79]) );
  XOR U5084 ( .A(n3955), .B(z[1]), .Z(z[7]) );
  XOR U5085 ( .A(n3957), .B(n3956), .Z(z[80]) );
  XOR U5086 ( .A(n3957), .B(z[82]), .Z(z[84]) );
  XOR U5087 ( .A(n3958), .B(z[81]), .Z(z[87]) );
  XOR U5088 ( .A(n3962), .B(n3959), .Z(z[88]) );
  XOR U5089 ( .A(n3961), .B(n3960), .Z(z[8]) );
  XOR U5090 ( .A(n3962), .B(z[90]), .Z(z[92]) );
  XOR U5091 ( .A(n3963), .B(z[89]), .Z(z[95]) );
  XOR U5092 ( .A(n3965), .B(n3964), .Z(z[96]) );
endmodule


module aes_comb ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [1279:0] key;
  output [127:0] out;
  input clk, rst;
  wire   \w1[9][127] , \w1[9][126] , \w1[9][125] , \w1[9][124] , \w1[9][123] ,
         \w1[9][122] , \w1[9][121] , \w1[9][120] , \w1[9][119] , \w1[9][118] ,
         \w1[9][117] , \w1[9][116] , \w1[9][115] , \w1[9][114] , \w1[9][113] ,
         \w1[9][112] , \w1[9][111] , \w1[9][110] , \w1[9][109] , \w1[9][108] ,
         \w1[9][107] , \w1[9][106] , \w1[9][105] , \w1[9][104] , \w1[9][103] ,
         \w1[9][102] , \w1[9][101] , \w1[9][100] , \w1[9][99] , \w1[9][98] ,
         \w1[9][97] , \w1[9][96] , \w1[9][95] , \w1[9][94] , \w1[9][93] ,
         \w1[9][92] , \w1[9][91] , \w1[9][90] , \w1[9][89] , \w1[9][88] ,
         \w1[9][87] , \w1[9][86] , \w1[9][85] , \w1[9][84] , \w1[9][83] ,
         \w1[9][82] , \w1[9][81] , \w1[9][80] , \w1[9][79] , \w1[9][78] ,
         \w1[9][77] , \w1[9][76] , \w1[9][75] , \w1[9][74] , \w1[9][73] ,
         \w1[9][72] , \w1[9][71] , \w1[9][70] , \w1[9][69] , \w1[9][68] ,
         \w1[9][67] , \w1[9][66] , \w1[9][65] , \w1[9][64] , \w1[9][63] ,
         \w1[9][62] , \w1[9][61] , \w1[9][60] , \w1[9][59] , \w1[9][58] ,
         \w1[9][57] , \w1[9][56] , \w1[9][55] , \w1[9][54] , \w1[9][53] ,
         \w1[9][52] , \w1[9][51] , \w1[9][50] , \w1[9][49] , \w1[9][48] ,
         \w1[9][47] , \w1[9][46] , \w1[9][45] , \w1[9][44] , \w1[9][43] ,
         \w1[9][42] , \w1[9][41] , \w1[9][40] , \w1[9][39] , \w1[9][38] ,
         \w1[9][37] , \w1[9][36] , \w1[9][35] , \w1[9][34] , \w1[9][33] ,
         \w1[9][32] , \w1[9][31] , \w1[9][30] , \w1[9][29] , \w1[9][28] ,
         \w1[9][27] , \w1[9][26] , \w1[9][25] , \w1[9][24] , \w1[9][23] ,
         \w1[9][22] , \w1[9][21] , \w1[9][20] , \w1[9][19] , \w1[9][18] ,
         \w1[9][17] , \w1[9][16] , \w1[9][15] , \w1[9][14] , \w1[9][13] ,
         \w1[9][12] , \w1[9][11] , \w1[9][10] , \w1[9][9] , \w1[9][8] ,
         \w1[9][7] , \w1[9][6] , \w1[9][5] , \w1[9][4] , \w1[9][3] ,
         \w1[9][2] , \w1[9][1] , \w1[9][0] , \w1[8][127] , \w1[8][126] ,
         \w1[8][125] , \w1[8][124] , \w1[8][123] , \w1[8][122] , \w1[8][121] ,
         \w1[8][120] , \w1[8][119] , \w1[8][118] , \w1[8][117] , \w1[8][116] ,
         \w1[8][115] , \w1[8][114] , \w1[8][113] , \w1[8][112] , \w1[8][111] ,
         \w1[8][110] , \w1[8][109] , \w1[8][108] , \w1[8][107] , \w1[8][106] ,
         \w1[8][105] , \w1[8][104] , \w1[8][103] , \w1[8][102] , \w1[8][101] ,
         \w1[8][100] , \w1[8][99] , \w1[8][98] , \w1[8][97] , \w1[8][96] ,
         \w1[8][95] , \w1[8][94] , \w1[8][93] , \w1[8][92] , \w1[8][91] ,
         \w1[8][90] , \w1[8][89] , \w1[8][88] , \w1[8][87] , \w1[8][86] ,
         \w1[8][85] , \w1[8][84] , \w1[8][83] , \w1[8][82] , \w1[8][81] ,
         \w1[8][80] , \w1[8][79] , \w1[8][78] , \w1[8][77] , \w1[8][76] ,
         \w1[8][75] , \w1[8][74] , \w1[8][73] , \w1[8][72] , \w1[8][71] ,
         \w1[8][70] , \w1[8][69] , \w1[8][68] , \w1[8][67] , \w1[8][66] ,
         \w1[8][65] , \w1[8][64] , \w1[8][63] , \w1[8][62] , \w1[8][61] ,
         \w1[8][60] , \w1[8][59] , \w1[8][58] , \w1[8][57] , \w1[8][56] ,
         \w1[8][55] , \w1[8][54] , \w1[8][53] , \w1[8][52] , \w1[8][51] ,
         \w1[8][50] , \w1[8][49] , \w1[8][48] , \w1[8][47] , \w1[8][46] ,
         \w1[8][45] , \w1[8][44] , \w1[8][43] , \w1[8][42] , \w1[8][41] ,
         \w1[8][40] , \w1[8][39] , \w1[8][38] , \w1[8][37] , \w1[8][36] ,
         \w1[8][35] , \w1[8][34] , \w1[8][33] , \w1[8][32] , \w1[8][31] ,
         \w1[8][30] , \w1[8][29] , \w1[8][28] , \w1[8][27] , \w1[8][26] ,
         \w1[8][25] , \w1[8][24] , \w1[8][23] , \w1[8][22] , \w1[8][21] ,
         \w1[8][20] , \w1[8][19] , \w1[8][18] , \w1[8][17] , \w1[8][16] ,
         \w1[8][15] , \w1[8][14] , \w1[8][13] , \w1[8][12] , \w1[8][11] ,
         \w1[8][10] , \w1[8][9] , \w1[8][8] , \w1[8][7] , \w1[8][6] ,
         \w1[8][5] , \w1[8][4] , \w1[8][3] , \w1[8][2] , \w1[8][1] ,
         \w1[8][0] , \w1[7][127] , \w1[7][126] , \w1[7][125] , \w1[7][124] ,
         \w1[7][123] , \w1[7][122] , \w1[7][121] , \w1[7][120] , \w1[7][119] ,
         \w1[7][118] , \w1[7][117] , \w1[7][116] , \w1[7][115] , \w1[7][114] ,
         \w1[7][113] , \w1[7][112] , \w1[7][111] , \w1[7][110] , \w1[7][109] ,
         \w1[7][108] , \w1[7][107] , \w1[7][106] , \w1[7][105] , \w1[7][104] ,
         \w1[7][103] , \w1[7][102] , \w1[7][101] , \w1[7][100] , \w1[7][99] ,
         \w1[7][98] , \w1[7][97] , \w1[7][96] , \w1[7][95] , \w1[7][94] ,
         \w1[7][93] , \w1[7][92] , \w1[7][91] , \w1[7][90] , \w1[7][89] ,
         \w1[7][88] , \w1[7][87] , \w1[7][86] , \w1[7][85] , \w1[7][84] ,
         \w1[7][83] , \w1[7][82] , \w1[7][81] , \w1[7][80] , \w1[7][79] ,
         \w1[7][78] , \w1[7][77] , \w1[7][76] , \w1[7][75] , \w1[7][74] ,
         \w1[7][73] , \w1[7][72] , \w1[7][71] , \w1[7][70] , \w1[7][69] ,
         \w1[7][68] , \w1[7][67] , \w1[7][66] , \w1[7][65] , \w1[7][64] ,
         \w1[7][63] , \w1[7][62] , \w1[7][61] , \w1[7][60] , \w1[7][59] ,
         \w1[7][58] , \w1[7][57] , \w1[7][56] , \w1[7][55] , \w1[7][54] ,
         \w1[7][53] , \w1[7][52] , \w1[7][51] , \w1[7][50] , \w1[7][49] ,
         \w1[7][48] , \w1[7][47] , \w1[7][46] , \w1[7][45] , \w1[7][44] ,
         \w1[7][43] , \w1[7][42] , \w1[7][41] , \w1[7][40] , \w1[7][39] ,
         \w1[7][38] , \w1[7][37] , \w1[7][36] , \w1[7][35] , \w1[7][34] ,
         \w1[7][33] , \w1[7][32] , \w1[7][31] , \w1[7][30] , \w1[7][29] ,
         \w1[7][28] , \w1[7][27] , \w1[7][26] , \w1[7][25] , \w1[7][24] ,
         \w1[7][23] , \w1[7][22] , \w1[7][21] , \w1[7][20] , \w1[7][19] ,
         \w1[7][18] , \w1[7][17] , \w1[7][16] , \w1[7][15] , \w1[7][14] ,
         \w1[7][13] , \w1[7][12] , \w1[7][11] , \w1[7][10] , \w1[7][9] ,
         \w1[7][8] , \w1[7][7] , \w1[7][6] , \w1[7][5] , \w1[7][4] ,
         \w1[7][3] , \w1[7][2] , \w1[7][1] , \w1[7][0] , \w1[6][127] ,
         \w1[6][126] , \w1[6][125] , \w1[6][124] , \w1[6][123] , \w1[6][122] ,
         \w1[6][121] , \w1[6][120] , \w1[6][119] , \w1[6][118] , \w1[6][117] ,
         \w1[6][116] , \w1[6][115] , \w1[6][114] , \w1[6][113] , \w1[6][112] ,
         \w1[6][111] , \w1[6][110] , \w1[6][109] , \w1[6][108] , \w1[6][107] ,
         \w1[6][106] , \w1[6][105] , \w1[6][104] , \w1[6][103] , \w1[6][102] ,
         \w1[6][101] , \w1[6][100] , \w1[6][99] , \w1[6][98] , \w1[6][97] ,
         \w1[6][96] , \w1[6][95] , \w1[6][94] , \w1[6][93] , \w1[6][92] ,
         \w1[6][91] , \w1[6][90] , \w1[6][89] , \w1[6][88] , \w1[6][87] ,
         \w1[6][86] , \w1[6][85] , \w1[6][84] , \w1[6][83] , \w1[6][82] ,
         \w1[6][81] , \w1[6][80] , \w1[6][79] , \w1[6][78] , \w1[6][77] ,
         \w1[6][76] , \w1[6][75] , \w1[6][74] , \w1[6][73] , \w1[6][72] ,
         \w1[6][71] , \w1[6][70] , \w1[6][69] , \w1[6][68] , \w1[6][67] ,
         \w1[6][66] , \w1[6][65] , \w1[6][64] , \w1[6][63] , \w1[6][62] ,
         \w1[6][61] , \w1[6][60] , \w1[6][59] , \w1[6][58] , \w1[6][57] ,
         \w1[6][56] , \w1[6][55] , \w1[6][54] , \w1[6][53] , \w1[6][52] ,
         \w1[6][51] , \w1[6][50] , \w1[6][49] , \w1[6][48] , \w1[6][47] ,
         \w1[6][46] , \w1[6][45] , \w1[6][44] , \w1[6][43] , \w1[6][42] ,
         \w1[6][41] , \w1[6][40] , \w1[6][39] , \w1[6][38] , \w1[6][37] ,
         \w1[6][36] , \w1[6][35] , \w1[6][34] , \w1[6][33] , \w1[6][32] ,
         \w1[6][31] , \w1[6][30] , \w1[6][29] , \w1[6][28] , \w1[6][27] ,
         \w1[6][26] , \w1[6][25] , \w1[6][24] , \w1[6][23] , \w1[6][22] ,
         \w1[6][21] , \w1[6][20] , \w1[6][19] , \w1[6][18] , \w1[6][17] ,
         \w1[6][16] , \w1[6][15] , \w1[6][14] , \w1[6][13] , \w1[6][12] ,
         \w1[6][11] , \w1[6][10] , \w1[6][9] , \w1[6][8] , \w1[6][7] ,
         \w1[6][6] , \w1[6][5] , \w1[6][4] , \w1[6][3] , \w1[6][2] ,
         \w1[6][1] , \w1[6][0] , \w1[5][127] , \w1[5][126] , \w1[5][125] ,
         \w1[5][124] , \w1[5][123] , \w1[5][122] , \w1[5][121] , \w1[5][120] ,
         \w1[5][119] , \w1[5][118] , \w1[5][117] , \w1[5][116] , \w1[5][115] ,
         \w1[5][114] , \w1[5][113] , \w1[5][112] , \w1[5][111] , \w1[5][110] ,
         \w1[5][109] , \w1[5][108] , \w1[5][107] , \w1[5][106] , \w1[5][105] ,
         \w1[5][104] , \w1[5][103] , \w1[5][102] , \w1[5][101] , \w1[5][100] ,
         \w1[5][99] , \w1[5][98] , \w1[5][97] , \w1[5][96] , \w1[5][95] ,
         \w1[5][94] , \w1[5][93] , \w1[5][92] , \w1[5][91] , \w1[5][90] ,
         \w1[5][89] , \w1[5][88] , \w1[5][87] , \w1[5][86] , \w1[5][85] ,
         \w1[5][84] , \w1[5][83] , \w1[5][82] , \w1[5][81] , \w1[5][80] ,
         \w1[5][79] , \w1[5][78] , \w1[5][77] , \w1[5][76] , \w1[5][75] ,
         \w1[5][74] , \w1[5][73] , \w1[5][72] , \w1[5][71] , \w1[5][70] ,
         \w1[5][69] , \w1[5][68] , \w1[5][67] , \w1[5][66] , \w1[5][65] ,
         \w1[5][64] , \w1[5][63] , \w1[5][62] , \w1[5][61] , \w1[5][60] ,
         \w1[5][59] , \w1[5][58] , \w1[5][57] , \w1[5][56] , \w1[5][55] ,
         \w1[5][54] , \w1[5][53] , \w1[5][52] , \w1[5][51] , \w1[5][50] ,
         \w1[5][49] , \w1[5][48] , \w1[5][47] , \w1[5][46] , \w1[5][45] ,
         \w1[5][44] , \w1[5][43] , \w1[5][42] , \w1[5][41] , \w1[5][40] ,
         \w1[5][39] , \w1[5][38] , \w1[5][37] , \w1[5][36] , \w1[5][35] ,
         \w1[5][34] , \w1[5][33] , \w1[5][32] , \w1[5][31] , \w1[5][30] ,
         \w1[5][29] , \w1[5][28] , \w1[5][27] , \w1[5][26] , \w1[5][25] ,
         \w1[5][24] , \w1[5][23] , \w1[5][22] , \w1[5][21] , \w1[5][20] ,
         \w1[5][19] , \w1[5][18] , \w1[5][17] , \w1[5][16] , \w1[5][15] ,
         \w1[5][14] , \w1[5][13] , \w1[5][12] , \w1[5][11] , \w1[5][10] ,
         \w1[5][9] , \w1[5][8] , \w1[5][7] , \w1[5][6] , \w1[5][5] ,
         \w1[5][4] , \w1[5][3] , \w1[5][2] , \w1[5][1] , \w1[5][0] ,
         \w1[4][127] , \w1[4][126] , \w1[4][125] , \w1[4][124] , \w1[4][123] ,
         \w1[4][122] , \w1[4][121] , \w1[4][120] , \w1[4][119] , \w1[4][118] ,
         \w1[4][117] , \w1[4][116] , \w1[4][115] , \w1[4][114] , \w1[4][113] ,
         \w1[4][112] , \w1[4][111] , \w1[4][110] , \w1[4][109] , \w1[4][108] ,
         \w1[4][107] , \w1[4][106] , \w1[4][105] , \w1[4][104] , \w1[4][103] ,
         \w1[4][102] , \w1[4][101] , \w1[4][100] , \w1[4][99] , \w1[4][98] ,
         \w1[4][97] , \w1[4][96] , \w1[4][95] , \w1[4][94] , \w1[4][93] ,
         \w1[4][92] , \w1[4][91] , \w1[4][90] , \w1[4][89] , \w1[4][88] ,
         \w1[4][87] , \w1[4][86] , \w1[4][85] , \w1[4][84] , \w1[4][83] ,
         \w1[4][82] , \w1[4][81] , \w1[4][80] , \w1[4][79] , \w1[4][78] ,
         \w1[4][77] , \w1[4][76] , \w1[4][75] , \w1[4][74] , \w1[4][73] ,
         \w1[4][72] , \w1[4][71] , \w1[4][70] , \w1[4][69] , \w1[4][68] ,
         \w1[4][67] , \w1[4][66] , \w1[4][65] , \w1[4][64] , \w1[4][63] ,
         \w1[4][62] , \w1[4][61] , \w1[4][60] , \w1[4][59] , \w1[4][58] ,
         \w1[4][57] , \w1[4][56] , \w1[4][55] , \w1[4][54] , \w1[4][53] ,
         \w1[4][52] , \w1[4][51] , \w1[4][50] , \w1[4][49] , \w1[4][48] ,
         \w1[4][47] , \w1[4][46] , \w1[4][45] , \w1[4][44] , \w1[4][43] ,
         \w1[4][42] , \w1[4][41] , \w1[4][40] , \w1[4][39] , \w1[4][38] ,
         \w1[4][37] , \w1[4][36] , \w1[4][35] , \w1[4][34] , \w1[4][33] ,
         \w1[4][32] , \w1[4][31] , \w1[4][30] , \w1[4][29] , \w1[4][28] ,
         \w1[4][27] , \w1[4][26] , \w1[4][25] , \w1[4][24] , \w1[4][23] ,
         \w1[4][22] , \w1[4][21] , \w1[4][20] , \w1[4][19] , \w1[4][18] ,
         \w1[4][17] , \w1[4][16] , \w1[4][15] , \w1[4][14] , \w1[4][13] ,
         \w1[4][12] , \w1[4][11] , \w1[4][10] , \w1[4][9] , \w1[4][8] ,
         \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , \w1[4][3] ,
         \w1[4][2] , \w1[4][1] , \w1[4][0] , \w1[3][127] , \w1[3][126] ,
         \w1[3][125] , \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] ,
         \w1[3][120] , \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] ,
         \w1[3][115] , \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] ,
         \w1[3][110] , \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] ,
         \w1[3][105] , \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] ,
         \w1[3][100] , \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] ,
         \w1[3][95] , \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] ,
         \w1[3][90] , \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] ,
         \w1[3][85] , \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] ,
         \w1[3][80] , \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] ,
         \w1[3][75] , \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] ,
         \w1[3][70] , \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] ,
         \w1[3][65] , \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] ,
         \w1[3][60] , \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] ,
         \w1[3][55] , \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] ,
         \w1[3][50] , \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] ,
         \w1[3][45] , \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] ,
         \w1[3][40] , \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] ,
         \w1[3][35] , \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] ,
         \w1[3][30] , \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] ,
         \w1[3][25] , \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] ,
         \w1[3][20] , \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] ,
         \w1[3][15] , \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] ,
         \w1[3][10] , \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] ,
         \w1[3][5] , \w1[3][4] , \w1[3][3] , \w1[3][2] , \w1[3][1] ,
         \w1[3][0] , \w1[2][127] , \w1[2][126] , \w1[2][125] , \w1[2][124] ,
         \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , \w1[2][119] ,
         \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , \w1[2][114] ,
         \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , \w1[2][109] ,
         \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , \w1[2][104] ,
         \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , \w1[2][99] ,
         \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , \w1[2][94] ,
         \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , \w1[2][89] ,
         \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , \w1[2][84] ,
         \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , \w1[2][79] ,
         \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , \w1[2][74] ,
         \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , \w1[2][69] ,
         \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , \w1[2][64] ,
         \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , \w1[2][59] ,
         \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , \w1[2][54] ,
         \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , \w1[2][49] ,
         \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , \w1[2][44] ,
         \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , \w1[2][39] ,
         \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , \w1[2][34] ,
         \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , \w1[2][29] ,
         \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , \w1[2][24] ,
         \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , \w1[2][19] ,
         \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , \w1[2][14] ,
         \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , \w1[2][9] ,
         \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] ,
         \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] , \w1[1][127] ,
         \w1[1][126] , \w1[1][125] , \w1[1][124] , \w1[1][123] , \w1[1][122] ,
         \w1[1][121] , \w1[1][120] , \w1[1][119] , \w1[1][118] , \w1[1][117] ,
         \w1[1][116] , \w1[1][115] , \w1[1][114] , \w1[1][113] , \w1[1][112] ,
         \w1[1][111] , \w1[1][110] , \w1[1][109] , \w1[1][108] , \w1[1][107] ,
         \w1[1][106] , \w1[1][105] , \w1[1][104] , \w1[1][103] , \w1[1][102] ,
         \w1[1][101] , \w1[1][100] , \w1[1][99] , \w1[1][98] , \w1[1][97] ,
         \w1[1][96] , \w1[1][95] , \w1[1][94] , \w1[1][93] , \w1[1][92] ,
         \w1[1][91] , \w1[1][90] , \w1[1][89] , \w1[1][88] , \w1[1][87] ,
         \w1[1][86] , \w1[1][85] , \w1[1][84] , \w1[1][83] , \w1[1][82] ,
         \w1[1][81] , \w1[1][80] , \w1[1][79] , \w1[1][78] , \w1[1][77] ,
         \w1[1][76] , \w1[1][75] , \w1[1][74] , \w1[1][73] , \w1[1][72] ,
         \w1[1][71] , \w1[1][70] , \w1[1][69] , \w1[1][68] , \w1[1][67] ,
         \w1[1][66] , \w1[1][65] , \w1[1][64] , \w1[1][63] , \w1[1][62] ,
         \w1[1][61] , \w1[1][60] , \w1[1][59] , \w1[1][58] , \w1[1][57] ,
         \w1[1][56] , \w1[1][55] , \w1[1][54] , \w1[1][53] , \w1[1][52] ,
         \w1[1][51] , \w1[1][50] , \w1[1][49] , \w1[1][48] , \w1[1][47] ,
         \w1[1][46] , \w1[1][45] , \w1[1][44] , \w1[1][43] , \w1[1][42] ,
         \w1[1][41] , \w1[1][40] , \w1[1][39] , \w1[1][38] , \w1[1][37] ,
         \w1[1][36] , \w1[1][35] , \w1[1][34] , \w1[1][33] , \w1[1][32] ,
         \w1[1][31] , \w1[1][30] , \w1[1][29] , \w1[1][28] , \w1[1][27] ,
         \w1[1][26] , \w1[1][25] , \w1[1][24] , \w1[1][23] , \w1[1][22] ,
         \w1[1][21] , \w1[1][20] , \w1[1][19] , \w1[1][18] , \w1[1][17] ,
         \w1[1][16] , \w1[1][15] , \w1[1][14] , \w1[1][13] , \w1[1][12] ,
         \w1[1][11] , \w1[1][10] , \w1[1][9] , \w1[1][8] , \w1[1][7] ,
         \w1[1][6] , \w1[1][5] , \w1[1][4] , \w1[1][3] , \w1[1][2] ,
         \w1[1][1] , \w1[1][0] , \w1[0][127] , \w1[0][126] , \w1[0][125] ,
         \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] ,
         \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] ,
         \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] ,
         \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] ,
         \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] ,
         \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] ,
         \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] ,
         \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] ,
         \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] ,
         \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] ,
         \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] ,
         \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] ,
         \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] ,
         \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] ,
         \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] ,
         \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] ,
         \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] ,
         \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] ,
         \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] ,
         \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] ,
         \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] ,
         \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] ,
         \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] ,
         \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] ,
         \w1[0][4] , \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] ,
         \w3[9][127] , \w3[9][126] , \w3[9][125] , \w3[9][124] , \w3[9][123] ,
         \w3[9][122] , \w3[9][121] , \w3[9][120] , \w3[9][119] , \w3[9][118] ,
         \w3[9][117] , \w3[9][116] , \w3[9][115] , \w3[9][114] , \w3[9][113] ,
         \w3[9][112] , \w3[9][111] , \w3[9][110] , \w3[9][109] , \w3[9][108] ,
         \w3[9][107] , \w3[9][106] , \w3[9][105] , \w3[9][104] , \w3[9][103] ,
         \w3[9][102] , \w3[9][101] , \w3[9][100] , \w3[9][99] , \w3[9][98] ,
         \w3[9][97] , \w3[9][96] , \w3[9][95] , \w3[9][94] , \w3[9][93] ,
         \w3[9][92] , \w3[9][91] , \w3[9][90] , \w3[9][89] , \w3[9][88] ,
         \w3[9][87] , \w3[9][86] , \w3[9][85] , \w3[9][84] , \w3[9][83] ,
         \w3[9][82] , \w3[9][81] , \w3[9][80] , \w3[9][79] , \w3[9][78] ,
         \w3[9][77] , \w3[9][76] , \w3[9][75] , \w3[9][74] , \w3[9][73] ,
         \w3[9][72] , \w3[9][71] , \w3[9][70] , \w3[9][69] , \w3[9][68] ,
         \w3[9][67] , \w3[9][66] , \w3[9][65] , \w3[9][64] , \w3[9][63] ,
         \w3[9][62] , \w3[9][61] , \w3[9][60] , \w3[9][59] , \w3[9][58] ,
         \w3[9][57] , \w3[9][56] , \w3[9][55] , \w3[9][54] , \w3[9][53] ,
         \w3[9][52] , \w3[9][51] , \w3[9][50] , \w3[9][49] , \w3[9][48] ,
         \w3[9][47] , \w3[9][46] , \w3[9][45] , \w3[9][44] , \w3[9][43] ,
         \w3[9][42] , \w3[9][41] , \w3[9][40] , \w3[9][39] , \w3[9][38] ,
         \w3[9][37] , \w3[9][36] , \w3[9][35] , \w3[9][34] , \w3[9][33] ,
         \w3[9][32] , \w3[9][31] , \w3[9][30] , \w3[9][29] , \w3[9][28] ,
         \w3[9][27] , \w3[9][26] , \w3[9][25] , \w3[9][24] , \w3[9][23] ,
         \w3[9][22] , \w3[9][21] , \w3[9][20] , \w3[9][19] , \w3[9][18] ,
         \w3[9][17] , \w3[9][16] , \w3[9][15] , \w3[9][14] , \w3[9][13] ,
         \w3[9][12] , \w3[9][11] , \w3[9][10] , \w3[9][9] , \w3[9][8] ,
         \w3[9][7] , \w3[9][6] , \w3[9][5] , \w3[9][4] , \w3[9][3] ,
         \w3[9][2] , \w3[9][1] , \w3[9][0] , \w3[8][127] , \w3[8][126] ,
         \w3[8][125] , \w3[8][124] , \w3[8][123] , \w3[8][122] , \w3[8][121] ,
         \w3[8][120] , \w3[8][119] , \w3[8][118] , \w3[8][117] , \w3[8][116] ,
         \w3[8][115] , \w3[8][114] , \w3[8][113] , \w3[8][112] , \w3[8][111] ,
         \w3[8][110] , \w3[8][109] , \w3[8][108] , \w3[8][107] , \w3[8][106] ,
         \w3[8][105] , \w3[8][104] , \w3[8][103] , \w3[8][102] , \w3[8][101] ,
         \w3[8][100] , \w3[8][99] , \w3[8][98] , \w3[8][97] , \w3[8][96] ,
         \w3[8][95] , \w3[8][94] , \w3[8][93] , \w3[8][92] , \w3[8][91] ,
         \w3[8][90] , \w3[8][89] , \w3[8][88] , \w3[8][87] , \w3[8][86] ,
         \w3[8][85] , \w3[8][84] , \w3[8][83] , \w3[8][82] , \w3[8][81] ,
         \w3[8][80] , \w3[8][79] , \w3[8][78] , \w3[8][77] , \w3[8][76] ,
         \w3[8][75] , \w3[8][74] , \w3[8][73] , \w3[8][72] , \w3[8][71] ,
         \w3[8][70] , \w3[8][69] , \w3[8][68] , \w3[8][67] , \w3[8][66] ,
         \w3[8][65] , \w3[8][64] , \w3[8][63] , \w3[8][62] , \w3[8][61] ,
         \w3[8][60] , \w3[8][59] , \w3[8][58] , \w3[8][57] , \w3[8][56] ,
         \w3[8][55] , \w3[8][54] , \w3[8][53] , \w3[8][52] , \w3[8][51] ,
         \w3[8][50] , \w3[8][49] , \w3[8][48] , \w3[8][47] , \w3[8][46] ,
         \w3[8][45] , \w3[8][44] , \w3[8][43] , \w3[8][42] , \w3[8][41] ,
         \w3[8][40] , \w3[8][39] , \w3[8][38] , \w3[8][37] , \w3[8][36] ,
         \w3[8][35] , \w3[8][34] , \w3[8][33] , \w3[8][32] , \w3[8][31] ,
         \w3[8][30] , \w3[8][29] , \w3[8][28] , \w3[8][27] , \w3[8][26] ,
         \w3[8][25] , \w3[8][24] , \w3[8][23] , \w3[8][22] , \w3[8][21] ,
         \w3[8][20] , \w3[8][19] , \w3[8][18] , \w3[8][17] , \w3[8][16] ,
         \w3[8][15] , \w3[8][14] , \w3[8][13] , \w3[8][12] , \w3[8][11] ,
         \w3[8][10] , \w3[8][9] , \w3[8][8] , \w3[8][7] , \w3[8][6] ,
         \w3[8][5] , \w3[8][4] , \w3[8][3] , \w3[8][2] , \w3[8][1] ,
         \w3[8][0] , \w3[7][127] , \w3[7][126] , \w3[7][125] , \w3[7][124] ,
         \w3[7][123] , \w3[7][122] , \w3[7][121] , \w3[7][120] , \w3[7][119] ,
         \w3[7][118] , \w3[7][117] , \w3[7][116] , \w3[7][115] , \w3[7][114] ,
         \w3[7][113] , \w3[7][112] , \w3[7][111] , \w3[7][110] , \w3[7][109] ,
         \w3[7][108] , \w3[7][107] , \w3[7][106] , \w3[7][105] , \w3[7][104] ,
         \w3[7][103] , \w3[7][102] , \w3[7][101] , \w3[7][100] , \w3[7][99] ,
         \w3[7][98] , \w3[7][97] , \w3[7][96] , \w3[7][95] , \w3[7][94] ,
         \w3[7][93] , \w3[7][92] , \w3[7][91] , \w3[7][90] , \w3[7][89] ,
         \w3[7][88] , \w3[7][87] , \w3[7][86] , \w3[7][85] , \w3[7][84] ,
         \w3[7][83] , \w3[7][82] , \w3[7][81] , \w3[7][80] , \w3[7][79] ,
         \w3[7][78] , \w3[7][77] , \w3[7][76] , \w3[7][75] , \w3[7][74] ,
         \w3[7][73] , \w3[7][72] , \w3[7][71] , \w3[7][70] , \w3[7][69] ,
         \w3[7][68] , \w3[7][67] , \w3[7][66] , \w3[7][65] , \w3[7][64] ,
         \w3[7][63] , \w3[7][62] , \w3[7][61] , \w3[7][60] , \w3[7][59] ,
         \w3[7][58] , \w3[7][57] , \w3[7][56] , \w3[7][55] , \w3[7][54] ,
         \w3[7][53] , \w3[7][52] , \w3[7][51] , \w3[7][50] , \w3[7][49] ,
         \w3[7][48] , \w3[7][47] , \w3[7][46] , \w3[7][45] , \w3[7][44] ,
         \w3[7][43] , \w3[7][42] , \w3[7][41] , \w3[7][40] , \w3[7][39] ,
         \w3[7][38] , \w3[7][37] , \w3[7][36] , \w3[7][35] , \w3[7][34] ,
         \w3[7][33] , \w3[7][32] , \w3[7][31] , \w3[7][30] , \w3[7][29] ,
         \w3[7][28] , \w3[7][27] , \w3[7][26] , \w3[7][25] , \w3[7][24] ,
         \w3[7][23] , \w3[7][22] , \w3[7][21] , \w3[7][20] , \w3[7][19] ,
         \w3[7][18] , \w3[7][17] , \w3[7][16] , \w3[7][15] , \w3[7][14] ,
         \w3[7][13] , \w3[7][12] , \w3[7][11] , \w3[7][10] , \w3[7][9] ,
         \w3[7][8] , \w3[7][7] , \w3[7][6] , \w3[7][5] , \w3[7][4] ,
         \w3[7][3] , \w3[7][2] , \w3[7][1] , \w3[7][0] , \w3[6][127] ,
         \w3[6][126] , \w3[6][125] , \w3[6][124] , \w3[6][123] , \w3[6][122] ,
         \w3[6][121] , \w3[6][120] , \w3[6][119] , \w3[6][118] , \w3[6][117] ,
         \w3[6][116] , \w3[6][115] , \w3[6][114] , \w3[6][113] , \w3[6][112] ,
         \w3[6][111] , \w3[6][110] , \w3[6][109] , \w3[6][108] , \w3[6][107] ,
         \w3[6][106] , \w3[6][105] , \w3[6][104] , \w3[6][103] , \w3[6][102] ,
         \w3[6][101] , \w3[6][100] , \w3[6][99] , \w3[6][98] , \w3[6][97] ,
         \w3[6][96] , \w3[6][95] , \w3[6][94] , \w3[6][93] , \w3[6][92] ,
         \w3[6][91] , \w3[6][90] , \w3[6][89] , \w3[6][88] , \w3[6][87] ,
         \w3[6][86] , \w3[6][85] , \w3[6][84] , \w3[6][83] , \w3[6][82] ,
         \w3[6][81] , \w3[6][80] , \w3[6][79] , \w3[6][78] , \w3[6][77] ,
         \w3[6][76] , \w3[6][75] , \w3[6][74] , \w3[6][73] , \w3[6][72] ,
         \w3[6][71] , \w3[6][70] , \w3[6][69] , \w3[6][68] , \w3[6][67] ,
         \w3[6][66] , \w3[6][65] , \w3[6][64] , \w3[6][63] , \w3[6][62] ,
         \w3[6][61] , \w3[6][60] , \w3[6][59] , \w3[6][58] , \w3[6][57] ,
         \w3[6][56] , \w3[6][55] , \w3[6][54] , \w3[6][53] , \w3[6][52] ,
         \w3[6][51] , \w3[6][50] , \w3[6][49] , \w3[6][48] , \w3[6][47] ,
         \w3[6][46] , \w3[6][45] , \w3[6][44] , \w3[6][43] , \w3[6][42] ,
         \w3[6][41] , \w3[6][40] , \w3[6][39] , \w3[6][38] , \w3[6][37] ,
         \w3[6][36] , \w3[6][35] , \w3[6][34] , \w3[6][33] , \w3[6][32] ,
         \w3[6][31] , \w3[6][30] , \w3[6][29] , \w3[6][28] , \w3[6][27] ,
         \w3[6][26] , \w3[6][25] , \w3[6][24] , \w3[6][23] , \w3[6][22] ,
         \w3[6][21] , \w3[6][20] , \w3[6][19] , \w3[6][18] , \w3[6][17] ,
         \w3[6][16] , \w3[6][15] , \w3[6][14] , \w3[6][13] , \w3[6][12] ,
         \w3[6][11] , \w3[6][10] , \w3[6][9] , \w3[6][8] , \w3[6][7] ,
         \w3[6][6] , \w3[6][5] , \w3[6][4] , \w3[6][3] , \w3[6][2] ,
         \w3[6][1] , \w3[6][0] , \w3[5][127] , \w3[5][126] , \w3[5][125] ,
         \w3[5][124] , \w3[5][123] , \w3[5][122] , \w3[5][121] , \w3[5][120] ,
         \w3[5][119] , \w3[5][118] , \w3[5][117] , \w3[5][116] , \w3[5][115] ,
         \w3[5][114] , \w3[5][113] , \w3[5][112] , \w3[5][111] , \w3[5][110] ,
         \w3[5][109] , \w3[5][108] , \w3[5][107] , \w3[5][106] , \w3[5][105] ,
         \w3[5][104] , \w3[5][103] , \w3[5][102] , \w3[5][101] , \w3[5][100] ,
         \w3[5][99] , \w3[5][98] , \w3[5][97] , \w3[5][96] , \w3[5][95] ,
         \w3[5][94] , \w3[5][93] , \w3[5][92] , \w3[5][91] , \w3[5][90] ,
         \w3[5][89] , \w3[5][88] , \w3[5][87] , \w3[5][86] , \w3[5][85] ,
         \w3[5][84] , \w3[5][83] , \w3[5][82] , \w3[5][81] , \w3[5][80] ,
         \w3[5][79] , \w3[5][78] , \w3[5][77] , \w3[5][76] , \w3[5][75] ,
         \w3[5][74] , \w3[5][73] , \w3[5][72] , \w3[5][71] , \w3[5][70] ,
         \w3[5][69] , \w3[5][68] , \w3[5][67] , \w3[5][66] , \w3[5][65] ,
         \w3[5][64] , \w3[5][63] , \w3[5][62] , \w3[5][61] , \w3[5][60] ,
         \w3[5][59] , \w3[5][58] , \w3[5][57] , \w3[5][56] , \w3[5][55] ,
         \w3[5][54] , \w3[5][53] , \w3[5][52] , \w3[5][51] , \w3[5][50] ,
         \w3[5][49] , \w3[5][48] , \w3[5][47] , \w3[5][46] , \w3[5][45] ,
         \w3[5][44] , \w3[5][43] , \w3[5][42] , \w3[5][41] , \w3[5][40] ,
         \w3[5][39] , \w3[5][38] , \w3[5][37] , \w3[5][36] , \w3[5][35] ,
         \w3[5][34] , \w3[5][33] , \w3[5][32] , \w3[5][31] , \w3[5][30] ,
         \w3[5][29] , \w3[5][28] , \w3[5][27] , \w3[5][26] , \w3[5][25] ,
         \w3[5][24] , \w3[5][23] , \w3[5][22] , \w3[5][21] , \w3[5][20] ,
         \w3[5][19] , \w3[5][18] , \w3[5][17] , \w3[5][16] , \w3[5][15] ,
         \w3[5][14] , \w3[5][13] , \w3[5][12] , \w3[5][11] , \w3[5][10] ,
         \w3[5][9] , \w3[5][8] , \w3[5][7] , \w3[5][6] , \w3[5][5] ,
         \w3[5][4] , \w3[5][3] , \w3[5][2] , \w3[5][1] , \w3[5][0] ,
         \w3[4][127] , \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] ,
         \w3[4][122] , \w3[4][121] , \w3[4][120] , \w3[4][119] , \w3[4][118] ,
         \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , \w3[4][113] ,
         \w3[4][112] , \w3[4][111] , \w3[4][110] , \w3[4][109] , \w3[4][108] ,
         \w3[4][107] , \w3[4][106] , \w3[4][105] , \w3[4][104] , \w3[4][103] ,
         \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] ,
         \w3[4][97] , \w3[4][96] , \w3[4][95] , \w3[4][94] , \w3[4][93] ,
         \w3[4][92] , \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] ,
         \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , \w3[4][83] ,
         \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][79] , \w3[4][78] ,
         \w3[4][77] , \w3[4][76] , \w3[4][75] , \w3[4][74] , \w3[4][73] ,
         \w3[4][72] , \w3[4][71] , \w3[4][70] , \w3[4][69] , \w3[4][68] ,
         \w3[4][67] , \w3[4][66] , \w3[4][65] , \w3[4][64] , \w3[4][63] ,
         \w3[4][62] , \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] ,
         \w3[4][57] , \w3[4][56] , \w3[4][55] , \w3[4][54] , \w3[4][53] ,
         \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , \w3[4][48] ,
         \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] ,
         \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][39] , \w3[4][38] ,
         \w3[4][37] , \w3[4][36] , \w3[4][35] , \w3[4][34] , \w3[4][33] ,
         \w3[4][32] , \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] ,
         \w3[4][27] , \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][23] ,
         \w3[4][22] , \w3[4][21] , \w3[4][20] , \w3[4][19] , \w3[4][18] ,
         \w3[4][17] , \w3[4][16] , \w3[4][15] , \w3[4][14] , \w3[4][13] ,
         \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] ,
         \w3[4][7] , \w3[4][6] , \w3[4][5] , \w3[4][4] , \w3[4][3] ,
         \w3[4][2] , \w3[4][1] , \w3[4][0] , \w3[3][127] , \w3[3][126] ,
         \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , \w3[3][121] ,
         \w3[3][120] , \w3[3][119] , \w3[3][118] , \w3[3][117] , \w3[3][116] ,
         \w3[3][115] , \w3[3][114] , \w3[3][113] , \w3[3][112] , \w3[3][111] ,
         \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] ,
         \w3[3][105] , \w3[3][104] , \w3[3][103] , \w3[3][102] , \w3[3][101] ,
         \w3[3][100] , \w3[3][99] , \w3[3][98] , \w3[3][97] , \w3[3][96] ,
         \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , \w3[3][91] ,
         \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][87] , \w3[3][86] ,
         \w3[3][85] , \w3[3][84] , \w3[3][83] , \w3[3][82] , \w3[3][81] ,
         \w3[3][80] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] ,
         \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][71] ,
         \w3[3][70] , \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] ,
         \w3[3][65] , \w3[3][64] , \w3[3][63] , \w3[3][62] , \w3[3][61] ,
         \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , \w3[3][56] ,
         \w3[3][55] , \w3[3][54] , \w3[3][53] , \w3[3][52] , \w3[3][51] ,
         \w3[3][50] , \w3[3][49] , \w3[3][48] , \w3[3][47] , \w3[3][46] ,
         \w3[3][45] , \w3[3][44] , \w3[3][43] , \w3[3][42] , \w3[3][41] ,
         \w3[3][40] , \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] ,
         \w3[3][35] , \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][31] ,
         \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , \w3[3][26] ,
         \w3[3][25] , \w3[3][24] , \w3[3][23] , \w3[3][22] , \w3[3][21] ,
         \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] ,
         \w3[3][15] , \w3[3][14] , \w3[3][13] , \w3[3][12] , \w3[3][11] ,
         \w3[3][10] , \w3[3][9] , \w3[3][8] , \w3[3][7] , \w3[3][6] ,
         \w3[3][5] , \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] ,
         \w3[3][0] , \w3[2][127] , \w3[2][126] , \w3[2][125] , \w3[2][124] ,
         \w3[2][123] , \w3[2][122] , \w3[2][121] , \w3[2][120] , \w3[2][119] ,
         \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] ,
         \w3[2][113] , \w3[2][112] , \w3[2][111] , \w3[2][110] , \w3[2][109] ,
         \w3[2][108] , \w3[2][107] , \w3[2][106] , \w3[2][105] , \w3[2][104] ,
         \w3[2][103] , \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] ,
         \w3[2][98] , \w3[2][97] , \w3[2][96] , \w3[2][95] , \w3[2][94] ,
         \w3[2][93] , \w3[2][92] , \w3[2][91] , \w3[2][90] , \w3[2][89] ,
         \w3[2][88] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] ,
         \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][79] ,
         \w3[2][78] , \w3[2][77] , \w3[2][76] , \w3[2][75] , \w3[2][74] ,
         \w3[2][73] , \w3[2][72] , \w3[2][71] , \w3[2][70] , \w3[2][69] ,
         \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , \w3[2][64] ,
         \w3[2][63] , \w3[2][62] , \w3[2][61] , \w3[2][60] , \w3[2][59] ,
         \w3[2][58] , \w3[2][57] , \w3[2][56] , \w3[2][55] , \w3[2][54] ,
         \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] ,
         \w3[2][48] , \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] ,
         \w3[2][43] , \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][39] ,
         \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , \w3[2][34] ,
         \w3[2][33] , \w3[2][32] , \w3[2][31] , \w3[2][30] , \w3[2][29] ,
         \w3[2][28] , \w3[2][27] , \w3[2][26] , \w3[2][25] , \w3[2][24] ,
         \w3[2][23] , \w3[2][22] , \w3[2][21] , \w3[2][20] , \w3[2][19] ,
         \w3[2][18] , \w3[2][17] , \w3[2][16] , \w3[2][15] , \w3[2][14] ,
         \w3[2][13] , \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] ,
         \w3[2][8] , \w3[2][7] , \w3[2][6] , \w3[2][5] , \w3[2][4] ,
         \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , \w3[1][127] ,
         \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] ,
         \w3[1][121] , \w3[1][120] , \w3[1][119] , \w3[1][118] , \w3[1][117] ,
         \w3[1][116] , \w3[1][115] , \w3[1][114] , \w3[1][113] , \w3[1][112] ,
         \w3[1][111] , \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] ,
         \w3[1][106] , \w3[1][105] , \w3[1][104] , \w3[1][103] , \w3[1][102] ,
         \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , \w3[1][97] ,
         \w3[1][96] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] ,
         \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][87] ,
         \w3[1][86] , \w3[1][85] , \w3[1][84] , \w3[1][83] , \w3[1][82] ,
         \w3[1][81] , \w3[1][80] , \w3[1][79] , \w3[1][78] , \w3[1][77] ,
         \w3[1][76] , \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] ,
         \w3[1][71] , \w3[1][70] , \w3[1][69] , \w3[1][68] , \w3[1][67] ,
         \w3[1][66] , \w3[1][65] , \w3[1][64] , \w3[1][63] , \w3[1][62] ,
         \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] ,
         \w3[1][56] , \w3[1][55] , \w3[1][54] , \w3[1][53] , \w3[1][52] ,
         \w3[1][51] , \w3[1][50] , \w3[1][49] , \w3[1][48] , \w3[1][47] ,
         \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , \w3[1][42] ,
         \w3[1][41] , \w3[1][40] , \w3[1][39] , \w3[1][38] , \w3[1][37] ,
         \w3[1][36] , \w3[1][35] , \w3[1][34] , \w3[1][33] , \w3[1][32] ,
         \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] ,
         \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][23] , \w3[1][22] ,
         \w3[1][21] , \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] ,
         \w3[1][16] , \w3[1][15] , \w3[1][14] , \w3[1][13] , \w3[1][12] ,
         \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , \w3[1][7] ,
         \w3[1][6] , \w3[1][5] , \w3[1][4] , \w3[1][3] , \w3[1][2] ,
         \w3[1][1] , \w3[1][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] ,
         \w3[0][124] , \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] ,
         \w3[0][119] , \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] ,
         \w3[0][114] , \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] ,
         \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] ,
         \w3[0][104] , \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] ,
         \w3[0][99] , \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] ,
         \w3[0][94] , \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] ,
         \w3[0][89] , \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] ,
         \w3[0][84] , \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] ,
         \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] ,
         \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] ,
         \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] ,
         \w3[0][64] , \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] ,
         \w3[0][59] , \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] ,
         \w3[0][54] , \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] ,
         \w3[0][49] , \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] ,
         \w3[0][44] , \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] ,
         \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] ,
         \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] ,
         \w3[0][29] , \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] ,
         \w3[0][24] , \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] ,
         \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] ,
         \w3[0][14] , \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] ,
         \w3[0][9] , \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] ,
         \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632;

  SubBytes_0 \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  SubBytes_9 \SUBBYTES[1].a  ( .x({\w1[1][127] , \w1[1][126] , \w1[1][125] , 
        \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , 
        \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , 
        \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , 
        \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , 
        \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , 
        \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , 
        \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , 
        \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , 
        \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , 
        \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , 
        \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , 
        \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , 
        \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , 
        \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , 
        \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , 
        \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , 
        \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , 
        \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , 
        \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , 
        \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , 
        \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , 
        \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , 
        \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , 
        \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] , 
        \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] }), .z({\w3[1][127] , 
        \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , 
        \w3[1][121] , \w3[1][120] , \w3[1][23] , \w3[1][22] , \w3[1][21] , 
        \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] , 
        \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , 
        \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][71] , \w3[1][70] , 
        \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] , \w3[1][65] , 
        \w3[1][64] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , 
        \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][119] , 
        \w3[1][118] , \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , 
        \w3[1][113] , \w3[1][112] , \w3[1][15] , \w3[1][14] , \w3[1][13] , 
        \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , 
        \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] , \w3[1][35] , 
        \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][63] , \w3[1][62] , 
        \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , 
        \w3[1][56] , \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , 
        \w3[1][83] , \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][111] , 
        \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] , 
        \w3[1][105] , \w3[1][104] , \w3[1][7] , \w3[1][6] , \w3[1][5] , 
        \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] , \w3[1][0] , 
        \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , 
        \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][55] , \w3[1][54] , 
        \w3[1][53] , \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , 
        \w3[1][48] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] , 
        \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][103] , 
        \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , 
        \w3[1][97] , \w3[1][96] }) );
  SubBytes_8 \SUBBYTES[2].a  ( .x({\w1[2][127] , \w1[2][126] , \w1[2][125] , 
        \w1[2][124] , \w1[2][123] , \w1[2][122] , \w1[2][121] , \w1[2][120] , 
        \w1[2][119] , \w1[2][118] , \w1[2][117] , \w1[2][116] , \w1[2][115] , 
        \w1[2][114] , \w1[2][113] , \w1[2][112] , \w1[2][111] , \w1[2][110] , 
        \w1[2][109] , \w1[2][108] , \w1[2][107] , \w1[2][106] , \w1[2][105] , 
        \w1[2][104] , \w1[2][103] , \w1[2][102] , \w1[2][101] , \w1[2][100] , 
        \w1[2][99] , \w1[2][98] , \w1[2][97] , \w1[2][96] , \w1[2][95] , 
        \w1[2][94] , \w1[2][93] , \w1[2][92] , \w1[2][91] , \w1[2][90] , 
        \w1[2][89] , \w1[2][88] , \w1[2][87] , \w1[2][86] , \w1[2][85] , 
        \w1[2][84] , \w1[2][83] , \w1[2][82] , \w1[2][81] , \w1[2][80] , 
        \w1[2][79] , \w1[2][78] , \w1[2][77] , \w1[2][76] , \w1[2][75] , 
        \w1[2][74] , \w1[2][73] , \w1[2][72] , \w1[2][71] , \w1[2][70] , 
        \w1[2][69] , \w1[2][68] , \w1[2][67] , \w1[2][66] , \w1[2][65] , 
        \w1[2][64] , \w1[2][63] , \w1[2][62] , \w1[2][61] , \w1[2][60] , 
        \w1[2][59] , \w1[2][58] , \w1[2][57] , \w1[2][56] , \w1[2][55] , 
        \w1[2][54] , \w1[2][53] , \w1[2][52] , \w1[2][51] , \w1[2][50] , 
        \w1[2][49] , \w1[2][48] , \w1[2][47] , \w1[2][46] , \w1[2][45] , 
        \w1[2][44] , \w1[2][43] , \w1[2][42] , \w1[2][41] , \w1[2][40] , 
        \w1[2][39] , \w1[2][38] , \w1[2][37] , \w1[2][36] , \w1[2][35] , 
        \w1[2][34] , \w1[2][33] , \w1[2][32] , \w1[2][31] , \w1[2][30] , 
        \w1[2][29] , \w1[2][28] , \w1[2][27] , \w1[2][26] , \w1[2][25] , 
        \w1[2][24] , \w1[2][23] , \w1[2][22] , \w1[2][21] , \w1[2][20] , 
        \w1[2][19] , \w1[2][18] , \w1[2][17] , \w1[2][16] , \w1[2][15] , 
        \w1[2][14] , \w1[2][13] , \w1[2][12] , \w1[2][11] , \w1[2][10] , 
        \w1[2][9] , \w1[2][8] , \w1[2][7] , \w1[2][6] , \w1[2][5] , \w1[2][4] , 
        \w1[2][3] , \w1[2][2] , \w1[2][1] , \w1[2][0] }), .z({\w3[2][127] , 
        \w3[2][126] , \w3[2][125] , \w3[2][124] , \w3[2][123] , \w3[2][122] , 
        \w3[2][121] , \w3[2][120] , \w3[2][23] , \w3[2][22] , \w3[2][21] , 
        \w3[2][20] , \w3[2][19] , \w3[2][18] , \w3[2][17] , \w3[2][16] , 
        \w3[2][47] , \w3[2][46] , \w3[2][45] , \w3[2][44] , \w3[2][43] , 
        \w3[2][42] , \w3[2][41] , \w3[2][40] , \w3[2][71] , \w3[2][70] , 
        \w3[2][69] , \w3[2][68] , \w3[2][67] , \w3[2][66] , \w3[2][65] , 
        \w3[2][64] , \w3[2][95] , \w3[2][94] , \w3[2][93] , \w3[2][92] , 
        \w3[2][91] , \w3[2][90] , \w3[2][89] , \w3[2][88] , \w3[2][119] , 
        \w3[2][118] , \w3[2][117] , \w3[2][116] , \w3[2][115] , \w3[2][114] , 
        \w3[2][113] , \w3[2][112] , \w3[2][15] , \w3[2][14] , \w3[2][13] , 
        \w3[2][12] , \w3[2][11] , \w3[2][10] , \w3[2][9] , \w3[2][8] , 
        \w3[2][39] , \w3[2][38] , \w3[2][37] , \w3[2][36] , \w3[2][35] , 
        \w3[2][34] , \w3[2][33] , \w3[2][32] , \w3[2][63] , \w3[2][62] , 
        \w3[2][61] , \w3[2][60] , \w3[2][59] , \w3[2][58] , \w3[2][57] , 
        \w3[2][56] , \w3[2][87] , \w3[2][86] , \w3[2][85] , \w3[2][84] , 
        \w3[2][83] , \w3[2][82] , \w3[2][81] , \w3[2][80] , \w3[2][111] , 
        \w3[2][110] , \w3[2][109] , \w3[2][108] , \w3[2][107] , \w3[2][106] , 
        \w3[2][105] , \w3[2][104] , \w3[2][7] , \w3[2][6] , \w3[2][5] , 
        \w3[2][4] , \w3[2][3] , \w3[2][2] , \w3[2][1] , \w3[2][0] , 
        \w3[2][31] , \w3[2][30] , \w3[2][29] , \w3[2][28] , \w3[2][27] , 
        \w3[2][26] , \w3[2][25] , \w3[2][24] , \w3[2][55] , \w3[2][54] , 
        \w3[2][53] , \w3[2][52] , \w3[2][51] , \w3[2][50] , \w3[2][49] , 
        \w3[2][48] , \w3[2][79] , \w3[2][78] , \w3[2][77] , \w3[2][76] , 
        \w3[2][75] , \w3[2][74] , \w3[2][73] , \w3[2][72] , \w3[2][103] , 
        \w3[2][102] , \w3[2][101] , \w3[2][100] , \w3[2][99] , \w3[2][98] , 
        \w3[2][97] , \w3[2][96] }) );
  SubBytes_7 \SUBBYTES[3].a  ( .x({\w1[3][127] , \w1[3][126] , \w1[3][125] , 
        \w1[3][124] , \w1[3][123] , \w1[3][122] , \w1[3][121] , \w1[3][120] , 
        \w1[3][119] , \w1[3][118] , \w1[3][117] , \w1[3][116] , \w1[3][115] , 
        \w1[3][114] , \w1[3][113] , \w1[3][112] , \w1[3][111] , \w1[3][110] , 
        \w1[3][109] , \w1[3][108] , \w1[3][107] , \w1[3][106] , \w1[3][105] , 
        \w1[3][104] , \w1[3][103] , \w1[3][102] , \w1[3][101] , \w1[3][100] , 
        \w1[3][99] , \w1[3][98] , \w1[3][97] , \w1[3][96] , \w1[3][95] , 
        \w1[3][94] , \w1[3][93] , \w1[3][92] , \w1[3][91] , \w1[3][90] , 
        \w1[3][89] , \w1[3][88] , \w1[3][87] , \w1[3][86] , \w1[3][85] , 
        \w1[3][84] , \w1[3][83] , \w1[3][82] , \w1[3][81] , \w1[3][80] , 
        \w1[3][79] , \w1[3][78] , \w1[3][77] , \w1[3][76] , \w1[3][75] , 
        \w1[3][74] , \w1[3][73] , \w1[3][72] , \w1[3][71] , \w1[3][70] , 
        \w1[3][69] , \w1[3][68] , \w1[3][67] , \w1[3][66] , \w1[3][65] , 
        \w1[3][64] , \w1[3][63] , \w1[3][62] , \w1[3][61] , \w1[3][60] , 
        \w1[3][59] , \w1[3][58] , \w1[3][57] , \w1[3][56] , \w1[3][55] , 
        \w1[3][54] , \w1[3][53] , \w1[3][52] , \w1[3][51] , \w1[3][50] , 
        \w1[3][49] , \w1[3][48] , \w1[3][47] , \w1[3][46] , \w1[3][45] , 
        \w1[3][44] , \w1[3][43] , \w1[3][42] , \w1[3][41] , \w1[3][40] , 
        \w1[3][39] , \w1[3][38] , \w1[3][37] , \w1[3][36] , \w1[3][35] , 
        \w1[3][34] , \w1[3][33] , \w1[3][32] , \w1[3][31] , \w1[3][30] , 
        \w1[3][29] , \w1[3][28] , \w1[3][27] , \w1[3][26] , \w1[3][25] , 
        \w1[3][24] , \w1[3][23] , \w1[3][22] , \w1[3][21] , \w1[3][20] , 
        \w1[3][19] , \w1[3][18] , \w1[3][17] , \w1[3][16] , \w1[3][15] , 
        \w1[3][14] , \w1[3][13] , \w1[3][12] , \w1[3][11] , \w1[3][10] , 
        \w1[3][9] , \w1[3][8] , \w1[3][7] , \w1[3][6] , \w1[3][5] , \w1[3][4] , 
        \w1[3][3] , \w1[3][2] , \w1[3][1] , \w1[3][0] }), .z({\w3[3][127] , 
        \w3[3][126] , \w3[3][125] , \w3[3][124] , \w3[3][123] , \w3[3][122] , 
        \w3[3][121] , \w3[3][120] , \w3[3][23] , \w3[3][22] , \w3[3][21] , 
        \w3[3][20] , \w3[3][19] , \w3[3][18] , \w3[3][17] , \w3[3][16] , 
        \w3[3][47] , \w3[3][46] , \w3[3][45] , \w3[3][44] , \w3[3][43] , 
        \w3[3][42] , \w3[3][41] , \w3[3][40] , \w3[3][71] , \w3[3][70] , 
        \w3[3][69] , \w3[3][68] , \w3[3][67] , \w3[3][66] , \w3[3][65] , 
        \w3[3][64] , \w3[3][95] , \w3[3][94] , \w3[3][93] , \w3[3][92] , 
        \w3[3][91] , \w3[3][90] , \w3[3][89] , \w3[3][88] , \w3[3][119] , 
        \w3[3][118] , \w3[3][117] , \w3[3][116] , \w3[3][115] , \w3[3][114] , 
        \w3[3][113] , \w3[3][112] , \w3[3][15] , \w3[3][14] , \w3[3][13] , 
        \w3[3][12] , \w3[3][11] , \w3[3][10] , \w3[3][9] , \w3[3][8] , 
        \w3[3][39] , \w3[3][38] , \w3[3][37] , \w3[3][36] , \w3[3][35] , 
        \w3[3][34] , \w3[3][33] , \w3[3][32] , \w3[3][63] , \w3[3][62] , 
        \w3[3][61] , \w3[3][60] , \w3[3][59] , \w3[3][58] , \w3[3][57] , 
        \w3[3][56] , \w3[3][87] , \w3[3][86] , \w3[3][85] , \w3[3][84] , 
        \w3[3][83] , \w3[3][82] , \w3[3][81] , \w3[3][80] , \w3[3][111] , 
        \w3[3][110] , \w3[3][109] , \w3[3][108] , \w3[3][107] , \w3[3][106] , 
        \w3[3][105] , \w3[3][104] , \w3[3][7] , \w3[3][6] , \w3[3][5] , 
        \w3[3][4] , \w3[3][3] , \w3[3][2] , \w3[3][1] , \w3[3][0] , 
        \w3[3][31] , \w3[3][30] , \w3[3][29] , \w3[3][28] , \w3[3][27] , 
        \w3[3][26] , \w3[3][25] , \w3[3][24] , \w3[3][55] , \w3[3][54] , 
        \w3[3][53] , \w3[3][52] , \w3[3][51] , \w3[3][50] , \w3[3][49] , 
        \w3[3][48] , \w3[3][79] , \w3[3][78] , \w3[3][77] , \w3[3][76] , 
        \w3[3][75] , \w3[3][74] , \w3[3][73] , \w3[3][72] , \w3[3][103] , 
        \w3[3][102] , \w3[3][101] , \w3[3][100] , \w3[3][99] , \w3[3][98] , 
        \w3[3][97] , \w3[3][96] }) );
  SubBytes_6 \SUBBYTES[4].a  ( .x({\w1[4][127] , \w1[4][126] , \w1[4][125] , 
        \w1[4][124] , \w1[4][123] , \w1[4][122] , \w1[4][121] , \w1[4][120] , 
        \w1[4][119] , \w1[4][118] , \w1[4][117] , \w1[4][116] , \w1[4][115] , 
        \w1[4][114] , \w1[4][113] , \w1[4][112] , \w1[4][111] , \w1[4][110] , 
        \w1[4][109] , \w1[4][108] , \w1[4][107] , \w1[4][106] , \w1[4][105] , 
        \w1[4][104] , \w1[4][103] , \w1[4][102] , \w1[4][101] , \w1[4][100] , 
        \w1[4][99] , \w1[4][98] , \w1[4][97] , \w1[4][96] , \w1[4][95] , 
        \w1[4][94] , \w1[4][93] , \w1[4][92] , \w1[4][91] , \w1[4][90] , 
        \w1[4][89] , \w1[4][88] , \w1[4][87] , \w1[4][86] , \w1[4][85] , 
        \w1[4][84] , \w1[4][83] , \w1[4][82] , \w1[4][81] , \w1[4][80] , 
        \w1[4][79] , \w1[4][78] , \w1[4][77] , \w1[4][76] , \w1[4][75] , 
        \w1[4][74] , \w1[4][73] , \w1[4][72] , \w1[4][71] , \w1[4][70] , 
        \w1[4][69] , \w1[4][68] , \w1[4][67] , \w1[4][66] , \w1[4][65] , 
        \w1[4][64] , \w1[4][63] , \w1[4][62] , \w1[4][61] , \w1[4][60] , 
        \w1[4][59] , \w1[4][58] , \w1[4][57] , \w1[4][56] , \w1[4][55] , 
        \w1[4][54] , \w1[4][53] , \w1[4][52] , \w1[4][51] , \w1[4][50] , 
        \w1[4][49] , \w1[4][48] , \w1[4][47] , \w1[4][46] , \w1[4][45] , 
        \w1[4][44] , \w1[4][43] , \w1[4][42] , \w1[4][41] , \w1[4][40] , 
        \w1[4][39] , \w1[4][38] , \w1[4][37] , \w1[4][36] , \w1[4][35] , 
        \w1[4][34] , \w1[4][33] , \w1[4][32] , \w1[4][31] , \w1[4][30] , 
        \w1[4][29] , \w1[4][28] , \w1[4][27] , \w1[4][26] , \w1[4][25] , 
        \w1[4][24] , \w1[4][23] , \w1[4][22] , \w1[4][21] , \w1[4][20] , 
        \w1[4][19] , \w1[4][18] , \w1[4][17] , \w1[4][16] , \w1[4][15] , 
        \w1[4][14] , \w1[4][13] , \w1[4][12] , \w1[4][11] , \w1[4][10] , 
        \w1[4][9] , \w1[4][8] , \w1[4][7] , \w1[4][6] , \w1[4][5] , \w1[4][4] , 
        \w1[4][3] , \w1[4][2] , \w1[4][1] , \w1[4][0] }), .z({\w3[4][127] , 
        \w3[4][126] , \w3[4][125] , \w3[4][124] , \w3[4][123] , \w3[4][122] , 
        \w3[4][121] , \w3[4][120] , \w3[4][23] , \w3[4][22] , \w3[4][21] , 
        \w3[4][20] , \w3[4][19] , \w3[4][18] , \w3[4][17] , \w3[4][16] , 
        \w3[4][47] , \w3[4][46] , \w3[4][45] , \w3[4][44] , \w3[4][43] , 
        \w3[4][42] , \w3[4][41] , \w3[4][40] , \w3[4][71] , \w3[4][70] , 
        \w3[4][69] , \w3[4][68] , \w3[4][67] , \w3[4][66] , \w3[4][65] , 
        \w3[4][64] , \w3[4][95] , \w3[4][94] , \w3[4][93] , \w3[4][92] , 
        \w3[4][91] , \w3[4][90] , \w3[4][89] , \w3[4][88] , \w3[4][119] , 
        \w3[4][118] , \w3[4][117] , \w3[4][116] , \w3[4][115] , \w3[4][114] , 
        \w3[4][113] , \w3[4][112] , \w3[4][15] , \w3[4][14] , \w3[4][13] , 
        \w3[4][12] , \w3[4][11] , \w3[4][10] , \w3[4][9] , \w3[4][8] , 
        \w3[4][39] , \w3[4][38] , \w3[4][37] , \w3[4][36] , \w3[4][35] , 
        \w3[4][34] , \w3[4][33] , \w3[4][32] , \w3[4][63] , \w3[4][62] , 
        \w3[4][61] , \w3[4][60] , \w3[4][59] , \w3[4][58] , \w3[4][57] , 
        \w3[4][56] , \w3[4][87] , \w3[4][86] , \w3[4][85] , \w3[4][84] , 
        \w3[4][83] , \w3[4][82] , \w3[4][81] , \w3[4][80] , \w3[4][111] , 
        \w3[4][110] , \w3[4][109] , \w3[4][108] , \w3[4][107] , \w3[4][106] , 
        \w3[4][105] , \w3[4][104] , \w3[4][7] , \w3[4][6] , \w3[4][5] , 
        \w3[4][4] , \w3[4][3] , \w3[4][2] , \w3[4][1] , \w3[4][0] , 
        \w3[4][31] , \w3[4][30] , \w3[4][29] , \w3[4][28] , \w3[4][27] , 
        \w3[4][26] , \w3[4][25] , \w3[4][24] , \w3[4][55] , \w3[4][54] , 
        \w3[4][53] , \w3[4][52] , \w3[4][51] , \w3[4][50] , \w3[4][49] , 
        \w3[4][48] , \w3[4][79] , \w3[4][78] , \w3[4][77] , \w3[4][76] , 
        \w3[4][75] , \w3[4][74] , \w3[4][73] , \w3[4][72] , \w3[4][103] , 
        \w3[4][102] , \w3[4][101] , \w3[4][100] , \w3[4][99] , \w3[4][98] , 
        \w3[4][97] , \w3[4][96] }) );
  SubBytes_5 \SUBBYTES[5].a  ( .x({\w1[5][127] , \w1[5][126] , \w1[5][125] , 
        \w1[5][124] , \w1[5][123] , \w1[5][122] , \w1[5][121] , \w1[5][120] , 
        \w1[5][119] , \w1[5][118] , \w1[5][117] , \w1[5][116] , \w1[5][115] , 
        \w1[5][114] , \w1[5][113] , \w1[5][112] , \w1[5][111] , \w1[5][110] , 
        \w1[5][109] , \w1[5][108] , \w1[5][107] , \w1[5][106] , \w1[5][105] , 
        \w1[5][104] , \w1[5][103] , \w1[5][102] , \w1[5][101] , \w1[5][100] , 
        \w1[5][99] , \w1[5][98] , \w1[5][97] , \w1[5][96] , \w1[5][95] , 
        \w1[5][94] , \w1[5][93] , \w1[5][92] , \w1[5][91] , \w1[5][90] , 
        \w1[5][89] , \w1[5][88] , \w1[5][87] , \w1[5][86] , \w1[5][85] , 
        \w1[5][84] , \w1[5][83] , \w1[5][82] , \w1[5][81] , \w1[5][80] , 
        \w1[5][79] , \w1[5][78] , \w1[5][77] , \w1[5][76] , \w1[5][75] , 
        \w1[5][74] , \w1[5][73] , \w1[5][72] , \w1[5][71] , \w1[5][70] , 
        \w1[5][69] , \w1[5][68] , \w1[5][67] , \w1[5][66] , \w1[5][65] , 
        \w1[5][64] , \w1[5][63] , \w1[5][62] , \w1[5][61] , \w1[5][60] , 
        \w1[5][59] , \w1[5][58] , \w1[5][57] , \w1[5][56] , \w1[5][55] , 
        \w1[5][54] , \w1[5][53] , \w1[5][52] , \w1[5][51] , \w1[5][50] , 
        \w1[5][49] , \w1[5][48] , \w1[5][47] , \w1[5][46] , \w1[5][45] , 
        \w1[5][44] , \w1[5][43] , \w1[5][42] , \w1[5][41] , \w1[5][40] , 
        \w1[5][39] , \w1[5][38] , \w1[5][37] , \w1[5][36] , \w1[5][35] , 
        \w1[5][34] , \w1[5][33] , \w1[5][32] , \w1[5][31] , \w1[5][30] , 
        \w1[5][29] , \w1[5][28] , \w1[5][27] , \w1[5][26] , \w1[5][25] , 
        \w1[5][24] , \w1[5][23] , \w1[5][22] , \w1[5][21] , \w1[5][20] , 
        \w1[5][19] , \w1[5][18] , \w1[5][17] , \w1[5][16] , \w1[5][15] , 
        \w1[5][14] , \w1[5][13] , \w1[5][12] , \w1[5][11] , \w1[5][10] , 
        \w1[5][9] , \w1[5][8] , \w1[5][7] , \w1[5][6] , \w1[5][5] , \w1[5][4] , 
        \w1[5][3] , \w1[5][2] , \w1[5][1] , \w1[5][0] }), .z({\w3[5][127] , 
        \w3[5][126] , \w3[5][125] , \w3[5][124] , \w3[5][123] , \w3[5][122] , 
        \w3[5][121] , \w3[5][120] , \w3[5][23] , \w3[5][22] , \w3[5][21] , 
        \w3[5][20] , \w3[5][19] , \w3[5][18] , \w3[5][17] , \w3[5][16] , 
        \w3[5][47] , \w3[5][46] , \w3[5][45] , \w3[5][44] , \w3[5][43] , 
        \w3[5][42] , \w3[5][41] , \w3[5][40] , \w3[5][71] , \w3[5][70] , 
        \w3[5][69] , \w3[5][68] , \w3[5][67] , \w3[5][66] , \w3[5][65] , 
        \w3[5][64] , \w3[5][95] , \w3[5][94] , \w3[5][93] , \w3[5][92] , 
        \w3[5][91] , \w3[5][90] , \w3[5][89] , \w3[5][88] , \w3[5][119] , 
        \w3[5][118] , \w3[5][117] , \w3[5][116] , \w3[5][115] , \w3[5][114] , 
        \w3[5][113] , \w3[5][112] , \w3[5][15] , \w3[5][14] , \w3[5][13] , 
        \w3[5][12] , \w3[5][11] , \w3[5][10] , \w3[5][9] , \w3[5][8] , 
        \w3[5][39] , \w3[5][38] , \w3[5][37] , \w3[5][36] , \w3[5][35] , 
        \w3[5][34] , \w3[5][33] , \w3[5][32] , \w3[5][63] , \w3[5][62] , 
        \w3[5][61] , \w3[5][60] , \w3[5][59] , \w3[5][58] , \w3[5][57] , 
        \w3[5][56] , \w3[5][87] , \w3[5][86] , \w3[5][85] , \w3[5][84] , 
        \w3[5][83] , \w3[5][82] , \w3[5][81] , \w3[5][80] , \w3[5][111] , 
        \w3[5][110] , \w3[5][109] , \w3[5][108] , \w3[5][107] , \w3[5][106] , 
        \w3[5][105] , \w3[5][104] , \w3[5][7] , \w3[5][6] , \w3[5][5] , 
        \w3[5][4] , \w3[5][3] , \w3[5][2] , \w3[5][1] , \w3[5][0] , 
        \w3[5][31] , \w3[5][30] , \w3[5][29] , \w3[5][28] , \w3[5][27] , 
        \w3[5][26] , \w3[5][25] , \w3[5][24] , \w3[5][55] , \w3[5][54] , 
        \w3[5][53] , \w3[5][52] , \w3[5][51] , \w3[5][50] , \w3[5][49] , 
        \w3[5][48] , \w3[5][79] , \w3[5][78] , \w3[5][77] , \w3[5][76] , 
        \w3[5][75] , \w3[5][74] , \w3[5][73] , \w3[5][72] , \w3[5][103] , 
        \w3[5][102] , \w3[5][101] , \w3[5][100] , \w3[5][99] , \w3[5][98] , 
        \w3[5][97] , \w3[5][96] }) );
  SubBytes_4 \SUBBYTES[6].a  ( .x({\w1[6][127] , \w1[6][126] , \w1[6][125] , 
        \w1[6][124] , \w1[6][123] , \w1[6][122] , \w1[6][121] , \w1[6][120] , 
        \w1[6][119] , \w1[6][118] , \w1[6][117] , \w1[6][116] , \w1[6][115] , 
        \w1[6][114] , \w1[6][113] , \w1[6][112] , \w1[6][111] , \w1[6][110] , 
        \w1[6][109] , \w1[6][108] , \w1[6][107] , \w1[6][106] , \w1[6][105] , 
        \w1[6][104] , \w1[6][103] , \w1[6][102] , \w1[6][101] , \w1[6][100] , 
        \w1[6][99] , \w1[6][98] , \w1[6][97] , \w1[6][96] , \w1[6][95] , 
        \w1[6][94] , \w1[6][93] , \w1[6][92] , \w1[6][91] , \w1[6][90] , 
        \w1[6][89] , \w1[6][88] , \w1[6][87] , \w1[6][86] , \w1[6][85] , 
        \w1[6][84] , \w1[6][83] , \w1[6][82] , \w1[6][81] , \w1[6][80] , 
        \w1[6][79] , \w1[6][78] , \w1[6][77] , \w1[6][76] , \w1[6][75] , 
        \w1[6][74] , \w1[6][73] , \w1[6][72] , \w1[6][71] , \w1[6][70] , 
        \w1[6][69] , \w1[6][68] , \w1[6][67] , \w1[6][66] , \w1[6][65] , 
        \w1[6][64] , \w1[6][63] , \w1[6][62] , \w1[6][61] , \w1[6][60] , 
        \w1[6][59] , \w1[6][58] , \w1[6][57] , \w1[6][56] , \w1[6][55] , 
        \w1[6][54] , \w1[6][53] , \w1[6][52] , \w1[6][51] , \w1[6][50] , 
        \w1[6][49] , \w1[6][48] , \w1[6][47] , \w1[6][46] , \w1[6][45] , 
        \w1[6][44] , \w1[6][43] , \w1[6][42] , \w1[6][41] , \w1[6][40] , 
        \w1[6][39] , \w1[6][38] , \w1[6][37] , \w1[6][36] , \w1[6][35] , 
        \w1[6][34] , \w1[6][33] , \w1[6][32] , \w1[6][31] , \w1[6][30] , 
        \w1[6][29] , \w1[6][28] , \w1[6][27] , \w1[6][26] , \w1[6][25] , 
        \w1[6][24] , \w1[6][23] , \w1[6][22] , \w1[6][21] , \w1[6][20] , 
        \w1[6][19] , \w1[6][18] , \w1[6][17] , \w1[6][16] , \w1[6][15] , 
        \w1[6][14] , \w1[6][13] , \w1[6][12] , \w1[6][11] , \w1[6][10] , 
        \w1[6][9] , \w1[6][8] , \w1[6][7] , \w1[6][6] , \w1[6][5] , \w1[6][4] , 
        \w1[6][3] , \w1[6][2] , \w1[6][1] , \w1[6][0] }), .z({\w3[6][127] , 
        \w3[6][126] , \w3[6][125] , \w3[6][124] , \w3[6][123] , \w3[6][122] , 
        \w3[6][121] , \w3[6][120] , \w3[6][23] , \w3[6][22] , \w3[6][21] , 
        \w3[6][20] , \w3[6][19] , \w3[6][18] , \w3[6][17] , \w3[6][16] , 
        \w3[6][47] , \w3[6][46] , \w3[6][45] , \w3[6][44] , \w3[6][43] , 
        \w3[6][42] , \w3[6][41] , \w3[6][40] , \w3[6][71] , \w3[6][70] , 
        \w3[6][69] , \w3[6][68] , \w3[6][67] , \w3[6][66] , \w3[6][65] , 
        \w3[6][64] , \w3[6][95] , \w3[6][94] , \w3[6][93] , \w3[6][92] , 
        \w3[6][91] , \w3[6][90] , \w3[6][89] , \w3[6][88] , \w3[6][119] , 
        \w3[6][118] , \w3[6][117] , \w3[6][116] , \w3[6][115] , \w3[6][114] , 
        \w3[6][113] , \w3[6][112] , \w3[6][15] , \w3[6][14] , \w3[6][13] , 
        \w3[6][12] , \w3[6][11] , \w3[6][10] , \w3[6][9] , \w3[6][8] , 
        \w3[6][39] , \w3[6][38] , \w3[6][37] , \w3[6][36] , \w3[6][35] , 
        \w3[6][34] , \w3[6][33] , \w3[6][32] , \w3[6][63] , \w3[6][62] , 
        \w3[6][61] , \w3[6][60] , \w3[6][59] , \w3[6][58] , \w3[6][57] , 
        \w3[6][56] , \w3[6][87] , \w3[6][86] , \w3[6][85] , \w3[6][84] , 
        \w3[6][83] , \w3[6][82] , \w3[6][81] , \w3[6][80] , \w3[6][111] , 
        \w3[6][110] , \w3[6][109] , \w3[6][108] , \w3[6][107] , \w3[6][106] , 
        \w3[6][105] , \w3[6][104] , \w3[6][7] , \w3[6][6] , \w3[6][5] , 
        \w3[6][4] , \w3[6][3] , \w3[6][2] , \w3[6][1] , \w3[6][0] , 
        \w3[6][31] , \w3[6][30] , \w3[6][29] , \w3[6][28] , \w3[6][27] , 
        \w3[6][26] , \w3[6][25] , \w3[6][24] , \w3[6][55] , \w3[6][54] , 
        \w3[6][53] , \w3[6][52] , \w3[6][51] , \w3[6][50] , \w3[6][49] , 
        \w3[6][48] , \w3[6][79] , \w3[6][78] , \w3[6][77] , \w3[6][76] , 
        \w3[6][75] , \w3[6][74] , \w3[6][73] , \w3[6][72] , \w3[6][103] , 
        \w3[6][102] , \w3[6][101] , \w3[6][100] , \w3[6][99] , \w3[6][98] , 
        \w3[6][97] , \w3[6][96] }) );
  SubBytes_3 \SUBBYTES[7].a  ( .x({\w1[7][127] , \w1[7][126] , \w1[7][125] , 
        \w1[7][124] , \w1[7][123] , \w1[7][122] , \w1[7][121] , \w1[7][120] , 
        \w1[7][119] , \w1[7][118] , \w1[7][117] , \w1[7][116] , \w1[7][115] , 
        \w1[7][114] , \w1[7][113] , \w1[7][112] , \w1[7][111] , \w1[7][110] , 
        \w1[7][109] , \w1[7][108] , \w1[7][107] , \w1[7][106] , \w1[7][105] , 
        \w1[7][104] , \w1[7][103] , \w1[7][102] , \w1[7][101] , \w1[7][100] , 
        \w1[7][99] , \w1[7][98] , \w1[7][97] , \w1[7][96] , \w1[7][95] , 
        \w1[7][94] , \w1[7][93] , \w1[7][92] , \w1[7][91] , \w1[7][90] , 
        \w1[7][89] , \w1[7][88] , \w1[7][87] , \w1[7][86] , \w1[7][85] , 
        \w1[7][84] , \w1[7][83] , \w1[7][82] , \w1[7][81] , \w1[7][80] , 
        \w1[7][79] , \w1[7][78] , \w1[7][77] , \w1[7][76] , \w1[7][75] , 
        \w1[7][74] , \w1[7][73] , \w1[7][72] , \w1[7][71] , \w1[7][70] , 
        \w1[7][69] , \w1[7][68] , \w1[7][67] , \w1[7][66] , \w1[7][65] , 
        \w1[7][64] , \w1[7][63] , \w1[7][62] , \w1[7][61] , \w1[7][60] , 
        \w1[7][59] , \w1[7][58] , \w1[7][57] , \w1[7][56] , \w1[7][55] , 
        \w1[7][54] , \w1[7][53] , \w1[7][52] , \w1[7][51] , \w1[7][50] , 
        \w1[7][49] , \w1[7][48] , \w1[7][47] , \w1[7][46] , \w1[7][45] , 
        \w1[7][44] , \w1[7][43] , \w1[7][42] , \w1[7][41] , \w1[7][40] , 
        \w1[7][39] , \w1[7][38] , \w1[7][37] , \w1[7][36] , \w1[7][35] , 
        \w1[7][34] , \w1[7][33] , \w1[7][32] , \w1[7][31] , \w1[7][30] , 
        \w1[7][29] , \w1[7][28] , \w1[7][27] , \w1[7][26] , \w1[7][25] , 
        \w1[7][24] , \w1[7][23] , \w1[7][22] , \w1[7][21] , \w1[7][20] , 
        \w1[7][19] , \w1[7][18] , \w1[7][17] , \w1[7][16] , \w1[7][15] , 
        \w1[7][14] , \w1[7][13] , \w1[7][12] , \w1[7][11] , \w1[7][10] , 
        \w1[7][9] , \w1[7][8] , \w1[7][7] , \w1[7][6] , \w1[7][5] , \w1[7][4] , 
        \w1[7][3] , \w1[7][2] , \w1[7][1] , \w1[7][0] }), .z({\w3[7][127] , 
        \w3[7][126] , \w3[7][125] , \w3[7][124] , \w3[7][123] , \w3[7][122] , 
        \w3[7][121] , \w3[7][120] , \w3[7][23] , \w3[7][22] , \w3[7][21] , 
        \w3[7][20] , \w3[7][19] , \w3[7][18] , \w3[7][17] , \w3[7][16] , 
        \w3[7][47] , \w3[7][46] , \w3[7][45] , \w3[7][44] , \w3[7][43] , 
        \w3[7][42] , \w3[7][41] , \w3[7][40] , \w3[7][71] , \w3[7][70] , 
        \w3[7][69] , \w3[7][68] , \w3[7][67] , \w3[7][66] , \w3[7][65] , 
        \w3[7][64] , \w3[7][95] , \w3[7][94] , \w3[7][93] , \w3[7][92] , 
        \w3[7][91] , \w3[7][90] , \w3[7][89] , \w3[7][88] , \w3[7][119] , 
        \w3[7][118] , \w3[7][117] , \w3[7][116] , \w3[7][115] , \w3[7][114] , 
        \w3[7][113] , \w3[7][112] , \w3[7][15] , \w3[7][14] , \w3[7][13] , 
        \w3[7][12] , \w3[7][11] , \w3[7][10] , \w3[7][9] , \w3[7][8] , 
        \w3[7][39] , \w3[7][38] , \w3[7][37] , \w3[7][36] , \w3[7][35] , 
        \w3[7][34] , \w3[7][33] , \w3[7][32] , \w3[7][63] , \w3[7][62] , 
        \w3[7][61] , \w3[7][60] , \w3[7][59] , \w3[7][58] , \w3[7][57] , 
        \w3[7][56] , \w3[7][87] , \w3[7][86] , \w3[7][85] , \w3[7][84] , 
        \w3[7][83] , \w3[7][82] , \w3[7][81] , \w3[7][80] , \w3[7][111] , 
        \w3[7][110] , \w3[7][109] , \w3[7][108] , \w3[7][107] , \w3[7][106] , 
        \w3[7][105] , \w3[7][104] , \w3[7][7] , \w3[7][6] , \w3[7][5] , 
        \w3[7][4] , \w3[7][3] , \w3[7][2] , \w3[7][1] , \w3[7][0] , 
        \w3[7][31] , \w3[7][30] , \w3[7][29] , \w3[7][28] , \w3[7][27] , 
        \w3[7][26] , \w3[7][25] , \w3[7][24] , \w3[7][55] , \w3[7][54] , 
        \w3[7][53] , \w3[7][52] , \w3[7][51] , \w3[7][50] , \w3[7][49] , 
        \w3[7][48] , \w3[7][79] , \w3[7][78] , \w3[7][77] , \w3[7][76] , 
        \w3[7][75] , \w3[7][74] , \w3[7][73] , \w3[7][72] , \w3[7][103] , 
        \w3[7][102] , \w3[7][101] , \w3[7][100] , \w3[7][99] , \w3[7][98] , 
        \w3[7][97] , \w3[7][96] }) );
  SubBytes_2 \SUBBYTES[8].a  ( .x({\w1[8][127] , \w1[8][126] , \w1[8][125] , 
        \w1[8][124] , \w1[8][123] , \w1[8][122] , \w1[8][121] , \w1[8][120] , 
        \w1[8][119] , \w1[8][118] , \w1[8][117] , \w1[8][116] , \w1[8][115] , 
        \w1[8][114] , \w1[8][113] , \w1[8][112] , \w1[8][111] , \w1[8][110] , 
        \w1[8][109] , \w1[8][108] , \w1[8][107] , \w1[8][106] , \w1[8][105] , 
        \w1[8][104] , \w1[8][103] , \w1[8][102] , \w1[8][101] , \w1[8][100] , 
        \w1[8][99] , \w1[8][98] , \w1[8][97] , \w1[8][96] , \w1[8][95] , 
        \w1[8][94] , \w1[8][93] , \w1[8][92] , \w1[8][91] , \w1[8][90] , 
        \w1[8][89] , \w1[8][88] , \w1[8][87] , \w1[8][86] , \w1[8][85] , 
        \w1[8][84] , \w1[8][83] , \w1[8][82] , \w1[8][81] , \w1[8][80] , 
        \w1[8][79] , \w1[8][78] , \w1[8][77] , \w1[8][76] , \w1[8][75] , 
        \w1[8][74] , \w1[8][73] , \w1[8][72] , \w1[8][71] , \w1[8][70] , 
        \w1[8][69] , \w1[8][68] , \w1[8][67] , \w1[8][66] , \w1[8][65] , 
        \w1[8][64] , \w1[8][63] , \w1[8][62] , \w1[8][61] , \w1[8][60] , 
        \w1[8][59] , \w1[8][58] , \w1[8][57] , \w1[8][56] , \w1[8][55] , 
        \w1[8][54] , \w1[8][53] , \w1[8][52] , \w1[8][51] , \w1[8][50] , 
        \w1[8][49] , \w1[8][48] , \w1[8][47] , \w1[8][46] , \w1[8][45] , 
        \w1[8][44] , \w1[8][43] , \w1[8][42] , \w1[8][41] , \w1[8][40] , 
        \w1[8][39] , \w1[8][38] , \w1[8][37] , \w1[8][36] , \w1[8][35] , 
        \w1[8][34] , \w1[8][33] , \w1[8][32] , \w1[8][31] , \w1[8][30] , 
        \w1[8][29] , \w1[8][28] , \w1[8][27] , \w1[8][26] , \w1[8][25] , 
        \w1[8][24] , \w1[8][23] , \w1[8][22] , \w1[8][21] , \w1[8][20] , 
        \w1[8][19] , \w1[8][18] , \w1[8][17] , \w1[8][16] , \w1[8][15] , 
        \w1[8][14] , \w1[8][13] , \w1[8][12] , \w1[8][11] , \w1[8][10] , 
        \w1[8][9] , \w1[8][8] , \w1[8][7] , \w1[8][6] , \w1[8][5] , \w1[8][4] , 
        \w1[8][3] , \w1[8][2] , \w1[8][1] , \w1[8][0] }), .z({\w3[8][127] , 
        \w3[8][126] , \w3[8][125] , \w3[8][124] , \w3[8][123] , \w3[8][122] , 
        \w3[8][121] , \w3[8][120] , \w3[8][23] , \w3[8][22] , \w3[8][21] , 
        \w3[8][20] , \w3[8][19] , \w3[8][18] , \w3[8][17] , \w3[8][16] , 
        \w3[8][47] , \w3[8][46] , \w3[8][45] , \w3[8][44] , \w3[8][43] , 
        \w3[8][42] , \w3[8][41] , \w3[8][40] , \w3[8][71] , \w3[8][70] , 
        \w3[8][69] , \w3[8][68] , \w3[8][67] , \w3[8][66] , \w3[8][65] , 
        \w3[8][64] , \w3[8][95] , \w3[8][94] , \w3[8][93] , \w3[8][92] , 
        \w3[8][91] , \w3[8][90] , \w3[8][89] , \w3[8][88] , \w3[8][119] , 
        \w3[8][118] , \w3[8][117] , \w3[8][116] , \w3[8][115] , \w3[8][114] , 
        \w3[8][113] , \w3[8][112] , \w3[8][15] , \w3[8][14] , \w3[8][13] , 
        \w3[8][12] , \w3[8][11] , \w3[8][10] , \w3[8][9] , \w3[8][8] , 
        \w3[8][39] , \w3[8][38] , \w3[8][37] , \w3[8][36] , \w3[8][35] , 
        \w3[8][34] , \w3[8][33] , \w3[8][32] , \w3[8][63] , \w3[8][62] , 
        \w3[8][61] , \w3[8][60] , \w3[8][59] , \w3[8][58] , \w3[8][57] , 
        \w3[8][56] , \w3[8][87] , \w3[8][86] , \w3[8][85] , \w3[8][84] , 
        \w3[8][83] , \w3[8][82] , \w3[8][81] , \w3[8][80] , \w3[8][111] , 
        \w3[8][110] , \w3[8][109] , \w3[8][108] , \w3[8][107] , \w3[8][106] , 
        \w3[8][105] , \w3[8][104] , \w3[8][7] , \w3[8][6] , \w3[8][5] , 
        \w3[8][4] , \w3[8][3] , \w3[8][2] , \w3[8][1] , \w3[8][0] , 
        \w3[8][31] , \w3[8][30] , \w3[8][29] , \w3[8][28] , \w3[8][27] , 
        \w3[8][26] , \w3[8][25] , \w3[8][24] , \w3[8][55] , \w3[8][54] , 
        \w3[8][53] , \w3[8][52] , \w3[8][51] , \w3[8][50] , \w3[8][49] , 
        \w3[8][48] , \w3[8][79] , \w3[8][78] , \w3[8][77] , \w3[8][76] , 
        \w3[8][75] , \w3[8][74] , \w3[8][73] , \w3[8][72] , \w3[8][103] , 
        \w3[8][102] , \w3[8][101] , \w3[8][100] , \w3[8][99] , \w3[8][98] , 
        \w3[8][97] , \w3[8][96] }) );
  SubBytes_1 \SUBBYTES[9].a  ( .x({\w1[9][127] , \w1[9][126] , \w1[9][125] , 
        \w1[9][124] , \w1[9][123] , \w1[9][122] , \w1[9][121] , \w1[9][120] , 
        \w1[9][119] , \w1[9][118] , \w1[9][117] , \w1[9][116] , \w1[9][115] , 
        \w1[9][114] , \w1[9][113] , \w1[9][112] , \w1[9][111] , \w1[9][110] , 
        \w1[9][109] , \w1[9][108] , \w1[9][107] , \w1[9][106] , \w1[9][105] , 
        \w1[9][104] , \w1[9][103] , \w1[9][102] , \w1[9][101] , \w1[9][100] , 
        \w1[9][99] , \w1[9][98] , \w1[9][97] , \w1[9][96] , \w1[9][95] , 
        \w1[9][94] , \w1[9][93] , \w1[9][92] , \w1[9][91] , \w1[9][90] , 
        \w1[9][89] , \w1[9][88] , \w1[9][87] , \w1[9][86] , \w1[9][85] , 
        \w1[9][84] , \w1[9][83] , \w1[9][82] , \w1[9][81] , \w1[9][80] , 
        \w1[9][79] , \w1[9][78] , \w1[9][77] , \w1[9][76] , \w1[9][75] , 
        \w1[9][74] , \w1[9][73] , \w1[9][72] , \w1[9][71] , \w1[9][70] , 
        \w1[9][69] , \w1[9][68] , \w1[9][67] , \w1[9][66] , \w1[9][65] , 
        \w1[9][64] , \w1[9][63] , \w1[9][62] , \w1[9][61] , \w1[9][60] , 
        \w1[9][59] , \w1[9][58] , \w1[9][57] , \w1[9][56] , \w1[9][55] , 
        \w1[9][54] , \w1[9][53] , \w1[9][52] , \w1[9][51] , \w1[9][50] , 
        \w1[9][49] , \w1[9][48] , \w1[9][47] , \w1[9][46] , \w1[9][45] , 
        \w1[9][44] , \w1[9][43] , \w1[9][42] , \w1[9][41] , \w1[9][40] , 
        \w1[9][39] , \w1[9][38] , \w1[9][37] , \w1[9][36] , \w1[9][35] , 
        \w1[9][34] , \w1[9][33] , \w1[9][32] , \w1[9][31] , \w1[9][30] , 
        \w1[9][29] , \w1[9][28] , \w1[9][27] , \w1[9][26] , \w1[9][25] , 
        \w1[9][24] , \w1[9][23] , \w1[9][22] , \w1[9][21] , \w1[9][20] , 
        \w1[9][19] , \w1[9][18] , \w1[9][17] , \w1[9][16] , \w1[9][15] , 
        \w1[9][14] , \w1[9][13] , \w1[9][12] , \w1[9][11] , \w1[9][10] , 
        \w1[9][9] , \w1[9][8] , \w1[9][7] , \w1[9][6] , \w1[9][5] , \w1[9][4] , 
        \w1[9][3] , \w1[9][2] , \w1[9][1] , \w1[9][0] }), .z({\w3[9][127] , 
        \w3[9][126] , \w3[9][125] , \w3[9][124] , \w3[9][123] , \w3[9][122] , 
        \w3[9][121] , \w3[9][120] , \w3[9][23] , \w3[9][22] , \w3[9][21] , 
        \w3[9][20] , \w3[9][19] , \w3[9][18] , \w3[9][17] , \w3[9][16] , 
        \w3[9][47] , \w3[9][46] , \w3[9][45] , \w3[9][44] , \w3[9][43] , 
        \w3[9][42] , \w3[9][41] , \w3[9][40] , \w3[9][71] , \w3[9][70] , 
        \w3[9][69] , \w3[9][68] , \w3[9][67] , \w3[9][66] , \w3[9][65] , 
        \w3[9][64] , \w3[9][95] , \w3[9][94] , \w3[9][93] , \w3[9][92] , 
        \w3[9][91] , \w3[9][90] , \w3[9][89] , \w3[9][88] , \w3[9][119] , 
        \w3[9][118] , \w3[9][117] , \w3[9][116] , \w3[9][115] , \w3[9][114] , 
        \w3[9][113] , \w3[9][112] , \w3[9][15] , \w3[9][14] , \w3[9][13] , 
        \w3[9][12] , \w3[9][11] , \w3[9][10] , \w3[9][9] , \w3[9][8] , 
        \w3[9][39] , \w3[9][38] , \w3[9][37] , \w3[9][36] , \w3[9][35] , 
        \w3[9][34] , \w3[9][33] , \w3[9][32] , \w3[9][63] , \w3[9][62] , 
        \w3[9][61] , \w3[9][60] , \w3[9][59] , \w3[9][58] , \w3[9][57] , 
        \w3[9][56] , \w3[9][87] , \w3[9][86] , \w3[9][85] , \w3[9][84] , 
        \w3[9][83] , \w3[9][82] , \w3[9][81] , \w3[9][80] , \w3[9][111] , 
        \w3[9][110] , \w3[9][109] , \w3[9][108] , \w3[9][107] , \w3[9][106] , 
        \w3[9][105] , \w3[9][104] , \w3[9][7] , \w3[9][6] , \w3[9][5] , 
        \w3[9][4] , \w3[9][3] , \w3[9][2] , \w3[9][1] , \w3[9][0] , 
        \w3[9][31] , \w3[9][30] , \w3[9][29] , \w3[9][28] , \w3[9][27] , 
        \w3[9][26] , \w3[9][25] , \w3[9][24] , \w3[9][55] , \w3[9][54] , 
        \w3[9][53] , \w3[9][52] , \w3[9][51] , \w3[9][50] , \w3[9][49] , 
        \w3[9][48] , \w3[9][79] , \w3[9][78] , \w3[9][77] , \w3[9][76] , 
        \w3[9][75] , \w3[9][74] , \w3[9][73] , \w3[9][72] , \w3[9][103] , 
        \w3[9][102] , \w3[9][101] , \w3[9][100] , \w3[9][99] , \w3[9][98] , 
        \w3[9][97] , \w3[9][96] }) );
  XOR U5225 ( .A(key[1152]), .B(\w3[9][0] ), .Z(out[0]) );
  XOR U5226 ( .A(key[1252]), .B(\w3[9][100] ), .Z(out[100]) );
  XOR U5227 ( .A(key[1253]), .B(\w3[9][101] ), .Z(out[101]) );
  XOR U5228 ( .A(key[1254]), .B(\w3[9][102] ), .Z(out[102]) );
  XOR U5229 ( .A(key[1255]), .B(\w3[9][103] ), .Z(out[103]) );
  XOR U5230 ( .A(key[1256]), .B(\w3[9][104] ), .Z(out[104]) );
  XOR U5231 ( .A(key[1257]), .B(\w3[9][105] ), .Z(out[105]) );
  XOR U5232 ( .A(key[1258]), .B(\w3[9][106] ), .Z(out[106]) );
  XOR U5233 ( .A(key[1259]), .B(\w3[9][107] ), .Z(out[107]) );
  XOR U5234 ( .A(key[1260]), .B(\w3[9][108] ), .Z(out[108]) );
  XOR U5235 ( .A(key[1261]), .B(\w3[9][109] ), .Z(out[109]) );
  XOR U5236 ( .A(key[1162]), .B(\w3[9][10] ), .Z(out[10]) );
  XOR U5237 ( .A(key[1262]), .B(\w3[9][110] ), .Z(out[110]) );
  XOR U5238 ( .A(key[1263]), .B(\w3[9][111] ), .Z(out[111]) );
  XOR U5239 ( .A(key[1264]), .B(\w3[9][112] ), .Z(out[112]) );
  XOR U5240 ( .A(key[1265]), .B(\w3[9][113] ), .Z(out[113]) );
  XOR U5241 ( .A(key[1266]), .B(\w3[9][114] ), .Z(out[114]) );
  XOR U5242 ( .A(key[1267]), .B(\w3[9][115] ), .Z(out[115]) );
  XOR U5243 ( .A(key[1268]), .B(\w3[9][116] ), .Z(out[116]) );
  XOR U5244 ( .A(key[1269]), .B(\w3[9][117] ), .Z(out[117]) );
  XOR U5245 ( .A(key[1270]), .B(\w3[9][118] ), .Z(out[118]) );
  XOR U5246 ( .A(key[1271]), .B(\w3[9][119] ), .Z(out[119]) );
  XOR U5247 ( .A(key[1163]), .B(\w3[9][11] ), .Z(out[11]) );
  XOR U5248 ( .A(key[1272]), .B(\w3[9][120] ), .Z(out[120]) );
  XOR U5249 ( .A(key[1273]), .B(\w3[9][121] ), .Z(out[121]) );
  XOR U5250 ( .A(key[1274]), .B(\w3[9][122] ), .Z(out[122]) );
  XOR U5251 ( .A(key[1275]), .B(\w3[9][123] ), .Z(out[123]) );
  XOR U5252 ( .A(key[1276]), .B(\w3[9][124] ), .Z(out[124]) );
  XOR U5253 ( .A(key[1277]), .B(\w3[9][125] ), .Z(out[125]) );
  XOR U5254 ( .A(key[1278]), .B(\w3[9][126] ), .Z(out[126]) );
  XOR U5255 ( .A(key[1279]), .B(\w3[9][127] ), .Z(out[127]) );
  XOR U5256 ( .A(key[1164]), .B(\w3[9][12] ), .Z(out[12]) );
  XOR U5257 ( .A(key[1165]), .B(\w3[9][13] ), .Z(out[13]) );
  XOR U5258 ( .A(key[1166]), .B(\w3[9][14] ), .Z(out[14]) );
  XOR U5259 ( .A(key[1167]), .B(\w3[9][15] ), .Z(out[15]) );
  XOR U5260 ( .A(key[1168]), .B(\w3[9][16] ), .Z(out[16]) );
  XOR U5261 ( .A(key[1169]), .B(\w3[9][17] ), .Z(out[17]) );
  XOR U5262 ( .A(key[1170]), .B(\w3[9][18] ), .Z(out[18]) );
  XOR U5263 ( .A(key[1171]), .B(\w3[9][19] ), .Z(out[19]) );
  XOR U5264 ( .A(key[1153]), .B(\w3[9][1] ), .Z(out[1]) );
  XOR U5265 ( .A(key[1172]), .B(\w3[9][20] ), .Z(out[20]) );
  XOR U5266 ( .A(key[1173]), .B(\w3[9][21] ), .Z(out[21]) );
  XOR U5267 ( .A(key[1174]), .B(\w3[9][22] ), .Z(out[22]) );
  XOR U5268 ( .A(key[1175]), .B(\w3[9][23] ), .Z(out[23]) );
  XOR U5269 ( .A(key[1176]), .B(\w3[9][24] ), .Z(out[24]) );
  XOR U5270 ( .A(key[1177]), .B(\w3[9][25] ), .Z(out[25]) );
  XOR U5271 ( .A(key[1178]), .B(\w3[9][26] ), .Z(out[26]) );
  XOR U5272 ( .A(key[1179]), .B(\w3[9][27] ), .Z(out[27]) );
  XOR U5273 ( .A(key[1180]), .B(\w3[9][28] ), .Z(out[28]) );
  XOR U5274 ( .A(key[1181]), .B(\w3[9][29] ), .Z(out[29]) );
  XOR U5275 ( .A(key[1154]), .B(\w3[9][2] ), .Z(out[2]) );
  XOR U5276 ( .A(key[1182]), .B(\w3[9][30] ), .Z(out[30]) );
  XOR U5277 ( .A(key[1183]), .B(\w3[9][31] ), .Z(out[31]) );
  XOR U5278 ( .A(key[1184]), .B(\w3[9][32] ), .Z(out[32]) );
  XOR U5279 ( .A(key[1185]), .B(\w3[9][33] ), .Z(out[33]) );
  XOR U5280 ( .A(key[1186]), .B(\w3[9][34] ), .Z(out[34]) );
  XOR U5281 ( .A(key[1187]), .B(\w3[9][35] ), .Z(out[35]) );
  XOR U5282 ( .A(key[1188]), .B(\w3[9][36] ), .Z(out[36]) );
  XOR U5283 ( .A(key[1189]), .B(\w3[9][37] ), .Z(out[37]) );
  XOR U5284 ( .A(key[1190]), .B(\w3[9][38] ), .Z(out[38]) );
  XOR U5285 ( .A(key[1191]), .B(\w3[9][39] ), .Z(out[39]) );
  XOR U5286 ( .A(key[1155]), .B(\w3[9][3] ), .Z(out[3]) );
  XOR U5287 ( .A(key[1192]), .B(\w3[9][40] ), .Z(out[40]) );
  XOR U5288 ( .A(key[1193]), .B(\w3[9][41] ), .Z(out[41]) );
  XOR U5289 ( .A(key[1194]), .B(\w3[9][42] ), .Z(out[42]) );
  XOR U5290 ( .A(key[1195]), .B(\w3[9][43] ), .Z(out[43]) );
  XOR U5291 ( .A(key[1196]), .B(\w3[9][44] ), .Z(out[44]) );
  XOR U5292 ( .A(key[1197]), .B(\w3[9][45] ), .Z(out[45]) );
  XOR U5293 ( .A(key[1198]), .B(\w3[9][46] ), .Z(out[46]) );
  XOR U5294 ( .A(key[1199]), .B(\w3[9][47] ), .Z(out[47]) );
  XOR U5295 ( .A(key[1200]), .B(\w3[9][48] ), .Z(out[48]) );
  XOR U5296 ( .A(key[1201]), .B(\w3[9][49] ), .Z(out[49]) );
  XOR U5297 ( .A(key[1156]), .B(\w3[9][4] ), .Z(out[4]) );
  XOR U5298 ( .A(key[1202]), .B(\w3[9][50] ), .Z(out[50]) );
  XOR U5299 ( .A(key[1203]), .B(\w3[9][51] ), .Z(out[51]) );
  XOR U5300 ( .A(key[1204]), .B(\w3[9][52] ), .Z(out[52]) );
  XOR U5301 ( .A(key[1205]), .B(\w3[9][53] ), .Z(out[53]) );
  XOR U5302 ( .A(key[1206]), .B(\w3[9][54] ), .Z(out[54]) );
  XOR U5303 ( .A(key[1207]), .B(\w3[9][55] ), .Z(out[55]) );
  XOR U5304 ( .A(key[1208]), .B(\w3[9][56] ), .Z(out[56]) );
  XOR U5305 ( .A(key[1209]), .B(\w3[9][57] ), .Z(out[57]) );
  XOR U5306 ( .A(key[1210]), .B(\w3[9][58] ), .Z(out[58]) );
  XOR U5307 ( .A(key[1211]), .B(\w3[9][59] ), .Z(out[59]) );
  XOR U5308 ( .A(key[1157]), .B(\w3[9][5] ), .Z(out[5]) );
  XOR U5309 ( .A(key[1212]), .B(\w3[9][60] ), .Z(out[60]) );
  XOR U5310 ( .A(key[1213]), .B(\w3[9][61] ), .Z(out[61]) );
  XOR U5311 ( .A(key[1214]), .B(\w3[9][62] ), .Z(out[62]) );
  XOR U5312 ( .A(key[1215]), .B(\w3[9][63] ), .Z(out[63]) );
  XOR U5313 ( .A(key[1216]), .B(\w3[9][64] ), .Z(out[64]) );
  XOR U5314 ( .A(key[1217]), .B(\w3[9][65] ), .Z(out[65]) );
  XOR U5315 ( .A(key[1218]), .B(\w3[9][66] ), .Z(out[66]) );
  XOR U5316 ( .A(key[1219]), .B(\w3[9][67] ), .Z(out[67]) );
  XOR U5317 ( .A(key[1220]), .B(\w3[9][68] ), .Z(out[68]) );
  XOR U5318 ( .A(key[1221]), .B(\w3[9][69] ), .Z(out[69]) );
  XOR U5319 ( .A(key[1158]), .B(\w3[9][6] ), .Z(out[6]) );
  XOR U5320 ( .A(key[1222]), .B(\w3[9][70] ), .Z(out[70]) );
  XOR U5321 ( .A(key[1223]), .B(\w3[9][71] ), .Z(out[71]) );
  XOR U5322 ( .A(key[1224]), .B(\w3[9][72] ), .Z(out[72]) );
  XOR U5323 ( .A(key[1225]), .B(\w3[9][73] ), .Z(out[73]) );
  XOR U5324 ( .A(key[1226]), .B(\w3[9][74] ), .Z(out[74]) );
  XOR U5325 ( .A(key[1227]), .B(\w3[9][75] ), .Z(out[75]) );
  XOR U5326 ( .A(key[1228]), .B(\w3[9][76] ), .Z(out[76]) );
  XOR U5327 ( .A(key[1229]), .B(\w3[9][77] ), .Z(out[77]) );
  XOR U5328 ( .A(key[1230]), .B(\w3[9][78] ), .Z(out[78]) );
  XOR U5329 ( .A(key[1231]), .B(\w3[9][79] ), .Z(out[79]) );
  XOR U5330 ( .A(key[1159]), .B(\w3[9][7] ), .Z(out[7]) );
  XOR U5331 ( .A(key[1232]), .B(\w3[9][80] ), .Z(out[80]) );
  XOR U5332 ( .A(key[1233]), .B(\w3[9][81] ), .Z(out[81]) );
  XOR U5333 ( .A(key[1234]), .B(\w3[9][82] ), .Z(out[82]) );
  XOR U5334 ( .A(key[1235]), .B(\w3[9][83] ), .Z(out[83]) );
  XOR U5335 ( .A(key[1236]), .B(\w3[9][84] ), .Z(out[84]) );
  XOR U5336 ( .A(key[1237]), .B(\w3[9][85] ), .Z(out[85]) );
  XOR U5337 ( .A(key[1238]), .B(\w3[9][86] ), .Z(out[86]) );
  XOR U5338 ( .A(key[1239]), .B(\w3[9][87] ), .Z(out[87]) );
  XOR U5339 ( .A(key[1240]), .B(\w3[9][88] ), .Z(out[88]) );
  XOR U5340 ( .A(key[1241]), .B(\w3[9][89] ), .Z(out[89]) );
  XOR U5341 ( .A(key[1160]), .B(\w3[9][8] ), .Z(out[8]) );
  XOR U5342 ( .A(key[1242]), .B(\w3[9][90] ), .Z(out[90]) );
  XOR U5343 ( .A(key[1243]), .B(\w3[9][91] ), .Z(out[91]) );
  XOR U5344 ( .A(key[1244]), .B(\w3[9][92] ), .Z(out[92]) );
  XOR U5345 ( .A(key[1245]), .B(\w3[9][93] ), .Z(out[93]) );
  XOR U5346 ( .A(key[1246]), .B(\w3[9][94] ), .Z(out[94]) );
  XOR U5347 ( .A(key[1247]), .B(\w3[9][95] ), .Z(out[95]) );
  XOR U5348 ( .A(key[1248]), .B(\w3[9][96] ), .Z(out[96]) );
  XOR U5349 ( .A(key[1249]), .B(\w3[9][97] ), .Z(out[97]) );
  XOR U5350 ( .A(key[1250]), .B(\w3[9][98] ), .Z(out[98]) );
  XOR U5351 ( .A(key[1251]), .B(\w3[9][99] ), .Z(out[99]) );
  XOR U5352 ( .A(key[1161]), .B(\w3[9][9] ), .Z(out[9]) );
  XOR U5353 ( .A(key[0]), .B(msg[0]), .Z(\w1[0][0] ) );
  XOR U5354 ( .A(key[100]), .B(msg[100]), .Z(\w1[0][100] ) );
  XOR U5355 ( .A(key[101]), .B(msg[101]), .Z(\w1[0][101] ) );
  XOR U5356 ( .A(key[102]), .B(msg[102]), .Z(\w1[0][102] ) );
  XOR U5357 ( .A(key[103]), .B(msg[103]), .Z(\w1[0][103] ) );
  XOR U5358 ( .A(key[104]), .B(msg[104]), .Z(\w1[0][104] ) );
  XOR U5359 ( .A(key[105]), .B(msg[105]), .Z(\w1[0][105] ) );
  XOR U5360 ( .A(key[106]), .B(msg[106]), .Z(\w1[0][106] ) );
  XOR U5361 ( .A(key[107]), .B(msg[107]), .Z(\w1[0][107] ) );
  XOR U5362 ( .A(key[108]), .B(msg[108]), .Z(\w1[0][108] ) );
  XOR U5363 ( .A(key[109]), .B(msg[109]), .Z(\w1[0][109] ) );
  XOR U5364 ( .A(key[10]), .B(msg[10]), .Z(\w1[0][10] ) );
  XOR U5365 ( .A(key[110]), .B(msg[110]), .Z(\w1[0][110] ) );
  XOR U5366 ( .A(key[111]), .B(msg[111]), .Z(\w1[0][111] ) );
  XOR U5367 ( .A(key[112]), .B(msg[112]), .Z(\w1[0][112] ) );
  XOR U5368 ( .A(key[113]), .B(msg[113]), .Z(\w1[0][113] ) );
  XOR U5369 ( .A(key[114]), .B(msg[114]), .Z(\w1[0][114] ) );
  XOR U5370 ( .A(key[115]), .B(msg[115]), .Z(\w1[0][115] ) );
  XOR U5371 ( .A(key[116]), .B(msg[116]), .Z(\w1[0][116] ) );
  XOR U5372 ( .A(key[117]), .B(msg[117]), .Z(\w1[0][117] ) );
  XOR U5373 ( .A(key[118]), .B(msg[118]), .Z(\w1[0][118] ) );
  XOR U5374 ( .A(key[119]), .B(msg[119]), .Z(\w1[0][119] ) );
  XOR U5375 ( .A(key[11]), .B(msg[11]), .Z(\w1[0][11] ) );
  XOR U5376 ( .A(key[120]), .B(msg[120]), .Z(\w1[0][120] ) );
  XOR U5377 ( .A(key[121]), .B(msg[121]), .Z(\w1[0][121] ) );
  XOR U5378 ( .A(key[122]), .B(msg[122]), .Z(\w1[0][122] ) );
  XOR U5379 ( .A(key[123]), .B(msg[123]), .Z(\w1[0][123] ) );
  XOR U5380 ( .A(key[124]), .B(msg[124]), .Z(\w1[0][124] ) );
  XOR U5381 ( .A(key[125]), .B(msg[125]), .Z(\w1[0][125] ) );
  XOR U5382 ( .A(key[126]), .B(msg[126]), .Z(\w1[0][126] ) );
  XOR U5383 ( .A(key[127]), .B(msg[127]), .Z(\w1[0][127] ) );
  XOR U5384 ( .A(key[12]), .B(msg[12]), .Z(\w1[0][12] ) );
  XOR U5385 ( .A(key[13]), .B(msg[13]), .Z(\w1[0][13] ) );
  XOR U5386 ( .A(key[14]), .B(msg[14]), .Z(\w1[0][14] ) );
  XOR U5387 ( .A(key[15]), .B(msg[15]), .Z(\w1[0][15] ) );
  XOR U5388 ( .A(key[16]), .B(msg[16]), .Z(\w1[0][16] ) );
  XOR U5389 ( .A(key[17]), .B(msg[17]), .Z(\w1[0][17] ) );
  XOR U5390 ( .A(key[18]), .B(msg[18]), .Z(\w1[0][18] ) );
  XOR U5391 ( .A(key[19]), .B(msg[19]), .Z(\w1[0][19] ) );
  XOR U5392 ( .A(key[1]), .B(msg[1]), .Z(\w1[0][1] ) );
  XOR U5393 ( .A(key[20]), .B(msg[20]), .Z(\w1[0][20] ) );
  XOR U5394 ( .A(key[21]), .B(msg[21]), .Z(\w1[0][21] ) );
  XOR U5395 ( .A(key[22]), .B(msg[22]), .Z(\w1[0][22] ) );
  XOR U5396 ( .A(key[23]), .B(msg[23]), .Z(\w1[0][23] ) );
  XOR U5397 ( .A(key[24]), .B(msg[24]), .Z(\w1[0][24] ) );
  XOR U5398 ( .A(key[25]), .B(msg[25]), .Z(\w1[0][25] ) );
  XOR U5399 ( .A(key[26]), .B(msg[26]), .Z(\w1[0][26] ) );
  XOR U5400 ( .A(key[27]), .B(msg[27]), .Z(\w1[0][27] ) );
  XOR U5401 ( .A(key[28]), .B(msg[28]), .Z(\w1[0][28] ) );
  XOR U5402 ( .A(key[29]), .B(msg[29]), .Z(\w1[0][29] ) );
  XOR U5403 ( .A(key[2]), .B(msg[2]), .Z(\w1[0][2] ) );
  XOR U5404 ( .A(key[30]), .B(msg[30]), .Z(\w1[0][30] ) );
  XOR U5405 ( .A(key[31]), .B(msg[31]), .Z(\w1[0][31] ) );
  XOR U5406 ( .A(key[32]), .B(msg[32]), .Z(\w1[0][32] ) );
  XOR U5407 ( .A(key[33]), .B(msg[33]), .Z(\w1[0][33] ) );
  XOR U5408 ( .A(key[34]), .B(msg[34]), .Z(\w1[0][34] ) );
  XOR U5409 ( .A(key[35]), .B(msg[35]), .Z(\w1[0][35] ) );
  XOR U5410 ( .A(key[36]), .B(msg[36]), .Z(\w1[0][36] ) );
  XOR U5411 ( .A(key[37]), .B(msg[37]), .Z(\w1[0][37] ) );
  XOR U5412 ( .A(key[38]), .B(msg[38]), .Z(\w1[0][38] ) );
  XOR U5413 ( .A(key[39]), .B(msg[39]), .Z(\w1[0][39] ) );
  XOR U5414 ( .A(key[3]), .B(msg[3]), .Z(\w1[0][3] ) );
  XOR U5415 ( .A(key[40]), .B(msg[40]), .Z(\w1[0][40] ) );
  XOR U5416 ( .A(key[41]), .B(msg[41]), .Z(\w1[0][41] ) );
  XOR U5417 ( .A(key[42]), .B(msg[42]), .Z(\w1[0][42] ) );
  XOR U5418 ( .A(key[43]), .B(msg[43]), .Z(\w1[0][43] ) );
  XOR U5419 ( .A(key[44]), .B(msg[44]), .Z(\w1[0][44] ) );
  XOR U5420 ( .A(key[45]), .B(msg[45]), .Z(\w1[0][45] ) );
  XOR U5421 ( .A(key[46]), .B(msg[46]), .Z(\w1[0][46] ) );
  XOR U5422 ( .A(key[47]), .B(msg[47]), .Z(\w1[0][47] ) );
  XOR U5423 ( .A(key[48]), .B(msg[48]), .Z(\w1[0][48] ) );
  XOR U5424 ( .A(key[49]), .B(msg[49]), .Z(\w1[0][49] ) );
  XOR U5425 ( .A(key[4]), .B(msg[4]), .Z(\w1[0][4] ) );
  XOR U5426 ( .A(key[50]), .B(msg[50]), .Z(\w1[0][50] ) );
  XOR U5427 ( .A(key[51]), .B(msg[51]), .Z(\w1[0][51] ) );
  XOR U5428 ( .A(key[52]), .B(msg[52]), .Z(\w1[0][52] ) );
  XOR U5429 ( .A(key[53]), .B(msg[53]), .Z(\w1[0][53] ) );
  XOR U5430 ( .A(key[54]), .B(msg[54]), .Z(\w1[0][54] ) );
  XOR U5431 ( .A(key[55]), .B(msg[55]), .Z(\w1[0][55] ) );
  XOR U5432 ( .A(key[56]), .B(msg[56]), .Z(\w1[0][56] ) );
  XOR U5433 ( .A(key[57]), .B(msg[57]), .Z(\w1[0][57] ) );
  XOR U5434 ( .A(key[58]), .B(msg[58]), .Z(\w1[0][58] ) );
  XOR U5435 ( .A(key[59]), .B(msg[59]), .Z(\w1[0][59] ) );
  XOR U5436 ( .A(key[5]), .B(msg[5]), .Z(\w1[0][5] ) );
  XOR U5437 ( .A(key[60]), .B(msg[60]), .Z(\w1[0][60] ) );
  XOR U5438 ( .A(key[61]), .B(msg[61]), .Z(\w1[0][61] ) );
  XOR U5439 ( .A(key[62]), .B(msg[62]), .Z(\w1[0][62] ) );
  XOR U5440 ( .A(key[63]), .B(msg[63]), .Z(\w1[0][63] ) );
  XOR U5441 ( .A(key[64]), .B(msg[64]), .Z(\w1[0][64] ) );
  XOR U5442 ( .A(key[65]), .B(msg[65]), .Z(\w1[0][65] ) );
  XOR U5443 ( .A(key[66]), .B(msg[66]), .Z(\w1[0][66] ) );
  XOR U5444 ( .A(key[67]), .B(msg[67]), .Z(\w1[0][67] ) );
  XOR U5445 ( .A(key[68]), .B(msg[68]), .Z(\w1[0][68] ) );
  XOR U5446 ( .A(key[69]), .B(msg[69]), .Z(\w1[0][69] ) );
  XOR U5447 ( .A(key[6]), .B(msg[6]), .Z(\w1[0][6] ) );
  XOR U5448 ( .A(key[70]), .B(msg[70]), .Z(\w1[0][70] ) );
  XOR U5449 ( .A(key[71]), .B(msg[71]), .Z(\w1[0][71] ) );
  XOR U5450 ( .A(key[72]), .B(msg[72]), .Z(\w1[0][72] ) );
  XOR U5451 ( .A(key[73]), .B(msg[73]), .Z(\w1[0][73] ) );
  XOR U5452 ( .A(key[74]), .B(msg[74]), .Z(\w1[0][74] ) );
  XOR U5453 ( .A(key[75]), .B(msg[75]), .Z(\w1[0][75] ) );
  XOR U5454 ( .A(key[76]), .B(msg[76]), .Z(\w1[0][76] ) );
  XOR U5455 ( .A(key[77]), .B(msg[77]), .Z(\w1[0][77] ) );
  XOR U5456 ( .A(key[78]), .B(msg[78]), .Z(\w1[0][78] ) );
  XOR U5457 ( .A(key[79]), .B(msg[79]), .Z(\w1[0][79] ) );
  XOR U5458 ( .A(key[7]), .B(msg[7]), .Z(\w1[0][7] ) );
  XOR U5459 ( .A(key[80]), .B(msg[80]), .Z(\w1[0][80] ) );
  XOR U5460 ( .A(key[81]), .B(msg[81]), .Z(\w1[0][81] ) );
  XOR U5461 ( .A(key[82]), .B(msg[82]), .Z(\w1[0][82] ) );
  XOR U5462 ( .A(key[83]), .B(msg[83]), .Z(\w1[0][83] ) );
  XOR U5463 ( .A(key[84]), .B(msg[84]), .Z(\w1[0][84] ) );
  XOR U5464 ( .A(key[85]), .B(msg[85]), .Z(\w1[0][85] ) );
  XOR U5465 ( .A(key[86]), .B(msg[86]), .Z(\w1[0][86] ) );
  XOR U5466 ( .A(key[87]), .B(msg[87]), .Z(\w1[0][87] ) );
  XOR U5467 ( .A(key[88]), .B(msg[88]), .Z(\w1[0][88] ) );
  XOR U5468 ( .A(key[89]), .B(msg[89]), .Z(\w1[0][89] ) );
  XOR U5469 ( .A(key[8]), .B(msg[8]), .Z(\w1[0][8] ) );
  XOR U5470 ( .A(key[90]), .B(msg[90]), .Z(\w1[0][90] ) );
  XOR U5471 ( .A(key[91]), .B(msg[91]), .Z(\w1[0][91] ) );
  XOR U5472 ( .A(key[92]), .B(msg[92]), .Z(\w1[0][92] ) );
  XOR U5473 ( .A(key[93]), .B(msg[93]), .Z(\w1[0][93] ) );
  XOR U5474 ( .A(key[94]), .B(msg[94]), .Z(\w1[0][94] ) );
  XOR U5475 ( .A(key[95]), .B(msg[95]), .Z(\w1[0][95] ) );
  XOR U5476 ( .A(key[96]), .B(msg[96]), .Z(\w1[0][96] ) );
  XOR U5477 ( .A(key[97]), .B(msg[97]), .Z(\w1[0][97] ) );
  XOR U5478 ( .A(key[98]), .B(msg[98]), .Z(\w1[0][98] ) );
  XOR U5479 ( .A(key[99]), .B(msg[99]), .Z(\w1[0][99] ) );
  XOR U5480 ( .A(key[9]), .B(msg[9]), .Z(\w1[0][9] ) );
  XOR U5481 ( .A(\w3[0][8] ), .B(key[128]), .Z(n3818) );
  XOR U5482 ( .A(\w3[0][1] ), .B(\w3[0][25] ), .Z(n4240) );
  XOR U5483 ( .A(\w3[0][16] ), .B(\w3[0][24] ), .Z(n4196) );
  XNOR U5484 ( .A(n4240), .B(n4196), .Z(n3817) );
  XNOR U5485 ( .A(n3818), .B(n3817), .Z(\w1[1][0] ) );
  XOR U5486 ( .A(\w3[0][96] ), .B(\w3[0][101] ), .Z(n3844) );
  XOR U5487 ( .A(n3844), .B(key[228]), .Z(n3822) );
  XOR U5488 ( .A(\w3[0][116] ), .B(\w3[0][125] ), .Z(n3820) );
  XNOR U5489 ( .A(\w3[0][120] ), .B(\w3[0][108] ), .Z(n3819) );
  XNOR U5490 ( .A(n3820), .B(n3819), .Z(n3901) );
  XNOR U5491 ( .A(\w3[0][124] ), .B(n3901), .Z(n3821) );
  XNOR U5492 ( .A(n3822), .B(n3821), .Z(\w1[1][100] ) );
  XOR U5493 ( .A(\w3[0][102] ), .B(\w3[0][126] ), .Z(n3853) );
  XOR U5494 ( .A(n3853), .B(key[229]), .Z(n3824) );
  XOR U5495 ( .A(\w3[0][109] ), .B(\w3[0][117] ), .Z(n3904) );
  XNOR U5496 ( .A(\w3[0][125] ), .B(n3904), .Z(n3823) );
  XNOR U5497 ( .A(n3824), .B(n3823), .Z(\w1[1][101] ) );
  XOR U5498 ( .A(\w3[0][96] ), .B(\w3[0][103] ), .Z(n3854) );
  XOR U5499 ( .A(n3854), .B(key[230]), .Z(n3826) );
  XOR U5500 ( .A(\w3[0][110] ), .B(\w3[0][118] ), .Z(n3872) );
  XNOR U5501 ( .A(\w3[0][120] ), .B(\w3[0][127] ), .Z(n3828) );
  XNOR U5502 ( .A(n3872), .B(n3828), .Z(n3909) );
  XNOR U5503 ( .A(\w3[0][126] ), .B(n3909), .Z(n3825) );
  XNOR U5504 ( .A(n3826), .B(n3825), .Z(\w1[1][102] ) );
  XOR U5505 ( .A(\w3[0][111] ), .B(\w3[0][119] ), .Z(n3912) );
  XNOR U5506 ( .A(n3912), .B(key[231]), .Z(n3827) );
  XNOR U5507 ( .A(n3828), .B(n3827), .Z(n3829) );
  XNOR U5508 ( .A(\w3[0][96] ), .B(n3829), .Z(\w1[1][103] ) );
  XOR U5509 ( .A(key[232]), .B(\w3[0][105] ), .Z(n3831) );
  XNOR U5510 ( .A(\w3[0][96] ), .B(\w3[0][97] ), .Z(n3830) );
  XNOR U5511 ( .A(n3831), .B(n3830), .Z(n3832) );
  XNOR U5512 ( .A(\w3[0][120] ), .B(\w3[0][112] ), .Z(n4222) );
  XNOR U5513 ( .A(n3832), .B(n4222), .Z(\w1[1][104] ) );
  XOR U5514 ( .A(\w3[0][106] ), .B(\w3[0][113] ), .Z(n3834) );
  XOR U5515 ( .A(\w3[0][97] ), .B(\w3[0][121] ), .Z(n4221) );
  XNOR U5516 ( .A(n4221), .B(key[233]), .Z(n3833) );
  XNOR U5517 ( .A(n3834), .B(n3833), .Z(n3835) );
  XOR U5518 ( .A(\w3[0][98] ), .B(n3835), .Z(\w1[1][105] ) );
  XOR U5519 ( .A(\w3[0][107] ), .B(\w3[0][114] ), .Z(n3837) );
  XOR U5520 ( .A(\w3[0][98] ), .B(\w3[0][122] ), .Z(n4226) );
  XNOR U5521 ( .A(n4226), .B(key[234]), .Z(n3836) );
  XNOR U5522 ( .A(n3837), .B(n3836), .Z(n3838) );
  XOR U5523 ( .A(\w3[0][99] ), .B(n3838), .Z(\w1[1][106] ) );
  XOR U5524 ( .A(\w3[0][99] ), .B(\w3[0][123] ), .Z(n4230) );
  XNOR U5525 ( .A(\w3[0][108] ), .B(n4230), .Z(n3839) );
  XNOR U5526 ( .A(\w3[0][104] ), .B(n3839), .Z(n3865) );
  XOR U5527 ( .A(n3865), .B(key[235]), .Z(n3841) );
  XOR U5528 ( .A(\w3[0][96] ), .B(\w3[0][100] ), .Z(n4234) );
  XNOR U5529 ( .A(\w3[0][115] ), .B(n4234), .Z(n3840) );
  XNOR U5530 ( .A(n3841), .B(n3840), .Z(\w1[1][107] ) );
  XOR U5531 ( .A(\w3[0][100] ), .B(\w3[0][104] ), .Z(n3843) );
  XNOR U5532 ( .A(\w3[0][124] ), .B(\w3[0][109] ), .Z(n3842) );
  XNOR U5533 ( .A(n3843), .B(n3842), .Z(n3868) );
  XOR U5534 ( .A(n3868), .B(key[236]), .Z(n3846) );
  XNOR U5535 ( .A(\w3[0][116] ), .B(n3844), .Z(n3845) );
  XNOR U5536 ( .A(n3846), .B(n3845), .Z(\w1[1][108] ) );
  XOR U5537 ( .A(\w3[0][125] ), .B(\w3[0][101] ), .Z(n3871) );
  XOR U5538 ( .A(n3871), .B(key[237]), .Z(n3848) );
  XNOR U5539 ( .A(\w3[0][102] ), .B(\w3[0][110] ), .Z(n3847) );
  XNOR U5540 ( .A(n3848), .B(n3847), .Z(n3849) );
  XOR U5541 ( .A(\w3[0][117] ), .B(n3849), .Z(\w1[1][109] ) );
  XOR U5542 ( .A(\w3[0][11] ), .B(\w3[0][18] ), .Z(n3851) );
  XOR U5543 ( .A(\w3[0][2] ), .B(\w3[0][26] ), .Z(n3935) );
  XNOR U5544 ( .A(n3935), .B(key[138]), .Z(n3850) );
  XNOR U5545 ( .A(n3851), .B(n3850), .Z(n3852) );
  XOR U5546 ( .A(\w3[0][3] ), .B(n3852), .Z(\w1[1][10] ) );
  XNOR U5547 ( .A(\w3[0][111] ), .B(\w3[0][104] ), .Z(n3880) );
  XNOR U5548 ( .A(n3853), .B(n3880), .Z(n3875) );
  XOR U5549 ( .A(n3875), .B(key[238]), .Z(n3856) );
  XNOR U5550 ( .A(\w3[0][118] ), .B(n3854), .Z(n3855) );
  XNOR U5551 ( .A(n3856), .B(n3855), .Z(\w1[1][110] ) );
  XOR U5552 ( .A(\w3[0][127] ), .B(\w3[0][103] ), .Z(n3878) );
  XOR U5553 ( .A(n3878), .B(key[239]), .Z(n3858) );
  XOR U5554 ( .A(\w3[0][96] ), .B(\w3[0][104] ), .Z(n3885) );
  XNOR U5555 ( .A(\w3[0][119] ), .B(n3885), .Z(n3857) );
  XNOR U5556 ( .A(n3858), .B(n3857), .Z(\w1[1][111] ) );
  XOR U5557 ( .A(\w3[0][105] ), .B(\w3[0][113] ), .Z(n4225) );
  XOR U5558 ( .A(n4225), .B(key[240]), .Z(n3860) );
  XNOR U5559 ( .A(\w3[0][120] ), .B(n3885), .Z(n3859) );
  XNOR U5560 ( .A(n3860), .B(n3859), .Z(\w1[1][112] ) );
  XOR U5561 ( .A(\w3[0][106] ), .B(\w3[0][114] ), .Z(n4229) );
  XOR U5562 ( .A(n4229), .B(key[241]), .Z(n3862) );
  XNOR U5563 ( .A(\w3[0][105] ), .B(n4221), .Z(n3861) );
  XNOR U5564 ( .A(n3862), .B(n3861), .Z(\w1[1][113] ) );
  XOR U5565 ( .A(\w3[0][107] ), .B(\w3[0][115] ), .Z(n3896) );
  XOR U5566 ( .A(n3896), .B(key[242]), .Z(n3864) );
  XNOR U5567 ( .A(\w3[0][106] ), .B(n4226), .Z(n3863) );
  XNOR U5568 ( .A(n3864), .B(n3863), .Z(\w1[1][114] ) );
  XOR U5569 ( .A(\w3[0][116] ), .B(\w3[0][112] ), .Z(n3897) );
  XOR U5570 ( .A(n3897), .B(key[243]), .Z(n3867) );
  XNOR U5571 ( .A(\w3[0][107] ), .B(n3865), .Z(n3866) );
  XNOR U5572 ( .A(n3867), .B(n3866), .Z(\w1[1][115] ) );
  XOR U5573 ( .A(\w3[0][117] ), .B(\w3[0][112] ), .Z(n3900) );
  XOR U5574 ( .A(n3900), .B(key[244]), .Z(n3870) );
  XNOR U5575 ( .A(\w3[0][108] ), .B(n3868), .Z(n3869) );
  XNOR U5576 ( .A(n3870), .B(n3869), .Z(\w1[1][116] ) );
  XOR U5577 ( .A(n3871), .B(key[245]), .Z(n3874) );
  XNOR U5578 ( .A(\w3[0][109] ), .B(n3872), .Z(n3873) );
  XNOR U5579 ( .A(n3874), .B(n3873), .Z(\w1[1][117] ) );
  XOR U5580 ( .A(\w3[0][119] ), .B(\w3[0][112] ), .Z(n3908) );
  XOR U5581 ( .A(n3908), .B(key[246]), .Z(n3877) );
  XNOR U5582 ( .A(\w3[0][110] ), .B(n3875), .Z(n3876) );
  XNOR U5583 ( .A(n3877), .B(n3876), .Z(\w1[1][118] ) );
  XNOR U5584 ( .A(n3878), .B(key[247]), .Z(n3879) );
  XNOR U5585 ( .A(n3880), .B(n3879), .Z(n3881) );
  XNOR U5586 ( .A(\w3[0][112] ), .B(n3881), .Z(\w1[1][119] ) );
  XOR U5587 ( .A(\w3[0][3] ), .B(\w3[0][27] ), .Z(n3976) );
  XNOR U5588 ( .A(\w3[0][8] ), .B(\w3[0][12] ), .Z(n3882) );
  XNOR U5589 ( .A(n3976), .B(n3882), .Z(n3932) );
  XOR U5590 ( .A(n3932), .B(key[139]), .Z(n3884) );
  XOR U5591 ( .A(\w3[0][0] ), .B(\w3[0][4] ), .Z(n4006) );
  XNOR U5592 ( .A(\w3[0][19] ), .B(n4006), .Z(n3883) );
  XNOR U5593 ( .A(n3884), .B(n3883), .Z(\w1[1][11] ) );
  XOR U5594 ( .A(n3885), .B(key[248]), .Z(n3887) );
  XNOR U5595 ( .A(\w3[0][121] ), .B(\w3[0][113] ), .Z(n3886) );
  XNOR U5596 ( .A(n3887), .B(n3886), .Z(n3888) );
  XOR U5597 ( .A(\w3[0][112] ), .B(n3888), .Z(\w1[1][120] ) );
  XOR U5598 ( .A(n4225), .B(key[249]), .Z(n3890) );
  XNOR U5599 ( .A(\w3[0][122] ), .B(\w3[0][114] ), .Z(n3889) );
  XNOR U5600 ( .A(n3890), .B(n3889), .Z(n3891) );
  XOR U5601 ( .A(\w3[0][97] ), .B(n3891), .Z(\w1[1][121] ) );
  XOR U5602 ( .A(n4229), .B(key[250]), .Z(n3893) );
  XNOR U5603 ( .A(\w3[0][115] ), .B(\w3[0][123] ), .Z(n3892) );
  XNOR U5604 ( .A(n3893), .B(n3892), .Z(n3894) );
  XOR U5605 ( .A(\w3[0][98] ), .B(n3894), .Z(\w1[1][122] ) );
  XNOR U5606 ( .A(\w3[0][124] ), .B(\w3[0][120] ), .Z(n3895) );
  XNOR U5607 ( .A(n3896), .B(n3895), .Z(n4233) );
  XOR U5608 ( .A(n4233), .B(key[251]), .Z(n3899) );
  XNOR U5609 ( .A(\w3[0][99] ), .B(n3897), .Z(n3898) );
  XNOR U5610 ( .A(n3899), .B(n3898), .Z(\w1[1][123] ) );
  XOR U5611 ( .A(n3900), .B(key[252]), .Z(n3903) );
  XNOR U5612 ( .A(n3901), .B(\w3[0][100] ), .Z(n3902) );
  XNOR U5613 ( .A(n3903), .B(n3902), .Z(\w1[1][124] ) );
  XOR U5614 ( .A(\w3[0][118] ), .B(key[253]), .Z(n3906) );
  XNOR U5615 ( .A(n3904), .B(\w3[0][126] ), .Z(n3905) );
  XNOR U5616 ( .A(n3906), .B(n3905), .Z(n3907) );
  XOR U5617 ( .A(\w3[0][101] ), .B(n3907), .Z(\w1[1][125] ) );
  XOR U5618 ( .A(n3908), .B(key[254]), .Z(n3911) );
  XNOR U5619 ( .A(\w3[0][102] ), .B(n3909), .Z(n3910) );
  XNOR U5620 ( .A(n3911), .B(n3910), .Z(\w1[1][126] ) );
  XNOR U5621 ( .A(n3912), .B(key[255]), .Z(n3913) );
  XNOR U5622 ( .A(n4222), .B(n3913), .Z(n3914) );
  XNOR U5623 ( .A(\w3[0][103] ), .B(n3914), .Z(\w1[1][127] ) );
  XOR U5624 ( .A(\w3[0][13] ), .B(\w3[0][28] ), .Z(n3916) );
  XNOR U5625 ( .A(\w3[0][8] ), .B(\w3[0][4] ), .Z(n3915) );
  XNOR U5626 ( .A(n3916), .B(n3915), .Z(n3938) );
  XOR U5627 ( .A(n3938), .B(key[140]), .Z(n3918) );
  XOR U5628 ( .A(\w3[0][0] ), .B(\w3[0][5] ), .Z(n4043) );
  XNOR U5629 ( .A(\w3[0][20] ), .B(n4043), .Z(n3917) );
  XNOR U5630 ( .A(n3918), .B(n3917), .Z(\w1[1][12] ) );
  XOR U5631 ( .A(\w3[0][14] ), .B(\w3[0][6] ), .Z(n3920) );
  XOR U5632 ( .A(\w3[0][5] ), .B(\w3[0][29] ), .Z(n3941) );
  XNOR U5633 ( .A(n3941), .B(key[141]), .Z(n3919) );
  XNOR U5634 ( .A(n3920), .B(n3919), .Z(n3921) );
  XOR U5635 ( .A(\w3[0][21] ), .B(n3921), .Z(\w1[1][13] ) );
  XOR U5636 ( .A(\w3[0][6] ), .B(\w3[0][30] ), .Z(n4084) );
  XNOR U5637 ( .A(\w3[0][8] ), .B(\w3[0][15] ), .Z(n3949) );
  XNOR U5638 ( .A(n4084), .B(n3949), .Z(n3944) );
  XOR U5639 ( .A(n3944), .B(key[142]), .Z(n3923) );
  XOR U5640 ( .A(\w3[0][0] ), .B(\w3[0][7] ), .Z(n4119) );
  XNOR U5641 ( .A(\w3[0][22] ), .B(n4119), .Z(n3922) );
  XNOR U5642 ( .A(n3923), .B(n3922), .Z(\w1[1][14] ) );
  XOR U5643 ( .A(\w3[0][7] ), .B(\w3[0][31] ), .Z(n3947) );
  XOR U5644 ( .A(n3947), .B(key[143]), .Z(n3925) );
  XOR U5645 ( .A(\w3[0][8] ), .B(\w3[0][0] ), .Z(n3951) );
  XNOR U5646 ( .A(\w3[0][23] ), .B(n3951), .Z(n3924) );
  XNOR U5647 ( .A(n3925), .B(n3924), .Z(\w1[1][15] ) );
  XOR U5648 ( .A(\w3[0][17] ), .B(\w3[0][9] ), .Z(n3955) );
  XOR U5649 ( .A(n3955), .B(key[144]), .Z(n3927) );
  XNOR U5650 ( .A(\w3[0][24] ), .B(n3951), .Z(n3926) );
  XNOR U5651 ( .A(n3927), .B(n3926), .Z(\w1[1][16] ) );
  XOR U5652 ( .A(\w3[0][18] ), .B(\w3[0][10] ), .Z(n3975) );
  XOR U5653 ( .A(n3975), .B(key[145]), .Z(n3929) );
  XNOR U5654 ( .A(n4240), .B(\w3[0][9] ), .Z(n3928) );
  XNOR U5655 ( .A(n3929), .B(n3928), .Z(\w1[1][17] ) );
  XOR U5656 ( .A(\w3[0][11] ), .B(\w3[0][19] ), .Z(n3963) );
  XOR U5657 ( .A(n3963), .B(key[146]), .Z(n3931) );
  XNOR U5658 ( .A(n3935), .B(\w3[0][10] ), .Z(n3930) );
  XNOR U5659 ( .A(n3931), .B(n3930), .Z(\w1[1][18] ) );
  XOR U5660 ( .A(\w3[0][16] ), .B(\w3[0][20] ), .Z(n3964) );
  XOR U5661 ( .A(n3964), .B(key[147]), .Z(n3934) );
  XNOR U5662 ( .A(\w3[0][11] ), .B(n3932), .Z(n3933) );
  XNOR U5663 ( .A(n3934), .B(n3933), .Z(\w1[1][19] ) );
  XOR U5664 ( .A(n3955), .B(key[129]), .Z(n3937) );
  XNOR U5665 ( .A(\w3[0][25] ), .B(n3935), .Z(n3936) );
  XNOR U5666 ( .A(n3937), .B(n3936), .Z(\w1[1][1] ) );
  XOR U5667 ( .A(\w3[0][16] ), .B(\w3[0][21] ), .Z(n3969) );
  XOR U5668 ( .A(n3969), .B(key[148]), .Z(n3940) );
  XNOR U5669 ( .A(\w3[0][12] ), .B(n3938), .Z(n3939) );
  XNOR U5670 ( .A(n3940), .B(n3939), .Z(\w1[1][20] ) );
  XOR U5671 ( .A(\w3[0][14] ), .B(\w3[0][22] ), .Z(n3979) );
  XOR U5672 ( .A(n3979), .B(key[149]), .Z(n3943) );
  XNOR U5673 ( .A(\w3[0][13] ), .B(n3941), .Z(n3942) );
  XNOR U5674 ( .A(n3943), .B(n3942), .Z(\w1[1][21] ) );
  XOR U5675 ( .A(\w3[0][16] ), .B(\w3[0][23] ), .Z(n3980) );
  XOR U5676 ( .A(n3980), .B(key[150]), .Z(n3946) );
  XNOR U5677 ( .A(\w3[0][14] ), .B(n3944), .Z(n3945) );
  XNOR U5678 ( .A(n3946), .B(n3945), .Z(\w1[1][22] ) );
  XNOR U5679 ( .A(n3947), .B(key[151]), .Z(n3948) );
  XNOR U5680 ( .A(n3949), .B(n3948), .Z(n3950) );
  XNOR U5681 ( .A(\w3[0][16] ), .B(n3950), .Z(\w1[1][23] ) );
  XOR U5682 ( .A(\w3[0][17] ), .B(key[152]), .Z(n3953) );
  XNOR U5683 ( .A(\w3[0][25] ), .B(n3951), .Z(n3952) );
  XNOR U5684 ( .A(n3953), .B(n3952), .Z(n3954) );
  XOR U5685 ( .A(\w3[0][16] ), .B(n3954), .Z(\w1[1][24] ) );
  XOR U5686 ( .A(n3955), .B(key[153]), .Z(n3957) );
  XNOR U5687 ( .A(\w3[0][1] ), .B(\w3[0][26] ), .Z(n3956) );
  XNOR U5688 ( .A(n3957), .B(n3956), .Z(n3958) );
  XOR U5689 ( .A(\w3[0][18] ), .B(n3958), .Z(\w1[1][25] ) );
  XOR U5690 ( .A(n3975), .B(key[154]), .Z(n3960) );
  XNOR U5691 ( .A(\w3[0][2] ), .B(\w3[0][19] ), .Z(n3959) );
  XNOR U5692 ( .A(n3960), .B(n3959), .Z(n3961) );
  XOR U5693 ( .A(\w3[0][27] ), .B(n3961), .Z(\w1[1][26] ) );
  XNOR U5694 ( .A(\w3[0][24] ), .B(\w3[0][28] ), .Z(n3962) );
  XNOR U5695 ( .A(n3963), .B(n3962), .Z(n4005) );
  XOR U5696 ( .A(n4005), .B(key[155]), .Z(n3966) );
  XNOR U5697 ( .A(\w3[0][3] ), .B(n3964), .Z(n3965) );
  XNOR U5698 ( .A(n3966), .B(n3965), .Z(\w1[1][27] ) );
  XOR U5699 ( .A(\w3[0][20] ), .B(\w3[0][29] ), .Z(n3968) );
  XNOR U5700 ( .A(\w3[0][24] ), .B(\w3[0][12] ), .Z(n3967) );
  XNOR U5701 ( .A(n3968), .B(n3967), .Z(n4042) );
  XOR U5702 ( .A(n4042), .B(key[156]), .Z(n3971) );
  XNOR U5703 ( .A(\w3[0][4] ), .B(n3969), .Z(n3970) );
  XNOR U5704 ( .A(n3971), .B(n3970), .Z(\w1[1][28] ) );
  XOR U5705 ( .A(\w3[0][13] ), .B(\w3[0][21] ), .Z(n4083) );
  XOR U5706 ( .A(n4083), .B(key[157]), .Z(n3973) );
  XNOR U5707 ( .A(\w3[0][22] ), .B(\w3[0][30] ), .Z(n3972) );
  XNOR U5708 ( .A(n3973), .B(n3972), .Z(n3974) );
  XOR U5709 ( .A(\w3[0][5] ), .B(n3974), .Z(\w1[1][29] ) );
  XOR U5710 ( .A(n3975), .B(key[130]), .Z(n3978) );
  XNOR U5711 ( .A(\w3[0][26] ), .B(n3976), .Z(n3977) );
  XNOR U5712 ( .A(n3978), .B(n3977), .Z(\w1[1][2] ) );
  XNOR U5713 ( .A(\w3[0][24] ), .B(\w3[0][31] ), .Z(n4157) );
  XNOR U5714 ( .A(n3979), .B(n4157), .Z(n4118) );
  XOR U5715 ( .A(n4118), .B(key[158]), .Z(n3982) );
  XNOR U5716 ( .A(\w3[0][6] ), .B(n3980), .Z(n3981) );
  XNOR U5717 ( .A(n3982), .B(n3981), .Z(\w1[1][30] ) );
  XOR U5718 ( .A(\w3[0][15] ), .B(\w3[0][23] ), .Z(n4155) );
  XOR U5719 ( .A(n4155), .B(key[159]), .Z(n3984) );
  XNOR U5720 ( .A(n4196), .B(\w3[0][7] ), .Z(n3983) );
  XNOR U5721 ( .A(n3984), .B(n3983), .Z(\w1[1][31] ) );
  XOR U5722 ( .A(\w3[0][33] ), .B(\w3[0][57] ), .Z(n4039) );
  XOR U5723 ( .A(n4039), .B(key[160]), .Z(n3986) );
  XOR U5724 ( .A(\w3[0][48] ), .B(\w3[0][56] ), .Z(n4100) );
  XNOR U5725 ( .A(n4100), .B(\w3[0][40] ), .Z(n3985) );
  XNOR U5726 ( .A(n3986), .B(n3985), .Z(\w1[1][32] ) );
  XOR U5727 ( .A(\w3[0][34] ), .B(\w3[0][58] ), .Z(n4047) );
  XOR U5728 ( .A(n4047), .B(key[161]), .Z(n3988) );
  XOR U5729 ( .A(\w3[0][41] ), .B(\w3[0][49] ), .Z(n4071) );
  XNOR U5730 ( .A(\w3[0][57] ), .B(n4071), .Z(n3987) );
  XNOR U5731 ( .A(n3988), .B(n3987), .Z(\w1[1][33] ) );
  XOR U5732 ( .A(\w3[0][35] ), .B(\w3[0][59] ), .Z(n4018) );
  XOR U5733 ( .A(n4018), .B(key[162]), .Z(n3990) );
  XOR U5734 ( .A(\w3[0][42] ), .B(\w3[0][50] ), .Z(n4075) );
  XNOR U5735 ( .A(\w3[0][58] ), .B(n4075), .Z(n3989) );
  XNOR U5736 ( .A(n3990), .B(n3989), .Z(\w1[1][34] ) );
  XOR U5737 ( .A(\w3[0][36] ), .B(\w3[0][32] ), .Z(n4020) );
  XOR U5738 ( .A(n4020), .B(key[163]), .Z(n3993) );
  XOR U5739 ( .A(\w3[0][43] ), .B(\w3[0][51] ), .Z(n4046) );
  XNOR U5740 ( .A(\w3[0][56] ), .B(n4046), .Z(n3991) );
  XNOR U5741 ( .A(\w3[0][60] ), .B(n3991), .Z(n4080) );
  XNOR U5742 ( .A(\w3[0][59] ), .B(n4080), .Z(n3992) );
  XNOR U5743 ( .A(n3993), .B(n3992), .Z(\w1[1][35] ) );
  XOR U5744 ( .A(\w3[0][32] ), .B(\w3[0][37] ), .Z(n4025) );
  XOR U5745 ( .A(n4025), .B(key[164]), .Z(n3997) );
  XOR U5746 ( .A(\w3[0][52] ), .B(\w3[0][61] ), .Z(n3995) );
  XNOR U5747 ( .A(\w3[0][56] ), .B(\w3[0][44] ), .Z(n3994) );
  XNOR U5748 ( .A(n3995), .B(n3994), .Z(n4088) );
  XNOR U5749 ( .A(\w3[0][60] ), .B(n4088), .Z(n3996) );
  XNOR U5750 ( .A(n3997), .B(n3996), .Z(\w1[1][36] ) );
  XOR U5751 ( .A(\w3[0][38] ), .B(\w3[0][62] ), .Z(n4031) );
  XOR U5752 ( .A(n4031), .B(key[165]), .Z(n3999) );
  XOR U5753 ( .A(\w3[0][45] ), .B(\w3[0][53] ), .Z(n4091) );
  XNOR U5754 ( .A(\w3[0][61] ), .B(n4091), .Z(n3998) );
  XNOR U5755 ( .A(n3999), .B(n3998), .Z(\w1[1][37] ) );
  XOR U5756 ( .A(\w3[0][32] ), .B(\w3[0][39] ), .Z(n4032) );
  XOR U5757 ( .A(n4032), .B(key[166]), .Z(n4001) );
  XOR U5758 ( .A(\w3[0][46] ), .B(\w3[0][54] ), .Z(n4057) );
  XNOR U5759 ( .A(\w3[0][56] ), .B(\w3[0][63] ), .Z(n4003) );
  XNOR U5760 ( .A(n4057), .B(n4003), .Z(n4096) );
  XNOR U5761 ( .A(\w3[0][62] ), .B(n4096), .Z(n4000) );
  XNOR U5762 ( .A(n4001), .B(n4000), .Z(\w1[1][38] ) );
  XOR U5763 ( .A(\w3[0][47] ), .B(\w3[0][55] ), .Z(n4099) );
  XNOR U5764 ( .A(n4099), .B(key[167]), .Z(n4002) );
  XNOR U5765 ( .A(n4003), .B(n4002), .Z(n4004) );
  XNOR U5766 ( .A(\w3[0][32] ), .B(n4004), .Z(\w1[1][39] ) );
  XOR U5767 ( .A(n4005), .B(key[131]), .Z(n4008) );
  XNOR U5768 ( .A(n4006), .B(\w3[0][27] ), .Z(n4007) );
  XNOR U5769 ( .A(n4008), .B(n4007), .Z(\w1[1][3] ) );
  XOR U5770 ( .A(\w3[0][32] ), .B(key[168]), .Z(n4010) );
  XNOR U5771 ( .A(\w3[0][33] ), .B(\w3[0][41] ), .Z(n4009) );
  XNOR U5772 ( .A(n4010), .B(n4009), .Z(n4011) );
  XOR U5773 ( .A(n4100), .B(n4011), .Z(\w1[1][40] ) );
  XOR U5774 ( .A(\w3[0][42] ), .B(key[169]), .Z(n4013) );
  XNOR U5775 ( .A(\w3[0][49] ), .B(\w3[0][34] ), .Z(n4012) );
  XNOR U5776 ( .A(n4013), .B(n4012), .Z(n4014) );
  XOR U5777 ( .A(n4039), .B(n4014), .Z(\w1[1][41] ) );
  XOR U5778 ( .A(\w3[0][43] ), .B(key[170]), .Z(n4016) );
  XNOR U5779 ( .A(\w3[0][50] ), .B(\w3[0][35] ), .Z(n4015) );
  XNOR U5780 ( .A(n4016), .B(n4015), .Z(n4017) );
  XOR U5781 ( .A(n4047), .B(n4017), .Z(\w1[1][42] ) );
  XNOR U5782 ( .A(\w3[0][40] ), .B(n4018), .Z(n4019) );
  XNOR U5783 ( .A(\w3[0][44] ), .B(n4019), .Z(n4050) );
  XOR U5784 ( .A(n4050), .B(key[171]), .Z(n4022) );
  XNOR U5785 ( .A(\w3[0][51] ), .B(n4020), .Z(n4021) );
  XNOR U5786 ( .A(n4022), .B(n4021), .Z(\w1[1][43] ) );
  XOR U5787 ( .A(\w3[0][36] ), .B(\w3[0][45] ), .Z(n4024) );
  XNOR U5788 ( .A(\w3[0][40] ), .B(\w3[0][60] ), .Z(n4023) );
  XNOR U5789 ( .A(n4024), .B(n4023), .Z(n4053) );
  XOR U5790 ( .A(n4053), .B(key[172]), .Z(n4027) );
  XNOR U5791 ( .A(\w3[0][52] ), .B(n4025), .Z(n4026) );
  XNOR U5792 ( .A(n4027), .B(n4026), .Z(\w1[1][44] ) );
  XOR U5793 ( .A(\w3[0][61] ), .B(\w3[0][37] ), .Z(n4056) );
  XOR U5794 ( .A(n4056), .B(key[173]), .Z(n4029) );
  XNOR U5795 ( .A(\w3[0][38] ), .B(\w3[0][46] ), .Z(n4028) );
  XNOR U5796 ( .A(n4029), .B(n4028), .Z(n4030) );
  XOR U5797 ( .A(\w3[0][53] ), .B(n4030), .Z(\w1[1][45] ) );
  XNOR U5798 ( .A(\w3[0][40] ), .B(\w3[0][47] ), .Z(n4065) );
  XNOR U5799 ( .A(n4031), .B(n4065), .Z(n4060) );
  XOR U5800 ( .A(n4060), .B(key[174]), .Z(n4034) );
  XNOR U5801 ( .A(\w3[0][54] ), .B(n4032), .Z(n4033) );
  XNOR U5802 ( .A(n4034), .B(n4033), .Z(\w1[1][46] ) );
  XOR U5803 ( .A(\w3[0][63] ), .B(\w3[0][39] ), .Z(n4063) );
  XOR U5804 ( .A(n4063), .B(key[175]), .Z(n4036) );
  XOR U5805 ( .A(\w3[0][40] ), .B(\w3[0][32] ), .Z(n4067) );
  XNOR U5806 ( .A(\w3[0][55] ), .B(n4067), .Z(n4035) );
  XNOR U5807 ( .A(n4036), .B(n4035), .Z(\w1[1][47] ) );
  XOR U5808 ( .A(n4067), .B(key[176]), .Z(n4038) );
  XNOR U5809 ( .A(\w3[0][56] ), .B(n4071), .Z(n4037) );
  XNOR U5810 ( .A(n4038), .B(n4037), .Z(\w1[1][48] ) );
  XOR U5811 ( .A(n4075), .B(key[177]), .Z(n4041) );
  XNOR U5812 ( .A(n4039), .B(\w3[0][41] ), .Z(n4040) );
  XNOR U5813 ( .A(n4041), .B(n4040), .Z(\w1[1][49] ) );
  XOR U5814 ( .A(n4042), .B(key[132]), .Z(n4045) );
  XNOR U5815 ( .A(n4043), .B(\w3[0][28] ), .Z(n4044) );
  XNOR U5816 ( .A(n4045), .B(n4044), .Z(\w1[1][4] ) );
  XOR U5817 ( .A(n4046), .B(key[178]), .Z(n4049) );
  XNOR U5818 ( .A(n4047), .B(\w3[0][42] ), .Z(n4048) );
  XNOR U5819 ( .A(n4049), .B(n4048), .Z(\w1[1][50] ) );
  XOR U5820 ( .A(\w3[0][48] ), .B(\w3[0][52] ), .Z(n4079) );
  XOR U5821 ( .A(n4079), .B(key[179]), .Z(n4052) );
  XNOR U5822 ( .A(\w3[0][43] ), .B(n4050), .Z(n4051) );
  XNOR U5823 ( .A(n4052), .B(n4051), .Z(\w1[1][51] ) );
  XOR U5824 ( .A(\w3[0][48] ), .B(\w3[0][53] ), .Z(n4087) );
  XOR U5825 ( .A(n4087), .B(key[180]), .Z(n4055) );
  XNOR U5826 ( .A(\w3[0][44] ), .B(n4053), .Z(n4054) );
  XNOR U5827 ( .A(n4055), .B(n4054), .Z(\w1[1][52] ) );
  XOR U5828 ( .A(n4056), .B(key[181]), .Z(n4059) );
  XNOR U5829 ( .A(\w3[0][45] ), .B(n4057), .Z(n4058) );
  XNOR U5830 ( .A(n4059), .B(n4058), .Z(\w1[1][53] ) );
  XOR U5831 ( .A(\w3[0][48] ), .B(\w3[0][55] ), .Z(n4095) );
  XOR U5832 ( .A(n4095), .B(key[182]), .Z(n4062) );
  XNOR U5833 ( .A(\w3[0][46] ), .B(n4060), .Z(n4061) );
  XNOR U5834 ( .A(n4062), .B(n4061), .Z(\w1[1][54] ) );
  XNOR U5835 ( .A(n4063), .B(key[183]), .Z(n4064) );
  XNOR U5836 ( .A(n4065), .B(n4064), .Z(n4066) );
  XNOR U5837 ( .A(\w3[0][48] ), .B(n4066), .Z(\w1[1][55] ) );
  XOR U5838 ( .A(n4067), .B(key[184]), .Z(n4069) );
  XNOR U5839 ( .A(\w3[0][48] ), .B(\w3[0][49] ), .Z(n4068) );
  XNOR U5840 ( .A(n4069), .B(n4068), .Z(n4070) );
  XOR U5841 ( .A(\w3[0][57] ), .B(n4070), .Z(\w1[1][56] ) );
  XOR U5842 ( .A(\w3[0][50] ), .B(key[185]), .Z(n4073) );
  XNOR U5843 ( .A(n4071), .B(\w3[0][58] ), .Z(n4072) );
  XNOR U5844 ( .A(n4073), .B(n4072), .Z(n4074) );
  XOR U5845 ( .A(\w3[0][33] ), .B(n4074), .Z(\w1[1][57] ) );
  XOR U5846 ( .A(\w3[0][51] ), .B(key[186]), .Z(n4077) );
  XNOR U5847 ( .A(n4075), .B(\w3[0][59] ), .Z(n4076) );
  XNOR U5848 ( .A(n4077), .B(n4076), .Z(n4078) );
  XOR U5849 ( .A(\w3[0][34] ), .B(n4078), .Z(\w1[1][58] ) );
  XOR U5850 ( .A(n4079), .B(key[187]), .Z(n4082) );
  XNOR U5851 ( .A(\w3[0][35] ), .B(n4080), .Z(n4081) );
  XNOR U5852 ( .A(n4082), .B(n4081), .Z(\w1[1][59] ) );
  XOR U5853 ( .A(n4083), .B(key[133]), .Z(n4086) );
  XNOR U5854 ( .A(\w3[0][29] ), .B(n4084), .Z(n4085) );
  XNOR U5855 ( .A(n4086), .B(n4085), .Z(\w1[1][5] ) );
  XOR U5856 ( .A(n4087), .B(key[188]), .Z(n4090) );
  XNOR U5857 ( .A(\w3[0][36] ), .B(n4088), .Z(n4089) );
  XNOR U5858 ( .A(n4090), .B(n4089), .Z(\w1[1][60] ) );
  XOR U5859 ( .A(\w3[0][54] ), .B(key[189]), .Z(n4093) );
  XNOR U5860 ( .A(n4091), .B(\w3[0][62] ), .Z(n4092) );
  XNOR U5861 ( .A(n4093), .B(n4092), .Z(n4094) );
  XOR U5862 ( .A(\w3[0][37] ), .B(n4094), .Z(\w1[1][61] ) );
  XOR U5863 ( .A(n4095), .B(key[190]), .Z(n4098) );
  XNOR U5864 ( .A(\w3[0][38] ), .B(n4096), .Z(n4097) );
  XNOR U5865 ( .A(n4098), .B(n4097), .Z(\w1[1][62] ) );
  XOR U5866 ( .A(n4099), .B(key[191]), .Z(n4102) );
  XNOR U5867 ( .A(n4100), .B(\w3[0][39] ), .Z(n4101) );
  XNOR U5868 ( .A(n4102), .B(n4101), .Z(\w1[1][63] ) );
  XOR U5869 ( .A(\w3[0][65] ), .B(\w3[0][89] ), .Z(n4161) );
  XOR U5870 ( .A(n4161), .B(key[192]), .Z(n4104) );
  XOR U5871 ( .A(\w3[0][80] ), .B(\w3[0][88] ), .Z(n4218) );
  XNOR U5872 ( .A(n4218), .B(\w3[0][72] ), .Z(n4103) );
  XNOR U5873 ( .A(n4104), .B(n4103), .Z(\w1[1][64] ) );
  XOR U5874 ( .A(\w3[0][66] ), .B(\w3[0][90] ), .Z(n4165) );
  XOR U5875 ( .A(n4165), .B(key[193]), .Z(n4106) );
  XOR U5876 ( .A(\w3[0][73] ), .B(\w3[0][81] ), .Z(n4189) );
  XNOR U5877 ( .A(\w3[0][89] ), .B(n4189), .Z(n4105) );
  XNOR U5878 ( .A(n4106), .B(n4105), .Z(\w1[1][65] ) );
  XOR U5879 ( .A(\w3[0][67] ), .B(\w3[0][91] ), .Z(n4136) );
  XOR U5880 ( .A(n4136), .B(key[194]), .Z(n4108) );
  XOR U5881 ( .A(\w3[0][74] ), .B(\w3[0][82] ), .Z(n4197) );
  XNOR U5882 ( .A(\w3[0][90] ), .B(n4197), .Z(n4107) );
  XNOR U5883 ( .A(n4108), .B(n4107), .Z(\w1[1][66] ) );
  XOR U5884 ( .A(\w3[0][68] ), .B(\w3[0][64] ), .Z(n4138) );
  XOR U5885 ( .A(n4138), .B(key[195]), .Z(n4111) );
  XOR U5886 ( .A(\w3[0][75] ), .B(\w3[0][83] ), .Z(n4164) );
  XNOR U5887 ( .A(\w3[0][88] ), .B(n4164), .Z(n4109) );
  XNOR U5888 ( .A(\w3[0][92] ), .B(n4109), .Z(n4202) );
  XNOR U5889 ( .A(\w3[0][91] ), .B(n4202), .Z(n4110) );
  XNOR U5890 ( .A(n4111), .B(n4110), .Z(\w1[1][67] ) );
  XOR U5891 ( .A(\w3[0][64] ), .B(\w3[0][69] ), .Z(n4143) );
  XOR U5892 ( .A(n4143), .B(key[196]), .Z(n4115) );
  XOR U5893 ( .A(\w3[0][84] ), .B(\w3[0][93] ), .Z(n4113) );
  XNOR U5894 ( .A(\w3[0][88] ), .B(\w3[0][76] ), .Z(n4112) );
  XNOR U5895 ( .A(n4113), .B(n4112), .Z(n4206) );
  XNOR U5896 ( .A(\w3[0][92] ), .B(n4206), .Z(n4114) );
  XNOR U5897 ( .A(n4115), .B(n4114), .Z(\w1[1][68] ) );
  XOR U5898 ( .A(\w3[0][70] ), .B(\w3[0][94] ), .Z(n4149) );
  XOR U5899 ( .A(n4149), .B(key[197]), .Z(n4117) );
  XOR U5900 ( .A(\w3[0][77] ), .B(\w3[0][85] ), .Z(n4209) );
  XNOR U5901 ( .A(\w3[0][93] ), .B(n4209), .Z(n4116) );
  XNOR U5902 ( .A(n4117), .B(n4116), .Z(\w1[1][69] ) );
  XOR U5903 ( .A(n4118), .B(key[134]), .Z(n4121) );
  XNOR U5904 ( .A(n4119), .B(\w3[0][30] ), .Z(n4120) );
  XNOR U5905 ( .A(n4121), .B(n4120), .Z(\w1[1][6] ) );
  XOR U5906 ( .A(\w3[0][64] ), .B(\w3[0][71] ), .Z(n4150) );
  XOR U5907 ( .A(n4150), .B(key[198]), .Z(n4123) );
  XOR U5908 ( .A(\w3[0][78] ), .B(\w3[0][86] ), .Z(n4175) );
  XNOR U5909 ( .A(\w3[0][88] ), .B(\w3[0][95] ), .Z(n4125) );
  XNOR U5910 ( .A(n4175), .B(n4125), .Z(n4214) );
  XNOR U5911 ( .A(\w3[0][94] ), .B(n4214), .Z(n4122) );
  XNOR U5912 ( .A(n4123), .B(n4122), .Z(\w1[1][70] ) );
  XOR U5913 ( .A(\w3[0][79] ), .B(\w3[0][87] ), .Z(n4217) );
  XNOR U5914 ( .A(n4217), .B(key[199]), .Z(n4124) );
  XNOR U5915 ( .A(n4125), .B(n4124), .Z(n4126) );
  XNOR U5916 ( .A(\w3[0][64] ), .B(n4126), .Z(\w1[1][71] ) );
  XOR U5917 ( .A(\w3[0][64] ), .B(key[200]), .Z(n4128) );
  XNOR U5918 ( .A(\w3[0][65] ), .B(\w3[0][73] ), .Z(n4127) );
  XNOR U5919 ( .A(n4128), .B(n4127), .Z(n4129) );
  XOR U5920 ( .A(n4218), .B(n4129), .Z(\w1[1][72] ) );
  XOR U5921 ( .A(\w3[0][74] ), .B(key[201]), .Z(n4131) );
  XNOR U5922 ( .A(\w3[0][81] ), .B(\w3[0][66] ), .Z(n4130) );
  XNOR U5923 ( .A(n4131), .B(n4130), .Z(n4132) );
  XOR U5924 ( .A(n4161), .B(n4132), .Z(\w1[1][73] ) );
  XOR U5925 ( .A(\w3[0][75] ), .B(key[202]), .Z(n4134) );
  XNOR U5926 ( .A(\w3[0][82] ), .B(\w3[0][67] ), .Z(n4133) );
  XNOR U5927 ( .A(n4134), .B(n4133), .Z(n4135) );
  XOR U5928 ( .A(n4165), .B(n4135), .Z(\w1[1][74] ) );
  XNOR U5929 ( .A(\w3[0][72] ), .B(n4136), .Z(n4137) );
  XNOR U5930 ( .A(\w3[0][76] ), .B(n4137), .Z(n4168) );
  XOR U5931 ( .A(n4168), .B(key[203]), .Z(n4140) );
  XNOR U5932 ( .A(\w3[0][83] ), .B(n4138), .Z(n4139) );
  XNOR U5933 ( .A(n4140), .B(n4139), .Z(\w1[1][75] ) );
  XOR U5934 ( .A(\w3[0][68] ), .B(\w3[0][77] ), .Z(n4142) );
  XNOR U5935 ( .A(\w3[0][72] ), .B(\w3[0][92] ), .Z(n4141) );
  XNOR U5936 ( .A(n4142), .B(n4141), .Z(n4171) );
  XOR U5937 ( .A(n4171), .B(key[204]), .Z(n4145) );
  XNOR U5938 ( .A(\w3[0][84] ), .B(n4143), .Z(n4144) );
  XNOR U5939 ( .A(n4145), .B(n4144), .Z(\w1[1][76] ) );
  XOR U5940 ( .A(\w3[0][93] ), .B(\w3[0][69] ), .Z(n4174) );
  XOR U5941 ( .A(n4174), .B(key[205]), .Z(n4147) );
  XNOR U5942 ( .A(\w3[0][70] ), .B(\w3[0][78] ), .Z(n4146) );
  XNOR U5943 ( .A(n4147), .B(n4146), .Z(n4148) );
  XOR U5944 ( .A(\w3[0][85] ), .B(n4148), .Z(\w1[1][77] ) );
  XNOR U5945 ( .A(\w3[0][72] ), .B(\w3[0][79] ), .Z(n4183) );
  XNOR U5946 ( .A(n4149), .B(n4183), .Z(n4178) );
  XOR U5947 ( .A(n4178), .B(key[206]), .Z(n4152) );
  XNOR U5948 ( .A(\w3[0][86] ), .B(n4150), .Z(n4151) );
  XNOR U5949 ( .A(n4152), .B(n4151), .Z(\w1[1][78] ) );
  XOR U5950 ( .A(\w3[0][95] ), .B(\w3[0][71] ), .Z(n4181) );
  XOR U5951 ( .A(n4181), .B(key[207]), .Z(n4154) );
  XOR U5952 ( .A(\w3[0][72] ), .B(\w3[0][64] ), .Z(n4185) );
  XNOR U5953 ( .A(\w3[0][87] ), .B(n4185), .Z(n4153) );
  XNOR U5954 ( .A(n4154), .B(n4153), .Z(\w1[1][79] ) );
  XNOR U5955 ( .A(n4155), .B(key[135]), .Z(n4156) );
  XNOR U5956 ( .A(n4157), .B(n4156), .Z(n4158) );
  XNOR U5957 ( .A(\w3[0][0] ), .B(n4158), .Z(\w1[1][7] ) );
  XOR U5958 ( .A(n4185), .B(key[208]), .Z(n4160) );
  XNOR U5959 ( .A(\w3[0][88] ), .B(n4189), .Z(n4159) );
  XNOR U5960 ( .A(n4160), .B(n4159), .Z(\w1[1][80] ) );
  XOR U5961 ( .A(n4197), .B(key[209]), .Z(n4163) );
  XNOR U5962 ( .A(n4161), .B(\w3[0][73] ), .Z(n4162) );
  XNOR U5963 ( .A(n4163), .B(n4162), .Z(\w1[1][81] ) );
  XOR U5964 ( .A(n4164), .B(key[210]), .Z(n4167) );
  XNOR U5965 ( .A(n4165), .B(\w3[0][74] ), .Z(n4166) );
  XNOR U5966 ( .A(n4167), .B(n4166), .Z(\w1[1][82] ) );
  XOR U5967 ( .A(\w3[0][80] ), .B(\w3[0][84] ), .Z(n4201) );
  XOR U5968 ( .A(n4201), .B(key[211]), .Z(n4170) );
  XNOR U5969 ( .A(\w3[0][75] ), .B(n4168), .Z(n4169) );
  XNOR U5970 ( .A(n4170), .B(n4169), .Z(\w1[1][83] ) );
  XOR U5971 ( .A(\w3[0][80] ), .B(\w3[0][85] ), .Z(n4205) );
  XOR U5972 ( .A(n4205), .B(key[212]), .Z(n4173) );
  XNOR U5973 ( .A(\w3[0][76] ), .B(n4171), .Z(n4172) );
  XNOR U5974 ( .A(n4173), .B(n4172), .Z(\w1[1][84] ) );
  XOR U5975 ( .A(n4174), .B(key[213]), .Z(n4177) );
  XNOR U5976 ( .A(\w3[0][77] ), .B(n4175), .Z(n4176) );
  XNOR U5977 ( .A(n4177), .B(n4176), .Z(\w1[1][85] ) );
  XOR U5978 ( .A(\w3[0][80] ), .B(\w3[0][87] ), .Z(n4213) );
  XOR U5979 ( .A(n4213), .B(key[214]), .Z(n4180) );
  XNOR U5980 ( .A(\w3[0][78] ), .B(n4178), .Z(n4179) );
  XNOR U5981 ( .A(n4180), .B(n4179), .Z(\w1[1][86] ) );
  XNOR U5982 ( .A(n4181), .B(key[215]), .Z(n4182) );
  XNOR U5983 ( .A(n4183), .B(n4182), .Z(n4184) );
  XNOR U5984 ( .A(\w3[0][80] ), .B(n4184), .Z(\w1[1][87] ) );
  XOR U5985 ( .A(n4185), .B(key[216]), .Z(n4187) );
  XNOR U5986 ( .A(\w3[0][80] ), .B(\w3[0][81] ), .Z(n4186) );
  XNOR U5987 ( .A(n4187), .B(n4186), .Z(n4188) );
  XOR U5988 ( .A(\w3[0][89] ), .B(n4188), .Z(\w1[1][88] ) );
  XOR U5989 ( .A(\w3[0][82] ), .B(key[217]), .Z(n4191) );
  XNOR U5990 ( .A(n4189), .B(\w3[0][90] ), .Z(n4190) );
  XNOR U5991 ( .A(n4191), .B(n4190), .Z(n4192) );
  XOR U5992 ( .A(\w3[0][65] ), .B(n4192), .Z(\w1[1][89] ) );
  XOR U5993 ( .A(\w3[0][9] ), .B(key[136]), .Z(n4194) );
  XNOR U5994 ( .A(\w3[0][1] ), .B(\w3[0][0] ), .Z(n4193) );
  XNOR U5995 ( .A(n4194), .B(n4193), .Z(n4195) );
  XOR U5996 ( .A(n4196), .B(n4195), .Z(\w1[1][8] ) );
  XOR U5997 ( .A(\w3[0][83] ), .B(key[218]), .Z(n4199) );
  XNOR U5998 ( .A(n4197), .B(\w3[0][91] ), .Z(n4198) );
  XNOR U5999 ( .A(n4199), .B(n4198), .Z(n4200) );
  XOR U6000 ( .A(\w3[0][66] ), .B(n4200), .Z(\w1[1][90] ) );
  XOR U6001 ( .A(n4201), .B(key[219]), .Z(n4204) );
  XNOR U6002 ( .A(\w3[0][67] ), .B(n4202), .Z(n4203) );
  XNOR U6003 ( .A(n4204), .B(n4203), .Z(\w1[1][91] ) );
  XOR U6004 ( .A(n4205), .B(key[220]), .Z(n4208) );
  XNOR U6005 ( .A(\w3[0][68] ), .B(n4206), .Z(n4207) );
  XNOR U6006 ( .A(n4208), .B(n4207), .Z(\w1[1][92] ) );
  XOR U6007 ( .A(\w3[0][86] ), .B(key[221]), .Z(n4211) );
  XNOR U6008 ( .A(n4209), .B(\w3[0][94] ), .Z(n4210) );
  XNOR U6009 ( .A(n4211), .B(n4210), .Z(n4212) );
  XOR U6010 ( .A(\w3[0][69] ), .B(n4212), .Z(\w1[1][93] ) );
  XOR U6011 ( .A(n4213), .B(key[222]), .Z(n4216) );
  XNOR U6012 ( .A(\w3[0][70] ), .B(n4214), .Z(n4215) );
  XNOR U6013 ( .A(n4216), .B(n4215), .Z(\w1[1][94] ) );
  XOR U6014 ( .A(n4217), .B(key[223]), .Z(n4220) );
  XNOR U6015 ( .A(n4218), .B(\w3[0][71] ), .Z(n4219) );
  XNOR U6016 ( .A(n4220), .B(n4219), .Z(\w1[1][95] ) );
  XOR U6017 ( .A(\w3[0][104] ), .B(key[224]), .Z(n4224) );
  XOR U6018 ( .A(n4222), .B(n4221), .Z(n4223) );
  XNOR U6019 ( .A(n4224), .B(n4223), .Z(\w1[1][96] ) );
  XOR U6020 ( .A(n4225), .B(key[225]), .Z(n4228) );
  XNOR U6021 ( .A(\w3[0][121] ), .B(n4226), .Z(n4227) );
  XNOR U6022 ( .A(n4228), .B(n4227), .Z(\w1[1][97] ) );
  XOR U6023 ( .A(n4229), .B(key[226]), .Z(n4232) );
  XNOR U6024 ( .A(\w3[0][122] ), .B(n4230), .Z(n4231) );
  XNOR U6025 ( .A(n4232), .B(n4231), .Z(\w1[1][98] ) );
  XOR U6026 ( .A(n4233), .B(key[227]), .Z(n4236) );
  XNOR U6027 ( .A(n4234), .B(\w3[0][123] ), .Z(n4235) );
  XNOR U6028 ( .A(n4236), .B(n4235), .Z(\w1[1][99] ) );
  XOR U6029 ( .A(\w3[0][10] ), .B(key[137]), .Z(n4238) );
  XNOR U6030 ( .A(\w3[0][2] ), .B(\w3[0][17] ), .Z(n4237) );
  XNOR U6031 ( .A(n4238), .B(n4237), .Z(n4239) );
  XOR U6032 ( .A(n4240), .B(n4239), .Z(\w1[1][9] ) );
  XOR U6033 ( .A(\w3[1][8] ), .B(key[256]), .Z(n4242) );
  XOR U6034 ( .A(\w3[1][1] ), .B(\w3[1][25] ), .Z(n4664) );
  XOR U6035 ( .A(\w3[1][16] ), .B(\w3[1][24] ), .Z(n4620) );
  XNOR U6036 ( .A(n4664), .B(n4620), .Z(n4241) );
  XNOR U6037 ( .A(n4242), .B(n4241), .Z(\w1[2][0] ) );
  XOR U6038 ( .A(\w3[1][96] ), .B(\w3[1][101] ), .Z(n4267) );
  XOR U6039 ( .A(n4267), .B(key[356]), .Z(n4246) );
  XOR U6040 ( .A(\w3[1][116] ), .B(\w3[1][125] ), .Z(n4244) );
  XNOR U6041 ( .A(\w3[1][120] ), .B(\w3[1][108] ), .Z(n4243) );
  XNOR U6042 ( .A(n4244), .B(n4243), .Z(n4325) );
  XNOR U6043 ( .A(\w3[1][124] ), .B(n4325), .Z(n4245) );
  XNOR U6044 ( .A(n4246), .B(n4245), .Z(\w1[2][100] ) );
  XOR U6045 ( .A(\w3[1][102] ), .B(\w3[1][126] ), .Z(n4276) );
  XOR U6046 ( .A(n4276), .B(key[357]), .Z(n4248) );
  XOR U6047 ( .A(\w3[1][109] ), .B(\w3[1][117] ), .Z(n4328) );
  XNOR U6048 ( .A(\w3[1][125] ), .B(n4328), .Z(n4247) );
  XNOR U6049 ( .A(n4248), .B(n4247), .Z(\w1[2][101] ) );
  XOR U6050 ( .A(\w3[1][96] ), .B(\w3[1][103] ), .Z(n4277) );
  XOR U6051 ( .A(n4277), .B(key[358]), .Z(n4250) );
  XOR U6052 ( .A(\w3[1][110] ), .B(\w3[1][118] ), .Z(n4295) );
  XNOR U6053 ( .A(\w3[1][120] ), .B(\w3[1][127] ), .Z(n4252) );
  XNOR U6054 ( .A(n4295), .B(n4252), .Z(n4333) );
  XNOR U6055 ( .A(\w3[1][126] ), .B(n4333), .Z(n4249) );
  XNOR U6056 ( .A(n4250), .B(n4249), .Z(\w1[2][102] ) );
  XOR U6057 ( .A(\w3[1][111] ), .B(\w3[1][119] ), .Z(n4336) );
  XNOR U6058 ( .A(n4336), .B(key[359]), .Z(n4251) );
  XNOR U6059 ( .A(n4252), .B(n4251), .Z(n4253) );
  XNOR U6060 ( .A(\w3[1][96] ), .B(n4253), .Z(\w1[2][103] ) );
  XOR U6061 ( .A(\w3[1][105] ), .B(\w3[1][97] ), .Z(n4315) );
  XOR U6062 ( .A(n4315), .B(key[360]), .Z(n4255) );
  XOR U6063 ( .A(\w3[1][120] ), .B(\w3[1][112] ), .Z(n4646) );
  XNOR U6064 ( .A(\w3[1][96] ), .B(n4646), .Z(n4254) );
  XNOR U6065 ( .A(n4255), .B(n4254), .Z(\w1[2][104] ) );
  XOR U6066 ( .A(\w3[1][106] ), .B(\w3[1][113] ), .Z(n4257) );
  XOR U6067 ( .A(\w3[1][97] ), .B(\w3[1][121] ), .Z(n4645) );
  XNOR U6068 ( .A(n4645), .B(key[361]), .Z(n4256) );
  XNOR U6069 ( .A(n4257), .B(n4256), .Z(n4258) );
  XOR U6070 ( .A(\w3[1][98] ), .B(n4258), .Z(\w1[2][105] ) );
  XOR U6071 ( .A(\w3[1][107] ), .B(\w3[1][99] ), .Z(n4260) );
  XOR U6072 ( .A(\w3[1][98] ), .B(\w3[1][122] ), .Z(n4650) );
  XNOR U6073 ( .A(n4650), .B(key[362]), .Z(n4259) );
  XNOR U6074 ( .A(n4260), .B(n4259), .Z(n4261) );
  XOR U6075 ( .A(\w3[1][114] ), .B(n4261), .Z(\w1[2][106] ) );
  XOR U6076 ( .A(\w3[1][99] ), .B(\w3[1][123] ), .Z(n4654) );
  XNOR U6077 ( .A(\w3[1][108] ), .B(n4654), .Z(n4262) );
  XNOR U6078 ( .A(\w3[1][104] ), .B(n4262), .Z(n4288) );
  XOR U6079 ( .A(n4288), .B(key[363]), .Z(n4264) );
  XOR U6080 ( .A(\w3[1][96] ), .B(\w3[1][100] ), .Z(n4658) );
  XNOR U6081 ( .A(\w3[1][115] ), .B(n4658), .Z(n4263) );
  XNOR U6082 ( .A(n4264), .B(n4263), .Z(\w1[2][107] ) );
  XOR U6083 ( .A(\w3[1][100] ), .B(\w3[1][104] ), .Z(n4266) );
  XNOR U6084 ( .A(\w3[1][124] ), .B(\w3[1][109] ), .Z(n4265) );
  XNOR U6085 ( .A(n4266), .B(n4265), .Z(n4291) );
  XOR U6086 ( .A(n4291), .B(key[364]), .Z(n4269) );
  XNOR U6087 ( .A(\w3[1][116] ), .B(n4267), .Z(n4268) );
  XNOR U6088 ( .A(n4269), .B(n4268), .Z(\w1[2][108] ) );
  XOR U6089 ( .A(\w3[1][125] ), .B(\w3[1][101] ), .Z(n4294) );
  XOR U6090 ( .A(n4294), .B(key[365]), .Z(n4271) );
  XNOR U6091 ( .A(\w3[1][102] ), .B(\w3[1][110] ), .Z(n4270) );
  XNOR U6092 ( .A(n4271), .B(n4270), .Z(n4272) );
  XOR U6093 ( .A(\w3[1][117] ), .B(n4272), .Z(\w1[2][109] ) );
  XOR U6094 ( .A(\w3[1][11] ), .B(\w3[1][3] ), .Z(n4274) );
  XOR U6095 ( .A(\w3[1][2] ), .B(\w3[1][26] ), .Z(n4359) );
  XNOR U6096 ( .A(n4359), .B(key[266]), .Z(n4273) );
  XNOR U6097 ( .A(n4274), .B(n4273), .Z(n4275) );
  XOR U6098 ( .A(\w3[1][18] ), .B(n4275), .Z(\w1[2][10] ) );
  XNOR U6099 ( .A(\w3[1][111] ), .B(\w3[1][104] ), .Z(n4303) );
  XNOR U6100 ( .A(n4276), .B(n4303), .Z(n4298) );
  XOR U6101 ( .A(n4298), .B(key[366]), .Z(n4279) );
  XNOR U6102 ( .A(\w3[1][118] ), .B(n4277), .Z(n4278) );
  XNOR U6103 ( .A(n4279), .B(n4278), .Z(\w1[2][110] ) );
  XOR U6104 ( .A(\w3[1][127] ), .B(\w3[1][103] ), .Z(n4301) );
  XOR U6105 ( .A(n4301), .B(key[367]), .Z(n4281) );
  XOR U6106 ( .A(\w3[1][96] ), .B(\w3[1][104] ), .Z(n4308) );
  XNOR U6107 ( .A(\w3[1][119] ), .B(n4308), .Z(n4280) );
  XNOR U6108 ( .A(n4281), .B(n4280), .Z(\w1[2][111] ) );
  XOR U6109 ( .A(\w3[1][105] ), .B(\w3[1][113] ), .Z(n4649) );
  XOR U6110 ( .A(n4649), .B(key[368]), .Z(n4283) );
  XNOR U6111 ( .A(\w3[1][120] ), .B(n4308), .Z(n4282) );
  XNOR U6112 ( .A(n4283), .B(n4282), .Z(\w1[2][112] ) );
  XOR U6113 ( .A(\w3[1][106] ), .B(\w3[1][114] ), .Z(n4653) );
  XOR U6114 ( .A(n4653), .B(key[369]), .Z(n4285) );
  XNOR U6115 ( .A(n4315), .B(\w3[1][121] ), .Z(n4284) );
  XNOR U6116 ( .A(n4285), .B(n4284), .Z(\w1[2][113] ) );
  XOR U6117 ( .A(\w3[1][107] ), .B(\w3[1][115] ), .Z(n4320) );
  XOR U6118 ( .A(n4320), .B(key[370]), .Z(n4287) );
  XNOR U6119 ( .A(\w3[1][106] ), .B(n4650), .Z(n4286) );
  XNOR U6120 ( .A(n4287), .B(n4286), .Z(\w1[2][114] ) );
  XOR U6121 ( .A(\w3[1][116] ), .B(\w3[1][112] ), .Z(n4321) );
  XOR U6122 ( .A(n4321), .B(key[371]), .Z(n4290) );
  XNOR U6123 ( .A(\w3[1][107] ), .B(n4288), .Z(n4289) );
  XNOR U6124 ( .A(n4290), .B(n4289), .Z(\w1[2][115] ) );
  XOR U6125 ( .A(\w3[1][117] ), .B(\w3[1][112] ), .Z(n4324) );
  XOR U6126 ( .A(n4324), .B(key[372]), .Z(n4293) );
  XNOR U6127 ( .A(\w3[1][108] ), .B(n4291), .Z(n4292) );
  XNOR U6128 ( .A(n4293), .B(n4292), .Z(\w1[2][116] ) );
  XOR U6129 ( .A(n4294), .B(key[373]), .Z(n4297) );
  XNOR U6130 ( .A(\w3[1][109] ), .B(n4295), .Z(n4296) );
  XNOR U6131 ( .A(n4297), .B(n4296), .Z(\w1[2][117] ) );
  XOR U6132 ( .A(\w3[1][119] ), .B(\w3[1][112] ), .Z(n4332) );
  XOR U6133 ( .A(n4332), .B(key[374]), .Z(n4300) );
  XNOR U6134 ( .A(\w3[1][110] ), .B(n4298), .Z(n4299) );
  XNOR U6135 ( .A(n4300), .B(n4299), .Z(\w1[2][118] ) );
  XNOR U6136 ( .A(n4301), .B(key[375]), .Z(n4302) );
  XNOR U6137 ( .A(n4303), .B(n4302), .Z(n4304) );
  XNOR U6138 ( .A(\w3[1][112] ), .B(n4304), .Z(\w1[2][119] ) );
  XOR U6139 ( .A(\w3[1][3] ), .B(\w3[1][27] ), .Z(n4400) );
  XNOR U6140 ( .A(\w3[1][8] ), .B(\w3[1][12] ), .Z(n4305) );
  XNOR U6141 ( .A(n4400), .B(n4305), .Z(n4356) );
  XOR U6142 ( .A(n4356), .B(key[267]), .Z(n4307) );
  XOR U6143 ( .A(\w3[1][0] ), .B(\w3[1][4] ), .Z(n4430) );
  XNOR U6144 ( .A(\w3[1][19] ), .B(n4430), .Z(n4306) );
  XNOR U6145 ( .A(n4307), .B(n4306), .Z(\w1[2][11] ) );
  XOR U6146 ( .A(n4308), .B(key[376]), .Z(n4310) );
  XNOR U6147 ( .A(\w3[1][121] ), .B(\w3[1][113] ), .Z(n4309) );
  XNOR U6148 ( .A(n4310), .B(n4309), .Z(n4311) );
  XOR U6149 ( .A(\w3[1][112] ), .B(n4311), .Z(\w1[2][120] ) );
  XOR U6150 ( .A(\w3[1][122] ), .B(key[377]), .Z(n4313) );
  XNOR U6151 ( .A(\w3[1][113] ), .B(\w3[1][114] ), .Z(n4312) );
  XNOR U6152 ( .A(n4313), .B(n4312), .Z(n4314) );
  XOR U6153 ( .A(n4315), .B(n4314), .Z(\w1[2][121] ) );
  XOR U6154 ( .A(n4653), .B(key[378]), .Z(n4317) );
  XNOR U6155 ( .A(\w3[1][115] ), .B(\w3[1][123] ), .Z(n4316) );
  XNOR U6156 ( .A(n4317), .B(n4316), .Z(n4318) );
  XOR U6157 ( .A(\w3[1][98] ), .B(n4318), .Z(\w1[2][122] ) );
  XNOR U6158 ( .A(\w3[1][124] ), .B(\w3[1][120] ), .Z(n4319) );
  XNOR U6159 ( .A(n4320), .B(n4319), .Z(n4657) );
  XOR U6160 ( .A(n4657), .B(key[379]), .Z(n4323) );
  XNOR U6161 ( .A(\w3[1][99] ), .B(n4321), .Z(n4322) );
  XNOR U6162 ( .A(n4323), .B(n4322), .Z(\w1[2][123] ) );
  XOR U6163 ( .A(n4324), .B(key[380]), .Z(n4327) );
  XNOR U6164 ( .A(n4325), .B(\w3[1][100] ), .Z(n4326) );
  XNOR U6165 ( .A(n4327), .B(n4326), .Z(\w1[2][124] ) );
  XOR U6166 ( .A(\w3[1][118] ), .B(key[381]), .Z(n4330) );
  XNOR U6167 ( .A(n4328), .B(\w3[1][126] ), .Z(n4329) );
  XNOR U6168 ( .A(n4330), .B(n4329), .Z(n4331) );
  XOR U6169 ( .A(\w3[1][101] ), .B(n4331), .Z(\w1[2][125] ) );
  XOR U6170 ( .A(n4332), .B(key[382]), .Z(n4335) );
  XNOR U6171 ( .A(\w3[1][102] ), .B(n4333), .Z(n4334) );
  XNOR U6172 ( .A(n4335), .B(n4334), .Z(\w1[2][126] ) );
  XOR U6173 ( .A(n4646), .B(key[383]), .Z(n4338) );
  XNOR U6174 ( .A(\w3[1][103] ), .B(n4336), .Z(n4337) );
  XNOR U6175 ( .A(n4338), .B(n4337), .Z(\w1[2][127] ) );
  XOR U6176 ( .A(\w3[1][13] ), .B(\w3[1][28] ), .Z(n4340) );
  XNOR U6177 ( .A(\w3[1][8] ), .B(\w3[1][4] ), .Z(n4339) );
  XNOR U6178 ( .A(n4340), .B(n4339), .Z(n4362) );
  XOR U6179 ( .A(n4362), .B(key[268]), .Z(n4342) );
  XOR U6180 ( .A(\w3[1][0] ), .B(\w3[1][5] ), .Z(n4467) );
  XNOR U6181 ( .A(\w3[1][20] ), .B(n4467), .Z(n4341) );
  XNOR U6182 ( .A(n4342), .B(n4341), .Z(\w1[2][12] ) );
  XOR U6183 ( .A(\w3[1][14] ), .B(\w3[1][6] ), .Z(n4344) );
  XOR U6184 ( .A(\w3[1][5] ), .B(\w3[1][29] ), .Z(n4365) );
  XNOR U6185 ( .A(n4365), .B(key[269]), .Z(n4343) );
  XNOR U6186 ( .A(n4344), .B(n4343), .Z(n4345) );
  XOR U6187 ( .A(\w3[1][21] ), .B(n4345), .Z(\w1[2][13] ) );
  XOR U6188 ( .A(\w3[1][6] ), .B(\w3[1][30] ), .Z(n4508) );
  XNOR U6189 ( .A(\w3[1][8] ), .B(\w3[1][15] ), .Z(n4373) );
  XNOR U6190 ( .A(n4508), .B(n4373), .Z(n4368) );
  XOR U6191 ( .A(n4368), .B(key[270]), .Z(n4347) );
  XOR U6192 ( .A(\w3[1][0] ), .B(\w3[1][7] ), .Z(n4543) );
  XNOR U6193 ( .A(\w3[1][22] ), .B(n4543), .Z(n4346) );
  XNOR U6194 ( .A(n4347), .B(n4346), .Z(\w1[2][14] ) );
  XOR U6195 ( .A(\w3[1][7] ), .B(\w3[1][31] ), .Z(n4371) );
  XOR U6196 ( .A(n4371), .B(key[271]), .Z(n4349) );
  XOR U6197 ( .A(\w3[1][8] ), .B(\w3[1][0] ), .Z(n4375) );
  XNOR U6198 ( .A(\w3[1][23] ), .B(n4375), .Z(n4348) );
  XNOR U6199 ( .A(n4349), .B(n4348), .Z(\w1[2][15] ) );
  XOR U6200 ( .A(\w3[1][17] ), .B(\w3[1][9] ), .Z(n4379) );
  XOR U6201 ( .A(n4379), .B(key[272]), .Z(n4351) );
  XNOR U6202 ( .A(\w3[1][24] ), .B(n4375), .Z(n4350) );
  XNOR U6203 ( .A(n4351), .B(n4350), .Z(\w1[2][16] ) );
  XOR U6204 ( .A(\w3[1][18] ), .B(\w3[1][10] ), .Z(n4399) );
  XOR U6205 ( .A(n4399), .B(key[273]), .Z(n4353) );
  XNOR U6206 ( .A(n4664), .B(\w3[1][9] ), .Z(n4352) );
  XNOR U6207 ( .A(n4353), .B(n4352), .Z(\w1[2][17] ) );
  XOR U6208 ( .A(\w3[1][11] ), .B(\w3[1][19] ), .Z(n4387) );
  XOR U6209 ( .A(n4387), .B(key[274]), .Z(n4355) );
  XNOR U6210 ( .A(n4359), .B(\w3[1][10] ), .Z(n4354) );
  XNOR U6211 ( .A(n4355), .B(n4354), .Z(\w1[2][18] ) );
  XOR U6212 ( .A(\w3[1][16] ), .B(\w3[1][20] ), .Z(n4388) );
  XOR U6213 ( .A(n4388), .B(key[275]), .Z(n4358) );
  XNOR U6214 ( .A(\w3[1][11] ), .B(n4356), .Z(n4357) );
  XNOR U6215 ( .A(n4358), .B(n4357), .Z(\w1[2][19] ) );
  XOR U6216 ( .A(n4379), .B(key[257]), .Z(n4361) );
  XNOR U6217 ( .A(\w3[1][25] ), .B(n4359), .Z(n4360) );
  XNOR U6218 ( .A(n4361), .B(n4360), .Z(\w1[2][1] ) );
  XOR U6219 ( .A(\w3[1][16] ), .B(\w3[1][21] ), .Z(n4393) );
  XOR U6220 ( .A(n4393), .B(key[276]), .Z(n4364) );
  XNOR U6221 ( .A(\w3[1][12] ), .B(n4362), .Z(n4363) );
  XNOR U6222 ( .A(n4364), .B(n4363), .Z(\w1[2][20] ) );
  XOR U6223 ( .A(\w3[1][14] ), .B(\w3[1][22] ), .Z(n4403) );
  XOR U6224 ( .A(n4403), .B(key[277]), .Z(n4367) );
  XNOR U6225 ( .A(\w3[1][13] ), .B(n4365), .Z(n4366) );
  XNOR U6226 ( .A(n4367), .B(n4366), .Z(\w1[2][21] ) );
  XOR U6227 ( .A(\w3[1][16] ), .B(\w3[1][23] ), .Z(n4404) );
  XOR U6228 ( .A(n4404), .B(key[278]), .Z(n4370) );
  XNOR U6229 ( .A(\w3[1][14] ), .B(n4368), .Z(n4369) );
  XNOR U6230 ( .A(n4370), .B(n4369), .Z(\w1[2][22] ) );
  XNOR U6231 ( .A(n4371), .B(key[279]), .Z(n4372) );
  XNOR U6232 ( .A(n4373), .B(n4372), .Z(n4374) );
  XNOR U6233 ( .A(\w3[1][16] ), .B(n4374), .Z(\w1[2][23] ) );
  XOR U6234 ( .A(\w3[1][17] ), .B(key[280]), .Z(n4377) );
  XNOR U6235 ( .A(\w3[1][25] ), .B(n4375), .Z(n4376) );
  XNOR U6236 ( .A(n4377), .B(n4376), .Z(n4378) );
  XOR U6237 ( .A(\w3[1][16] ), .B(n4378), .Z(\w1[2][24] ) );
  XOR U6238 ( .A(n4379), .B(key[281]), .Z(n4381) );
  XNOR U6239 ( .A(\w3[1][1] ), .B(\w3[1][26] ), .Z(n4380) );
  XNOR U6240 ( .A(n4381), .B(n4380), .Z(n4382) );
  XOR U6241 ( .A(\w3[1][18] ), .B(n4382), .Z(\w1[2][25] ) );
  XOR U6242 ( .A(n4399), .B(key[282]), .Z(n4384) );
  XNOR U6243 ( .A(\w3[1][2] ), .B(\w3[1][19] ), .Z(n4383) );
  XNOR U6244 ( .A(n4384), .B(n4383), .Z(n4385) );
  XOR U6245 ( .A(\w3[1][27] ), .B(n4385), .Z(\w1[2][26] ) );
  XNOR U6246 ( .A(\w3[1][24] ), .B(\w3[1][28] ), .Z(n4386) );
  XNOR U6247 ( .A(n4387), .B(n4386), .Z(n4429) );
  XOR U6248 ( .A(n4429), .B(key[283]), .Z(n4390) );
  XNOR U6249 ( .A(\w3[1][3] ), .B(n4388), .Z(n4389) );
  XNOR U6250 ( .A(n4390), .B(n4389), .Z(\w1[2][27] ) );
  XOR U6251 ( .A(\w3[1][20] ), .B(\w3[1][29] ), .Z(n4392) );
  XNOR U6252 ( .A(\w3[1][24] ), .B(\w3[1][12] ), .Z(n4391) );
  XNOR U6253 ( .A(n4392), .B(n4391), .Z(n4466) );
  XOR U6254 ( .A(n4466), .B(key[284]), .Z(n4395) );
  XNOR U6255 ( .A(\w3[1][4] ), .B(n4393), .Z(n4394) );
  XNOR U6256 ( .A(n4395), .B(n4394), .Z(\w1[2][28] ) );
  XOR U6257 ( .A(\w3[1][13] ), .B(\w3[1][21] ), .Z(n4507) );
  XOR U6258 ( .A(n4507), .B(key[285]), .Z(n4397) );
  XNOR U6259 ( .A(\w3[1][22] ), .B(\w3[1][30] ), .Z(n4396) );
  XNOR U6260 ( .A(n4397), .B(n4396), .Z(n4398) );
  XOR U6261 ( .A(\w3[1][5] ), .B(n4398), .Z(\w1[2][29] ) );
  XOR U6262 ( .A(n4399), .B(key[258]), .Z(n4402) );
  XNOR U6263 ( .A(\w3[1][26] ), .B(n4400), .Z(n4401) );
  XNOR U6264 ( .A(n4402), .B(n4401), .Z(\w1[2][2] ) );
  XNOR U6265 ( .A(\w3[1][24] ), .B(\w3[1][31] ), .Z(n4581) );
  XNOR U6266 ( .A(n4403), .B(n4581), .Z(n4542) );
  XOR U6267 ( .A(n4542), .B(key[286]), .Z(n4406) );
  XNOR U6268 ( .A(\w3[1][6] ), .B(n4404), .Z(n4405) );
  XNOR U6269 ( .A(n4406), .B(n4405), .Z(\w1[2][30] ) );
  XOR U6270 ( .A(\w3[1][15] ), .B(\w3[1][23] ), .Z(n4579) );
  XOR U6271 ( .A(n4579), .B(key[287]), .Z(n4408) );
  XNOR U6272 ( .A(n4620), .B(\w3[1][7] ), .Z(n4407) );
  XNOR U6273 ( .A(n4408), .B(n4407), .Z(\w1[2][31] ) );
  XOR U6274 ( .A(\w3[1][33] ), .B(\w3[1][57] ), .Z(n4463) );
  XOR U6275 ( .A(n4463), .B(key[288]), .Z(n4410) );
  XOR U6276 ( .A(\w3[1][48] ), .B(\w3[1][56] ), .Z(n4524) );
  XNOR U6277 ( .A(n4524), .B(\w3[1][40] ), .Z(n4409) );
  XNOR U6278 ( .A(n4410), .B(n4409), .Z(\w1[2][32] ) );
  XOR U6279 ( .A(\w3[1][34] ), .B(\w3[1][58] ), .Z(n4471) );
  XOR U6280 ( .A(n4471), .B(key[289]), .Z(n4412) );
  XOR U6281 ( .A(\w3[1][41] ), .B(\w3[1][49] ), .Z(n4495) );
  XNOR U6282 ( .A(\w3[1][57] ), .B(n4495), .Z(n4411) );
  XNOR U6283 ( .A(n4412), .B(n4411), .Z(\w1[2][33] ) );
  XOR U6284 ( .A(\w3[1][35] ), .B(\w3[1][59] ), .Z(n4442) );
  XOR U6285 ( .A(n4442), .B(key[290]), .Z(n4414) );
  XOR U6286 ( .A(\w3[1][42] ), .B(\w3[1][50] ), .Z(n4499) );
  XNOR U6287 ( .A(\w3[1][58] ), .B(n4499), .Z(n4413) );
  XNOR U6288 ( .A(n4414), .B(n4413), .Z(\w1[2][34] ) );
  XOR U6289 ( .A(\w3[1][36] ), .B(\w3[1][32] ), .Z(n4444) );
  XOR U6290 ( .A(n4444), .B(key[291]), .Z(n4417) );
  XOR U6291 ( .A(\w3[1][43] ), .B(\w3[1][51] ), .Z(n4470) );
  XNOR U6292 ( .A(\w3[1][56] ), .B(n4470), .Z(n4415) );
  XNOR U6293 ( .A(\w3[1][60] ), .B(n4415), .Z(n4504) );
  XNOR U6294 ( .A(\w3[1][59] ), .B(n4504), .Z(n4416) );
  XNOR U6295 ( .A(n4417), .B(n4416), .Z(\w1[2][35] ) );
  XOR U6296 ( .A(\w3[1][32] ), .B(\w3[1][37] ), .Z(n4449) );
  XOR U6297 ( .A(n4449), .B(key[292]), .Z(n4421) );
  XOR U6298 ( .A(\w3[1][52] ), .B(\w3[1][61] ), .Z(n4419) );
  XNOR U6299 ( .A(\w3[1][56] ), .B(\w3[1][44] ), .Z(n4418) );
  XNOR U6300 ( .A(n4419), .B(n4418), .Z(n4512) );
  XNOR U6301 ( .A(\w3[1][60] ), .B(n4512), .Z(n4420) );
  XNOR U6302 ( .A(n4421), .B(n4420), .Z(\w1[2][36] ) );
  XOR U6303 ( .A(\w3[1][38] ), .B(\w3[1][62] ), .Z(n4455) );
  XOR U6304 ( .A(n4455), .B(key[293]), .Z(n4423) );
  XOR U6305 ( .A(\w3[1][45] ), .B(\w3[1][53] ), .Z(n4515) );
  XNOR U6306 ( .A(\w3[1][61] ), .B(n4515), .Z(n4422) );
  XNOR U6307 ( .A(n4423), .B(n4422), .Z(\w1[2][37] ) );
  XOR U6308 ( .A(\w3[1][32] ), .B(\w3[1][39] ), .Z(n4456) );
  XOR U6309 ( .A(n4456), .B(key[294]), .Z(n4425) );
  XOR U6310 ( .A(\w3[1][46] ), .B(\w3[1][54] ), .Z(n4481) );
  XNOR U6311 ( .A(\w3[1][56] ), .B(\w3[1][63] ), .Z(n4427) );
  XNOR U6312 ( .A(n4481), .B(n4427), .Z(n4520) );
  XNOR U6313 ( .A(\w3[1][62] ), .B(n4520), .Z(n4424) );
  XNOR U6314 ( .A(n4425), .B(n4424), .Z(\w1[2][38] ) );
  XOR U6315 ( .A(\w3[1][47] ), .B(\w3[1][55] ), .Z(n4523) );
  XNOR U6316 ( .A(n4523), .B(key[295]), .Z(n4426) );
  XNOR U6317 ( .A(n4427), .B(n4426), .Z(n4428) );
  XNOR U6318 ( .A(\w3[1][32] ), .B(n4428), .Z(\w1[2][39] ) );
  XOR U6319 ( .A(n4429), .B(key[259]), .Z(n4432) );
  XNOR U6320 ( .A(n4430), .B(\w3[1][27] ), .Z(n4431) );
  XNOR U6321 ( .A(n4432), .B(n4431), .Z(\w1[2][3] ) );
  XOR U6322 ( .A(\w3[1][32] ), .B(key[296]), .Z(n4434) );
  XNOR U6323 ( .A(\w3[1][33] ), .B(\w3[1][41] ), .Z(n4433) );
  XNOR U6324 ( .A(n4434), .B(n4433), .Z(n4435) );
  XOR U6325 ( .A(n4524), .B(n4435), .Z(\w1[2][40] ) );
  XOR U6326 ( .A(\w3[1][42] ), .B(key[297]), .Z(n4437) );
  XNOR U6327 ( .A(\w3[1][49] ), .B(\w3[1][34] ), .Z(n4436) );
  XNOR U6328 ( .A(n4437), .B(n4436), .Z(n4438) );
  XOR U6329 ( .A(n4463), .B(n4438), .Z(\w1[2][41] ) );
  XOR U6330 ( .A(\w3[1][43] ), .B(key[298]), .Z(n4440) );
  XNOR U6331 ( .A(\w3[1][50] ), .B(\w3[1][35] ), .Z(n4439) );
  XNOR U6332 ( .A(n4440), .B(n4439), .Z(n4441) );
  XOR U6333 ( .A(n4471), .B(n4441), .Z(\w1[2][42] ) );
  XNOR U6334 ( .A(\w3[1][40] ), .B(n4442), .Z(n4443) );
  XNOR U6335 ( .A(\w3[1][44] ), .B(n4443), .Z(n4474) );
  XOR U6336 ( .A(n4474), .B(key[299]), .Z(n4446) );
  XNOR U6337 ( .A(\w3[1][51] ), .B(n4444), .Z(n4445) );
  XNOR U6338 ( .A(n4446), .B(n4445), .Z(\w1[2][43] ) );
  XOR U6339 ( .A(\w3[1][36] ), .B(\w3[1][45] ), .Z(n4448) );
  XNOR U6340 ( .A(\w3[1][40] ), .B(\w3[1][60] ), .Z(n4447) );
  XNOR U6341 ( .A(n4448), .B(n4447), .Z(n4477) );
  XOR U6342 ( .A(n4477), .B(key[300]), .Z(n4451) );
  XNOR U6343 ( .A(\w3[1][52] ), .B(n4449), .Z(n4450) );
  XNOR U6344 ( .A(n4451), .B(n4450), .Z(\w1[2][44] ) );
  XOR U6345 ( .A(\w3[1][61] ), .B(\w3[1][37] ), .Z(n4480) );
  XOR U6346 ( .A(n4480), .B(key[301]), .Z(n4453) );
  XNOR U6347 ( .A(\w3[1][38] ), .B(\w3[1][46] ), .Z(n4452) );
  XNOR U6348 ( .A(n4453), .B(n4452), .Z(n4454) );
  XOR U6349 ( .A(\w3[1][53] ), .B(n4454), .Z(\w1[2][45] ) );
  XNOR U6350 ( .A(\w3[1][40] ), .B(\w3[1][47] ), .Z(n4489) );
  XNOR U6351 ( .A(n4455), .B(n4489), .Z(n4484) );
  XOR U6352 ( .A(n4484), .B(key[302]), .Z(n4458) );
  XNOR U6353 ( .A(\w3[1][54] ), .B(n4456), .Z(n4457) );
  XNOR U6354 ( .A(n4458), .B(n4457), .Z(\w1[2][46] ) );
  XOR U6355 ( .A(\w3[1][63] ), .B(\w3[1][39] ), .Z(n4487) );
  XOR U6356 ( .A(n4487), .B(key[303]), .Z(n4460) );
  XOR U6357 ( .A(\w3[1][40] ), .B(\w3[1][32] ), .Z(n4491) );
  XNOR U6358 ( .A(\w3[1][55] ), .B(n4491), .Z(n4459) );
  XNOR U6359 ( .A(n4460), .B(n4459), .Z(\w1[2][47] ) );
  XOR U6360 ( .A(n4491), .B(key[304]), .Z(n4462) );
  XNOR U6361 ( .A(\w3[1][56] ), .B(n4495), .Z(n4461) );
  XNOR U6362 ( .A(n4462), .B(n4461), .Z(\w1[2][48] ) );
  XOR U6363 ( .A(n4499), .B(key[305]), .Z(n4465) );
  XNOR U6364 ( .A(n4463), .B(\w3[1][41] ), .Z(n4464) );
  XNOR U6365 ( .A(n4465), .B(n4464), .Z(\w1[2][49] ) );
  XOR U6366 ( .A(n4466), .B(key[260]), .Z(n4469) );
  XNOR U6367 ( .A(n4467), .B(\w3[1][28] ), .Z(n4468) );
  XNOR U6368 ( .A(n4469), .B(n4468), .Z(\w1[2][4] ) );
  XOR U6369 ( .A(n4470), .B(key[306]), .Z(n4473) );
  XNOR U6370 ( .A(n4471), .B(\w3[1][42] ), .Z(n4472) );
  XNOR U6371 ( .A(n4473), .B(n4472), .Z(\w1[2][50] ) );
  XOR U6372 ( .A(\w3[1][48] ), .B(\w3[1][52] ), .Z(n4503) );
  XOR U6373 ( .A(n4503), .B(key[307]), .Z(n4476) );
  XNOR U6374 ( .A(\w3[1][43] ), .B(n4474), .Z(n4475) );
  XNOR U6375 ( .A(n4476), .B(n4475), .Z(\w1[2][51] ) );
  XOR U6376 ( .A(\w3[1][48] ), .B(\w3[1][53] ), .Z(n4511) );
  XOR U6377 ( .A(n4511), .B(key[308]), .Z(n4479) );
  XNOR U6378 ( .A(\w3[1][44] ), .B(n4477), .Z(n4478) );
  XNOR U6379 ( .A(n4479), .B(n4478), .Z(\w1[2][52] ) );
  XOR U6380 ( .A(n4480), .B(key[309]), .Z(n4483) );
  XNOR U6381 ( .A(\w3[1][45] ), .B(n4481), .Z(n4482) );
  XNOR U6382 ( .A(n4483), .B(n4482), .Z(\w1[2][53] ) );
  XOR U6383 ( .A(\w3[1][48] ), .B(\w3[1][55] ), .Z(n4519) );
  XOR U6384 ( .A(n4519), .B(key[310]), .Z(n4486) );
  XNOR U6385 ( .A(\w3[1][46] ), .B(n4484), .Z(n4485) );
  XNOR U6386 ( .A(n4486), .B(n4485), .Z(\w1[2][54] ) );
  XNOR U6387 ( .A(n4487), .B(key[311]), .Z(n4488) );
  XNOR U6388 ( .A(n4489), .B(n4488), .Z(n4490) );
  XNOR U6389 ( .A(\w3[1][48] ), .B(n4490), .Z(\w1[2][55] ) );
  XOR U6390 ( .A(n4491), .B(key[312]), .Z(n4493) );
  XNOR U6391 ( .A(\w3[1][48] ), .B(\w3[1][49] ), .Z(n4492) );
  XNOR U6392 ( .A(n4493), .B(n4492), .Z(n4494) );
  XOR U6393 ( .A(\w3[1][57] ), .B(n4494), .Z(\w1[2][56] ) );
  XOR U6394 ( .A(\w3[1][50] ), .B(key[313]), .Z(n4497) );
  XNOR U6395 ( .A(n4495), .B(\w3[1][58] ), .Z(n4496) );
  XNOR U6396 ( .A(n4497), .B(n4496), .Z(n4498) );
  XOR U6397 ( .A(\w3[1][33] ), .B(n4498), .Z(\w1[2][57] ) );
  XOR U6398 ( .A(\w3[1][51] ), .B(key[314]), .Z(n4501) );
  XNOR U6399 ( .A(n4499), .B(\w3[1][59] ), .Z(n4500) );
  XNOR U6400 ( .A(n4501), .B(n4500), .Z(n4502) );
  XOR U6401 ( .A(\w3[1][34] ), .B(n4502), .Z(\w1[2][58] ) );
  XOR U6402 ( .A(n4503), .B(key[315]), .Z(n4506) );
  XNOR U6403 ( .A(\w3[1][35] ), .B(n4504), .Z(n4505) );
  XNOR U6404 ( .A(n4506), .B(n4505), .Z(\w1[2][59] ) );
  XOR U6405 ( .A(n4507), .B(key[261]), .Z(n4510) );
  XNOR U6406 ( .A(\w3[1][29] ), .B(n4508), .Z(n4509) );
  XNOR U6407 ( .A(n4510), .B(n4509), .Z(\w1[2][5] ) );
  XOR U6408 ( .A(n4511), .B(key[316]), .Z(n4514) );
  XNOR U6409 ( .A(\w3[1][36] ), .B(n4512), .Z(n4513) );
  XNOR U6410 ( .A(n4514), .B(n4513), .Z(\w1[2][60] ) );
  XOR U6411 ( .A(\w3[1][54] ), .B(key[317]), .Z(n4517) );
  XNOR U6412 ( .A(n4515), .B(\w3[1][62] ), .Z(n4516) );
  XNOR U6413 ( .A(n4517), .B(n4516), .Z(n4518) );
  XOR U6414 ( .A(\w3[1][37] ), .B(n4518), .Z(\w1[2][61] ) );
  XOR U6415 ( .A(n4519), .B(key[318]), .Z(n4522) );
  XNOR U6416 ( .A(\w3[1][38] ), .B(n4520), .Z(n4521) );
  XNOR U6417 ( .A(n4522), .B(n4521), .Z(\w1[2][62] ) );
  XOR U6418 ( .A(n4523), .B(key[319]), .Z(n4526) );
  XNOR U6419 ( .A(n4524), .B(\w3[1][39] ), .Z(n4525) );
  XNOR U6420 ( .A(n4526), .B(n4525), .Z(\w1[2][63] ) );
  XOR U6421 ( .A(\w3[1][65] ), .B(\w3[1][89] ), .Z(n4585) );
  XOR U6422 ( .A(n4585), .B(key[320]), .Z(n4528) );
  XOR U6423 ( .A(\w3[1][80] ), .B(\w3[1][88] ), .Z(n4642) );
  XNOR U6424 ( .A(n4642), .B(\w3[1][72] ), .Z(n4527) );
  XNOR U6425 ( .A(n4528), .B(n4527), .Z(\w1[2][64] ) );
  XOR U6426 ( .A(\w3[1][66] ), .B(\w3[1][90] ), .Z(n4589) );
  XOR U6427 ( .A(n4589), .B(key[321]), .Z(n4530) );
  XOR U6428 ( .A(\w3[1][73] ), .B(\w3[1][81] ), .Z(n4613) );
  XNOR U6429 ( .A(\w3[1][89] ), .B(n4613), .Z(n4529) );
  XNOR U6430 ( .A(n4530), .B(n4529), .Z(\w1[2][65] ) );
  XOR U6431 ( .A(\w3[1][67] ), .B(\w3[1][91] ), .Z(n4560) );
  XOR U6432 ( .A(n4560), .B(key[322]), .Z(n4532) );
  XOR U6433 ( .A(\w3[1][74] ), .B(\w3[1][82] ), .Z(n4621) );
  XNOR U6434 ( .A(\w3[1][90] ), .B(n4621), .Z(n4531) );
  XNOR U6435 ( .A(n4532), .B(n4531), .Z(\w1[2][66] ) );
  XOR U6436 ( .A(\w3[1][68] ), .B(\w3[1][64] ), .Z(n4562) );
  XOR U6437 ( .A(n4562), .B(key[323]), .Z(n4535) );
  XOR U6438 ( .A(\w3[1][75] ), .B(\w3[1][83] ), .Z(n4588) );
  XNOR U6439 ( .A(\w3[1][88] ), .B(n4588), .Z(n4533) );
  XNOR U6440 ( .A(\w3[1][92] ), .B(n4533), .Z(n4626) );
  XNOR U6441 ( .A(\w3[1][91] ), .B(n4626), .Z(n4534) );
  XNOR U6442 ( .A(n4535), .B(n4534), .Z(\w1[2][67] ) );
  XOR U6443 ( .A(\w3[1][64] ), .B(\w3[1][69] ), .Z(n4567) );
  XOR U6444 ( .A(n4567), .B(key[324]), .Z(n4539) );
  XOR U6445 ( .A(\w3[1][84] ), .B(\w3[1][93] ), .Z(n4537) );
  XNOR U6446 ( .A(\w3[1][88] ), .B(\w3[1][76] ), .Z(n4536) );
  XNOR U6447 ( .A(n4537), .B(n4536), .Z(n4630) );
  XNOR U6448 ( .A(\w3[1][92] ), .B(n4630), .Z(n4538) );
  XNOR U6449 ( .A(n4539), .B(n4538), .Z(\w1[2][68] ) );
  XOR U6450 ( .A(\w3[1][70] ), .B(\w3[1][94] ), .Z(n4573) );
  XOR U6451 ( .A(n4573), .B(key[325]), .Z(n4541) );
  XOR U6452 ( .A(\w3[1][77] ), .B(\w3[1][85] ), .Z(n4633) );
  XNOR U6453 ( .A(\w3[1][93] ), .B(n4633), .Z(n4540) );
  XNOR U6454 ( .A(n4541), .B(n4540), .Z(\w1[2][69] ) );
  XOR U6455 ( .A(n4542), .B(key[262]), .Z(n4545) );
  XNOR U6456 ( .A(n4543), .B(\w3[1][30] ), .Z(n4544) );
  XNOR U6457 ( .A(n4545), .B(n4544), .Z(\w1[2][6] ) );
  XOR U6458 ( .A(\w3[1][64] ), .B(\w3[1][71] ), .Z(n4574) );
  XOR U6459 ( .A(n4574), .B(key[326]), .Z(n4547) );
  XOR U6460 ( .A(\w3[1][78] ), .B(\w3[1][86] ), .Z(n4599) );
  XNOR U6461 ( .A(\w3[1][88] ), .B(\w3[1][95] ), .Z(n4549) );
  XNOR U6462 ( .A(n4599), .B(n4549), .Z(n4638) );
  XNOR U6463 ( .A(\w3[1][94] ), .B(n4638), .Z(n4546) );
  XNOR U6464 ( .A(n4547), .B(n4546), .Z(\w1[2][70] ) );
  XOR U6465 ( .A(\w3[1][79] ), .B(\w3[1][87] ), .Z(n4641) );
  XNOR U6466 ( .A(n4641), .B(key[327]), .Z(n4548) );
  XNOR U6467 ( .A(n4549), .B(n4548), .Z(n4550) );
  XNOR U6468 ( .A(\w3[1][64] ), .B(n4550), .Z(\w1[2][71] ) );
  XOR U6469 ( .A(\w3[1][64] ), .B(key[328]), .Z(n4552) );
  XNOR U6470 ( .A(\w3[1][65] ), .B(\w3[1][73] ), .Z(n4551) );
  XNOR U6471 ( .A(n4552), .B(n4551), .Z(n4553) );
  XOR U6472 ( .A(n4642), .B(n4553), .Z(\w1[2][72] ) );
  XOR U6473 ( .A(\w3[1][74] ), .B(key[329]), .Z(n4555) );
  XNOR U6474 ( .A(\w3[1][81] ), .B(\w3[1][66] ), .Z(n4554) );
  XNOR U6475 ( .A(n4555), .B(n4554), .Z(n4556) );
  XOR U6476 ( .A(n4585), .B(n4556), .Z(\w1[2][73] ) );
  XOR U6477 ( .A(\w3[1][75] ), .B(key[330]), .Z(n4558) );
  XNOR U6478 ( .A(\w3[1][82] ), .B(\w3[1][67] ), .Z(n4557) );
  XNOR U6479 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U6480 ( .A(n4589), .B(n4559), .Z(\w1[2][74] ) );
  XNOR U6481 ( .A(\w3[1][72] ), .B(n4560), .Z(n4561) );
  XNOR U6482 ( .A(\w3[1][76] ), .B(n4561), .Z(n4592) );
  XOR U6483 ( .A(n4592), .B(key[331]), .Z(n4564) );
  XNOR U6484 ( .A(\w3[1][83] ), .B(n4562), .Z(n4563) );
  XNOR U6485 ( .A(n4564), .B(n4563), .Z(\w1[2][75] ) );
  XOR U6486 ( .A(\w3[1][68] ), .B(\w3[1][77] ), .Z(n4566) );
  XNOR U6487 ( .A(\w3[1][72] ), .B(\w3[1][92] ), .Z(n4565) );
  XNOR U6488 ( .A(n4566), .B(n4565), .Z(n4595) );
  XOR U6489 ( .A(n4595), .B(key[332]), .Z(n4569) );
  XNOR U6490 ( .A(\w3[1][84] ), .B(n4567), .Z(n4568) );
  XNOR U6491 ( .A(n4569), .B(n4568), .Z(\w1[2][76] ) );
  XOR U6492 ( .A(\w3[1][93] ), .B(\w3[1][69] ), .Z(n4598) );
  XOR U6493 ( .A(n4598), .B(key[333]), .Z(n4571) );
  XNOR U6494 ( .A(\w3[1][70] ), .B(\w3[1][78] ), .Z(n4570) );
  XNOR U6495 ( .A(n4571), .B(n4570), .Z(n4572) );
  XOR U6496 ( .A(\w3[1][85] ), .B(n4572), .Z(\w1[2][77] ) );
  XNOR U6497 ( .A(\w3[1][72] ), .B(\w3[1][79] ), .Z(n4607) );
  XNOR U6498 ( .A(n4573), .B(n4607), .Z(n4602) );
  XOR U6499 ( .A(n4602), .B(key[334]), .Z(n4576) );
  XNOR U6500 ( .A(\w3[1][86] ), .B(n4574), .Z(n4575) );
  XNOR U6501 ( .A(n4576), .B(n4575), .Z(\w1[2][78] ) );
  XOR U6502 ( .A(\w3[1][95] ), .B(\w3[1][71] ), .Z(n4605) );
  XOR U6503 ( .A(n4605), .B(key[335]), .Z(n4578) );
  XOR U6504 ( .A(\w3[1][72] ), .B(\w3[1][64] ), .Z(n4609) );
  XNOR U6505 ( .A(\w3[1][87] ), .B(n4609), .Z(n4577) );
  XNOR U6506 ( .A(n4578), .B(n4577), .Z(\w1[2][79] ) );
  XNOR U6507 ( .A(n4579), .B(key[263]), .Z(n4580) );
  XNOR U6508 ( .A(n4581), .B(n4580), .Z(n4582) );
  XNOR U6509 ( .A(\w3[1][0] ), .B(n4582), .Z(\w1[2][7] ) );
  XOR U6510 ( .A(n4609), .B(key[336]), .Z(n4584) );
  XNOR U6511 ( .A(\w3[1][88] ), .B(n4613), .Z(n4583) );
  XNOR U6512 ( .A(n4584), .B(n4583), .Z(\w1[2][80] ) );
  XOR U6513 ( .A(n4621), .B(key[337]), .Z(n4587) );
  XNOR U6514 ( .A(n4585), .B(\w3[1][73] ), .Z(n4586) );
  XNOR U6515 ( .A(n4587), .B(n4586), .Z(\w1[2][81] ) );
  XOR U6516 ( .A(n4588), .B(key[338]), .Z(n4591) );
  XNOR U6517 ( .A(n4589), .B(\w3[1][74] ), .Z(n4590) );
  XNOR U6518 ( .A(n4591), .B(n4590), .Z(\w1[2][82] ) );
  XOR U6519 ( .A(\w3[1][80] ), .B(\w3[1][84] ), .Z(n4625) );
  XOR U6520 ( .A(n4625), .B(key[339]), .Z(n4594) );
  XNOR U6521 ( .A(\w3[1][75] ), .B(n4592), .Z(n4593) );
  XNOR U6522 ( .A(n4594), .B(n4593), .Z(\w1[2][83] ) );
  XOR U6523 ( .A(\w3[1][80] ), .B(\w3[1][85] ), .Z(n4629) );
  XOR U6524 ( .A(n4629), .B(key[340]), .Z(n4597) );
  XNOR U6525 ( .A(\w3[1][76] ), .B(n4595), .Z(n4596) );
  XNOR U6526 ( .A(n4597), .B(n4596), .Z(\w1[2][84] ) );
  XOR U6527 ( .A(n4598), .B(key[341]), .Z(n4601) );
  XNOR U6528 ( .A(\w3[1][77] ), .B(n4599), .Z(n4600) );
  XNOR U6529 ( .A(n4601), .B(n4600), .Z(\w1[2][85] ) );
  XOR U6530 ( .A(\w3[1][80] ), .B(\w3[1][87] ), .Z(n4637) );
  XOR U6531 ( .A(n4637), .B(key[342]), .Z(n4604) );
  XNOR U6532 ( .A(\w3[1][78] ), .B(n4602), .Z(n4603) );
  XNOR U6533 ( .A(n4604), .B(n4603), .Z(\w1[2][86] ) );
  XNOR U6534 ( .A(n4605), .B(key[343]), .Z(n4606) );
  XNOR U6535 ( .A(n4607), .B(n4606), .Z(n4608) );
  XNOR U6536 ( .A(\w3[1][80] ), .B(n4608), .Z(\w1[2][87] ) );
  XOR U6537 ( .A(n4609), .B(key[344]), .Z(n4611) );
  XNOR U6538 ( .A(\w3[1][80] ), .B(\w3[1][81] ), .Z(n4610) );
  XNOR U6539 ( .A(n4611), .B(n4610), .Z(n4612) );
  XOR U6540 ( .A(\w3[1][89] ), .B(n4612), .Z(\w1[2][88] ) );
  XOR U6541 ( .A(\w3[1][82] ), .B(key[345]), .Z(n4615) );
  XNOR U6542 ( .A(n4613), .B(\w3[1][90] ), .Z(n4614) );
  XNOR U6543 ( .A(n4615), .B(n4614), .Z(n4616) );
  XOR U6544 ( .A(\w3[1][65] ), .B(n4616), .Z(\w1[2][89] ) );
  XOR U6545 ( .A(\w3[1][9] ), .B(key[264]), .Z(n4618) );
  XNOR U6546 ( .A(\w3[1][1] ), .B(\w3[1][0] ), .Z(n4617) );
  XNOR U6547 ( .A(n4618), .B(n4617), .Z(n4619) );
  XOR U6548 ( .A(n4620), .B(n4619), .Z(\w1[2][8] ) );
  XOR U6549 ( .A(\w3[1][83] ), .B(key[346]), .Z(n4623) );
  XNOR U6550 ( .A(n4621), .B(\w3[1][91] ), .Z(n4622) );
  XNOR U6551 ( .A(n4623), .B(n4622), .Z(n4624) );
  XOR U6552 ( .A(\w3[1][66] ), .B(n4624), .Z(\w1[2][90] ) );
  XOR U6553 ( .A(n4625), .B(key[347]), .Z(n4628) );
  XNOR U6554 ( .A(\w3[1][67] ), .B(n4626), .Z(n4627) );
  XNOR U6555 ( .A(n4628), .B(n4627), .Z(\w1[2][91] ) );
  XOR U6556 ( .A(n4629), .B(key[348]), .Z(n4632) );
  XNOR U6557 ( .A(\w3[1][68] ), .B(n4630), .Z(n4631) );
  XNOR U6558 ( .A(n4632), .B(n4631), .Z(\w1[2][92] ) );
  XOR U6559 ( .A(\w3[1][86] ), .B(key[349]), .Z(n4635) );
  XNOR U6560 ( .A(n4633), .B(\w3[1][94] ), .Z(n4634) );
  XNOR U6561 ( .A(n4635), .B(n4634), .Z(n4636) );
  XOR U6562 ( .A(\w3[1][69] ), .B(n4636), .Z(\w1[2][93] ) );
  XOR U6563 ( .A(n4637), .B(key[350]), .Z(n4640) );
  XNOR U6564 ( .A(\w3[1][70] ), .B(n4638), .Z(n4639) );
  XNOR U6565 ( .A(n4640), .B(n4639), .Z(\w1[2][94] ) );
  XOR U6566 ( .A(n4641), .B(key[351]), .Z(n4644) );
  XNOR U6567 ( .A(n4642), .B(\w3[1][71] ), .Z(n4643) );
  XNOR U6568 ( .A(n4644), .B(n4643), .Z(\w1[2][95] ) );
  XOR U6569 ( .A(\w3[1][104] ), .B(key[352]), .Z(n4648) );
  XNOR U6570 ( .A(n4646), .B(n4645), .Z(n4647) );
  XNOR U6571 ( .A(n4648), .B(n4647), .Z(\w1[2][96] ) );
  XOR U6572 ( .A(n4649), .B(key[353]), .Z(n4652) );
  XNOR U6573 ( .A(\w3[1][121] ), .B(n4650), .Z(n4651) );
  XNOR U6574 ( .A(n4652), .B(n4651), .Z(\w1[2][97] ) );
  XOR U6575 ( .A(n4653), .B(key[354]), .Z(n4656) );
  XNOR U6576 ( .A(\w3[1][122] ), .B(n4654), .Z(n4655) );
  XNOR U6577 ( .A(n4656), .B(n4655), .Z(\w1[2][98] ) );
  XOR U6578 ( .A(n4657), .B(key[355]), .Z(n4660) );
  XNOR U6579 ( .A(n4658), .B(\w3[1][123] ), .Z(n4659) );
  XNOR U6580 ( .A(n4660), .B(n4659), .Z(\w1[2][99] ) );
  XOR U6581 ( .A(\w3[1][10] ), .B(key[265]), .Z(n4662) );
  XNOR U6582 ( .A(\w3[1][2] ), .B(\w3[1][17] ), .Z(n4661) );
  XNOR U6583 ( .A(n4662), .B(n4661), .Z(n4663) );
  XOR U6584 ( .A(n4664), .B(n4663), .Z(\w1[2][9] ) );
  XOR U6585 ( .A(\w3[2][8] ), .B(key[384]), .Z(n4666) );
  XOR U6586 ( .A(\w3[2][1] ), .B(\w3[2][25] ), .Z(n5088) );
  XOR U6587 ( .A(\w3[2][16] ), .B(\w3[2][24] ), .Z(n5044) );
  XNOR U6588 ( .A(n5088), .B(n5044), .Z(n4665) );
  XNOR U6589 ( .A(n4666), .B(n4665), .Z(\w1[3][0] ) );
  XOR U6590 ( .A(\w3[2][96] ), .B(\w3[2][101] ), .Z(n4690) );
  XOR U6591 ( .A(n4690), .B(key[484]), .Z(n4670) );
  XOR U6592 ( .A(\w3[2][116] ), .B(\w3[2][125] ), .Z(n4668) );
  XNOR U6593 ( .A(\w3[2][120] ), .B(\w3[2][108] ), .Z(n4667) );
  XNOR U6594 ( .A(n4668), .B(n4667), .Z(n4749) );
  XNOR U6595 ( .A(\w3[2][124] ), .B(n4749), .Z(n4669) );
  XNOR U6596 ( .A(n4670), .B(n4669), .Z(\w1[3][100] ) );
  XOR U6597 ( .A(\w3[2][102] ), .B(\w3[2][126] ), .Z(n4699) );
  XOR U6598 ( .A(n4699), .B(key[485]), .Z(n4672) );
  XOR U6599 ( .A(\w3[2][109] ), .B(\w3[2][117] ), .Z(n4752) );
  XNOR U6600 ( .A(\w3[2][125] ), .B(n4752), .Z(n4671) );
  XNOR U6601 ( .A(n4672), .B(n4671), .Z(\w1[3][101] ) );
  XOR U6602 ( .A(\w3[2][96] ), .B(\w3[2][103] ), .Z(n4700) );
  XOR U6603 ( .A(n4700), .B(key[486]), .Z(n4674) );
  XOR U6604 ( .A(\w3[2][110] ), .B(\w3[2][118] ), .Z(n4718) );
  XNOR U6605 ( .A(\w3[2][120] ), .B(\w3[2][127] ), .Z(n4676) );
  XNOR U6606 ( .A(n4718), .B(n4676), .Z(n4757) );
  XNOR U6607 ( .A(\w3[2][126] ), .B(n4757), .Z(n4673) );
  XNOR U6608 ( .A(n4674), .B(n4673), .Z(\w1[3][102] ) );
  XOR U6609 ( .A(\w3[2][111] ), .B(\w3[2][119] ), .Z(n4760) );
  XNOR U6610 ( .A(n4760), .B(key[487]), .Z(n4675) );
  XNOR U6611 ( .A(n4676), .B(n4675), .Z(n4677) );
  XNOR U6612 ( .A(\w3[2][96] ), .B(n4677), .Z(\w1[3][103] ) );
  XOR U6613 ( .A(\w3[2][105] ), .B(\w3[2][97] ), .Z(n4738) );
  XOR U6614 ( .A(n4738), .B(key[488]), .Z(n4679) );
  XOR U6615 ( .A(\w3[2][120] ), .B(\w3[2][112] ), .Z(n5070) );
  XNOR U6616 ( .A(\w3[2][96] ), .B(n5070), .Z(n4678) );
  XNOR U6617 ( .A(n4679), .B(n4678), .Z(\w1[3][104] ) );
  XOR U6618 ( .A(\w3[2][106] ), .B(\w3[2][98] ), .Z(n4742) );
  XOR U6619 ( .A(n4742), .B(key[489]), .Z(n4681) );
  XOR U6620 ( .A(\w3[2][97] ), .B(\w3[2][121] ), .Z(n5069) );
  XNOR U6621 ( .A(\w3[2][113] ), .B(n5069), .Z(n4680) );
  XNOR U6622 ( .A(n4681), .B(n4680), .Z(\w1[3][105] ) );
  XOR U6623 ( .A(\w3[2][107] ), .B(\w3[2][99] ), .Z(n4683) );
  XOR U6624 ( .A(\w3[2][98] ), .B(\w3[2][122] ), .Z(n5074) );
  XNOR U6625 ( .A(n5074), .B(key[490]), .Z(n4682) );
  XNOR U6626 ( .A(n4683), .B(n4682), .Z(n4684) );
  XOR U6627 ( .A(\w3[2][114] ), .B(n4684), .Z(\w1[3][106] ) );
  XOR U6628 ( .A(\w3[2][99] ), .B(\w3[2][123] ), .Z(n5078) );
  XNOR U6629 ( .A(\w3[2][108] ), .B(n5078), .Z(n4685) );
  XNOR U6630 ( .A(\w3[2][104] ), .B(n4685), .Z(n4711) );
  XOR U6631 ( .A(n4711), .B(key[491]), .Z(n4687) );
  XOR U6632 ( .A(\w3[2][96] ), .B(\w3[2][100] ), .Z(n5082) );
  XNOR U6633 ( .A(\w3[2][115] ), .B(n5082), .Z(n4686) );
  XNOR U6634 ( .A(n4687), .B(n4686), .Z(\w1[3][107] ) );
  XOR U6635 ( .A(\w3[2][100] ), .B(\w3[2][104] ), .Z(n4689) );
  XNOR U6636 ( .A(\w3[2][124] ), .B(\w3[2][109] ), .Z(n4688) );
  XNOR U6637 ( .A(n4689), .B(n4688), .Z(n4714) );
  XOR U6638 ( .A(n4714), .B(key[492]), .Z(n4692) );
  XNOR U6639 ( .A(\w3[2][116] ), .B(n4690), .Z(n4691) );
  XNOR U6640 ( .A(n4692), .B(n4691), .Z(\w1[3][108] ) );
  XOR U6641 ( .A(\w3[2][125] ), .B(\w3[2][101] ), .Z(n4717) );
  XOR U6642 ( .A(n4717), .B(key[493]), .Z(n4694) );
  XNOR U6643 ( .A(\w3[2][102] ), .B(\w3[2][110] ), .Z(n4693) );
  XNOR U6644 ( .A(n4694), .B(n4693), .Z(n4695) );
  XOR U6645 ( .A(\w3[2][117] ), .B(n4695), .Z(\w1[3][109] ) );
  XOR U6646 ( .A(\w3[2][11] ), .B(\w3[2][18] ), .Z(n4697) );
  XOR U6647 ( .A(\w3[2][2] ), .B(\w3[2][26] ), .Z(n4783) );
  XNOR U6648 ( .A(n4783), .B(key[394]), .Z(n4696) );
  XNOR U6649 ( .A(n4697), .B(n4696), .Z(n4698) );
  XOR U6650 ( .A(\w3[2][3] ), .B(n4698), .Z(\w1[3][10] ) );
  XNOR U6651 ( .A(\w3[2][111] ), .B(\w3[2][104] ), .Z(n4726) );
  XNOR U6652 ( .A(n4699), .B(n4726), .Z(n4721) );
  XOR U6653 ( .A(n4721), .B(key[494]), .Z(n4702) );
  XNOR U6654 ( .A(\w3[2][118] ), .B(n4700), .Z(n4701) );
  XNOR U6655 ( .A(n4702), .B(n4701), .Z(\w1[3][110] ) );
  XOR U6656 ( .A(\w3[2][127] ), .B(\w3[2][103] ), .Z(n4724) );
  XOR U6657 ( .A(n4724), .B(key[495]), .Z(n4704) );
  XOR U6658 ( .A(\w3[2][96] ), .B(\w3[2][104] ), .Z(n4731) );
  XNOR U6659 ( .A(\w3[2][119] ), .B(n4731), .Z(n4703) );
  XNOR U6660 ( .A(n4704), .B(n4703), .Z(\w1[3][111] ) );
  XOR U6661 ( .A(\w3[2][105] ), .B(\w3[2][113] ), .Z(n5073) );
  XOR U6662 ( .A(n5073), .B(key[496]), .Z(n4706) );
  XNOR U6663 ( .A(\w3[2][120] ), .B(n4731), .Z(n4705) );
  XNOR U6664 ( .A(n4706), .B(n4705), .Z(\w1[3][112] ) );
  XOR U6665 ( .A(\w3[2][106] ), .B(\w3[2][114] ), .Z(n5077) );
  XOR U6666 ( .A(n5077), .B(key[497]), .Z(n4708) );
  XNOR U6667 ( .A(\w3[2][105] ), .B(n5069), .Z(n4707) );
  XNOR U6668 ( .A(n4708), .B(n4707), .Z(\w1[3][113] ) );
  XOR U6669 ( .A(\w3[2][107] ), .B(\w3[2][115] ), .Z(n4744) );
  XOR U6670 ( .A(n4744), .B(key[498]), .Z(n4710) );
  XNOR U6671 ( .A(n4742), .B(\w3[2][122] ), .Z(n4709) );
  XNOR U6672 ( .A(n4710), .B(n4709), .Z(\w1[3][114] ) );
  XOR U6673 ( .A(\w3[2][116] ), .B(\w3[2][112] ), .Z(n4745) );
  XOR U6674 ( .A(n4745), .B(key[499]), .Z(n4713) );
  XNOR U6675 ( .A(\w3[2][107] ), .B(n4711), .Z(n4712) );
  XNOR U6676 ( .A(n4713), .B(n4712), .Z(\w1[3][115] ) );
  XOR U6677 ( .A(\w3[2][117] ), .B(\w3[2][112] ), .Z(n4748) );
  XOR U6678 ( .A(n4748), .B(key[500]), .Z(n4716) );
  XNOR U6679 ( .A(\w3[2][108] ), .B(n4714), .Z(n4715) );
  XNOR U6680 ( .A(n4716), .B(n4715), .Z(\w1[3][116] ) );
  XOR U6681 ( .A(n4717), .B(key[501]), .Z(n4720) );
  XNOR U6682 ( .A(\w3[2][109] ), .B(n4718), .Z(n4719) );
  XNOR U6683 ( .A(n4720), .B(n4719), .Z(\w1[3][117] ) );
  XOR U6684 ( .A(\w3[2][119] ), .B(\w3[2][112] ), .Z(n4756) );
  XOR U6685 ( .A(n4756), .B(key[502]), .Z(n4723) );
  XNOR U6686 ( .A(\w3[2][110] ), .B(n4721), .Z(n4722) );
  XNOR U6687 ( .A(n4723), .B(n4722), .Z(\w1[3][118] ) );
  XNOR U6688 ( .A(n4724), .B(key[503]), .Z(n4725) );
  XNOR U6689 ( .A(n4726), .B(n4725), .Z(n4727) );
  XNOR U6690 ( .A(\w3[2][112] ), .B(n4727), .Z(\w1[3][119] ) );
  XOR U6691 ( .A(\w3[2][3] ), .B(\w3[2][27] ), .Z(n4824) );
  XNOR U6692 ( .A(\w3[2][8] ), .B(\w3[2][12] ), .Z(n4728) );
  XNOR U6693 ( .A(n4824), .B(n4728), .Z(n4780) );
  XOR U6694 ( .A(n4780), .B(key[395]), .Z(n4730) );
  XOR U6695 ( .A(\w3[2][0] ), .B(\w3[2][4] ), .Z(n4854) );
  XNOR U6696 ( .A(\w3[2][19] ), .B(n4854), .Z(n4729) );
  XNOR U6697 ( .A(n4730), .B(n4729), .Z(\w1[3][11] ) );
  XOR U6698 ( .A(n4731), .B(key[504]), .Z(n4733) );
  XNOR U6699 ( .A(\w3[2][113] ), .B(\w3[2][121] ), .Z(n4732) );
  XNOR U6700 ( .A(n4733), .B(n4732), .Z(n4734) );
  XOR U6701 ( .A(\w3[2][112] ), .B(n4734), .Z(\w1[3][120] ) );
  XOR U6702 ( .A(\w3[2][122] ), .B(key[505]), .Z(n4736) );
  XNOR U6703 ( .A(\w3[2][113] ), .B(\w3[2][114] ), .Z(n4735) );
  XNOR U6704 ( .A(n4736), .B(n4735), .Z(n4737) );
  XOR U6705 ( .A(n4738), .B(n4737), .Z(\w1[3][121] ) );
  XOR U6706 ( .A(\w3[2][123] ), .B(key[506]), .Z(n4740) );
  XNOR U6707 ( .A(\w3[2][114] ), .B(\w3[2][115] ), .Z(n4739) );
  XNOR U6708 ( .A(n4740), .B(n4739), .Z(n4741) );
  XOR U6709 ( .A(n4742), .B(n4741), .Z(\w1[3][122] ) );
  XNOR U6710 ( .A(\w3[2][124] ), .B(\w3[2][120] ), .Z(n4743) );
  XNOR U6711 ( .A(n4744), .B(n4743), .Z(n5081) );
  XOR U6712 ( .A(n5081), .B(key[507]), .Z(n4747) );
  XNOR U6713 ( .A(\w3[2][99] ), .B(n4745), .Z(n4746) );
  XNOR U6714 ( .A(n4747), .B(n4746), .Z(\w1[3][123] ) );
  XOR U6715 ( .A(n4748), .B(key[508]), .Z(n4751) );
  XNOR U6716 ( .A(n4749), .B(\w3[2][100] ), .Z(n4750) );
  XNOR U6717 ( .A(n4751), .B(n4750), .Z(\w1[3][124] ) );
  XOR U6718 ( .A(\w3[2][118] ), .B(key[509]), .Z(n4754) );
  XNOR U6719 ( .A(n4752), .B(\w3[2][126] ), .Z(n4753) );
  XNOR U6720 ( .A(n4754), .B(n4753), .Z(n4755) );
  XOR U6721 ( .A(\w3[2][101] ), .B(n4755), .Z(\w1[3][125] ) );
  XOR U6722 ( .A(n4756), .B(key[510]), .Z(n4759) );
  XNOR U6723 ( .A(\w3[2][102] ), .B(n4757), .Z(n4758) );
  XNOR U6724 ( .A(n4759), .B(n4758), .Z(\w1[3][126] ) );
  XOR U6725 ( .A(n5070), .B(key[511]), .Z(n4762) );
  XNOR U6726 ( .A(\w3[2][103] ), .B(n4760), .Z(n4761) );
  XNOR U6727 ( .A(n4762), .B(n4761), .Z(\w1[3][127] ) );
  XOR U6728 ( .A(\w3[2][13] ), .B(\w3[2][28] ), .Z(n4764) );
  XNOR U6729 ( .A(\w3[2][8] ), .B(\w3[2][4] ), .Z(n4763) );
  XNOR U6730 ( .A(n4764), .B(n4763), .Z(n4786) );
  XOR U6731 ( .A(n4786), .B(key[396]), .Z(n4766) );
  XOR U6732 ( .A(\w3[2][0] ), .B(\w3[2][5] ), .Z(n4891) );
  XNOR U6733 ( .A(\w3[2][20] ), .B(n4891), .Z(n4765) );
  XNOR U6734 ( .A(n4766), .B(n4765), .Z(\w1[3][12] ) );
  XOR U6735 ( .A(\w3[2][14] ), .B(\w3[2][21] ), .Z(n4768) );
  XOR U6736 ( .A(\w3[2][5] ), .B(\w3[2][29] ), .Z(n4789) );
  XNOR U6737 ( .A(n4789), .B(key[397]), .Z(n4767) );
  XNOR U6738 ( .A(n4768), .B(n4767), .Z(n4769) );
  XOR U6739 ( .A(\w3[2][6] ), .B(n4769), .Z(\w1[3][13] ) );
  XOR U6740 ( .A(\w3[2][6] ), .B(\w3[2][30] ), .Z(n4932) );
  XNOR U6741 ( .A(\w3[2][8] ), .B(\w3[2][15] ), .Z(n4797) );
  XNOR U6742 ( .A(n4932), .B(n4797), .Z(n4792) );
  XOR U6743 ( .A(n4792), .B(key[398]), .Z(n4771) );
  XOR U6744 ( .A(\w3[2][0] ), .B(\w3[2][7] ), .Z(n4967) );
  XNOR U6745 ( .A(\w3[2][22] ), .B(n4967), .Z(n4770) );
  XNOR U6746 ( .A(n4771), .B(n4770), .Z(\w1[3][14] ) );
  XOR U6747 ( .A(\w3[2][7] ), .B(\w3[2][31] ), .Z(n4795) );
  XOR U6748 ( .A(n4795), .B(key[399]), .Z(n4773) );
  XOR U6749 ( .A(\w3[2][8] ), .B(\w3[2][0] ), .Z(n4799) );
  XNOR U6750 ( .A(\w3[2][23] ), .B(n4799), .Z(n4772) );
  XNOR U6751 ( .A(n4773), .B(n4772), .Z(\w1[3][15] ) );
  XOR U6752 ( .A(\w3[2][17] ), .B(\w3[2][9] ), .Z(n4803) );
  XOR U6753 ( .A(n4803), .B(key[400]), .Z(n4775) );
  XNOR U6754 ( .A(\w3[2][24] ), .B(n4799), .Z(n4774) );
  XNOR U6755 ( .A(n4775), .B(n4774), .Z(\w1[3][16] ) );
  XOR U6756 ( .A(\w3[2][18] ), .B(\w3[2][10] ), .Z(n4823) );
  XOR U6757 ( .A(n4823), .B(key[401]), .Z(n4777) );
  XNOR U6758 ( .A(n5088), .B(\w3[2][9] ), .Z(n4776) );
  XNOR U6759 ( .A(n4777), .B(n4776), .Z(\w1[3][17] ) );
  XOR U6760 ( .A(\w3[2][11] ), .B(\w3[2][19] ), .Z(n4811) );
  XOR U6761 ( .A(n4811), .B(key[402]), .Z(n4779) );
  XNOR U6762 ( .A(n4783), .B(\w3[2][10] ), .Z(n4778) );
  XNOR U6763 ( .A(n4779), .B(n4778), .Z(\w1[3][18] ) );
  XOR U6764 ( .A(\w3[2][16] ), .B(\w3[2][20] ), .Z(n4812) );
  XOR U6765 ( .A(n4812), .B(key[403]), .Z(n4782) );
  XNOR U6766 ( .A(\w3[2][11] ), .B(n4780), .Z(n4781) );
  XNOR U6767 ( .A(n4782), .B(n4781), .Z(\w1[3][19] ) );
  XOR U6768 ( .A(n4803), .B(key[385]), .Z(n4785) );
  XNOR U6769 ( .A(\w3[2][25] ), .B(n4783), .Z(n4784) );
  XNOR U6770 ( .A(n4785), .B(n4784), .Z(\w1[3][1] ) );
  XOR U6771 ( .A(\w3[2][16] ), .B(\w3[2][21] ), .Z(n4817) );
  XOR U6772 ( .A(n4817), .B(key[404]), .Z(n4788) );
  XNOR U6773 ( .A(\w3[2][12] ), .B(n4786), .Z(n4787) );
  XNOR U6774 ( .A(n4788), .B(n4787), .Z(\w1[3][20] ) );
  XOR U6775 ( .A(\w3[2][14] ), .B(\w3[2][22] ), .Z(n4827) );
  XOR U6776 ( .A(n4827), .B(key[405]), .Z(n4791) );
  XNOR U6777 ( .A(\w3[2][13] ), .B(n4789), .Z(n4790) );
  XNOR U6778 ( .A(n4791), .B(n4790), .Z(\w1[3][21] ) );
  XOR U6779 ( .A(\w3[2][16] ), .B(\w3[2][23] ), .Z(n4828) );
  XOR U6780 ( .A(n4828), .B(key[406]), .Z(n4794) );
  XNOR U6781 ( .A(\w3[2][14] ), .B(n4792), .Z(n4793) );
  XNOR U6782 ( .A(n4794), .B(n4793), .Z(\w1[3][22] ) );
  XNOR U6783 ( .A(n4795), .B(key[407]), .Z(n4796) );
  XNOR U6784 ( .A(n4797), .B(n4796), .Z(n4798) );
  XNOR U6785 ( .A(\w3[2][16] ), .B(n4798), .Z(\w1[3][23] ) );
  XOR U6786 ( .A(\w3[2][17] ), .B(key[408]), .Z(n4801) );
  XNOR U6787 ( .A(\w3[2][25] ), .B(n4799), .Z(n4800) );
  XNOR U6788 ( .A(n4801), .B(n4800), .Z(n4802) );
  XOR U6789 ( .A(\w3[2][16] ), .B(n4802), .Z(\w1[3][24] ) );
  XOR U6790 ( .A(n4803), .B(key[409]), .Z(n4805) );
  XNOR U6791 ( .A(\w3[2][1] ), .B(\w3[2][26] ), .Z(n4804) );
  XNOR U6792 ( .A(n4805), .B(n4804), .Z(n4806) );
  XOR U6793 ( .A(\w3[2][18] ), .B(n4806), .Z(\w1[3][25] ) );
  XOR U6794 ( .A(n4823), .B(key[410]), .Z(n4808) );
  XNOR U6795 ( .A(\w3[2][2] ), .B(\w3[2][19] ), .Z(n4807) );
  XNOR U6796 ( .A(n4808), .B(n4807), .Z(n4809) );
  XOR U6797 ( .A(\w3[2][27] ), .B(n4809), .Z(\w1[3][26] ) );
  XNOR U6798 ( .A(\w3[2][24] ), .B(\w3[2][28] ), .Z(n4810) );
  XNOR U6799 ( .A(n4811), .B(n4810), .Z(n4853) );
  XOR U6800 ( .A(n4853), .B(key[411]), .Z(n4814) );
  XNOR U6801 ( .A(\w3[2][3] ), .B(n4812), .Z(n4813) );
  XNOR U6802 ( .A(n4814), .B(n4813), .Z(\w1[3][27] ) );
  XOR U6803 ( .A(\w3[2][20] ), .B(\w3[2][29] ), .Z(n4816) );
  XNOR U6804 ( .A(\w3[2][24] ), .B(\w3[2][12] ), .Z(n4815) );
  XNOR U6805 ( .A(n4816), .B(n4815), .Z(n4890) );
  XOR U6806 ( .A(n4890), .B(key[412]), .Z(n4819) );
  XNOR U6807 ( .A(\w3[2][4] ), .B(n4817), .Z(n4818) );
  XNOR U6808 ( .A(n4819), .B(n4818), .Z(\w1[3][28] ) );
  XOR U6809 ( .A(\w3[2][13] ), .B(\w3[2][21] ), .Z(n4931) );
  XOR U6810 ( .A(n4931), .B(key[413]), .Z(n4821) );
  XNOR U6811 ( .A(\w3[2][22] ), .B(\w3[2][30] ), .Z(n4820) );
  XNOR U6812 ( .A(n4821), .B(n4820), .Z(n4822) );
  XOR U6813 ( .A(\w3[2][5] ), .B(n4822), .Z(\w1[3][29] ) );
  XOR U6814 ( .A(n4823), .B(key[386]), .Z(n4826) );
  XNOR U6815 ( .A(\w3[2][26] ), .B(n4824), .Z(n4825) );
  XNOR U6816 ( .A(n4826), .B(n4825), .Z(\w1[3][2] ) );
  XNOR U6817 ( .A(\w3[2][24] ), .B(\w3[2][31] ), .Z(n5005) );
  XNOR U6818 ( .A(n4827), .B(n5005), .Z(n4966) );
  XOR U6819 ( .A(n4966), .B(key[414]), .Z(n4830) );
  XNOR U6820 ( .A(\w3[2][6] ), .B(n4828), .Z(n4829) );
  XNOR U6821 ( .A(n4830), .B(n4829), .Z(\w1[3][30] ) );
  XOR U6822 ( .A(\w3[2][15] ), .B(\w3[2][23] ), .Z(n5003) );
  XOR U6823 ( .A(n5003), .B(key[415]), .Z(n4832) );
  XNOR U6824 ( .A(n5044), .B(\w3[2][7] ), .Z(n4831) );
  XNOR U6825 ( .A(n4832), .B(n4831), .Z(\w1[3][31] ) );
  XOR U6826 ( .A(\w3[2][33] ), .B(\w3[2][57] ), .Z(n4887) );
  XOR U6827 ( .A(n4887), .B(key[416]), .Z(n4834) );
  XOR U6828 ( .A(\w3[2][48] ), .B(\w3[2][56] ), .Z(n4948) );
  XNOR U6829 ( .A(n4948), .B(\w3[2][40] ), .Z(n4833) );
  XNOR U6830 ( .A(n4834), .B(n4833), .Z(\w1[3][32] ) );
  XOR U6831 ( .A(\w3[2][34] ), .B(\w3[2][58] ), .Z(n4895) );
  XOR U6832 ( .A(n4895), .B(key[417]), .Z(n4836) );
  XOR U6833 ( .A(\w3[2][41] ), .B(\w3[2][49] ), .Z(n4919) );
  XNOR U6834 ( .A(\w3[2][57] ), .B(n4919), .Z(n4835) );
  XNOR U6835 ( .A(n4836), .B(n4835), .Z(\w1[3][33] ) );
  XOR U6836 ( .A(\w3[2][35] ), .B(\w3[2][59] ), .Z(n4866) );
  XOR U6837 ( .A(n4866), .B(key[418]), .Z(n4838) );
  XOR U6838 ( .A(\w3[2][42] ), .B(\w3[2][50] ), .Z(n4923) );
  XNOR U6839 ( .A(\w3[2][58] ), .B(n4923), .Z(n4837) );
  XNOR U6840 ( .A(n4838), .B(n4837), .Z(\w1[3][34] ) );
  XOR U6841 ( .A(\w3[2][36] ), .B(\w3[2][32] ), .Z(n4868) );
  XOR U6842 ( .A(n4868), .B(key[419]), .Z(n4841) );
  XOR U6843 ( .A(\w3[2][43] ), .B(\w3[2][51] ), .Z(n4894) );
  XNOR U6844 ( .A(\w3[2][56] ), .B(n4894), .Z(n4839) );
  XNOR U6845 ( .A(\w3[2][60] ), .B(n4839), .Z(n4928) );
  XNOR U6846 ( .A(\w3[2][59] ), .B(n4928), .Z(n4840) );
  XNOR U6847 ( .A(n4841), .B(n4840), .Z(\w1[3][35] ) );
  XOR U6848 ( .A(\w3[2][32] ), .B(\w3[2][37] ), .Z(n4873) );
  XOR U6849 ( .A(n4873), .B(key[420]), .Z(n4845) );
  XOR U6850 ( .A(\w3[2][52] ), .B(\w3[2][61] ), .Z(n4843) );
  XNOR U6851 ( .A(\w3[2][56] ), .B(\w3[2][44] ), .Z(n4842) );
  XNOR U6852 ( .A(n4843), .B(n4842), .Z(n4936) );
  XNOR U6853 ( .A(\w3[2][60] ), .B(n4936), .Z(n4844) );
  XNOR U6854 ( .A(n4845), .B(n4844), .Z(\w1[3][36] ) );
  XOR U6855 ( .A(\w3[2][38] ), .B(\w3[2][62] ), .Z(n4879) );
  XOR U6856 ( .A(n4879), .B(key[421]), .Z(n4847) );
  XOR U6857 ( .A(\w3[2][45] ), .B(\w3[2][53] ), .Z(n4939) );
  XNOR U6858 ( .A(\w3[2][61] ), .B(n4939), .Z(n4846) );
  XNOR U6859 ( .A(n4847), .B(n4846), .Z(\w1[3][37] ) );
  XOR U6860 ( .A(\w3[2][32] ), .B(\w3[2][39] ), .Z(n4880) );
  XOR U6861 ( .A(n4880), .B(key[422]), .Z(n4849) );
  XOR U6862 ( .A(\w3[2][46] ), .B(\w3[2][54] ), .Z(n4905) );
  XNOR U6863 ( .A(\w3[2][56] ), .B(\w3[2][63] ), .Z(n4851) );
  XNOR U6864 ( .A(n4905), .B(n4851), .Z(n4944) );
  XNOR U6865 ( .A(\w3[2][62] ), .B(n4944), .Z(n4848) );
  XNOR U6866 ( .A(n4849), .B(n4848), .Z(\w1[3][38] ) );
  XOR U6867 ( .A(\w3[2][47] ), .B(\w3[2][55] ), .Z(n4947) );
  XNOR U6868 ( .A(n4947), .B(key[423]), .Z(n4850) );
  XNOR U6869 ( .A(n4851), .B(n4850), .Z(n4852) );
  XNOR U6870 ( .A(\w3[2][32] ), .B(n4852), .Z(\w1[3][39] ) );
  XOR U6871 ( .A(n4853), .B(key[387]), .Z(n4856) );
  XNOR U6872 ( .A(n4854), .B(\w3[2][27] ), .Z(n4855) );
  XNOR U6873 ( .A(n4856), .B(n4855), .Z(\w1[3][3] ) );
  XOR U6874 ( .A(\w3[2][32] ), .B(key[424]), .Z(n4858) );
  XNOR U6875 ( .A(\w3[2][33] ), .B(\w3[2][41] ), .Z(n4857) );
  XNOR U6876 ( .A(n4858), .B(n4857), .Z(n4859) );
  XOR U6877 ( .A(n4948), .B(n4859), .Z(\w1[3][40] ) );
  XOR U6878 ( .A(\w3[2][42] ), .B(key[425]), .Z(n4861) );
  XNOR U6879 ( .A(\w3[2][49] ), .B(\w3[2][34] ), .Z(n4860) );
  XNOR U6880 ( .A(n4861), .B(n4860), .Z(n4862) );
  XOR U6881 ( .A(n4887), .B(n4862), .Z(\w1[3][41] ) );
  XOR U6882 ( .A(\w3[2][43] ), .B(key[426]), .Z(n4864) );
  XNOR U6883 ( .A(\w3[2][50] ), .B(\w3[2][35] ), .Z(n4863) );
  XNOR U6884 ( .A(n4864), .B(n4863), .Z(n4865) );
  XOR U6885 ( .A(n4895), .B(n4865), .Z(\w1[3][42] ) );
  XNOR U6886 ( .A(\w3[2][40] ), .B(n4866), .Z(n4867) );
  XNOR U6887 ( .A(\w3[2][44] ), .B(n4867), .Z(n4898) );
  XOR U6888 ( .A(n4898), .B(key[427]), .Z(n4870) );
  XNOR U6889 ( .A(\w3[2][51] ), .B(n4868), .Z(n4869) );
  XNOR U6890 ( .A(n4870), .B(n4869), .Z(\w1[3][43] ) );
  XOR U6891 ( .A(\w3[2][36] ), .B(\w3[2][45] ), .Z(n4872) );
  XNOR U6892 ( .A(\w3[2][40] ), .B(\w3[2][60] ), .Z(n4871) );
  XNOR U6893 ( .A(n4872), .B(n4871), .Z(n4901) );
  XOR U6894 ( .A(n4901), .B(key[428]), .Z(n4875) );
  XNOR U6895 ( .A(\w3[2][52] ), .B(n4873), .Z(n4874) );
  XNOR U6896 ( .A(n4875), .B(n4874), .Z(\w1[3][44] ) );
  XOR U6897 ( .A(\w3[2][61] ), .B(\w3[2][37] ), .Z(n4904) );
  XOR U6898 ( .A(n4904), .B(key[429]), .Z(n4877) );
  XNOR U6899 ( .A(\w3[2][38] ), .B(\w3[2][46] ), .Z(n4876) );
  XNOR U6900 ( .A(n4877), .B(n4876), .Z(n4878) );
  XOR U6901 ( .A(\w3[2][53] ), .B(n4878), .Z(\w1[3][45] ) );
  XNOR U6902 ( .A(\w3[2][40] ), .B(\w3[2][47] ), .Z(n4913) );
  XNOR U6903 ( .A(n4879), .B(n4913), .Z(n4908) );
  XOR U6904 ( .A(n4908), .B(key[430]), .Z(n4882) );
  XNOR U6905 ( .A(\w3[2][54] ), .B(n4880), .Z(n4881) );
  XNOR U6906 ( .A(n4882), .B(n4881), .Z(\w1[3][46] ) );
  XOR U6907 ( .A(\w3[2][63] ), .B(\w3[2][39] ), .Z(n4911) );
  XOR U6908 ( .A(n4911), .B(key[431]), .Z(n4884) );
  XOR U6909 ( .A(\w3[2][40] ), .B(\w3[2][32] ), .Z(n4915) );
  XNOR U6910 ( .A(\w3[2][55] ), .B(n4915), .Z(n4883) );
  XNOR U6911 ( .A(n4884), .B(n4883), .Z(\w1[3][47] ) );
  XOR U6912 ( .A(n4915), .B(key[432]), .Z(n4886) );
  XNOR U6913 ( .A(\w3[2][56] ), .B(n4919), .Z(n4885) );
  XNOR U6914 ( .A(n4886), .B(n4885), .Z(\w1[3][48] ) );
  XOR U6915 ( .A(n4923), .B(key[433]), .Z(n4889) );
  XNOR U6916 ( .A(n4887), .B(\w3[2][41] ), .Z(n4888) );
  XNOR U6917 ( .A(n4889), .B(n4888), .Z(\w1[3][49] ) );
  XOR U6918 ( .A(n4890), .B(key[388]), .Z(n4893) );
  XNOR U6919 ( .A(n4891), .B(\w3[2][28] ), .Z(n4892) );
  XNOR U6920 ( .A(n4893), .B(n4892), .Z(\w1[3][4] ) );
  XOR U6921 ( .A(n4894), .B(key[434]), .Z(n4897) );
  XNOR U6922 ( .A(n4895), .B(\w3[2][42] ), .Z(n4896) );
  XNOR U6923 ( .A(n4897), .B(n4896), .Z(\w1[3][50] ) );
  XOR U6924 ( .A(\w3[2][48] ), .B(\w3[2][52] ), .Z(n4927) );
  XOR U6925 ( .A(n4927), .B(key[435]), .Z(n4900) );
  XNOR U6926 ( .A(\w3[2][43] ), .B(n4898), .Z(n4899) );
  XNOR U6927 ( .A(n4900), .B(n4899), .Z(\w1[3][51] ) );
  XOR U6928 ( .A(\w3[2][48] ), .B(\w3[2][53] ), .Z(n4935) );
  XOR U6929 ( .A(n4935), .B(key[436]), .Z(n4903) );
  XNOR U6930 ( .A(\w3[2][44] ), .B(n4901), .Z(n4902) );
  XNOR U6931 ( .A(n4903), .B(n4902), .Z(\w1[3][52] ) );
  XOR U6932 ( .A(n4904), .B(key[437]), .Z(n4907) );
  XNOR U6933 ( .A(\w3[2][45] ), .B(n4905), .Z(n4906) );
  XNOR U6934 ( .A(n4907), .B(n4906), .Z(\w1[3][53] ) );
  XOR U6935 ( .A(\w3[2][48] ), .B(\w3[2][55] ), .Z(n4943) );
  XOR U6936 ( .A(n4943), .B(key[438]), .Z(n4910) );
  XNOR U6937 ( .A(\w3[2][46] ), .B(n4908), .Z(n4909) );
  XNOR U6938 ( .A(n4910), .B(n4909), .Z(\w1[3][54] ) );
  XNOR U6939 ( .A(n4911), .B(key[439]), .Z(n4912) );
  XNOR U6940 ( .A(n4913), .B(n4912), .Z(n4914) );
  XNOR U6941 ( .A(\w3[2][48] ), .B(n4914), .Z(\w1[3][55] ) );
  XOR U6942 ( .A(n4915), .B(key[440]), .Z(n4917) );
  XNOR U6943 ( .A(\w3[2][48] ), .B(\w3[2][49] ), .Z(n4916) );
  XNOR U6944 ( .A(n4917), .B(n4916), .Z(n4918) );
  XOR U6945 ( .A(\w3[2][57] ), .B(n4918), .Z(\w1[3][56] ) );
  XOR U6946 ( .A(\w3[2][50] ), .B(key[441]), .Z(n4921) );
  XNOR U6947 ( .A(n4919), .B(\w3[2][58] ), .Z(n4920) );
  XNOR U6948 ( .A(n4921), .B(n4920), .Z(n4922) );
  XOR U6949 ( .A(\w3[2][33] ), .B(n4922), .Z(\w1[3][57] ) );
  XOR U6950 ( .A(\w3[2][51] ), .B(key[442]), .Z(n4925) );
  XNOR U6951 ( .A(n4923), .B(\w3[2][59] ), .Z(n4924) );
  XNOR U6952 ( .A(n4925), .B(n4924), .Z(n4926) );
  XOR U6953 ( .A(\w3[2][34] ), .B(n4926), .Z(\w1[3][58] ) );
  XOR U6954 ( .A(n4927), .B(key[443]), .Z(n4930) );
  XNOR U6955 ( .A(\w3[2][35] ), .B(n4928), .Z(n4929) );
  XNOR U6956 ( .A(n4930), .B(n4929), .Z(\w1[3][59] ) );
  XOR U6957 ( .A(n4931), .B(key[389]), .Z(n4934) );
  XNOR U6958 ( .A(\w3[2][29] ), .B(n4932), .Z(n4933) );
  XNOR U6959 ( .A(n4934), .B(n4933), .Z(\w1[3][5] ) );
  XOR U6960 ( .A(n4935), .B(key[444]), .Z(n4938) );
  XNOR U6961 ( .A(\w3[2][36] ), .B(n4936), .Z(n4937) );
  XNOR U6962 ( .A(n4938), .B(n4937), .Z(\w1[3][60] ) );
  XOR U6963 ( .A(\w3[2][54] ), .B(key[445]), .Z(n4941) );
  XNOR U6964 ( .A(n4939), .B(\w3[2][62] ), .Z(n4940) );
  XNOR U6965 ( .A(n4941), .B(n4940), .Z(n4942) );
  XOR U6966 ( .A(\w3[2][37] ), .B(n4942), .Z(\w1[3][61] ) );
  XOR U6967 ( .A(n4943), .B(key[446]), .Z(n4946) );
  XNOR U6968 ( .A(\w3[2][38] ), .B(n4944), .Z(n4945) );
  XNOR U6969 ( .A(n4946), .B(n4945), .Z(\w1[3][62] ) );
  XOR U6970 ( .A(n4947), .B(key[447]), .Z(n4950) );
  XNOR U6971 ( .A(n4948), .B(\w3[2][39] ), .Z(n4949) );
  XNOR U6972 ( .A(n4950), .B(n4949), .Z(\w1[3][63] ) );
  XOR U6973 ( .A(\w3[2][65] ), .B(\w3[2][89] ), .Z(n5009) );
  XOR U6974 ( .A(n5009), .B(key[448]), .Z(n4952) );
  XOR U6975 ( .A(\w3[2][80] ), .B(\w3[2][88] ), .Z(n5066) );
  XNOR U6976 ( .A(n5066), .B(\w3[2][72] ), .Z(n4951) );
  XNOR U6977 ( .A(n4952), .B(n4951), .Z(\w1[3][64] ) );
  XOR U6978 ( .A(\w3[2][66] ), .B(\w3[2][90] ), .Z(n5013) );
  XOR U6979 ( .A(n5013), .B(key[449]), .Z(n4954) );
  XOR U6980 ( .A(\w3[2][73] ), .B(\w3[2][81] ), .Z(n5037) );
  XNOR U6981 ( .A(\w3[2][89] ), .B(n5037), .Z(n4953) );
  XNOR U6982 ( .A(n4954), .B(n4953), .Z(\w1[3][65] ) );
  XOR U6983 ( .A(\w3[2][67] ), .B(\w3[2][91] ), .Z(n4984) );
  XOR U6984 ( .A(n4984), .B(key[450]), .Z(n4956) );
  XOR U6985 ( .A(\w3[2][74] ), .B(\w3[2][82] ), .Z(n5045) );
  XNOR U6986 ( .A(\w3[2][90] ), .B(n5045), .Z(n4955) );
  XNOR U6987 ( .A(n4956), .B(n4955), .Z(\w1[3][66] ) );
  XOR U6988 ( .A(\w3[2][68] ), .B(\w3[2][64] ), .Z(n4986) );
  XOR U6989 ( .A(n4986), .B(key[451]), .Z(n4959) );
  XOR U6990 ( .A(\w3[2][75] ), .B(\w3[2][83] ), .Z(n5012) );
  XNOR U6991 ( .A(\w3[2][88] ), .B(n5012), .Z(n4957) );
  XNOR U6992 ( .A(\w3[2][92] ), .B(n4957), .Z(n5050) );
  XNOR U6993 ( .A(\w3[2][91] ), .B(n5050), .Z(n4958) );
  XNOR U6994 ( .A(n4959), .B(n4958), .Z(\w1[3][67] ) );
  XOR U6995 ( .A(\w3[2][64] ), .B(\w3[2][69] ), .Z(n4991) );
  XOR U6996 ( .A(n4991), .B(key[452]), .Z(n4963) );
  XOR U6997 ( .A(\w3[2][84] ), .B(\w3[2][93] ), .Z(n4961) );
  XNOR U6998 ( .A(\w3[2][88] ), .B(\w3[2][76] ), .Z(n4960) );
  XNOR U6999 ( .A(n4961), .B(n4960), .Z(n5054) );
  XNOR U7000 ( .A(\w3[2][92] ), .B(n5054), .Z(n4962) );
  XNOR U7001 ( .A(n4963), .B(n4962), .Z(\w1[3][68] ) );
  XOR U7002 ( .A(\w3[2][70] ), .B(\w3[2][94] ), .Z(n4997) );
  XOR U7003 ( .A(n4997), .B(key[453]), .Z(n4965) );
  XOR U7004 ( .A(\w3[2][77] ), .B(\w3[2][85] ), .Z(n5057) );
  XNOR U7005 ( .A(\w3[2][93] ), .B(n5057), .Z(n4964) );
  XNOR U7006 ( .A(n4965), .B(n4964), .Z(\w1[3][69] ) );
  XOR U7007 ( .A(n4966), .B(key[390]), .Z(n4969) );
  XNOR U7008 ( .A(n4967), .B(\w3[2][30] ), .Z(n4968) );
  XNOR U7009 ( .A(n4969), .B(n4968), .Z(\w1[3][6] ) );
  XOR U7010 ( .A(\w3[2][64] ), .B(\w3[2][71] ), .Z(n4998) );
  XOR U7011 ( .A(n4998), .B(key[454]), .Z(n4971) );
  XOR U7012 ( .A(\w3[2][78] ), .B(\w3[2][86] ), .Z(n5023) );
  XNOR U7013 ( .A(\w3[2][88] ), .B(\w3[2][95] ), .Z(n4973) );
  XNOR U7014 ( .A(n5023), .B(n4973), .Z(n5062) );
  XNOR U7015 ( .A(\w3[2][94] ), .B(n5062), .Z(n4970) );
  XNOR U7016 ( .A(n4971), .B(n4970), .Z(\w1[3][70] ) );
  XOR U7017 ( .A(\w3[2][79] ), .B(\w3[2][87] ), .Z(n5065) );
  XNOR U7018 ( .A(n5065), .B(key[455]), .Z(n4972) );
  XNOR U7019 ( .A(n4973), .B(n4972), .Z(n4974) );
  XNOR U7020 ( .A(\w3[2][64] ), .B(n4974), .Z(\w1[3][71] ) );
  XOR U7021 ( .A(\w3[2][64] ), .B(key[456]), .Z(n4976) );
  XNOR U7022 ( .A(\w3[2][65] ), .B(\w3[2][73] ), .Z(n4975) );
  XNOR U7023 ( .A(n4976), .B(n4975), .Z(n4977) );
  XOR U7024 ( .A(n5066), .B(n4977), .Z(\w1[3][72] ) );
  XOR U7025 ( .A(\w3[2][74] ), .B(key[457]), .Z(n4979) );
  XNOR U7026 ( .A(\w3[2][81] ), .B(\w3[2][66] ), .Z(n4978) );
  XNOR U7027 ( .A(n4979), .B(n4978), .Z(n4980) );
  XOR U7028 ( .A(n5009), .B(n4980), .Z(\w1[3][73] ) );
  XOR U7029 ( .A(\w3[2][75] ), .B(key[458]), .Z(n4982) );
  XNOR U7030 ( .A(\w3[2][82] ), .B(\w3[2][67] ), .Z(n4981) );
  XNOR U7031 ( .A(n4982), .B(n4981), .Z(n4983) );
  XOR U7032 ( .A(n5013), .B(n4983), .Z(\w1[3][74] ) );
  XNOR U7033 ( .A(\w3[2][72] ), .B(n4984), .Z(n4985) );
  XNOR U7034 ( .A(\w3[2][76] ), .B(n4985), .Z(n5016) );
  XOR U7035 ( .A(n5016), .B(key[459]), .Z(n4988) );
  XNOR U7036 ( .A(\w3[2][83] ), .B(n4986), .Z(n4987) );
  XNOR U7037 ( .A(n4988), .B(n4987), .Z(\w1[3][75] ) );
  XOR U7038 ( .A(\w3[2][68] ), .B(\w3[2][77] ), .Z(n4990) );
  XNOR U7039 ( .A(\w3[2][72] ), .B(\w3[2][92] ), .Z(n4989) );
  XNOR U7040 ( .A(n4990), .B(n4989), .Z(n5019) );
  XOR U7041 ( .A(n5019), .B(key[460]), .Z(n4993) );
  XNOR U7042 ( .A(\w3[2][84] ), .B(n4991), .Z(n4992) );
  XNOR U7043 ( .A(n4993), .B(n4992), .Z(\w1[3][76] ) );
  XOR U7044 ( .A(\w3[2][93] ), .B(\w3[2][69] ), .Z(n5022) );
  XOR U7045 ( .A(n5022), .B(key[461]), .Z(n4995) );
  XNOR U7046 ( .A(\w3[2][70] ), .B(\w3[2][78] ), .Z(n4994) );
  XNOR U7047 ( .A(n4995), .B(n4994), .Z(n4996) );
  XOR U7048 ( .A(\w3[2][85] ), .B(n4996), .Z(\w1[3][77] ) );
  XNOR U7049 ( .A(\w3[2][72] ), .B(\w3[2][79] ), .Z(n5031) );
  XNOR U7050 ( .A(n4997), .B(n5031), .Z(n5026) );
  XOR U7051 ( .A(n5026), .B(key[462]), .Z(n5000) );
  XNOR U7052 ( .A(\w3[2][86] ), .B(n4998), .Z(n4999) );
  XNOR U7053 ( .A(n5000), .B(n4999), .Z(\w1[3][78] ) );
  XOR U7054 ( .A(\w3[2][95] ), .B(\w3[2][71] ), .Z(n5029) );
  XOR U7055 ( .A(n5029), .B(key[463]), .Z(n5002) );
  XOR U7056 ( .A(\w3[2][72] ), .B(\w3[2][64] ), .Z(n5033) );
  XNOR U7057 ( .A(\w3[2][87] ), .B(n5033), .Z(n5001) );
  XNOR U7058 ( .A(n5002), .B(n5001), .Z(\w1[3][79] ) );
  XNOR U7059 ( .A(n5003), .B(key[391]), .Z(n5004) );
  XNOR U7060 ( .A(n5005), .B(n5004), .Z(n5006) );
  XNOR U7061 ( .A(\w3[2][0] ), .B(n5006), .Z(\w1[3][7] ) );
  XOR U7062 ( .A(n5033), .B(key[464]), .Z(n5008) );
  XNOR U7063 ( .A(\w3[2][88] ), .B(n5037), .Z(n5007) );
  XNOR U7064 ( .A(n5008), .B(n5007), .Z(\w1[3][80] ) );
  XOR U7065 ( .A(n5045), .B(key[465]), .Z(n5011) );
  XNOR U7066 ( .A(n5009), .B(\w3[2][73] ), .Z(n5010) );
  XNOR U7067 ( .A(n5011), .B(n5010), .Z(\w1[3][81] ) );
  XOR U7068 ( .A(n5012), .B(key[466]), .Z(n5015) );
  XNOR U7069 ( .A(n5013), .B(\w3[2][74] ), .Z(n5014) );
  XNOR U7070 ( .A(n5015), .B(n5014), .Z(\w1[3][82] ) );
  XOR U7071 ( .A(\w3[2][80] ), .B(\w3[2][84] ), .Z(n5049) );
  XOR U7072 ( .A(n5049), .B(key[467]), .Z(n5018) );
  XNOR U7073 ( .A(\w3[2][75] ), .B(n5016), .Z(n5017) );
  XNOR U7074 ( .A(n5018), .B(n5017), .Z(\w1[3][83] ) );
  XOR U7075 ( .A(\w3[2][80] ), .B(\w3[2][85] ), .Z(n5053) );
  XOR U7076 ( .A(n5053), .B(key[468]), .Z(n5021) );
  XNOR U7077 ( .A(\w3[2][76] ), .B(n5019), .Z(n5020) );
  XNOR U7078 ( .A(n5021), .B(n5020), .Z(\w1[3][84] ) );
  XOR U7079 ( .A(n5022), .B(key[469]), .Z(n5025) );
  XNOR U7080 ( .A(\w3[2][77] ), .B(n5023), .Z(n5024) );
  XNOR U7081 ( .A(n5025), .B(n5024), .Z(\w1[3][85] ) );
  XOR U7082 ( .A(\w3[2][80] ), .B(\w3[2][87] ), .Z(n5061) );
  XOR U7083 ( .A(n5061), .B(key[470]), .Z(n5028) );
  XNOR U7084 ( .A(\w3[2][78] ), .B(n5026), .Z(n5027) );
  XNOR U7085 ( .A(n5028), .B(n5027), .Z(\w1[3][86] ) );
  XNOR U7086 ( .A(n5029), .B(key[471]), .Z(n5030) );
  XNOR U7087 ( .A(n5031), .B(n5030), .Z(n5032) );
  XNOR U7088 ( .A(\w3[2][80] ), .B(n5032), .Z(\w1[3][87] ) );
  XOR U7089 ( .A(n5033), .B(key[472]), .Z(n5035) );
  XNOR U7090 ( .A(\w3[2][80] ), .B(\w3[2][81] ), .Z(n5034) );
  XNOR U7091 ( .A(n5035), .B(n5034), .Z(n5036) );
  XOR U7092 ( .A(\w3[2][89] ), .B(n5036), .Z(\w1[3][88] ) );
  XOR U7093 ( .A(\w3[2][82] ), .B(key[473]), .Z(n5039) );
  XNOR U7094 ( .A(n5037), .B(\w3[2][90] ), .Z(n5038) );
  XNOR U7095 ( .A(n5039), .B(n5038), .Z(n5040) );
  XOR U7096 ( .A(\w3[2][65] ), .B(n5040), .Z(\w1[3][89] ) );
  XOR U7097 ( .A(\w3[2][9] ), .B(key[392]), .Z(n5042) );
  XNOR U7098 ( .A(\w3[2][1] ), .B(\w3[2][0] ), .Z(n5041) );
  XNOR U7099 ( .A(n5042), .B(n5041), .Z(n5043) );
  XOR U7100 ( .A(n5044), .B(n5043), .Z(\w1[3][8] ) );
  XOR U7101 ( .A(\w3[2][83] ), .B(key[474]), .Z(n5047) );
  XNOR U7102 ( .A(n5045), .B(\w3[2][91] ), .Z(n5046) );
  XNOR U7103 ( .A(n5047), .B(n5046), .Z(n5048) );
  XOR U7104 ( .A(\w3[2][66] ), .B(n5048), .Z(\w1[3][90] ) );
  XOR U7105 ( .A(n5049), .B(key[475]), .Z(n5052) );
  XNOR U7106 ( .A(\w3[2][67] ), .B(n5050), .Z(n5051) );
  XNOR U7107 ( .A(n5052), .B(n5051), .Z(\w1[3][91] ) );
  XOR U7108 ( .A(n5053), .B(key[476]), .Z(n5056) );
  XNOR U7109 ( .A(\w3[2][68] ), .B(n5054), .Z(n5055) );
  XNOR U7110 ( .A(n5056), .B(n5055), .Z(\w1[3][92] ) );
  XOR U7111 ( .A(\w3[2][86] ), .B(key[477]), .Z(n5059) );
  XNOR U7112 ( .A(n5057), .B(\w3[2][94] ), .Z(n5058) );
  XNOR U7113 ( .A(n5059), .B(n5058), .Z(n5060) );
  XOR U7114 ( .A(\w3[2][69] ), .B(n5060), .Z(\w1[3][93] ) );
  XOR U7115 ( .A(n5061), .B(key[478]), .Z(n5064) );
  XNOR U7116 ( .A(\w3[2][70] ), .B(n5062), .Z(n5063) );
  XNOR U7117 ( .A(n5064), .B(n5063), .Z(\w1[3][94] ) );
  XOR U7118 ( .A(n5065), .B(key[479]), .Z(n5068) );
  XNOR U7119 ( .A(n5066), .B(\w3[2][71] ), .Z(n5067) );
  XNOR U7120 ( .A(n5068), .B(n5067), .Z(\w1[3][95] ) );
  XOR U7121 ( .A(\w3[2][104] ), .B(key[480]), .Z(n5072) );
  XNOR U7122 ( .A(n5070), .B(n5069), .Z(n5071) );
  XNOR U7123 ( .A(n5072), .B(n5071), .Z(\w1[3][96] ) );
  XOR U7124 ( .A(n5073), .B(key[481]), .Z(n5076) );
  XNOR U7125 ( .A(\w3[2][121] ), .B(n5074), .Z(n5075) );
  XNOR U7126 ( .A(n5076), .B(n5075), .Z(\w1[3][97] ) );
  XOR U7127 ( .A(n5077), .B(key[482]), .Z(n5080) );
  XNOR U7128 ( .A(\w3[2][122] ), .B(n5078), .Z(n5079) );
  XNOR U7129 ( .A(n5080), .B(n5079), .Z(\w1[3][98] ) );
  XOR U7130 ( .A(n5081), .B(key[483]), .Z(n5084) );
  XNOR U7131 ( .A(n5082), .B(\w3[2][123] ), .Z(n5083) );
  XNOR U7132 ( .A(n5084), .B(n5083), .Z(\w1[3][99] ) );
  XOR U7133 ( .A(\w3[2][10] ), .B(key[393]), .Z(n5086) );
  XNOR U7134 ( .A(\w3[2][2] ), .B(\w3[2][17] ), .Z(n5085) );
  XNOR U7135 ( .A(n5086), .B(n5085), .Z(n5087) );
  XOR U7136 ( .A(n5088), .B(n5087), .Z(\w1[3][9] ) );
  XOR U7137 ( .A(\w3[3][8] ), .B(key[512]), .Z(n5090) );
  XOR U7138 ( .A(\w3[3][1] ), .B(\w3[3][25] ), .Z(n5512) );
  XOR U7139 ( .A(\w3[3][16] ), .B(\w3[3][24] ), .Z(n5468) );
  XNOR U7140 ( .A(n5512), .B(n5468), .Z(n5089) );
  XNOR U7141 ( .A(n5090), .B(n5089), .Z(\w1[4][0] ) );
  XOR U7142 ( .A(\w3[3][96] ), .B(\w3[3][101] ), .Z(n5115) );
  XOR U7143 ( .A(n5115), .B(key[612]), .Z(n5094) );
  XOR U7144 ( .A(\w3[3][116] ), .B(\w3[3][125] ), .Z(n5092) );
  XNOR U7145 ( .A(\w3[3][120] ), .B(\w3[3][108] ), .Z(n5091) );
  XNOR U7146 ( .A(n5092), .B(n5091), .Z(n5173) );
  XNOR U7147 ( .A(\w3[3][124] ), .B(n5173), .Z(n5093) );
  XNOR U7148 ( .A(n5094), .B(n5093), .Z(\w1[4][100] ) );
  XOR U7149 ( .A(\w3[3][102] ), .B(\w3[3][126] ), .Z(n5124) );
  XOR U7150 ( .A(n5124), .B(key[613]), .Z(n5096) );
  XOR U7151 ( .A(\w3[3][109] ), .B(\w3[3][117] ), .Z(n5176) );
  XNOR U7152 ( .A(\w3[3][125] ), .B(n5176), .Z(n5095) );
  XNOR U7153 ( .A(n5096), .B(n5095), .Z(\w1[4][101] ) );
  XOR U7154 ( .A(\w3[3][96] ), .B(\w3[3][103] ), .Z(n5125) );
  XOR U7155 ( .A(n5125), .B(key[614]), .Z(n5098) );
  XOR U7156 ( .A(\w3[3][110] ), .B(\w3[3][118] ), .Z(n5143) );
  XNOR U7157 ( .A(\w3[3][120] ), .B(\w3[3][127] ), .Z(n5100) );
  XNOR U7158 ( .A(n5143), .B(n5100), .Z(n5181) );
  XNOR U7159 ( .A(\w3[3][126] ), .B(n5181), .Z(n5097) );
  XNOR U7160 ( .A(n5098), .B(n5097), .Z(\w1[4][102] ) );
  XOR U7161 ( .A(\w3[3][111] ), .B(\w3[3][119] ), .Z(n5184) );
  XNOR U7162 ( .A(n5184), .B(key[615]), .Z(n5099) );
  XNOR U7163 ( .A(n5100), .B(n5099), .Z(n5101) );
  XNOR U7164 ( .A(\w3[3][96] ), .B(n5101), .Z(\w1[4][103] ) );
  XOR U7165 ( .A(key[616]), .B(\w3[3][105] ), .Z(n5103) );
  XOR U7166 ( .A(\w3[3][120] ), .B(\w3[3][112] ), .Z(n5494) );
  XNOR U7167 ( .A(\w3[3][96] ), .B(n5494), .Z(n5102) );
  XNOR U7168 ( .A(n5103), .B(n5102), .Z(n5104) );
  XOR U7169 ( .A(\w3[3][97] ), .B(n5104), .Z(\w1[4][104] ) );
  XOR U7170 ( .A(\w3[3][106] ), .B(\w3[3][98] ), .Z(n5166) );
  XOR U7171 ( .A(n5166), .B(key[617]), .Z(n5106) );
  XOR U7172 ( .A(\w3[3][97] ), .B(\w3[3][121] ), .Z(n5493) );
  XNOR U7173 ( .A(\w3[3][113] ), .B(n5493), .Z(n5105) );
  XNOR U7174 ( .A(n5106), .B(n5105), .Z(\w1[4][105] ) );
  XOR U7175 ( .A(\w3[3][107] ), .B(\w3[3][114] ), .Z(n5108) );
  XOR U7176 ( .A(\w3[3][98] ), .B(\w3[3][122] ), .Z(n5498) );
  XNOR U7177 ( .A(n5498), .B(key[618]), .Z(n5107) );
  XNOR U7178 ( .A(n5108), .B(n5107), .Z(n5109) );
  XOR U7179 ( .A(\w3[3][99] ), .B(n5109), .Z(\w1[4][106] ) );
  XOR U7180 ( .A(\w3[3][99] ), .B(\w3[3][123] ), .Z(n5502) );
  XNOR U7181 ( .A(\w3[3][108] ), .B(n5502), .Z(n5110) );
  XNOR U7182 ( .A(\w3[3][104] ), .B(n5110), .Z(n5136) );
  XOR U7183 ( .A(n5136), .B(key[619]), .Z(n5112) );
  XOR U7184 ( .A(\w3[3][96] ), .B(\w3[3][100] ), .Z(n5506) );
  XNOR U7185 ( .A(\w3[3][115] ), .B(n5506), .Z(n5111) );
  XNOR U7186 ( .A(n5112), .B(n5111), .Z(\w1[4][107] ) );
  XOR U7187 ( .A(\w3[3][100] ), .B(\w3[3][104] ), .Z(n5114) );
  XNOR U7188 ( .A(\w3[3][124] ), .B(\w3[3][109] ), .Z(n5113) );
  XNOR U7189 ( .A(n5114), .B(n5113), .Z(n5139) );
  XOR U7190 ( .A(n5139), .B(key[620]), .Z(n5117) );
  XNOR U7191 ( .A(\w3[3][116] ), .B(n5115), .Z(n5116) );
  XNOR U7192 ( .A(n5117), .B(n5116), .Z(\w1[4][108] ) );
  XOR U7193 ( .A(\w3[3][125] ), .B(\w3[3][101] ), .Z(n5142) );
  XOR U7194 ( .A(n5142), .B(key[621]), .Z(n5119) );
  XNOR U7195 ( .A(\w3[3][102] ), .B(\w3[3][110] ), .Z(n5118) );
  XNOR U7196 ( .A(n5119), .B(n5118), .Z(n5120) );
  XOR U7197 ( .A(\w3[3][117] ), .B(n5120), .Z(\w1[4][109] ) );
  XOR U7198 ( .A(\w3[3][11] ), .B(\w3[3][18] ), .Z(n5122) );
  XOR U7199 ( .A(\w3[3][2] ), .B(\w3[3][26] ), .Z(n5207) );
  XNOR U7200 ( .A(n5207), .B(key[522]), .Z(n5121) );
  XNOR U7201 ( .A(n5122), .B(n5121), .Z(n5123) );
  XOR U7202 ( .A(\w3[3][3] ), .B(n5123), .Z(\w1[4][10] ) );
  XNOR U7203 ( .A(\w3[3][111] ), .B(\w3[3][104] ), .Z(n5151) );
  XNOR U7204 ( .A(n5124), .B(n5151), .Z(n5146) );
  XOR U7205 ( .A(n5146), .B(key[622]), .Z(n5127) );
  XNOR U7206 ( .A(\w3[3][118] ), .B(n5125), .Z(n5126) );
  XNOR U7207 ( .A(n5127), .B(n5126), .Z(\w1[4][110] ) );
  XOR U7208 ( .A(\w3[3][127] ), .B(\w3[3][103] ), .Z(n5149) );
  XOR U7209 ( .A(n5149), .B(key[623]), .Z(n5129) );
  XOR U7210 ( .A(\w3[3][96] ), .B(\w3[3][104] ), .Z(n5156) );
  XNOR U7211 ( .A(\w3[3][119] ), .B(n5156), .Z(n5128) );
  XNOR U7212 ( .A(n5129), .B(n5128), .Z(\w1[4][111] ) );
  XOR U7213 ( .A(\w3[3][105] ), .B(\w3[3][113] ), .Z(n5497) );
  XOR U7214 ( .A(n5497), .B(key[624]), .Z(n5131) );
  XNOR U7215 ( .A(\w3[3][120] ), .B(n5156), .Z(n5130) );
  XNOR U7216 ( .A(n5131), .B(n5130), .Z(\w1[4][112] ) );
  XOR U7217 ( .A(\w3[3][106] ), .B(\w3[3][114] ), .Z(n5501) );
  XOR U7218 ( .A(n5501), .B(key[625]), .Z(n5133) );
  XNOR U7219 ( .A(\w3[3][105] ), .B(n5493), .Z(n5132) );
  XNOR U7220 ( .A(n5133), .B(n5132), .Z(\w1[4][113] ) );
  XOR U7221 ( .A(\w3[3][107] ), .B(\w3[3][115] ), .Z(n5168) );
  XOR U7222 ( .A(n5168), .B(key[626]), .Z(n5135) );
  XNOR U7223 ( .A(n5166), .B(\w3[3][122] ), .Z(n5134) );
  XNOR U7224 ( .A(n5135), .B(n5134), .Z(\w1[4][114] ) );
  XOR U7225 ( .A(\w3[3][116] ), .B(\w3[3][112] ), .Z(n5169) );
  XOR U7226 ( .A(n5169), .B(key[627]), .Z(n5138) );
  XNOR U7227 ( .A(\w3[3][107] ), .B(n5136), .Z(n5137) );
  XNOR U7228 ( .A(n5138), .B(n5137), .Z(\w1[4][115] ) );
  XOR U7229 ( .A(\w3[3][117] ), .B(\w3[3][112] ), .Z(n5172) );
  XOR U7230 ( .A(n5172), .B(key[628]), .Z(n5141) );
  XNOR U7231 ( .A(\w3[3][108] ), .B(n5139), .Z(n5140) );
  XNOR U7232 ( .A(n5141), .B(n5140), .Z(\w1[4][116] ) );
  XOR U7233 ( .A(n5142), .B(key[629]), .Z(n5145) );
  XNOR U7234 ( .A(\w3[3][109] ), .B(n5143), .Z(n5144) );
  XNOR U7235 ( .A(n5145), .B(n5144), .Z(\w1[4][117] ) );
  XOR U7236 ( .A(\w3[3][119] ), .B(\w3[3][112] ), .Z(n5180) );
  XOR U7237 ( .A(n5180), .B(key[630]), .Z(n5148) );
  XNOR U7238 ( .A(\w3[3][110] ), .B(n5146), .Z(n5147) );
  XNOR U7239 ( .A(n5148), .B(n5147), .Z(\w1[4][118] ) );
  XNOR U7240 ( .A(n5149), .B(key[631]), .Z(n5150) );
  XNOR U7241 ( .A(n5151), .B(n5150), .Z(n5152) );
  XNOR U7242 ( .A(\w3[3][112] ), .B(n5152), .Z(\w1[4][119] ) );
  XOR U7243 ( .A(\w3[3][3] ), .B(\w3[3][27] ), .Z(n5248) );
  XNOR U7244 ( .A(\w3[3][8] ), .B(\w3[3][12] ), .Z(n5153) );
  XNOR U7245 ( .A(n5248), .B(n5153), .Z(n5204) );
  XOR U7246 ( .A(n5204), .B(key[523]), .Z(n5155) );
  XOR U7247 ( .A(\w3[3][0] ), .B(\w3[3][4] ), .Z(n5278) );
  XNOR U7248 ( .A(\w3[3][19] ), .B(n5278), .Z(n5154) );
  XNOR U7249 ( .A(n5155), .B(n5154), .Z(\w1[4][11] ) );
  XOR U7250 ( .A(n5156), .B(key[632]), .Z(n5158) );
  XNOR U7251 ( .A(\w3[3][113] ), .B(\w3[3][121] ), .Z(n5157) );
  XNOR U7252 ( .A(n5158), .B(n5157), .Z(n5159) );
  XOR U7253 ( .A(\w3[3][112] ), .B(n5159), .Z(\w1[4][120] ) );
  XOR U7254 ( .A(n5497), .B(key[633]), .Z(n5161) );
  XNOR U7255 ( .A(\w3[3][122] ), .B(\w3[3][114] ), .Z(n5160) );
  XNOR U7256 ( .A(n5161), .B(n5160), .Z(n5162) );
  XOR U7257 ( .A(\w3[3][97] ), .B(n5162), .Z(\w1[4][121] ) );
  XOR U7258 ( .A(\w3[3][123] ), .B(key[634]), .Z(n5164) );
  XNOR U7259 ( .A(\w3[3][114] ), .B(\w3[3][115] ), .Z(n5163) );
  XNOR U7260 ( .A(n5164), .B(n5163), .Z(n5165) );
  XOR U7261 ( .A(n5166), .B(n5165), .Z(\w1[4][122] ) );
  XNOR U7262 ( .A(\w3[3][124] ), .B(\w3[3][120] ), .Z(n5167) );
  XNOR U7263 ( .A(n5168), .B(n5167), .Z(n5505) );
  XOR U7264 ( .A(n5505), .B(key[635]), .Z(n5171) );
  XNOR U7265 ( .A(\w3[3][99] ), .B(n5169), .Z(n5170) );
  XNOR U7266 ( .A(n5171), .B(n5170), .Z(\w1[4][123] ) );
  XOR U7267 ( .A(n5172), .B(key[636]), .Z(n5175) );
  XNOR U7268 ( .A(n5173), .B(\w3[3][100] ), .Z(n5174) );
  XNOR U7269 ( .A(n5175), .B(n5174), .Z(\w1[4][124] ) );
  XOR U7270 ( .A(\w3[3][118] ), .B(key[637]), .Z(n5178) );
  XNOR U7271 ( .A(n5176), .B(\w3[3][126] ), .Z(n5177) );
  XNOR U7272 ( .A(n5178), .B(n5177), .Z(n5179) );
  XOR U7273 ( .A(\w3[3][101] ), .B(n5179), .Z(\w1[4][125] ) );
  XOR U7274 ( .A(n5180), .B(key[638]), .Z(n5183) );
  XNOR U7275 ( .A(\w3[3][102] ), .B(n5181), .Z(n5182) );
  XNOR U7276 ( .A(n5183), .B(n5182), .Z(\w1[4][126] ) );
  XOR U7277 ( .A(n5494), .B(key[639]), .Z(n5186) );
  XNOR U7278 ( .A(\w3[3][103] ), .B(n5184), .Z(n5185) );
  XNOR U7279 ( .A(n5186), .B(n5185), .Z(\w1[4][127] ) );
  XOR U7280 ( .A(\w3[3][13] ), .B(\w3[3][28] ), .Z(n5188) );
  XNOR U7281 ( .A(\w3[3][8] ), .B(\w3[3][4] ), .Z(n5187) );
  XNOR U7282 ( .A(n5188), .B(n5187), .Z(n5210) );
  XOR U7283 ( .A(n5210), .B(key[524]), .Z(n5190) );
  XOR U7284 ( .A(\w3[3][0] ), .B(\w3[3][5] ), .Z(n5315) );
  XNOR U7285 ( .A(\w3[3][20] ), .B(n5315), .Z(n5189) );
  XNOR U7286 ( .A(n5190), .B(n5189), .Z(\w1[4][12] ) );
  XOR U7287 ( .A(\w3[3][14] ), .B(\w3[3][6] ), .Z(n5192) );
  XOR U7288 ( .A(\w3[3][5] ), .B(\w3[3][29] ), .Z(n5213) );
  XNOR U7289 ( .A(n5213), .B(key[525]), .Z(n5191) );
  XNOR U7290 ( .A(n5192), .B(n5191), .Z(n5193) );
  XOR U7291 ( .A(\w3[3][21] ), .B(n5193), .Z(\w1[4][13] ) );
  XOR U7292 ( .A(\w3[3][6] ), .B(\w3[3][30] ), .Z(n5356) );
  XNOR U7293 ( .A(\w3[3][8] ), .B(\w3[3][15] ), .Z(n5221) );
  XNOR U7294 ( .A(n5356), .B(n5221), .Z(n5216) );
  XOR U7295 ( .A(n5216), .B(key[526]), .Z(n5195) );
  XOR U7296 ( .A(\w3[3][0] ), .B(\w3[3][7] ), .Z(n5391) );
  XNOR U7297 ( .A(\w3[3][22] ), .B(n5391), .Z(n5194) );
  XNOR U7298 ( .A(n5195), .B(n5194), .Z(\w1[4][14] ) );
  XOR U7299 ( .A(\w3[3][7] ), .B(\w3[3][31] ), .Z(n5219) );
  XOR U7300 ( .A(n5219), .B(key[527]), .Z(n5197) );
  XOR U7301 ( .A(\w3[3][8] ), .B(\w3[3][0] ), .Z(n5223) );
  XNOR U7302 ( .A(\w3[3][23] ), .B(n5223), .Z(n5196) );
  XNOR U7303 ( .A(n5197), .B(n5196), .Z(\w1[4][15] ) );
  XOR U7304 ( .A(\w3[3][17] ), .B(\w3[3][9] ), .Z(n5227) );
  XOR U7305 ( .A(n5227), .B(key[528]), .Z(n5199) );
  XNOR U7306 ( .A(\w3[3][24] ), .B(n5223), .Z(n5198) );
  XNOR U7307 ( .A(n5199), .B(n5198), .Z(\w1[4][16] ) );
  XOR U7308 ( .A(\w3[3][18] ), .B(\w3[3][10] ), .Z(n5247) );
  XOR U7309 ( .A(n5247), .B(key[529]), .Z(n5201) );
  XNOR U7310 ( .A(n5512), .B(\w3[3][9] ), .Z(n5200) );
  XNOR U7311 ( .A(n5201), .B(n5200), .Z(\w1[4][17] ) );
  XOR U7312 ( .A(\w3[3][11] ), .B(\w3[3][19] ), .Z(n5235) );
  XOR U7313 ( .A(n5235), .B(key[530]), .Z(n5203) );
  XNOR U7314 ( .A(n5207), .B(\w3[3][10] ), .Z(n5202) );
  XNOR U7315 ( .A(n5203), .B(n5202), .Z(\w1[4][18] ) );
  XOR U7316 ( .A(\w3[3][16] ), .B(\w3[3][20] ), .Z(n5236) );
  XOR U7317 ( .A(n5236), .B(key[531]), .Z(n5206) );
  XNOR U7318 ( .A(\w3[3][11] ), .B(n5204), .Z(n5205) );
  XNOR U7319 ( .A(n5206), .B(n5205), .Z(\w1[4][19] ) );
  XOR U7320 ( .A(n5227), .B(key[513]), .Z(n5209) );
  XNOR U7321 ( .A(\w3[3][25] ), .B(n5207), .Z(n5208) );
  XNOR U7322 ( .A(n5209), .B(n5208), .Z(\w1[4][1] ) );
  XOR U7323 ( .A(\w3[3][16] ), .B(\w3[3][21] ), .Z(n5241) );
  XOR U7324 ( .A(n5241), .B(key[532]), .Z(n5212) );
  XNOR U7325 ( .A(\w3[3][12] ), .B(n5210), .Z(n5211) );
  XNOR U7326 ( .A(n5212), .B(n5211), .Z(\w1[4][20] ) );
  XOR U7327 ( .A(\w3[3][14] ), .B(\w3[3][22] ), .Z(n5251) );
  XOR U7328 ( .A(n5251), .B(key[533]), .Z(n5215) );
  XNOR U7329 ( .A(\w3[3][13] ), .B(n5213), .Z(n5214) );
  XNOR U7330 ( .A(n5215), .B(n5214), .Z(\w1[4][21] ) );
  XOR U7331 ( .A(\w3[3][16] ), .B(\w3[3][23] ), .Z(n5252) );
  XOR U7332 ( .A(n5252), .B(key[534]), .Z(n5218) );
  XNOR U7333 ( .A(\w3[3][14] ), .B(n5216), .Z(n5217) );
  XNOR U7334 ( .A(n5218), .B(n5217), .Z(\w1[4][22] ) );
  XNOR U7335 ( .A(n5219), .B(key[535]), .Z(n5220) );
  XNOR U7336 ( .A(n5221), .B(n5220), .Z(n5222) );
  XNOR U7337 ( .A(\w3[3][16] ), .B(n5222), .Z(\w1[4][23] ) );
  XOR U7338 ( .A(\w3[3][17] ), .B(key[536]), .Z(n5225) );
  XNOR U7339 ( .A(\w3[3][25] ), .B(n5223), .Z(n5224) );
  XNOR U7340 ( .A(n5225), .B(n5224), .Z(n5226) );
  XOR U7341 ( .A(\w3[3][16] ), .B(n5226), .Z(\w1[4][24] ) );
  XOR U7342 ( .A(n5227), .B(key[537]), .Z(n5229) );
  XNOR U7343 ( .A(\w3[3][1] ), .B(\w3[3][26] ), .Z(n5228) );
  XNOR U7344 ( .A(n5229), .B(n5228), .Z(n5230) );
  XOR U7345 ( .A(\w3[3][18] ), .B(n5230), .Z(\w1[4][25] ) );
  XOR U7346 ( .A(n5247), .B(key[538]), .Z(n5232) );
  XNOR U7347 ( .A(\w3[3][2] ), .B(\w3[3][19] ), .Z(n5231) );
  XNOR U7348 ( .A(n5232), .B(n5231), .Z(n5233) );
  XOR U7349 ( .A(\w3[3][27] ), .B(n5233), .Z(\w1[4][26] ) );
  XNOR U7350 ( .A(\w3[3][24] ), .B(\w3[3][28] ), .Z(n5234) );
  XNOR U7351 ( .A(n5235), .B(n5234), .Z(n5277) );
  XOR U7352 ( .A(n5277), .B(key[539]), .Z(n5238) );
  XNOR U7353 ( .A(\w3[3][3] ), .B(n5236), .Z(n5237) );
  XNOR U7354 ( .A(n5238), .B(n5237), .Z(\w1[4][27] ) );
  XOR U7355 ( .A(\w3[3][20] ), .B(\w3[3][29] ), .Z(n5240) );
  XNOR U7356 ( .A(\w3[3][24] ), .B(\w3[3][12] ), .Z(n5239) );
  XNOR U7357 ( .A(n5240), .B(n5239), .Z(n5314) );
  XOR U7358 ( .A(n5314), .B(key[540]), .Z(n5243) );
  XNOR U7359 ( .A(\w3[3][4] ), .B(n5241), .Z(n5242) );
  XNOR U7360 ( .A(n5243), .B(n5242), .Z(\w1[4][28] ) );
  XOR U7361 ( .A(\w3[3][13] ), .B(\w3[3][21] ), .Z(n5355) );
  XOR U7362 ( .A(n5355), .B(key[541]), .Z(n5245) );
  XNOR U7363 ( .A(\w3[3][22] ), .B(\w3[3][30] ), .Z(n5244) );
  XNOR U7364 ( .A(n5245), .B(n5244), .Z(n5246) );
  XOR U7365 ( .A(\w3[3][5] ), .B(n5246), .Z(\w1[4][29] ) );
  XOR U7366 ( .A(n5247), .B(key[514]), .Z(n5250) );
  XNOR U7367 ( .A(\w3[3][26] ), .B(n5248), .Z(n5249) );
  XNOR U7368 ( .A(n5250), .B(n5249), .Z(\w1[4][2] ) );
  XNOR U7369 ( .A(\w3[3][24] ), .B(\w3[3][31] ), .Z(n5429) );
  XNOR U7370 ( .A(n5251), .B(n5429), .Z(n5390) );
  XOR U7371 ( .A(n5390), .B(key[542]), .Z(n5254) );
  XNOR U7372 ( .A(\w3[3][6] ), .B(n5252), .Z(n5253) );
  XNOR U7373 ( .A(n5254), .B(n5253), .Z(\w1[4][30] ) );
  XOR U7374 ( .A(\w3[3][15] ), .B(\w3[3][23] ), .Z(n5427) );
  XOR U7375 ( .A(n5427), .B(key[543]), .Z(n5256) );
  XNOR U7376 ( .A(n5468), .B(\w3[3][7] ), .Z(n5255) );
  XNOR U7377 ( .A(n5256), .B(n5255), .Z(\w1[4][31] ) );
  XOR U7378 ( .A(\w3[3][33] ), .B(\w3[3][57] ), .Z(n5311) );
  XOR U7379 ( .A(n5311), .B(key[544]), .Z(n5258) );
  XOR U7380 ( .A(\w3[3][48] ), .B(\w3[3][56] ), .Z(n5372) );
  XNOR U7381 ( .A(n5372), .B(\w3[3][40] ), .Z(n5257) );
  XNOR U7382 ( .A(n5258), .B(n5257), .Z(\w1[4][32] ) );
  XOR U7383 ( .A(\w3[3][34] ), .B(\w3[3][58] ), .Z(n5319) );
  XOR U7384 ( .A(n5319), .B(key[545]), .Z(n5260) );
  XOR U7385 ( .A(\w3[3][41] ), .B(\w3[3][49] ), .Z(n5343) );
  XNOR U7386 ( .A(\w3[3][57] ), .B(n5343), .Z(n5259) );
  XNOR U7387 ( .A(n5260), .B(n5259), .Z(\w1[4][33] ) );
  XOR U7388 ( .A(\w3[3][35] ), .B(\w3[3][59] ), .Z(n5290) );
  XOR U7389 ( .A(n5290), .B(key[546]), .Z(n5262) );
  XOR U7390 ( .A(\w3[3][42] ), .B(\w3[3][50] ), .Z(n5347) );
  XNOR U7391 ( .A(\w3[3][58] ), .B(n5347), .Z(n5261) );
  XNOR U7392 ( .A(n5262), .B(n5261), .Z(\w1[4][34] ) );
  XOR U7393 ( .A(\w3[3][36] ), .B(\w3[3][32] ), .Z(n5292) );
  XOR U7394 ( .A(n5292), .B(key[547]), .Z(n5265) );
  XOR U7395 ( .A(\w3[3][43] ), .B(\w3[3][51] ), .Z(n5318) );
  XNOR U7396 ( .A(\w3[3][56] ), .B(n5318), .Z(n5263) );
  XNOR U7397 ( .A(\w3[3][60] ), .B(n5263), .Z(n5352) );
  XNOR U7398 ( .A(\w3[3][59] ), .B(n5352), .Z(n5264) );
  XNOR U7399 ( .A(n5265), .B(n5264), .Z(\w1[4][35] ) );
  XOR U7400 ( .A(\w3[3][32] ), .B(\w3[3][37] ), .Z(n5297) );
  XOR U7401 ( .A(n5297), .B(key[548]), .Z(n5269) );
  XOR U7402 ( .A(\w3[3][52] ), .B(\w3[3][61] ), .Z(n5267) );
  XNOR U7403 ( .A(\w3[3][56] ), .B(\w3[3][44] ), .Z(n5266) );
  XNOR U7404 ( .A(n5267), .B(n5266), .Z(n5360) );
  XNOR U7405 ( .A(\w3[3][60] ), .B(n5360), .Z(n5268) );
  XNOR U7406 ( .A(n5269), .B(n5268), .Z(\w1[4][36] ) );
  XOR U7407 ( .A(\w3[3][38] ), .B(\w3[3][62] ), .Z(n5303) );
  XOR U7408 ( .A(n5303), .B(key[549]), .Z(n5271) );
  XOR U7409 ( .A(\w3[3][45] ), .B(\w3[3][53] ), .Z(n5363) );
  XNOR U7410 ( .A(\w3[3][61] ), .B(n5363), .Z(n5270) );
  XNOR U7411 ( .A(n5271), .B(n5270), .Z(\w1[4][37] ) );
  XOR U7412 ( .A(\w3[3][32] ), .B(\w3[3][39] ), .Z(n5304) );
  XOR U7413 ( .A(n5304), .B(key[550]), .Z(n5273) );
  XOR U7414 ( .A(\w3[3][46] ), .B(\w3[3][54] ), .Z(n5329) );
  XNOR U7415 ( .A(\w3[3][56] ), .B(\w3[3][63] ), .Z(n5275) );
  XNOR U7416 ( .A(n5329), .B(n5275), .Z(n5368) );
  XNOR U7417 ( .A(\w3[3][62] ), .B(n5368), .Z(n5272) );
  XNOR U7418 ( .A(n5273), .B(n5272), .Z(\w1[4][38] ) );
  XOR U7419 ( .A(\w3[3][47] ), .B(\w3[3][55] ), .Z(n5371) );
  XNOR U7420 ( .A(n5371), .B(key[551]), .Z(n5274) );
  XNOR U7421 ( .A(n5275), .B(n5274), .Z(n5276) );
  XNOR U7422 ( .A(\w3[3][32] ), .B(n5276), .Z(\w1[4][39] ) );
  XOR U7423 ( .A(n5277), .B(key[515]), .Z(n5280) );
  XNOR U7424 ( .A(n5278), .B(\w3[3][27] ), .Z(n5279) );
  XNOR U7425 ( .A(n5280), .B(n5279), .Z(\w1[4][3] ) );
  XOR U7426 ( .A(\w3[3][32] ), .B(key[552]), .Z(n5282) );
  XNOR U7427 ( .A(\w3[3][33] ), .B(\w3[3][41] ), .Z(n5281) );
  XNOR U7428 ( .A(n5282), .B(n5281), .Z(n5283) );
  XOR U7429 ( .A(n5372), .B(n5283), .Z(\w1[4][40] ) );
  XOR U7430 ( .A(\w3[3][42] ), .B(key[553]), .Z(n5285) );
  XNOR U7431 ( .A(\w3[3][49] ), .B(\w3[3][34] ), .Z(n5284) );
  XNOR U7432 ( .A(n5285), .B(n5284), .Z(n5286) );
  XOR U7433 ( .A(n5311), .B(n5286), .Z(\w1[4][41] ) );
  XOR U7434 ( .A(\w3[3][43] ), .B(key[554]), .Z(n5288) );
  XNOR U7435 ( .A(\w3[3][50] ), .B(\w3[3][35] ), .Z(n5287) );
  XNOR U7436 ( .A(n5288), .B(n5287), .Z(n5289) );
  XOR U7437 ( .A(n5319), .B(n5289), .Z(\w1[4][42] ) );
  XNOR U7438 ( .A(\w3[3][40] ), .B(n5290), .Z(n5291) );
  XNOR U7439 ( .A(\w3[3][44] ), .B(n5291), .Z(n5322) );
  XOR U7440 ( .A(n5322), .B(key[555]), .Z(n5294) );
  XNOR U7441 ( .A(\w3[3][51] ), .B(n5292), .Z(n5293) );
  XNOR U7442 ( .A(n5294), .B(n5293), .Z(\w1[4][43] ) );
  XOR U7443 ( .A(\w3[3][36] ), .B(\w3[3][45] ), .Z(n5296) );
  XNOR U7444 ( .A(\w3[3][40] ), .B(\w3[3][60] ), .Z(n5295) );
  XNOR U7445 ( .A(n5296), .B(n5295), .Z(n5325) );
  XOR U7446 ( .A(n5325), .B(key[556]), .Z(n5299) );
  XNOR U7447 ( .A(\w3[3][52] ), .B(n5297), .Z(n5298) );
  XNOR U7448 ( .A(n5299), .B(n5298), .Z(\w1[4][44] ) );
  XOR U7449 ( .A(\w3[3][61] ), .B(\w3[3][37] ), .Z(n5328) );
  XOR U7450 ( .A(n5328), .B(key[557]), .Z(n5301) );
  XNOR U7451 ( .A(\w3[3][38] ), .B(\w3[3][46] ), .Z(n5300) );
  XNOR U7452 ( .A(n5301), .B(n5300), .Z(n5302) );
  XOR U7453 ( .A(\w3[3][53] ), .B(n5302), .Z(\w1[4][45] ) );
  XNOR U7454 ( .A(\w3[3][40] ), .B(\w3[3][47] ), .Z(n5337) );
  XNOR U7455 ( .A(n5303), .B(n5337), .Z(n5332) );
  XOR U7456 ( .A(n5332), .B(key[558]), .Z(n5306) );
  XNOR U7457 ( .A(\w3[3][54] ), .B(n5304), .Z(n5305) );
  XNOR U7458 ( .A(n5306), .B(n5305), .Z(\w1[4][46] ) );
  XOR U7459 ( .A(\w3[3][63] ), .B(\w3[3][39] ), .Z(n5335) );
  XOR U7460 ( .A(n5335), .B(key[559]), .Z(n5308) );
  XOR U7461 ( .A(\w3[3][40] ), .B(\w3[3][32] ), .Z(n5339) );
  XNOR U7462 ( .A(\w3[3][55] ), .B(n5339), .Z(n5307) );
  XNOR U7463 ( .A(n5308), .B(n5307), .Z(\w1[4][47] ) );
  XOR U7464 ( .A(n5339), .B(key[560]), .Z(n5310) );
  XNOR U7465 ( .A(\w3[3][56] ), .B(n5343), .Z(n5309) );
  XNOR U7466 ( .A(n5310), .B(n5309), .Z(\w1[4][48] ) );
  XOR U7467 ( .A(n5347), .B(key[561]), .Z(n5313) );
  XNOR U7468 ( .A(n5311), .B(\w3[3][41] ), .Z(n5312) );
  XNOR U7469 ( .A(n5313), .B(n5312), .Z(\w1[4][49] ) );
  XOR U7470 ( .A(n5314), .B(key[516]), .Z(n5317) );
  XNOR U7471 ( .A(n5315), .B(\w3[3][28] ), .Z(n5316) );
  XNOR U7472 ( .A(n5317), .B(n5316), .Z(\w1[4][4] ) );
  XOR U7473 ( .A(n5318), .B(key[562]), .Z(n5321) );
  XNOR U7474 ( .A(n5319), .B(\w3[3][42] ), .Z(n5320) );
  XNOR U7475 ( .A(n5321), .B(n5320), .Z(\w1[4][50] ) );
  XOR U7476 ( .A(\w3[3][48] ), .B(\w3[3][52] ), .Z(n5351) );
  XOR U7477 ( .A(n5351), .B(key[563]), .Z(n5324) );
  XNOR U7478 ( .A(\w3[3][43] ), .B(n5322), .Z(n5323) );
  XNOR U7479 ( .A(n5324), .B(n5323), .Z(\w1[4][51] ) );
  XOR U7480 ( .A(\w3[3][48] ), .B(\w3[3][53] ), .Z(n5359) );
  XOR U7481 ( .A(n5359), .B(key[564]), .Z(n5327) );
  XNOR U7482 ( .A(\w3[3][44] ), .B(n5325), .Z(n5326) );
  XNOR U7483 ( .A(n5327), .B(n5326), .Z(\w1[4][52] ) );
  XOR U7484 ( .A(n5328), .B(key[565]), .Z(n5331) );
  XNOR U7485 ( .A(\w3[3][45] ), .B(n5329), .Z(n5330) );
  XNOR U7486 ( .A(n5331), .B(n5330), .Z(\w1[4][53] ) );
  XOR U7487 ( .A(\w3[3][48] ), .B(\w3[3][55] ), .Z(n5367) );
  XOR U7488 ( .A(n5367), .B(key[566]), .Z(n5334) );
  XNOR U7489 ( .A(\w3[3][46] ), .B(n5332), .Z(n5333) );
  XNOR U7490 ( .A(n5334), .B(n5333), .Z(\w1[4][54] ) );
  XNOR U7491 ( .A(n5335), .B(key[567]), .Z(n5336) );
  XNOR U7492 ( .A(n5337), .B(n5336), .Z(n5338) );
  XNOR U7493 ( .A(\w3[3][48] ), .B(n5338), .Z(\w1[4][55] ) );
  XOR U7494 ( .A(n5339), .B(key[568]), .Z(n5341) );
  XNOR U7495 ( .A(\w3[3][48] ), .B(\w3[3][49] ), .Z(n5340) );
  XNOR U7496 ( .A(n5341), .B(n5340), .Z(n5342) );
  XOR U7497 ( .A(\w3[3][57] ), .B(n5342), .Z(\w1[4][56] ) );
  XOR U7498 ( .A(\w3[3][50] ), .B(key[569]), .Z(n5345) );
  XNOR U7499 ( .A(n5343), .B(\w3[3][58] ), .Z(n5344) );
  XNOR U7500 ( .A(n5345), .B(n5344), .Z(n5346) );
  XOR U7501 ( .A(\w3[3][33] ), .B(n5346), .Z(\w1[4][57] ) );
  XOR U7502 ( .A(\w3[3][51] ), .B(key[570]), .Z(n5349) );
  XNOR U7503 ( .A(n5347), .B(\w3[3][59] ), .Z(n5348) );
  XNOR U7504 ( .A(n5349), .B(n5348), .Z(n5350) );
  XOR U7505 ( .A(\w3[3][34] ), .B(n5350), .Z(\w1[4][58] ) );
  XOR U7506 ( .A(n5351), .B(key[571]), .Z(n5354) );
  XNOR U7507 ( .A(\w3[3][35] ), .B(n5352), .Z(n5353) );
  XNOR U7508 ( .A(n5354), .B(n5353), .Z(\w1[4][59] ) );
  XOR U7509 ( .A(n5355), .B(key[517]), .Z(n5358) );
  XNOR U7510 ( .A(\w3[3][29] ), .B(n5356), .Z(n5357) );
  XNOR U7511 ( .A(n5358), .B(n5357), .Z(\w1[4][5] ) );
  XOR U7512 ( .A(n5359), .B(key[572]), .Z(n5362) );
  XNOR U7513 ( .A(\w3[3][36] ), .B(n5360), .Z(n5361) );
  XNOR U7514 ( .A(n5362), .B(n5361), .Z(\w1[4][60] ) );
  XOR U7515 ( .A(\w3[3][54] ), .B(key[573]), .Z(n5365) );
  XNOR U7516 ( .A(n5363), .B(\w3[3][62] ), .Z(n5364) );
  XNOR U7517 ( .A(n5365), .B(n5364), .Z(n5366) );
  XOR U7518 ( .A(\w3[3][37] ), .B(n5366), .Z(\w1[4][61] ) );
  XOR U7519 ( .A(n5367), .B(key[574]), .Z(n5370) );
  XNOR U7520 ( .A(\w3[3][38] ), .B(n5368), .Z(n5369) );
  XNOR U7521 ( .A(n5370), .B(n5369), .Z(\w1[4][62] ) );
  XOR U7522 ( .A(n5371), .B(key[575]), .Z(n5374) );
  XNOR U7523 ( .A(n5372), .B(\w3[3][39] ), .Z(n5373) );
  XNOR U7524 ( .A(n5374), .B(n5373), .Z(\w1[4][63] ) );
  XOR U7525 ( .A(\w3[3][65] ), .B(\w3[3][89] ), .Z(n5433) );
  XOR U7526 ( .A(n5433), .B(key[576]), .Z(n5376) );
  XOR U7527 ( .A(\w3[3][80] ), .B(\w3[3][88] ), .Z(n5490) );
  XNOR U7528 ( .A(n5490), .B(\w3[3][72] ), .Z(n5375) );
  XNOR U7529 ( .A(n5376), .B(n5375), .Z(\w1[4][64] ) );
  XOR U7530 ( .A(\w3[3][66] ), .B(\w3[3][90] ), .Z(n5437) );
  XOR U7531 ( .A(n5437), .B(key[577]), .Z(n5378) );
  XOR U7532 ( .A(\w3[3][73] ), .B(\w3[3][81] ), .Z(n5461) );
  XNOR U7533 ( .A(\w3[3][89] ), .B(n5461), .Z(n5377) );
  XNOR U7534 ( .A(n5378), .B(n5377), .Z(\w1[4][65] ) );
  XOR U7535 ( .A(\w3[3][67] ), .B(\w3[3][91] ), .Z(n5408) );
  XOR U7536 ( .A(n5408), .B(key[578]), .Z(n5380) );
  XOR U7537 ( .A(\w3[3][74] ), .B(\w3[3][82] ), .Z(n5469) );
  XNOR U7538 ( .A(\w3[3][90] ), .B(n5469), .Z(n5379) );
  XNOR U7539 ( .A(n5380), .B(n5379), .Z(\w1[4][66] ) );
  XOR U7540 ( .A(\w3[3][68] ), .B(\w3[3][64] ), .Z(n5410) );
  XOR U7541 ( .A(n5410), .B(key[579]), .Z(n5383) );
  XOR U7542 ( .A(\w3[3][75] ), .B(\w3[3][83] ), .Z(n5436) );
  XNOR U7543 ( .A(\w3[3][88] ), .B(n5436), .Z(n5381) );
  XNOR U7544 ( .A(\w3[3][92] ), .B(n5381), .Z(n5474) );
  XNOR U7545 ( .A(\w3[3][91] ), .B(n5474), .Z(n5382) );
  XNOR U7546 ( .A(n5383), .B(n5382), .Z(\w1[4][67] ) );
  XOR U7547 ( .A(\w3[3][64] ), .B(\w3[3][69] ), .Z(n5415) );
  XOR U7548 ( .A(n5415), .B(key[580]), .Z(n5387) );
  XOR U7549 ( .A(\w3[3][84] ), .B(\w3[3][93] ), .Z(n5385) );
  XNOR U7550 ( .A(\w3[3][88] ), .B(\w3[3][76] ), .Z(n5384) );
  XNOR U7551 ( .A(n5385), .B(n5384), .Z(n5478) );
  XNOR U7552 ( .A(\w3[3][92] ), .B(n5478), .Z(n5386) );
  XNOR U7553 ( .A(n5387), .B(n5386), .Z(\w1[4][68] ) );
  XOR U7554 ( .A(\w3[3][70] ), .B(\w3[3][94] ), .Z(n5421) );
  XOR U7555 ( .A(n5421), .B(key[581]), .Z(n5389) );
  XOR U7556 ( .A(\w3[3][77] ), .B(\w3[3][85] ), .Z(n5481) );
  XNOR U7557 ( .A(\w3[3][93] ), .B(n5481), .Z(n5388) );
  XNOR U7558 ( .A(n5389), .B(n5388), .Z(\w1[4][69] ) );
  XOR U7559 ( .A(n5390), .B(key[518]), .Z(n5393) );
  XNOR U7560 ( .A(n5391), .B(\w3[3][30] ), .Z(n5392) );
  XNOR U7561 ( .A(n5393), .B(n5392), .Z(\w1[4][6] ) );
  XOR U7562 ( .A(\w3[3][64] ), .B(\w3[3][71] ), .Z(n5422) );
  XOR U7563 ( .A(n5422), .B(key[582]), .Z(n5395) );
  XOR U7564 ( .A(\w3[3][78] ), .B(\w3[3][86] ), .Z(n5447) );
  XNOR U7565 ( .A(\w3[3][88] ), .B(\w3[3][95] ), .Z(n5397) );
  XNOR U7566 ( .A(n5447), .B(n5397), .Z(n5486) );
  XNOR U7567 ( .A(\w3[3][94] ), .B(n5486), .Z(n5394) );
  XNOR U7568 ( .A(n5395), .B(n5394), .Z(\w1[4][70] ) );
  XOR U7569 ( .A(\w3[3][79] ), .B(\w3[3][87] ), .Z(n5489) );
  XNOR U7570 ( .A(n5489), .B(key[583]), .Z(n5396) );
  XNOR U7571 ( .A(n5397), .B(n5396), .Z(n5398) );
  XNOR U7572 ( .A(\w3[3][64] ), .B(n5398), .Z(\w1[4][71] ) );
  XOR U7573 ( .A(\w3[3][64] ), .B(key[584]), .Z(n5400) );
  XNOR U7574 ( .A(\w3[3][65] ), .B(\w3[3][73] ), .Z(n5399) );
  XNOR U7575 ( .A(n5400), .B(n5399), .Z(n5401) );
  XOR U7576 ( .A(n5490), .B(n5401), .Z(\w1[4][72] ) );
  XOR U7577 ( .A(\w3[3][74] ), .B(key[585]), .Z(n5403) );
  XNOR U7578 ( .A(\w3[3][81] ), .B(\w3[3][66] ), .Z(n5402) );
  XNOR U7579 ( .A(n5403), .B(n5402), .Z(n5404) );
  XOR U7580 ( .A(n5433), .B(n5404), .Z(\w1[4][73] ) );
  XOR U7581 ( .A(\w3[3][75] ), .B(key[586]), .Z(n5406) );
  XNOR U7582 ( .A(\w3[3][82] ), .B(\w3[3][67] ), .Z(n5405) );
  XNOR U7583 ( .A(n5406), .B(n5405), .Z(n5407) );
  XOR U7584 ( .A(n5437), .B(n5407), .Z(\w1[4][74] ) );
  XNOR U7585 ( .A(\w3[3][72] ), .B(n5408), .Z(n5409) );
  XNOR U7586 ( .A(\w3[3][76] ), .B(n5409), .Z(n5440) );
  XOR U7587 ( .A(n5440), .B(key[587]), .Z(n5412) );
  XNOR U7588 ( .A(\w3[3][83] ), .B(n5410), .Z(n5411) );
  XNOR U7589 ( .A(n5412), .B(n5411), .Z(\w1[4][75] ) );
  XOR U7590 ( .A(\w3[3][68] ), .B(\w3[3][77] ), .Z(n5414) );
  XNOR U7591 ( .A(\w3[3][72] ), .B(\w3[3][92] ), .Z(n5413) );
  XNOR U7592 ( .A(n5414), .B(n5413), .Z(n5443) );
  XOR U7593 ( .A(n5443), .B(key[588]), .Z(n5417) );
  XNOR U7594 ( .A(\w3[3][84] ), .B(n5415), .Z(n5416) );
  XNOR U7595 ( .A(n5417), .B(n5416), .Z(\w1[4][76] ) );
  XOR U7596 ( .A(\w3[3][93] ), .B(\w3[3][69] ), .Z(n5446) );
  XOR U7597 ( .A(n5446), .B(key[589]), .Z(n5419) );
  XNOR U7598 ( .A(\w3[3][70] ), .B(\w3[3][78] ), .Z(n5418) );
  XNOR U7599 ( .A(n5419), .B(n5418), .Z(n5420) );
  XOR U7600 ( .A(\w3[3][85] ), .B(n5420), .Z(\w1[4][77] ) );
  XNOR U7601 ( .A(\w3[3][72] ), .B(\w3[3][79] ), .Z(n5455) );
  XNOR U7602 ( .A(n5421), .B(n5455), .Z(n5450) );
  XOR U7603 ( .A(n5450), .B(key[590]), .Z(n5424) );
  XNOR U7604 ( .A(\w3[3][86] ), .B(n5422), .Z(n5423) );
  XNOR U7605 ( .A(n5424), .B(n5423), .Z(\w1[4][78] ) );
  XOR U7606 ( .A(\w3[3][95] ), .B(\w3[3][71] ), .Z(n5453) );
  XOR U7607 ( .A(n5453), .B(key[591]), .Z(n5426) );
  XOR U7608 ( .A(\w3[3][72] ), .B(\w3[3][64] ), .Z(n5457) );
  XNOR U7609 ( .A(\w3[3][87] ), .B(n5457), .Z(n5425) );
  XNOR U7610 ( .A(n5426), .B(n5425), .Z(\w1[4][79] ) );
  XNOR U7611 ( .A(n5427), .B(key[519]), .Z(n5428) );
  XNOR U7612 ( .A(n5429), .B(n5428), .Z(n5430) );
  XNOR U7613 ( .A(\w3[3][0] ), .B(n5430), .Z(\w1[4][7] ) );
  XOR U7614 ( .A(n5457), .B(key[592]), .Z(n5432) );
  XNOR U7615 ( .A(\w3[3][88] ), .B(n5461), .Z(n5431) );
  XNOR U7616 ( .A(n5432), .B(n5431), .Z(\w1[4][80] ) );
  XOR U7617 ( .A(n5469), .B(key[593]), .Z(n5435) );
  XNOR U7618 ( .A(n5433), .B(\w3[3][73] ), .Z(n5434) );
  XNOR U7619 ( .A(n5435), .B(n5434), .Z(\w1[4][81] ) );
  XOR U7620 ( .A(n5436), .B(key[594]), .Z(n5439) );
  XNOR U7621 ( .A(n5437), .B(\w3[3][74] ), .Z(n5438) );
  XNOR U7622 ( .A(n5439), .B(n5438), .Z(\w1[4][82] ) );
  XOR U7623 ( .A(\w3[3][80] ), .B(\w3[3][84] ), .Z(n5473) );
  XOR U7624 ( .A(n5473), .B(key[595]), .Z(n5442) );
  XNOR U7625 ( .A(\w3[3][75] ), .B(n5440), .Z(n5441) );
  XNOR U7626 ( .A(n5442), .B(n5441), .Z(\w1[4][83] ) );
  XOR U7627 ( .A(\w3[3][80] ), .B(\w3[3][85] ), .Z(n5477) );
  XOR U7628 ( .A(n5477), .B(key[596]), .Z(n5445) );
  XNOR U7629 ( .A(\w3[3][76] ), .B(n5443), .Z(n5444) );
  XNOR U7630 ( .A(n5445), .B(n5444), .Z(\w1[4][84] ) );
  XOR U7631 ( .A(n5446), .B(key[597]), .Z(n5449) );
  XNOR U7632 ( .A(\w3[3][77] ), .B(n5447), .Z(n5448) );
  XNOR U7633 ( .A(n5449), .B(n5448), .Z(\w1[4][85] ) );
  XOR U7634 ( .A(\w3[3][80] ), .B(\w3[3][87] ), .Z(n5485) );
  XOR U7635 ( .A(n5485), .B(key[598]), .Z(n5452) );
  XNOR U7636 ( .A(\w3[3][78] ), .B(n5450), .Z(n5451) );
  XNOR U7637 ( .A(n5452), .B(n5451), .Z(\w1[4][86] ) );
  XNOR U7638 ( .A(n5453), .B(key[599]), .Z(n5454) );
  XNOR U7639 ( .A(n5455), .B(n5454), .Z(n5456) );
  XNOR U7640 ( .A(\w3[3][80] ), .B(n5456), .Z(\w1[4][87] ) );
  XOR U7641 ( .A(n5457), .B(key[600]), .Z(n5459) );
  XNOR U7642 ( .A(\w3[3][80] ), .B(\w3[3][81] ), .Z(n5458) );
  XNOR U7643 ( .A(n5459), .B(n5458), .Z(n5460) );
  XOR U7644 ( .A(\w3[3][89] ), .B(n5460), .Z(\w1[4][88] ) );
  XOR U7645 ( .A(\w3[3][82] ), .B(key[601]), .Z(n5463) );
  XNOR U7646 ( .A(n5461), .B(\w3[3][90] ), .Z(n5462) );
  XNOR U7647 ( .A(n5463), .B(n5462), .Z(n5464) );
  XOR U7648 ( .A(\w3[3][65] ), .B(n5464), .Z(\w1[4][89] ) );
  XOR U7649 ( .A(\w3[3][9] ), .B(key[520]), .Z(n5466) );
  XNOR U7650 ( .A(\w3[3][1] ), .B(\w3[3][0] ), .Z(n5465) );
  XNOR U7651 ( .A(n5466), .B(n5465), .Z(n5467) );
  XOR U7652 ( .A(n5468), .B(n5467), .Z(\w1[4][8] ) );
  XOR U7653 ( .A(\w3[3][83] ), .B(key[602]), .Z(n5471) );
  XNOR U7654 ( .A(n5469), .B(\w3[3][91] ), .Z(n5470) );
  XNOR U7655 ( .A(n5471), .B(n5470), .Z(n5472) );
  XOR U7656 ( .A(\w3[3][66] ), .B(n5472), .Z(\w1[4][90] ) );
  XOR U7657 ( .A(n5473), .B(key[603]), .Z(n5476) );
  XNOR U7658 ( .A(\w3[3][67] ), .B(n5474), .Z(n5475) );
  XNOR U7659 ( .A(n5476), .B(n5475), .Z(\w1[4][91] ) );
  XOR U7660 ( .A(n5477), .B(key[604]), .Z(n5480) );
  XNOR U7661 ( .A(\w3[3][68] ), .B(n5478), .Z(n5479) );
  XNOR U7662 ( .A(n5480), .B(n5479), .Z(\w1[4][92] ) );
  XOR U7663 ( .A(\w3[3][86] ), .B(key[605]), .Z(n5483) );
  XNOR U7664 ( .A(n5481), .B(\w3[3][94] ), .Z(n5482) );
  XNOR U7665 ( .A(n5483), .B(n5482), .Z(n5484) );
  XOR U7666 ( .A(\w3[3][69] ), .B(n5484), .Z(\w1[4][93] ) );
  XOR U7667 ( .A(n5485), .B(key[606]), .Z(n5488) );
  XNOR U7668 ( .A(\w3[3][70] ), .B(n5486), .Z(n5487) );
  XNOR U7669 ( .A(n5488), .B(n5487), .Z(\w1[4][94] ) );
  XOR U7670 ( .A(n5489), .B(key[607]), .Z(n5492) );
  XNOR U7671 ( .A(n5490), .B(\w3[3][71] ), .Z(n5491) );
  XNOR U7672 ( .A(n5492), .B(n5491), .Z(\w1[4][95] ) );
  XOR U7673 ( .A(\w3[3][104] ), .B(key[608]), .Z(n5496) );
  XNOR U7674 ( .A(n5494), .B(n5493), .Z(n5495) );
  XNOR U7675 ( .A(n5496), .B(n5495), .Z(\w1[4][96] ) );
  XOR U7676 ( .A(n5497), .B(key[609]), .Z(n5500) );
  XNOR U7677 ( .A(\w3[3][121] ), .B(n5498), .Z(n5499) );
  XNOR U7678 ( .A(n5500), .B(n5499), .Z(\w1[4][97] ) );
  XOR U7679 ( .A(n5501), .B(key[610]), .Z(n5504) );
  XNOR U7680 ( .A(\w3[3][122] ), .B(n5502), .Z(n5503) );
  XNOR U7681 ( .A(n5504), .B(n5503), .Z(\w1[4][98] ) );
  XOR U7682 ( .A(n5505), .B(key[611]), .Z(n5508) );
  XNOR U7683 ( .A(n5506), .B(\w3[3][123] ), .Z(n5507) );
  XNOR U7684 ( .A(n5508), .B(n5507), .Z(\w1[4][99] ) );
  XOR U7685 ( .A(\w3[3][10] ), .B(key[521]), .Z(n5510) );
  XNOR U7686 ( .A(\w3[3][2] ), .B(\w3[3][17] ), .Z(n5509) );
  XNOR U7687 ( .A(n5510), .B(n5509), .Z(n5511) );
  XOR U7688 ( .A(n5512), .B(n5511), .Z(\w1[4][9] ) );
  XOR U7689 ( .A(\w3[4][8] ), .B(key[640]), .Z(n5514) );
  XOR U7690 ( .A(\w3[4][1] ), .B(\w3[4][25] ), .Z(n5936) );
  XOR U7691 ( .A(\w3[4][16] ), .B(\w3[4][24] ), .Z(n5892) );
  XNOR U7692 ( .A(n5936), .B(n5892), .Z(n5513) );
  XNOR U7693 ( .A(n5514), .B(n5513), .Z(\w1[5][0] ) );
  XOR U7694 ( .A(\w3[4][96] ), .B(\w3[4][101] ), .Z(n5540) );
  XOR U7695 ( .A(n5540), .B(key[740]), .Z(n5518) );
  XOR U7696 ( .A(\w3[4][116] ), .B(\w3[4][125] ), .Z(n5516) );
  XNOR U7697 ( .A(\w3[4][120] ), .B(\w3[4][108] ), .Z(n5515) );
  XNOR U7698 ( .A(n5516), .B(n5515), .Z(n5597) );
  XNOR U7699 ( .A(\w3[4][124] ), .B(n5597), .Z(n5517) );
  XNOR U7700 ( .A(n5518), .B(n5517), .Z(\w1[5][100] ) );
  XOR U7701 ( .A(\w3[4][102] ), .B(\w3[4][126] ), .Z(n5549) );
  XOR U7702 ( .A(n5549), .B(key[741]), .Z(n5520) );
  XOR U7703 ( .A(\w3[4][109] ), .B(\w3[4][117] ), .Z(n5600) );
  XNOR U7704 ( .A(\w3[4][125] ), .B(n5600), .Z(n5519) );
  XNOR U7705 ( .A(n5520), .B(n5519), .Z(\w1[5][101] ) );
  XOR U7706 ( .A(\w3[4][96] ), .B(\w3[4][103] ), .Z(n5550) );
  XOR U7707 ( .A(n5550), .B(key[742]), .Z(n5522) );
  XOR U7708 ( .A(\w3[4][110] ), .B(\w3[4][118] ), .Z(n5568) );
  XNOR U7709 ( .A(\w3[4][120] ), .B(\w3[4][127] ), .Z(n5524) );
  XNOR U7710 ( .A(n5568), .B(n5524), .Z(n5605) );
  XNOR U7711 ( .A(\w3[4][126] ), .B(n5605), .Z(n5521) );
  XNOR U7712 ( .A(n5522), .B(n5521), .Z(\w1[5][102] ) );
  XOR U7713 ( .A(\w3[4][111] ), .B(\w3[4][119] ), .Z(n5608) );
  XNOR U7714 ( .A(n5608), .B(key[743]), .Z(n5523) );
  XNOR U7715 ( .A(n5524), .B(n5523), .Z(n5525) );
  XNOR U7716 ( .A(\w3[4][96] ), .B(n5525), .Z(\w1[5][103] ) );
  XOR U7717 ( .A(key[744]), .B(\w3[4][105] ), .Z(n5527) );
  XNOR U7718 ( .A(\w3[4][96] ), .B(\w3[4][97] ), .Z(n5526) );
  XNOR U7719 ( .A(n5527), .B(n5526), .Z(n5528) );
  XNOR U7720 ( .A(\w3[4][120] ), .B(\w3[4][112] ), .Z(n5918) );
  XNOR U7721 ( .A(n5528), .B(n5918), .Z(\w1[5][104] ) );
  XOR U7722 ( .A(\w3[4][106] ), .B(\w3[4][98] ), .Z(n5530) );
  XOR U7723 ( .A(\w3[4][97] ), .B(\w3[4][121] ), .Z(n5917) );
  XNOR U7724 ( .A(n5917), .B(key[745]), .Z(n5529) );
  XNOR U7725 ( .A(n5530), .B(n5529), .Z(n5531) );
  XOR U7726 ( .A(\w3[4][113] ), .B(n5531), .Z(\w1[5][105] ) );
  XOR U7727 ( .A(\w3[4][107] ), .B(\w3[4][99] ), .Z(n5533) );
  XOR U7728 ( .A(\w3[4][98] ), .B(\w3[4][122] ), .Z(n5922) );
  XNOR U7729 ( .A(n5922), .B(key[746]), .Z(n5532) );
  XNOR U7730 ( .A(n5533), .B(n5532), .Z(n5534) );
  XOR U7731 ( .A(\w3[4][114] ), .B(n5534), .Z(\w1[5][106] ) );
  XOR U7732 ( .A(\w3[4][99] ), .B(\w3[4][123] ), .Z(n5926) );
  XNOR U7733 ( .A(\w3[4][108] ), .B(n5926), .Z(n5535) );
  XNOR U7734 ( .A(\w3[4][104] ), .B(n5535), .Z(n5561) );
  XOR U7735 ( .A(n5561), .B(key[747]), .Z(n5537) );
  XOR U7736 ( .A(\w3[4][96] ), .B(\w3[4][100] ), .Z(n5930) );
  XNOR U7737 ( .A(\w3[4][115] ), .B(n5930), .Z(n5536) );
  XNOR U7738 ( .A(n5537), .B(n5536), .Z(\w1[5][107] ) );
  XOR U7739 ( .A(\w3[4][100] ), .B(\w3[4][104] ), .Z(n5539) );
  XNOR U7740 ( .A(\w3[4][124] ), .B(\w3[4][109] ), .Z(n5538) );
  XNOR U7741 ( .A(n5539), .B(n5538), .Z(n5564) );
  XOR U7742 ( .A(n5564), .B(key[748]), .Z(n5542) );
  XNOR U7743 ( .A(\w3[4][116] ), .B(n5540), .Z(n5541) );
  XNOR U7744 ( .A(n5542), .B(n5541), .Z(\w1[5][108] ) );
  XOR U7745 ( .A(\w3[4][125] ), .B(\w3[4][101] ), .Z(n5567) );
  XOR U7746 ( .A(n5567), .B(key[749]), .Z(n5544) );
  XNOR U7747 ( .A(\w3[4][102] ), .B(\w3[4][110] ), .Z(n5543) );
  XNOR U7748 ( .A(n5544), .B(n5543), .Z(n5545) );
  XOR U7749 ( .A(\w3[4][117] ), .B(n5545), .Z(\w1[5][109] ) );
  XOR U7750 ( .A(\w3[4][11] ), .B(\w3[4][18] ), .Z(n5547) );
  XOR U7751 ( .A(\w3[4][2] ), .B(\w3[4][26] ), .Z(n5631) );
  XNOR U7752 ( .A(n5631), .B(key[650]), .Z(n5546) );
  XNOR U7753 ( .A(n5547), .B(n5546), .Z(n5548) );
  XOR U7754 ( .A(\w3[4][3] ), .B(n5548), .Z(\w1[5][10] ) );
  XNOR U7755 ( .A(\w3[4][111] ), .B(\w3[4][104] ), .Z(n5576) );
  XNOR U7756 ( .A(n5549), .B(n5576), .Z(n5571) );
  XOR U7757 ( .A(n5571), .B(key[750]), .Z(n5552) );
  XNOR U7758 ( .A(\w3[4][118] ), .B(n5550), .Z(n5551) );
  XNOR U7759 ( .A(n5552), .B(n5551), .Z(\w1[5][110] ) );
  XOR U7760 ( .A(\w3[4][127] ), .B(\w3[4][103] ), .Z(n5574) );
  XOR U7761 ( .A(n5574), .B(key[751]), .Z(n5554) );
  XOR U7762 ( .A(\w3[4][96] ), .B(\w3[4][104] ), .Z(n5581) );
  XNOR U7763 ( .A(\w3[4][119] ), .B(n5581), .Z(n5553) );
  XNOR U7764 ( .A(n5554), .B(n5553), .Z(\w1[5][111] ) );
  XOR U7765 ( .A(\w3[4][105] ), .B(\w3[4][113] ), .Z(n5921) );
  XOR U7766 ( .A(n5921), .B(key[752]), .Z(n5556) );
  XNOR U7767 ( .A(\w3[4][120] ), .B(n5581), .Z(n5555) );
  XNOR U7768 ( .A(n5556), .B(n5555), .Z(\w1[5][112] ) );
  XOR U7769 ( .A(\w3[4][106] ), .B(\w3[4][114] ), .Z(n5925) );
  XOR U7770 ( .A(n5925), .B(key[753]), .Z(n5558) );
  XNOR U7771 ( .A(\w3[4][105] ), .B(n5917), .Z(n5557) );
  XNOR U7772 ( .A(n5558), .B(n5557), .Z(\w1[5][113] ) );
  XOR U7773 ( .A(\w3[4][107] ), .B(\w3[4][115] ), .Z(n5592) );
  XOR U7774 ( .A(n5592), .B(key[754]), .Z(n5560) );
  XNOR U7775 ( .A(\w3[4][106] ), .B(n5922), .Z(n5559) );
  XNOR U7776 ( .A(n5560), .B(n5559), .Z(\w1[5][114] ) );
  XOR U7777 ( .A(\w3[4][116] ), .B(\w3[4][112] ), .Z(n5593) );
  XOR U7778 ( .A(n5593), .B(key[755]), .Z(n5563) );
  XNOR U7779 ( .A(\w3[4][107] ), .B(n5561), .Z(n5562) );
  XNOR U7780 ( .A(n5563), .B(n5562), .Z(\w1[5][115] ) );
  XOR U7781 ( .A(\w3[4][117] ), .B(\w3[4][112] ), .Z(n5596) );
  XOR U7782 ( .A(n5596), .B(key[756]), .Z(n5566) );
  XNOR U7783 ( .A(\w3[4][108] ), .B(n5564), .Z(n5565) );
  XNOR U7784 ( .A(n5566), .B(n5565), .Z(\w1[5][116] ) );
  XOR U7785 ( .A(n5567), .B(key[757]), .Z(n5570) );
  XNOR U7786 ( .A(\w3[4][109] ), .B(n5568), .Z(n5569) );
  XNOR U7787 ( .A(n5570), .B(n5569), .Z(\w1[5][117] ) );
  XOR U7788 ( .A(\w3[4][119] ), .B(\w3[4][112] ), .Z(n5604) );
  XOR U7789 ( .A(n5604), .B(key[758]), .Z(n5573) );
  XNOR U7790 ( .A(\w3[4][110] ), .B(n5571), .Z(n5572) );
  XNOR U7791 ( .A(n5573), .B(n5572), .Z(\w1[5][118] ) );
  XNOR U7792 ( .A(n5574), .B(key[759]), .Z(n5575) );
  XNOR U7793 ( .A(n5576), .B(n5575), .Z(n5577) );
  XNOR U7794 ( .A(\w3[4][112] ), .B(n5577), .Z(\w1[5][119] ) );
  XOR U7795 ( .A(\w3[4][3] ), .B(\w3[4][27] ), .Z(n5672) );
  XNOR U7796 ( .A(\w3[4][8] ), .B(\w3[4][12] ), .Z(n5578) );
  XNOR U7797 ( .A(n5672), .B(n5578), .Z(n5628) );
  XOR U7798 ( .A(n5628), .B(key[651]), .Z(n5580) );
  XOR U7799 ( .A(\w3[4][0] ), .B(\w3[4][4] ), .Z(n5702) );
  XNOR U7800 ( .A(\w3[4][19] ), .B(n5702), .Z(n5579) );
  XNOR U7801 ( .A(n5580), .B(n5579), .Z(\w1[5][11] ) );
  XOR U7802 ( .A(n5581), .B(key[760]), .Z(n5583) );
  XNOR U7803 ( .A(\w3[4][113] ), .B(\w3[4][121] ), .Z(n5582) );
  XNOR U7804 ( .A(n5583), .B(n5582), .Z(n5584) );
  XOR U7805 ( .A(\w3[4][112] ), .B(n5584), .Z(\w1[5][120] ) );
  XOR U7806 ( .A(n5921), .B(key[761]), .Z(n5586) );
  XNOR U7807 ( .A(\w3[4][114] ), .B(\w3[4][122] ), .Z(n5585) );
  XNOR U7808 ( .A(n5586), .B(n5585), .Z(n5587) );
  XOR U7809 ( .A(\w3[4][97] ), .B(n5587), .Z(\w1[5][121] ) );
  XOR U7810 ( .A(n5925), .B(key[762]), .Z(n5589) );
  XNOR U7811 ( .A(\w3[4][115] ), .B(\w3[4][123] ), .Z(n5588) );
  XNOR U7812 ( .A(n5589), .B(n5588), .Z(n5590) );
  XOR U7813 ( .A(\w3[4][98] ), .B(n5590), .Z(\w1[5][122] ) );
  XNOR U7814 ( .A(\w3[4][124] ), .B(\w3[4][120] ), .Z(n5591) );
  XNOR U7815 ( .A(n5592), .B(n5591), .Z(n5929) );
  XOR U7816 ( .A(n5929), .B(key[763]), .Z(n5595) );
  XNOR U7817 ( .A(\w3[4][99] ), .B(n5593), .Z(n5594) );
  XNOR U7818 ( .A(n5595), .B(n5594), .Z(\w1[5][123] ) );
  XOR U7819 ( .A(n5596), .B(key[764]), .Z(n5599) );
  XNOR U7820 ( .A(n5597), .B(\w3[4][100] ), .Z(n5598) );
  XNOR U7821 ( .A(n5599), .B(n5598), .Z(\w1[5][124] ) );
  XOR U7822 ( .A(\w3[4][118] ), .B(key[765]), .Z(n5602) );
  XNOR U7823 ( .A(n5600), .B(\w3[4][126] ), .Z(n5601) );
  XNOR U7824 ( .A(n5602), .B(n5601), .Z(n5603) );
  XOR U7825 ( .A(\w3[4][101] ), .B(n5603), .Z(\w1[5][125] ) );
  XOR U7826 ( .A(n5604), .B(key[766]), .Z(n5607) );
  XNOR U7827 ( .A(\w3[4][102] ), .B(n5605), .Z(n5606) );
  XNOR U7828 ( .A(n5607), .B(n5606), .Z(\w1[5][126] ) );
  XNOR U7829 ( .A(n5608), .B(key[767]), .Z(n5609) );
  XNOR U7830 ( .A(n5918), .B(n5609), .Z(n5610) );
  XNOR U7831 ( .A(\w3[4][103] ), .B(n5610), .Z(\w1[5][127] ) );
  XOR U7832 ( .A(\w3[4][13] ), .B(\w3[4][28] ), .Z(n5612) );
  XNOR U7833 ( .A(\w3[4][8] ), .B(\w3[4][4] ), .Z(n5611) );
  XNOR U7834 ( .A(n5612), .B(n5611), .Z(n5634) );
  XOR U7835 ( .A(n5634), .B(key[652]), .Z(n5614) );
  XOR U7836 ( .A(\w3[4][0] ), .B(\w3[4][5] ), .Z(n5739) );
  XNOR U7837 ( .A(\w3[4][20] ), .B(n5739), .Z(n5613) );
  XNOR U7838 ( .A(n5614), .B(n5613), .Z(\w1[5][12] ) );
  XOR U7839 ( .A(\w3[4][14] ), .B(\w3[4][6] ), .Z(n5616) );
  XOR U7840 ( .A(\w3[4][5] ), .B(\w3[4][29] ), .Z(n5637) );
  XNOR U7841 ( .A(n5637), .B(key[653]), .Z(n5615) );
  XNOR U7842 ( .A(n5616), .B(n5615), .Z(n5617) );
  XOR U7843 ( .A(\w3[4][21] ), .B(n5617), .Z(\w1[5][13] ) );
  XOR U7844 ( .A(\w3[4][6] ), .B(\w3[4][30] ), .Z(n5780) );
  XNOR U7845 ( .A(\w3[4][8] ), .B(\w3[4][15] ), .Z(n5645) );
  XNOR U7846 ( .A(n5780), .B(n5645), .Z(n5640) );
  XOR U7847 ( .A(n5640), .B(key[654]), .Z(n5619) );
  XOR U7848 ( .A(\w3[4][0] ), .B(\w3[4][7] ), .Z(n5815) );
  XNOR U7849 ( .A(\w3[4][22] ), .B(n5815), .Z(n5618) );
  XNOR U7850 ( .A(n5619), .B(n5618), .Z(\w1[5][14] ) );
  XOR U7851 ( .A(\w3[4][7] ), .B(\w3[4][31] ), .Z(n5643) );
  XOR U7852 ( .A(n5643), .B(key[655]), .Z(n5621) );
  XOR U7853 ( .A(\w3[4][8] ), .B(\w3[4][0] ), .Z(n5647) );
  XNOR U7854 ( .A(\w3[4][23] ), .B(n5647), .Z(n5620) );
  XNOR U7855 ( .A(n5621), .B(n5620), .Z(\w1[5][15] ) );
  XOR U7856 ( .A(\w3[4][17] ), .B(\w3[4][9] ), .Z(n5651) );
  XOR U7857 ( .A(n5651), .B(key[656]), .Z(n5623) );
  XNOR U7858 ( .A(\w3[4][24] ), .B(n5647), .Z(n5622) );
  XNOR U7859 ( .A(n5623), .B(n5622), .Z(\w1[5][16] ) );
  XOR U7860 ( .A(\w3[4][18] ), .B(\w3[4][10] ), .Z(n5671) );
  XOR U7861 ( .A(n5671), .B(key[657]), .Z(n5625) );
  XNOR U7862 ( .A(n5936), .B(\w3[4][9] ), .Z(n5624) );
  XNOR U7863 ( .A(n5625), .B(n5624), .Z(\w1[5][17] ) );
  XOR U7864 ( .A(\w3[4][11] ), .B(\w3[4][19] ), .Z(n5659) );
  XOR U7865 ( .A(n5659), .B(key[658]), .Z(n5627) );
  XNOR U7866 ( .A(n5631), .B(\w3[4][10] ), .Z(n5626) );
  XNOR U7867 ( .A(n5627), .B(n5626), .Z(\w1[5][18] ) );
  XOR U7868 ( .A(\w3[4][16] ), .B(\w3[4][20] ), .Z(n5660) );
  XOR U7869 ( .A(n5660), .B(key[659]), .Z(n5630) );
  XNOR U7870 ( .A(\w3[4][11] ), .B(n5628), .Z(n5629) );
  XNOR U7871 ( .A(n5630), .B(n5629), .Z(\w1[5][19] ) );
  XOR U7872 ( .A(n5651), .B(key[641]), .Z(n5633) );
  XNOR U7873 ( .A(\w3[4][25] ), .B(n5631), .Z(n5632) );
  XNOR U7874 ( .A(n5633), .B(n5632), .Z(\w1[5][1] ) );
  XOR U7875 ( .A(\w3[4][16] ), .B(\w3[4][21] ), .Z(n5665) );
  XOR U7876 ( .A(n5665), .B(key[660]), .Z(n5636) );
  XNOR U7877 ( .A(\w3[4][12] ), .B(n5634), .Z(n5635) );
  XNOR U7878 ( .A(n5636), .B(n5635), .Z(\w1[5][20] ) );
  XOR U7879 ( .A(\w3[4][14] ), .B(\w3[4][22] ), .Z(n5675) );
  XOR U7880 ( .A(n5675), .B(key[661]), .Z(n5639) );
  XNOR U7881 ( .A(\w3[4][13] ), .B(n5637), .Z(n5638) );
  XNOR U7882 ( .A(n5639), .B(n5638), .Z(\w1[5][21] ) );
  XOR U7883 ( .A(\w3[4][16] ), .B(\w3[4][23] ), .Z(n5676) );
  XOR U7884 ( .A(n5676), .B(key[662]), .Z(n5642) );
  XNOR U7885 ( .A(\w3[4][14] ), .B(n5640), .Z(n5641) );
  XNOR U7886 ( .A(n5642), .B(n5641), .Z(\w1[5][22] ) );
  XNOR U7887 ( .A(n5643), .B(key[663]), .Z(n5644) );
  XNOR U7888 ( .A(n5645), .B(n5644), .Z(n5646) );
  XNOR U7889 ( .A(\w3[4][16] ), .B(n5646), .Z(\w1[5][23] ) );
  XOR U7890 ( .A(\w3[4][17] ), .B(key[664]), .Z(n5649) );
  XNOR U7891 ( .A(\w3[4][25] ), .B(n5647), .Z(n5648) );
  XNOR U7892 ( .A(n5649), .B(n5648), .Z(n5650) );
  XOR U7893 ( .A(\w3[4][16] ), .B(n5650), .Z(\w1[5][24] ) );
  XOR U7894 ( .A(n5651), .B(key[665]), .Z(n5653) );
  XNOR U7895 ( .A(\w3[4][1] ), .B(\w3[4][26] ), .Z(n5652) );
  XNOR U7896 ( .A(n5653), .B(n5652), .Z(n5654) );
  XOR U7897 ( .A(\w3[4][18] ), .B(n5654), .Z(\w1[5][25] ) );
  XOR U7898 ( .A(n5671), .B(key[666]), .Z(n5656) );
  XNOR U7899 ( .A(\w3[4][2] ), .B(\w3[4][19] ), .Z(n5655) );
  XNOR U7900 ( .A(n5656), .B(n5655), .Z(n5657) );
  XOR U7901 ( .A(\w3[4][27] ), .B(n5657), .Z(\w1[5][26] ) );
  XNOR U7902 ( .A(\w3[4][24] ), .B(\w3[4][28] ), .Z(n5658) );
  XNOR U7903 ( .A(n5659), .B(n5658), .Z(n5701) );
  XOR U7904 ( .A(n5701), .B(key[667]), .Z(n5662) );
  XNOR U7905 ( .A(\w3[4][3] ), .B(n5660), .Z(n5661) );
  XNOR U7906 ( .A(n5662), .B(n5661), .Z(\w1[5][27] ) );
  XOR U7907 ( .A(\w3[4][20] ), .B(\w3[4][29] ), .Z(n5664) );
  XNOR U7908 ( .A(\w3[4][24] ), .B(\w3[4][12] ), .Z(n5663) );
  XNOR U7909 ( .A(n5664), .B(n5663), .Z(n5738) );
  XOR U7910 ( .A(n5738), .B(key[668]), .Z(n5667) );
  XNOR U7911 ( .A(\w3[4][4] ), .B(n5665), .Z(n5666) );
  XNOR U7912 ( .A(n5667), .B(n5666), .Z(\w1[5][28] ) );
  XOR U7913 ( .A(\w3[4][13] ), .B(\w3[4][21] ), .Z(n5779) );
  XOR U7914 ( .A(n5779), .B(key[669]), .Z(n5669) );
  XNOR U7915 ( .A(\w3[4][22] ), .B(\w3[4][30] ), .Z(n5668) );
  XNOR U7916 ( .A(n5669), .B(n5668), .Z(n5670) );
  XOR U7917 ( .A(\w3[4][5] ), .B(n5670), .Z(\w1[5][29] ) );
  XOR U7918 ( .A(n5671), .B(key[642]), .Z(n5674) );
  XNOR U7919 ( .A(\w3[4][26] ), .B(n5672), .Z(n5673) );
  XNOR U7920 ( .A(n5674), .B(n5673), .Z(\w1[5][2] ) );
  XNOR U7921 ( .A(\w3[4][24] ), .B(\w3[4][31] ), .Z(n5853) );
  XNOR U7922 ( .A(n5675), .B(n5853), .Z(n5814) );
  XOR U7923 ( .A(n5814), .B(key[670]), .Z(n5678) );
  XNOR U7924 ( .A(\w3[4][6] ), .B(n5676), .Z(n5677) );
  XNOR U7925 ( .A(n5678), .B(n5677), .Z(\w1[5][30] ) );
  XOR U7926 ( .A(\w3[4][15] ), .B(\w3[4][23] ), .Z(n5851) );
  XOR U7927 ( .A(n5851), .B(key[671]), .Z(n5680) );
  XNOR U7928 ( .A(n5892), .B(\w3[4][7] ), .Z(n5679) );
  XNOR U7929 ( .A(n5680), .B(n5679), .Z(\w1[5][31] ) );
  XOR U7930 ( .A(\w3[4][33] ), .B(\w3[4][57] ), .Z(n5735) );
  XOR U7931 ( .A(n5735), .B(key[672]), .Z(n5682) );
  XOR U7932 ( .A(\w3[4][48] ), .B(\w3[4][56] ), .Z(n5796) );
  XNOR U7933 ( .A(n5796), .B(\w3[4][40] ), .Z(n5681) );
  XNOR U7934 ( .A(n5682), .B(n5681), .Z(\w1[5][32] ) );
  XOR U7935 ( .A(\w3[4][34] ), .B(\w3[4][58] ), .Z(n5743) );
  XOR U7936 ( .A(n5743), .B(key[673]), .Z(n5684) );
  XOR U7937 ( .A(\w3[4][41] ), .B(\w3[4][49] ), .Z(n5767) );
  XNOR U7938 ( .A(\w3[4][57] ), .B(n5767), .Z(n5683) );
  XNOR U7939 ( .A(n5684), .B(n5683), .Z(\w1[5][33] ) );
  XOR U7940 ( .A(\w3[4][35] ), .B(\w3[4][59] ), .Z(n5714) );
  XOR U7941 ( .A(n5714), .B(key[674]), .Z(n5686) );
  XOR U7942 ( .A(\w3[4][42] ), .B(\w3[4][50] ), .Z(n5771) );
  XNOR U7943 ( .A(\w3[4][58] ), .B(n5771), .Z(n5685) );
  XNOR U7944 ( .A(n5686), .B(n5685), .Z(\w1[5][34] ) );
  XOR U7945 ( .A(\w3[4][36] ), .B(\w3[4][32] ), .Z(n5716) );
  XOR U7946 ( .A(n5716), .B(key[675]), .Z(n5689) );
  XOR U7947 ( .A(\w3[4][43] ), .B(\w3[4][51] ), .Z(n5742) );
  XNOR U7948 ( .A(\w3[4][56] ), .B(n5742), .Z(n5687) );
  XNOR U7949 ( .A(\w3[4][60] ), .B(n5687), .Z(n5776) );
  XNOR U7950 ( .A(\w3[4][59] ), .B(n5776), .Z(n5688) );
  XNOR U7951 ( .A(n5689), .B(n5688), .Z(\w1[5][35] ) );
  XOR U7952 ( .A(\w3[4][32] ), .B(\w3[4][37] ), .Z(n5721) );
  XOR U7953 ( .A(n5721), .B(key[676]), .Z(n5693) );
  XOR U7954 ( .A(\w3[4][52] ), .B(\w3[4][61] ), .Z(n5691) );
  XNOR U7955 ( .A(\w3[4][56] ), .B(\w3[4][44] ), .Z(n5690) );
  XNOR U7956 ( .A(n5691), .B(n5690), .Z(n5784) );
  XNOR U7957 ( .A(\w3[4][60] ), .B(n5784), .Z(n5692) );
  XNOR U7958 ( .A(n5693), .B(n5692), .Z(\w1[5][36] ) );
  XOR U7959 ( .A(\w3[4][38] ), .B(\w3[4][62] ), .Z(n5727) );
  XOR U7960 ( .A(n5727), .B(key[677]), .Z(n5695) );
  XOR U7961 ( .A(\w3[4][45] ), .B(\w3[4][53] ), .Z(n5787) );
  XNOR U7962 ( .A(\w3[4][61] ), .B(n5787), .Z(n5694) );
  XNOR U7963 ( .A(n5695), .B(n5694), .Z(\w1[5][37] ) );
  XOR U7964 ( .A(\w3[4][32] ), .B(\w3[4][39] ), .Z(n5728) );
  XOR U7965 ( .A(n5728), .B(key[678]), .Z(n5697) );
  XOR U7966 ( .A(\w3[4][46] ), .B(\w3[4][54] ), .Z(n5753) );
  XNOR U7967 ( .A(\w3[4][56] ), .B(\w3[4][63] ), .Z(n5699) );
  XNOR U7968 ( .A(n5753), .B(n5699), .Z(n5792) );
  XNOR U7969 ( .A(\w3[4][62] ), .B(n5792), .Z(n5696) );
  XNOR U7970 ( .A(n5697), .B(n5696), .Z(\w1[5][38] ) );
  XOR U7971 ( .A(\w3[4][47] ), .B(\w3[4][55] ), .Z(n5795) );
  XNOR U7972 ( .A(n5795), .B(key[679]), .Z(n5698) );
  XNOR U7973 ( .A(n5699), .B(n5698), .Z(n5700) );
  XNOR U7974 ( .A(\w3[4][32] ), .B(n5700), .Z(\w1[5][39] ) );
  XOR U7975 ( .A(n5701), .B(key[643]), .Z(n5704) );
  XNOR U7976 ( .A(n5702), .B(\w3[4][27] ), .Z(n5703) );
  XNOR U7977 ( .A(n5704), .B(n5703), .Z(\w1[5][3] ) );
  XOR U7978 ( .A(\w3[4][32] ), .B(key[680]), .Z(n5706) );
  XNOR U7979 ( .A(\w3[4][33] ), .B(\w3[4][41] ), .Z(n5705) );
  XNOR U7980 ( .A(n5706), .B(n5705), .Z(n5707) );
  XOR U7981 ( .A(n5796), .B(n5707), .Z(\w1[5][40] ) );
  XOR U7982 ( .A(\w3[4][42] ), .B(key[681]), .Z(n5709) );
  XNOR U7983 ( .A(\w3[4][49] ), .B(\w3[4][34] ), .Z(n5708) );
  XNOR U7984 ( .A(n5709), .B(n5708), .Z(n5710) );
  XOR U7985 ( .A(n5735), .B(n5710), .Z(\w1[5][41] ) );
  XOR U7986 ( .A(\w3[4][43] ), .B(key[682]), .Z(n5712) );
  XNOR U7987 ( .A(\w3[4][50] ), .B(\w3[4][35] ), .Z(n5711) );
  XNOR U7988 ( .A(n5712), .B(n5711), .Z(n5713) );
  XOR U7989 ( .A(n5743), .B(n5713), .Z(\w1[5][42] ) );
  XNOR U7990 ( .A(\w3[4][40] ), .B(n5714), .Z(n5715) );
  XNOR U7991 ( .A(\w3[4][44] ), .B(n5715), .Z(n5746) );
  XOR U7992 ( .A(n5746), .B(key[683]), .Z(n5718) );
  XNOR U7993 ( .A(\w3[4][51] ), .B(n5716), .Z(n5717) );
  XNOR U7994 ( .A(n5718), .B(n5717), .Z(\w1[5][43] ) );
  XOR U7995 ( .A(\w3[4][36] ), .B(\w3[4][45] ), .Z(n5720) );
  XNOR U7996 ( .A(\w3[4][40] ), .B(\w3[4][60] ), .Z(n5719) );
  XNOR U7997 ( .A(n5720), .B(n5719), .Z(n5749) );
  XOR U7998 ( .A(n5749), .B(key[684]), .Z(n5723) );
  XNOR U7999 ( .A(\w3[4][52] ), .B(n5721), .Z(n5722) );
  XNOR U8000 ( .A(n5723), .B(n5722), .Z(\w1[5][44] ) );
  XOR U8001 ( .A(\w3[4][61] ), .B(\w3[4][37] ), .Z(n5752) );
  XOR U8002 ( .A(n5752), .B(key[685]), .Z(n5725) );
  XNOR U8003 ( .A(\w3[4][38] ), .B(\w3[4][46] ), .Z(n5724) );
  XNOR U8004 ( .A(n5725), .B(n5724), .Z(n5726) );
  XOR U8005 ( .A(\w3[4][53] ), .B(n5726), .Z(\w1[5][45] ) );
  XNOR U8006 ( .A(\w3[4][40] ), .B(\w3[4][47] ), .Z(n5761) );
  XNOR U8007 ( .A(n5727), .B(n5761), .Z(n5756) );
  XOR U8008 ( .A(n5756), .B(key[686]), .Z(n5730) );
  XNOR U8009 ( .A(\w3[4][54] ), .B(n5728), .Z(n5729) );
  XNOR U8010 ( .A(n5730), .B(n5729), .Z(\w1[5][46] ) );
  XOR U8011 ( .A(\w3[4][63] ), .B(\w3[4][39] ), .Z(n5759) );
  XOR U8012 ( .A(n5759), .B(key[687]), .Z(n5732) );
  XOR U8013 ( .A(\w3[4][40] ), .B(\w3[4][32] ), .Z(n5763) );
  XNOR U8014 ( .A(\w3[4][55] ), .B(n5763), .Z(n5731) );
  XNOR U8015 ( .A(n5732), .B(n5731), .Z(\w1[5][47] ) );
  XOR U8016 ( .A(n5763), .B(key[688]), .Z(n5734) );
  XNOR U8017 ( .A(\w3[4][56] ), .B(n5767), .Z(n5733) );
  XNOR U8018 ( .A(n5734), .B(n5733), .Z(\w1[5][48] ) );
  XOR U8019 ( .A(n5771), .B(key[689]), .Z(n5737) );
  XNOR U8020 ( .A(n5735), .B(\w3[4][41] ), .Z(n5736) );
  XNOR U8021 ( .A(n5737), .B(n5736), .Z(\w1[5][49] ) );
  XOR U8022 ( .A(n5738), .B(key[644]), .Z(n5741) );
  XNOR U8023 ( .A(n5739), .B(\w3[4][28] ), .Z(n5740) );
  XNOR U8024 ( .A(n5741), .B(n5740), .Z(\w1[5][4] ) );
  XOR U8025 ( .A(n5742), .B(key[690]), .Z(n5745) );
  XNOR U8026 ( .A(n5743), .B(\w3[4][42] ), .Z(n5744) );
  XNOR U8027 ( .A(n5745), .B(n5744), .Z(\w1[5][50] ) );
  XOR U8028 ( .A(\w3[4][48] ), .B(\w3[4][52] ), .Z(n5775) );
  XOR U8029 ( .A(n5775), .B(key[691]), .Z(n5748) );
  XNOR U8030 ( .A(\w3[4][43] ), .B(n5746), .Z(n5747) );
  XNOR U8031 ( .A(n5748), .B(n5747), .Z(\w1[5][51] ) );
  XOR U8032 ( .A(\w3[4][48] ), .B(\w3[4][53] ), .Z(n5783) );
  XOR U8033 ( .A(n5783), .B(key[692]), .Z(n5751) );
  XNOR U8034 ( .A(\w3[4][44] ), .B(n5749), .Z(n5750) );
  XNOR U8035 ( .A(n5751), .B(n5750), .Z(\w1[5][52] ) );
  XOR U8036 ( .A(n5752), .B(key[693]), .Z(n5755) );
  XNOR U8037 ( .A(\w3[4][45] ), .B(n5753), .Z(n5754) );
  XNOR U8038 ( .A(n5755), .B(n5754), .Z(\w1[5][53] ) );
  XOR U8039 ( .A(\w3[4][48] ), .B(\w3[4][55] ), .Z(n5791) );
  XOR U8040 ( .A(n5791), .B(key[694]), .Z(n5758) );
  XNOR U8041 ( .A(\w3[4][46] ), .B(n5756), .Z(n5757) );
  XNOR U8042 ( .A(n5758), .B(n5757), .Z(\w1[5][54] ) );
  XNOR U8043 ( .A(n5759), .B(key[695]), .Z(n5760) );
  XNOR U8044 ( .A(n5761), .B(n5760), .Z(n5762) );
  XNOR U8045 ( .A(\w3[4][48] ), .B(n5762), .Z(\w1[5][55] ) );
  XOR U8046 ( .A(n5763), .B(key[696]), .Z(n5765) );
  XNOR U8047 ( .A(\w3[4][48] ), .B(\w3[4][49] ), .Z(n5764) );
  XNOR U8048 ( .A(n5765), .B(n5764), .Z(n5766) );
  XOR U8049 ( .A(\w3[4][57] ), .B(n5766), .Z(\w1[5][56] ) );
  XOR U8050 ( .A(\w3[4][50] ), .B(key[697]), .Z(n5769) );
  XNOR U8051 ( .A(n5767), .B(\w3[4][58] ), .Z(n5768) );
  XNOR U8052 ( .A(n5769), .B(n5768), .Z(n5770) );
  XOR U8053 ( .A(\w3[4][33] ), .B(n5770), .Z(\w1[5][57] ) );
  XOR U8054 ( .A(\w3[4][51] ), .B(key[698]), .Z(n5773) );
  XNOR U8055 ( .A(n5771), .B(\w3[4][59] ), .Z(n5772) );
  XNOR U8056 ( .A(n5773), .B(n5772), .Z(n5774) );
  XOR U8057 ( .A(\w3[4][34] ), .B(n5774), .Z(\w1[5][58] ) );
  XOR U8058 ( .A(n5775), .B(key[699]), .Z(n5778) );
  XNOR U8059 ( .A(\w3[4][35] ), .B(n5776), .Z(n5777) );
  XNOR U8060 ( .A(n5778), .B(n5777), .Z(\w1[5][59] ) );
  XOR U8061 ( .A(n5779), .B(key[645]), .Z(n5782) );
  XNOR U8062 ( .A(\w3[4][29] ), .B(n5780), .Z(n5781) );
  XNOR U8063 ( .A(n5782), .B(n5781), .Z(\w1[5][5] ) );
  XOR U8064 ( .A(n5783), .B(key[700]), .Z(n5786) );
  XNOR U8065 ( .A(\w3[4][36] ), .B(n5784), .Z(n5785) );
  XNOR U8066 ( .A(n5786), .B(n5785), .Z(\w1[5][60] ) );
  XOR U8067 ( .A(\w3[4][54] ), .B(key[701]), .Z(n5789) );
  XNOR U8068 ( .A(n5787), .B(\w3[4][62] ), .Z(n5788) );
  XNOR U8069 ( .A(n5789), .B(n5788), .Z(n5790) );
  XOR U8070 ( .A(\w3[4][37] ), .B(n5790), .Z(\w1[5][61] ) );
  XOR U8071 ( .A(n5791), .B(key[702]), .Z(n5794) );
  XNOR U8072 ( .A(\w3[4][38] ), .B(n5792), .Z(n5793) );
  XNOR U8073 ( .A(n5794), .B(n5793), .Z(\w1[5][62] ) );
  XOR U8074 ( .A(n5795), .B(key[703]), .Z(n5798) );
  XNOR U8075 ( .A(n5796), .B(\w3[4][39] ), .Z(n5797) );
  XNOR U8076 ( .A(n5798), .B(n5797), .Z(\w1[5][63] ) );
  XOR U8077 ( .A(\w3[4][65] ), .B(\w3[4][89] ), .Z(n5857) );
  XOR U8078 ( .A(n5857), .B(key[704]), .Z(n5800) );
  XOR U8079 ( .A(\w3[4][80] ), .B(\w3[4][88] ), .Z(n5914) );
  XNOR U8080 ( .A(n5914), .B(\w3[4][72] ), .Z(n5799) );
  XNOR U8081 ( .A(n5800), .B(n5799), .Z(\w1[5][64] ) );
  XOR U8082 ( .A(\w3[4][66] ), .B(\w3[4][90] ), .Z(n5861) );
  XOR U8083 ( .A(n5861), .B(key[705]), .Z(n5802) );
  XOR U8084 ( .A(\w3[4][73] ), .B(\w3[4][81] ), .Z(n5885) );
  XNOR U8085 ( .A(\w3[4][89] ), .B(n5885), .Z(n5801) );
  XNOR U8086 ( .A(n5802), .B(n5801), .Z(\w1[5][65] ) );
  XOR U8087 ( .A(\w3[4][67] ), .B(\w3[4][91] ), .Z(n5832) );
  XOR U8088 ( .A(n5832), .B(key[706]), .Z(n5804) );
  XOR U8089 ( .A(\w3[4][74] ), .B(\w3[4][82] ), .Z(n5893) );
  XNOR U8090 ( .A(\w3[4][90] ), .B(n5893), .Z(n5803) );
  XNOR U8091 ( .A(n5804), .B(n5803), .Z(\w1[5][66] ) );
  XOR U8092 ( .A(\w3[4][68] ), .B(\w3[4][64] ), .Z(n5834) );
  XOR U8093 ( .A(n5834), .B(key[707]), .Z(n5807) );
  XOR U8094 ( .A(\w3[4][75] ), .B(\w3[4][83] ), .Z(n5860) );
  XNOR U8095 ( .A(\w3[4][88] ), .B(n5860), .Z(n5805) );
  XNOR U8096 ( .A(\w3[4][92] ), .B(n5805), .Z(n5898) );
  XNOR U8097 ( .A(\w3[4][91] ), .B(n5898), .Z(n5806) );
  XNOR U8098 ( .A(n5807), .B(n5806), .Z(\w1[5][67] ) );
  XOR U8099 ( .A(\w3[4][64] ), .B(\w3[4][69] ), .Z(n5839) );
  XOR U8100 ( .A(n5839), .B(key[708]), .Z(n5811) );
  XOR U8101 ( .A(\w3[4][84] ), .B(\w3[4][93] ), .Z(n5809) );
  XNOR U8102 ( .A(\w3[4][88] ), .B(\w3[4][76] ), .Z(n5808) );
  XNOR U8103 ( .A(n5809), .B(n5808), .Z(n5902) );
  XNOR U8104 ( .A(\w3[4][92] ), .B(n5902), .Z(n5810) );
  XNOR U8105 ( .A(n5811), .B(n5810), .Z(\w1[5][68] ) );
  XOR U8106 ( .A(\w3[4][70] ), .B(\w3[4][94] ), .Z(n5845) );
  XOR U8107 ( .A(n5845), .B(key[709]), .Z(n5813) );
  XOR U8108 ( .A(\w3[4][77] ), .B(\w3[4][85] ), .Z(n5905) );
  XNOR U8109 ( .A(\w3[4][93] ), .B(n5905), .Z(n5812) );
  XNOR U8110 ( .A(n5813), .B(n5812), .Z(\w1[5][69] ) );
  XOR U8111 ( .A(n5814), .B(key[646]), .Z(n5817) );
  XNOR U8112 ( .A(n5815), .B(\w3[4][30] ), .Z(n5816) );
  XNOR U8113 ( .A(n5817), .B(n5816), .Z(\w1[5][6] ) );
  XOR U8114 ( .A(\w3[4][64] ), .B(\w3[4][71] ), .Z(n5846) );
  XOR U8115 ( .A(n5846), .B(key[710]), .Z(n5819) );
  XOR U8116 ( .A(\w3[4][78] ), .B(\w3[4][86] ), .Z(n5871) );
  XNOR U8117 ( .A(\w3[4][88] ), .B(\w3[4][95] ), .Z(n5821) );
  XNOR U8118 ( .A(n5871), .B(n5821), .Z(n5910) );
  XNOR U8119 ( .A(\w3[4][94] ), .B(n5910), .Z(n5818) );
  XNOR U8120 ( .A(n5819), .B(n5818), .Z(\w1[5][70] ) );
  XOR U8121 ( .A(\w3[4][79] ), .B(\w3[4][87] ), .Z(n5913) );
  XNOR U8122 ( .A(n5913), .B(key[711]), .Z(n5820) );
  XNOR U8123 ( .A(n5821), .B(n5820), .Z(n5822) );
  XNOR U8124 ( .A(\w3[4][64] ), .B(n5822), .Z(\w1[5][71] ) );
  XOR U8125 ( .A(\w3[4][64] ), .B(key[712]), .Z(n5824) );
  XNOR U8126 ( .A(\w3[4][65] ), .B(\w3[4][73] ), .Z(n5823) );
  XNOR U8127 ( .A(n5824), .B(n5823), .Z(n5825) );
  XOR U8128 ( .A(n5914), .B(n5825), .Z(\w1[5][72] ) );
  XOR U8129 ( .A(\w3[4][74] ), .B(key[713]), .Z(n5827) );
  XNOR U8130 ( .A(\w3[4][81] ), .B(\w3[4][66] ), .Z(n5826) );
  XNOR U8131 ( .A(n5827), .B(n5826), .Z(n5828) );
  XOR U8132 ( .A(n5857), .B(n5828), .Z(\w1[5][73] ) );
  XOR U8133 ( .A(\w3[4][75] ), .B(key[714]), .Z(n5830) );
  XNOR U8134 ( .A(\w3[4][82] ), .B(\w3[4][67] ), .Z(n5829) );
  XNOR U8135 ( .A(n5830), .B(n5829), .Z(n5831) );
  XOR U8136 ( .A(n5861), .B(n5831), .Z(\w1[5][74] ) );
  XNOR U8137 ( .A(\w3[4][72] ), .B(n5832), .Z(n5833) );
  XNOR U8138 ( .A(\w3[4][76] ), .B(n5833), .Z(n5864) );
  XOR U8139 ( .A(n5864), .B(key[715]), .Z(n5836) );
  XNOR U8140 ( .A(\w3[4][83] ), .B(n5834), .Z(n5835) );
  XNOR U8141 ( .A(n5836), .B(n5835), .Z(\w1[5][75] ) );
  XOR U8142 ( .A(\w3[4][68] ), .B(\w3[4][77] ), .Z(n5838) );
  XNOR U8143 ( .A(\w3[4][72] ), .B(\w3[4][92] ), .Z(n5837) );
  XNOR U8144 ( .A(n5838), .B(n5837), .Z(n5867) );
  XOR U8145 ( .A(n5867), .B(key[716]), .Z(n5841) );
  XNOR U8146 ( .A(\w3[4][84] ), .B(n5839), .Z(n5840) );
  XNOR U8147 ( .A(n5841), .B(n5840), .Z(\w1[5][76] ) );
  XOR U8148 ( .A(\w3[4][93] ), .B(\w3[4][69] ), .Z(n5870) );
  XOR U8149 ( .A(n5870), .B(key[717]), .Z(n5843) );
  XNOR U8150 ( .A(\w3[4][70] ), .B(\w3[4][78] ), .Z(n5842) );
  XNOR U8151 ( .A(n5843), .B(n5842), .Z(n5844) );
  XOR U8152 ( .A(\w3[4][85] ), .B(n5844), .Z(\w1[5][77] ) );
  XNOR U8153 ( .A(\w3[4][72] ), .B(\w3[4][79] ), .Z(n5879) );
  XNOR U8154 ( .A(n5845), .B(n5879), .Z(n5874) );
  XOR U8155 ( .A(n5874), .B(key[718]), .Z(n5848) );
  XNOR U8156 ( .A(\w3[4][86] ), .B(n5846), .Z(n5847) );
  XNOR U8157 ( .A(n5848), .B(n5847), .Z(\w1[5][78] ) );
  XOR U8158 ( .A(\w3[4][95] ), .B(\w3[4][71] ), .Z(n5877) );
  XOR U8159 ( .A(n5877), .B(key[719]), .Z(n5850) );
  XOR U8160 ( .A(\w3[4][72] ), .B(\w3[4][64] ), .Z(n5881) );
  XNOR U8161 ( .A(\w3[4][87] ), .B(n5881), .Z(n5849) );
  XNOR U8162 ( .A(n5850), .B(n5849), .Z(\w1[5][79] ) );
  XNOR U8163 ( .A(n5851), .B(key[647]), .Z(n5852) );
  XNOR U8164 ( .A(n5853), .B(n5852), .Z(n5854) );
  XNOR U8165 ( .A(\w3[4][0] ), .B(n5854), .Z(\w1[5][7] ) );
  XOR U8166 ( .A(n5881), .B(key[720]), .Z(n5856) );
  XNOR U8167 ( .A(\w3[4][88] ), .B(n5885), .Z(n5855) );
  XNOR U8168 ( .A(n5856), .B(n5855), .Z(\w1[5][80] ) );
  XOR U8169 ( .A(n5893), .B(key[721]), .Z(n5859) );
  XNOR U8170 ( .A(n5857), .B(\w3[4][73] ), .Z(n5858) );
  XNOR U8171 ( .A(n5859), .B(n5858), .Z(\w1[5][81] ) );
  XOR U8172 ( .A(n5860), .B(key[722]), .Z(n5863) );
  XNOR U8173 ( .A(n5861), .B(\w3[4][74] ), .Z(n5862) );
  XNOR U8174 ( .A(n5863), .B(n5862), .Z(\w1[5][82] ) );
  XOR U8175 ( .A(\w3[4][80] ), .B(\w3[4][84] ), .Z(n5897) );
  XOR U8176 ( .A(n5897), .B(key[723]), .Z(n5866) );
  XNOR U8177 ( .A(\w3[4][75] ), .B(n5864), .Z(n5865) );
  XNOR U8178 ( .A(n5866), .B(n5865), .Z(\w1[5][83] ) );
  XOR U8179 ( .A(\w3[4][80] ), .B(\w3[4][85] ), .Z(n5901) );
  XOR U8180 ( .A(n5901), .B(key[724]), .Z(n5869) );
  XNOR U8181 ( .A(\w3[4][76] ), .B(n5867), .Z(n5868) );
  XNOR U8182 ( .A(n5869), .B(n5868), .Z(\w1[5][84] ) );
  XOR U8183 ( .A(n5870), .B(key[725]), .Z(n5873) );
  XNOR U8184 ( .A(\w3[4][77] ), .B(n5871), .Z(n5872) );
  XNOR U8185 ( .A(n5873), .B(n5872), .Z(\w1[5][85] ) );
  XOR U8186 ( .A(\w3[4][80] ), .B(\w3[4][87] ), .Z(n5909) );
  XOR U8187 ( .A(n5909), .B(key[726]), .Z(n5876) );
  XNOR U8188 ( .A(\w3[4][78] ), .B(n5874), .Z(n5875) );
  XNOR U8189 ( .A(n5876), .B(n5875), .Z(\w1[5][86] ) );
  XNOR U8190 ( .A(n5877), .B(key[727]), .Z(n5878) );
  XNOR U8191 ( .A(n5879), .B(n5878), .Z(n5880) );
  XNOR U8192 ( .A(\w3[4][80] ), .B(n5880), .Z(\w1[5][87] ) );
  XOR U8193 ( .A(n5881), .B(key[728]), .Z(n5883) );
  XNOR U8194 ( .A(\w3[4][80] ), .B(\w3[4][81] ), .Z(n5882) );
  XNOR U8195 ( .A(n5883), .B(n5882), .Z(n5884) );
  XOR U8196 ( .A(\w3[4][89] ), .B(n5884), .Z(\w1[5][88] ) );
  XOR U8197 ( .A(\w3[4][82] ), .B(key[729]), .Z(n5887) );
  XNOR U8198 ( .A(n5885), .B(\w3[4][90] ), .Z(n5886) );
  XNOR U8199 ( .A(n5887), .B(n5886), .Z(n5888) );
  XOR U8200 ( .A(\w3[4][65] ), .B(n5888), .Z(\w1[5][89] ) );
  XOR U8201 ( .A(\w3[4][9] ), .B(key[648]), .Z(n5890) );
  XNOR U8202 ( .A(\w3[4][1] ), .B(\w3[4][0] ), .Z(n5889) );
  XNOR U8203 ( .A(n5890), .B(n5889), .Z(n5891) );
  XOR U8204 ( .A(n5892), .B(n5891), .Z(\w1[5][8] ) );
  XOR U8205 ( .A(\w3[4][83] ), .B(key[730]), .Z(n5895) );
  XNOR U8206 ( .A(n5893), .B(\w3[4][91] ), .Z(n5894) );
  XNOR U8207 ( .A(n5895), .B(n5894), .Z(n5896) );
  XOR U8208 ( .A(\w3[4][66] ), .B(n5896), .Z(\w1[5][90] ) );
  XOR U8209 ( .A(n5897), .B(key[731]), .Z(n5900) );
  XNOR U8210 ( .A(\w3[4][67] ), .B(n5898), .Z(n5899) );
  XNOR U8211 ( .A(n5900), .B(n5899), .Z(\w1[5][91] ) );
  XOR U8212 ( .A(n5901), .B(key[732]), .Z(n5904) );
  XNOR U8213 ( .A(\w3[4][68] ), .B(n5902), .Z(n5903) );
  XNOR U8214 ( .A(n5904), .B(n5903), .Z(\w1[5][92] ) );
  XOR U8215 ( .A(\w3[4][86] ), .B(key[733]), .Z(n5907) );
  XNOR U8216 ( .A(n5905), .B(\w3[4][94] ), .Z(n5906) );
  XNOR U8217 ( .A(n5907), .B(n5906), .Z(n5908) );
  XOR U8218 ( .A(\w3[4][69] ), .B(n5908), .Z(\w1[5][93] ) );
  XOR U8219 ( .A(n5909), .B(key[734]), .Z(n5912) );
  XNOR U8220 ( .A(\w3[4][70] ), .B(n5910), .Z(n5911) );
  XNOR U8221 ( .A(n5912), .B(n5911), .Z(\w1[5][94] ) );
  XOR U8222 ( .A(n5913), .B(key[735]), .Z(n5916) );
  XNOR U8223 ( .A(n5914), .B(\w3[4][71] ), .Z(n5915) );
  XNOR U8224 ( .A(n5916), .B(n5915), .Z(\w1[5][95] ) );
  XOR U8225 ( .A(\w3[4][104] ), .B(key[736]), .Z(n5920) );
  XOR U8226 ( .A(n5918), .B(n5917), .Z(n5919) );
  XNOR U8227 ( .A(n5920), .B(n5919), .Z(\w1[5][96] ) );
  XOR U8228 ( .A(n5921), .B(key[737]), .Z(n5924) );
  XNOR U8229 ( .A(\w3[4][121] ), .B(n5922), .Z(n5923) );
  XNOR U8230 ( .A(n5924), .B(n5923), .Z(\w1[5][97] ) );
  XOR U8231 ( .A(n5925), .B(key[738]), .Z(n5928) );
  XNOR U8232 ( .A(\w3[4][122] ), .B(n5926), .Z(n5927) );
  XNOR U8233 ( .A(n5928), .B(n5927), .Z(\w1[5][98] ) );
  XOR U8234 ( .A(n5929), .B(key[739]), .Z(n5932) );
  XNOR U8235 ( .A(n5930), .B(\w3[4][123] ), .Z(n5931) );
  XNOR U8236 ( .A(n5932), .B(n5931), .Z(\w1[5][99] ) );
  XOR U8237 ( .A(\w3[4][10] ), .B(key[649]), .Z(n5934) );
  XNOR U8238 ( .A(\w3[4][2] ), .B(\w3[4][17] ), .Z(n5933) );
  XNOR U8239 ( .A(n5934), .B(n5933), .Z(n5935) );
  XOR U8240 ( .A(n5936), .B(n5935), .Z(\w1[5][9] ) );
  XOR U8241 ( .A(\w3[5][8] ), .B(key[768]), .Z(n5938) );
  XOR U8242 ( .A(\w3[5][1] ), .B(\w3[5][25] ), .Z(n6360) );
  XOR U8243 ( .A(\w3[5][16] ), .B(\w3[5][24] ), .Z(n6316) );
  XNOR U8244 ( .A(n6360), .B(n6316), .Z(n5937) );
  XNOR U8245 ( .A(n5938), .B(n5937), .Z(\w1[6][0] ) );
  XOR U8246 ( .A(\w3[5][96] ), .B(\w3[5][101] ), .Z(n5963) );
  XOR U8247 ( .A(n5963), .B(key[868]), .Z(n5942) );
  XOR U8248 ( .A(\w3[5][116] ), .B(\w3[5][125] ), .Z(n5940) );
  XNOR U8249 ( .A(\w3[5][120] ), .B(\w3[5][108] ), .Z(n5939) );
  XNOR U8250 ( .A(n5940), .B(n5939), .Z(n6021) );
  XNOR U8251 ( .A(\w3[5][124] ), .B(n6021), .Z(n5941) );
  XNOR U8252 ( .A(n5942), .B(n5941), .Z(\w1[6][100] ) );
  XOR U8253 ( .A(\w3[5][102] ), .B(\w3[5][126] ), .Z(n5972) );
  XOR U8254 ( .A(n5972), .B(key[869]), .Z(n5944) );
  XOR U8255 ( .A(\w3[5][109] ), .B(\w3[5][117] ), .Z(n6024) );
  XNOR U8256 ( .A(\w3[5][125] ), .B(n6024), .Z(n5943) );
  XNOR U8257 ( .A(n5944), .B(n5943), .Z(\w1[6][101] ) );
  XOR U8258 ( .A(\w3[5][96] ), .B(\w3[5][103] ), .Z(n5973) );
  XOR U8259 ( .A(n5973), .B(key[870]), .Z(n5946) );
  XOR U8260 ( .A(\w3[5][110] ), .B(\w3[5][118] ), .Z(n5992) );
  XNOR U8261 ( .A(\w3[5][120] ), .B(\w3[5][127] ), .Z(n5948) );
  XNOR U8262 ( .A(n5992), .B(n5948), .Z(n6029) );
  XNOR U8263 ( .A(\w3[5][126] ), .B(n6029), .Z(n5945) );
  XNOR U8264 ( .A(n5946), .B(n5945), .Z(\w1[6][102] ) );
  XOR U8265 ( .A(\w3[5][111] ), .B(\w3[5][119] ), .Z(n6032) );
  XNOR U8266 ( .A(n6032), .B(key[871]), .Z(n5947) );
  XNOR U8267 ( .A(n5948), .B(n5947), .Z(n5949) );
  XNOR U8268 ( .A(\w3[5][96] ), .B(n5949), .Z(\w1[6][103] ) );
  XOR U8269 ( .A(\w3[5][105] ), .B(\w3[5][97] ), .Z(n5980) );
  XOR U8270 ( .A(n5980), .B(key[872]), .Z(n5951) );
  XOR U8271 ( .A(\w3[5][120] ), .B(\w3[5][112] ), .Z(n6342) );
  XNOR U8272 ( .A(\w3[5][96] ), .B(n6342), .Z(n5950) );
  XNOR U8273 ( .A(n5951), .B(n5950), .Z(\w1[6][104] ) );
  XOR U8274 ( .A(\w3[5][106] ), .B(\w3[5][98] ), .Z(n5953) );
  XOR U8275 ( .A(\w3[5][97] ), .B(\w3[5][121] ), .Z(n6341) );
  XNOR U8276 ( .A(n6341), .B(key[873]), .Z(n5952) );
  XNOR U8277 ( .A(n5953), .B(n5952), .Z(n5954) );
  XOR U8278 ( .A(\w3[5][113] ), .B(n5954), .Z(\w1[6][105] ) );
  XOR U8279 ( .A(\w3[5][107] ), .B(\w3[5][114] ), .Z(n5956) );
  XOR U8280 ( .A(\w3[5][98] ), .B(\w3[5][122] ), .Z(n6346) );
  XNOR U8281 ( .A(n6346), .B(key[874]), .Z(n5955) );
  XNOR U8282 ( .A(n5956), .B(n5955), .Z(n5957) );
  XOR U8283 ( .A(\w3[5][99] ), .B(n5957), .Z(\w1[6][106] ) );
  XOR U8284 ( .A(\w3[5][99] ), .B(\w3[5][123] ), .Z(n6350) );
  XNOR U8285 ( .A(\w3[5][108] ), .B(n6350), .Z(n5958) );
  XNOR U8286 ( .A(\w3[5][104] ), .B(n5958), .Z(n5985) );
  XOR U8287 ( .A(n5985), .B(key[875]), .Z(n5960) );
  XOR U8288 ( .A(\w3[5][96] ), .B(\w3[5][100] ), .Z(n6354) );
  XNOR U8289 ( .A(\w3[5][115] ), .B(n6354), .Z(n5959) );
  XNOR U8290 ( .A(n5960), .B(n5959), .Z(\w1[6][107] ) );
  XOR U8291 ( .A(\w3[5][100] ), .B(\w3[5][104] ), .Z(n5962) );
  XNOR U8292 ( .A(\w3[5][124] ), .B(\w3[5][109] ), .Z(n5961) );
  XNOR U8293 ( .A(n5962), .B(n5961), .Z(n5988) );
  XOR U8294 ( .A(n5988), .B(key[876]), .Z(n5965) );
  XNOR U8295 ( .A(\w3[5][116] ), .B(n5963), .Z(n5964) );
  XNOR U8296 ( .A(n5965), .B(n5964), .Z(\w1[6][108] ) );
  XOR U8297 ( .A(\w3[5][125] ), .B(\w3[5][101] ), .Z(n5991) );
  XOR U8298 ( .A(n5991), .B(key[877]), .Z(n5967) );
  XNOR U8299 ( .A(\w3[5][102] ), .B(\w3[5][110] ), .Z(n5966) );
  XNOR U8300 ( .A(n5967), .B(n5966), .Z(n5968) );
  XOR U8301 ( .A(\w3[5][117] ), .B(n5968), .Z(\w1[6][109] ) );
  XOR U8302 ( .A(\w3[5][11] ), .B(\w3[5][18] ), .Z(n5970) );
  XOR U8303 ( .A(\w3[5][2] ), .B(\w3[5][26] ), .Z(n6055) );
  XNOR U8304 ( .A(n6055), .B(key[778]), .Z(n5969) );
  XNOR U8305 ( .A(n5970), .B(n5969), .Z(n5971) );
  XOR U8306 ( .A(\w3[5][3] ), .B(n5971), .Z(\w1[6][10] ) );
  XNOR U8307 ( .A(\w3[5][111] ), .B(\w3[5][104] ), .Z(n6000) );
  XNOR U8308 ( .A(n5972), .B(n6000), .Z(n5995) );
  XOR U8309 ( .A(n5995), .B(key[878]), .Z(n5975) );
  XNOR U8310 ( .A(\w3[5][118] ), .B(n5973), .Z(n5974) );
  XNOR U8311 ( .A(n5975), .B(n5974), .Z(\w1[6][110] ) );
  XOR U8312 ( .A(\w3[5][127] ), .B(\w3[5][103] ), .Z(n5998) );
  XOR U8313 ( .A(n5998), .B(key[879]), .Z(n5977) );
  XOR U8314 ( .A(\w3[5][96] ), .B(\w3[5][104] ), .Z(n6005) );
  XNOR U8315 ( .A(\w3[5][119] ), .B(n6005), .Z(n5976) );
  XNOR U8316 ( .A(n5977), .B(n5976), .Z(\w1[6][111] ) );
  XOR U8317 ( .A(\w3[5][105] ), .B(\w3[5][113] ), .Z(n6345) );
  XOR U8318 ( .A(n6345), .B(key[880]), .Z(n5979) );
  XNOR U8319 ( .A(\w3[5][120] ), .B(n6005), .Z(n5978) );
  XNOR U8320 ( .A(n5979), .B(n5978), .Z(\w1[6][112] ) );
  XOR U8321 ( .A(\w3[5][106] ), .B(\w3[5][114] ), .Z(n6349) );
  XOR U8322 ( .A(n6349), .B(key[881]), .Z(n5982) );
  XNOR U8323 ( .A(n5980), .B(\w3[5][121] ), .Z(n5981) );
  XNOR U8324 ( .A(n5982), .B(n5981), .Z(\w1[6][113] ) );
  XOR U8325 ( .A(\w3[5][107] ), .B(\w3[5][115] ), .Z(n6016) );
  XOR U8326 ( .A(n6016), .B(key[882]), .Z(n5984) );
  XNOR U8327 ( .A(\w3[5][106] ), .B(n6346), .Z(n5983) );
  XNOR U8328 ( .A(n5984), .B(n5983), .Z(\w1[6][114] ) );
  XOR U8329 ( .A(\w3[5][116] ), .B(\w3[5][112] ), .Z(n6017) );
  XOR U8330 ( .A(n6017), .B(key[883]), .Z(n5987) );
  XNOR U8331 ( .A(\w3[5][107] ), .B(n5985), .Z(n5986) );
  XNOR U8332 ( .A(n5987), .B(n5986), .Z(\w1[6][115] ) );
  XOR U8333 ( .A(\w3[5][117] ), .B(\w3[5][112] ), .Z(n6020) );
  XOR U8334 ( .A(n6020), .B(key[884]), .Z(n5990) );
  XNOR U8335 ( .A(\w3[5][108] ), .B(n5988), .Z(n5989) );
  XNOR U8336 ( .A(n5990), .B(n5989), .Z(\w1[6][116] ) );
  XOR U8337 ( .A(n5991), .B(key[885]), .Z(n5994) );
  XNOR U8338 ( .A(\w3[5][109] ), .B(n5992), .Z(n5993) );
  XNOR U8339 ( .A(n5994), .B(n5993), .Z(\w1[6][117] ) );
  XOR U8340 ( .A(\w3[5][119] ), .B(\w3[5][112] ), .Z(n6028) );
  XOR U8341 ( .A(n6028), .B(key[886]), .Z(n5997) );
  XNOR U8342 ( .A(\w3[5][110] ), .B(n5995), .Z(n5996) );
  XNOR U8343 ( .A(n5997), .B(n5996), .Z(\w1[6][118] ) );
  XNOR U8344 ( .A(n5998), .B(key[887]), .Z(n5999) );
  XNOR U8345 ( .A(n6000), .B(n5999), .Z(n6001) );
  XNOR U8346 ( .A(\w3[5][112] ), .B(n6001), .Z(\w1[6][119] ) );
  XOR U8347 ( .A(\w3[5][3] ), .B(\w3[5][27] ), .Z(n6096) );
  XNOR U8348 ( .A(\w3[5][8] ), .B(\w3[5][12] ), .Z(n6002) );
  XNOR U8349 ( .A(n6096), .B(n6002), .Z(n6052) );
  XOR U8350 ( .A(n6052), .B(key[779]), .Z(n6004) );
  XOR U8351 ( .A(\w3[5][0] ), .B(\w3[5][4] ), .Z(n6126) );
  XNOR U8352 ( .A(\w3[5][19] ), .B(n6126), .Z(n6003) );
  XNOR U8353 ( .A(n6004), .B(n6003), .Z(\w1[6][11] ) );
  XOR U8354 ( .A(n6005), .B(key[888]), .Z(n6007) );
  XNOR U8355 ( .A(\w3[5][113] ), .B(\w3[5][121] ), .Z(n6006) );
  XNOR U8356 ( .A(n6007), .B(n6006), .Z(n6008) );
  XOR U8357 ( .A(\w3[5][112] ), .B(n6008), .Z(\w1[6][120] ) );
  XOR U8358 ( .A(n6345), .B(key[889]), .Z(n6010) );
  XNOR U8359 ( .A(\w3[5][122] ), .B(\w3[5][114] ), .Z(n6009) );
  XNOR U8360 ( .A(n6010), .B(n6009), .Z(n6011) );
  XOR U8361 ( .A(\w3[5][97] ), .B(n6011), .Z(\w1[6][121] ) );
  XOR U8362 ( .A(n6349), .B(key[890]), .Z(n6013) );
  XNOR U8363 ( .A(\w3[5][115] ), .B(\w3[5][123] ), .Z(n6012) );
  XNOR U8364 ( .A(n6013), .B(n6012), .Z(n6014) );
  XOR U8365 ( .A(\w3[5][98] ), .B(n6014), .Z(\w1[6][122] ) );
  XNOR U8366 ( .A(\w3[5][124] ), .B(\w3[5][120] ), .Z(n6015) );
  XNOR U8367 ( .A(n6016), .B(n6015), .Z(n6353) );
  XOR U8368 ( .A(n6353), .B(key[891]), .Z(n6019) );
  XNOR U8369 ( .A(\w3[5][99] ), .B(n6017), .Z(n6018) );
  XNOR U8370 ( .A(n6019), .B(n6018), .Z(\w1[6][123] ) );
  XOR U8371 ( .A(n6020), .B(key[892]), .Z(n6023) );
  XNOR U8372 ( .A(n6021), .B(\w3[5][100] ), .Z(n6022) );
  XNOR U8373 ( .A(n6023), .B(n6022), .Z(\w1[6][124] ) );
  XOR U8374 ( .A(\w3[5][118] ), .B(key[893]), .Z(n6026) );
  XNOR U8375 ( .A(n6024), .B(\w3[5][126] ), .Z(n6025) );
  XNOR U8376 ( .A(n6026), .B(n6025), .Z(n6027) );
  XOR U8377 ( .A(\w3[5][101] ), .B(n6027), .Z(\w1[6][125] ) );
  XOR U8378 ( .A(n6028), .B(key[894]), .Z(n6031) );
  XNOR U8379 ( .A(\w3[5][102] ), .B(n6029), .Z(n6030) );
  XNOR U8380 ( .A(n6031), .B(n6030), .Z(\w1[6][126] ) );
  XOR U8381 ( .A(n6342), .B(key[895]), .Z(n6034) );
  XNOR U8382 ( .A(\w3[5][103] ), .B(n6032), .Z(n6033) );
  XNOR U8383 ( .A(n6034), .B(n6033), .Z(\w1[6][127] ) );
  XOR U8384 ( .A(\w3[5][13] ), .B(\w3[5][28] ), .Z(n6036) );
  XNOR U8385 ( .A(\w3[5][8] ), .B(\w3[5][4] ), .Z(n6035) );
  XNOR U8386 ( .A(n6036), .B(n6035), .Z(n6058) );
  XOR U8387 ( .A(n6058), .B(key[780]), .Z(n6038) );
  XOR U8388 ( .A(\w3[5][0] ), .B(\w3[5][5] ), .Z(n6163) );
  XNOR U8389 ( .A(\w3[5][20] ), .B(n6163), .Z(n6037) );
  XNOR U8390 ( .A(n6038), .B(n6037), .Z(\w1[6][12] ) );
  XOR U8391 ( .A(\w3[5][14] ), .B(\w3[5][6] ), .Z(n6040) );
  XOR U8392 ( .A(\w3[5][5] ), .B(\w3[5][29] ), .Z(n6061) );
  XNOR U8393 ( .A(n6061), .B(key[781]), .Z(n6039) );
  XNOR U8394 ( .A(n6040), .B(n6039), .Z(n6041) );
  XOR U8395 ( .A(\w3[5][21] ), .B(n6041), .Z(\w1[6][13] ) );
  XOR U8396 ( .A(\w3[5][6] ), .B(\w3[5][30] ), .Z(n6204) );
  XNOR U8397 ( .A(\w3[5][8] ), .B(\w3[5][15] ), .Z(n6069) );
  XNOR U8398 ( .A(n6204), .B(n6069), .Z(n6064) );
  XOR U8399 ( .A(n6064), .B(key[782]), .Z(n6043) );
  XOR U8400 ( .A(\w3[5][0] ), .B(\w3[5][7] ), .Z(n6239) );
  XNOR U8401 ( .A(\w3[5][22] ), .B(n6239), .Z(n6042) );
  XNOR U8402 ( .A(n6043), .B(n6042), .Z(\w1[6][14] ) );
  XOR U8403 ( .A(\w3[5][7] ), .B(\w3[5][31] ), .Z(n6067) );
  XOR U8404 ( .A(n6067), .B(key[783]), .Z(n6045) );
  XOR U8405 ( .A(\w3[5][8] ), .B(\w3[5][0] ), .Z(n6071) );
  XNOR U8406 ( .A(\w3[5][23] ), .B(n6071), .Z(n6044) );
  XNOR U8407 ( .A(n6045), .B(n6044), .Z(\w1[6][15] ) );
  XOR U8408 ( .A(\w3[5][17] ), .B(\w3[5][9] ), .Z(n6075) );
  XOR U8409 ( .A(n6075), .B(key[784]), .Z(n6047) );
  XNOR U8410 ( .A(\w3[5][24] ), .B(n6071), .Z(n6046) );
  XNOR U8411 ( .A(n6047), .B(n6046), .Z(\w1[6][16] ) );
  XOR U8412 ( .A(\w3[5][18] ), .B(\w3[5][10] ), .Z(n6095) );
  XOR U8413 ( .A(n6095), .B(key[785]), .Z(n6049) );
  XNOR U8414 ( .A(n6360), .B(\w3[5][9] ), .Z(n6048) );
  XNOR U8415 ( .A(n6049), .B(n6048), .Z(\w1[6][17] ) );
  XOR U8416 ( .A(\w3[5][11] ), .B(\w3[5][19] ), .Z(n6083) );
  XOR U8417 ( .A(n6083), .B(key[786]), .Z(n6051) );
  XNOR U8418 ( .A(n6055), .B(\w3[5][10] ), .Z(n6050) );
  XNOR U8419 ( .A(n6051), .B(n6050), .Z(\w1[6][18] ) );
  XOR U8420 ( .A(\w3[5][16] ), .B(\w3[5][20] ), .Z(n6084) );
  XOR U8421 ( .A(n6084), .B(key[787]), .Z(n6054) );
  XNOR U8422 ( .A(\w3[5][11] ), .B(n6052), .Z(n6053) );
  XNOR U8423 ( .A(n6054), .B(n6053), .Z(\w1[6][19] ) );
  XOR U8424 ( .A(n6075), .B(key[769]), .Z(n6057) );
  XNOR U8425 ( .A(\w3[5][25] ), .B(n6055), .Z(n6056) );
  XNOR U8426 ( .A(n6057), .B(n6056), .Z(\w1[6][1] ) );
  XOR U8427 ( .A(\w3[5][16] ), .B(\w3[5][21] ), .Z(n6089) );
  XOR U8428 ( .A(n6089), .B(key[788]), .Z(n6060) );
  XNOR U8429 ( .A(\w3[5][12] ), .B(n6058), .Z(n6059) );
  XNOR U8430 ( .A(n6060), .B(n6059), .Z(\w1[6][20] ) );
  XOR U8431 ( .A(\w3[5][14] ), .B(\w3[5][22] ), .Z(n6099) );
  XOR U8432 ( .A(n6099), .B(key[789]), .Z(n6063) );
  XNOR U8433 ( .A(\w3[5][13] ), .B(n6061), .Z(n6062) );
  XNOR U8434 ( .A(n6063), .B(n6062), .Z(\w1[6][21] ) );
  XOR U8435 ( .A(\w3[5][16] ), .B(\w3[5][23] ), .Z(n6100) );
  XOR U8436 ( .A(n6100), .B(key[790]), .Z(n6066) );
  XNOR U8437 ( .A(\w3[5][14] ), .B(n6064), .Z(n6065) );
  XNOR U8438 ( .A(n6066), .B(n6065), .Z(\w1[6][22] ) );
  XNOR U8439 ( .A(n6067), .B(key[791]), .Z(n6068) );
  XNOR U8440 ( .A(n6069), .B(n6068), .Z(n6070) );
  XNOR U8441 ( .A(\w3[5][16] ), .B(n6070), .Z(\w1[6][23] ) );
  XOR U8442 ( .A(\w3[5][17] ), .B(key[792]), .Z(n6073) );
  XNOR U8443 ( .A(\w3[5][25] ), .B(n6071), .Z(n6072) );
  XNOR U8444 ( .A(n6073), .B(n6072), .Z(n6074) );
  XOR U8445 ( .A(\w3[5][16] ), .B(n6074), .Z(\w1[6][24] ) );
  XOR U8446 ( .A(n6075), .B(key[793]), .Z(n6077) );
  XNOR U8447 ( .A(\w3[5][1] ), .B(\w3[5][26] ), .Z(n6076) );
  XNOR U8448 ( .A(n6077), .B(n6076), .Z(n6078) );
  XOR U8449 ( .A(\w3[5][18] ), .B(n6078), .Z(\w1[6][25] ) );
  XOR U8450 ( .A(n6095), .B(key[794]), .Z(n6080) );
  XNOR U8451 ( .A(\w3[5][2] ), .B(\w3[5][19] ), .Z(n6079) );
  XNOR U8452 ( .A(n6080), .B(n6079), .Z(n6081) );
  XOR U8453 ( .A(\w3[5][27] ), .B(n6081), .Z(\w1[6][26] ) );
  XNOR U8454 ( .A(\w3[5][24] ), .B(\w3[5][28] ), .Z(n6082) );
  XNOR U8455 ( .A(n6083), .B(n6082), .Z(n6125) );
  XOR U8456 ( .A(n6125), .B(key[795]), .Z(n6086) );
  XNOR U8457 ( .A(\w3[5][3] ), .B(n6084), .Z(n6085) );
  XNOR U8458 ( .A(n6086), .B(n6085), .Z(\w1[6][27] ) );
  XOR U8459 ( .A(\w3[5][20] ), .B(\w3[5][29] ), .Z(n6088) );
  XNOR U8460 ( .A(\w3[5][24] ), .B(\w3[5][12] ), .Z(n6087) );
  XNOR U8461 ( .A(n6088), .B(n6087), .Z(n6162) );
  XOR U8462 ( .A(n6162), .B(key[796]), .Z(n6091) );
  XNOR U8463 ( .A(\w3[5][4] ), .B(n6089), .Z(n6090) );
  XNOR U8464 ( .A(n6091), .B(n6090), .Z(\w1[6][28] ) );
  XOR U8465 ( .A(\w3[5][13] ), .B(\w3[5][21] ), .Z(n6203) );
  XOR U8466 ( .A(n6203), .B(key[797]), .Z(n6093) );
  XNOR U8467 ( .A(\w3[5][22] ), .B(\w3[5][30] ), .Z(n6092) );
  XNOR U8468 ( .A(n6093), .B(n6092), .Z(n6094) );
  XOR U8469 ( .A(\w3[5][5] ), .B(n6094), .Z(\w1[6][29] ) );
  XOR U8470 ( .A(n6095), .B(key[770]), .Z(n6098) );
  XNOR U8471 ( .A(\w3[5][26] ), .B(n6096), .Z(n6097) );
  XNOR U8472 ( .A(n6098), .B(n6097), .Z(\w1[6][2] ) );
  XNOR U8473 ( .A(\w3[5][24] ), .B(\w3[5][31] ), .Z(n6277) );
  XNOR U8474 ( .A(n6099), .B(n6277), .Z(n6238) );
  XOR U8475 ( .A(n6238), .B(key[798]), .Z(n6102) );
  XNOR U8476 ( .A(\w3[5][6] ), .B(n6100), .Z(n6101) );
  XNOR U8477 ( .A(n6102), .B(n6101), .Z(\w1[6][30] ) );
  XOR U8478 ( .A(\w3[5][15] ), .B(\w3[5][23] ), .Z(n6275) );
  XOR U8479 ( .A(n6275), .B(key[799]), .Z(n6104) );
  XNOR U8480 ( .A(n6316), .B(\w3[5][7] ), .Z(n6103) );
  XNOR U8481 ( .A(n6104), .B(n6103), .Z(\w1[6][31] ) );
  XOR U8482 ( .A(\w3[5][33] ), .B(\w3[5][57] ), .Z(n6159) );
  XOR U8483 ( .A(n6159), .B(key[800]), .Z(n6106) );
  XOR U8484 ( .A(\w3[5][48] ), .B(\w3[5][56] ), .Z(n6220) );
  XNOR U8485 ( .A(n6220), .B(\w3[5][40] ), .Z(n6105) );
  XNOR U8486 ( .A(n6106), .B(n6105), .Z(\w1[6][32] ) );
  XOR U8487 ( .A(\w3[5][34] ), .B(\w3[5][58] ), .Z(n6167) );
  XOR U8488 ( .A(n6167), .B(key[801]), .Z(n6108) );
  XOR U8489 ( .A(\w3[5][41] ), .B(\w3[5][49] ), .Z(n6191) );
  XNOR U8490 ( .A(\w3[5][57] ), .B(n6191), .Z(n6107) );
  XNOR U8491 ( .A(n6108), .B(n6107), .Z(\w1[6][33] ) );
  XOR U8492 ( .A(\w3[5][35] ), .B(\w3[5][59] ), .Z(n6138) );
  XOR U8493 ( .A(n6138), .B(key[802]), .Z(n6110) );
  XOR U8494 ( .A(\w3[5][42] ), .B(\w3[5][50] ), .Z(n6195) );
  XNOR U8495 ( .A(\w3[5][58] ), .B(n6195), .Z(n6109) );
  XNOR U8496 ( .A(n6110), .B(n6109), .Z(\w1[6][34] ) );
  XOR U8497 ( .A(\w3[5][36] ), .B(\w3[5][32] ), .Z(n6140) );
  XOR U8498 ( .A(n6140), .B(key[803]), .Z(n6113) );
  XOR U8499 ( .A(\w3[5][43] ), .B(\w3[5][51] ), .Z(n6166) );
  XNOR U8500 ( .A(\w3[5][56] ), .B(n6166), .Z(n6111) );
  XNOR U8501 ( .A(\w3[5][60] ), .B(n6111), .Z(n6200) );
  XNOR U8502 ( .A(\w3[5][59] ), .B(n6200), .Z(n6112) );
  XNOR U8503 ( .A(n6113), .B(n6112), .Z(\w1[6][35] ) );
  XOR U8504 ( .A(\w3[5][32] ), .B(\w3[5][37] ), .Z(n6145) );
  XOR U8505 ( .A(n6145), .B(key[804]), .Z(n6117) );
  XOR U8506 ( .A(\w3[5][52] ), .B(\w3[5][61] ), .Z(n6115) );
  XNOR U8507 ( .A(\w3[5][56] ), .B(\w3[5][44] ), .Z(n6114) );
  XNOR U8508 ( .A(n6115), .B(n6114), .Z(n6208) );
  XNOR U8509 ( .A(\w3[5][60] ), .B(n6208), .Z(n6116) );
  XNOR U8510 ( .A(n6117), .B(n6116), .Z(\w1[6][36] ) );
  XOR U8511 ( .A(\w3[5][38] ), .B(\w3[5][62] ), .Z(n6151) );
  XOR U8512 ( .A(n6151), .B(key[805]), .Z(n6119) );
  XOR U8513 ( .A(\w3[5][45] ), .B(\w3[5][53] ), .Z(n6211) );
  XNOR U8514 ( .A(\w3[5][61] ), .B(n6211), .Z(n6118) );
  XNOR U8515 ( .A(n6119), .B(n6118), .Z(\w1[6][37] ) );
  XOR U8516 ( .A(\w3[5][32] ), .B(\w3[5][39] ), .Z(n6152) );
  XOR U8517 ( .A(n6152), .B(key[806]), .Z(n6121) );
  XOR U8518 ( .A(\w3[5][46] ), .B(\w3[5][54] ), .Z(n6177) );
  XNOR U8519 ( .A(\w3[5][56] ), .B(\w3[5][63] ), .Z(n6123) );
  XNOR U8520 ( .A(n6177), .B(n6123), .Z(n6216) );
  XNOR U8521 ( .A(\w3[5][62] ), .B(n6216), .Z(n6120) );
  XNOR U8522 ( .A(n6121), .B(n6120), .Z(\w1[6][38] ) );
  XOR U8523 ( .A(\w3[5][47] ), .B(\w3[5][55] ), .Z(n6219) );
  XNOR U8524 ( .A(n6219), .B(key[807]), .Z(n6122) );
  XNOR U8525 ( .A(n6123), .B(n6122), .Z(n6124) );
  XNOR U8526 ( .A(\w3[5][32] ), .B(n6124), .Z(\w1[6][39] ) );
  XOR U8527 ( .A(n6125), .B(key[771]), .Z(n6128) );
  XNOR U8528 ( .A(n6126), .B(\w3[5][27] ), .Z(n6127) );
  XNOR U8529 ( .A(n6128), .B(n6127), .Z(\w1[6][3] ) );
  XOR U8530 ( .A(\w3[5][32] ), .B(key[808]), .Z(n6130) );
  XNOR U8531 ( .A(\w3[5][33] ), .B(\w3[5][41] ), .Z(n6129) );
  XNOR U8532 ( .A(n6130), .B(n6129), .Z(n6131) );
  XOR U8533 ( .A(n6220), .B(n6131), .Z(\w1[6][40] ) );
  XOR U8534 ( .A(\w3[5][42] ), .B(key[809]), .Z(n6133) );
  XNOR U8535 ( .A(\w3[5][49] ), .B(\w3[5][34] ), .Z(n6132) );
  XNOR U8536 ( .A(n6133), .B(n6132), .Z(n6134) );
  XOR U8537 ( .A(n6159), .B(n6134), .Z(\w1[6][41] ) );
  XOR U8538 ( .A(\w3[5][43] ), .B(key[810]), .Z(n6136) );
  XNOR U8539 ( .A(\w3[5][50] ), .B(\w3[5][35] ), .Z(n6135) );
  XNOR U8540 ( .A(n6136), .B(n6135), .Z(n6137) );
  XOR U8541 ( .A(n6167), .B(n6137), .Z(\w1[6][42] ) );
  XNOR U8542 ( .A(\w3[5][40] ), .B(n6138), .Z(n6139) );
  XNOR U8543 ( .A(\w3[5][44] ), .B(n6139), .Z(n6170) );
  XOR U8544 ( .A(n6170), .B(key[811]), .Z(n6142) );
  XNOR U8545 ( .A(\w3[5][51] ), .B(n6140), .Z(n6141) );
  XNOR U8546 ( .A(n6142), .B(n6141), .Z(\w1[6][43] ) );
  XOR U8547 ( .A(\w3[5][36] ), .B(\w3[5][45] ), .Z(n6144) );
  XNOR U8548 ( .A(\w3[5][40] ), .B(\w3[5][60] ), .Z(n6143) );
  XNOR U8549 ( .A(n6144), .B(n6143), .Z(n6173) );
  XOR U8550 ( .A(n6173), .B(key[812]), .Z(n6147) );
  XNOR U8551 ( .A(\w3[5][52] ), .B(n6145), .Z(n6146) );
  XNOR U8552 ( .A(n6147), .B(n6146), .Z(\w1[6][44] ) );
  XOR U8553 ( .A(\w3[5][61] ), .B(\w3[5][37] ), .Z(n6176) );
  XOR U8554 ( .A(n6176), .B(key[813]), .Z(n6149) );
  XNOR U8555 ( .A(\w3[5][38] ), .B(\w3[5][46] ), .Z(n6148) );
  XNOR U8556 ( .A(n6149), .B(n6148), .Z(n6150) );
  XOR U8557 ( .A(\w3[5][53] ), .B(n6150), .Z(\w1[6][45] ) );
  XNOR U8558 ( .A(\w3[5][40] ), .B(\w3[5][47] ), .Z(n6185) );
  XNOR U8559 ( .A(n6151), .B(n6185), .Z(n6180) );
  XOR U8560 ( .A(n6180), .B(key[814]), .Z(n6154) );
  XNOR U8561 ( .A(\w3[5][54] ), .B(n6152), .Z(n6153) );
  XNOR U8562 ( .A(n6154), .B(n6153), .Z(\w1[6][46] ) );
  XOR U8563 ( .A(\w3[5][63] ), .B(\w3[5][39] ), .Z(n6183) );
  XOR U8564 ( .A(n6183), .B(key[815]), .Z(n6156) );
  XOR U8565 ( .A(\w3[5][40] ), .B(\w3[5][32] ), .Z(n6187) );
  XNOR U8566 ( .A(\w3[5][55] ), .B(n6187), .Z(n6155) );
  XNOR U8567 ( .A(n6156), .B(n6155), .Z(\w1[6][47] ) );
  XOR U8568 ( .A(n6187), .B(key[816]), .Z(n6158) );
  XNOR U8569 ( .A(\w3[5][56] ), .B(n6191), .Z(n6157) );
  XNOR U8570 ( .A(n6158), .B(n6157), .Z(\w1[6][48] ) );
  XOR U8571 ( .A(n6195), .B(key[817]), .Z(n6161) );
  XNOR U8572 ( .A(n6159), .B(\w3[5][41] ), .Z(n6160) );
  XNOR U8573 ( .A(n6161), .B(n6160), .Z(\w1[6][49] ) );
  XOR U8574 ( .A(n6162), .B(key[772]), .Z(n6165) );
  XNOR U8575 ( .A(n6163), .B(\w3[5][28] ), .Z(n6164) );
  XNOR U8576 ( .A(n6165), .B(n6164), .Z(\w1[6][4] ) );
  XOR U8577 ( .A(n6166), .B(key[818]), .Z(n6169) );
  XNOR U8578 ( .A(n6167), .B(\w3[5][42] ), .Z(n6168) );
  XNOR U8579 ( .A(n6169), .B(n6168), .Z(\w1[6][50] ) );
  XOR U8580 ( .A(\w3[5][48] ), .B(\w3[5][52] ), .Z(n6199) );
  XOR U8581 ( .A(n6199), .B(key[819]), .Z(n6172) );
  XNOR U8582 ( .A(\w3[5][43] ), .B(n6170), .Z(n6171) );
  XNOR U8583 ( .A(n6172), .B(n6171), .Z(\w1[6][51] ) );
  XOR U8584 ( .A(\w3[5][48] ), .B(\w3[5][53] ), .Z(n6207) );
  XOR U8585 ( .A(n6207), .B(key[820]), .Z(n6175) );
  XNOR U8586 ( .A(\w3[5][44] ), .B(n6173), .Z(n6174) );
  XNOR U8587 ( .A(n6175), .B(n6174), .Z(\w1[6][52] ) );
  XOR U8588 ( .A(n6176), .B(key[821]), .Z(n6179) );
  XNOR U8589 ( .A(\w3[5][45] ), .B(n6177), .Z(n6178) );
  XNOR U8590 ( .A(n6179), .B(n6178), .Z(\w1[6][53] ) );
  XOR U8591 ( .A(\w3[5][48] ), .B(\w3[5][55] ), .Z(n6215) );
  XOR U8592 ( .A(n6215), .B(key[822]), .Z(n6182) );
  XNOR U8593 ( .A(\w3[5][46] ), .B(n6180), .Z(n6181) );
  XNOR U8594 ( .A(n6182), .B(n6181), .Z(\w1[6][54] ) );
  XNOR U8595 ( .A(n6183), .B(key[823]), .Z(n6184) );
  XNOR U8596 ( .A(n6185), .B(n6184), .Z(n6186) );
  XNOR U8597 ( .A(\w3[5][48] ), .B(n6186), .Z(\w1[6][55] ) );
  XOR U8598 ( .A(n6187), .B(key[824]), .Z(n6189) );
  XNOR U8599 ( .A(\w3[5][48] ), .B(\w3[5][49] ), .Z(n6188) );
  XNOR U8600 ( .A(n6189), .B(n6188), .Z(n6190) );
  XOR U8601 ( .A(\w3[5][57] ), .B(n6190), .Z(\w1[6][56] ) );
  XOR U8602 ( .A(\w3[5][50] ), .B(key[825]), .Z(n6193) );
  XNOR U8603 ( .A(n6191), .B(\w3[5][58] ), .Z(n6192) );
  XNOR U8604 ( .A(n6193), .B(n6192), .Z(n6194) );
  XOR U8605 ( .A(\w3[5][33] ), .B(n6194), .Z(\w1[6][57] ) );
  XOR U8606 ( .A(\w3[5][51] ), .B(key[826]), .Z(n6197) );
  XNOR U8607 ( .A(n6195), .B(\w3[5][59] ), .Z(n6196) );
  XNOR U8608 ( .A(n6197), .B(n6196), .Z(n6198) );
  XOR U8609 ( .A(\w3[5][34] ), .B(n6198), .Z(\w1[6][58] ) );
  XOR U8610 ( .A(n6199), .B(key[827]), .Z(n6202) );
  XNOR U8611 ( .A(\w3[5][35] ), .B(n6200), .Z(n6201) );
  XNOR U8612 ( .A(n6202), .B(n6201), .Z(\w1[6][59] ) );
  XOR U8613 ( .A(n6203), .B(key[773]), .Z(n6206) );
  XNOR U8614 ( .A(\w3[5][29] ), .B(n6204), .Z(n6205) );
  XNOR U8615 ( .A(n6206), .B(n6205), .Z(\w1[6][5] ) );
  XOR U8616 ( .A(n6207), .B(key[828]), .Z(n6210) );
  XNOR U8617 ( .A(\w3[5][36] ), .B(n6208), .Z(n6209) );
  XNOR U8618 ( .A(n6210), .B(n6209), .Z(\w1[6][60] ) );
  XOR U8619 ( .A(\w3[5][54] ), .B(key[829]), .Z(n6213) );
  XNOR U8620 ( .A(n6211), .B(\w3[5][62] ), .Z(n6212) );
  XNOR U8621 ( .A(n6213), .B(n6212), .Z(n6214) );
  XOR U8622 ( .A(\w3[5][37] ), .B(n6214), .Z(\w1[6][61] ) );
  XOR U8623 ( .A(n6215), .B(key[830]), .Z(n6218) );
  XNOR U8624 ( .A(\w3[5][38] ), .B(n6216), .Z(n6217) );
  XNOR U8625 ( .A(n6218), .B(n6217), .Z(\w1[6][62] ) );
  XOR U8626 ( .A(n6219), .B(key[831]), .Z(n6222) );
  XNOR U8627 ( .A(n6220), .B(\w3[5][39] ), .Z(n6221) );
  XNOR U8628 ( .A(n6222), .B(n6221), .Z(\w1[6][63] ) );
  XOR U8629 ( .A(\w3[5][65] ), .B(\w3[5][89] ), .Z(n6281) );
  XOR U8630 ( .A(n6281), .B(key[832]), .Z(n6224) );
  XOR U8631 ( .A(\w3[5][80] ), .B(\w3[5][88] ), .Z(n6338) );
  XNOR U8632 ( .A(n6338), .B(\w3[5][72] ), .Z(n6223) );
  XNOR U8633 ( .A(n6224), .B(n6223), .Z(\w1[6][64] ) );
  XOR U8634 ( .A(\w3[5][66] ), .B(\w3[5][90] ), .Z(n6285) );
  XOR U8635 ( .A(n6285), .B(key[833]), .Z(n6226) );
  XOR U8636 ( .A(\w3[5][73] ), .B(\w3[5][81] ), .Z(n6309) );
  XNOR U8637 ( .A(\w3[5][89] ), .B(n6309), .Z(n6225) );
  XNOR U8638 ( .A(n6226), .B(n6225), .Z(\w1[6][65] ) );
  XOR U8639 ( .A(\w3[5][67] ), .B(\w3[5][91] ), .Z(n6256) );
  XOR U8640 ( .A(n6256), .B(key[834]), .Z(n6228) );
  XOR U8641 ( .A(\w3[5][74] ), .B(\w3[5][82] ), .Z(n6317) );
  XNOR U8642 ( .A(\w3[5][90] ), .B(n6317), .Z(n6227) );
  XNOR U8643 ( .A(n6228), .B(n6227), .Z(\w1[6][66] ) );
  XOR U8644 ( .A(\w3[5][68] ), .B(\w3[5][64] ), .Z(n6258) );
  XOR U8645 ( .A(n6258), .B(key[835]), .Z(n6231) );
  XOR U8646 ( .A(\w3[5][75] ), .B(\w3[5][83] ), .Z(n6284) );
  XNOR U8647 ( .A(\w3[5][88] ), .B(n6284), .Z(n6229) );
  XNOR U8648 ( .A(\w3[5][92] ), .B(n6229), .Z(n6322) );
  XNOR U8649 ( .A(\w3[5][91] ), .B(n6322), .Z(n6230) );
  XNOR U8650 ( .A(n6231), .B(n6230), .Z(\w1[6][67] ) );
  XOR U8651 ( .A(\w3[5][64] ), .B(\w3[5][69] ), .Z(n6263) );
  XOR U8652 ( .A(n6263), .B(key[836]), .Z(n6235) );
  XOR U8653 ( .A(\w3[5][84] ), .B(\w3[5][93] ), .Z(n6233) );
  XNOR U8654 ( .A(\w3[5][88] ), .B(\w3[5][76] ), .Z(n6232) );
  XNOR U8655 ( .A(n6233), .B(n6232), .Z(n6326) );
  XNOR U8656 ( .A(\w3[5][92] ), .B(n6326), .Z(n6234) );
  XNOR U8657 ( .A(n6235), .B(n6234), .Z(\w1[6][68] ) );
  XOR U8658 ( .A(\w3[5][70] ), .B(\w3[5][94] ), .Z(n6269) );
  XOR U8659 ( .A(n6269), .B(key[837]), .Z(n6237) );
  XOR U8660 ( .A(\w3[5][77] ), .B(\w3[5][85] ), .Z(n6329) );
  XNOR U8661 ( .A(\w3[5][93] ), .B(n6329), .Z(n6236) );
  XNOR U8662 ( .A(n6237), .B(n6236), .Z(\w1[6][69] ) );
  XOR U8663 ( .A(n6238), .B(key[774]), .Z(n6241) );
  XNOR U8664 ( .A(n6239), .B(\w3[5][30] ), .Z(n6240) );
  XNOR U8665 ( .A(n6241), .B(n6240), .Z(\w1[6][6] ) );
  XOR U8666 ( .A(\w3[5][64] ), .B(\w3[5][71] ), .Z(n6270) );
  XOR U8667 ( .A(n6270), .B(key[838]), .Z(n6243) );
  XOR U8668 ( .A(\w3[5][78] ), .B(\w3[5][86] ), .Z(n6295) );
  XNOR U8669 ( .A(\w3[5][88] ), .B(\w3[5][95] ), .Z(n6245) );
  XNOR U8670 ( .A(n6295), .B(n6245), .Z(n6334) );
  XNOR U8671 ( .A(\w3[5][94] ), .B(n6334), .Z(n6242) );
  XNOR U8672 ( .A(n6243), .B(n6242), .Z(\w1[6][70] ) );
  XOR U8673 ( .A(\w3[5][79] ), .B(\w3[5][87] ), .Z(n6337) );
  XNOR U8674 ( .A(n6337), .B(key[839]), .Z(n6244) );
  XNOR U8675 ( .A(n6245), .B(n6244), .Z(n6246) );
  XNOR U8676 ( .A(\w3[5][64] ), .B(n6246), .Z(\w1[6][71] ) );
  XOR U8677 ( .A(\w3[5][64] ), .B(key[840]), .Z(n6248) );
  XNOR U8678 ( .A(\w3[5][65] ), .B(\w3[5][73] ), .Z(n6247) );
  XNOR U8679 ( .A(n6248), .B(n6247), .Z(n6249) );
  XOR U8680 ( .A(n6338), .B(n6249), .Z(\w1[6][72] ) );
  XOR U8681 ( .A(\w3[5][74] ), .B(key[841]), .Z(n6251) );
  XNOR U8682 ( .A(\w3[5][81] ), .B(\w3[5][66] ), .Z(n6250) );
  XNOR U8683 ( .A(n6251), .B(n6250), .Z(n6252) );
  XOR U8684 ( .A(n6281), .B(n6252), .Z(\w1[6][73] ) );
  XOR U8685 ( .A(\w3[5][75] ), .B(key[842]), .Z(n6254) );
  XNOR U8686 ( .A(\w3[5][82] ), .B(\w3[5][67] ), .Z(n6253) );
  XNOR U8687 ( .A(n6254), .B(n6253), .Z(n6255) );
  XOR U8688 ( .A(n6285), .B(n6255), .Z(\w1[6][74] ) );
  XNOR U8689 ( .A(\w3[5][72] ), .B(n6256), .Z(n6257) );
  XNOR U8690 ( .A(\w3[5][76] ), .B(n6257), .Z(n6288) );
  XOR U8691 ( .A(n6288), .B(key[843]), .Z(n6260) );
  XNOR U8692 ( .A(\w3[5][83] ), .B(n6258), .Z(n6259) );
  XNOR U8693 ( .A(n6260), .B(n6259), .Z(\w1[6][75] ) );
  XOR U8694 ( .A(\w3[5][68] ), .B(\w3[5][77] ), .Z(n6262) );
  XNOR U8695 ( .A(\w3[5][72] ), .B(\w3[5][92] ), .Z(n6261) );
  XNOR U8696 ( .A(n6262), .B(n6261), .Z(n6291) );
  XOR U8697 ( .A(n6291), .B(key[844]), .Z(n6265) );
  XNOR U8698 ( .A(\w3[5][84] ), .B(n6263), .Z(n6264) );
  XNOR U8699 ( .A(n6265), .B(n6264), .Z(\w1[6][76] ) );
  XOR U8700 ( .A(\w3[5][93] ), .B(\w3[5][69] ), .Z(n6294) );
  XOR U8701 ( .A(n6294), .B(key[845]), .Z(n6267) );
  XNOR U8702 ( .A(\w3[5][70] ), .B(\w3[5][78] ), .Z(n6266) );
  XNOR U8703 ( .A(n6267), .B(n6266), .Z(n6268) );
  XOR U8704 ( .A(\w3[5][85] ), .B(n6268), .Z(\w1[6][77] ) );
  XNOR U8705 ( .A(\w3[5][72] ), .B(\w3[5][79] ), .Z(n6303) );
  XNOR U8706 ( .A(n6269), .B(n6303), .Z(n6298) );
  XOR U8707 ( .A(n6298), .B(key[846]), .Z(n6272) );
  XNOR U8708 ( .A(\w3[5][86] ), .B(n6270), .Z(n6271) );
  XNOR U8709 ( .A(n6272), .B(n6271), .Z(\w1[6][78] ) );
  XOR U8710 ( .A(\w3[5][95] ), .B(\w3[5][71] ), .Z(n6301) );
  XOR U8711 ( .A(n6301), .B(key[847]), .Z(n6274) );
  XOR U8712 ( .A(\w3[5][72] ), .B(\w3[5][64] ), .Z(n6305) );
  XNOR U8713 ( .A(\w3[5][87] ), .B(n6305), .Z(n6273) );
  XNOR U8714 ( .A(n6274), .B(n6273), .Z(\w1[6][79] ) );
  XNOR U8715 ( .A(n6275), .B(key[775]), .Z(n6276) );
  XNOR U8716 ( .A(n6277), .B(n6276), .Z(n6278) );
  XNOR U8717 ( .A(\w3[5][0] ), .B(n6278), .Z(\w1[6][7] ) );
  XOR U8718 ( .A(n6305), .B(key[848]), .Z(n6280) );
  XNOR U8719 ( .A(\w3[5][88] ), .B(n6309), .Z(n6279) );
  XNOR U8720 ( .A(n6280), .B(n6279), .Z(\w1[6][80] ) );
  XOR U8721 ( .A(n6317), .B(key[849]), .Z(n6283) );
  XNOR U8722 ( .A(n6281), .B(\w3[5][73] ), .Z(n6282) );
  XNOR U8723 ( .A(n6283), .B(n6282), .Z(\w1[6][81] ) );
  XOR U8724 ( .A(n6284), .B(key[850]), .Z(n6287) );
  XNOR U8725 ( .A(n6285), .B(\w3[5][74] ), .Z(n6286) );
  XNOR U8726 ( .A(n6287), .B(n6286), .Z(\w1[6][82] ) );
  XOR U8727 ( .A(\w3[5][80] ), .B(\w3[5][84] ), .Z(n6321) );
  XOR U8728 ( .A(n6321), .B(key[851]), .Z(n6290) );
  XNOR U8729 ( .A(\w3[5][75] ), .B(n6288), .Z(n6289) );
  XNOR U8730 ( .A(n6290), .B(n6289), .Z(\w1[6][83] ) );
  XOR U8731 ( .A(\w3[5][80] ), .B(\w3[5][85] ), .Z(n6325) );
  XOR U8732 ( .A(n6325), .B(key[852]), .Z(n6293) );
  XNOR U8733 ( .A(\w3[5][76] ), .B(n6291), .Z(n6292) );
  XNOR U8734 ( .A(n6293), .B(n6292), .Z(\w1[6][84] ) );
  XOR U8735 ( .A(n6294), .B(key[853]), .Z(n6297) );
  XNOR U8736 ( .A(\w3[5][77] ), .B(n6295), .Z(n6296) );
  XNOR U8737 ( .A(n6297), .B(n6296), .Z(\w1[6][85] ) );
  XOR U8738 ( .A(\w3[5][80] ), .B(\w3[5][87] ), .Z(n6333) );
  XOR U8739 ( .A(n6333), .B(key[854]), .Z(n6300) );
  XNOR U8740 ( .A(\w3[5][78] ), .B(n6298), .Z(n6299) );
  XNOR U8741 ( .A(n6300), .B(n6299), .Z(\w1[6][86] ) );
  XNOR U8742 ( .A(n6301), .B(key[855]), .Z(n6302) );
  XNOR U8743 ( .A(n6303), .B(n6302), .Z(n6304) );
  XNOR U8744 ( .A(\w3[5][80] ), .B(n6304), .Z(\w1[6][87] ) );
  XOR U8745 ( .A(n6305), .B(key[856]), .Z(n6307) );
  XNOR U8746 ( .A(\w3[5][80] ), .B(\w3[5][81] ), .Z(n6306) );
  XNOR U8747 ( .A(n6307), .B(n6306), .Z(n6308) );
  XOR U8748 ( .A(\w3[5][89] ), .B(n6308), .Z(\w1[6][88] ) );
  XOR U8749 ( .A(\w3[5][82] ), .B(key[857]), .Z(n6311) );
  XNOR U8750 ( .A(n6309), .B(\w3[5][90] ), .Z(n6310) );
  XNOR U8751 ( .A(n6311), .B(n6310), .Z(n6312) );
  XOR U8752 ( .A(\w3[5][65] ), .B(n6312), .Z(\w1[6][89] ) );
  XOR U8753 ( .A(\w3[5][9] ), .B(key[776]), .Z(n6314) );
  XNOR U8754 ( .A(\w3[5][1] ), .B(\w3[5][0] ), .Z(n6313) );
  XNOR U8755 ( .A(n6314), .B(n6313), .Z(n6315) );
  XOR U8756 ( .A(n6316), .B(n6315), .Z(\w1[6][8] ) );
  XOR U8757 ( .A(\w3[5][83] ), .B(key[858]), .Z(n6319) );
  XNOR U8758 ( .A(n6317), .B(\w3[5][91] ), .Z(n6318) );
  XNOR U8759 ( .A(n6319), .B(n6318), .Z(n6320) );
  XOR U8760 ( .A(\w3[5][66] ), .B(n6320), .Z(\w1[6][90] ) );
  XOR U8761 ( .A(n6321), .B(key[859]), .Z(n6324) );
  XNOR U8762 ( .A(\w3[5][67] ), .B(n6322), .Z(n6323) );
  XNOR U8763 ( .A(n6324), .B(n6323), .Z(\w1[6][91] ) );
  XOR U8764 ( .A(n6325), .B(key[860]), .Z(n6328) );
  XNOR U8765 ( .A(\w3[5][68] ), .B(n6326), .Z(n6327) );
  XNOR U8766 ( .A(n6328), .B(n6327), .Z(\w1[6][92] ) );
  XOR U8767 ( .A(\w3[5][86] ), .B(key[861]), .Z(n6331) );
  XNOR U8768 ( .A(n6329), .B(\w3[5][94] ), .Z(n6330) );
  XNOR U8769 ( .A(n6331), .B(n6330), .Z(n6332) );
  XOR U8770 ( .A(\w3[5][69] ), .B(n6332), .Z(\w1[6][93] ) );
  XOR U8771 ( .A(n6333), .B(key[862]), .Z(n6336) );
  XNOR U8772 ( .A(\w3[5][70] ), .B(n6334), .Z(n6335) );
  XNOR U8773 ( .A(n6336), .B(n6335), .Z(\w1[6][94] ) );
  XOR U8774 ( .A(n6337), .B(key[863]), .Z(n6340) );
  XNOR U8775 ( .A(n6338), .B(\w3[5][71] ), .Z(n6339) );
  XNOR U8776 ( .A(n6340), .B(n6339), .Z(\w1[6][95] ) );
  XOR U8777 ( .A(\w3[5][104] ), .B(key[864]), .Z(n6344) );
  XNOR U8778 ( .A(n6342), .B(n6341), .Z(n6343) );
  XNOR U8779 ( .A(n6344), .B(n6343), .Z(\w1[6][96] ) );
  XOR U8780 ( .A(n6345), .B(key[865]), .Z(n6348) );
  XNOR U8781 ( .A(\w3[5][121] ), .B(n6346), .Z(n6347) );
  XNOR U8782 ( .A(n6348), .B(n6347), .Z(\w1[6][97] ) );
  XOR U8783 ( .A(n6349), .B(key[866]), .Z(n6352) );
  XNOR U8784 ( .A(\w3[5][122] ), .B(n6350), .Z(n6351) );
  XNOR U8785 ( .A(n6352), .B(n6351), .Z(\w1[6][98] ) );
  XOR U8786 ( .A(n6353), .B(key[867]), .Z(n6356) );
  XNOR U8787 ( .A(n6354), .B(\w3[5][123] ), .Z(n6355) );
  XNOR U8788 ( .A(n6356), .B(n6355), .Z(\w1[6][99] ) );
  XOR U8789 ( .A(\w3[5][10] ), .B(key[777]), .Z(n6358) );
  XNOR U8790 ( .A(\w3[5][2] ), .B(\w3[5][17] ), .Z(n6357) );
  XNOR U8791 ( .A(n6358), .B(n6357), .Z(n6359) );
  XOR U8792 ( .A(n6360), .B(n6359), .Z(\w1[6][9] ) );
  XOR U8793 ( .A(\w3[6][8] ), .B(key[896]), .Z(n6362) );
  XOR U8794 ( .A(\w3[6][1] ), .B(\w3[6][25] ), .Z(n6784) );
  XOR U8795 ( .A(\w3[6][16] ), .B(\w3[6][24] ), .Z(n6740) );
  XNOR U8796 ( .A(n6784), .B(n6740), .Z(n6361) );
  XNOR U8797 ( .A(n6362), .B(n6361), .Z(\w1[7][0] ) );
  XOR U8798 ( .A(\w3[6][96] ), .B(\w3[6][101] ), .Z(n6387) );
  XOR U8799 ( .A(n6387), .B(key[996]), .Z(n6366) );
  XOR U8800 ( .A(\w3[6][116] ), .B(\w3[6][125] ), .Z(n6364) );
  XNOR U8801 ( .A(\w3[6][120] ), .B(\w3[6][108] ), .Z(n6363) );
  XNOR U8802 ( .A(n6364), .B(n6363), .Z(n6445) );
  XNOR U8803 ( .A(\w3[6][124] ), .B(n6445), .Z(n6365) );
  XNOR U8804 ( .A(n6366), .B(n6365), .Z(\w1[7][100] ) );
  XOR U8805 ( .A(\w3[6][102] ), .B(\w3[6][126] ), .Z(n6396) );
  XOR U8806 ( .A(n6396), .B(key[997]), .Z(n6368) );
  XOR U8807 ( .A(\w3[6][109] ), .B(\w3[6][117] ), .Z(n6448) );
  XNOR U8808 ( .A(\w3[6][125] ), .B(n6448), .Z(n6367) );
  XNOR U8809 ( .A(n6368), .B(n6367), .Z(\w1[7][101] ) );
  XOR U8810 ( .A(\w3[6][96] ), .B(\w3[6][103] ), .Z(n6397) );
  XOR U8811 ( .A(n6397), .B(key[998]), .Z(n6370) );
  XOR U8812 ( .A(\w3[6][110] ), .B(\w3[6][118] ), .Z(n6415) );
  XNOR U8813 ( .A(\w3[6][120] ), .B(\w3[6][127] ), .Z(n6372) );
  XNOR U8814 ( .A(n6415), .B(n6372), .Z(n6453) );
  XNOR U8815 ( .A(\w3[6][126] ), .B(n6453), .Z(n6369) );
  XNOR U8816 ( .A(n6370), .B(n6369), .Z(\w1[7][102] ) );
  XOR U8817 ( .A(\w3[6][111] ), .B(\w3[6][119] ), .Z(n6456) );
  XNOR U8818 ( .A(n6456), .B(key[999]), .Z(n6371) );
  XNOR U8819 ( .A(n6372), .B(n6371), .Z(n6373) );
  XNOR U8820 ( .A(\w3[6][96] ), .B(n6373), .Z(\w1[7][103] ) );
  XOR U8821 ( .A(\w3[6][105] ), .B(\w3[6][97] ), .Z(n6435) );
  XOR U8822 ( .A(n6435), .B(key[1000]), .Z(n6375) );
  XOR U8823 ( .A(\w3[6][120] ), .B(\w3[6][112] ), .Z(n6766) );
  XNOR U8824 ( .A(\w3[6][96] ), .B(n6766), .Z(n6374) );
  XNOR U8825 ( .A(n6375), .B(n6374), .Z(\w1[7][104] ) );
  XOR U8826 ( .A(\w3[6][106] ), .B(\w3[6][113] ), .Z(n6377) );
  XOR U8827 ( .A(\w3[6][97] ), .B(\w3[6][121] ), .Z(n6765) );
  XNOR U8828 ( .A(n6765), .B(key[1001]), .Z(n6376) );
  XNOR U8829 ( .A(n6377), .B(n6376), .Z(n6378) );
  XOR U8830 ( .A(\w3[6][98] ), .B(n6378), .Z(\w1[7][105] ) );
  XOR U8831 ( .A(\w3[6][107] ), .B(\w3[6][114] ), .Z(n6380) );
  XOR U8832 ( .A(\w3[6][98] ), .B(\w3[6][122] ), .Z(n6770) );
  XNOR U8833 ( .A(n6770), .B(key[1002]), .Z(n6379) );
  XNOR U8834 ( .A(n6380), .B(n6379), .Z(n6381) );
  XOR U8835 ( .A(\w3[6][99] ), .B(n6381), .Z(\w1[7][106] ) );
  XOR U8836 ( .A(\w3[6][99] ), .B(\w3[6][123] ), .Z(n6774) );
  XNOR U8837 ( .A(\w3[6][108] ), .B(n6774), .Z(n6382) );
  XNOR U8838 ( .A(\w3[6][104] ), .B(n6382), .Z(n6408) );
  XOR U8839 ( .A(n6408), .B(key[1003]), .Z(n6384) );
  XOR U8840 ( .A(\w3[6][96] ), .B(\w3[6][100] ), .Z(n6778) );
  XNOR U8841 ( .A(\w3[6][115] ), .B(n6778), .Z(n6383) );
  XNOR U8842 ( .A(n6384), .B(n6383), .Z(\w1[7][107] ) );
  XOR U8843 ( .A(\w3[6][100] ), .B(\w3[6][104] ), .Z(n6386) );
  XNOR U8844 ( .A(\w3[6][124] ), .B(\w3[6][109] ), .Z(n6385) );
  XNOR U8845 ( .A(n6386), .B(n6385), .Z(n6411) );
  XOR U8846 ( .A(n6411), .B(key[1004]), .Z(n6389) );
  XNOR U8847 ( .A(\w3[6][116] ), .B(n6387), .Z(n6388) );
  XNOR U8848 ( .A(n6389), .B(n6388), .Z(\w1[7][108] ) );
  XOR U8849 ( .A(\w3[6][125] ), .B(\w3[6][101] ), .Z(n6414) );
  XOR U8850 ( .A(n6414), .B(key[1005]), .Z(n6391) );
  XNOR U8851 ( .A(\w3[6][102] ), .B(\w3[6][110] ), .Z(n6390) );
  XNOR U8852 ( .A(n6391), .B(n6390), .Z(n6392) );
  XOR U8853 ( .A(\w3[6][117] ), .B(n6392), .Z(\w1[7][109] ) );
  XOR U8854 ( .A(\w3[6][11] ), .B(\w3[6][18] ), .Z(n6394) );
  XOR U8855 ( .A(\w3[6][2] ), .B(\w3[6][26] ), .Z(n6479) );
  XNOR U8856 ( .A(n6479), .B(key[906]), .Z(n6393) );
  XNOR U8857 ( .A(n6394), .B(n6393), .Z(n6395) );
  XOR U8858 ( .A(\w3[6][3] ), .B(n6395), .Z(\w1[7][10] ) );
  XNOR U8859 ( .A(\w3[6][111] ), .B(\w3[6][104] ), .Z(n6423) );
  XNOR U8860 ( .A(n6396), .B(n6423), .Z(n6418) );
  XOR U8861 ( .A(n6418), .B(key[1006]), .Z(n6399) );
  XNOR U8862 ( .A(\w3[6][118] ), .B(n6397), .Z(n6398) );
  XNOR U8863 ( .A(n6399), .B(n6398), .Z(\w1[7][110] ) );
  XOR U8864 ( .A(\w3[6][127] ), .B(\w3[6][103] ), .Z(n6421) );
  XOR U8865 ( .A(n6421), .B(key[1007]), .Z(n6401) );
  XOR U8866 ( .A(\w3[6][96] ), .B(\w3[6][104] ), .Z(n6428) );
  XNOR U8867 ( .A(\w3[6][119] ), .B(n6428), .Z(n6400) );
  XNOR U8868 ( .A(n6401), .B(n6400), .Z(\w1[7][111] ) );
  XOR U8869 ( .A(\w3[6][105] ), .B(\w3[6][113] ), .Z(n6769) );
  XOR U8870 ( .A(n6769), .B(key[1008]), .Z(n6403) );
  XNOR U8871 ( .A(\w3[6][120] ), .B(n6428), .Z(n6402) );
  XNOR U8872 ( .A(n6403), .B(n6402), .Z(\w1[7][112] ) );
  XOR U8873 ( .A(\w3[6][106] ), .B(\w3[6][114] ), .Z(n6773) );
  XOR U8874 ( .A(n6773), .B(key[1009]), .Z(n6405) );
  XNOR U8875 ( .A(n6435), .B(\w3[6][121] ), .Z(n6404) );
  XNOR U8876 ( .A(n6405), .B(n6404), .Z(\w1[7][113] ) );
  XOR U8877 ( .A(\w3[6][107] ), .B(\w3[6][115] ), .Z(n6440) );
  XOR U8878 ( .A(n6440), .B(key[1010]), .Z(n6407) );
  XNOR U8879 ( .A(\w3[6][106] ), .B(n6770), .Z(n6406) );
  XNOR U8880 ( .A(n6407), .B(n6406), .Z(\w1[7][114] ) );
  XOR U8881 ( .A(\w3[6][116] ), .B(\w3[6][112] ), .Z(n6441) );
  XOR U8882 ( .A(n6441), .B(key[1011]), .Z(n6410) );
  XNOR U8883 ( .A(\w3[6][107] ), .B(n6408), .Z(n6409) );
  XNOR U8884 ( .A(n6410), .B(n6409), .Z(\w1[7][115] ) );
  XOR U8885 ( .A(\w3[6][117] ), .B(\w3[6][112] ), .Z(n6444) );
  XOR U8886 ( .A(n6444), .B(key[1012]), .Z(n6413) );
  XNOR U8887 ( .A(\w3[6][108] ), .B(n6411), .Z(n6412) );
  XNOR U8888 ( .A(n6413), .B(n6412), .Z(\w1[7][116] ) );
  XOR U8889 ( .A(n6414), .B(key[1013]), .Z(n6417) );
  XNOR U8890 ( .A(\w3[6][109] ), .B(n6415), .Z(n6416) );
  XNOR U8891 ( .A(n6417), .B(n6416), .Z(\w1[7][117] ) );
  XOR U8892 ( .A(\w3[6][119] ), .B(\w3[6][112] ), .Z(n6452) );
  XOR U8893 ( .A(n6452), .B(key[1014]), .Z(n6420) );
  XNOR U8894 ( .A(\w3[6][110] ), .B(n6418), .Z(n6419) );
  XNOR U8895 ( .A(n6420), .B(n6419), .Z(\w1[7][118] ) );
  XNOR U8896 ( .A(n6421), .B(key[1015]), .Z(n6422) );
  XNOR U8897 ( .A(n6423), .B(n6422), .Z(n6424) );
  XNOR U8898 ( .A(\w3[6][112] ), .B(n6424), .Z(\w1[7][119] ) );
  XOR U8899 ( .A(\w3[6][3] ), .B(\w3[6][27] ), .Z(n6520) );
  XNOR U8900 ( .A(\w3[6][8] ), .B(\w3[6][12] ), .Z(n6425) );
  XNOR U8901 ( .A(n6520), .B(n6425), .Z(n6476) );
  XOR U8902 ( .A(n6476), .B(key[907]), .Z(n6427) );
  XOR U8903 ( .A(\w3[6][0] ), .B(\w3[6][4] ), .Z(n6550) );
  XNOR U8904 ( .A(\w3[6][19] ), .B(n6550), .Z(n6426) );
  XNOR U8905 ( .A(n6427), .B(n6426), .Z(\w1[7][11] ) );
  XOR U8906 ( .A(n6428), .B(key[1016]), .Z(n6430) );
  XNOR U8907 ( .A(\w3[6][121] ), .B(\w3[6][113] ), .Z(n6429) );
  XNOR U8908 ( .A(n6430), .B(n6429), .Z(n6431) );
  XOR U8909 ( .A(\w3[6][112] ), .B(n6431), .Z(\w1[7][120] ) );
  XOR U8910 ( .A(\w3[6][114] ), .B(key[1017]), .Z(n6433) );
  XNOR U8911 ( .A(\w3[6][113] ), .B(\w3[6][122] ), .Z(n6432) );
  XNOR U8912 ( .A(n6433), .B(n6432), .Z(n6434) );
  XOR U8913 ( .A(n6435), .B(n6434), .Z(\w1[7][121] ) );
  XOR U8914 ( .A(n6773), .B(key[1018]), .Z(n6437) );
  XNOR U8915 ( .A(\w3[6][115] ), .B(\w3[6][123] ), .Z(n6436) );
  XNOR U8916 ( .A(n6437), .B(n6436), .Z(n6438) );
  XOR U8917 ( .A(\w3[6][98] ), .B(n6438), .Z(\w1[7][122] ) );
  XNOR U8918 ( .A(\w3[6][124] ), .B(\w3[6][120] ), .Z(n6439) );
  XNOR U8919 ( .A(n6440), .B(n6439), .Z(n6777) );
  XOR U8920 ( .A(n6777), .B(key[1019]), .Z(n6443) );
  XNOR U8921 ( .A(\w3[6][99] ), .B(n6441), .Z(n6442) );
  XNOR U8922 ( .A(n6443), .B(n6442), .Z(\w1[7][123] ) );
  XOR U8923 ( .A(n6444), .B(key[1020]), .Z(n6447) );
  XNOR U8924 ( .A(n6445), .B(\w3[6][100] ), .Z(n6446) );
  XNOR U8925 ( .A(n6447), .B(n6446), .Z(\w1[7][124] ) );
  XOR U8926 ( .A(\w3[6][118] ), .B(key[1021]), .Z(n6450) );
  XNOR U8927 ( .A(n6448), .B(\w3[6][126] ), .Z(n6449) );
  XNOR U8928 ( .A(n6450), .B(n6449), .Z(n6451) );
  XOR U8929 ( .A(\w3[6][101] ), .B(n6451), .Z(\w1[7][125] ) );
  XOR U8930 ( .A(n6452), .B(key[1022]), .Z(n6455) );
  XNOR U8931 ( .A(\w3[6][102] ), .B(n6453), .Z(n6454) );
  XNOR U8932 ( .A(n6455), .B(n6454), .Z(\w1[7][126] ) );
  XOR U8933 ( .A(n6766), .B(key[1023]), .Z(n6458) );
  XNOR U8934 ( .A(\w3[6][103] ), .B(n6456), .Z(n6457) );
  XNOR U8935 ( .A(n6458), .B(n6457), .Z(\w1[7][127] ) );
  XOR U8936 ( .A(\w3[6][13] ), .B(\w3[6][28] ), .Z(n6460) );
  XNOR U8937 ( .A(\w3[6][8] ), .B(\w3[6][4] ), .Z(n6459) );
  XNOR U8938 ( .A(n6460), .B(n6459), .Z(n6482) );
  XOR U8939 ( .A(n6482), .B(key[908]), .Z(n6462) );
  XOR U8940 ( .A(\w3[6][0] ), .B(\w3[6][5] ), .Z(n6587) );
  XNOR U8941 ( .A(\w3[6][20] ), .B(n6587), .Z(n6461) );
  XNOR U8942 ( .A(n6462), .B(n6461), .Z(\w1[7][12] ) );
  XOR U8943 ( .A(\w3[6][14] ), .B(\w3[6][21] ), .Z(n6464) );
  XOR U8944 ( .A(\w3[6][5] ), .B(\w3[6][29] ), .Z(n6485) );
  XNOR U8945 ( .A(n6485), .B(key[909]), .Z(n6463) );
  XNOR U8946 ( .A(n6464), .B(n6463), .Z(n6465) );
  XOR U8947 ( .A(\w3[6][6] ), .B(n6465), .Z(\w1[7][13] ) );
  XOR U8948 ( .A(\w3[6][6] ), .B(\w3[6][30] ), .Z(n6628) );
  XNOR U8949 ( .A(\w3[6][8] ), .B(\w3[6][15] ), .Z(n6493) );
  XNOR U8950 ( .A(n6628), .B(n6493), .Z(n6488) );
  XOR U8951 ( .A(n6488), .B(key[910]), .Z(n6467) );
  XOR U8952 ( .A(\w3[6][0] ), .B(\w3[6][7] ), .Z(n6663) );
  XNOR U8953 ( .A(\w3[6][22] ), .B(n6663), .Z(n6466) );
  XNOR U8954 ( .A(n6467), .B(n6466), .Z(\w1[7][14] ) );
  XOR U8955 ( .A(\w3[6][7] ), .B(\w3[6][31] ), .Z(n6491) );
  XOR U8956 ( .A(n6491), .B(key[911]), .Z(n6469) );
  XOR U8957 ( .A(\w3[6][8] ), .B(\w3[6][0] ), .Z(n6495) );
  XNOR U8958 ( .A(\w3[6][23] ), .B(n6495), .Z(n6468) );
  XNOR U8959 ( .A(n6469), .B(n6468), .Z(\w1[7][15] ) );
  XOR U8960 ( .A(\w3[6][17] ), .B(\w3[6][9] ), .Z(n6499) );
  XOR U8961 ( .A(n6499), .B(key[912]), .Z(n6471) );
  XNOR U8962 ( .A(\w3[6][24] ), .B(n6495), .Z(n6470) );
  XNOR U8963 ( .A(n6471), .B(n6470), .Z(\w1[7][16] ) );
  XOR U8964 ( .A(\w3[6][18] ), .B(\w3[6][10] ), .Z(n6519) );
  XOR U8965 ( .A(n6519), .B(key[913]), .Z(n6473) );
  XNOR U8966 ( .A(n6784), .B(\w3[6][9] ), .Z(n6472) );
  XNOR U8967 ( .A(n6473), .B(n6472), .Z(\w1[7][17] ) );
  XOR U8968 ( .A(\w3[6][11] ), .B(\w3[6][19] ), .Z(n6507) );
  XOR U8969 ( .A(n6507), .B(key[914]), .Z(n6475) );
  XNOR U8970 ( .A(n6479), .B(\w3[6][10] ), .Z(n6474) );
  XNOR U8971 ( .A(n6475), .B(n6474), .Z(\w1[7][18] ) );
  XOR U8972 ( .A(\w3[6][16] ), .B(\w3[6][20] ), .Z(n6508) );
  XOR U8973 ( .A(n6508), .B(key[915]), .Z(n6478) );
  XNOR U8974 ( .A(\w3[6][11] ), .B(n6476), .Z(n6477) );
  XNOR U8975 ( .A(n6478), .B(n6477), .Z(\w1[7][19] ) );
  XOR U8976 ( .A(n6499), .B(key[897]), .Z(n6481) );
  XNOR U8977 ( .A(\w3[6][25] ), .B(n6479), .Z(n6480) );
  XNOR U8978 ( .A(n6481), .B(n6480), .Z(\w1[7][1] ) );
  XOR U8979 ( .A(\w3[6][16] ), .B(\w3[6][21] ), .Z(n6513) );
  XOR U8980 ( .A(n6513), .B(key[916]), .Z(n6484) );
  XNOR U8981 ( .A(\w3[6][12] ), .B(n6482), .Z(n6483) );
  XNOR U8982 ( .A(n6484), .B(n6483), .Z(\w1[7][20] ) );
  XOR U8983 ( .A(\w3[6][14] ), .B(\w3[6][22] ), .Z(n6523) );
  XOR U8984 ( .A(n6523), .B(key[917]), .Z(n6487) );
  XNOR U8985 ( .A(\w3[6][13] ), .B(n6485), .Z(n6486) );
  XNOR U8986 ( .A(n6487), .B(n6486), .Z(\w1[7][21] ) );
  XOR U8987 ( .A(\w3[6][16] ), .B(\w3[6][23] ), .Z(n6524) );
  XOR U8988 ( .A(n6524), .B(key[918]), .Z(n6490) );
  XNOR U8989 ( .A(\w3[6][14] ), .B(n6488), .Z(n6489) );
  XNOR U8990 ( .A(n6490), .B(n6489), .Z(\w1[7][22] ) );
  XNOR U8991 ( .A(n6491), .B(key[919]), .Z(n6492) );
  XNOR U8992 ( .A(n6493), .B(n6492), .Z(n6494) );
  XNOR U8993 ( .A(\w3[6][16] ), .B(n6494), .Z(\w1[7][23] ) );
  XOR U8994 ( .A(\w3[6][17] ), .B(key[920]), .Z(n6497) );
  XNOR U8995 ( .A(\w3[6][25] ), .B(n6495), .Z(n6496) );
  XNOR U8996 ( .A(n6497), .B(n6496), .Z(n6498) );
  XOR U8997 ( .A(\w3[6][16] ), .B(n6498), .Z(\w1[7][24] ) );
  XOR U8998 ( .A(n6499), .B(key[921]), .Z(n6501) );
  XNOR U8999 ( .A(\w3[6][1] ), .B(\w3[6][26] ), .Z(n6500) );
  XNOR U9000 ( .A(n6501), .B(n6500), .Z(n6502) );
  XOR U9001 ( .A(\w3[6][18] ), .B(n6502), .Z(\w1[7][25] ) );
  XOR U9002 ( .A(n6519), .B(key[922]), .Z(n6504) );
  XNOR U9003 ( .A(\w3[6][2] ), .B(\w3[6][19] ), .Z(n6503) );
  XNOR U9004 ( .A(n6504), .B(n6503), .Z(n6505) );
  XOR U9005 ( .A(\w3[6][27] ), .B(n6505), .Z(\w1[7][26] ) );
  XNOR U9006 ( .A(\w3[6][24] ), .B(\w3[6][28] ), .Z(n6506) );
  XNOR U9007 ( .A(n6507), .B(n6506), .Z(n6549) );
  XOR U9008 ( .A(n6549), .B(key[923]), .Z(n6510) );
  XNOR U9009 ( .A(\w3[6][3] ), .B(n6508), .Z(n6509) );
  XNOR U9010 ( .A(n6510), .B(n6509), .Z(\w1[7][27] ) );
  XOR U9011 ( .A(\w3[6][20] ), .B(\w3[6][29] ), .Z(n6512) );
  XNOR U9012 ( .A(\w3[6][24] ), .B(\w3[6][12] ), .Z(n6511) );
  XNOR U9013 ( .A(n6512), .B(n6511), .Z(n6586) );
  XOR U9014 ( .A(n6586), .B(key[924]), .Z(n6515) );
  XNOR U9015 ( .A(\w3[6][4] ), .B(n6513), .Z(n6514) );
  XNOR U9016 ( .A(n6515), .B(n6514), .Z(\w1[7][28] ) );
  XOR U9017 ( .A(\w3[6][13] ), .B(\w3[6][21] ), .Z(n6627) );
  XOR U9018 ( .A(n6627), .B(key[925]), .Z(n6517) );
  XNOR U9019 ( .A(\w3[6][22] ), .B(\w3[6][30] ), .Z(n6516) );
  XNOR U9020 ( .A(n6517), .B(n6516), .Z(n6518) );
  XOR U9021 ( .A(\w3[6][5] ), .B(n6518), .Z(\w1[7][29] ) );
  XOR U9022 ( .A(n6519), .B(key[898]), .Z(n6522) );
  XNOR U9023 ( .A(\w3[6][26] ), .B(n6520), .Z(n6521) );
  XNOR U9024 ( .A(n6522), .B(n6521), .Z(\w1[7][2] ) );
  XNOR U9025 ( .A(\w3[6][24] ), .B(\w3[6][31] ), .Z(n6701) );
  XNOR U9026 ( .A(n6523), .B(n6701), .Z(n6662) );
  XOR U9027 ( .A(n6662), .B(key[926]), .Z(n6526) );
  XNOR U9028 ( .A(\w3[6][6] ), .B(n6524), .Z(n6525) );
  XNOR U9029 ( .A(n6526), .B(n6525), .Z(\w1[7][30] ) );
  XOR U9030 ( .A(\w3[6][15] ), .B(\w3[6][23] ), .Z(n6699) );
  XOR U9031 ( .A(n6699), .B(key[927]), .Z(n6528) );
  XNOR U9032 ( .A(n6740), .B(\w3[6][7] ), .Z(n6527) );
  XNOR U9033 ( .A(n6528), .B(n6527), .Z(\w1[7][31] ) );
  XOR U9034 ( .A(\w3[6][33] ), .B(\w3[6][57] ), .Z(n6583) );
  XOR U9035 ( .A(n6583), .B(key[928]), .Z(n6530) );
  XOR U9036 ( .A(\w3[6][48] ), .B(\w3[6][56] ), .Z(n6644) );
  XNOR U9037 ( .A(n6644), .B(\w3[6][40] ), .Z(n6529) );
  XNOR U9038 ( .A(n6530), .B(n6529), .Z(\w1[7][32] ) );
  XOR U9039 ( .A(\w3[6][34] ), .B(\w3[6][58] ), .Z(n6591) );
  XOR U9040 ( .A(n6591), .B(key[929]), .Z(n6532) );
  XOR U9041 ( .A(\w3[6][41] ), .B(\w3[6][49] ), .Z(n6615) );
  XNOR U9042 ( .A(\w3[6][57] ), .B(n6615), .Z(n6531) );
  XNOR U9043 ( .A(n6532), .B(n6531), .Z(\w1[7][33] ) );
  XOR U9044 ( .A(\w3[6][35] ), .B(\w3[6][59] ), .Z(n6562) );
  XOR U9045 ( .A(n6562), .B(key[930]), .Z(n6534) );
  XOR U9046 ( .A(\w3[6][42] ), .B(\w3[6][50] ), .Z(n6619) );
  XNOR U9047 ( .A(\w3[6][58] ), .B(n6619), .Z(n6533) );
  XNOR U9048 ( .A(n6534), .B(n6533), .Z(\w1[7][34] ) );
  XOR U9049 ( .A(\w3[6][36] ), .B(\w3[6][32] ), .Z(n6564) );
  XOR U9050 ( .A(n6564), .B(key[931]), .Z(n6537) );
  XOR U9051 ( .A(\w3[6][43] ), .B(\w3[6][51] ), .Z(n6590) );
  XNOR U9052 ( .A(\w3[6][56] ), .B(n6590), .Z(n6535) );
  XNOR U9053 ( .A(\w3[6][60] ), .B(n6535), .Z(n6624) );
  XNOR U9054 ( .A(\w3[6][59] ), .B(n6624), .Z(n6536) );
  XNOR U9055 ( .A(n6537), .B(n6536), .Z(\w1[7][35] ) );
  XOR U9056 ( .A(\w3[6][32] ), .B(\w3[6][37] ), .Z(n6569) );
  XOR U9057 ( .A(n6569), .B(key[932]), .Z(n6541) );
  XOR U9058 ( .A(\w3[6][52] ), .B(\w3[6][61] ), .Z(n6539) );
  XNOR U9059 ( .A(\w3[6][56] ), .B(\w3[6][44] ), .Z(n6538) );
  XNOR U9060 ( .A(n6539), .B(n6538), .Z(n6632) );
  XNOR U9061 ( .A(\w3[6][60] ), .B(n6632), .Z(n6540) );
  XNOR U9062 ( .A(n6541), .B(n6540), .Z(\w1[7][36] ) );
  XOR U9063 ( .A(\w3[6][38] ), .B(\w3[6][62] ), .Z(n6575) );
  XOR U9064 ( .A(n6575), .B(key[933]), .Z(n6543) );
  XOR U9065 ( .A(\w3[6][45] ), .B(\w3[6][53] ), .Z(n6635) );
  XNOR U9066 ( .A(\w3[6][61] ), .B(n6635), .Z(n6542) );
  XNOR U9067 ( .A(n6543), .B(n6542), .Z(\w1[7][37] ) );
  XOR U9068 ( .A(\w3[6][32] ), .B(\w3[6][39] ), .Z(n6576) );
  XOR U9069 ( .A(n6576), .B(key[934]), .Z(n6545) );
  XOR U9070 ( .A(\w3[6][46] ), .B(\w3[6][54] ), .Z(n6601) );
  XNOR U9071 ( .A(\w3[6][56] ), .B(\w3[6][63] ), .Z(n6547) );
  XNOR U9072 ( .A(n6601), .B(n6547), .Z(n6640) );
  XNOR U9073 ( .A(\w3[6][62] ), .B(n6640), .Z(n6544) );
  XNOR U9074 ( .A(n6545), .B(n6544), .Z(\w1[7][38] ) );
  XOR U9075 ( .A(\w3[6][47] ), .B(\w3[6][55] ), .Z(n6643) );
  XNOR U9076 ( .A(n6643), .B(key[935]), .Z(n6546) );
  XNOR U9077 ( .A(n6547), .B(n6546), .Z(n6548) );
  XNOR U9078 ( .A(\w3[6][32] ), .B(n6548), .Z(\w1[7][39] ) );
  XOR U9079 ( .A(n6549), .B(key[899]), .Z(n6552) );
  XNOR U9080 ( .A(n6550), .B(\w3[6][27] ), .Z(n6551) );
  XNOR U9081 ( .A(n6552), .B(n6551), .Z(\w1[7][3] ) );
  XOR U9082 ( .A(\w3[6][32] ), .B(key[936]), .Z(n6554) );
  XNOR U9083 ( .A(\w3[6][33] ), .B(\w3[6][41] ), .Z(n6553) );
  XNOR U9084 ( .A(n6554), .B(n6553), .Z(n6555) );
  XOR U9085 ( .A(n6644), .B(n6555), .Z(\w1[7][40] ) );
  XOR U9086 ( .A(\w3[6][42] ), .B(key[937]), .Z(n6557) );
  XNOR U9087 ( .A(\w3[6][49] ), .B(\w3[6][34] ), .Z(n6556) );
  XNOR U9088 ( .A(n6557), .B(n6556), .Z(n6558) );
  XOR U9089 ( .A(n6583), .B(n6558), .Z(\w1[7][41] ) );
  XOR U9090 ( .A(\w3[6][43] ), .B(key[938]), .Z(n6560) );
  XNOR U9091 ( .A(\w3[6][50] ), .B(\w3[6][35] ), .Z(n6559) );
  XNOR U9092 ( .A(n6560), .B(n6559), .Z(n6561) );
  XOR U9093 ( .A(n6591), .B(n6561), .Z(\w1[7][42] ) );
  XNOR U9094 ( .A(\w3[6][40] ), .B(n6562), .Z(n6563) );
  XNOR U9095 ( .A(\w3[6][44] ), .B(n6563), .Z(n6594) );
  XOR U9096 ( .A(n6594), .B(key[939]), .Z(n6566) );
  XNOR U9097 ( .A(\w3[6][51] ), .B(n6564), .Z(n6565) );
  XNOR U9098 ( .A(n6566), .B(n6565), .Z(\w1[7][43] ) );
  XOR U9099 ( .A(\w3[6][36] ), .B(\w3[6][45] ), .Z(n6568) );
  XNOR U9100 ( .A(\w3[6][40] ), .B(\w3[6][60] ), .Z(n6567) );
  XNOR U9101 ( .A(n6568), .B(n6567), .Z(n6597) );
  XOR U9102 ( .A(n6597), .B(key[940]), .Z(n6571) );
  XNOR U9103 ( .A(\w3[6][52] ), .B(n6569), .Z(n6570) );
  XNOR U9104 ( .A(n6571), .B(n6570), .Z(\w1[7][44] ) );
  XOR U9105 ( .A(\w3[6][61] ), .B(\w3[6][37] ), .Z(n6600) );
  XOR U9106 ( .A(n6600), .B(key[941]), .Z(n6573) );
  XNOR U9107 ( .A(\w3[6][38] ), .B(\w3[6][46] ), .Z(n6572) );
  XNOR U9108 ( .A(n6573), .B(n6572), .Z(n6574) );
  XOR U9109 ( .A(\w3[6][53] ), .B(n6574), .Z(\w1[7][45] ) );
  XNOR U9110 ( .A(\w3[6][40] ), .B(\w3[6][47] ), .Z(n6609) );
  XNOR U9111 ( .A(n6575), .B(n6609), .Z(n6604) );
  XOR U9112 ( .A(n6604), .B(key[942]), .Z(n6578) );
  XNOR U9113 ( .A(\w3[6][54] ), .B(n6576), .Z(n6577) );
  XNOR U9114 ( .A(n6578), .B(n6577), .Z(\w1[7][46] ) );
  XOR U9115 ( .A(\w3[6][63] ), .B(\w3[6][39] ), .Z(n6607) );
  XOR U9116 ( .A(n6607), .B(key[943]), .Z(n6580) );
  XOR U9117 ( .A(\w3[6][40] ), .B(\w3[6][32] ), .Z(n6611) );
  XNOR U9118 ( .A(\w3[6][55] ), .B(n6611), .Z(n6579) );
  XNOR U9119 ( .A(n6580), .B(n6579), .Z(\w1[7][47] ) );
  XOR U9120 ( .A(n6611), .B(key[944]), .Z(n6582) );
  XNOR U9121 ( .A(\w3[6][56] ), .B(n6615), .Z(n6581) );
  XNOR U9122 ( .A(n6582), .B(n6581), .Z(\w1[7][48] ) );
  XOR U9123 ( .A(n6619), .B(key[945]), .Z(n6585) );
  XNOR U9124 ( .A(n6583), .B(\w3[6][41] ), .Z(n6584) );
  XNOR U9125 ( .A(n6585), .B(n6584), .Z(\w1[7][49] ) );
  XOR U9126 ( .A(n6586), .B(key[900]), .Z(n6589) );
  XNOR U9127 ( .A(n6587), .B(\w3[6][28] ), .Z(n6588) );
  XNOR U9128 ( .A(n6589), .B(n6588), .Z(\w1[7][4] ) );
  XOR U9129 ( .A(n6590), .B(key[946]), .Z(n6593) );
  XNOR U9130 ( .A(n6591), .B(\w3[6][42] ), .Z(n6592) );
  XNOR U9131 ( .A(n6593), .B(n6592), .Z(\w1[7][50] ) );
  XOR U9132 ( .A(\w3[6][48] ), .B(\w3[6][52] ), .Z(n6623) );
  XOR U9133 ( .A(n6623), .B(key[947]), .Z(n6596) );
  XNOR U9134 ( .A(\w3[6][43] ), .B(n6594), .Z(n6595) );
  XNOR U9135 ( .A(n6596), .B(n6595), .Z(\w1[7][51] ) );
  XOR U9136 ( .A(\w3[6][48] ), .B(\w3[6][53] ), .Z(n6631) );
  XOR U9137 ( .A(n6631), .B(key[948]), .Z(n6599) );
  XNOR U9138 ( .A(\w3[6][44] ), .B(n6597), .Z(n6598) );
  XNOR U9139 ( .A(n6599), .B(n6598), .Z(\w1[7][52] ) );
  XOR U9140 ( .A(n6600), .B(key[949]), .Z(n6603) );
  XNOR U9141 ( .A(\w3[6][45] ), .B(n6601), .Z(n6602) );
  XNOR U9142 ( .A(n6603), .B(n6602), .Z(\w1[7][53] ) );
  XOR U9143 ( .A(\w3[6][48] ), .B(\w3[6][55] ), .Z(n6639) );
  XOR U9144 ( .A(n6639), .B(key[950]), .Z(n6606) );
  XNOR U9145 ( .A(\w3[6][46] ), .B(n6604), .Z(n6605) );
  XNOR U9146 ( .A(n6606), .B(n6605), .Z(\w1[7][54] ) );
  XNOR U9147 ( .A(n6607), .B(key[951]), .Z(n6608) );
  XNOR U9148 ( .A(n6609), .B(n6608), .Z(n6610) );
  XNOR U9149 ( .A(\w3[6][48] ), .B(n6610), .Z(\w1[7][55] ) );
  XOR U9150 ( .A(n6611), .B(key[952]), .Z(n6613) );
  XNOR U9151 ( .A(\w3[6][48] ), .B(\w3[6][49] ), .Z(n6612) );
  XNOR U9152 ( .A(n6613), .B(n6612), .Z(n6614) );
  XOR U9153 ( .A(\w3[6][57] ), .B(n6614), .Z(\w1[7][56] ) );
  XOR U9154 ( .A(\w3[6][50] ), .B(key[953]), .Z(n6617) );
  XNOR U9155 ( .A(n6615), .B(\w3[6][58] ), .Z(n6616) );
  XNOR U9156 ( .A(n6617), .B(n6616), .Z(n6618) );
  XOR U9157 ( .A(\w3[6][33] ), .B(n6618), .Z(\w1[7][57] ) );
  XOR U9158 ( .A(\w3[6][51] ), .B(key[954]), .Z(n6621) );
  XNOR U9159 ( .A(n6619), .B(\w3[6][59] ), .Z(n6620) );
  XNOR U9160 ( .A(n6621), .B(n6620), .Z(n6622) );
  XOR U9161 ( .A(\w3[6][34] ), .B(n6622), .Z(\w1[7][58] ) );
  XOR U9162 ( .A(n6623), .B(key[955]), .Z(n6626) );
  XNOR U9163 ( .A(\w3[6][35] ), .B(n6624), .Z(n6625) );
  XNOR U9164 ( .A(n6626), .B(n6625), .Z(\w1[7][59] ) );
  XOR U9165 ( .A(n6627), .B(key[901]), .Z(n6630) );
  XNOR U9166 ( .A(\w3[6][29] ), .B(n6628), .Z(n6629) );
  XNOR U9167 ( .A(n6630), .B(n6629), .Z(\w1[7][5] ) );
  XOR U9168 ( .A(n6631), .B(key[956]), .Z(n6634) );
  XNOR U9169 ( .A(\w3[6][36] ), .B(n6632), .Z(n6633) );
  XNOR U9170 ( .A(n6634), .B(n6633), .Z(\w1[7][60] ) );
  XOR U9171 ( .A(\w3[6][54] ), .B(key[957]), .Z(n6637) );
  XNOR U9172 ( .A(n6635), .B(\w3[6][62] ), .Z(n6636) );
  XNOR U9173 ( .A(n6637), .B(n6636), .Z(n6638) );
  XOR U9174 ( .A(\w3[6][37] ), .B(n6638), .Z(\w1[7][61] ) );
  XOR U9175 ( .A(n6639), .B(key[958]), .Z(n6642) );
  XNOR U9176 ( .A(\w3[6][38] ), .B(n6640), .Z(n6641) );
  XNOR U9177 ( .A(n6642), .B(n6641), .Z(\w1[7][62] ) );
  XOR U9178 ( .A(n6643), .B(key[959]), .Z(n6646) );
  XNOR U9179 ( .A(n6644), .B(\w3[6][39] ), .Z(n6645) );
  XNOR U9180 ( .A(n6646), .B(n6645), .Z(\w1[7][63] ) );
  XOR U9181 ( .A(\w3[6][65] ), .B(\w3[6][89] ), .Z(n6705) );
  XOR U9182 ( .A(n6705), .B(key[960]), .Z(n6648) );
  XOR U9183 ( .A(\w3[6][80] ), .B(\w3[6][88] ), .Z(n6762) );
  XNOR U9184 ( .A(n6762), .B(\w3[6][72] ), .Z(n6647) );
  XNOR U9185 ( .A(n6648), .B(n6647), .Z(\w1[7][64] ) );
  XOR U9186 ( .A(\w3[6][66] ), .B(\w3[6][90] ), .Z(n6709) );
  XOR U9187 ( .A(n6709), .B(key[961]), .Z(n6650) );
  XOR U9188 ( .A(\w3[6][73] ), .B(\w3[6][81] ), .Z(n6733) );
  XNOR U9189 ( .A(\w3[6][89] ), .B(n6733), .Z(n6649) );
  XNOR U9190 ( .A(n6650), .B(n6649), .Z(\w1[7][65] ) );
  XOR U9191 ( .A(\w3[6][67] ), .B(\w3[6][91] ), .Z(n6680) );
  XOR U9192 ( .A(n6680), .B(key[962]), .Z(n6652) );
  XOR U9193 ( .A(\w3[6][74] ), .B(\w3[6][82] ), .Z(n6741) );
  XNOR U9194 ( .A(\w3[6][90] ), .B(n6741), .Z(n6651) );
  XNOR U9195 ( .A(n6652), .B(n6651), .Z(\w1[7][66] ) );
  XOR U9196 ( .A(\w3[6][68] ), .B(\w3[6][64] ), .Z(n6682) );
  XOR U9197 ( .A(n6682), .B(key[963]), .Z(n6655) );
  XOR U9198 ( .A(\w3[6][75] ), .B(\w3[6][83] ), .Z(n6708) );
  XNOR U9199 ( .A(\w3[6][88] ), .B(n6708), .Z(n6653) );
  XNOR U9200 ( .A(\w3[6][92] ), .B(n6653), .Z(n6746) );
  XNOR U9201 ( .A(\w3[6][91] ), .B(n6746), .Z(n6654) );
  XNOR U9202 ( .A(n6655), .B(n6654), .Z(\w1[7][67] ) );
  XOR U9203 ( .A(\w3[6][64] ), .B(\w3[6][69] ), .Z(n6687) );
  XOR U9204 ( .A(n6687), .B(key[964]), .Z(n6659) );
  XOR U9205 ( .A(\w3[6][84] ), .B(\w3[6][93] ), .Z(n6657) );
  XNOR U9206 ( .A(\w3[6][88] ), .B(\w3[6][76] ), .Z(n6656) );
  XNOR U9207 ( .A(n6657), .B(n6656), .Z(n6750) );
  XNOR U9208 ( .A(\w3[6][92] ), .B(n6750), .Z(n6658) );
  XNOR U9209 ( .A(n6659), .B(n6658), .Z(\w1[7][68] ) );
  XOR U9210 ( .A(\w3[6][70] ), .B(\w3[6][94] ), .Z(n6693) );
  XOR U9211 ( .A(n6693), .B(key[965]), .Z(n6661) );
  XOR U9212 ( .A(\w3[6][77] ), .B(\w3[6][85] ), .Z(n6753) );
  XNOR U9213 ( .A(\w3[6][93] ), .B(n6753), .Z(n6660) );
  XNOR U9214 ( .A(n6661), .B(n6660), .Z(\w1[7][69] ) );
  XOR U9215 ( .A(n6662), .B(key[902]), .Z(n6665) );
  XNOR U9216 ( .A(n6663), .B(\w3[6][30] ), .Z(n6664) );
  XNOR U9217 ( .A(n6665), .B(n6664), .Z(\w1[7][6] ) );
  XOR U9218 ( .A(\w3[6][64] ), .B(\w3[6][71] ), .Z(n6694) );
  XOR U9219 ( .A(n6694), .B(key[966]), .Z(n6667) );
  XOR U9220 ( .A(\w3[6][78] ), .B(\w3[6][86] ), .Z(n6719) );
  XNOR U9221 ( .A(\w3[6][88] ), .B(\w3[6][95] ), .Z(n6669) );
  XNOR U9222 ( .A(n6719), .B(n6669), .Z(n6758) );
  XNOR U9223 ( .A(\w3[6][94] ), .B(n6758), .Z(n6666) );
  XNOR U9224 ( .A(n6667), .B(n6666), .Z(\w1[7][70] ) );
  XOR U9225 ( .A(\w3[6][79] ), .B(\w3[6][87] ), .Z(n6761) );
  XNOR U9226 ( .A(n6761), .B(key[967]), .Z(n6668) );
  XNOR U9227 ( .A(n6669), .B(n6668), .Z(n6670) );
  XNOR U9228 ( .A(\w3[6][64] ), .B(n6670), .Z(\w1[7][71] ) );
  XOR U9229 ( .A(\w3[6][64] ), .B(key[968]), .Z(n6672) );
  XNOR U9230 ( .A(\w3[6][65] ), .B(\w3[6][73] ), .Z(n6671) );
  XNOR U9231 ( .A(n6672), .B(n6671), .Z(n6673) );
  XOR U9232 ( .A(n6762), .B(n6673), .Z(\w1[7][72] ) );
  XOR U9233 ( .A(\w3[6][74] ), .B(key[969]), .Z(n6675) );
  XNOR U9234 ( .A(\w3[6][81] ), .B(\w3[6][66] ), .Z(n6674) );
  XNOR U9235 ( .A(n6675), .B(n6674), .Z(n6676) );
  XOR U9236 ( .A(n6705), .B(n6676), .Z(\w1[7][73] ) );
  XOR U9237 ( .A(\w3[6][75] ), .B(key[970]), .Z(n6678) );
  XNOR U9238 ( .A(\w3[6][82] ), .B(\w3[6][67] ), .Z(n6677) );
  XNOR U9239 ( .A(n6678), .B(n6677), .Z(n6679) );
  XOR U9240 ( .A(n6709), .B(n6679), .Z(\w1[7][74] ) );
  XNOR U9241 ( .A(\w3[6][72] ), .B(n6680), .Z(n6681) );
  XNOR U9242 ( .A(\w3[6][76] ), .B(n6681), .Z(n6712) );
  XOR U9243 ( .A(n6712), .B(key[971]), .Z(n6684) );
  XNOR U9244 ( .A(\w3[6][83] ), .B(n6682), .Z(n6683) );
  XNOR U9245 ( .A(n6684), .B(n6683), .Z(\w1[7][75] ) );
  XOR U9246 ( .A(\w3[6][68] ), .B(\w3[6][77] ), .Z(n6686) );
  XNOR U9247 ( .A(\w3[6][72] ), .B(\w3[6][92] ), .Z(n6685) );
  XNOR U9248 ( .A(n6686), .B(n6685), .Z(n6715) );
  XOR U9249 ( .A(n6715), .B(key[972]), .Z(n6689) );
  XNOR U9250 ( .A(\w3[6][84] ), .B(n6687), .Z(n6688) );
  XNOR U9251 ( .A(n6689), .B(n6688), .Z(\w1[7][76] ) );
  XOR U9252 ( .A(\w3[6][93] ), .B(\w3[6][69] ), .Z(n6718) );
  XOR U9253 ( .A(n6718), .B(key[973]), .Z(n6691) );
  XNOR U9254 ( .A(\w3[6][70] ), .B(\w3[6][78] ), .Z(n6690) );
  XNOR U9255 ( .A(n6691), .B(n6690), .Z(n6692) );
  XOR U9256 ( .A(\w3[6][85] ), .B(n6692), .Z(\w1[7][77] ) );
  XNOR U9257 ( .A(\w3[6][72] ), .B(\w3[6][79] ), .Z(n6727) );
  XNOR U9258 ( .A(n6693), .B(n6727), .Z(n6722) );
  XOR U9259 ( .A(n6722), .B(key[974]), .Z(n6696) );
  XNOR U9260 ( .A(\w3[6][86] ), .B(n6694), .Z(n6695) );
  XNOR U9261 ( .A(n6696), .B(n6695), .Z(\w1[7][78] ) );
  XOR U9262 ( .A(\w3[6][95] ), .B(\w3[6][71] ), .Z(n6725) );
  XOR U9263 ( .A(n6725), .B(key[975]), .Z(n6698) );
  XOR U9264 ( .A(\w3[6][72] ), .B(\w3[6][64] ), .Z(n6729) );
  XNOR U9265 ( .A(\w3[6][87] ), .B(n6729), .Z(n6697) );
  XNOR U9266 ( .A(n6698), .B(n6697), .Z(\w1[7][79] ) );
  XNOR U9267 ( .A(n6699), .B(key[903]), .Z(n6700) );
  XNOR U9268 ( .A(n6701), .B(n6700), .Z(n6702) );
  XNOR U9269 ( .A(\w3[6][0] ), .B(n6702), .Z(\w1[7][7] ) );
  XOR U9270 ( .A(n6729), .B(key[976]), .Z(n6704) );
  XNOR U9271 ( .A(\w3[6][88] ), .B(n6733), .Z(n6703) );
  XNOR U9272 ( .A(n6704), .B(n6703), .Z(\w1[7][80] ) );
  XOR U9273 ( .A(n6741), .B(key[977]), .Z(n6707) );
  XNOR U9274 ( .A(n6705), .B(\w3[6][73] ), .Z(n6706) );
  XNOR U9275 ( .A(n6707), .B(n6706), .Z(\w1[7][81] ) );
  XOR U9276 ( .A(n6708), .B(key[978]), .Z(n6711) );
  XNOR U9277 ( .A(n6709), .B(\w3[6][74] ), .Z(n6710) );
  XNOR U9278 ( .A(n6711), .B(n6710), .Z(\w1[7][82] ) );
  XOR U9279 ( .A(\w3[6][80] ), .B(\w3[6][84] ), .Z(n6745) );
  XOR U9280 ( .A(n6745), .B(key[979]), .Z(n6714) );
  XNOR U9281 ( .A(\w3[6][75] ), .B(n6712), .Z(n6713) );
  XNOR U9282 ( .A(n6714), .B(n6713), .Z(\w1[7][83] ) );
  XOR U9283 ( .A(\w3[6][80] ), .B(\w3[6][85] ), .Z(n6749) );
  XOR U9284 ( .A(n6749), .B(key[980]), .Z(n6717) );
  XNOR U9285 ( .A(\w3[6][76] ), .B(n6715), .Z(n6716) );
  XNOR U9286 ( .A(n6717), .B(n6716), .Z(\w1[7][84] ) );
  XOR U9287 ( .A(n6718), .B(key[981]), .Z(n6721) );
  XNOR U9288 ( .A(\w3[6][77] ), .B(n6719), .Z(n6720) );
  XNOR U9289 ( .A(n6721), .B(n6720), .Z(\w1[7][85] ) );
  XOR U9290 ( .A(\w3[6][80] ), .B(\w3[6][87] ), .Z(n6757) );
  XOR U9291 ( .A(n6757), .B(key[982]), .Z(n6724) );
  XNOR U9292 ( .A(\w3[6][78] ), .B(n6722), .Z(n6723) );
  XNOR U9293 ( .A(n6724), .B(n6723), .Z(\w1[7][86] ) );
  XNOR U9294 ( .A(n6725), .B(key[983]), .Z(n6726) );
  XNOR U9295 ( .A(n6727), .B(n6726), .Z(n6728) );
  XNOR U9296 ( .A(\w3[6][80] ), .B(n6728), .Z(\w1[7][87] ) );
  XOR U9297 ( .A(n6729), .B(key[984]), .Z(n6731) );
  XNOR U9298 ( .A(\w3[6][80] ), .B(\w3[6][81] ), .Z(n6730) );
  XNOR U9299 ( .A(n6731), .B(n6730), .Z(n6732) );
  XOR U9300 ( .A(\w3[6][89] ), .B(n6732), .Z(\w1[7][88] ) );
  XOR U9301 ( .A(\w3[6][82] ), .B(key[985]), .Z(n6735) );
  XNOR U9302 ( .A(n6733), .B(\w3[6][90] ), .Z(n6734) );
  XNOR U9303 ( .A(n6735), .B(n6734), .Z(n6736) );
  XOR U9304 ( .A(\w3[6][65] ), .B(n6736), .Z(\w1[7][89] ) );
  XOR U9305 ( .A(\w3[6][9] ), .B(key[904]), .Z(n6738) );
  XNOR U9306 ( .A(\w3[6][1] ), .B(\w3[6][0] ), .Z(n6737) );
  XNOR U9307 ( .A(n6738), .B(n6737), .Z(n6739) );
  XOR U9308 ( .A(n6740), .B(n6739), .Z(\w1[7][8] ) );
  XOR U9309 ( .A(\w3[6][83] ), .B(key[986]), .Z(n6743) );
  XNOR U9310 ( .A(n6741), .B(\w3[6][91] ), .Z(n6742) );
  XNOR U9311 ( .A(n6743), .B(n6742), .Z(n6744) );
  XOR U9312 ( .A(\w3[6][66] ), .B(n6744), .Z(\w1[7][90] ) );
  XOR U9313 ( .A(n6745), .B(key[987]), .Z(n6748) );
  XNOR U9314 ( .A(\w3[6][67] ), .B(n6746), .Z(n6747) );
  XNOR U9315 ( .A(n6748), .B(n6747), .Z(\w1[7][91] ) );
  XOR U9316 ( .A(n6749), .B(key[988]), .Z(n6752) );
  XNOR U9317 ( .A(\w3[6][68] ), .B(n6750), .Z(n6751) );
  XNOR U9318 ( .A(n6752), .B(n6751), .Z(\w1[7][92] ) );
  XOR U9319 ( .A(\w3[6][86] ), .B(key[989]), .Z(n6755) );
  XNOR U9320 ( .A(n6753), .B(\w3[6][94] ), .Z(n6754) );
  XNOR U9321 ( .A(n6755), .B(n6754), .Z(n6756) );
  XOR U9322 ( .A(\w3[6][69] ), .B(n6756), .Z(\w1[7][93] ) );
  XOR U9323 ( .A(n6757), .B(key[990]), .Z(n6760) );
  XNOR U9324 ( .A(\w3[6][70] ), .B(n6758), .Z(n6759) );
  XNOR U9325 ( .A(n6760), .B(n6759), .Z(\w1[7][94] ) );
  XOR U9326 ( .A(n6761), .B(key[991]), .Z(n6764) );
  XNOR U9327 ( .A(n6762), .B(\w3[6][71] ), .Z(n6763) );
  XNOR U9328 ( .A(n6764), .B(n6763), .Z(\w1[7][95] ) );
  XOR U9329 ( .A(\w3[6][104] ), .B(key[992]), .Z(n6768) );
  XNOR U9330 ( .A(n6766), .B(n6765), .Z(n6767) );
  XNOR U9331 ( .A(n6768), .B(n6767), .Z(\w1[7][96] ) );
  XOR U9332 ( .A(n6769), .B(key[993]), .Z(n6772) );
  XNOR U9333 ( .A(\w3[6][121] ), .B(n6770), .Z(n6771) );
  XNOR U9334 ( .A(n6772), .B(n6771), .Z(\w1[7][97] ) );
  XOR U9335 ( .A(n6773), .B(key[994]), .Z(n6776) );
  XNOR U9336 ( .A(\w3[6][122] ), .B(n6774), .Z(n6775) );
  XNOR U9337 ( .A(n6776), .B(n6775), .Z(\w1[7][98] ) );
  XOR U9338 ( .A(n6777), .B(key[995]), .Z(n6780) );
  XNOR U9339 ( .A(n6778), .B(\w3[6][123] ), .Z(n6779) );
  XNOR U9340 ( .A(n6780), .B(n6779), .Z(\w1[7][99] ) );
  XOR U9341 ( .A(\w3[6][10] ), .B(key[905]), .Z(n6782) );
  XNOR U9342 ( .A(\w3[6][2] ), .B(\w3[6][17] ), .Z(n6781) );
  XNOR U9343 ( .A(n6782), .B(n6781), .Z(n6783) );
  XOR U9344 ( .A(n6784), .B(n6783), .Z(\w1[7][9] ) );
  XOR U9345 ( .A(\w3[7][8] ), .B(key[1024]), .Z(n6786) );
  XOR U9346 ( .A(\w3[7][1] ), .B(\w3[7][25] ), .Z(n7208) );
  XOR U9347 ( .A(\w3[7][16] ), .B(\w3[7][24] ), .Z(n7164) );
  XNOR U9348 ( .A(n7208), .B(n7164), .Z(n6785) );
  XNOR U9349 ( .A(n6786), .B(n6785), .Z(\w1[8][0] ) );
  XOR U9350 ( .A(\w3[7][96] ), .B(\w3[7][101] ), .Z(n6812) );
  XOR U9351 ( .A(n6812), .B(key[1124]), .Z(n6790) );
  XOR U9352 ( .A(\w3[7][116] ), .B(\w3[7][125] ), .Z(n6788) );
  XNOR U9353 ( .A(\w3[7][120] ), .B(\w3[7][108] ), .Z(n6787) );
  XNOR U9354 ( .A(n6788), .B(n6787), .Z(n6869) );
  XNOR U9355 ( .A(\w3[7][124] ), .B(n6869), .Z(n6789) );
  XNOR U9356 ( .A(n6790), .B(n6789), .Z(\w1[8][100] ) );
  XOR U9357 ( .A(\w3[7][102] ), .B(\w3[7][126] ), .Z(n6821) );
  XOR U9358 ( .A(n6821), .B(key[1125]), .Z(n6792) );
  XOR U9359 ( .A(\w3[7][109] ), .B(\w3[7][117] ), .Z(n6872) );
  XNOR U9360 ( .A(\w3[7][125] ), .B(n6872), .Z(n6791) );
  XNOR U9361 ( .A(n6792), .B(n6791), .Z(\w1[8][101] ) );
  XOR U9362 ( .A(\w3[7][96] ), .B(\w3[7][103] ), .Z(n6822) );
  XOR U9363 ( .A(n6822), .B(key[1126]), .Z(n6794) );
  XOR U9364 ( .A(\w3[7][110] ), .B(\w3[7][118] ), .Z(n6840) );
  XNOR U9365 ( .A(\w3[7][120] ), .B(\w3[7][127] ), .Z(n6796) );
  XNOR U9366 ( .A(n6840), .B(n6796), .Z(n6877) );
  XNOR U9367 ( .A(\w3[7][126] ), .B(n6877), .Z(n6793) );
  XNOR U9368 ( .A(n6794), .B(n6793), .Z(\w1[8][102] ) );
  XOR U9369 ( .A(\w3[7][111] ), .B(\w3[7][119] ), .Z(n6880) );
  XNOR U9370 ( .A(n6880), .B(key[1127]), .Z(n6795) );
  XNOR U9371 ( .A(n6796), .B(n6795), .Z(n6797) );
  XNOR U9372 ( .A(\w3[7][96] ), .B(n6797), .Z(\w1[8][103] ) );
  XOR U9373 ( .A(key[1128]), .B(\w3[7][105] ), .Z(n6799) );
  XNOR U9374 ( .A(\w3[7][96] ), .B(\w3[7][97] ), .Z(n6798) );
  XNOR U9375 ( .A(n6799), .B(n6798), .Z(n6800) );
  XNOR U9376 ( .A(\w3[7][120] ), .B(\w3[7][112] ), .Z(n7190) );
  XNOR U9377 ( .A(n6800), .B(n7190), .Z(\w1[8][104] ) );
  XOR U9378 ( .A(\w3[7][106] ), .B(\w3[7][98] ), .Z(n6802) );
  XOR U9379 ( .A(\w3[7][121] ), .B(\w3[7][113] ), .Z(n6854) );
  XNOR U9380 ( .A(n6854), .B(key[1129]), .Z(n6801) );
  XNOR U9381 ( .A(n6802), .B(n6801), .Z(n6803) );
  XOR U9382 ( .A(\w3[7][97] ), .B(n6803), .Z(\w1[8][105] ) );
  XOR U9383 ( .A(\w3[7][107] ), .B(\w3[7][99] ), .Z(n6805) );
  XOR U9384 ( .A(\w3[7][98] ), .B(\w3[7][122] ), .Z(n7194) );
  XNOR U9385 ( .A(n7194), .B(key[1130]), .Z(n6804) );
  XNOR U9386 ( .A(n6805), .B(n6804), .Z(n6806) );
  XOR U9387 ( .A(\w3[7][114] ), .B(n6806), .Z(\w1[8][106] ) );
  XOR U9388 ( .A(\w3[7][99] ), .B(\w3[7][123] ), .Z(n7198) );
  XNOR U9389 ( .A(\w3[7][108] ), .B(n7198), .Z(n6807) );
  XNOR U9390 ( .A(\w3[7][104] ), .B(n6807), .Z(n6833) );
  XOR U9391 ( .A(n6833), .B(key[1131]), .Z(n6809) );
  XOR U9392 ( .A(\w3[7][96] ), .B(\w3[7][100] ), .Z(n7202) );
  XNOR U9393 ( .A(\w3[7][115] ), .B(n7202), .Z(n6808) );
  XNOR U9394 ( .A(n6809), .B(n6808), .Z(\w1[8][107] ) );
  XOR U9395 ( .A(\w3[7][100] ), .B(\w3[7][104] ), .Z(n6811) );
  XNOR U9396 ( .A(\w3[7][124] ), .B(\w3[7][109] ), .Z(n6810) );
  XNOR U9397 ( .A(n6811), .B(n6810), .Z(n6836) );
  XOR U9398 ( .A(n6836), .B(key[1132]), .Z(n6814) );
  XNOR U9399 ( .A(\w3[7][116] ), .B(n6812), .Z(n6813) );
  XNOR U9400 ( .A(n6814), .B(n6813), .Z(\w1[8][108] ) );
  XOR U9401 ( .A(\w3[7][125] ), .B(\w3[7][101] ), .Z(n6839) );
  XOR U9402 ( .A(n6839), .B(key[1133]), .Z(n6816) );
  XNOR U9403 ( .A(\w3[7][102] ), .B(\w3[7][110] ), .Z(n6815) );
  XNOR U9404 ( .A(n6816), .B(n6815), .Z(n6817) );
  XOR U9405 ( .A(\w3[7][117] ), .B(n6817), .Z(\w1[8][109] ) );
  XOR U9406 ( .A(\w3[7][11] ), .B(\w3[7][18] ), .Z(n6819) );
  XOR U9407 ( .A(\w3[7][2] ), .B(\w3[7][26] ), .Z(n6903) );
  XNOR U9408 ( .A(n6903), .B(key[1034]), .Z(n6818) );
  XNOR U9409 ( .A(n6819), .B(n6818), .Z(n6820) );
  XOR U9410 ( .A(\w3[7][3] ), .B(n6820), .Z(\w1[8][10] ) );
  XNOR U9411 ( .A(\w3[7][111] ), .B(\w3[7][104] ), .Z(n6848) );
  XNOR U9412 ( .A(n6821), .B(n6848), .Z(n6843) );
  XOR U9413 ( .A(n6843), .B(key[1134]), .Z(n6824) );
  XNOR U9414 ( .A(\w3[7][118] ), .B(n6822), .Z(n6823) );
  XNOR U9415 ( .A(n6824), .B(n6823), .Z(\w1[8][110] ) );
  XOR U9416 ( .A(\w3[7][127] ), .B(\w3[7][103] ), .Z(n6846) );
  XOR U9417 ( .A(n6846), .B(key[1135]), .Z(n6826) );
  XOR U9418 ( .A(\w3[7][96] ), .B(\w3[7][104] ), .Z(n6853) );
  XNOR U9419 ( .A(\w3[7][119] ), .B(n6853), .Z(n6825) );
  XNOR U9420 ( .A(n6826), .B(n6825), .Z(\w1[8][111] ) );
  XOR U9421 ( .A(\w3[7][105] ), .B(\w3[7][113] ), .Z(n7193) );
  XOR U9422 ( .A(n7193), .B(key[1136]), .Z(n6828) );
  XNOR U9423 ( .A(\w3[7][120] ), .B(n6853), .Z(n6827) );
  XNOR U9424 ( .A(n6828), .B(n6827), .Z(\w1[8][112] ) );
  XOR U9425 ( .A(\w3[7][97] ), .B(\w3[7][121] ), .Z(n7189) );
  XOR U9426 ( .A(n7189), .B(key[1137]), .Z(n6830) );
  XOR U9427 ( .A(\w3[7][106] ), .B(\w3[7][114] ), .Z(n7197) );
  XNOR U9428 ( .A(\w3[7][105] ), .B(n7197), .Z(n6829) );
  XNOR U9429 ( .A(n6830), .B(n6829), .Z(\w1[8][113] ) );
  XOR U9430 ( .A(\w3[7][107] ), .B(\w3[7][115] ), .Z(n6864) );
  XOR U9431 ( .A(n6864), .B(key[1138]), .Z(n6832) );
  XNOR U9432 ( .A(\w3[7][106] ), .B(n7194), .Z(n6831) );
  XNOR U9433 ( .A(n6832), .B(n6831), .Z(\w1[8][114] ) );
  XOR U9434 ( .A(\w3[7][116] ), .B(\w3[7][112] ), .Z(n6865) );
  XOR U9435 ( .A(n6865), .B(key[1139]), .Z(n6835) );
  XNOR U9436 ( .A(\w3[7][107] ), .B(n6833), .Z(n6834) );
  XNOR U9437 ( .A(n6835), .B(n6834), .Z(\w1[8][115] ) );
  XOR U9438 ( .A(\w3[7][117] ), .B(\w3[7][112] ), .Z(n6868) );
  XOR U9439 ( .A(n6868), .B(key[1140]), .Z(n6838) );
  XNOR U9440 ( .A(\w3[7][108] ), .B(n6836), .Z(n6837) );
  XNOR U9441 ( .A(n6838), .B(n6837), .Z(\w1[8][116] ) );
  XOR U9442 ( .A(n6839), .B(key[1141]), .Z(n6842) );
  XNOR U9443 ( .A(\w3[7][109] ), .B(n6840), .Z(n6841) );
  XNOR U9444 ( .A(n6842), .B(n6841), .Z(\w1[8][117] ) );
  XOR U9445 ( .A(\w3[7][119] ), .B(\w3[7][112] ), .Z(n6876) );
  XOR U9446 ( .A(n6876), .B(key[1142]), .Z(n6845) );
  XNOR U9447 ( .A(\w3[7][110] ), .B(n6843), .Z(n6844) );
  XNOR U9448 ( .A(n6845), .B(n6844), .Z(\w1[8][118] ) );
  XNOR U9449 ( .A(n6846), .B(key[1143]), .Z(n6847) );
  XNOR U9450 ( .A(n6848), .B(n6847), .Z(n6849) );
  XNOR U9451 ( .A(\w3[7][112] ), .B(n6849), .Z(\w1[8][119] ) );
  XOR U9452 ( .A(\w3[7][3] ), .B(\w3[7][27] ), .Z(n6944) );
  XNOR U9453 ( .A(\w3[7][8] ), .B(\w3[7][12] ), .Z(n6850) );
  XNOR U9454 ( .A(n6944), .B(n6850), .Z(n6900) );
  XOR U9455 ( .A(n6900), .B(key[1035]), .Z(n6852) );
  XOR U9456 ( .A(\w3[7][0] ), .B(\w3[7][4] ), .Z(n6974) );
  XNOR U9457 ( .A(\w3[7][19] ), .B(n6974), .Z(n6851) );
  XNOR U9458 ( .A(n6852), .B(n6851), .Z(\w1[8][11] ) );
  XOR U9459 ( .A(n6853), .B(key[1144]), .Z(n6856) );
  XNOR U9460 ( .A(\w3[7][112] ), .B(n6854), .Z(n6855) );
  XNOR U9461 ( .A(n6856), .B(n6855), .Z(\w1[8][120] ) );
  XOR U9462 ( .A(n7193), .B(key[1145]), .Z(n6858) );
  XNOR U9463 ( .A(\w3[7][114] ), .B(\w3[7][122] ), .Z(n6857) );
  XNOR U9464 ( .A(n6858), .B(n6857), .Z(n6859) );
  XOR U9465 ( .A(\w3[7][97] ), .B(n6859), .Z(\w1[8][121] ) );
  XOR U9466 ( .A(n7197), .B(key[1146]), .Z(n6861) );
  XNOR U9467 ( .A(\w3[7][115] ), .B(\w3[7][123] ), .Z(n6860) );
  XNOR U9468 ( .A(n6861), .B(n6860), .Z(n6862) );
  XOR U9469 ( .A(\w3[7][98] ), .B(n6862), .Z(\w1[8][122] ) );
  XNOR U9470 ( .A(\w3[7][124] ), .B(\w3[7][120] ), .Z(n6863) );
  XNOR U9471 ( .A(n6864), .B(n6863), .Z(n7201) );
  XOR U9472 ( .A(n7201), .B(key[1147]), .Z(n6867) );
  XNOR U9473 ( .A(\w3[7][99] ), .B(n6865), .Z(n6866) );
  XNOR U9474 ( .A(n6867), .B(n6866), .Z(\w1[8][123] ) );
  XOR U9475 ( .A(n6868), .B(key[1148]), .Z(n6871) );
  XNOR U9476 ( .A(n6869), .B(\w3[7][100] ), .Z(n6870) );
  XNOR U9477 ( .A(n6871), .B(n6870), .Z(\w1[8][124] ) );
  XOR U9478 ( .A(\w3[7][118] ), .B(key[1149]), .Z(n6874) );
  XNOR U9479 ( .A(n6872), .B(\w3[7][126] ), .Z(n6873) );
  XNOR U9480 ( .A(n6874), .B(n6873), .Z(n6875) );
  XOR U9481 ( .A(\w3[7][101] ), .B(n6875), .Z(\w1[8][125] ) );
  XOR U9482 ( .A(n6876), .B(key[1150]), .Z(n6879) );
  XNOR U9483 ( .A(\w3[7][102] ), .B(n6877), .Z(n6878) );
  XNOR U9484 ( .A(n6879), .B(n6878), .Z(\w1[8][126] ) );
  XNOR U9485 ( .A(n6880), .B(key[1151]), .Z(n6881) );
  XNOR U9486 ( .A(n7190), .B(n6881), .Z(n6882) );
  XNOR U9487 ( .A(\w3[7][103] ), .B(n6882), .Z(\w1[8][127] ) );
  XOR U9488 ( .A(\w3[7][13] ), .B(\w3[7][28] ), .Z(n6884) );
  XNOR U9489 ( .A(\w3[7][8] ), .B(\w3[7][4] ), .Z(n6883) );
  XNOR U9490 ( .A(n6884), .B(n6883), .Z(n6906) );
  XOR U9491 ( .A(n6906), .B(key[1036]), .Z(n6886) );
  XOR U9492 ( .A(\w3[7][0] ), .B(\w3[7][5] ), .Z(n7011) );
  XNOR U9493 ( .A(\w3[7][20] ), .B(n7011), .Z(n6885) );
  XNOR U9494 ( .A(n6886), .B(n6885), .Z(\w1[8][12] ) );
  XOR U9495 ( .A(\w3[7][14] ), .B(\w3[7][21] ), .Z(n6888) );
  XOR U9496 ( .A(\w3[7][5] ), .B(\w3[7][29] ), .Z(n6909) );
  XNOR U9497 ( .A(n6909), .B(key[1037]), .Z(n6887) );
  XNOR U9498 ( .A(n6888), .B(n6887), .Z(n6889) );
  XOR U9499 ( .A(\w3[7][6] ), .B(n6889), .Z(\w1[8][13] ) );
  XOR U9500 ( .A(\w3[7][6] ), .B(\w3[7][30] ), .Z(n7052) );
  XNOR U9501 ( .A(\w3[7][8] ), .B(\w3[7][15] ), .Z(n6917) );
  XNOR U9502 ( .A(n7052), .B(n6917), .Z(n6912) );
  XOR U9503 ( .A(n6912), .B(key[1038]), .Z(n6891) );
  XOR U9504 ( .A(\w3[7][0] ), .B(\w3[7][7] ), .Z(n7087) );
  XNOR U9505 ( .A(\w3[7][22] ), .B(n7087), .Z(n6890) );
  XNOR U9506 ( .A(n6891), .B(n6890), .Z(\w1[8][14] ) );
  XOR U9507 ( .A(\w3[7][7] ), .B(\w3[7][31] ), .Z(n6915) );
  XOR U9508 ( .A(n6915), .B(key[1039]), .Z(n6893) );
  XOR U9509 ( .A(\w3[7][8] ), .B(\w3[7][0] ), .Z(n6919) );
  XNOR U9510 ( .A(\w3[7][23] ), .B(n6919), .Z(n6892) );
  XNOR U9511 ( .A(n6893), .B(n6892), .Z(\w1[8][15] ) );
  XOR U9512 ( .A(\w3[7][17] ), .B(\w3[7][9] ), .Z(n6923) );
  XOR U9513 ( .A(n6923), .B(key[1040]), .Z(n6895) );
  XNOR U9514 ( .A(\w3[7][24] ), .B(n6919), .Z(n6894) );
  XNOR U9515 ( .A(n6895), .B(n6894), .Z(\w1[8][16] ) );
  XOR U9516 ( .A(\w3[7][18] ), .B(\w3[7][10] ), .Z(n6943) );
  XOR U9517 ( .A(n6943), .B(key[1041]), .Z(n6897) );
  XNOR U9518 ( .A(n7208), .B(\w3[7][9] ), .Z(n6896) );
  XNOR U9519 ( .A(n6897), .B(n6896), .Z(\w1[8][17] ) );
  XOR U9520 ( .A(\w3[7][11] ), .B(\w3[7][19] ), .Z(n6931) );
  XOR U9521 ( .A(n6931), .B(key[1042]), .Z(n6899) );
  XNOR U9522 ( .A(n6903), .B(\w3[7][10] ), .Z(n6898) );
  XNOR U9523 ( .A(n6899), .B(n6898), .Z(\w1[8][18] ) );
  XOR U9524 ( .A(\w3[7][16] ), .B(\w3[7][20] ), .Z(n6932) );
  XOR U9525 ( .A(n6932), .B(key[1043]), .Z(n6902) );
  XNOR U9526 ( .A(\w3[7][11] ), .B(n6900), .Z(n6901) );
  XNOR U9527 ( .A(n6902), .B(n6901), .Z(\w1[8][19] ) );
  XOR U9528 ( .A(n6923), .B(key[1025]), .Z(n6905) );
  XNOR U9529 ( .A(\w3[7][25] ), .B(n6903), .Z(n6904) );
  XNOR U9530 ( .A(n6905), .B(n6904), .Z(\w1[8][1] ) );
  XOR U9531 ( .A(\w3[7][16] ), .B(\w3[7][21] ), .Z(n6937) );
  XOR U9532 ( .A(n6937), .B(key[1044]), .Z(n6908) );
  XNOR U9533 ( .A(\w3[7][12] ), .B(n6906), .Z(n6907) );
  XNOR U9534 ( .A(n6908), .B(n6907), .Z(\w1[8][20] ) );
  XOR U9535 ( .A(\w3[7][14] ), .B(\w3[7][22] ), .Z(n6947) );
  XOR U9536 ( .A(n6947), .B(key[1045]), .Z(n6911) );
  XNOR U9537 ( .A(\w3[7][13] ), .B(n6909), .Z(n6910) );
  XNOR U9538 ( .A(n6911), .B(n6910), .Z(\w1[8][21] ) );
  XOR U9539 ( .A(\w3[7][16] ), .B(\w3[7][23] ), .Z(n6948) );
  XOR U9540 ( .A(n6948), .B(key[1046]), .Z(n6914) );
  XNOR U9541 ( .A(\w3[7][14] ), .B(n6912), .Z(n6913) );
  XNOR U9542 ( .A(n6914), .B(n6913), .Z(\w1[8][22] ) );
  XNOR U9543 ( .A(n6915), .B(key[1047]), .Z(n6916) );
  XNOR U9544 ( .A(n6917), .B(n6916), .Z(n6918) );
  XNOR U9545 ( .A(\w3[7][16] ), .B(n6918), .Z(\w1[8][23] ) );
  XOR U9546 ( .A(\w3[7][17] ), .B(key[1048]), .Z(n6921) );
  XNOR U9547 ( .A(\w3[7][25] ), .B(n6919), .Z(n6920) );
  XNOR U9548 ( .A(n6921), .B(n6920), .Z(n6922) );
  XOR U9549 ( .A(\w3[7][16] ), .B(n6922), .Z(\w1[8][24] ) );
  XOR U9550 ( .A(n6923), .B(key[1049]), .Z(n6925) );
  XNOR U9551 ( .A(\w3[7][1] ), .B(\w3[7][26] ), .Z(n6924) );
  XNOR U9552 ( .A(n6925), .B(n6924), .Z(n6926) );
  XOR U9553 ( .A(\w3[7][18] ), .B(n6926), .Z(\w1[8][25] ) );
  XOR U9554 ( .A(n6943), .B(key[1050]), .Z(n6928) );
  XNOR U9555 ( .A(\w3[7][2] ), .B(\w3[7][19] ), .Z(n6927) );
  XNOR U9556 ( .A(n6928), .B(n6927), .Z(n6929) );
  XOR U9557 ( .A(\w3[7][27] ), .B(n6929), .Z(\w1[8][26] ) );
  XNOR U9558 ( .A(\w3[7][24] ), .B(\w3[7][28] ), .Z(n6930) );
  XNOR U9559 ( .A(n6931), .B(n6930), .Z(n6973) );
  XOR U9560 ( .A(n6973), .B(key[1051]), .Z(n6934) );
  XNOR U9561 ( .A(\w3[7][3] ), .B(n6932), .Z(n6933) );
  XNOR U9562 ( .A(n6934), .B(n6933), .Z(\w1[8][27] ) );
  XOR U9563 ( .A(\w3[7][20] ), .B(\w3[7][29] ), .Z(n6936) );
  XNOR U9564 ( .A(\w3[7][24] ), .B(\w3[7][12] ), .Z(n6935) );
  XNOR U9565 ( .A(n6936), .B(n6935), .Z(n7010) );
  XOR U9566 ( .A(n7010), .B(key[1052]), .Z(n6939) );
  XNOR U9567 ( .A(\w3[7][4] ), .B(n6937), .Z(n6938) );
  XNOR U9568 ( .A(n6939), .B(n6938), .Z(\w1[8][28] ) );
  XOR U9569 ( .A(\w3[7][13] ), .B(\w3[7][21] ), .Z(n7051) );
  XOR U9570 ( .A(n7051), .B(key[1053]), .Z(n6941) );
  XNOR U9571 ( .A(\w3[7][22] ), .B(\w3[7][30] ), .Z(n6940) );
  XNOR U9572 ( .A(n6941), .B(n6940), .Z(n6942) );
  XOR U9573 ( .A(\w3[7][5] ), .B(n6942), .Z(\w1[8][29] ) );
  XOR U9574 ( .A(n6943), .B(key[1026]), .Z(n6946) );
  XNOR U9575 ( .A(\w3[7][26] ), .B(n6944), .Z(n6945) );
  XNOR U9576 ( .A(n6946), .B(n6945), .Z(\w1[8][2] ) );
  XNOR U9577 ( .A(\w3[7][24] ), .B(\w3[7][31] ), .Z(n7125) );
  XNOR U9578 ( .A(n6947), .B(n7125), .Z(n7086) );
  XOR U9579 ( .A(n7086), .B(key[1054]), .Z(n6950) );
  XNOR U9580 ( .A(\w3[7][6] ), .B(n6948), .Z(n6949) );
  XNOR U9581 ( .A(n6950), .B(n6949), .Z(\w1[8][30] ) );
  XOR U9582 ( .A(\w3[7][15] ), .B(\w3[7][23] ), .Z(n7123) );
  XOR U9583 ( .A(n7123), .B(key[1055]), .Z(n6952) );
  XNOR U9584 ( .A(n7164), .B(\w3[7][7] ), .Z(n6951) );
  XNOR U9585 ( .A(n6952), .B(n6951), .Z(\w1[8][31] ) );
  XOR U9586 ( .A(\w3[7][33] ), .B(\w3[7][57] ), .Z(n7007) );
  XOR U9587 ( .A(n7007), .B(key[1056]), .Z(n6954) );
  XOR U9588 ( .A(\w3[7][48] ), .B(\w3[7][56] ), .Z(n7068) );
  XNOR U9589 ( .A(n7068), .B(\w3[7][40] ), .Z(n6953) );
  XNOR U9590 ( .A(n6954), .B(n6953), .Z(\w1[8][32] ) );
  XOR U9591 ( .A(\w3[7][34] ), .B(\w3[7][58] ), .Z(n7015) );
  XOR U9592 ( .A(n7015), .B(key[1057]), .Z(n6956) );
  XOR U9593 ( .A(\w3[7][41] ), .B(\w3[7][49] ), .Z(n7039) );
  XNOR U9594 ( .A(\w3[7][57] ), .B(n7039), .Z(n6955) );
  XNOR U9595 ( .A(n6956), .B(n6955), .Z(\w1[8][33] ) );
  XOR U9596 ( .A(\w3[7][35] ), .B(\w3[7][59] ), .Z(n6986) );
  XOR U9597 ( .A(n6986), .B(key[1058]), .Z(n6958) );
  XOR U9598 ( .A(\w3[7][42] ), .B(\w3[7][50] ), .Z(n7043) );
  XNOR U9599 ( .A(\w3[7][58] ), .B(n7043), .Z(n6957) );
  XNOR U9600 ( .A(n6958), .B(n6957), .Z(\w1[8][34] ) );
  XOR U9601 ( .A(\w3[7][36] ), .B(\w3[7][32] ), .Z(n6988) );
  XOR U9602 ( .A(n6988), .B(key[1059]), .Z(n6961) );
  XOR U9603 ( .A(\w3[7][43] ), .B(\w3[7][51] ), .Z(n7014) );
  XNOR U9604 ( .A(\w3[7][56] ), .B(n7014), .Z(n6959) );
  XNOR U9605 ( .A(\w3[7][60] ), .B(n6959), .Z(n7048) );
  XNOR U9606 ( .A(\w3[7][59] ), .B(n7048), .Z(n6960) );
  XNOR U9607 ( .A(n6961), .B(n6960), .Z(\w1[8][35] ) );
  XOR U9608 ( .A(\w3[7][32] ), .B(\w3[7][37] ), .Z(n6993) );
  XOR U9609 ( .A(n6993), .B(key[1060]), .Z(n6965) );
  XOR U9610 ( .A(\w3[7][52] ), .B(\w3[7][61] ), .Z(n6963) );
  XNOR U9611 ( .A(\w3[7][56] ), .B(\w3[7][44] ), .Z(n6962) );
  XNOR U9612 ( .A(n6963), .B(n6962), .Z(n7056) );
  XNOR U9613 ( .A(\w3[7][60] ), .B(n7056), .Z(n6964) );
  XNOR U9614 ( .A(n6965), .B(n6964), .Z(\w1[8][36] ) );
  XOR U9615 ( .A(\w3[7][38] ), .B(\w3[7][62] ), .Z(n6999) );
  XOR U9616 ( .A(n6999), .B(key[1061]), .Z(n6967) );
  XOR U9617 ( .A(\w3[7][45] ), .B(\w3[7][53] ), .Z(n7059) );
  XNOR U9618 ( .A(\w3[7][61] ), .B(n7059), .Z(n6966) );
  XNOR U9619 ( .A(n6967), .B(n6966), .Z(\w1[8][37] ) );
  XOR U9620 ( .A(\w3[7][32] ), .B(\w3[7][39] ), .Z(n7000) );
  XOR U9621 ( .A(n7000), .B(key[1062]), .Z(n6969) );
  XOR U9622 ( .A(\w3[7][46] ), .B(\w3[7][54] ), .Z(n7025) );
  XNOR U9623 ( .A(\w3[7][56] ), .B(\w3[7][63] ), .Z(n6971) );
  XNOR U9624 ( .A(n7025), .B(n6971), .Z(n7064) );
  XNOR U9625 ( .A(\w3[7][62] ), .B(n7064), .Z(n6968) );
  XNOR U9626 ( .A(n6969), .B(n6968), .Z(\w1[8][38] ) );
  XOR U9627 ( .A(\w3[7][47] ), .B(\w3[7][55] ), .Z(n7067) );
  XNOR U9628 ( .A(n7067), .B(key[1063]), .Z(n6970) );
  XNOR U9629 ( .A(n6971), .B(n6970), .Z(n6972) );
  XNOR U9630 ( .A(\w3[7][32] ), .B(n6972), .Z(\w1[8][39] ) );
  XOR U9631 ( .A(n6973), .B(key[1027]), .Z(n6976) );
  XNOR U9632 ( .A(n6974), .B(\w3[7][27] ), .Z(n6975) );
  XNOR U9633 ( .A(n6976), .B(n6975), .Z(\w1[8][3] ) );
  XOR U9634 ( .A(\w3[7][32] ), .B(key[1064]), .Z(n6978) );
  XNOR U9635 ( .A(\w3[7][33] ), .B(\w3[7][41] ), .Z(n6977) );
  XNOR U9636 ( .A(n6978), .B(n6977), .Z(n6979) );
  XOR U9637 ( .A(n7068), .B(n6979), .Z(\w1[8][40] ) );
  XOR U9638 ( .A(\w3[7][42] ), .B(key[1065]), .Z(n6981) );
  XNOR U9639 ( .A(\w3[7][49] ), .B(\w3[7][34] ), .Z(n6980) );
  XNOR U9640 ( .A(n6981), .B(n6980), .Z(n6982) );
  XOR U9641 ( .A(n7007), .B(n6982), .Z(\w1[8][41] ) );
  XOR U9642 ( .A(\w3[7][43] ), .B(key[1066]), .Z(n6984) );
  XNOR U9643 ( .A(\w3[7][50] ), .B(\w3[7][35] ), .Z(n6983) );
  XNOR U9644 ( .A(n6984), .B(n6983), .Z(n6985) );
  XOR U9645 ( .A(n7015), .B(n6985), .Z(\w1[8][42] ) );
  XNOR U9646 ( .A(\w3[7][40] ), .B(n6986), .Z(n6987) );
  XNOR U9647 ( .A(\w3[7][44] ), .B(n6987), .Z(n7018) );
  XOR U9648 ( .A(n7018), .B(key[1067]), .Z(n6990) );
  XNOR U9649 ( .A(\w3[7][51] ), .B(n6988), .Z(n6989) );
  XNOR U9650 ( .A(n6990), .B(n6989), .Z(\w1[8][43] ) );
  XOR U9651 ( .A(\w3[7][36] ), .B(\w3[7][45] ), .Z(n6992) );
  XNOR U9652 ( .A(\w3[7][40] ), .B(\w3[7][60] ), .Z(n6991) );
  XNOR U9653 ( .A(n6992), .B(n6991), .Z(n7021) );
  XOR U9654 ( .A(n7021), .B(key[1068]), .Z(n6995) );
  XNOR U9655 ( .A(\w3[7][52] ), .B(n6993), .Z(n6994) );
  XNOR U9656 ( .A(n6995), .B(n6994), .Z(\w1[8][44] ) );
  XOR U9657 ( .A(\w3[7][61] ), .B(\w3[7][37] ), .Z(n7024) );
  XOR U9658 ( .A(n7024), .B(key[1069]), .Z(n6997) );
  XNOR U9659 ( .A(\w3[7][38] ), .B(\w3[7][46] ), .Z(n6996) );
  XNOR U9660 ( .A(n6997), .B(n6996), .Z(n6998) );
  XOR U9661 ( .A(\w3[7][53] ), .B(n6998), .Z(\w1[8][45] ) );
  XNOR U9662 ( .A(\w3[7][40] ), .B(\w3[7][47] ), .Z(n7033) );
  XNOR U9663 ( .A(n6999), .B(n7033), .Z(n7028) );
  XOR U9664 ( .A(n7028), .B(key[1070]), .Z(n7002) );
  XNOR U9665 ( .A(\w3[7][54] ), .B(n7000), .Z(n7001) );
  XNOR U9666 ( .A(n7002), .B(n7001), .Z(\w1[8][46] ) );
  XOR U9667 ( .A(\w3[7][63] ), .B(\w3[7][39] ), .Z(n7031) );
  XOR U9668 ( .A(n7031), .B(key[1071]), .Z(n7004) );
  XOR U9669 ( .A(\w3[7][40] ), .B(\w3[7][32] ), .Z(n7035) );
  XNOR U9670 ( .A(\w3[7][55] ), .B(n7035), .Z(n7003) );
  XNOR U9671 ( .A(n7004), .B(n7003), .Z(\w1[8][47] ) );
  XOR U9672 ( .A(n7035), .B(key[1072]), .Z(n7006) );
  XNOR U9673 ( .A(\w3[7][56] ), .B(n7039), .Z(n7005) );
  XNOR U9674 ( .A(n7006), .B(n7005), .Z(\w1[8][48] ) );
  XOR U9675 ( .A(n7043), .B(key[1073]), .Z(n7009) );
  XNOR U9676 ( .A(n7007), .B(\w3[7][41] ), .Z(n7008) );
  XNOR U9677 ( .A(n7009), .B(n7008), .Z(\w1[8][49] ) );
  XOR U9678 ( .A(n7010), .B(key[1028]), .Z(n7013) );
  XNOR U9679 ( .A(n7011), .B(\w3[7][28] ), .Z(n7012) );
  XNOR U9680 ( .A(n7013), .B(n7012), .Z(\w1[8][4] ) );
  XOR U9681 ( .A(n7014), .B(key[1074]), .Z(n7017) );
  XNOR U9682 ( .A(n7015), .B(\w3[7][42] ), .Z(n7016) );
  XNOR U9683 ( .A(n7017), .B(n7016), .Z(\w1[8][50] ) );
  XOR U9684 ( .A(\w3[7][48] ), .B(\w3[7][52] ), .Z(n7047) );
  XOR U9685 ( .A(n7047), .B(key[1075]), .Z(n7020) );
  XNOR U9686 ( .A(\w3[7][43] ), .B(n7018), .Z(n7019) );
  XNOR U9687 ( .A(n7020), .B(n7019), .Z(\w1[8][51] ) );
  XOR U9688 ( .A(\w3[7][48] ), .B(\w3[7][53] ), .Z(n7055) );
  XOR U9689 ( .A(n7055), .B(key[1076]), .Z(n7023) );
  XNOR U9690 ( .A(\w3[7][44] ), .B(n7021), .Z(n7022) );
  XNOR U9691 ( .A(n7023), .B(n7022), .Z(\w1[8][52] ) );
  XOR U9692 ( .A(n7024), .B(key[1077]), .Z(n7027) );
  XNOR U9693 ( .A(\w3[7][45] ), .B(n7025), .Z(n7026) );
  XNOR U9694 ( .A(n7027), .B(n7026), .Z(\w1[8][53] ) );
  XOR U9695 ( .A(\w3[7][48] ), .B(\w3[7][55] ), .Z(n7063) );
  XOR U9696 ( .A(n7063), .B(key[1078]), .Z(n7030) );
  XNOR U9697 ( .A(\w3[7][46] ), .B(n7028), .Z(n7029) );
  XNOR U9698 ( .A(n7030), .B(n7029), .Z(\w1[8][54] ) );
  XNOR U9699 ( .A(n7031), .B(key[1079]), .Z(n7032) );
  XNOR U9700 ( .A(n7033), .B(n7032), .Z(n7034) );
  XNOR U9701 ( .A(\w3[7][48] ), .B(n7034), .Z(\w1[8][55] ) );
  XOR U9702 ( .A(n7035), .B(key[1080]), .Z(n7037) );
  XNOR U9703 ( .A(\w3[7][48] ), .B(\w3[7][49] ), .Z(n7036) );
  XNOR U9704 ( .A(n7037), .B(n7036), .Z(n7038) );
  XOR U9705 ( .A(\w3[7][57] ), .B(n7038), .Z(\w1[8][56] ) );
  XOR U9706 ( .A(\w3[7][50] ), .B(key[1081]), .Z(n7041) );
  XNOR U9707 ( .A(n7039), .B(\w3[7][58] ), .Z(n7040) );
  XNOR U9708 ( .A(n7041), .B(n7040), .Z(n7042) );
  XOR U9709 ( .A(\w3[7][33] ), .B(n7042), .Z(\w1[8][57] ) );
  XOR U9710 ( .A(\w3[7][51] ), .B(key[1082]), .Z(n7045) );
  XNOR U9711 ( .A(n7043), .B(\w3[7][59] ), .Z(n7044) );
  XNOR U9712 ( .A(n7045), .B(n7044), .Z(n7046) );
  XOR U9713 ( .A(\w3[7][34] ), .B(n7046), .Z(\w1[8][58] ) );
  XOR U9714 ( .A(n7047), .B(key[1083]), .Z(n7050) );
  XNOR U9715 ( .A(\w3[7][35] ), .B(n7048), .Z(n7049) );
  XNOR U9716 ( .A(n7050), .B(n7049), .Z(\w1[8][59] ) );
  XOR U9717 ( .A(n7051), .B(key[1029]), .Z(n7054) );
  XNOR U9718 ( .A(\w3[7][29] ), .B(n7052), .Z(n7053) );
  XNOR U9719 ( .A(n7054), .B(n7053), .Z(\w1[8][5] ) );
  XOR U9720 ( .A(n7055), .B(key[1084]), .Z(n7058) );
  XNOR U9721 ( .A(\w3[7][36] ), .B(n7056), .Z(n7057) );
  XNOR U9722 ( .A(n7058), .B(n7057), .Z(\w1[8][60] ) );
  XOR U9723 ( .A(\w3[7][54] ), .B(key[1085]), .Z(n7061) );
  XNOR U9724 ( .A(n7059), .B(\w3[7][62] ), .Z(n7060) );
  XNOR U9725 ( .A(n7061), .B(n7060), .Z(n7062) );
  XOR U9726 ( .A(\w3[7][37] ), .B(n7062), .Z(\w1[8][61] ) );
  XOR U9727 ( .A(n7063), .B(key[1086]), .Z(n7066) );
  XNOR U9728 ( .A(\w3[7][38] ), .B(n7064), .Z(n7065) );
  XNOR U9729 ( .A(n7066), .B(n7065), .Z(\w1[8][62] ) );
  XOR U9730 ( .A(n7067), .B(key[1087]), .Z(n7070) );
  XNOR U9731 ( .A(n7068), .B(\w3[7][39] ), .Z(n7069) );
  XNOR U9732 ( .A(n7070), .B(n7069), .Z(\w1[8][63] ) );
  XOR U9733 ( .A(\w3[7][65] ), .B(\w3[7][89] ), .Z(n7129) );
  XOR U9734 ( .A(n7129), .B(key[1088]), .Z(n7072) );
  XOR U9735 ( .A(\w3[7][80] ), .B(\w3[7][88] ), .Z(n7186) );
  XNOR U9736 ( .A(n7186), .B(\w3[7][72] ), .Z(n7071) );
  XNOR U9737 ( .A(n7072), .B(n7071), .Z(\w1[8][64] ) );
  XOR U9738 ( .A(\w3[7][66] ), .B(\w3[7][90] ), .Z(n7133) );
  XOR U9739 ( .A(n7133), .B(key[1089]), .Z(n7074) );
  XOR U9740 ( .A(\w3[7][73] ), .B(\w3[7][81] ), .Z(n7157) );
  XNOR U9741 ( .A(\w3[7][89] ), .B(n7157), .Z(n7073) );
  XNOR U9742 ( .A(n7074), .B(n7073), .Z(\w1[8][65] ) );
  XOR U9743 ( .A(\w3[7][67] ), .B(\w3[7][91] ), .Z(n7104) );
  XOR U9744 ( .A(n7104), .B(key[1090]), .Z(n7076) );
  XOR U9745 ( .A(\w3[7][74] ), .B(\w3[7][82] ), .Z(n7165) );
  XNOR U9746 ( .A(\w3[7][90] ), .B(n7165), .Z(n7075) );
  XNOR U9747 ( .A(n7076), .B(n7075), .Z(\w1[8][66] ) );
  XOR U9748 ( .A(\w3[7][68] ), .B(\w3[7][64] ), .Z(n7106) );
  XOR U9749 ( .A(n7106), .B(key[1091]), .Z(n7079) );
  XOR U9750 ( .A(\w3[7][75] ), .B(\w3[7][83] ), .Z(n7132) );
  XNOR U9751 ( .A(\w3[7][88] ), .B(n7132), .Z(n7077) );
  XNOR U9752 ( .A(\w3[7][92] ), .B(n7077), .Z(n7170) );
  XNOR U9753 ( .A(\w3[7][91] ), .B(n7170), .Z(n7078) );
  XNOR U9754 ( .A(n7079), .B(n7078), .Z(\w1[8][67] ) );
  XOR U9755 ( .A(\w3[7][64] ), .B(\w3[7][69] ), .Z(n7111) );
  XOR U9756 ( .A(n7111), .B(key[1092]), .Z(n7083) );
  XOR U9757 ( .A(\w3[7][84] ), .B(\w3[7][93] ), .Z(n7081) );
  XNOR U9758 ( .A(\w3[7][88] ), .B(\w3[7][76] ), .Z(n7080) );
  XNOR U9759 ( .A(n7081), .B(n7080), .Z(n7174) );
  XNOR U9760 ( .A(\w3[7][92] ), .B(n7174), .Z(n7082) );
  XNOR U9761 ( .A(n7083), .B(n7082), .Z(\w1[8][68] ) );
  XOR U9762 ( .A(\w3[7][70] ), .B(\w3[7][94] ), .Z(n7117) );
  XOR U9763 ( .A(n7117), .B(key[1093]), .Z(n7085) );
  XOR U9764 ( .A(\w3[7][77] ), .B(\w3[7][85] ), .Z(n7177) );
  XNOR U9765 ( .A(\w3[7][93] ), .B(n7177), .Z(n7084) );
  XNOR U9766 ( .A(n7085), .B(n7084), .Z(\w1[8][69] ) );
  XOR U9767 ( .A(n7086), .B(key[1030]), .Z(n7089) );
  XNOR U9768 ( .A(n7087), .B(\w3[7][30] ), .Z(n7088) );
  XNOR U9769 ( .A(n7089), .B(n7088), .Z(\w1[8][6] ) );
  XOR U9770 ( .A(\w3[7][64] ), .B(\w3[7][71] ), .Z(n7118) );
  XOR U9771 ( .A(n7118), .B(key[1094]), .Z(n7091) );
  XOR U9772 ( .A(\w3[7][78] ), .B(\w3[7][86] ), .Z(n7143) );
  XNOR U9773 ( .A(\w3[7][88] ), .B(\w3[7][95] ), .Z(n7093) );
  XNOR U9774 ( .A(n7143), .B(n7093), .Z(n7182) );
  XNOR U9775 ( .A(\w3[7][94] ), .B(n7182), .Z(n7090) );
  XNOR U9776 ( .A(n7091), .B(n7090), .Z(\w1[8][70] ) );
  XOR U9777 ( .A(\w3[7][79] ), .B(\w3[7][87] ), .Z(n7185) );
  XNOR U9778 ( .A(n7185), .B(key[1095]), .Z(n7092) );
  XNOR U9779 ( .A(n7093), .B(n7092), .Z(n7094) );
  XNOR U9780 ( .A(\w3[7][64] ), .B(n7094), .Z(\w1[8][71] ) );
  XOR U9781 ( .A(\w3[7][64] ), .B(key[1096]), .Z(n7096) );
  XNOR U9782 ( .A(\w3[7][65] ), .B(\w3[7][73] ), .Z(n7095) );
  XNOR U9783 ( .A(n7096), .B(n7095), .Z(n7097) );
  XOR U9784 ( .A(n7186), .B(n7097), .Z(\w1[8][72] ) );
  XOR U9785 ( .A(\w3[7][74] ), .B(key[1097]), .Z(n7099) );
  XNOR U9786 ( .A(\w3[7][81] ), .B(\w3[7][66] ), .Z(n7098) );
  XNOR U9787 ( .A(n7099), .B(n7098), .Z(n7100) );
  XOR U9788 ( .A(n7129), .B(n7100), .Z(\w1[8][73] ) );
  XOR U9789 ( .A(\w3[7][75] ), .B(key[1098]), .Z(n7102) );
  XNOR U9790 ( .A(\w3[7][82] ), .B(\w3[7][67] ), .Z(n7101) );
  XNOR U9791 ( .A(n7102), .B(n7101), .Z(n7103) );
  XOR U9792 ( .A(n7133), .B(n7103), .Z(\w1[8][74] ) );
  XNOR U9793 ( .A(\w3[7][72] ), .B(n7104), .Z(n7105) );
  XNOR U9794 ( .A(\w3[7][76] ), .B(n7105), .Z(n7136) );
  XOR U9795 ( .A(n7136), .B(key[1099]), .Z(n7108) );
  XNOR U9796 ( .A(\w3[7][83] ), .B(n7106), .Z(n7107) );
  XNOR U9797 ( .A(n7108), .B(n7107), .Z(\w1[8][75] ) );
  XOR U9798 ( .A(\w3[7][68] ), .B(\w3[7][77] ), .Z(n7110) );
  XNOR U9799 ( .A(\w3[7][72] ), .B(\w3[7][92] ), .Z(n7109) );
  XNOR U9800 ( .A(n7110), .B(n7109), .Z(n7139) );
  XOR U9801 ( .A(n7139), .B(key[1100]), .Z(n7113) );
  XNOR U9802 ( .A(\w3[7][84] ), .B(n7111), .Z(n7112) );
  XNOR U9803 ( .A(n7113), .B(n7112), .Z(\w1[8][76] ) );
  XOR U9804 ( .A(\w3[7][93] ), .B(\w3[7][69] ), .Z(n7142) );
  XOR U9805 ( .A(n7142), .B(key[1101]), .Z(n7115) );
  XNOR U9806 ( .A(\w3[7][70] ), .B(\w3[7][78] ), .Z(n7114) );
  XNOR U9807 ( .A(n7115), .B(n7114), .Z(n7116) );
  XOR U9808 ( .A(\w3[7][85] ), .B(n7116), .Z(\w1[8][77] ) );
  XNOR U9809 ( .A(\w3[7][72] ), .B(\w3[7][79] ), .Z(n7151) );
  XNOR U9810 ( .A(n7117), .B(n7151), .Z(n7146) );
  XOR U9811 ( .A(n7146), .B(key[1102]), .Z(n7120) );
  XNOR U9812 ( .A(\w3[7][86] ), .B(n7118), .Z(n7119) );
  XNOR U9813 ( .A(n7120), .B(n7119), .Z(\w1[8][78] ) );
  XOR U9814 ( .A(\w3[7][95] ), .B(\w3[7][71] ), .Z(n7149) );
  XOR U9815 ( .A(n7149), .B(key[1103]), .Z(n7122) );
  XOR U9816 ( .A(\w3[7][72] ), .B(\w3[7][64] ), .Z(n7153) );
  XNOR U9817 ( .A(\w3[7][87] ), .B(n7153), .Z(n7121) );
  XNOR U9818 ( .A(n7122), .B(n7121), .Z(\w1[8][79] ) );
  XNOR U9819 ( .A(n7123), .B(key[1031]), .Z(n7124) );
  XNOR U9820 ( .A(n7125), .B(n7124), .Z(n7126) );
  XNOR U9821 ( .A(\w3[7][0] ), .B(n7126), .Z(\w1[8][7] ) );
  XOR U9822 ( .A(n7153), .B(key[1104]), .Z(n7128) );
  XNOR U9823 ( .A(\w3[7][88] ), .B(n7157), .Z(n7127) );
  XNOR U9824 ( .A(n7128), .B(n7127), .Z(\w1[8][80] ) );
  XOR U9825 ( .A(n7165), .B(key[1105]), .Z(n7131) );
  XNOR U9826 ( .A(n7129), .B(\w3[7][73] ), .Z(n7130) );
  XNOR U9827 ( .A(n7131), .B(n7130), .Z(\w1[8][81] ) );
  XOR U9828 ( .A(n7132), .B(key[1106]), .Z(n7135) );
  XNOR U9829 ( .A(n7133), .B(\w3[7][74] ), .Z(n7134) );
  XNOR U9830 ( .A(n7135), .B(n7134), .Z(\w1[8][82] ) );
  XOR U9831 ( .A(\w3[7][80] ), .B(\w3[7][84] ), .Z(n7169) );
  XOR U9832 ( .A(n7169), .B(key[1107]), .Z(n7138) );
  XNOR U9833 ( .A(\w3[7][75] ), .B(n7136), .Z(n7137) );
  XNOR U9834 ( .A(n7138), .B(n7137), .Z(\w1[8][83] ) );
  XOR U9835 ( .A(\w3[7][80] ), .B(\w3[7][85] ), .Z(n7173) );
  XOR U9836 ( .A(n7173), .B(key[1108]), .Z(n7141) );
  XNOR U9837 ( .A(\w3[7][76] ), .B(n7139), .Z(n7140) );
  XNOR U9838 ( .A(n7141), .B(n7140), .Z(\w1[8][84] ) );
  XOR U9839 ( .A(n7142), .B(key[1109]), .Z(n7145) );
  XNOR U9840 ( .A(\w3[7][77] ), .B(n7143), .Z(n7144) );
  XNOR U9841 ( .A(n7145), .B(n7144), .Z(\w1[8][85] ) );
  XOR U9842 ( .A(\w3[7][80] ), .B(\w3[7][87] ), .Z(n7181) );
  XOR U9843 ( .A(n7181), .B(key[1110]), .Z(n7148) );
  XNOR U9844 ( .A(\w3[7][78] ), .B(n7146), .Z(n7147) );
  XNOR U9845 ( .A(n7148), .B(n7147), .Z(\w1[8][86] ) );
  XNOR U9846 ( .A(n7149), .B(key[1111]), .Z(n7150) );
  XNOR U9847 ( .A(n7151), .B(n7150), .Z(n7152) );
  XNOR U9848 ( .A(\w3[7][80] ), .B(n7152), .Z(\w1[8][87] ) );
  XOR U9849 ( .A(n7153), .B(key[1112]), .Z(n7155) );
  XNOR U9850 ( .A(\w3[7][80] ), .B(\w3[7][81] ), .Z(n7154) );
  XNOR U9851 ( .A(n7155), .B(n7154), .Z(n7156) );
  XOR U9852 ( .A(\w3[7][89] ), .B(n7156), .Z(\w1[8][88] ) );
  XOR U9853 ( .A(\w3[7][82] ), .B(key[1113]), .Z(n7159) );
  XNOR U9854 ( .A(n7157), .B(\w3[7][90] ), .Z(n7158) );
  XNOR U9855 ( .A(n7159), .B(n7158), .Z(n7160) );
  XOR U9856 ( .A(\w3[7][65] ), .B(n7160), .Z(\w1[8][89] ) );
  XOR U9857 ( .A(\w3[7][9] ), .B(key[1032]), .Z(n7162) );
  XNOR U9858 ( .A(\w3[7][1] ), .B(\w3[7][0] ), .Z(n7161) );
  XNOR U9859 ( .A(n7162), .B(n7161), .Z(n7163) );
  XOR U9860 ( .A(n7164), .B(n7163), .Z(\w1[8][8] ) );
  XOR U9861 ( .A(\w3[7][83] ), .B(key[1114]), .Z(n7167) );
  XNOR U9862 ( .A(n7165), .B(\w3[7][91] ), .Z(n7166) );
  XNOR U9863 ( .A(n7167), .B(n7166), .Z(n7168) );
  XOR U9864 ( .A(\w3[7][66] ), .B(n7168), .Z(\w1[8][90] ) );
  XOR U9865 ( .A(n7169), .B(key[1115]), .Z(n7172) );
  XNOR U9866 ( .A(\w3[7][67] ), .B(n7170), .Z(n7171) );
  XNOR U9867 ( .A(n7172), .B(n7171), .Z(\w1[8][91] ) );
  XOR U9868 ( .A(n7173), .B(key[1116]), .Z(n7176) );
  XNOR U9869 ( .A(\w3[7][68] ), .B(n7174), .Z(n7175) );
  XNOR U9870 ( .A(n7176), .B(n7175), .Z(\w1[8][92] ) );
  XOR U9871 ( .A(\w3[7][86] ), .B(key[1117]), .Z(n7179) );
  XNOR U9872 ( .A(n7177), .B(\w3[7][94] ), .Z(n7178) );
  XNOR U9873 ( .A(n7179), .B(n7178), .Z(n7180) );
  XOR U9874 ( .A(\w3[7][69] ), .B(n7180), .Z(\w1[8][93] ) );
  XOR U9875 ( .A(n7181), .B(key[1118]), .Z(n7184) );
  XNOR U9876 ( .A(\w3[7][70] ), .B(n7182), .Z(n7183) );
  XNOR U9877 ( .A(n7184), .B(n7183), .Z(\w1[8][94] ) );
  XOR U9878 ( .A(n7185), .B(key[1119]), .Z(n7188) );
  XNOR U9879 ( .A(n7186), .B(\w3[7][71] ), .Z(n7187) );
  XNOR U9880 ( .A(n7188), .B(n7187), .Z(\w1[8][95] ) );
  XOR U9881 ( .A(n7189), .B(key[1120]), .Z(n7192) );
  XOR U9882 ( .A(n7190), .B(\w3[7][104] ), .Z(n7191) );
  XNOR U9883 ( .A(n7192), .B(n7191), .Z(\w1[8][96] ) );
  XOR U9884 ( .A(n7193), .B(key[1121]), .Z(n7196) );
  XNOR U9885 ( .A(\w3[7][121] ), .B(n7194), .Z(n7195) );
  XNOR U9886 ( .A(n7196), .B(n7195), .Z(\w1[8][97] ) );
  XOR U9887 ( .A(n7197), .B(key[1122]), .Z(n7200) );
  XNOR U9888 ( .A(\w3[7][122] ), .B(n7198), .Z(n7199) );
  XNOR U9889 ( .A(n7200), .B(n7199), .Z(\w1[8][98] ) );
  XOR U9890 ( .A(n7201), .B(key[1123]), .Z(n7204) );
  XNOR U9891 ( .A(n7202), .B(\w3[7][123] ), .Z(n7203) );
  XNOR U9892 ( .A(n7204), .B(n7203), .Z(\w1[8][99] ) );
  XOR U9893 ( .A(\w3[7][10] ), .B(key[1033]), .Z(n7206) );
  XNOR U9894 ( .A(\w3[7][2] ), .B(\w3[7][17] ), .Z(n7205) );
  XNOR U9895 ( .A(n7206), .B(n7205), .Z(n7207) );
  XOR U9896 ( .A(n7208), .B(n7207), .Z(\w1[8][9] ) );
  XOR U9897 ( .A(\w3[8][8] ), .B(key[1152]), .Z(n7210) );
  XOR U9898 ( .A(\w3[8][1] ), .B(\w3[8][25] ), .Z(n7632) );
  XOR U9899 ( .A(\w3[8][16] ), .B(\w3[8][24] ), .Z(n7588) );
  XNOR U9900 ( .A(n7632), .B(n7588), .Z(n7209) );
  XNOR U9901 ( .A(n7210), .B(n7209), .Z(\w1[9][0] ) );
  XOR U9902 ( .A(\w3[8][96] ), .B(\w3[8][101] ), .Z(n7236) );
  XOR U9903 ( .A(n7236), .B(key[1252]), .Z(n7214) );
  XOR U9904 ( .A(\w3[8][116] ), .B(\w3[8][125] ), .Z(n7212) );
  XNOR U9905 ( .A(\w3[8][120] ), .B(\w3[8][108] ), .Z(n7211) );
  XNOR U9906 ( .A(n7212), .B(n7211), .Z(n7293) );
  XNOR U9907 ( .A(\w3[8][124] ), .B(n7293), .Z(n7213) );
  XNOR U9908 ( .A(n7214), .B(n7213), .Z(\w1[9][100] ) );
  XOR U9909 ( .A(\w3[8][102] ), .B(\w3[8][126] ), .Z(n7245) );
  XOR U9910 ( .A(n7245), .B(key[1253]), .Z(n7216) );
  XOR U9911 ( .A(\w3[8][109] ), .B(\w3[8][117] ), .Z(n7299) );
  XNOR U9912 ( .A(\w3[8][125] ), .B(n7299), .Z(n7215) );
  XNOR U9913 ( .A(n7216), .B(n7215), .Z(\w1[9][101] ) );
  XOR U9914 ( .A(\w3[8][96] ), .B(\w3[8][103] ), .Z(n7246) );
  XOR U9915 ( .A(n7246), .B(key[1254]), .Z(n7218) );
  XOR U9916 ( .A(\w3[8][110] ), .B(\w3[8][118] ), .Z(n7264) );
  XNOR U9917 ( .A(\w3[8][120] ), .B(\w3[8][127] ), .Z(n7220) );
  XNOR U9918 ( .A(n7264), .B(n7220), .Z(n7301) );
  XNOR U9919 ( .A(\w3[8][126] ), .B(n7301), .Z(n7217) );
  XNOR U9920 ( .A(n7218), .B(n7217), .Z(\w1[9][102] ) );
  XOR U9921 ( .A(\w3[8][111] ), .B(\w3[8][119] ), .Z(n7304) );
  XNOR U9922 ( .A(n7304), .B(key[1255]), .Z(n7219) );
  XNOR U9923 ( .A(n7220), .B(n7219), .Z(n7221) );
  XNOR U9924 ( .A(\w3[8][96] ), .B(n7221), .Z(\w1[9][103] ) );
  XOR U9925 ( .A(key[1256]), .B(\w3[8][105] ), .Z(n7223) );
  XNOR U9926 ( .A(\w3[8][96] ), .B(\w3[8][97] ), .Z(n7222) );
  XNOR U9927 ( .A(n7223), .B(n7222), .Z(n7224) );
  XNOR U9928 ( .A(\w3[8][120] ), .B(\w3[8][112] ), .Z(n7614) );
  XNOR U9929 ( .A(n7224), .B(n7614), .Z(\w1[9][104] ) );
  XOR U9930 ( .A(\w3[8][106] ), .B(\w3[8][98] ), .Z(n7226) );
  XOR U9931 ( .A(\w3[8][97] ), .B(\w3[8][121] ), .Z(n7613) );
  XNOR U9932 ( .A(n7613), .B(key[1257]), .Z(n7225) );
  XNOR U9933 ( .A(n7226), .B(n7225), .Z(n7227) );
  XOR U9934 ( .A(\w3[8][113] ), .B(n7227), .Z(\w1[9][105] ) );
  XOR U9935 ( .A(\w3[8][107] ), .B(\w3[8][114] ), .Z(n7229) );
  XOR U9936 ( .A(\w3[8][98] ), .B(\w3[8][122] ), .Z(n7618) );
  XNOR U9937 ( .A(n7618), .B(key[1258]), .Z(n7228) );
  XNOR U9938 ( .A(n7229), .B(n7228), .Z(n7230) );
  XOR U9939 ( .A(\w3[8][99] ), .B(n7230), .Z(\w1[9][106] ) );
  XOR U9940 ( .A(\w3[8][99] ), .B(\w3[8][123] ), .Z(n7622) );
  XNOR U9941 ( .A(\w3[8][108] ), .B(n7622), .Z(n7231) );
  XNOR U9942 ( .A(\w3[8][104] ), .B(n7231), .Z(n7257) );
  XOR U9943 ( .A(n7257), .B(key[1259]), .Z(n7233) );
  XOR U9944 ( .A(\w3[8][96] ), .B(\w3[8][100] ), .Z(n7626) );
  XNOR U9945 ( .A(\w3[8][115] ), .B(n7626), .Z(n7232) );
  XNOR U9946 ( .A(n7233), .B(n7232), .Z(\w1[9][107] ) );
  XOR U9947 ( .A(\w3[8][100] ), .B(\w3[8][104] ), .Z(n7235) );
  XNOR U9948 ( .A(\w3[8][124] ), .B(\w3[8][109] ), .Z(n7234) );
  XNOR U9949 ( .A(n7235), .B(n7234), .Z(n7260) );
  XOR U9950 ( .A(n7260), .B(key[1260]), .Z(n7238) );
  XNOR U9951 ( .A(\w3[8][116] ), .B(n7236), .Z(n7237) );
  XNOR U9952 ( .A(n7238), .B(n7237), .Z(\w1[9][108] ) );
  XOR U9953 ( .A(\w3[8][125] ), .B(\w3[8][101] ), .Z(n7263) );
  XOR U9954 ( .A(n7263), .B(key[1261]), .Z(n7240) );
  XNOR U9955 ( .A(\w3[8][102] ), .B(\w3[8][110] ), .Z(n7239) );
  XNOR U9956 ( .A(n7240), .B(n7239), .Z(n7241) );
  XOR U9957 ( .A(\w3[8][117] ), .B(n7241), .Z(\w1[9][109] ) );
  XOR U9958 ( .A(\w3[8][11] ), .B(\w3[8][3] ), .Z(n7243) );
  XOR U9959 ( .A(\w3[8][2] ), .B(\w3[8][26] ), .Z(n7327) );
  XNOR U9960 ( .A(n7327), .B(key[1162]), .Z(n7242) );
  XNOR U9961 ( .A(n7243), .B(n7242), .Z(n7244) );
  XOR U9962 ( .A(\w3[8][18] ), .B(n7244), .Z(\w1[9][10] ) );
  XNOR U9963 ( .A(\w3[8][111] ), .B(\w3[8][104] ), .Z(n7272) );
  XNOR U9964 ( .A(n7245), .B(n7272), .Z(n7267) );
  XOR U9965 ( .A(n7267), .B(key[1262]), .Z(n7248) );
  XNOR U9966 ( .A(\w3[8][118] ), .B(n7246), .Z(n7247) );
  XNOR U9967 ( .A(n7248), .B(n7247), .Z(\w1[9][110] ) );
  XOR U9968 ( .A(\w3[8][127] ), .B(\w3[8][103] ), .Z(n7270) );
  XOR U9969 ( .A(n7270), .B(key[1263]), .Z(n7250) );
  XOR U9970 ( .A(\w3[8][96] ), .B(\w3[8][104] ), .Z(n7277) );
  XNOR U9971 ( .A(\w3[8][119] ), .B(n7277), .Z(n7249) );
  XNOR U9972 ( .A(n7250), .B(n7249), .Z(\w1[9][111] ) );
  XOR U9973 ( .A(\w3[8][105] ), .B(\w3[8][113] ), .Z(n7280) );
  XOR U9974 ( .A(n7280), .B(key[1264]), .Z(n7252) );
  XNOR U9975 ( .A(\w3[8][120] ), .B(n7277), .Z(n7251) );
  XNOR U9976 ( .A(n7252), .B(n7251), .Z(\w1[9][112] ) );
  XOR U9977 ( .A(\w3[8][106] ), .B(\w3[8][114] ), .Z(n7283) );
  XOR U9978 ( .A(n7283), .B(key[1265]), .Z(n7254) );
  XNOR U9979 ( .A(\w3[8][105] ), .B(n7613), .Z(n7253) );
  XNOR U9980 ( .A(n7254), .B(n7253), .Z(\w1[9][113] ) );
  XOR U9981 ( .A(\w3[8][107] ), .B(\w3[8][115] ), .Z(n7288) );
  XOR U9982 ( .A(n7288), .B(key[1266]), .Z(n7256) );
  XNOR U9983 ( .A(\w3[8][106] ), .B(n7618), .Z(n7255) );
  XNOR U9984 ( .A(n7256), .B(n7255), .Z(\w1[9][114] ) );
  XOR U9985 ( .A(\w3[8][116] ), .B(\w3[8][112] ), .Z(n7289) );
  XOR U9986 ( .A(n7289), .B(key[1267]), .Z(n7259) );
  XNOR U9987 ( .A(\w3[8][107] ), .B(n7257), .Z(n7258) );
  XNOR U9988 ( .A(n7259), .B(n7258), .Z(\w1[9][115] ) );
  XOR U9989 ( .A(\w3[8][117] ), .B(\w3[8][112] ), .Z(n7292) );
  XOR U9990 ( .A(n7292), .B(key[1268]), .Z(n7262) );
  XNOR U9991 ( .A(\w3[8][108] ), .B(n7260), .Z(n7261) );
  XNOR U9992 ( .A(n7262), .B(n7261), .Z(\w1[9][116] ) );
  XOR U9993 ( .A(n7263), .B(key[1269]), .Z(n7266) );
  XNOR U9994 ( .A(\w3[8][109] ), .B(n7264), .Z(n7265) );
  XNOR U9995 ( .A(n7266), .B(n7265), .Z(\w1[9][117] ) );
  XOR U9996 ( .A(\w3[8][119] ), .B(\w3[8][112] ), .Z(n7300) );
  XOR U9997 ( .A(n7300), .B(key[1270]), .Z(n7269) );
  XNOR U9998 ( .A(\w3[8][110] ), .B(n7267), .Z(n7268) );
  XNOR U9999 ( .A(n7269), .B(n7268), .Z(\w1[9][118] ) );
  XNOR U10000 ( .A(n7270), .B(key[1271]), .Z(n7271) );
  XNOR U10001 ( .A(n7272), .B(n7271), .Z(n7273) );
  XNOR U10002 ( .A(\w3[8][112] ), .B(n7273), .Z(\w1[9][119] ) );
  XOR U10003 ( .A(\w3[8][3] ), .B(\w3[8][27] ), .Z(n7368) );
  XNOR U10004 ( .A(\w3[8][8] ), .B(\w3[8][12] ), .Z(n7274) );
  XNOR U10005 ( .A(n7368), .B(n7274), .Z(n7324) );
  XOR U10006 ( .A(n7324), .B(key[1163]), .Z(n7276) );
  XOR U10007 ( .A(\w3[8][0] ), .B(\w3[8][4] ), .Z(n7398) );
  XNOR U10008 ( .A(\w3[8][19] ), .B(n7398), .Z(n7275) );
  XNOR U10009 ( .A(n7276), .B(n7275), .Z(\w1[9][11] ) );
  XOR U10010 ( .A(\w3[8][113] ), .B(\w3[8][121] ), .Z(n7617) );
  XOR U10011 ( .A(n7617), .B(key[1272]), .Z(n7279) );
  XNOR U10012 ( .A(\w3[8][112] ), .B(n7277), .Z(n7278) );
  XNOR U10013 ( .A(n7279), .B(n7278), .Z(\w1[9][120] ) );
  XOR U10014 ( .A(\w3[8][122] ), .B(\w3[8][114] ), .Z(n7621) );
  XOR U10015 ( .A(n7621), .B(key[1273]), .Z(n7282) );
  XNOR U10016 ( .A(\w3[8][97] ), .B(n7280), .Z(n7281) );
  XNOR U10017 ( .A(n7282), .B(n7281), .Z(\w1[9][121] ) );
  XOR U10018 ( .A(n7283), .B(key[1274]), .Z(n7285) );
  XNOR U10019 ( .A(\w3[8][115] ), .B(\w3[8][123] ), .Z(n7284) );
  XNOR U10020 ( .A(n7285), .B(n7284), .Z(n7286) );
  XOR U10021 ( .A(\w3[8][98] ), .B(n7286), .Z(\w1[9][122] ) );
  XNOR U10022 ( .A(\w3[8][124] ), .B(\w3[8][120] ), .Z(n7287) );
  XNOR U10023 ( .A(n7288), .B(n7287), .Z(n7625) );
  XOR U10024 ( .A(n7625), .B(key[1275]), .Z(n7291) );
  XNOR U10025 ( .A(\w3[8][99] ), .B(n7289), .Z(n7290) );
  XNOR U10026 ( .A(n7291), .B(n7290), .Z(\w1[9][123] ) );
  XOR U10027 ( .A(n7292), .B(key[1276]), .Z(n7295) );
  XNOR U10028 ( .A(n7293), .B(\w3[8][100] ), .Z(n7294) );
  XNOR U10029 ( .A(n7295), .B(n7294), .Z(\w1[9][124] ) );
  XOR U10030 ( .A(\w3[8][118] ), .B(key[1277]), .Z(n7297) );
  XNOR U10031 ( .A(\w3[8][101] ), .B(\w3[8][126] ), .Z(n7296) );
  XNOR U10032 ( .A(n7297), .B(n7296), .Z(n7298) );
  XOR U10033 ( .A(n7299), .B(n7298), .Z(\w1[9][125] ) );
  XOR U10034 ( .A(n7300), .B(key[1278]), .Z(n7303) );
  XNOR U10035 ( .A(\w3[8][102] ), .B(n7301), .Z(n7302) );
  XNOR U10036 ( .A(n7303), .B(n7302), .Z(\w1[9][126] ) );
  XNOR U10037 ( .A(n7304), .B(key[1279]), .Z(n7305) );
  XNOR U10038 ( .A(n7614), .B(n7305), .Z(n7306) );
  XNOR U10039 ( .A(\w3[8][103] ), .B(n7306), .Z(\w1[9][127] ) );
  XOR U10040 ( .A(\w3[8][13] ), .B(\w3[8][28] ), .Z(n7308) );
  XNOR U10041 ( .A(\w3[8][8] ), .B(\w3[8][4] ), .Z(n7307) );
  XNOR U10042 ( .A(n7308), .B(n7307), .Z(n7330) );
  XOR U10043 ( .A(n7330), .B(key[1164]), .Z(n7310) );
  XOR U10044 ( .A(\w3[8][0] ), .B(\w3[8][5] ), .Z(n7435) );
  XNOR U10045 ( .A(\w3[8][20] ), .B(n7435), .Z(n7309) );
  XNOR U10046 ( .A(n7310), .B(n7309), .Z(\w1[9][12] ) );
  XOR U10047 ( .A(\w3[8][14] ), .B(\w3[8][6] ), .Z(n7312) );
  XOR U10048 ( .A(\w3[8][5] ), .B(\w3[8][29] ), .Z(n7333) );
  XNOR U10049 ( .A(n7333), .B(key[1165]), .Z(n7311) );
  XNOR U10050 ( .A(n7312), .B(n7311), .Z(n7313) );
  XOR U10051 ( .A(\w3[8][21] ), .B(n7313), .Z(\w1[9][13] ) );
  XOR U10052 ( .A(\w3[8][6] ), .B(\w3[8][30] ), .Z(n7476) );
  XNOR U10053 ( .A(\w3[8][8] ), .B(\w3[8][15] ), .Z(n7341) );
  XNOR U10054 ( .A(n7476), .B(n7341), .Z(n7336) );
  XOR U10055 ( .A(n7336), .B(key[1166]), .Z(n7315) );
  XOR U10056 ( .A(\w3[8][0] ), .B(\w3[8][7] ), .Z(n7511) );
  XNOR U10057 ( .A(\w3[8][22] ), .B(n7511), .Z(n7314) );
  XNOR U10058 ( .A(n7315), .B(n7314), .Z(\w1[9][14] ) );
  XOR U10059 ( .A(\w3[8][7] ), .B(\w3[8][31] ), .Z(n7339) );
  XOR U10060 ( .A(n7339), .B(key[1167]), .Z(n7317) );
  XOR U10061 ( .A(\w3[8][8] ), .B(\w3[8][0] ), .Z(n7343) );
  XNOR U10062 ( .A(\w3[8][23] ), .B(n7343), .Z(n7316) );
  XNOR U10063 ( .A(n7317), .B(n7316), .Z(\w1[9][15] ) );
  XOR U10064 ( .A(\w3[8][17] ), .B(\w3[8][9] ), .Z(n7347) );
  XOR U10065 ( .A(n7347), .B(key[1168]), .Z(n7319) );
  XNOR U10066 ( .A(\w3[8][24] ), .B(n7343), .Z(n7318) );
  XNOR U10067 ( .A(n7319), .B(n7318), .Z(\w1[9][16] ) );
  XOR U10068 ( .A(\w3[8][18] ), .B(\w3[8][10] ), .Z(n7367) );
  XOR U10069 ( .A(n7367), .B(key[1169]), .Z(n7321) );
  XNOR U10070 ( .A(n7632), .B(\w3[8][9] ), .Z(n7320) );
  XNOR U10071 ( .A(n7321), .B(n7320), .Z(\w1[9][17] ) );
  XOR U10072 ( .A(\w3[8][11] ), .B(\w3[8][19] ), .Z(n7355) );
  XOR U10073 ( .A(n7355), .B(key[1170]), .Z(n7323) );
  XNOR U10074 ( .A(n7327), .B(\w3[8][10] ), .Z(n7322) );
  XNOR U10075 ( .A(n7323), .B(n7322), .Z(\w1[9][18] ) );
  XOR U10076 ( .A(\w3[8][16] ), .B(\w3[8][20] ), .Z(n7356) );
  XOR U10077 ( .A(n7356), .B(key[1171]), .Z(n7326) );
  XNOR U10078 ( .A(\w3[8][11] ), .B(n7324), .Z(n7325) );
  XNOR U10079 ( .A(n7326), .B(n7325), .Z(\w1[9][19] ) );
  XOR U10080 ( .A(n7347), .B(key[1153]), .Z(n7329) );
  XNOR U10081 ( .A(\w3[8][25] ), .B(n7327), .Z(n7328) );
  XNOR U10082 ( .A(n7329), .B(n7328), .Z(\w1[9][1] ) );
  XOR U10083 ( .A(\w3[8][16] ), .B(\w3[8][21] ), .Z(n7361) );
  XOR U10084 ( .A(n7361), .B(key[1172]), .Z(n7332) );
  XNOR U10085 ( .A(\w3[8][12] ), .B(n7330), .Z(n7331) );
  XNOR U10086 ( .A(n7332), .B(n7331), .Z(\w1[9][20] ) );
  XOR U10087 ( .A(\w3[8][14] ), .B(\w3[8][22] ), .Z(n7371) );
  XOR U10088 ( .A(n7371), .B(key[1173]), .Z(n7335) );
  XNOR U10089 ( .A(\w3[8][13] ), .B(n7333), .Z(n7334) );
  XNOR U10090 ( .A(n7335), .B(n7334), .Z(\w1[9][21] ) );
  XOR U10091 ( .A(\w3[8][16] ), .B(\w3[8][23] ), .Z(n7372) );
  XOR U10092 ( .A(n7372), .B(key[1174]), .Z(n7338) );
  XNOR U10093 ( .A(\w3[8][14] ), .B(n7336), .Z(n7337) );
  XNOR U10094 ( .A(n7338), .B(n7337), .Z(\w1[9][22] ) );
  XNOR U10095 ( .A(n7339), .B(key[1175]), .Z(n7340) );
  XNOR U10096 ( .A(n7341), .B(n7340), .Z(n7342) );
  XNOR U10097 ( .A(\w3[8][16] ), .B(n7342), .Z(\w1[9][23] ) );
  XOR U10098 ( .A(\w3[8][17] ), .B(key[1176]), .Z(n7345) );
  XNOR U10099 ( .A(\w3[8][25] ), .B(n7343), .Z(n7344) );
  XNOR U10100 ( .A(n7345), .B(n7344), .Z(n7346) );
  XOR U10101 ( .A(\w3[8][16] ), .B(n7346), .Z(\w1[9][24] ) );
  XOR U10102 ( .A(n7347), .B(key[1177]), .Z(n7349) );
  XNOR U10103 ( .A(\w3[8][1] ), .B(\w3[8][26] ), .Z(n7348) );
  XNOR U10104 ( .A(n7349), .B(n7348), .Z(n7350) );
  XOR U10105 ( .A(\w3[8][18] ), .B(n7350), .Z(\w1[9][25] ) );
  XOR U10106 ( .A(n7367), .B(key[1178]), .Z(n7352) );
  XNOR U10107 ( .A(\w3[8][2] ), .B(\w3[8][19] ), .Z(n7351) );
  XNOR U10108 ( .A(n7352), .B(n7351), .Z(n7353) );
  XOR U10109 ( .A(\w3[8][27] ), .B(n7353), .Z(\w1[9][26] ) );
  XNOR U10110 ( .A(\w3[8][24] ), .B(\w3[8][28] ), .Z(n7354) );
  XNOR U10111 ( .A(n7355), .B(n7354), .Z(n7397) );
  XOR U10112 ( .A(n7397), .B(key[1179]), .Z(n7358) );
  XNOR U10113 ( .A(\w3[8][3] ), .B(n7356), .Z(n7357) );
  XNOR U10114 ( .A(n7358), .B(n7357), .Z(\w1[9][27] ) );
  XOR U10115 ( .A(\w3[8][20] ), .B(\w3[8][29] ), .Z(n7360) );
  XNOR U10116 ( .A(\w3[8][24] ), .B(\w3[8][12] ), .Z(n7359) );
  XNOR U10117 ( .A(n7360), .B(n7359), .Z(n7434) );
  XOR U10118 ( .A(n7434), .B(key[1180]), .Z(n7363) );
  XNOR U10119 ( .A(\w3[8][4] ), .B(n7361), .Z(n7362) );
  XNOR U10120 ( .A(n7363), .B(n7362), .Z(\w1[9][28] ) );
  XOR U10121 ( .A(\w3[8][13] ), .B(\w3[8][21] ), .Z(n7475) );
  XOR U10122 ( .A(n7475), .B(key[1181]), .Z(n7365) );
  XNOR U10123 ( .A(\w3[8][22] ), .B(\w3[8][30] ), .Z(n7364) );
  XNOR U10124 ( .A(n7365), .B(n7364), .Z(n7366) );
  XOR U10125 ( .A(\w3[8][5] ), .B(n7366), .Z(\w1[9][29] ) );
  XOR U10126 ( .A(n7367), .B(key[1154]), .Z(n7370) );
  XNOR U10127 ( .A(\w3[8][26] ), .B(n7368), .Z(n7369) );
  XNOR U10128 ( .A(n7370), .B(n7369), .Z(\w1[9][2] ) );
  XNOR U10129 ( .A(\w3[8][24] ), .B(\w3[8][31] ), .Z(n7549) );
  XNOR U10130 ( .A(n7371), .B(n7549), .Z(n7510) );
  XOR U10131 ( .A(n7510), .B(key[1182]), .Z(n7374) );
  XNOR U10132 ( .A(\w3[8][6] ), .B(n7372), .Z(n7373) );
  XNOR U10133 ( .A(n7374), .B(n7373), .Z(\w1[9][30] ) );
  XOR U10134 ( .A(\w3[8][15] ), .B(\w3[8][23] ), .Z(n7547) );
  XOR U10135 ( .A(n7547), .B(key[1183]), .Z(n7376) );
  XNOR U10136 ( .A(n7588), .B(\w3[8][7] ), .Z(n7375) );
  XNOR U10137 ( .A(n7376), .B(n7375), .Z(\w1[9][31] ) );
  XOR U10138 ( .A(\w3[8][33] ), .B(\w3[8][57] ), .Z(n7431) );
  XOR U10139 ( .A(n7431), .B(key[1184]), .Z(n7378) );
  XOR U10140 ( .A(\w3[8][48] ), .B(\w3[8][56] ), .Z(n7492) );
  XNOR U10141 ( .A(n7492), .B(\w3[8][40] ), .Z(n7377) );
  XNOR U10142 ( .A(n7378), .B(n7377), .Z(\w1[9][32] ) );
  XOR U10143 ( .A(\w3[8][34] ), .B(\w3[8][58] ), .Z(n7439) );
  XOR U10144 ( .A(n7439), .B(key[1185]), .Z(n7380) );
  XOR U10145 ( .A(\w3[8][41] ), .B(\w3[8][49] ), .Z(n7466) );
  XNOR U10146 ( .A(\w3[8][57] ), .B(n7466), .Z(n7379) );
  XNOR U10147 ( .A(n7380), .B(n7379), .Z(\w1[9][33] ) );
  XOR U10148 ( .A(\w3[8][35] ), .B(\w3[8][59] ), .Z(n7410) );
  XOR U10149 ( .A(n7410), .B(key[1186]), .Z(n7382) );
  XOR U10150 ( .A(\w3[8][42] ), .B(\w3[8][50] ), .Z(n7470) );
  XNOR U10151 ( .A(\w3[8][58] ), .B(n7470), .Z(n7381) );
  XNOR U10152 ( .A(n7382), .B(n7381), .Z(\w1[9][34] ) );
  XOR U10153 ( .A(\w3[8][36] ), .B(\w3[8][32] ), .Z(n7412) );
  XOR U10154 ( .A(n7412), .B(key[1187]), .Z(n7385) );
  XOR U10155 ( .A(\w3[8][43] ), .B(\w3[8][51] ), .Z(n7438) );
  XNOR U10156 ( .A(\w3[8][56] ), .B(n7438), .Z(n7383) );
  XNOR U10157 ( .A(\w3[8][60] ), .B(n7383), .Z(n7472) );
  XNOR U10158 ( .A(\w3[8][59] ), .B(n7472), .Z(n7384) );
  XNOR U10159 ( .A(n7385), .B(n7384), .Z(\w1[9][35] ) );
  XOR U10160 ( .A(\w3[8][32] ), .B(\w3[8][37] ), .Z(n7417) );
  XOR U10161 ( .A(n7417), .B(key[1188]), .Z(n7389) );
  XOR U10162 ( .A(\w3[8][52] ), .B(\w3[8][61] ), .Z(n7387) );
  XNOR U10163 ( .A(\w3[8][56] ), .B(\w3[8][44] ), .Z(n7386) );
  XNOR U10164 ( .A(n7387), .B(n7386), .Z(n7480) );
  XNOR U10165 ( .A(\w3[8][60] ), .B(n7480), .Z(n7388) );
  XNOR U10166 ( .A(n7389), .B(n7388), .Z(\w1[9][36] ) );
  XOR U10167 ( .A(\w3[8][38] ), .B(\w3[8][62] ), .Z(n7423) );
  XOR U10168 ( .A(n7423), .B(key[1189]), .Z(n7391) );
  XOR U10169 ( .A(\w3[8][45] ), .B(\w3[8][53] ), .Z(n7486) );
  XNOR U10170 ( .A(\w3[8][61] ), .B(n7486), .Z(n7390) );
  XNOR U10171 ( .A(n7391), .B(n7390), .Z(\w1[9][37] ) );
  XOR U10172 ( .A(\w3[8][32] ), .B(\w3[8][39] ), .Z(n7424) );
  XOR U10173 ( .A(n7424), .B(key[1190]), .Z(n7393) );
  XOR U10174 ( .A(\w3[8][46] ), .B(\w3[8][54] ), .Z(n7449) );
  XNOR U10175 ( .A(\w3[8][56] ), .B(\w3[8][63] ), .Z(n7395) );
  XNOR U10176 ( .A(n7449), .B(n7395), .Z(n7488) );
  XNOR U10177 ( .A(\w3[8][62] ), .B(n7488), .Z(n7392) );
  XNOR U10178 ( .A(n7393), .B(n7392), .Z(\w1[9][38] ) );
  XOR U10179 ( .A(\w3[8][47] ), .B(\w3[8][55] ), .Z(n7491) );
  XNOR U10180 ( .A(n7491), .B(key[1191]), .Z(n7394) );
  XNOR U10181 ( .A(n7395), .B(n7394), .Z(n7396) );
  XNOR U10182 ( .A(\w3[8][32] ), .B(n7396), .Z(\w1[9][39] ) );
  XOR U10183 ( .A(n7397), .B(key[1155]), .Z(n7400) );
  XNOR U10184 ( .A(n7398), .B(\w3[8][27] ), .Z(n7399) );
  XNOR U10185 ( .A(n7400), .B(n7399), .Z(\w1[9][3] ) );
  XOR U10186 ( .A(\w3[8][32] ), .B(key[1192]), .Z(n7402) );
  XNOR U10187 ( .A(\w3[8][33] ), .B(\w3[8][41] ), .Z(n7401) );
  XNOR U10188 ( .A(n7402), .B(n7401), .Z(n7403) );
  XOR U10189 ( .A(n7492), .B(n7403), .Z(\w1[9][40] ) );
  XOR U10190 ( .A(\w3[8][42] ), .B(key[1193]), .Z(n7405) );
  XNOR U10191 ( .A(\w3[8][49] ), .B(\w3[8][34] ), .Z(n7404) );
  XNOR U10192 ( .A(n7405), .B(n7404), .Z(n7406) );
  XOR U10193 ( .A(n7431), .B(n7406), .Z(\w1[9][41] ) );
  XOR U10194 ( .A(\w3[8][43] ), .B(key[1194]), .Z(n7408) );
  XNOR U10195 ( .A(\w3[8][50] ), .B(\w3[8][35] ), .Z(n7407) );
  XNOR U10196 ( .A(n7408), .B(n7407), .Z(n7409) );
  XOR U10197 ( .A(n7439), .B(n7409), .Z(\w1[9][42] ) );
  XNOR U10198 ( .A(\w3[8][40] ), .B(n7410), .Z(n7411) );
  XNOR U10199 ( .A(\w3[8][44] ), .B(n7411), .Z(n7442) );
  XOR U10200 ( .A(n7442), .B(key[1195]), .Z(n7414) );
  XNOR U10201 ( .A(\w3[8][51] ), .B(n7412), .Z(n7413) );
  XNOR U10202 ( .A(n7414), .B(n7413), .Z(\w1[9][43] ) );
  XOR U10203 ( .A(\w3[8][36] ), .B(\w3[8][45] ), .Z(n7416) );
  XNOR U10204 ( .A(\w3[8][40] ), .B(\w3[8][60] ), .Z(n7415) );
  XNOR U10205 ( .A(n7416), .B(n7415), .Z(n7445) );
  XOR U10206 ( .A(n7445), .B(key[1196]), .Z(n7419) );
  XNOR U10207 ( .A(\w3[8][52] ), .B(n7417), .Z(n7418) );
  XNOR U10208 ( .A(n7419), .B(n7418), .Z(\w1[9][44] ) );
  XOR U10209 ( .A(\w3[8][61] ), .B(\w3[8][37] ), .Z(n7448) );
  XOR U10210 ( .A(n7448), .B(key[1197]), .Z(n7421) );
  XNOR U10211 ( .A(\w3[8][38] ), .B(\w3[8][46] ), .Z(n7420) );
  XNOR U10212 ( .A(n7421), .B(n7420), .Z(n7422) );
  XOR U10213 ( .A(\w3[8][53] ), .B(n7422), .Z(\w1[9][45] ) );
  XNOR U10214 ( .A(\w3[8][40] ), .B(\w3[8][47] ), .Z(n7457) );
  XNOR U10215 ( .A(n7423), .B(n7457), .Z(n7452) );
  XOR U10216 ( .A(n7452), .B(key[1198]), .Z(n7426) );
  XNOR U10217 ( .A(\w3[8][54] ), .B(n7424), .Z(n7425) );
  XNOR U10218 ( .A(n7426), .B(n7425), .Z(\w1[9][46] ) );
  XOR U10219 ( .A(\w3[8][63] ), .B(\w3[8][39] ), .Z(n7455) );
  XOR U10220 ( .A(n7455), .B(key[1199]), .Z(n7428) );
  XOR U10221 ( .A(\w3[8][40] ), .B(\w3[8][32] ), .Z(n7459) );
  XNOR U10222 ( .A(\w3[8][55] ), .B(n7459), .Z(n7427) );
  XNOR U10223 ( .A(n7428), .B(n7427), .Z(\w1[9][47] ) );
  XOR U10224 ( .A(n7459), .B(key[1200]), .Z(n7430) );
  XNOR U10225 ( .A(\w3[8][56] ), .B(n7466), .Z(n7429) );
  XNOR U10226 ( .A(n7430), .B(n7429), .Z(\w1[9][48] ) );
  XOR U10227 ( .A(n7470), .B(key[1201]), .Z(n7433) );
  XNOR U10228 ( .A(n7431), .B(\w3[8][41] ), .Z(n7432) );
  XNOR U10229 ( .A(n7433), .B(n7432), .Z(\w1[9][49] ) );
  XOR U10230 ( .A(n7434), .B(key[1156]), .Z(n7437) );
  XNOR U10231 ( .A(n7435), .B(\w3[8][28] ), .Z(n7436) );
  XNOR U10232 ( .A(n7437), .B(n7436), .Z(\w1[9][4] ) );
  XOR U10233 ( .A(n7438), .B(key[1202]), .Z(n7441) );
  XNOR U10234 ( .A(n7439), .B(\w3[8][42] ), .Z(n7440) );
  XNOR U10235 ( .A(n7441), .B(n7440), .Z(\w1[9][50] ) );
  XOR U10236 ( .A(\w3[8][48] ), .B(\w3[8][52] ), .Z(n7471) );
  XOR U10237 ( .A(n7471), .B(key[1203]), .Z(n7444) );
  XNOR U10238 ( .A(\w3[8][43] ), .B(n7442), .Z(n7443) );
  XNOR U10239 ( .A(n7444), .B(n7443), .Z(\w1[9][51] ) );
  XOR U10240 ( .A(\w3[8][48] ), .B(\w3[8][53] ), .Z(n7479) );
  XOR U10241 ( .A(n7479), .B(key[1204]), .Z(n7447) );
  XNOR U10242 ( .A(\w3[8][44] ), .B(n7445), .Z(n7446) );
  XNOR U10243 ( .A(n7447), .B(n7446), .Z(\w1[9][52] ) );
  XOR U10244 ( .A(n7448), .B(key[1205]), .Z(n7451) );
  XNOR U10245 ( .A(\w3[8][45] ), .B(n7449), .Z(n7450) );
  XNOR U10246 ( .A(n7451), .B(n7450), .Z(\w1[9][53] ) );
  XOR U10247 ( .A(\w3[8][48] ), .B(\w3[8][55] ), .Z(n7487) );
  XOR U10248 ( .A(n7487), .B(key[1206]), .Z(n7454) );
  XNOR U10249 ( .A(\w3[8][46] ), .B(n7452), .Z(n7453) );
  XNOR U10250 ( .A(n7454), .B(n7453), .Z(\w1[9][54] ) );
  XNOR U10251 ( .A(n7455), .B(key[1207]), .Z(n7456) );
  XNOR U10252 ( .A(n7457), .B(n7456), .Z(n7458) );
  XNOR U10253 ( .A(\w3[8][48] ), .B(n7458), .Z(\w1[9][55] ) );
  XOR U10254 ( .A(n7459), .B(key[1208]), .Z(n7461) );
  XNOR U10255 ( .A(\w3[8][48] ), .B(\w3[8][49] ), .Z(n7460) );
  XNOR U10256 ( .A(n7461), .B(n7460), .Z(n7462) );
  XOR U10257 ( .A(\w3[8][57] ), .B(n7462), .Z(\w1[9][56] ) );
  XOR U10258 ( .A(\w3[8][50] ), .B(key[1209]), .Z(n7464) );
  XNOR U10259 ( .A(\w3[8][33] ), .B(\w3[8][58] ), .Z(n7463) );
  XNOR U10260 ( .A(n7464), .B(n7463), .Z(n7465) );
  XOR U10261 ( .A(n7466), .B(n7465), .Z(\w1[9][57] ) );
  XOR U10262 ( .A(\w3[8][51] ), .B(key[1210]), .Z(n7468) );
  XNOR U10263 ( .A(\w3[8][34] ), .B(\w3[8][59] ), .Z(n7467) );
  XNOR U10264 ( .A(n7468), .B(n7467), .Z(n7469) );
  XOR U10265 ( .A(n7470), .B(n7469), .Z(\w1[9][58] ) );
  XOR U10266 ( .A(n7471), .B(key[1211]), .Z(n7474) );
  XNOR U10267 ( .A(\w3[8][35] ), .B(n7472), .Z(n7473) );
  XNOR U10268 ( .A(n7474), .B(n7473), .Z(\w1[9][59] ) );
  XOR U10269 ( .A(n7475), .B(key[1157]), .Z(n7478) );
  XNOR U10270 ( .A(\w3[8][29] ), .B(n7476), .Z(n7477) );
  XNOR U10271 ( .A(n7478), .B(n7477), .Z(\w1[9][5] ) );
  XOR U10272 ( .A(n7479), .B(key[1212]), .Z(n7482) );
  XNOR U10273 ( .A(\w3[8][36] ), .B(n7480), .Z(n7481) );
  XNOR U10274 ( .A(n7482), .B(n7481), .Z(\w1[9][60] ) );
  XOR U10275 ( .A(\w3[8][54] ), .B(key[1213]), .Z(n7484) );
  XNOR U10276 ( .A(\w3[8][37] ), .B(\w3[8][62] ), .Z(n7483) );
  XNOR U10277 ( .A(n7484), .B(n7483), .Z(n7485) );
  XOR U10278 ( .A(n7486), .B(n7485), .Z(\w1[9][61] ) );
  XOR U10279 ( .A(n7487), .B(key[1214]), .Z(n7490) );
  XNOR U10280 ( .A(\w3[8][38] ), .B(n7488), .Z(n7489) );
  XNOR U10281 ( .A(n7490), .B(n7489), .Z(\w1[9][62] ) );
  XOR U10282 ( .A(n7491), .B(key[1215]), .Z(n7494) );
  XNOR U10283 ( .A(n7492), .B(\w3[8][39] ), .Z(n7493) );
  XNOR U10284 ( .A(n7494), .B(n7493), .Z(\w1[9][63] ) );
  XOR U10285 ( .A(\w3[8][65] ), .B(\w3[8][89] ), .Z(n7553) );
  XOR U10286 ( .A(n7553), .B(key[1216]), .Z(n7496) );
  XOR U10287 ( .A(\w3[8][80] ), .B(\w3[8][88] ), .Z(n7610) );
  XNOR U10288 ( .A(n7610), .B(\w3[8][72] ), .Z(n7495) );
  XNOR U10289 ( .A(n7496), .B(n7495), .Z(\w1[9][64] ) );
  XOR U10290 ( .A(\w3[8][66] ), .B(\w3[8][90] ), .Z(n7557) );
  XOR U10291 ( .A(n7557), .B(key[1217]), .Z(n7498) );
  XOR U10292 ( .A(\w3[8][73] ), .B(\w3[8][81] ), .Z(n7584) );
  XNOR U10293 ( .A(\w3[8][89] ), .B(n7584), .Z(n7497) );
  XNOR U10294 ( .A(n7498), .B(n7497), .Z(\w1[9][65] ) );
  XOR U10295 ( .A(\w3[8][67] ), .B(\w3[8][91] ), .Z(n7528) );
  XOR U10296 ( .A(n7528), .B(key[1218]), .Z(n7500) );
  XOR U10297 ( .A(\w3[8][74] ), .B(\w3[8][82] ), .Z(n7592) );
  XNOR U10298 ( .A(\w3[8][90] ), .B(n7592), .Z(n7499) );
  XNOR U10299 ( .A(n7500), .B(n7499), .Z(\w1[9][66] ) );
  XOR U10300 ( .A(\w3[8][68] ), .B(\w3[8][64] ), .Z(n7530) );
  XOR U10301 ( .A(n7530), .B(key[1219]), .Z(n7503) );
  XOR U10302 ( .A(\w3[8][75] ), .B(\w3[8][83] ), .Z(n7556) );
  XNOR U10303 ( .A(\w3[8][88] ), .B(n7556), .Z(n7501) );
  XNOR U10304 ( .A(\w3[8][92] ), .B(n7501), .Z(n7594) );
  XNOR U10305 ( .A(\w3[8][91] ), .B(n7594), .Z(n7502) );
  XNOR U10306 ( .A(n7503), .B(n7502), .Z(\w1[9][67] ) );
  XOR U10307 ( .A(\w3[8][64] ), .B(\w3[8][69] ), .Z(n7535) );
  XOR U10308 ( .A(n7535), .B(key[1220]), .Z(n7507) );
  XOR U10309 ( .A(\w3[8][84] ), .B(\w3[8][93] ), .Z(n7505) );
  XNOR U10310 ( .A(\w3[8][88] ), .B(\w3[8][76] ), .Z(n7504) );
  XNOR U10311 ( .A(n7505), .B(n7504), .Z(n7598) );
  XNOR U10312 ( .A(\w3[8][92] ), .B(n7598), .Z(n7506) );
  XNOR U10313 ( .A(n7507), .B(n7506), .Z(\w1[9][68] ) );
  XOR U10314 ( .A(\w3[8][70] ), .B(\w3[8][94] ), .Z(n7541) );
  XOR U10315 ( .A(n7541), .B(key[1221]), .Z(n7509) );
  XOR U10316 ( .A(\w3[8][77] ), .B(\w3[8][85] ), .Z(n7604) );
  XNOR U10317 ( .A(\w3[8][93] ), .B(n7604), .Z(n7508) );
  XNOR U10318 ( .A(n7509), .B(n7508), .Z(\w1[9][69] ) );
  XOR U10319 ( .A(n7510), .B(key[1158]), .Z(n7513) );
  XNOR U10320 ( .A(n7511), .B(\w3[8][30] ), .Z(n7512) );
  XNOR U10321 ( .A(n7513), .B(n7512), .Z(\w1[9][6] ) );
  XOR U10322 ( .A(\w3[8][64] ), .B(\w3[8][71] ), .Z(n7542) );
  XOR U10323 ( .A(n7542), .B(key[1222]), .Z(n7515) );
  XOR U10324 ( .A(\w3[8][78] ), .B(\w3[8][86] ), .Z(n7567) );
  XNOR U10325 ( .A(\w3[8][88] ), .B(\w3[8][95] ), .Z(n7517) );
  XNOR U10326 ( .A(n7567), .B(n7517), .Z(n7606) );
  XNOR U10327 ( .A(\w3[8][94] ), .B(n7606), .Z(n7514) );
  XNOR U10328 ( .A(n7515), .B(n7514), .Z(\w1[9][70] ) );
  XOR U10329 ( .A(\w3[8][79] ), .B(\w3[8][87] ), .Z(n7609) );
  XNOR U10330 ( .A(n7609), .B(key[1223]), .Z(n7516) );
  XNOR U10331 ( .A(n7517), .B(n7516), .Z(n7518) );
  XNOR U10332 ( .A(\w3[8][64] ), .B(n7518), .Z(\w1[9][71] ) );
  XOR U10333 ( .A(\w3[8][64] ), .B(key[1224]), .Z(n7520) );
  XNOR U10334 ( .A(\w3[8][65] ), .B(\w3[8][73] ), .Z(n7519) );
  XNOR U10335 ( .A(n7520), .B(n7519), .Z(n7521) );
  XOR U10336 ( .A(n7610), .B(n7521), .Z(\w1[9][72] ) );
  XOR U10337 ( .A(\w3[8][74] ), .B(key[1225]), .Z(n7523) );
  XNOR U10338 ( .A(\w3[8][81] ), .B(\w3[8][66] ), .Z(n7522) );
  XNOR U10339 ( .A(n7523), .B(n7522), .Z(n7524) );
  XOR U10340 ( .A(n7553), .B(n7524), .Z(\w1[9][73] ) );
  XOR U10341 ( .A(\w3[8][75] ), .B(key[1226]), .Z(n7526) );
  XNOR U10342 ( .A(\w3[8][82] ), .B(\w3[8][67] ), .Z(n7525) );
  XNOR U10343 ( .A(n7526), .B(n7525), .Z(n7527) );
  XOR U10344 ( .A(n7557), .B(n7527), .Z(\w1[9][74] ) );
  XNOR U10345 ( .A(\w3[8][72] ), .B(n7528), .Z(n7529) );
  XNOR U10346 ( .A(\w3[8][76] ), .B(n7529), .Z(n7560) );
  XOR U10347 ( .A(n7560), .B(key[1227]), .Z(n7532) );
  XNOR U10348 ( .A(\w3[8][83] ), .B(n7530), .Z(n7531) );
  XNOR U10349 ( .A(n7532), .B(n7531), .Z(\w1[9][75] ) );
  XOR U10350 ( .A(\w3[8][68] ), .B(\w3[8][77] ), .Z(n7534) );
  XNOR U10351 ( .A(\w3[8][72] ), .B(\w3[8][92] ), .Z(n7533) );
  XNOR U10352 ( .A(n7534), .B(n7533), .Z(n7563) );
  XOR U10353 ( .A(n7563), .B(key[1228]), .Z(n7537) );
  XNOR U10354 ( .A(\w3[8][84] ), .B(n7535), .Z(n7536) );
  XNOR U10355 ( .A(n7537), .B(n7536), .Z(\w1[9][76] ) );
  XOR U10356 ( .A(\w3[8][93] ), .B(\w3[8][69] ), .Z(n7566) );
  XOR U10357 ( .A(n7566), .B(key[1229]), .Z(n7539) );
  XNOR U10358 ( .A(\w3[8][70] ), .B(\w3[8][78] ), .Z(n7538) );
  XNOR U10359 ( .A(n7539), .B(n7538), .Z(n7540) );
  XOR U10360 ( .A(\w3[8][85] ), .B(n7540), .Z(\w1[9][77] ) );
  XNOR U10361 ( .A(\w3[8][72] ), .B(\w3[8][79] ), .Z(n7575) );
  XNOR U10362 ( .A(n7541), .B(n7575), .Z(n7570) );
  XOR U10363 ( .A(n7570), .B(key[1230]), .Z(n7544) );
  XNOR U10364 ( .A(\w3[8][86] ), .B(n7542), .Z(n7543) );
  XNOR U10365 ( .A(n7544), .B(n7543), .Z(\w1[9][78] ) );
  XOR U10366 ( .A(\w3[8][95] ), .B(\w3[8][71] ), .Z(n7573) );
  XOR U10367 ( .A(n7573), .B(key[1231]), .Z(n7546) );
  XOR U10368 ( .A(\w3[8][72] ), .B(\w3[8][64] ), .Z(n7577) );
  XNOR U10369 ( .A(\w3[8][87] ), .B(n7577), .Z(n7545) );
  XNOR U10370 ( .A(n7546), .B(n7545), .Z(\w1[9][79] ) );
  XNOR U10371 ( .A(n7547), .B(key[1159]), .Z(n7548) );
  XNOR U10372 ( .A(n7549), .B(n7548), .Z(n7550) );
  XNOR U10373 ( .A(\w3[8][0] ), .B(n7550), .Z(\w1[9][7] ) );
  XOR U10374 ( .A(n7577), .B(key[1232]), .Z(n7552) );
  XNOR U10375 ( .A(\w3[8][88] ), .B(n7584), .Z(n7551) );
  XNOR U10376 ( .A(n7552), .B(n7551), .Z(\w1[9][80] ) );
  XOR U10377 ( .A(n7592), .B(key[1233]), .Z(n7555) );
  XNOR U10378 ( .A(n7553), .B(\w3[8][73] ), .Z(n7554) );
  XNOR U10379 ( .A(n7555), .B(n7554), .Z(\w1[9][81] ) );
  XOR U10380 ( .A(n7556), .B(key[1234]), .Z(n7559) );
  XNOR U10381 ( .A(n7557), .B(\w3[8][74] ), .Z(n7558) );
  XNOR U10382 ( .A(n7559), .B(n7558), .Z(\w1[9][82] ) );
  XOR U10383 ( .A(\w3[8][80] ), .B(\w3[8][84] ), .Z(n7593) );
  XOR U10384 ( .A(n7593), .B(key[1235]), .Z(n7562) );
  XNOR U10385 ( .A(\w3[8][75] ), .B(n7560), .Z(n7561) );
  XNOR U10386 ( .A(n7562), .B(n7561), .Z(\w1[9][83] ) );
  XOR U10387 ( .A(\w3[8][80] ), .B(\w3[8][85] ), .Z(n7597) );
  XOR U10388 ( .A(n7597), .B(key[1236]), .Z(n7565) );
  XNOR U10389 ( .A(\w3[8][76] ), .B(n7563), .Z(n7564) );
  XNOR U10390 ( .A(n7565), .B(n7564), .Z(\w1[9][84] ) );
  XOR U10391 ( .A(n7566), .B(key[1237]), .Z(n7569) );
  XNOR U10392 ( .A(\w3[8][77] ), .B(n7567), .Z(n7568) );
  XNOR U10393 ( .A(n7569), .B(n7568), .Z(\w1[9][85] ) );
  XOR U10394 ( .A(\w3[8][80] ), .B(\w3[8][87] ), .Z(n7605) );
  XOR U10395 ( .A(n7605), .B(key[1238]), .Z(n7572) );
  XNOR U10396 ( .A(\w3[8][78] ), .B(n7570), .Z(n7571) );
  XNOR U10397 ( .A(n7572), .B(n7571), .Z(\w1[9][86] ) );
  XNOR U10398 ( .A(n7573), .B(key[1239]), .Z(n7574) );
  XNOR U10399 ( .A(n7575), .B(n7574), .Z(n7576) );
  XNOR U10400 ( .A(\w3[8][80] ), .B(n7576), .Z(\w1[9][87] ) );
  XOR U10401 ( .A(n7577), .B(key[1240]), .Z(n7579) );
  XNOR U10402 ( .A(\w3[8][80] ), .B(\w3[8][81] ), .Z(n7578) );
  XNOR U10403 ( .A(n7579), .B(n7578), .Z(n7580) );
  XOR U10404 ( .A(\w3[8][89] ), .B(n7580), .Z(\w1[9][88] ) );
  XOR U10405 ( .A(\w3[8][82] ), .B(key[1241]), .Z(n7582) );
  XNOR U10406 ( .A(\w3[8][65] ), .B(\w3[8][90] ), .Z(n7581) );
  XNOR U10407 ( .A(n7582), .B(n7581), .Z(n7583) );
  XOR U10408 ( .A(n7584), .B(n7583), .Z(\w1[9][89] ) );
  XOR U10409 ( .A(\w3[8][9] ), .B(key[1160]), .Z(n7586) );
  XNOR U10410 ( .A(\w3[8][1] ), .B(\w3[8][0] ), .Z(n7585) );
  XNOR U10411 ( .A(n7586), .B(n7585), .Z(n7587) );
  XOR U10412 ( .A(n7588), .B(n7587), .Z(\w1[9][8] ) );
  XOR U10413 ( .A(\w3[8][83] ), .B(key[1242]), .Z(n7590) );
  XNOR U10414 ( .A(\w3[8][66] ), .B(\w3[8][91] ), .Z(n7589) );
  XNOR U10415 ( .A(n7590), .B(n7589), .Z(n7591) );
  XOR U10416 ( .A(n7592), .B(n7591), .Z(\w1[9][90] ) );
  XOR U10417 ( .A(n7593), .B(key[1243]), .Z(n7596) );
  XNOR U10418 ( .A(\w3[8][67] ), .B(n7594), .Z(n7595) );
  XNOR U10419 ( .A(n7596), .B(n7595), .Z(\w1[9][91] ) );
  XOR U10420 ( .A(n7597), .B(key[1244]), .Z(n7600) );
  XNOR U10421 ( .A(\w3[8][68] ), .B(n7598), .Z(n7599) );
  XNOR U10422 ( .A(n7600), .B(n7599), .Z(\w1[9][92] ) );
  XOR U10423 ( .A(\w3[8][86] ), .B(key[1245]), .Z(n7602) );
  XNOR U10424 ( .A(\w3[8][69] ), .B(\w3[8][94] ), .Z(n7601) );
  XNOR U10425 ( .A(n7602), .B(n7601), .Z(n7603) );
  XOR U10426 ( .A(n7604), .B(n7603), .Z(\w1[9][93] ) );
  XOR U10427 ( .A(n7605), .B(key[1246]), .Z(n7608) );
  XNOR U10428 ( .A(\w3[8][70] ), .B(n7606), .Z(n7607) );
  XNOR U10429 ( .A(n7608), .B(n7607), .Z(\w1[9][94] ) );
  XOR U10430 ( .A(n7609), .B(key[1247]), .Z(n7612) );
  XNOR U10431 ( .A(n7610), .B(\w3[8][71] ), .Z(n7611) );
  XNOR U10432 ( .A(n7612), .B(n7611), .Z(\w1[9][95] ) );
  XOR U10433 ( .A(\w3[8][104] ), .B(key[1248]), .Z(n7616) );
  XOR U10434 ( .A(n7614), .B(n7613), .Z(n7615) );
  XNOR U10435 ( .A(n7616), .B(n7615), .Z(\w1[9][96] ) );
  XOR U10436 ( .A(n7617), .B(key[1249]), .Z(n7620) );
  XNOR U10437 ( .A(\w3[8][105] ), .B(n7618), .Z(n7619) );
  XNOR U10438 ( .A(n7620), .B(n7619), .Z(\w1[9][97] ) );
  XOR U10439 ( .A(n7621), .B(key[1250]), .Z(n7624) );
  XNOR U10440 ( .A(\w3[8][106] ), .B(n7622), .Z(n7623) );
  XNOR U10441 ( .A(n7624), .B(n7623), .Z(\w1[9][98] ) );
  XOR U10442 ( .A(n7625), .B(key[1251]), .Z(n7628) );
  XNOR U10443 ( .A(n7626), .B(\w3[8][123] ), .Z(n7627) );
  XNOR U10444 ( .A(n7628), .B(n7627), .Z(\w1[9][99] ) );
  XOR U10445 ( .A(\w3[8][10] ), .B(key[1161]), .Z(n7630) );
  XNOR U10446 ( .A(\w3[8][2] ), .B(\w3[8][17] ), .Z(n7629) );
  XNOR U10447 ( .A(n7630), .B(n7629), .Z(n7631) );
  XOR U10448 ( .A(n7632), .B(n7631), .Z(\w1[9][9] ) );
endmodule

