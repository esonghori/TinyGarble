
module matrixMult_N_M_1_N3_M32 ( clk, rst, x, y, o );
  input [95:0] x;
  input [287:0] y;
  output [95:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  NAND U3 ( .A(n5150), .B(n5149), .Z(n1) );
  NAND U4 ( .A(n5147), .B(n5148), .Z(n2) );
  AND U5 ( .A(n1), .B(n2), .Z(n5201) );
  NAND U6 ( .A(n1146), .B(n1147), .Z(n3) );
  NANDN U7 ( .A(n1910), .B(n1304), .Z(n4) );
  NAND U8 ( .A(n3), .B(n4), .Z(n1221) );
  XNOR U9 ( .A(n8388), .B(n8387), .Z(n8390) );
  XNOR U10 ( .A(n5725), .B(n5724), .Z(n5693) );
  XNOR U11 ( .A(n5781), .B(n5780), .Z(n5679) );
  NAND U12 ( .A(n8575), .B(n8574), .Z(n5) );
  NANDN U13 ( .A(n8577), .B(n8576), .Z(n6) );
  AND U14 ( .A(n5), .B(n6), .Z(n9024) );
  NAND U15 ( .A(n5833), .B(n5834), .Z(n5838) );
  XNOR U16 ( .A(n5130), .B(n5129), .Z(n5131) );
  NAND U17 ( .A(n8051), .B(n8050), .Z(n7) );
  NAND U18 ( .A(n8049), .B(n8048), .Z(n8) );
  NAND U19 ( .A(n7), .B(n8), .Z(n8126) );
  NAND U20 ( .A(n7994), .B(n7993), .Z(n9) );
  NAND U21 ( .A(n7991), .B(n7992), .Z(n10) );
  AND U22 ( .A(n9), .B(n10), .Z(n8173) );
  XNOR U23 ( .A(n4304), .B(n4303), .Z(n4289) );
  NAND U24 ( .A(n1144), .B(n1145), .Z(n11) );
  NANDN U25 ( .A(n1241), .B(n1143), .Z(n12) );
  NAND U26 ( .A(n11), .B(n12), .Z(n1220) );
  XNOR U27 ( .A(n6486), .B(n6485), .Z(n6515) );
  XNOR U28 ( .A(n6920), .B(n6919), .Z(n6880) );
  XNOR U29 ( .A(n7047), .B(n7046), .Z(n7048) );
  NAND U30 ( .A(n8134), .B(n8133), .Z(n13) );
  NAND U31 ( .A(n8131), .B(n8132), .Z(n14) );
  NAND U32 ( .A(n13), .B(n14), .Z(n8383) );
  NAND U33 ( .A(n8178), .B(n8177), .Z(n15) );
  NAND U34 ( .A(n8176), .B(n8175), .Z(n16) );
  NAND U35 ( .A(n15), .B(n16), .Z(n8380) );
  XNOR U36 ( .A(n3389), .B(o[38]), .Z(n3381) );
  XNOR U37 ( .A(n3967), .B(n3966), .Z(n3958) );
  AND U38 ( .A(n4204), .B(n4203), .Z(n17) );
  AND U39 ( .A(n4548), .B(y[231]), .Z(n18) );
  NAND U40 ( .A(x[80]), .B(n18), .Z(n19) );
  NANDN U41 ( .A(n17), .B(n19), .Z(n4354) );
  NAND U42 ( .A(n5257), .B(n5256), .Z(n20) );
  NAND U43 ( .A(n5254), .B(n5255), .Z(n21) );
  NAND U44 ( .A(n20), .B(n21), .Z(n5463) );
  XNOR U45 ( .A(n1064), .B(n1063), .Z(n1055) );
  XNOR U46 ( .A(n1117), .B(n1116), .Z(n1118) );
  XNOR U47 ( .A(n1125), .B(n1124), .Z(n1089) );
  NAND U48 ( .A(n1215), .B(n1214), .Z(n22) );
  NAND U49 ( .A(n1212), .B(n1213), .Z(n23) );
  AND U50 ( .A(n22), .B(n23), .Z(n1343) );
  NAND U51 ( .A(n8334), .B(n8333), .Z(n24) );
  NAND U52 ( .A(n8332), .B(n8331), .Z(n25) );
  NAND U53 ( .A(n24), .B(n25), .Z(n8422) );
  NAND U54 ( .A(n8536), .B(n8535), .Z(n26) );
  NAND U55 ( .A(n8533), .B(n8534), .Z(n27) );
  NAND U56 ( .A(n26), .B(n27), .Z(n8663) );
  XNOR U57 ( .A(n8690), .B(n8689), .Z(n8581) );
  XOR U58 ( .A(n8585), .B(n8584), .Z(n8587) );
  XNOR U59 ( .A(n3987), .B(n3986), .Z(n3988) );
  OR U60 ( .A(n4364), .B(n4365), .Z(n28) );
  NAND U61 ( .A(n4363), .B(n4362), .Z(n29) );
  AND U62 ( .A(n28), .B(n29), .Z(n4494) );
  XNOR U63 ( .A(n5799), .B(n5798), .Z(n5689) );
  XOR U64 ( .A(n5693), .B(n5692), .Z(n5695) );
  XNOR U65 ( .A(n5826), .B(n5825), .Z(n5785) );
  NAND U66 ( .A(n5470), .B(n5469), .Z(n30) );
  NAND U67 ( .A(n5468), .B(n5467), .Z(n31) );
  NAND U68 ( .A(n30), .B(n31), .Z(n5645) );
  XNOR U69 ( .A(n832), .B(n831), .Z(n833) );
  XOR U70 ( .A(n1633), .B(n1632), .Z(n1626) );
  XNOR U71 ( .A(n8717), .B(n8716), .Z(n8676) );
  XNOR U72 ( .A(n8754), .B(n8753), .Z(n8750) );
  XNOR U73 ( .A(n3299), .B(o[35]), .Z(n3301) );
  XNOR U74 ( .A(n3456), .B(n3455), .Z(n3469) );
  XNOR U75 ( .A(n3518), .B(n3517), .Z(n3520) );
  XNOR U76 ( .A(n5842), .B(n5841), .Z(n5840) );
  NAND U77 ( .A(n5649), .B(n5648), .Z(n32) );
  NANDN U78 ( .A(n5651), .B(n5650), .Z(n33) );
  AND U79 ( .A(n32), .B(n33), .Z(n5662) );
  XNOR U80 ( .A(n382), .B(o[3]), .Z(n384) );
  NAND U81 ( .A(n2933), .B(n3112), .Z(n34) );
  XOR U82 ( .A(n2933), .B(n3112), .Z(n35) );
  NAND U83 ( .A(n35), .B(n2934), .Z(n36) );
  NAND U84 ( .A(n34), .B(n36), .Z(n2983) );
  XOR U85 ( .A(n8565), .B(n8566), .Z(n37) );
  NANDN U86 ( .A(n8567), .B(n37), .Z(n38) );
  NAND U87 ( .A(n8565), .B(n8566), .Z(n39) );
  AND U88 ( .A(n38), .B(n39), .Z(n9031) );
  NAND U89 ( .A(n3428), .B(n3429), .Z(n40) );
  XOR U90 ( .A(n3428), .B(n3429), .Z(n41) );
  NANDN U91 ( .A(n3427), .B(n41), .Z(n42) );
  NAND U92 ( .A(n40), .B(n42), .Z(n3465) );
  XNOR U93 ( .A(n5832), .B(n5831), .Z(n5829) );
  XNOR U94 ( .A(n3258), .B(n3257), .Z(n3255) );
  XNOR U95 ( .A(n1423), .B(n1422), .Z(n1404) );
  XNOR U96 ( .A(n6362), .B(o[73]), .Z(n6354) );
  XNOR U97 ( .A(n6789), .B(n6788), .Z(n6818) );
  XNOR U98 ( .A(n7165), .B(n7164), .Z(n7167) );
  XNOR U99 ( .A(n8366), .B(o[91]), .Z(n8377) );
  XOR U100 ( .A(n5245), .B(n5244), .Z(n5247) );
  XNOR U101 ( .A(n5235), .B(n5234), .Z(n5239) );
  XNOR U102 ( .A(n2369), .B(n2368), .Z(n2371) );
  XNOR U103 ( .A(n2359), .B(n2358), .Z(n2363) );
  XOR U104 ( .A(n6515), .B(n6514), .Z(n6517) );
  XOR U105 ( .A(n8394), .B(n8393), .Z(n8396) );
  NAND U106 ( .A(n8174), .B(n8173), .Z(n43) );
  NAND U107 ( .A(n8172), .B(n8171), .Z(n44) );
  NAND U108 ( .A(n43), .B(n44), .Z(n8381) );
  NAND U109 ( .A(n8317), .B(n8316), .Z(n45) );
  NAND U110 ( .A(n8315), .B(n8314), .Z(n46) );
  NAND U111 ( .A(n45), .B(n46), .Z(n8497) );
  XNOR U112 ( .A(n3688), .B(n3687), .Z(n3681) );
  XNOR U113 ( .A(n3965), .B(n3964), .Z(n3966) );
  NAND U114 ( .A(n4250), .B(n4249), .Z(n47) );
  NAND U115 ( .A(n4248), .B(n4247), .Z(n48) );
  NAND U116 ( .A(n47), .B(n48), .Z(n4363) );
  NAND U117 ( .A(n4196), .B(n4197), .Z(n49) );
  NANDN U118 ( .A(n4195), .B(n4194), .Z(n50) );
  NAND U119 ( .A(n49), .B(n50), .Z(n4287) );
  NAND U120 ( .A(n4293), .B(n4294), .Z(n51) );
  NANDN U121 ( .A(n4296), .B(n4295), .Z(n52) );
  NAND U122 ( .A(n51), .B(n52), .Z(n4388) );
  NAND U123 ( .A(n4350), .B(n4351), .Z(n53) );
  NANDN U124 ( .A(n4353), .B(n4352), .Z(n54) );
  NAND U125 ( .A(n53), .B(n54), .Z(n4484) );
  XOR U126 ( .A(n5593), .B(n5592), .Z(n5595) );
  XNOR U127 ( .A(n785), .B(n784), .Z(n778) );
  XNOR U128 ( .A(n1056), .B(n1055), .Z(n1057) );
  NAND U129 ( .A(n1098), .B(n1097), .Z(n55) );
  NAND U130 ( .A(n1095), .B(n1096), .Z(n56) );
  AND U131 ( .A(n55), .B(n56), .Z(n1254) );
  NAND U132 ( .A(n1218), .B(n1219), .Z(n57) );
  NAND U133 ( .A(n1216), .B(n1217), .Z(n58) );
  AND U134 ( .A(n57), .B(n58), .Z(n1342) );
  XNOR U135 ( .A(n6142), .B(o[67]), .Z(n6151) );
  XOR U136 ( .A(n7978), .B(n7977), .Z(n7971) );
  NAND U137 ( .A(n8386), .B(n8385), .Z(n59) );
  NAND U138 ( .A(n8384), .B(n8383), .Z(n60) );
  NAND U139 ( .A(n59), .B(n60), .Z(n8542) );
  NAND U140 ( .A(n8532), .B(n8531), .Z(n61) );
  NAND U141 ( .A(n8529), .B(n8530), .Z(n62) );
  NAND U142 ( .A(n61), .B(n62), .Z(n8664) );
  XNOR U143 ( .A(n8579), .B(n8578), .Z(n8580) );
  XNOR U144 ( .A(n8956), .B(n8955), .Z(n8953) );
  XNOR U145 ( .A(n8778), .B(n8777), .Z(n8775) );
  NAND U146 ( .A(n3340), .B(n3341), .Z(n63) );
  NAND U147 ( .A(n3568), .B(n3902), .Z(n64) );
  AND U148 ( .A(n63), .B(n64), .Z(n3371) );
  NAND U149 ( .A(n3380), .B(n3379), .Z(n65) );
  NANDN U150 ( .A(n3406), .B(n3407), .Z(n66) );
  AND U151 ( .A(n65), .B(n66), .Z(n3419) );
  XNOR U152 ( .A(n4183), .B(n4182), .Z(n4184) );
  NAND U153 ( .A(n4357), .B(n4356), .Z(n67) );
  NAND U154 ( .A(n4354), .B(n4355), .Z(n68) );
  AND U155 ( .A(n67), .B(n68), .Z(n4496) );
  XNOR U156 ( .A(n5486), .B(n5485), .Z(n5351) );
  XNOR U157 ( .A(n5689), .B(n5688), .Z(n5694) );
  XOR U158 ( .A(n5785), .B(n5784), .Z(n5787) );
  XNOR U159 ( .A(n1119), .B(n1118), .Z(n1091) );
  XNOR U160 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U161 ( .A(n1261), .B(n1260), .Z(n69) );
  NAND U162 ( .A(n1258), .B(n1259), .Z(n70) );
  NAND U163 ( .A(n69), .B(n70), .Z(n1273) );
  XNOR U164 ( .A(n2164), .B(n2163), .Z(n2304) );
  XNOR U165 ( .A(n2900), .B(n2899), .Z(n2815) );
  XOR U166 ( .A(n6965), .B(n6964), .Z(n7059) );
  XNOR U167 ( .A(n8672), .B(n8671), .Z(n8735) );
  XNOR U168 ( .A(n8978), .B(n8977), .Z(n8975) );
  XOR U169 ( .A(n3478), .B(n3477), .Z(n3519) );
  XNOR U170 ( .A(n3989), .B(n3988), .Z(n4077) );
  NAND U171 ( .A(n5518), .B(n5517), .Z(n71) );
  NANDN U172 ( .A(n5516), .B(n5515), .Z(n72) );
  AND U173 ( .A(n71), .B(n72), .Z(n5680) );
  XNOR U174 ( .A(n6072), .B(n6071), .Z(n6069) );
  XNOR U175 ( .A(n5848), .B(n5847), .Z(n5845) );
  XNOR U176 ( .A(n5836), .B(n5835), .Z(n5833) );
  NAND U177 ( .A(n5644), .B(n5645), .Z(n73) );
  NANDN U178 ( .A(n5647), .B(n5646), .Z(n74) );
  NAND U179 ( .A(n73), .B(n74), .Z(n5663) );
  XNOR U180 ( .A(n983), .B(n982), .Z(n985) );
  XOR U181 ( .A(n3246), .B(n3245), .Z(n3244) );
  XNOR U182 ( .A(n2984), .B(n2983), .Z(n2982) );
  NAND U183 ( .A(n9000), .B(n8999), .Z(n75) );
  NANDN U184 ( .A(n9002), .B(n9001), .Z(n76) );
  AND U185 ( .A(n75), .B(n76), .Z(n9010) );
  NAND U186 ( .A(n3286), .B(n3287), .Z(n77) );
  XOR U187 ( .A(n3286), .B(n3287), .Z(n78) );
  NANDN U188 ( .A(n3285), .B(n78), .Z(n79) );
  NAND U189 ( .A(n77), .B(n79), .Z(n3307) );
  NAND U190 ( .A(n3466), .B(n3467), .Z(n80) );
  XOR U191 ( .A(n3466), .B(n3467), .Z(n81) );
  NANDN U192 ( .A(n3465), .B(n81), .Z(n82) );
  NAND U193 ( .A(n80), .B(n82), .Z(n3524) );
  NAND U194 ( .A(n3983), .B(n3984), .Z(n83) );
  XOR U195 ( .A(n3983), .B(n3984), .Z(n84) );
  NANDN U196 ( .A(n3982), .B(n84), .Z(n85) );
  NAND U197 ( .A(n83), .B(n85), .Z(n4072) );
  XOR U198 ( .A(n4276), .B(n4275), .Z(n86) );
  NANDN U199 ( .A(n4277), .B(n86), .Z(n87) );
  NAND U200 ( .A(n4276), .B(n4275), .Z(n88) );
  AND U201 ( .A(n87), .B(n88), .Z(n4385) );
  NAND U202 ( .A(n4516), .B(n4517), .Z(n89) );
  XOR U203 ( .A(n4516), .B(n4517), .Z(n90) );
  NANDN U204 ( .A(n4515), .B(n90), .Z(n91) );
  NAND U205 ( .A(n89), .B(n91), .Z(n4758) );
  NAND U206 ( .A(n5654), .B(n5655), .Z(n92) );
  XOR U207 ( .A(n5654), .B(n5655), .Z(n93) );
  NANDN U208 ( .A(n5653), .B(n93), .Z(n94) );
  NAND U209 ( .A(n92), .B(n94), .Z(n6110) );
  NAND U210 ( .A(n369), .B(n370), .Z(n95) );
  XOR U211 ( .A(n369), .B(n370), .Z(n96) );
  NANDN U212 ( .A(n368), .B(n96), .Z(n97) );
  NAND U213 ( .A(n95), .B(n97), .Z(n390) );
  XOR U214 ( .A(n903), .B(n904), .Z(n98) );
  NANDN U215 ( .A(n905), .B(n98), .Z(n99) );
  NAND U216 ( .A(n903), .B(n904), .Z(n100) );
  AND U217 ( .A(n99), .B(n100), .Z(n989) );
  NAND U218 ( .A(n1614), .B(n1615), .Z(n101) );
  XOR U219 ( .A(n1614), .B(n1615), .Z(n102) );
  NANDN U220 ( .A(n1616), .B(n102), .Z(n103) );
  NAND U221 ( .A(n101), .B(n103), .Z(n1745) );
  NAND U222 ( .A(n1742), .B(n1743), .Z(n104) );
  NANDN U223 ( .A(n1741), .B(n1740), .Z(n105) );
  NAND U224 ( .A(n104), .B(n105), .Z(n1754) );
  XOR U225 ( .A(n2793), .B(n2794), .Z(n106) );
  NANDN U226 ( .A(n2795), .B(n106), .Z(n107) );
  NAND U227 ( .A(n2793), .B(n2794), .Z(n108) );
  AND U228 ( .A(n107), .B(n108), .Z(n2797) );
  XNOR U229 ( .A(n2971), .B(n2972), .Z(n2969) );
  XNOR U230 ( .A(n7244), .B(n7243), .Z(n7258) );
  XNOR U231 ( .A(n8039), .B(n8038), .Z(n8041) );
  XNOR U232 ( .A(n4096), .B(n4095), .Z(n4106) );
  XOR U233 ( .A(n5182), .B(n5181), .Z(n5184) );
  XNOR U234 ( .A(n1455), .B(n1454), .Z(n1405) );
  XNOR U235 ( .A(n1645), .B(n1644), .Z(n1662) );
  XNOR U236 ( .A(n6468), .B(n6467), .Z(n6486) );
  XNOR U237 ( .A(n7883), .B(n7882), .Z(n7884) );
  XNOR U238 ( .A(n8150), .B(n8149), .Z(n8131) );
  XNOR U239 ( .A(n8870), .B(o[94]), .Z(n8893) );
  XNOR U240 ( .A(n3862), .B(n3861), .Z(n3834) );
  NAND U241 ( .A(n4102), .B(n4103), .Z(n109) );
  NANDN U242 ( .A(n5092), .B(n4101), .Z(n110) );
  NAND U243 ( .A(n109), .B(n110), .Z(n4246) );
  XNOR U244 ( .A(n4336), .B(n4335), .Z(n4290) );
  XNOR U245 ( .A(n4963), .B(n4962), .Z(n4965) );
  XNOR U246 ( .A(n5144), .B(n5143), .Z(n5116) );
  XNOR U247 ( .A(n5239), .B(n5238), .Z(n5240) );
  NAND U248 ( .A(n5154), .B(n5153), .Z(n111) );
  NAND U249 ( .A(n5151), .B(n5152), .Z(n112) );
  AND U250 ( .A(n111), .B(n112), .Z(n5200) );
  NAND U251 ( .A(n5157), .B(n5156), .Z(n113) );
  NANDN U252 ( .A(n5159), .B(n5158), .Z(n114) );
  AND U253 ( .A(n113), .B(n114), .Z(n5256) );
  XNOR U254 ( .A(n967), .B(n966), .Z(n938) );
  XNOR U255 ( .A(n1044), .B(n1043), .Z(n1046) );
  XNOR U256 ( .A(n1131), .B(n1130), .Z(n1097) );
  XNOR U257 ( .A(n1123), .B(n1122), .Z(n1124) );
  NAND U258 ( .A(n1151), .B(n1150), .Z(n115) );
  NAND U259 ( .A(n1149), .B(n1148), .Z(n116) );
  NAND U260 ( .A(n115), .B(n116), .Z(n1219) );
  XNOR U261 ( .A(n1431), .B(n1430), .Z(n1469) );
  XNOR U262 ( .A(n2363), .B(n2362), .Z(n2365) );
  XNOR U263 ( .A(n2347), .B(n2346), .Z(n2328) );
  XNOR U264 ( .A(n6599), .B(n6598), .Z(n6601) );
  XNOR U265 ( .A(n7291), .B(n7290), .Z(n7294) );
  XOR U266 ( .A(n8496), .B(n8495), .Z(n8498) );
  NAND U267 ( .A(n8321), .B(n8320), .Z(n117) );
  NAND U268 ( .A(n8319), .B(n8318), .Z(n118) );
  NAND U269 ( .A(n117), .B(n118), .Z(n8503) );
  XOR U270 ( .A(n3444), .B(n4226), .Z(n3446) );
  XNOR U271 ( .A(n3698), .B(n3699), .Z(n3684) );
  XNOR U272 ( .A(n3959), .B(n3958), .Z(n3960) );
  XNOR U273 ( .A(n5885), .B(n5884), .Z(n5882) );
  NAND U274 ( .A(n5207), .B(n5206), .Z(n119) );
  NAND U275 ( .A(n5204), .B(n5205), .Z(n120) );
  NAND U276 ( .A(n119), .B(n120), .Z(n5467) );
  NAND U277 ( .A(n5253), .B(n5252), .Z(n121) );
  NAND U278 ( .A(n5251), .B(n5250), .Z(n122) );
  NAND U279 ( .A(n121), .B(n122), .Z(n5465) );
  XNOR U280 ( .A(n1062), .B(n1061), .Z(n1063) );
  NAND U281 ( .A(n1338), .B(n1339), .Z(n123) );
  NANDN U282 ( .A(n1341), .B(n1340), .Z(n124) );
  NAND U283 ( .A(n123), .B(n124), .Z(n1398) );
  XNOR U284 ( .A(n1538), .B(n1537), .Z(n1596) );
  XOR U285 ( .A(n2608), .B(n2607), .Z(n2610) );
  XNOR U286 ( .A(n6393), .B(n6392), .Z(n6394) );
  XNOR U287 ( .A(n6914), .B(n6913), .Z(n6882) );
  XOR U288 ( .A(n6824), .B(n6823), .Z(n6826) );
  XOR U289 ( .A(n7049), .B(n7048), .Z(n6963) );
  XNOR U290 ( .A(n7071), .B(n7070), .Z(n7173) );
  XNOR U291 ( .A(n8402), .B(n8401), .Z(n8281) );
  NAND U292 ( .A(n8338), .B(n8337), .Z(n125) );
  NANDN U293 ( .A(n8336), .B(n8335), .Z(n126) );
  AND U294 ( .A(n125), .B(n126), .Z(n8510) );
  NAND U295 ( .A(n8330), .B(n8329), .Z(n127) );
  NAND U296 ( .A(n8328), .B(n8327), .Z(n128) );
  NAND U297 ( .A(n127), .B(n128), .Z(n8423) );
  NAND U298 ( .A(n8379), .B(n8380), .Z(n129) );
  NANDN U299 ( .A(n8382), .B(n8381), .Z(n130) );
  NAND U300 ( .A(n129), .B(n130), .Z(n8541) );
  NAND U301 ( .A(n8528), .B(n8527), .Z(n131) );
  NAND U302 ( .A(n8525), .B(n8526), .Z(n132) );
  NAND U303 ( .A(n131), .B(n132), .Z(n8665) );
  XNOR U304 ( .A(n8581), .B(n8580), .Z(n8586) );
  XNOR U305 ( .A(n3392), .B(n3391), .Z(n3393) );
  XNOR U306 ( .A(n3418), .B(n3417), .Z(n3420) );
  XNOR U307 ( .A(n3454), .B(n3453), .Z(n3455) );
  XNOR U308 ( .A(n4189), .B(n4188), .Z(n4190) );
  NAND U309 ( .A(n4361), .B(n4360), .Z(n133) );
  NAND U310 ( .A(n4359), .B(n4358), .Z(n134) );
  NAND U311 ( .A(n133), .B(n134), .Z(n4493) );
  NAND U312 ( .A(n4287), .B(n4288), .Z(n135) );
  NANDN U313 ( .A(n4286), .B(n4285), .Z(n136) );
  NAND U314 ( .A(n135), .B(n136), .Z(n4491) );
  XNOR U315 ( .A(n5359), .B(n5358), .Z(n5341) );
  NAND U316 ( .A(n5424), .B(n5423), .Z(n137) );
  NANDN U317 ( .A(n5426), .B(n5425), .Z(n138) );
  AND U318 ( .A(n137), .B(n138), .Z(n5605) );
  XNOR U319 ( .A(n5687), .B(n5686), .Z(n5688) );
  XNOR U320 ( .A(n6038), .B(n6037), .Z(n6035) );
  XNOR U321 ( .A(n5504), .B(n5503), .Z(n5506) );
  XNOR U322 ( .A(n834), .B(n833), .Z(n837) );
  XOR U323 ( .A(n1177), .B(n1176), .Z(n1266) );
  XNOR U324 ( .A(n2898), .B(n2897), .Z(n2899) );
  XNOR U325 ( .A(n2948), .B(n2947), .Z(n2910) );
  XNOR U326 ( .A(n6137), .B(n6136), .Z(n6152) );
  XOR U327 ( .A(n6401), .B(n6400), .Z(n6451) );
  XNOR U328 ( .A(n6458), .B(n6457), .Z(n6459) );
  XNOR U329 ( .A(n8111), .B(n8110), .Z(n8113) );
  NAND U330 ( .A(n8421), .B(n8420), .Z(n139) );
  NANDN U331 ( .A(n8419), .B(n8418), .Z(n140) );
  AND U332 ( .A(n139), .B(n140), .Z(n8736) );
  XNOR U333 ( .A(n9002), .B(n9001), .Z(n8999) );
  XNOR U334 ( .A(n8766), .B(n8765), .Z(n8763) );
  XOR U335 ( .A(n3406), .B(n3338), .Z(n141) );
  NANDN U336 ( .A(n3339), .B(n141), .Z(n142) );
  NAND U337 ( .A(n3406), .B(n3338), .Z(n143) );
  AND U338 ( .A(n142), .B(n143), .Z(n3362) );
  NAND U339 ( .A(n3373), .B(n3372), .Z(n144) );
  NANDN U340 ( .A(n3371), .B(n3370), .Z(n145) );
  AND U341 ( .A(n144), .B(n145), .Z(n3426) );
  XNOR U342 ( .A(n3582), .B(n3581), .Z(n3584) );
  NAND U343 ( .A(n5625), .B(n5624), .Z(n146) );
  NAND U344 ( .A(n5622), .B(n5623), .Z(n147) );
  NAND U345 ( .A(n146), .B(n147), .Z(n5667) );
  XNOR U346 ( .A(n6092), .B(n6091), .Z(n6102) );
  XNOR U347 ( .A(n6060), .B(n6059), .Z(n6057) );
  XNOR U348 ( .A(n6088), .B(n6087), .Z(n6085) );
  XOR U349 ( .A(n507), .B(n421), .Z(n148) );
  NANDN U350 ( .A(n422), .B(n148), .Z(n149) );
  NAND U351 ( .A(n507), .B(n421), .Z(n150) );
  AND U352 ( .A(n149), .B(n150), .Z(n478) );
  XNOR U353 ( .A(n1086), .B(n1085), .Z(n1162) );
  XNOR U354 ( .A(n1374), .B(n1373), .Z(n1375) );
  NAND U355 ( .A(n1279), .B(n1278), .Z(n151) );
  NANDN U356 ( .A(n1277), .B(n1276), .Z(n152) );
  AND U357 ( .A(n151), .B(n152), .Z(n1495) );
  XNOR U358 ( .A(n1749), .B(n1748), .Z(n1750) );
  XOR U359 ( .A(n2479), .B(n2478), .Z(n2620) );
  XNOR U360 ( .A(n3200), .B(n3199), .Z(n3222) );
  XOR U361 ( .A(n3214), .B(n3213), .Z(n3212) );
  XOR U362 ( .A(n6382), .B(n6383), .Z(n153) );
  NANDN U363 ( .A(n6384), .B(n153), .Z(n154) );
  NAND U364 ( .A(n6382), .B(n6383), .Z(n155) );
  AND U365 ( .A(n154), .B(n155), .Z(n6444) );
  NAND U366 ( .A(n7065), .B(n7066), .Z(n156) );
  XOR U367 ( .A(n7065), .B(n7066), .Z(n157) );
  NANDN U368 ( .A(n7064), .B(n157), .Z(n158) );
  NAND U369 ( .A(n156), .B(n158), .Z(n7170) );
  XOR U370 ( .A(n7959), .B(n7960), .Z(n159) );
  NANDN U371 ( .A(n7961), .B(n159), .Z(n160) );
  NAND U372 ( .A(n7959), .B(n7960), .Z(n161) );
  AND U373 ( .A(n160), .B(n161), .Z(n8097) );
  NAND U374 ( .A(n8988), .B(n8987), .Z(n162) );
  NANDN U375 ( .A(n8990), .B(n8989), .Z(n163) );
  AND U376 ( .A(n162), .B(n163), .Z(n164) );
  NAND U377 ( .A(n8994), .B(n8993), .Z(n165) );
  NANDN U378 ( .A(n8992), .B(n8991), .Z(n166) );
  NAND U379 ( .A(n165), .B(n166), .Z(n167) );
  XNOR U380 ( .A(n164), .B(n167), .Z(n8995) );
  XOR U381 ( .A(n3324), .B(n3325), .Z(n168) );
  NANDN U382 ( .A(n3326), .B(n168), .Z(n169) );
  NAND U383 ( .A(n3324), .B(n3325), .Z(n170) );
  AND U384 ( .A(n169), .B(n170), .Z(n3354) );
  NAND U385 ( .A(n3524), .B(n3523), .Z(n171) );
  XOR U386 ( .A(n3524), .B(n3523), .Z(n172) );
  NANDN U387 ( .A(n3525), .B(n172), .Z(n173) );
  NAND U388 ( .A(n171), .B(n173), .Z(n3579) );
  XOR U389 ( .A(n4072), .B(n4073), .Z(n174) );
  NANDN U390 ( .A(n4074), .B(n174), .Z(n175) );
  NAND U391 ( .A(n4072), .B(n4073), .Z(n176) );
  AND U392 ( .A(n175), .B(n176), .Z(n4179) );
  XOR U393 ( .A(n4386), .B(n4385), .Z(n177) );
  NANDN U394 ( .A(n4384), .B(n177), .Z(n178) );
  NAND U395 ( .A(n4386), .B(n4385), .Z(n179) );
  AND U396 ( .A(n178), .B(n179), .Z(n4506) );
  XOR U397 ( .A(n4759), .B(n4758), .Z(n180) );
  NANDN U398 ( .A(n4760), .B(n180), .Z(n181) );
  NAND U399 ( .A(n4759), .B(n4758), .Z(n182) );
  AND U400 ( .A(n181), .B(n182), .Z(n4768) );
  XOR U401 ( .A(n5053), .B(n5054), .Z(n183) );
  NANDN U402 ( .A(n5055), .B(n183), .Z(n184) );
  NAND U403 ( .A(n5053), .B(n5054), .Z(n185) );
  AND U404 ( .A(n184), .B(n185), .Z(n5334) );
  NAND U405 ( .A(n5662), .B(n5663), .Z(n186) );
  NANDN U406 ( .A(n5665), .B(n5664), .Z(n187) );
  NAND U407 ( .A(n186), .B(n187), .Z(n6108) );
  NAND U408 ( .A(n390), .B(n391), .Z(n188) );
  XOR U409 ( .A(n390), .B(n391), .Z(n189) );
  NANDN U410 ( .A(n389), .B(n189), .Z(n190) );
  NAND U411 ( .A(n188), .B(n190), .Z(n407) );
  XOR U412 ( .A(n531), .B(n532), .Z(n191) );
  NANDN U413 ( .A(n533), .B(n191), .Z(n192) );
  NAND U414 ( .A(n531), .B(n532), .Z(n193) );
  AND U415 ( .A(n192), .B(n193), .Z(n621) );
  NAND U416 ( .A(n764), .B(n765), .Z(n194) );
  XOR U417 ( .A(n764), .B(n765), .Z(n195) );
  NANDN U418 ( .A(n763), .B(n195), .Z(n196) );
  NAND U419 ( .A(n194), .B(n196), .Z(n903) );
  XOR U420 ( .A(n1074), .B(n1073), .Z(n197) );
  NANDN U421 ( .A(n1075), .B(n197), .Z(n198) );
  NAND U422 ( .A(n1074), .B(n1073), .Z(n199) );
  AND U423 ( .A(n198), .B(n199), .Z(n1167) );
  NAND U424 ( .A(n1745), .B(n1746), .Z(n200) );
  XOR U425 ( .A(n1745), .B(n1746), .Z(n201) );
  NANDN U426 ( .A(n1744), .B(n201), .Z(n202) );
  NAND U427 ( .A(n200), .B(n202), .Z(n1755) );
  XOR U428 ( .A(n2300), .B(n2301), .Z(n203) );
  NANDN U429 ( .A(n2302), .B(n203), .Z(n204) );
  NAND U430 ( .A(n2300), .B(n2301), .Z(n205) );
  AND U431 ( .A(n204), .B(n205), .Z(n2464) );
  NAND U432 ( .A(n2797), .B(n2798), .Z(n206) );
  XOR U433 ( .A(n2797), .B(n2798), .Z(n207) );
  NANDN U434 ( .A(n2799), .B(n207), .Z(n208) );
  NAND U435 ( .A(n206), .B(n208), .Z(n3263) );
  XNOR U436 ( .A(n8057), .B(n8236), .Z(n7860) );
  XNOR U437 ( .A(n6976), .B(n6975), .Z(n7000) );
  XNOR U438 ( .A(n6990), .B(n6989), .Z(n6992) );
  XNOR U439 ( .A(n7229), .B(n7228), .Z(n7259) );
  XNOR U440 ( .A(n7642), .B(n7641), .Z(n7606) );
  XNOR U441 ( .A(n7706), .B(n7705), .Z(n7743) );
  XNOR U442 ( .A(n7782), .B(n7781), .Z(n7769) );
  XNOR U443 ( .A(n7895), .B(n7894), .Z(n7889) );
  XNOR U444 ( .A(n4927), .B(n4926), .Z(n4921) );
  XNOR U445 ( .A(n5132), .B(n5131), .Z(n5142) );
  XNOR U446 ( .A(n5176), .B(n5175), .Z(n5178) );
  XNOR U447 ( .A(n1241), .B(n1240), .Z(n1242) );
  XNOR U448 ( .A(n1662), .B(n1661), .Z(n1719) );
  XNOR U449 ( .A(n1910), .B(n1909), .Z(n1947) );
  XOR U450 ( .A(n2194), .B(n2193), .Z(n2200) );
  XNOR U451 ( .A(n6528), .B(n6527), .Z(n6530) );
  XOR U452 ( .A(n6550), .B(n6551), .Z(n6535) );
  XOR U453 ( .A(n6785), .B(n6784), .Z(n6819) );
  XNOR U454 ( .A(n6887), .B(n6886), .Z(n6889) );
  XNOR U455 ( .A(n7252), .B(n7251), .Z(n7199) );
  XNOR U456 ( .A(n7624), .B(n7623), .Z(n7581) );
  NAND U457 ( .A(n8065), .B(n8064), .Z(n209) );
  NAND U458 ( .A(n8062), .B(n8063), .Z(n210) );
  AND U459 ( .A(n209), .B(n210), .Z(n8133) );
  NAND U460 ( .A(n8047), .B(n8046), .Z(n211) );
  NAND U461 ( .A(n8044), .B(n8045), .Z(n212) );
  AND U462 ( .A(n211), .B(n212), .Z(n8125) );
  NAND U463 ( .A(n8056), .B(n8055), .Z(n213) );
  NAND U464 ( .A(n8053), .B(n8054), .Z(n214) );
  AND U465 ( .A(n213), .B(n214), .Z(n8177) );
  NAND U466 ( .A(n7990), .B(n7989), .Z(n215) );
  NAND U467 ( .A(n7987), .B(n7988), .Z(n216) );
  AND U468 ( .A(n215), .B(n216), .Z(n8171) );
  XNOR U469 ( .A(n8894), .B(n8893), .Z(n8891) );
  NAND U470 ( .A(n4107), .B(n4106), .Z(n217) );
  NANDN U471 ( .A(n4109), .B(n4108), .Z(n218) );
  AND U472 ( .A(n217), .B(n218), .Z(n4194) );
  XNOR U473 ( .A(n4312), .B(n4311), .Z(n4350) );
  XNOR U474 ( .A(n5284), .B(n5283), .Z(n5286) );
  NAND U475 ( .A(n5168), .B(n5167), .Z(n219) );
  NAND U476 ( .A(n5165), .B(n5166), .Z(n220) );
  AND U477 ( .A(n219), .B(n220), .Z(n5207) );
  XNOR U478 ( .A(n1155), .B(n1154), .Z(n1156) );
  XNOR U479 ( .A(n1464), .B(n1463), .Z(n1465) );
  XNOR U480 ( .A(n1502), .B(n1501), .Z(n1504) );
  XNOR U481 ( .A(n1974), .B(n1973), .Z(n1936) );
  NAND U482 ( .A(n2045), .B(n2044), .Z(n221) );
  NANDN U483 ( .A(n2047), .B(n2046), .Z(n222) );
  AND U484 ( .A(n221), .B(n222), .Z(n2206) );
  NAND U485 ( .A(n2065), .B(n2066), .Z(n223) );
  NANDN U486 ( .A(n2068), .B(n2067), .Z(n224) );
  NAND U487 ( .A(n223), .B(n224), .Z(n2215) );
  XNOR U488 ( .A(n6438), .B(n6437), .Z(n6439) );
  XNOR U489 ( .A(n6373), .B(n6372), .Z(n6374) );
  XOR U490 ( .A(n6379), .B(n6378), .Z(n6367) );
  XNOR U491 ( .A(n6918), .B(n6917), .Z(n6919) );
  XOR U492 ( .A(n6895), .B(n6894), .Z(n6911) );
  XOR U493 ( .A(n7055), .B(n7054), .Z(n6968) );
  XNOR U494 ( .A(n7075), .B(n7074), .Z(n7077) );
  XNOR U495 ( .A(n7289), .B(n7288), .Z(n7290) );
  XNOR U496 ( .A(n7976), .B(n7975), .Z(n7977) );
  NAND U497 ( .A(n8377), .B(n8378), .Z(n225) );
  NANDN U498 ( .A(n8376), .B(n8375), .Z(n226) );
  NAND U499 ( .A(n225), .B(n226), .Z(n8526) );
  XNOR U500 ( .A(n8932), .B(n8931), .Z(n8930) );
  XOR U501 ( .A(n3684), .B(n3683), .Z(n3678) );
  XNOR U502 ( .A(n3971), .B(n3970), .Z(n3973) );
  NAND U503 ( .A(n3914), .B(n4013), .Z(n227) );
  NANDN U504 ( .A(n3916), .B(n3915), .Z(n228) );
  AND U505 ( .A(n227), .B(n228), .Z(n3993) );
  NAND U506 ( .A(n4100), .B(n4099), .Z(n229) );
  NAND U507 ( .A(n4213), .B(n5093), .Z(n230) );
  NAND U508 ( .A(n229), .B(n230), .Z(n4263) );
  NAND U509 ( .A(n4246), .B(n4245), .Z(n231) );
  NAND U510 ( .A(n4243), .B(n4244), .Z(n232) );
  NAND U511 ( .A(n231), .B(n232), .Z(n4362) );
  NAND U512 ( .A(n4290), .B(n4289), .Z(n233) );
  NANDN U513 ( .A(n4292), .B(n4291), .Z(n234) );
  AND U514 ( .A(n233), .B(n234), .Z(n4389) );
  XNOR U515 ( .A(n5071), .B(n5070), .Z(n5074) );
  XNOR U516 ( .A(n5272), .B(n5271), .Z(n5274) );
  NAND U517 ( .A(n5461), .B(n5462), .Z(n235) );
  NANDN U518 ( .A(n5460), .B(n5459), .Z(n236) );
  NAND U519 ( .A(n235), .B(n236), .Z(n5626) );
  NAND U520 ( .A(n5395), .B(n5394), .Z(n237) );
  NAND U521 ( .A(n5392), .B(n5393), .Z(n238) );
  NAND U522 ( .A(n237), .B(n238), .Z(n5594) );
  XNOR U523 ( .A(n5911), .B(n5910), .Z(n5908) );
  XNOR U524 ( .A(n6006), .B(n6005), .Z(n6003) );
  NAND U525 ( .A(n5203), .B(n5202), .Z(n239) );
  NAND U526 ( .A(n5200), .B(n5201), .Z(n240) );
  NAND U527 ( .A(n239), .B(n240), .Z(n5469) );
  XNOR U528 ( .A(n605), .B(n604), .Z(n606) );
  XOR U529 ( .A(n796), .B(n795), .Z(n780) );
  XNOR U530 ( .A(n1068), .B(n1067), .Z(n1070) );
  NAND U531 ( .A(n1221), .B(n1220), .Z(n241) );
  NANDN U532 ( .A(n1223), .B(n1222), .Z(n242) );
  AND U533 ( .A(n241), .B(n242), .Z(n1344) );
  NAND U534 ( .A(n1335), .B(n1334), .Z(n243) );
  NANDN U535 ( .A(n1337), .B(n1336), .Z(n244) );
  AND U536 ( .A(n243), .B(n244), .Z(n1399) );
  XNOR U537 ( .A(n1472), .B(n1471), .Z(n1393) );
  XNOR U538 ( .A(n1407), .B(n1406), .Z(n1386) );
  XNOR U539 ( .A(n1597), .B(n1596), .Z(n1598) );
  XNOR U540 ( .A(n1631), .B(n1630), .Z(n1632) );
  XNOR U541 ( .A(n2016), .B(n2015), .Z(n2002) );
  NAND U542 ( .A(n2331), .B(n2330), .Z(n245) );
  NAND U543 ( .A(n2328), .B(n2329), .Z(n246) );
  AND U544 ( .A(n245), .B(n246), .Z(n2495) );
  NAND U545 ( .A(n2535), .B(n2534), .Z(n247) );
  NANDN U546 ( .A(n2533), .B(n2532), .Z(n248) );
  AND U547 ( .A(n247), .B(n248), .Z(n2736) );
  XNOR U548 ( .A(n6215), .B(n6214), .Z(n6217) );
  XOR U549 ( .A(n6267), .B(n6189), .Z(n249) );
  NANDN U550 ( .A(n6190), .B(n249), .Z(n250) );
  NAND U551 ( .A(n6267), .B(n6189), .Z(n251) );
  AND U552 ( .A(n250), .B(n251), .Z(n6245) );
  XNOR U553 ( .A(n6399), .B(n6398), .Z(n6400) );
  NAND U554 ( .A(n6311), .B(n7117), .Z(n252) );
  NANDN U555 ( .A(n6313), .B(n6312), .Z(n253) );
  AND U556 ( .A(n252), .B(n253), .Z(n6341) );
  XNOR U557 ( .A(n7069), .B(n7068), .Z(n7070) );
  XNOR U558 ( .A(n7422), .B(n7421), .Z(n7423) );
  XNOR U559 ( .A(n7970), .B(n7969), .Z(n7972) );
  XNOR U560 ( .A(n8281), .B(n8280), .Z(n8283) );
  NAND U561 ( .A(n8340), .B(n8339), .Z(n254) );
  NANDN U562 ( .A(n8342), .B(n8341), .Z(n255) );
  AND U563 ( .A(n254), .B(n255), .Z(n8508) );
  NAND U564 ( .A(n8307), .B(n8306), .Z(n256) );
  NAND U565 ( .A(n8304), .B(n8305), .Z(n257) );
  AND U566 ( .A(n256), .B(n257), .Z(n8520) );
  XNOR U567 ( .A(n8670), .B(n8669), .Z(n8671) );
  XOR U568 ( .A(n8694), .B(n8693), .Z(n8696) );
  XNOR U569 ( .A(n8950), .B(n8949), .Z(n8947) );
  XNOR U570 ( .A(n8786), .B(n8785), .Z(n8783) );
  XNOR U571 ( .A(n3460), .B(n3459), .Z(n3461) );
  XNOR U572 ( .A(n3961), .B(n3960), .Z(n3953) );
  XNOR U573 ( .A(n5351), .B(n5350), .Z(n5353) );
  NAND U574 ( .A(n5422), .B(n5421), .Z(n258) );
  NANDN U575 ( .A(n5420), .B(n5419), .Z(n259) );
  AND U576 ( .A(n258), .B(n259), .Z(n5607) );
  XNOR U577 ( .A(n5779), .B(n5778), .Z(n5780) );
  XNOR U578 ( .A(n5854), .B(n5853), .Z(n5851) );
  XOR U579 ( .A(n5803), .B(n5802), .Z(n5805) );
  XNOR U580 ( .A(n6032), .B(n6031), .Z(n6029) );
  XNOR U581 ( .A(n5860), .B(n5859), .Z(n5857) );
  NAND U582 ( .A(n5466), .B(n5465), .Z(n260) );
  NAND U583 ( .A(n5464), .B(n5463), .Z(n261) );
  NAND U584 ( .A(n260), .B(n261), .Z(n5644) );
  XNOR U585 ( .A(n838), .B(n837), .Z(n840) );
  XNOR U586 ( .A(n1058), .B(n1057), .Z(n1049) );
  XNOR U587 ( .A(n1090), .B(n1089), .Z(n1092) );
  XNOR U588 ( .A(n1175), .B(n1174), .Z(n1176) );
  XNOR U589 ( .A(n2471), .B(n2470), .Z(n2473) );
  XNOR U590 ( .A(n2678), .B(n2677), .Z(n2671) );
  XNOR U591 ( .A(n2924), .B(n2923), .Z(n2900) );
  XNOR U592 ( .A(n2910), .B(n2909), .Z(n2912) );
  XOR U593 ( .A(n2928), .B(n2927), .Z(n2929) );
  XOR U594 ( .A(n3010), .B(n3009), .Z(n3008) );
  XNOR U595 ( .A(n3002), .B(n3001), .Z(n2999) );
  XNOR U596 ( .A(n2996), .B(n2995), .Z(n2993) );
  XNOR U597 ( .A(n6208), .B(n6207), .Z(n6209) );
  XOR U598 ( .A(n6592), .B(n6591), .Z(n6594) );
  XNOR U599 ( .A(n6672), .B(n6671), .Z(n6674) );
  XNOR U600 ( .A(n6760), .B(n6759), .Z(n6762) );
  XNOR U601 ( .A(n6862), .B(n6861), .Z(n6863) );
  XNOR U602 ( .A(n8409), .B(n8408), .Z(n8553) );
  NAND U603 ( .A(n8540), .B(n8539), .Z(n262) );
  NAND U604 ( .A(n8537), .B(n8538), .Z(n263) );
  NAND U605 ( .A(n262), .B(n263), .Z(n8720) );
  XOR U606 ( .A(n8676), .B(n8675), .Z(n8678) );
  OR U607 ( .A(n8543), .B(n8544), .Z(n264) );
  NAND U608 ( .A(n8542), .B(n8541), .Z(n265) );
  AND U609 ( .A(n264), .B(n265), .Z(n8575) );
  XOR U610 ( .A(n9012), .B(n9011), .Z(n266) );
  XNOR U611 ( .A(n9013), .B(n266), .Z(n9000) );
  XNOR U612 ( .A(n8990), .B(n8989), .Z(n8987) );
  XNOR U613 ( .A(n8972), .B(n8971), .Z(n8970) );
  XOR U614 ( .A(n3469), .B(n3468), .Z(n3471) );
  XOR U615 ( .A(n4185), .B(n4184), .Z(n4279) );
  NAND U616 ( .A(n4492), .B(n4491), .Z(n267) );
  NAND U617 ( .A(n4489), .B(n4490), .Z(n268) );
  AND U618 ( .A(n267), .B(n268), .Z(n4510) );
  NAND U619 ( .A(n1272), .B(n1273), .Z(n269) );
  NANDN U620 ( .A(n1275), .B(n1274), .Z(n270) );
  NAND U621 ( .A(n269), .B(n270), .Z(n1496) );
  XOR U622 ( .A(n2304), .B(n2303), .Z(n2306) );
  XNOR U623 ( .A(n2632), .B(n2631), .Z(n2789) );
  XNOR U624 ( .A(n3240), .B(n3239), .Z(n3238) );
  XNOR U625 ( .A(n3225), .B(n3226), .Z(n3228) );
  XOR U626 ( .A(n2990), .B(n2989), .Z(n2988) );
  XOR U627 ( .A(n6126), .B(n6127), .Z(n271) );
  NANDN U628 ( .A(n6128), .B(n271), .Z(n272) );
  NAND U629 ( .A(n6126), .B(n6127), .Z(n273) );
  AND U630 ( .A(n272), .B(n273), .Z(n6146) );
  NAND U631 ( .A(n6331), .B(n6332), .Z(n274) );
  XOR U632 ( .A(n6331), .B(n6332), .Z(n275) );
  NANDN U633 ( .A(n6330), .B(n275), .Z(n276) );
  NAND U634 ( .A(n274), .B(n276), .Z(n6382) );
  XOR U635 ( .A(n6463), .B(n6464), .Z(n277) );
  NANDN U636 ( .A(n6465), .B(n277), .Z(n278) );
  NAND U637 ( .A(n6463), .B(n6464), .Z(n279) );
  AND U638 ( .A(n278), .B(n279), .Z(n6586) );
  XOR U639 ( .A(n7170), .B(n7171), .Z(n280) );
  NANDN U640 ( .A(n7172), .B(n280), .Z(n281) );
  NAND U641 ( .A(n7170), .B(n7171), .Z(n282) );
  AND U642 ( .A(n281), .B(n282), .Z(n7188) );
  XOR U643 ( .A(n7675), .B(n7676), .Z(n283) );
  NANDN U644 ( .A(n7677), .B(n283), .Z(n284) );
  NAND U645 ( .A(n7675), .B(n7676), .Z(n285) );
  AND U646 ( .A(n284), .B(n285), .Z(n7816) );
  XOR U647 ( .A(n8116), .B(n8117), .Z(n286) );
  NANDN U648 ( .A(n8118), .B(n286), .Z(n287) );
  NAND U649 ( .A(n8116), .B(n8117), .Z(n288) );
  AND U650 ( .A(n287), .B(n288), .Z(n8269) );
  XNOR U651 ( .A(n9032), .B(n9031), .Z(n9030) );
  NAND U652 ( .A(n3307), .B(n3308), .Z(n289) );
  XOR U653 ( .A(n3307), .B(n3308), .Z(n290) );
  NANDN U654 ( .A(n3306), .B(n290), .Z(n291) );
  NAND U655 ( .A(n289), .B(n291), .Z(n3324) );
  XOR U656 ( .A(n3367), .B(n3368), .Z(n292) );
  NANDN U657 ( .A(n3369), .B(n292), .Z(n293) );
  NAND U658 ( .A(n3367), .B(n3368), .Z(n294) );
  AND U659 ( .A(n293), .B(n294), .Z(n3428) );
  NAND U660 ( .A(n3426), .B(n3425), .Z(n295) );
  NAND U661 ( .A(n3423), .B(n3424), .Z(n296) );
  AND U662 ( .A(n295), .B(n296), .Z(n3466) );
  XOR U663 ( .A(n3579), .B(n3578), .Z(n297) );
  NANDN U664 ( .A(n3580), .B(n297), .Z(n298) );
  NAND U665 ( .A(n3579), .B(n3578), .Z(n299) );
  AND U666 ( .A(n298), .B(n299), .Z(n3644) );
  XOR U667 ( .A(n3739), .B(n3740), .Z(n300) );
  NANDN U668 ( .A(n3741), .B(n300), .Z(n301) );
  NAND U669 ( .A(n3739), .B(n3740), .Z(n302) );
  AND U670 ( .A(n301), .B(n302), .Z(n3816) );
  XOR U671 ( .A(n4180), .B(n4179), .Z(n303) );
  NANDN U672 ( .A(n4178), .B(n303), .Z(n304) );
  NAND U673 ( .A(n4180), .B(n4179), .Z(n305) );
  AND U674 ( .A(n304), .B(n305), .Z(n4276) );
  XOR U675 ( .A(n4506), .B(n4505), .Z(n306) );
  NANDN U676 ( .A(n4507), .B(n306), .Z(n307) );
  NAND U677 ( .A(n4506), .B(n4505), .Z(n308) );
  AND U678 ( .A(n307), .B(n308), .Z(n4516) );
  XOR U679 ( .A(n4768), .B(n4769), .Z(n309) );
  NANDN U680 ( .A(n4770), .B(n309), .Z(n310) );
  NAND U681 ( .A(n4768), .B(n4769), .Z(n311) );
  AND U682 ( .A(n310), .B(n311), .Z(n5040) );
  XOR U683 ( .A(n5347), .B(n5348), .Z(n312) );
  NANDN U684 ( .A(n5349), .B(n312), .Z(n313) );
  NAND U685 ( .A(n5347), .B(n5348), .Z(n314) );
  AND U686 ( .A(n313), .B(n314), .Z(n5497) );
  XOR U687 ( .A(n407), .B(n408), .Z(n315) );
  NANDN U688 ( .A(n409), .B(n315), .Z(n316) );
  NAND U689 ( .A(n407), .B(n408), .Z(n317) );
  AND U690 ( .A(n316), .B(n317), .Z(n434) );
  NAND U691 ( .A(n491), .B(n492), .Z(n318) );
  XOR U692 ( .A(n491), .B(n492), .Z(n319) );
  NANDN U693 ( .A(n490), .B(n319), .Z(n320) );
  NAND U694 ( .A(n318), .B(n320), .Z(n531) );
  XOR U695 ( .A(n634), .B(n635), .Z(n321) );
  NANDN U696 ( .A(n636), .B(n321), .Z(n322) );
  NAND U697 ( .A(n634), .B(n635), .Z(n323) );
  AND U698 ( .A(n322), .B(n323), .Z(n744) );
  XOR U699 ( .A(n990), .B(n989), .Z(n324) );
  NANDN U700 ( .A(n988), .B(n324), .Z(n325) );
  NAND U701 ( .A(n990), .B(n989), .Z(n326) );
  AND U702 ( .A(n325), .B(n326), .Z(n1074) );
  XOR U703 ( .A(n1262), .B(n1263), .Z(n327) );
  NANDN U704 ( .A(n1264), .B(n327), .Z(n328) );
  NAND U705 ( .A(n1262), .B(n1263), .Z(n329) );
  AND U706 ( .A(n328), .B(n329), .Z(n1368) );
  XOR U707 ( .A(n1754), .B(n1755), .Z(n330) );
  NANDN U708 ( .A(n1756), .B(n330), .Z(n331) );
  NAND U709 ( .A(n1754), .B(n1755), .Z(n332) );
  AND U710 ( .A(n331), .B(n332), .Z(n1884) );
  XOR U711 ( .A(n2625), .B(n2626), .Z(n333) );
  NANDN U712 ( .A(n2627), .B(n333), .Z(n334) );
  NAND U713 ( .A(n2625), .B(n2626), .Z(n335) );
  AND U714 ( .A(n334), .B(n335), .Z(n2794) );
  XNOR U715 ( .A(n3264), .B(n3263), .Z(n3262) );
  NAND U716 ( .A(n5829), .B(n5830), .Z(n336) );
  NANDN U717 ( .A(n5832), .B(n5831), .Z(n337) );
  AND U718 ( .A(n336), .B(n337), .Z(n338) );
  AND U719 ( .A(n6104), .B(n6103), .Z(n339) );
  XNOR U720 ( .A(n6098), .B(n6097), .Z(n340) );
  XNOR U721 ( .A(n339), .B(n340), .Z(n341) );
  AND U722 ( .A(n5838), .B(n5837), .Z(n342) );
  XNOR U723 ( .A(n6084), .B(n6083), .Z(n343) );
  XNOR U724 ( .A(n342), .B(n343), .Z(n344) );
  NANDN U725 ( .A(n6105), .B(n6106), .Z(n345) );
  NANDN U726 ( .A(n6107), .B(n6108), .Z(n346) );
  AND U727 ( .A(n345), .B(n346), .Z(n347) );
  NAND U728 ( .A(n6112), .B(n6111), .Z(n348) );
  NANDN U729 ( .A(n6110), .B(n6109), .Z(n349) );
  AND U730 ( .A(n348), .B(n349), .Z(n350) );
  XOR U731 ( .A(n347), .B(n350), .Z(n351) );
  XNOR U732 ( .A(n341), .B(n344), .Z(n352) );
  XNOR U733 ( .A(n351), .B(n352), .Z(n353) );
  XNOR U734 ( .A(n338), .B(n353), .Z(N128) );
  AND U735 ( .A(y[192]), .B(x[64]), .Z(n997) );
  XOR U736 ( .A(n997), .B(o[0]), .Z(N33) );
  AND U737 ( .A(x[65]), .B(y[192]), .Z(n363) );
  AND U738 ( .A(y[193]), .B(x[64]), .Z(n354) );
  XNOR U739 ( .A(n354), .B(o[1]), .Z(n357) );
  XNOR U740 ( .A(n363), .B(n357), .Z(n359) );
  NAND U741 ( .A(n997), .B(o[0]), .Z(n358) );
  XNOR U742 ( .A(n359), .B(n358), .Z(N34) );
  AND U743 ( .A(n354), .B(o[1]), .Z(n365) );
  AND U744 ( .A(x[66]), .B(y[192]), .Z(n356) );
  AND U745 ( .A(x[65]), .B(y[193]), .Z(n355) );
  XOR U746 ( .A(n356), .B(n355), .Z(n364) );
  XOR U747 ( .A(n365), .B(n364), .Z(n370) );
  NANDN U748 ( .A(n363), .B(n357), .Z(n361) );
  NAND U749 ( .A(n359), .B(n358), .Z(n360) );
  NAND U750 ( .A(n361), .B(n360), .Z(n368) );
  NAND U751 ( .A(y[194]), .B(x[64]), .Z(n373) );
  XNOR U752 ( .A(o[2]), .B(n373), .Z(n369) );
  XOR U753 ( .A(n368), .B(n369), .Z(n362) );
  XNOR U754 ( .A(n370), .B(n362), .Z(N35) );
  NAND U755 ( .A(y[193]), .B(x[66]), .Z(n382) );
  NANDN U756 ( .A(n382), .B(n363), .Z(n367) );
  NAND U757 ( .A(n365), .B(n364), .Z(n366) );
  AND U758 ( .A(n367), .B(n366), .Z(n389) );
  AND U759 ( .A(y[194]), .B(x[65]), .Z(n499) );
  XOR U760 ( .A(n499), .B(n384), .Z(n386) );
  AND U761 ( .A(x[67]), .B(y[192]), .Z(n372) );
  NAND U762 ( .A(x[64]), .B(y[195]), .Z(n371) );
  XNOR U763 ( .A(n372), .B(n371), .Z(n377) );
  ANDN U764 ( .B(o[2]), .A(n373), .Z(n376) );
  XOR U765 ( .A(n377), .B(n376), .Z(n385) );
  XOR U766 ( .A(n386), .B(n385), .Z(n391) );
  XNOR U767 ( .A(n390), .B(n391), .Z(n374) );
  XOR U768 ( .A(n389), .B(n374), .Z(N36) );
  AND U769 ( .A(y[195]), .B(x[67]), .Z(n375) );
  NAND U770 ( .A(n997), .B(n375), .Z(n379) );
  NAND U771 ( .A(n377), .B(n376), .Z(n378) );
  AND U772 ( .A(n379), .B(n378), .Z(n413) );
  AND U773 ( .A(y[196]), .B(x[64]), .Z(n381) );
  NAND U774 ( .A(y[192]), .B(x[68]), .Z(n380) );
  XNOR U775 ( .A(n381), .B(n380), .Z(n404) );
  ANDN U776 ( .B(o[3]), .A(n382), .Z(n403) );
  XOR U777 ( .A(n404), .B(n403), .Z(n411) );
  AND U778 ( .A(x[65]), .B(y[195]), .Z(n589) );
  NAND U779 ( .A(x[66]), .B(y[194]), .Z(n383) );
  XNOR U780 ( .A(n589), .B(n383), .Z(n400) );
  NAND U781 ( .A(y[193]), .B(x[67]), .Z(n395) );
  XNOR U782 ( .A(o[4]), .B(n395), .Z(n399) );
  XOR U783 ( .A(n400), .B(n399), .Z(n410) );
  XOR U784 ( .A(n411), .B(n410), .Z(n412) );
  XOR U785 ( .A(n413), .B(n412), .Z(n409) );
  NAND U786 ( .A(n499), .B(n384), .Z(n388) );
  NAND U787 ( .A(n386), .B(n385), .Z(n387) );
  NAND U788 ( .A(n388), .B(n387), .Z(n408) );
  XOR U789 ( .A(n408), .B(n407), .Z(n392) );
  XNOR U790 ( .A(n409), .B(n392), .Z(N37) );
  AND U791 ( .A(y[196]), .B(x[65]), .Z(n394) );
  NAND U792 ( .A(x[67]), .B(y[194]), .Z(n393) );
  XNOR U793 ( .A(n394), .B(n393), .Z(n418) );
  AND U794 ( .A(x[68]), .B(y[193]), .Z(n429) );
  XOR U795 ( .A(n429), .B(o[5]), .Z(n417) );
  XNOR U796 ( .A(n418), .B(n417), .Z(n421) );
  NAND U797 ( .A(y[195]), .B(x[66]), .Z(n507) );
  ANDN U798 ( .B(o[4]), .A(n395), .Z(n423) );
  AND U799 ( .A(y[197]), .B(x[64]), .Z(n397) );
  NAND U800 ( .A(y[192]), .B(x[69]), .Z(n396) );
  XOR U801 ( .A(n397), .B(n396), .Z(n424) );
  XNOR U802 ( .A(n423), .B(n424), .Z(n422) );
  XOR U803 ( .A(n507), .B(n422), .Z(n398) );
  XOR U804 ( .A(n421), .B(n398), .Z(n442) );
  NANDN U805 ( .A(n507), .B(n499), .Z(n402) );
  NAND U806 ( .A(n400), .B(n399), .Z(n401) );
  AND U807 ( .A(n402), .B(n401), .Z(n440) );
  AND U808 ( .A(x[68]), .B(y[196]), .Z(n1191) );
  NAND U809 ( .A(n1191), .B(n997), .Z(n406) );
  NAND U810 ( .A(n404), .B(n403), .Z(n405) );
  NAND U811 ( .A(n406), .B(n405), .Z(n439) );
  XNOR U812 ( .A(n440), .B(n439), .Z(n441) );
  XNOR U813 ( .A(n442), .B(n441), .Z(n436) );
  NAND U814 ( .A(n411), .B(n410), .Z(n415) );
  NANDN U815 ( .A(n413), .B(n412), .Z(n414) );
  NAND U816 ( .A(n415), .B(n414), .Z(n433) );
  IV U817 ( .A(n433), .Z(n432) );
  XOR U818 ( .A(n434), .B(n432), .Z(n416) );
  XNOR U819 ( .A(n436), .B(n416), .Z(N38) );
  AND U820 ( .A(x[67]), .B(y[196]), .Z(n508) );
  NAND U821 ( .A(n508), .B(n499), .Z(n420) );
  NAND U822 ( .A(n418), .B(n417), .Z(n419) );
  NAND U823 ( .A(n420), .B(n419), .Z(n477) );
  XOR U824 ( .A(n477), .B(n478), .Z(n480) );
  AND U825 ( .A(x[69]), .B(y[197]), .Z(n678) );
  NAND U826 ( .A(n997), .B(n678), .Z(n426) );
  NANDN U827 ( .A(n424), .B(n423), .Z(n425) );
  AND U828 ( .A(n426), .B(n425), .Z(n447) );
  AND U829 ( .A(y[198]), .B(x[64]), .Z(n428) );
  NAND U830 ( .A(x[70]), .B(y[192]), .Z(n427) );
  XNOR U831 ( .A(n428), .B(n427), .Z(n453) );
  NAND U832 ( .A(n429), .B(o[5]), .Z(n454) );
  XNOR U833 ( .A(n453), .B(n454), .Z(n446) );
  XNOR U834 ( .A(n447), .B(n446), .Z(n449) );
  AND U835 ( .A(y[196]), .B(x[66]), .Z(n960) );
  NAND U836 ( .A(x[67]), .B(y[195]), .Z(n430) );
  XNOR U837 ( .A(n960), .B(n430), .Z(n458) );
  AND U838 ( .A(y[197]), .B(x[65]), .Z(n704) );
  NAND U839 ( .A(y[194]), .B(x[68]), .Z(n431) );
  XNOR U840 ( .A(n704), .B(n431), .Z(n462) );
  NAND U841 ( .A(x[69]), .B(y[193]), .Z(n469) );
  XNOR U842 ( .A(o[6]), .B(n469), .Z(n461) );
  XOR U843 ( .A(n462), .B(n461), .Z(n457) );
  XOR U844 ( .A(n458), .B(n457), .Z(n448) );
  XOR U845 ( .A(n449), .B(n448), .Z(n479) );
  XOR U846 ( .A(n480), .B(n479), .Z(n473) );
  OR U847 ( .A(n434), .B(n432), .Z(n438) );
  ANDN U848 ( .B(n434), .A(n433), .Z(n435) );
  OR U849 ( .A(n436), .B(n435), .Z(n437) );
  AND U850 ( .A(n438), .B(n437), .Z(n471) );
  NANDN U851 ( .A(n440), .B(n439), .Z(n444) );
  NAND U852 ( .A(n442), .B(n441), .Z(n443) );
  AND U853 ( .A(n444), .B(n443), .Z(n472) );
  IV U854 ( .A(n472), .Z(n470) );
  XOR U855 ( .A(n471), .B(n470), .Z(n445) );
  XNOR U856 ( .A(n473), .B(n445), .Z(N39) );
  NANDN U857 ( .A(n447), .B(n446), .Z(n451) );
  NAND U858 ( .A(n449), .B(n448), .Z(n450) );
  AND U859 ( .A(n451), .B(n450), .Z(n487) );
  AND U860 ( .A(y[198]), .B(x[65]), .Z(n859) );
  NAND U861 ( .A(x[69]), .B(y[194]), .Z(n452) );
  XNOR U862 ( .A(n859), .B(n452), .Z(n501) );
  NAND U863 ( .A(y[193]), .B(x[70]), .Z(n505) );
  XNOR U864 ( .A(o[7]), .B(n505), .Z(n500) );
  XOR U865 ( .A(n501), .B(n500), .Z(n519) );
  AND U866 ( .A(x[70]), .B(y[198]), .Z(n718) );
  NAND U867 ( .A(n997), .B(n718), .Z(n456) );
  NANDN U868 ( .A(n454), .B(n453), .Z(n455) );
  AND U869 ( .A(n456), .B(n455), .Z(n518) );
  XNOR U870 ( .A(n519), .B(n518), .Z(n520) );
  NANDN U871 ( .A(n507), .B(n508), .Z(n460) );
  NAND U872 ( .A(n458), .B(n457), .Z(n459) );
  NAND U873 ( .A(n460), .B(n459), .Z(n521) );
  XNOR U874 ( .A(n520), .B(n521), .Z(n485) );
  AND U875 ( .A(x[68]), .B(y[197]), .Z(n1002) );
  NAND U876 ( .A(n1002), .B(n499), .Z(n464) );
  NAND U877 ( .A(n462), .B(n461), .Z(n463) );
  AND U878 ( .A(n464), .B(n463), .Z(n496) );
  AND U879 ( .A(y[197]), .B(x[66]), .Z(n466) );
  NAND U880 ( .A(y[195]), .B(x[68]), .Z(n465) );
  XNOR U881 ( .A(n466), .B(n465), .Z(n509) );
  XOR U882 ( .A(n509), .B(n508), .Z(n494) );
  AND U883 ( .A(y[199]), .B(x[64]), .Z(n468) );
  NAND U884 ( .A(x[71]), .B(y[192]), .Z(n467) );
  XNOR U885 ( .A(n468), .B(n467), .Z(n513) );
  ANDN U886 ( .B(o[6]), .A(n469), .Z(n512) );
  XNOR U887 ( .A(n513), .B(n512), .Z(n493) );
  XNOR U888 ( .A(n494), .B(n493), .Z(n495) );
  XOR U889 ( .A(n496), .B(n495), .Z(n484) );
  XOR U890 ( .A(n485), .B(n484), .Z(n486) );
  XNOR U891 ( .A(n487), .B(n486), .Z(n492) );
  NANDN U892 ( .A(n470), .B(n471), .Z(n476) );
  NOR U893 ( .A(n472), .B(n471), .Z(n474) );
  OR U894 ( .A(n474), .B(n473), .Z(n475) );
  AND U895 ( .A(n476), .B(n475), .Z(n491) );
  NAND U896 ( .A(n478), .B(n477), .Z(n482) );
  NAND U897 ( .A(n480), .B(n479), .Z(n481) );
  AND U898 ( .A(n482), .B(n481), .Z(n490) );
  XOR U899 ( .A(n491), .B(n490), .Z(n483) );
  XNOR U900 ( .A(n492), .B(n483), .Z(N40) );
  NAND U901 ( .A(n485), .B(n484), .Z(n489) );
  NAND U902 ( .A(n487), .B(n486), .Z(n488) );
  AND U903 ( .A(n489), .B(n488), .Z(n532) );
  NANDN U904 ( .A(n494), .B(n493), .Z(n498) );
  NAND U905 ( .A(n496), .B(n495), .Z(n497) );
  AND U906 ( .A(n498), .B(n497), .Z(n567) );
  AND U907 ( .A(x[69]), .B(y[198]), .Z(n670) );
  NAND U908 ( .A(n670), .B(n499), .Z(n503) );
  NAND U909 ( .A(n501), .B(n500), .Z(n502) );
  AND U910 ( .A(n503), .B(n502), .Z(n565) );
  AND U911 ( .A(y[199]), .B(x[65]), .Z(n992) );
  NAND U912 ( .A(y[195]), .B(x[69]), .Z(n504) );
  XNOR U913 ( .A(n992), .B(n504), .Z(n555) );
  ANDN U914 ( .B(o[7]), .A(n505), .Z(n554) );
  XOR U915 ( .A(n555), .B(n554), .Z(n540) );
  NAND U916 ( .A(x[67]), .B(y[197]), .Z(n1317) );
  AND U917 ( .A(y[198]), .B(x[66]), .Z(n1421) );
  NAND U918 ( .A(x[70]), .B(y[194]), .Z(n506) );
  XNOR U919 ( .A(n1421), .B(n506), .Z(n535) );
  XNOR U920 ( .A(n1191), .B(n535), .Z(n538) );
  XOR U921 ( .A(n1317), .B(n538), .Z(n539) );
  XOR U922 ( .A(n540), .B(n539), .Z(n564) );
  XNOR U923 ( .A(n565), .B(n564), .Z(n566) );
  XOR U924 ( .A(n567), .B(n566), .Z(n528) );
  NANDN U925 ( .A(n507), .B(n1002), .Z(n511) );
  NAND U926 ( .A(n509), .B(n508), .Z(n510) );
  AND U927 ( .A(n511), .B(n510), .Z(n561) );
  AND U928 ( .A(x[71]), .B(y[199]), .Z(n880) );
  NAND U929 ( .A(n997), .B(n880), .Z(n515) );
  NAND U930 ( .A(n513), .B(n512), .Z(n514) );
  AND U931 ( .A(n515), .B(n514), .Z(n559) );
  AND U932 ( .A(x[72]), .B(y[192]), .Z(n517) );
  NAND U933 ( .A(x[64]), .B(y[200]), .Z(n516) );
  XNOR U934 ( .A(n517), .B(n516), .Z(n545) );
  NAND U935 ( .A(y[193]), .B(x[71]), .Z(n550) );
  XNOR U936 ( .A(o[8]), .B(n550), .Z(n544) );
  XOR U937 ( .A(n545), .B(n544), .Z(n558) );
  XNOR U938 ( .A(n559), .B(n558), .Z(n560) );
  XOR U939 ( .A(n561), .B(n560), .Z(n526) );
  NANDN U940 ( .A(n519), .B(n518), .Z(n523) );
  NANDN U941 ( .A(n521), .B(n520), .Z(n522) );
  NAND U942 ( .A(n523), .B(n522), .Z(n525) );
  XOR U943 ( .A(n526), .B(n525), .Z(n527) );
  XNOR U944 ( .A(n528), .B(n527), .Z(n533) );
  XNOR U945 ( .A(n531), .B(n533), .Z(n524) );
  XOR U946 ( .A(n532), .B(n524), .Z(N41) );
  NAND U947 ( .A(n526), .B(n525), .Z(n530) );
  NANDN U948 ( .A(n528), .B(n527), .Z(n529) );
  NAND U949 ( .A(n530), .B(n529), .Z(n622) );
  IV U950 ( .A(n622), .Z(n620) );
  AND U951 ( .A(y[194]), .B(x[66]), .Z(n534) );
  NAND U952 ( .A(n718), .B(n534), .Z(n537) );
  NAND U953 ( .A(n1191), .B(n535), .Z(n536) );
  AND U954 ( .A(n537), .B(n536), .Z(n572) );
  NAND U955 ( .A(n1317), .B(n538), .Z(n542) );
  NANDN U956 ( .A(n540), .B(n539), .Z(n541) );
  AND U957 ( .A(n542), .B(n541), .Z(n571) );
  XNOR U958 ( .A(n572), .B(n571), .Z(n574) );
  AND U959 ( .A(y[200]), .B(x[72]), .Z(n543) );
  NAND U960 ( .A(n543), .B(n997), .Z(n547) );
  NAND U961 ( .A(n545), .B(n544), .Z(n546) );
  AND U962 ( .A(n547), .B(n546), .Z(n607) );
  AND U963 ( .A(y[196]), .B(x[69]), .Z(n549) );
  NAND U964 ( .A(x[71]), .B(y[194]), .Z(n548) );
  XNOR U965 ( .A(n549), .B(n548), .Z(n579) );
  ANDN U966 ( .B(o[8]), .A(n550), .Z(n578) );
  XOR U967 ( .A(n579), .B(n578), .Z(n605) );
  AND U968 ( .A(x[73]), .B(y[192]), .Z(n552) );
  NAND U969 ( .A(x[64]), .B(y[201]), .Z(n551) );
  XNOR U970 ( .A(n552), .B(n551), .Z(n586) );
  NAND U971 ( .A(y[193]), .B(x[72]), .Z(n596) );
  XNOR U972 ( .A(o[9]), .B(n596), .Z(n585) );
  XNOR U973 ( .A(n586), .B(n585), .Z(n604) );
  XOR U974 ( .A(n607), .B(n606), .Z(n601) );
  AND U975 ( .A(x[70]), .B(y[195]), .Z(n964) );
  NAND U976 ( .A(x[65]), .B(y[200]), .Z(n553) );
  XNOR U977 ( .A(n964), .B(n553), .Z(n591) );
  XNOR U978 ( .A(n1002), .B(n591), .Z(n610) );
  AND U979 ( .A(y[199]), .B(x[66]), .Z(n1233) );
  NAND U980 ( .A(x[67]), .B(y[198]), .Z(n917) );
  XOR U981 ( .A(n1233), .B(n917), .Z(n611) );
  XOR U982 ( .A(n610), .B(n611), .Z(n599) );
  NAND U983 ( .A(x[69]), .B(y[199]), .Z(n794) );
  NANDN U984 ( .A(n794), .B(n589), .Z(n557) );
  NAND U985 ( .A(n555), .B(n554), .Z(n556) );
  NAND U986 ( .A(n557), .B(n556), .Z(n598) );
  XOR U987 ( .A(n599), .B(n598), .Z(n600) );
  XNOR U988 ( .A(n601), .B(n600), .Z(n573) );
  XOR U989 ( .A(n574), .B(n573), .Z(n617) );
  NANDN U990 ( .A(n559), .B(n558), .Z(n563) );
  NANDN U991 ( .A(n561), .B(n560), .Z(n562) );
  AND U992 ( .A(n563), .B(n562), .Z(n615) );
  NANDN U993 ( .A(n565), .B(n564), .Z(n569) );
  NAND U994 ( .A(n567), .B(n566), .Z(n568) );
  NAND U995 ( .A(n569), .B(n568), .Z(n614) );
  XNOR U996 ( .A(n615), .B(n614), .Z(n616) );
  XOR U997 ( .A(n617), .B(n616), .Z(n623) );
  XNOR U998 ( .A(n621), .B(n623), .Z(n570) );
  XOR U999 ( .A(n620), .B(n570), .Z(N42) );
  NANDN U1000 ( .A(n572), .B(n571), .Z(n576) );
  NAND U1001 ( .A(n574), .B(n573), .Z(n575) );
  AND U1002 ( .A(n576), .B(n575), .Z(n631) );
  AND U1003 ( .A(x[71]), .B(y[196]), .Z(n672) );
  AND U1004 ( .A(y[194]), .B(x[69]), .Z(n577) );
  NAND U1005 ( .A(n672), .B(n577), .Z(n581) );
  NAND U1006 ( .A(n579), .B(n578), .Z(n580) );
  AND U1007 ( .A(n581), .B(n580), .Z(n685) );
  AND U1008 ( .A(x[71]), .B(y[195]), .Z(n583) );
  NAND U1009 ( .A(y[198]), .B(x[68]), .Z(n582) );
  XNOR U1010 ( .A(n583), .B(n582), .Z(n657) );
  AND U1011 ( .A(x[70]), .B(y[196]), .Z(n656) );
  XOR U1012 ( .A(n657), .B(n656), .Z(n683) );
  AND U1013 ( .A(y[194]), .B(x[72]), .Z(n855) );
  NAND U1014 ( .A(y[193]), .B(x[73]), .Z(n666) );
  XNOR U1015 ( .A(o[10]), .B(n666), .Z(n677) );
  XOR U1016 ( .A(n855), .B(n677), .Z(n679) );
  XNOR U1017 ( .A(n679), .B(n678), .Z(n682) );
  XNOR U1018 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U1019 ( .A(n685), .B(n684), .Z(n645) );
  AND U1020 ( .A(y[201]), .B(x[73]), .Z(n584) );
  NAND U1021 ( .A(n584), .B(n997), .Z(n588) );
  NAND U1022 ( .A(n586), .B(n585), .Z(n587) );
  NAND U1023 ( .A(n588), .B(n587), .Z(n643) );
  AND U1024 ( .A(y[200]), .B(x[70]), .Z(n590) );
  NAND U1025 ( .A(n590), .B(n589), .Z(n593) );
  NAND U1026 ( .A(n591), .B(n1002), .Z(n592) );
  AND U1027 ( .A(n593), .B(n592), .Z(n652) );
  AND U1028 ( .A(y[202]), .B(x[64]), .Z(n595) );
  NAND U1029 ( .A(x[74]), .B(y[192]), .Z(n594) );
  XNOR U1030 ( .A(n595), .B(n594), .Z(n661) );
  ANDN U1031 ( .B(o[9]), .A(n596), .Z(n660) );
  XOR U1032 ( .A(n661), .B(n660), .Z(n650) );
  AND U1033 ( .A(y[199]), .B(x[67]), .Z(n1552) );
  NAND U1034 ( .A(x[65]), .B(y[201]), .Z(n597) );
  XNOR U1035 ( .A(n1552), .B(n597), .Z(n673) );
  NAND U1036 ( .A(y[200]), .B(x[66]), .Z(n674) );
  XNOR U1037 ( .A(n673), .B(n674), .Z(n649) );
  XOR U1038 ( .A(n650), .B(n649), .Z(n651) );
  XOR U1039 ( .A(n652), .B(n651), .Z(n644) );
  XOR U1040 ( .A(n643), .B(n644), .Z(n646) );
  XOR U1041 ( .A(n645), .B(n646), .Z(n629) );
  NAND U1042 ( .A(n599), .B(n598), .Z(n603) );
  NANDN U1043 ( .A(n601), .B(n600), .Z(n602) );
  NAND U1044 ( .A(n603), .B(n602), .Z(n639) );
  NANDN U1045 ( .A(n605), .B(n604), .Z(n609) );
  NAND U1046 ( .A(n607), .B(n606), .Z(n608) );
  AND U1047 ( .A(n609), .B(n608), .Z(n638) );
  NANDN U1048 ( .A(n611), .B(n610), .Z(n613) );
  ANDN U1049 ( .B(n917), .A(n1233), .Z(n612) );
  ANDN U1050 ( .B(n613), .A(n612), .Z(n637) );
  XOR U1051 ( .A(n638), .B(n637), .Z(n640) );
  XNOR U1052 ( .A(n639), .B(n640), .Z(n628) );
  XOR U1053 ( .A(n629), .B(n628), .Z(n630) );
  XOR U1054 ( .A(n631), .B(n630), .Z(n636) );
  NANDN U1055 ( .A(n615), .B(n614), .Z(n619) );
  NAND U1056 ( .A(n617), .B(n616), .Z(n618) );
  NAND U1057 ( .A(n619), .B(n618), .Z(n635) );
  NANDN U1058 ( .A(n620), .B(n621), .Z(n626) );
  NOR U1059 ( .A(n622), .B(n621), .Z(n624) );
  OR U1060 ( .A(n624), .B(n623), .Z(n625) );
  AND U1061 ( .A(n626), .B(n625), .Z(n634) );
  XOR U1062 ( .A(n635), .B(n634), .Z(n627) );
  XNOR U1063 ( .A(n636), .B(n627), .Z(N43) );
  NAND U1064 ( .A(n629), .B(n628), .Z(n633) );
  NAND U1065 ( .A(n631), .B(n630), .Z(n632) );
  NAND U1066 ( .A(n633), .B(n632), .Z(n745) );
  IV U1067 ( .A(n745), .Z(n743) );
  NAND U1068 ( .A(n638), .B(n637), .Z(n642) );
  NAND U1069 ( .A(n640), .B(n639), .Z(n641) );
  NAND U1070 ( .A(n642), .B(n641), .Z(n752) );
  NANDN U1071 ( .A(n644), .B(n643), .Z(n648) );
  NANDN U1072 ( .A(n646), .B(n645), .Z(n647) );
  NAND U1073 ( .A(n648), .B(n647), .Z(n751) );
  NAND U1074 ( .A(n650), .B(n649), .Z(n654) );
  NANDN U1075 ( .A(n652), .B(n651), .Z(n653) );
  NAND U1076 ( .A(n654), .B(n653), .Z(n739) );
  AND U1077 ( .A(x[71]), .B(y[198]), .Z(n789) );
  AND U1078 ( .A(x[68]), .B(y[195]), .Z(n655) );
  NAND U1079 ( .A(n789), .B(n655), .Z(n659) );
  NAND U1080 ( .A(n657), .B(n656), .Z(n658) );
  NAND U1081 ( .A(n659), .B(n658), .Z(n737) );
  AND U1082 ( .A(y[202]), .B(x[74]), .Z(n1427) );
  NAND U1083 ( .A(n1427), .B(n997), .Z(n663) );
  NAND U1084 ( .A(n661), .B(n660), .Z(n662) );
  NAND U1085 ( .A(n663), .B(n662), .Z(n733) );
  AND U1086 ( .A(y[203]), .B(x[64]), .Z(n665) );
  NAND U1087 ( .A(x[75]), .B(y[192]), .Z(n664) );
  XNOR U1088 ( .A(n665), .B(n664), .Z(n710) );
  ANDN U1089 ( .B(o[10]), .A(n666), .Z(n709) );
  XOR U1090 ( .A(n710), .B(n709), .Z(n732) );
  AND U1091 ( .A(y[197]), .B(x[70]), .Z(n668) );
  NAND U1092 ( .A(y[202]), .B(x[65]), .Z(n667) );
  XNOR U1093 ( .A(n668), .B(n667), .Z(n706) );
  NAND U1094 ( .A(y[193]), .B(x[74]), .Z(n719) );
  XNOR U1095 ( .A(o[11]), .B(n719), .Z(n705) );
  XOR U1096 ( .A(n706), .B(n705), .Z(n731) );
  XOR U1097 ( .A(n732), .B(n731), .Z(n734) );
  XNOR U1098 ( .A(n733), .B(n734), .Z(n738) );
  XOR U1099 ( .A(n737), .B(n738), .Z(n740) );
  XOR U1100 ( .A(n739), .B(n740), .Z(n722) );
  NAND U1101 ( .A(y[200]), .B(x[67]), .Z(n1682) );
  NAND U1102 ( .A(x[66]), .B(y[201]), .Z(n669) );
  XNOR U1103 ( .A(n670), .B(n669), .Z(n701) );
  AND U1104 ( .A(x[68]), .B(y[199]), .Z(n700) );
  XNOR U1105 ( .A(n701), .B(n700), .Z(n726) );
  XOR U1106 ( .A(n1682), .B(n726), .Z(n728) );
  NAND U1107 ( .A(x[73]), .B(y[194]), .Z(n671) );
  XNOR U1108 ( .A(n672), .B(n671), .Z(n714) );
  AND U1109 ( .A(y[195]), .B(x[72]), .Z(n713) );
  XNOR U1110 ( .A(n714), .B(n713), .Z(n727) );
  XOR U1111 ( .A(n728), .B(n727), .Z(n692) );
  NAND U1112 ( .A(y[201]), .B(x[67]), .Z(n785) );
  NANDN U1113 ( .A(n785), .B(n992), .Z(n676) );
  NANDN U1114 ( .A(n674), .B(n673), .Z(n675) );
  AND U1115 ( .A(n676), .B(n675), .Z(n690) );
  NAND U1116 ( .A(n855), .B(n677), .Z(n681) );
  NAND U1117 ( .A(n679), .B(n678), .Z(n680) );
  NAND U1118 ( .A(n681), .B(n680), .Z(n689) );
  XNOR U1119 ( .A(n690), .B(n689), .Z(n691) );
  XOR U1120 ( .A(n692), .B(n691), .Z(n721) );
  NANDN U1121 ( .A(n683), .B(n682), .Z(n687) );
  NAND U1122 ( .A(n685), .B(n684), .Z(n686) );
  NAND U1123 ( .A(n687), .B(n686), .Z(n720) );
  XOR U1124 ( .A(n721), .B(n720), .Z(n723) );
  XNOR U1125 ( .A(n722), .B(n723), .Z(n750) );
  XOR U1126 ( .A(n751), .B(n750), .Z(n753) );
  XOR U1127 ( .A(n752), .B(n753), .Z(n746) );
  XNOR U1128 ( .A(n744), .B(n746), .Z(n688) );
  XOR U1129 ( .A(n743), .B(n688), .Z(N44) );
  NANDN U1130 ( .A(n690), .B(n689), .Z(n694) );
  NANDN U1131 ( .A(n692), .B(n691), .Z(n693) );
  NAND U1132 ( .A(n694), .B(n693), .Z(n826) );
  AND U1133 ( .A(y[195]), .B(x[73]), .Z(n1416) );
  AND U1134 ( .A(x[74]), .B(y[194]), .Z(n1458) );
  NAND U1135 ( .A(y[200]), .B(x[68]), .Z(n695) );
  XNOR U1136 ( .A(n1458), .B(n695), .Z(n817) );
  XOR U1137 ( .A(n1416), .B(n817), .Z(n796) );
  NAND U1138 ( .A(x[71]), .B(y[197]), .Z(n793) );
  XOR U1139 ( .A(n794), .B(n793), .Z(n795) );
  AND U1140 ( .A(x[76]), .B(y[192]), .Z(n697) );
  NAND U1141 ( .A(x[64]), .B(y[204]), .Z(n696) );
  XNOR U1142 ( .A(n697), .B(n696), .Z(n810) );
  NAND U1143 ( .A(y[193]), .B(x[75]), .Z(n790) );
  XNOR U1144 ( .A(o[12]), .B(n790), .Z(n809) );
  XOR U1145 ( .A(n810), .B(n809), .Z(n779) );
  AND U1146 ( .A(x[72]), .B(y[196]), .Z(n699) );
  NAND U1147 ( .A(x[66]), .B(y[202]), .Z(n698) );
  XNOR U1148 ( .A(n699), .B(n698), .Z(n784) );
  XOR U1149 ( .A(n779), .B(n778), .Z(n781) );
  XOR U1150 ( .A(n780), .B(n781), .Z(n775) );
  AND U1151 ( .A(y[201]), .B(x[69]), .Z(n1224) );
  NAND U1152 ( .A(n1421), .B(n1224), .Z(n703) );
  NAND U1153 ( .A(n701), .B(n700), .Z(n702) );
  AND U1154 ( .A(n703), .B(n702), .Z(n773) );
  AND U1155 ( .A(x[70]), .B(y[202]), .Z(n1008) );
  NAND U1156 ( .A(n1008), .B(n704), .Z(n708) );
  NAND U1157 ( .A(n706), .B(n705), .Z(n707) );
  NAND U1158 ( .A(n708), .B(n707), .Z(n772) );
  XNOR U1159 ( .A(n773), .B(n772), .Z(n774) );
  XOR U1160 ( .A(n775), .B(n774), .Z(n825) );
  AND U1161 ( .A(x[75]), .B(y[203]), .Z(n1808) );
  NAND U1162 ( .A(n1808), .B(n997), .Z(n712) );
  NAND U1163 ( .A(n710), .B(n709), .Z(n711) );
  AND U1164 ( .A(n712), .B(n711), .Z(n802) );
  AND U1165 ( .A(y[194]), .B(x[71]), .Z(n950) );
  AND U1166 ( .A(y[196]), .B(x[73]), .Z(n792) );
  NAND U1167 ( .A(n950), .B(n792), .Z(n716) );
  NAND U1168 ( .A(n714), .B(n713), .Z(n715) );
  AND U1169 ( .A(n716), .B(n715), .Z(n800) );
  NAND U1170 ( .A(y[203]), .B(x[65]), .Z(n717) );
  XNOR U1171 ( .A(n718), .B(n717), .Z(n806) );
  ANDN U1172 ( .B(o[11]), .A(n719), .Z(n805) );
  XOR U1173 ( .A(n806), .B(n805), .Z(n799) );
  XNOR U1174 ( .A(n800), .B(n799), .Z(n801) );
  XNOR U1175 ( .A(n802), .B(n801), .Z(n824) );
  XOR U1176 ( .A(n825), .B(n824), .Z(n827) );
  XNOR U1177 ( .A(n826), .B(n827), .Z(n758) );
  NAND U1178 ( .A(n721), .B(n720), .Z(n725) );
  NAND U1179 ( .A(n723), .B(n722), .Z(n724) );
  NAND U1180 ( .A(n725), .B(n724), .Z(n757) );
  XOR U1181 ( .A(n758), .B(n757), .Z(n760) );
  NAND U1182 ( .A(n1682), .B(n726), .Z(n730) );
  NAND U1183 ( .A(n728), .B(n727), .Z(n729) );
  NAND U1184 ( .A(n730), .B(n729), .Z(n766) );
  NAND U1185 ( .A(n732), .B(n731), .Z(n736) );
  NAND U1186 ( .A(n734), .B(n733), .Z(n735) );
  AND U1187 ( .A(n736), .B(n735), .Z(n767) );
  XOR U1188 ( .A(n766), .B(n767), .Z(n769) );
  NANDN U1189 ( .A(n738), .B(n737), .Z(n742) );
  NANDN U1190 ( .A(n740), .B(n739), .Z(n741) );
  AND U1191 ( .A(n742), .B(n741), .Z(n768) );
  XOR U1192 ( .A(n769), .B(n768), .Z(n759) );
  XNOR U1193 ( .A(n760), .B(n759), .Z(n765) );
  NANDN U1194 ( .A(n743), .B(n744), .Z(n749) );
  NOR U1195 ( .A(n745), .B(n744), .Z(n747) );
  OR U1196 ( .A(n747), .B(n746), .Z(n748) );
  AND U1197 ( .A(n749), .B(n748), .Z(n764) );
  NAND U1198 ( .A(n751), .B(n750), .Z(n755) );
  NAND U1199 ( .A(n753), .B(n752), .Z(n754) );
  AND U1200 ( .A(n755), .B(n754), .Z(n763) );
  XOR U1201 ( .A(n764), .B(n763), .Z(n756) );
  XNOR U1202 ( .A(n765), .B(n756), .Z(N45) );
  NAND U1203 ( .A(n758), .B(n757), .Z(n762) );
  NAND U1204 ( .A(n760), .B(n759), .Z(n761) );
  AND U1205 ( .A(n762), .B(n761), .Z(n904) );
  NAND U1206 ( .A(n767), .B(n766), .Z(n771) );
  NAND U1207 ( .A(n769), .B(n768), .Z(n770) );
  NAND U1208 ( .A(n771), .B(n770), .Z(n899) );
  NANDN U1209 ( .A(n773), .B(n772), .Z(n777) );
  NAND U1210 ( .A(n775), .B(n774), .Z(n776) );
  AND U1211 ( .A(n777), .B(n776), .Z(n838) );
  NAND U1212 ( .A(n779), .B(n778), .Z(n783) );
  NAND U1213 ( .A(n781), .B(n780), .Z(n782) );
  AND U1214 ( .A(n783), .B(n782), .Z(n834) );
  AND U1215 ( .A(x[72]), .B(y[202]), .Z(n2080) );
  NAND U1216 ( .A(n2080), .B(n960), .Z(n787) );
  NANDN U1217 ( .A(n785), .B(n784), .Z(n786) );
  AND U1218 ( .A(n787), .B(n786), .Z(n870) );
  NAND U1219 ( .A(x[65]), .B(y[204]), .Z(n788) );
  XNOR U1220 ( .A(n789), .B(n788), .Z(n861) );
  ANDN U1221 ( .B(o[12]), .A(n790), .Z(n860) );
  XOR U1222 ( .A(n861), .B(n860), .Z(n868) );
  AND U1223 ( .A(y[199]), .B(x[70]), .Z(n1846) );
  NAND U1224 ( .A(x[66]), .B(y[203]), .Z(n791) );
  XOR U1225 ( .A(n792), .B(n791), .Z(n873) );
  XNOR U1226 ( .A(n1846), .B(n873), .Z(n867) );
  XOR U1227 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1228 ( .A(n870), .B(n869), .Z(n831) );
  AND U1229 ( .A(n794), .B(n793), .Z(n798) );
  NANDN U1230 ( .A(n796), .B(n795), .Z(n797) );
  NANDN U1231 ( .A(n798), .B(n797), .Z(n832) );
  NANDN U1232 ( .A(n800), .B(n799), .Z(n804) );
  NANDN U1233 ( .A(n802), .B(n801), .Z(n803) );
  AND U1234 ( .A(n804), .B(n803), .Z(n846) );
  AND U1235 ( .A(x[70]), .B(y[203]), .Z(n1225) );
  NAND U1236 ( .A(n1225), .B(n859), .Z(n808) );
  NAND U1237 ( .A(n806), .B(n805), .Z(n807) );
  AND U1238 ( .A(n808), .B(n807), .Z(n852) );
  AND U1239 ( .A(y[204]), .B(x[76]), .Z(n2086) );
  NAND U1240 ( .A(n2086), .B(n997), .Z(n812) );
  NAND U1241 ( .A(n810), .B(n809), .Z(n811) );
  AND U1242 ( .A(n812), .B(n811), .Z(n850) );
  AND U1243 ( .A(y[195]), .B(x[74]), .Z(n1694) );
  AND U1244 ( .A(x[72]), .B(y[197]), .Z(n814) );
  NAND U1245 ( .A(x[75]), .B(y[194]), .Z(n813) );
  XOR U1246 ( .A(n814), .B(n813), .Z(n856) );
  XNOR U1247 ( .A(n1694), .B(n856), .Z(n849) );
  XNOR U1248 ( .A(n850), .B(n849), .Z(n851) );
  XNOR U1249 ( .A(n852), .B(n851), .Z(n844) );
  AND U1250 ( .A(y[200]), .B(x[74]), .Z(n816) );
  AND U1251 ( .A(x[68]), .B(y[194]), .Z(n815) );
  NAND U1252 ( .A(n816), .B(n815), .Z(n819) );
  NAND U1253 ( .A(n1416), .B(n817), .Z(n818) );
  AND U1254 ( .A(n819), .B(n818), .Z(n894) );
  AND U1255 ( .A(y[205]), .B(x[64]), .Z(n821) );
  NAND U1256 ( .A(x[77]), .B(y[192]), .Z(n820) );
  XNOR U1257 ( .A(n821), .B(n820), .Z(n886) );
  NAND U1258 ( .A(y[193]), .B(x[76]), .Z(n878) );
  XNOR U1259 ( .A(o[13]), .B(n878), .Z(n885) );
  XOR U1260 ( .A(n886), .B(n885), .Z(n892) );
  AND U1261 ( .A(y[202]), .B(x[67]), .Z(n823) );
  NAND U1262 ( .A(y[200]), .B(x[69]), .Z(n822) );
  XNOR U1263 ( .A(n823), .B(n822), .Z(n881) );
  NAND U1264 ( .A(x[68]), .B(y[201]), .Z(n882) );
  XNOR U1265 ( .A(n881), .B(n882), .Z(n891) );
  XOR U1266 ( .A(n892), .B(n891), .Z(n893) );
  XNOR U1267 ( .A(n894), .B(n893), .Z(n843) );
  XOR U1268 ( .A(n844), .B(n843), .Z(n845) );
  XNOR U1269 ( .A(n846), .B(n845), .Z(n839) );
  XOR U1270 ( .A(n840), .B(n839), .Z(n898) );
  NAND U1271 ( .A(n825), .B(n824), .Z(n829) );
  NAND U1272 ( .A(n827), .B(n826), .Z(n828) );
  AND U1273 ( .A(n829), .B(n828), .Z(n897) );
  XNOR U1274 ( .A(n898), .B(n897), .Z(n900) );
  XOR U1275 ( .A(n899), .B(n900), .Z(n905) );
  XNOR U1276 ( .A(n903), .B(n905), .Z(n830) );
  XOR U1277 ( .A(n904), .B(n830), .Z(N46) );
  NANDN U1278 ( .A(n832), .B(n831), .Z(n836) );
  NANDN U1279 ( .A(n834), .B(n833), .Z(n835) );
  AND U1280 ( .A(n836), .B(n835), .Z(n983) );
  NANDN U1281 ( .A(n838), .B(n837), .Z(n842) );
  NAND U1282 ( .A(n840), .B(n839), .Z(n841) );
  NAND U1283 ( .A(n842), .B(n841), .Z(n982) );
  NAND U1284 ( .A(n844), .B(n843), .Z(n848) );
  NANDN U1285 ( .A(n846), .B(n845), .Z(n847) );
  AND U1286 ( .A(n848), .B(n847), .Z(n910) );
  NANDN U1287 ( .A(n850), .B(n849), .Z(n854) );
  NANDN U1288 ( .A(n852), .B(n851), .Z(n853) );
  AND U1289 ( .A(n854), .B(n853), .Z(n973) );
  AND U1290 ( .A(x[75]), .B(y[197]), .Z(n1022) );
  NAND U1291 ( .A(n1022), .B(n855), .Z(n858) );
  NANDN U1292 ( .A(n856), .B(n1694), .Z(n857) );
  AND U1293 ( .A(n858), .B(n857), .Z(n933) );
  NAND U1294 ( .A(y[204]), .B(x[71]), .Z(n1431) );
  NANDN U1295 ( .A(n1431), .B(n859), .Z(n863) );
  NAND U1296 ( .A(n861), .B(n860), .Z(n862) );
  NAND U1297 ( .A(n863), .B(n862), .Z(n932) );
  XNOR U1298 ( .A(n933), .B(n932), .Z(n935) );
  AND U1299 ( .A(x[68]), .B(y[202]), .Z(n1326) );
  AND U1300 ( .A(x[72]), .B(y[198]), .Z(n865) );
  NAND U1301 ( .A(y[203]), .B(x[67]), .Z(n864) );
  XOR U1302 ( .A(n865), .B(n864), .Z(n918) );
  XNOR U1303 ( .A(n1224), .B(n918), .Z(n927) );
  XOR U1304 ( .A(n1326), .B(n927), .Z(n929) );
  AND U1305 ( .A(x[73]), .B(y[197]), .Z(n1517) );
  AND U1306 ( .A(x[74]), .B(y[196]), .Z(n1547) );
  AND U1307 ( .A(x[66]), .B(y[204]), .Z(n866) );
  XOR U1308 ( .A(n1547), .B(n866), .Z(n961) );
  XOR U1309 ( .A(n1517), .B(n961), .Z(n928) );
  XOR U1310 ( .A(n929), .B(n928), .Z(n934) );
  XOR U1311 ( .A(n935), .B(n934), .Z(n971) );
  NAND U1312 ( .A(n868), .B(n867), .Z(n872) );
  NANDN U1313 ( .A(n870), .B(n869), .Z(n871) );
  AND U1314 ( .A(n872), .B(n871), .Z(n970) );
  XNOR U1315 ( .A(n971), .B(n970), .Z(n972) );
  XOR U1316 ( .A(n973), .B(n972), .Z(n908) );
  AND U1317 ( .A(y[203]), .B(x[73]), .Z(n1429) );
  NAND U1318 ( .A(n1429), .B(n960), .Z(n875) );
  NANDN U1319 ( .A(n873), .B(n1846), .Z(n874) );
  AND U1320 ( .A(n875), .B(n874), .Z(n947) );
  AND U1321 ( .A(y[206]), .B(x[64]), .Z(n877) );
  NAND U1322 ( .A(y[192]), .B(x[78]), .Z(n876) );
  XNOR U1323 ( .A(n877), .B(n876), .Z(n914) );
  ANDN U1324 ( .B(o[13]), .A(n878), .Z(n913) );
  XOR U1325 ( .A(n914), .B(n913), .Z(n945) );
  NAND U1326 ( .A(x[76]), .B(y[194]), .Z(n879) );
  XNOR U1327 ( .A(n880), .B(n879), .Z(n951) );
  NAND U1328 ( .A(y[193]), .B(x[77]), .Z(n959) );
  XOR U1329 ( .A(o[14]), .B(n959), .Z(n952) );
  XNOR U1330 ( .A(n951), .B(n952), .Z(n944) );
  XOR U1331 ( .A(n945), .B(n944), .Z(n946) );
  XOR U1332 ( .A(n947), .B(n946), .Z(n977) );
  AND U1333 ( .A(x[69]), .B(y[202]), .Z(n1009) );
  NANDN U1334 ( .A(n1682), .B(n1009), .Z(n884) );
  NANDN U1335 ( .A(n882), .B(n881), .Z(n883) );
  AND U1336 ( .A(n884), .B(n883), .Z(n941) );
  AND U1337 ( .A(y[205]), .B(x[77]), .Z(n2426) );
  NAND U1338 ( .A(n2426), .B(n997), .Z(n888) );
  NAND U1339 ( .A(n886), .B(n885), .Z(n887) );
  AND U1340 ( .A(n888), .B(n887), .Z(n939) );
  AND U1341 ( .A(x[75]), .B(y[195]), .Z(n890) );
  NAND U1342 ( .A(x[70]), .B(y[200]), .Z(n889) );
  XNOR U1343 ( .A(n890), .B(n889), .Z(n966) );
  NAND U1344 ( .A(x[65]), .B(y[205]), .Z(n967) );
  XNOR U1345 ( .A(n939), .B(n938), .Z(n940) );
  XOR U1346 ( .A(n941), .B(n940), .Z(n976) );
  XOR U1347 ( .A(n977), .B(n976), .Z(n979) );
  NAND U1348 ( .A(n892), .B(n891), .Z(n896) );
  NANDN U1349 ( .A(n894), .B(n893), .Z(n895) );
  AND U1350 ( .A(n896), .B(n895), .Z(n978) );
  XNOR U1351 ( .A(n979), .B(n978), .Z(n907) );
  XNOR U1352 ( .A(n908), .B(n907), .Z(n909) );
  XNOR U1353 ( .A(n910), .B(n909), .Z(n984) );
  XNOR U1354 ( .A(n985), .B(n984), .Z(n990) );
  NANDN U1355 ( .A(n898), .B(n897), .Z(n902) );
  NAND U1356 ( .A(n900), .B(n899), .Z(n901) );
  AND U1357 ( .A(n902), .B(n901), .Z(n988) );
  XNOR U1358 ( .A(n988), .B(n989), .Z(n906) );
  XNOR U1359 ( .A(n990), .B(n906), .Z(N47) );
  NANDN U1360 ( .A(n908), .B(n907), .Z(n912) );
  NANDN U1361 ( .A(n910), .B(n909), .Z(n911) );
  AND U1362 ( .A(n912), .B(n911), .Z(n1079) );
  AND U1363 ( .A(x[78]), .B(y[206]), .Z(n2697) );
  NAND U1364 ( .A(n2697), .B(n997), .Z(n916) );
  NAND U1365 ( .A(n914), .B(n913), .Z(n915) );
  AND U1366 ( .A(n916), .B(n915), .Z(n1024) );
  AND U1367 ( .A(y[203]), .B(x[72]), .Z(n1301) );
  NANDN U1368 ( .A(n917), .B(n1301), .Z(n920) );
  NANDN U1369 ( .A(n918), .B(n1224), .Z(n919) );
  NAND U1370 ( .A(n920), .B(n919), .Z(n1023) );
  XNOR U1371 ( .A(n1024), .B(n1023), .Z(n1026) );
  AND U1372 ( .A(x[74]), .B(y[197]), .Z(n922) );
  NAND U1373 ( .A(y[203]), .B(x[68]), .Z(n921) );
  XNOR U1374 ( .A(n922), .B(n921), .Z(n1004) );
  AND U1375 ( .A(y[200]), .B(x[71]), .Z(n1003) );
  XOR U1376 ( .A(n1004), .B(n1003), .Z(n1011) );
  AND U1377 ( .A(y[201]), .B(x[70]), .Z(n1143) );
  XOR U1378 ( .A(n1143), .B(n1009), .Z(n1010) );
  XOR U1379 ( .A(n1011), .B(n1010), .Z(n1045) );
  AND U1380 ( .A(y[198]), .B(x[73]), .Z(n924) );
  NAND U1381 ( .A(x[66]), .B(y[205]), .Z(n923) );
  XNOR U1382 ( .A(n924), .B(n923), .Z(n1014) );
  NAND U1383 ( .A(y[204]), .B(x[67]), .Z(n1015) );
  XNOR U1384 ( .A(n1014), .B(n1015), .Z(n1043) );
  AND U1385 ( .A(x[72]), .B(y[199]), .Z(n926) );
  NAND U1386 ( .A(y[206]), .B(x[65]), .Z(n925) );
  XNOR U1387 ( .A(n926), .B(n925), .Z(n993) );
  NAND U1388 ( .A(y[193]), .B(x[78]), .Z(n1020) );
  XOR U1389 ( .A(o[15]), .B(n1020), .Z(n994) );
  XOR U1390 ( .A(n993), .B(n994), .Z(n1044) );
  XOR U1391 ( .A(n1045), .B(n1046), .Z(n1025) );
  XOR U1392 ( .A(n1026), .B(n1025), .Z(n1068) );
  NAND U1393 ( .A(n1326), .B(n927), .Z(n931) );
  NAND U1394 ( .A(n929), .B(n928), .Z(n930) );
  AND U1395 ( .A(n931), .B(n930), .Z(n1067) );
  NANDN U1396 ( .A(n933), .B(n932), .Z(n937) );
  NAND U1397 ( .A(n935), .B(n934), .Z(n936) );
  AND U1398 ( .A(n937), .B(n936), .Z(n1069) );
  XOR U1399 ( .A(n1070), .B(n1069), .Z(n1050) );
  NANDN U1400 ( .A(n939), .B(n938), .Z(n943) );
  NANDN U1401 ( .A(n941), .B(n940), .Z(n942) );
  AND U1402 ( .A(n943), .B(n942), .Z(n1058) );
  NAND U1403 ( .A(n945), .B(n944), .Z(n949) );
  NANDN U1404 ( .A(n947), .B(n946), .Z(n948) );
  AND U1405 ( .A(n949), .B(n948), .Z(n1056) );
  NAND U1406 ( .A(x[76]), .B(y[199]), .Z(n1423) );
  NANDN U1407 ( .A(n1423), .B(n950), .Z(n954) );
  NANDN U1408 ( .A(n952), .B(n951), .Z(n953) );
  AND U1409 ( .A(n954), .B(n953), .Z(n1032) );
  AND U1410 ( .A(y[196]), .B(x[75]), .Z(n956) );
  NAND U1411 ( .A(x[77]), .B(y[194]), .Z(n955) );
  XNOR U1412 ( .A(n956), .B(n955), .Z(n1036) );
  AND U1413 ( .A(y[195]), .B(x[76]), .Z(n1035) );
  XOR U1414 ( .A(n1036), .B(n1035), .Z(n1030) );
  AND U1415 ( .A(y[207]), .B(x[64]), .Z(n958) );
  NAND U1416 ( .A(x[79]), .B(y[192]), .Z(n957) );
  XNOR U1417 ( .A(n958), .B(n957), .Z(n999) );
  ANDN U1418 ( .B(o[14]), .A(n959), .Z(n998) );
  XNOR U1419 ( .A(n999), .B(n998), .Z(n1029) );
  XNOR U1420 ( .A(n1030), .B(n1029), .Z(n1031) );
  XOR U1421 ( .A(n1032), .B(n1031), .Z(n1064) );
  AND U1422 ( .A(y[204]), .B(x[74]), .Z(n1681) );
  IV U1423 ( .A(n1681), .Z(n1848) );
  NANDN U1424 ( .A(n1848), .B(n960), .Z(n963) );
  NAND U1425 ( .A(n1517), .B(n961), .Z(n962) );
  AND U1426 ( .A(n963), .B(n962), .Z(n1062) );
  AND U1427 ( .A(y[200]), .B(x[75]), .Z(n965) );
  NAND U1428 ( .A(n965), .B(n964), .Z(n969) );
  NANDN U1429 ( .A(n967), .B(n966), .Z(n968) );
  NAND U1430 ( .A(n969), .B(n968), .Z(n1061) );
  XNOR U1431 ( .A(n1050), .B(n1049), .Z(n1051) );
  NANDN U1432 ( .A(n971), .B(n970), .Z(n975) );
  NAND U1433 ( .A(n973), .B(n972), .Z(n974) );
  NAND U1434 ( .A(n975), .B(n974), .Z(n1052) );
  XNOR U1435 ( .A(n1051), .B(n1052), .Z(n1076) );
  NAND U1436 ( .A(n977), .B(n976), .Z(n981) );
  NAND U1437 ( .A(n979), .B(n978), .Z(n980) );
  NAND U1438 ( .A(n981), .B(n980), .Z(n1077) );
  XNOR U1439 ( .A(n1076), .B(n1077), .Z(n1078) );
  XOR U1440 ( .A(n1079), .B(n1078), .Z(n1075) );
  NANDN U1441 ( .A(n983), .B(n982), .Z(n987) );
  NAND U1442 ( .A(n985), .B(n984), .Z(n986) );
  NAND U1443 ( .A(n987), .B(n986), .Z(n1073) );
  XOR U1444 ( .A(n1073), .B(n1074), .Z(n991) );
  XNOR U1445 ( .A(n1075), .B(n991), .Z(N48) );
  AND U1446 ( .A(y[206]), .B(x[72]), .Z(n1703) );
  NAND U1447 ( .A(n1703), .B(n992), .Z(n996) );
  NANDN U1448 ( .A(n994), .B(n993), .Z(n995) );
  NAND U1449 ( .A(n996), .B(n995), .Z(n1095) );
  AND U1450 ( .A(y[207]), .B(x[79]), .Z(n3020) );
  NAND U1451 ( .A(n3020), .B(n997), .Z(n1001) );
  NAND U1452 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1453 ( .A(n1001), .B(n1000), .Z(n1096) );
  XOR U1454 ( .A(n1095), .B(n1096), .Z(n1098) );
  AND U1455 ( .A(y[203]), .B(x[74]), .Z(n1560) );
  NAND U1456 ( .A(n1560), .B(n1002), .Z(n1006) );
  NAND U1457 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1458 ( .A(n1006), .B(n1005), .Z(n1131) );
  AND U1459 ( .A(x[64]), .B(y[208]), .Z(n1149) );
  AND U1460 ( .A(x[80]), .B(y[192]), .Z(n1148) );
  XOR U1461 ( .A(n1149), .B(n1148), .Z(n1151) );
  AND U1462 ( .A(y[193]), .B(x[79]), .Z(n1140) );
  XOR U1463 ( .A(n1140), .B(o[16]), .Z(n1150) );
  XOR U1464 ( .A(n1151), .B(n1150), .Z(n1129) );
  NAND U1465 ( .A(x[71]), .B(y[201]), .Z(n1007) );
  XNOR U1466 ( .A(n1008), .B(n1007), .Z(n1145) );
  AND U1467 ( .A(y[198]), .B(x[74]), .Z(n1144) );
  XOR U1468 ( .A(n1145), .B(n1144), .Z(n1128) );
  XOR U1469 ( .A(n1129), .B(n1128), .Z(n1130) );
  XOR U1470 ( .A(n1098), .B(n1097), .Z(n1125) );
  OR U1471 ( .A(n1009), .B(n1143), .Z(n1013) );
  NANDN U1472 ( .A(n1011), .B(n1010), .Z(n1012) );
  AND U1473 ( .A(n1013), .B(n1012), .Z(n1123) );
  AND U1474 ( .A(y[205]), .B(x[73]), .Z(n1829) );
  NAND U1475 ( .A(n1829), .B(n1421), .Z(n1017) );
  NANDN U1476 ( .A(n1015), .B(n1014), .Z(n1016) );
  AND U1477 ( .A(n1017), .B(n1016), .Z(n1157) );
  AND U1478 ( .A(y[207]), .B(x[65]), .Z(n1019) );
  NAND U1479 ( .A(x[72]), .B(y[200]), .Z(n1018) );
  XNOR U1480 ( .A(n1019), .B(n1018), .Z(n1147) );
  ANDN U1481 ( .B(o[15]), .A(n1020), .Z(n1146) );
  XOR U1482 ( .A(n1147), .B(n1146), .Z(n1154) );
  NAND U1483 ( .A(x[78]), .B(y[194]), .Z(n1021) );
  XNOR U1484 ( .A(n1022), .B(n1021), .Z(n1105) );
  NAND U1485 ( .A(x[68]), .B(y[204]), .Z(n1106) );
  XOR U1486 ( .A(n1105), .B(n1106), .Z(n1155) );
  XOR U1487 ( .A(n1157), .B(n1156), .Z(n1122) );
  NANDN U1488 ( .A(n1024), .B(n1023), .Z(n1028) );
  NAND U1489 ( .A(n1026), .B(n1025), .Z(n1027) );
  NAND U1490 ( .A(n1028), .B(n1027), .Z(n1090) );
  NANDN U1491 ( .A(n1030), .B(n1029), .Z(n1034) );
  NAND U1492 ( .A(n1032), .B(n1031), .Z(n1033) );
  AND U1493 ( .A(n1034), .B(n1033), .Z(n1119) );
  AND U1494 ( .A(y[194]), .B(x[75]), .Z(n1654) );
  AND U1495 ( .A(y[196]), .B(x[77]), .Z(n1115) );
  NAND U1496 ( .A(n1654), .B(n1115), .Z(n1038) );
  NAND U1497 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1498 ( .A(n1038), .B(n1037), .Z(n1101) );
  AND U1499 ( .A(x[73]), .B(y[199]), .Z(n1040) );
  NAND U1500 ( .A(x[66]), .B(y[206]), .Z(n1039) );
  XNOR U1501 ( .A(n1040), .B(n1039), .Z(n1109) );
  NAND U1502 ( .A(y[205]), .B(x[67]), .Z(n1110) );
  XNOR U1503 ( .A(n1109), .B(n1110), .Z(n1099) );
  AND U1504 ( .A(x[76]), .B(y[196]), .Z(n1818) );
  AND U1505 ( .A(x[77]), .B(y[195]), .Z(n1042) );
  NAND U1506 ( .A(y[203]), .B(x[69]), .Z(n1041) );
  XOR U1507 ( .A(n1042), .B(n1041), .Z(n1135) );
  XOR U1508 ( .A(n1818), .B(n1135), .Z(n1100) );
  XOR U1509 ( .A(n1099), .B(n1100), .Z(n1102) );
  XOR U1510 ( .A(n1101), .B(n1102), .Z(n1117) );
  NANDN U1511 ( .A(n1044), .B(n1043), .Z(n1048) );
  NAND U1512 ( .A(n1046), .B(n1045), .Z(n1047) );
  AND U1513 ( .A(n1048), .B(n1047), .Z(n1116) );
  XOR U1514 ( .A(n1092), .B(n1091), .Z(n1161) );
  NANDN U1515 ( .A(n1050), .B(n1049), .Z(n1054) );
  NANDN U1516 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1517 ( .A(n1054), .B(n1053), .Z(n1160) );
  XNOR U1518 ( .A(n1161), .B(n1160), .Z(n1163) );
  NANDN U1519 ( .A(n1056), .B(n1055), .Z(n1060) );
  NANDN U1520 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U1521 ( .A(n1060), .B(n1059), .Z(n1086) );
  NANDN U1522 ( .A(n1062), .B(n1061), .Z(n1066) );
  NANDN U1523 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1524 ( .A(n1066), .B(n1065), .Z(n1084) );
  NANDN U1525 ( .A(n1068), .B(n1067), .Z(n1072) );
  NAND U1526 ( .A(n1070), .B(n1069), .Z(n1071) );
  AND U1527 ( .A(n1072), .B(n1071), .Z(n1083) );
  XOR U1528 ( .A(n1163), .B(n1162), .Z(n1169) );
  NANDN U1529 ( .A(n1077), .B(n1076), .Z(n1081) );
  NANDN U1530 ( .A(n1079), .B(n1078), .Z(n1080) );
  AND U1531 ( .A(n1081), .B(n1080), .Z(n1168) );
  IV U1532 ( .A(n1168), .Z(n1166) );
  XOR U1533 ( .A(n1167), .B(n1166), .Z(n1082) );
  XNOR U1534 ( .A(n1169), .B(n1082), .Z(N49) );
  NANDN U1535 ( .A(n1084), .B(n1083), .Z(n1088) );
  NANDN U1536 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U1537 ( .A(n1088), .B(n1087), .Z(n1268) );
  NANDN U1538 ( .A(n1090), .B(n1089), .Z(n1094) );
  NAND U1539 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U1540 ( .A(n1094), .B(n1093), .Z(n1177) );
  NANDN U1541 ( .A(n1100), .B(n1099), .Z(n1104) );
  OR U1542 ( .A(n1102), .B(n1101), .Z(n1103) );
  AND U1543 ( .A(n1104), .B(n1103), .Z(n1253) );
  NAND U1544 ( .A(x[78]), .B(y[197]), .Z(n1455) );
  NANDN U1545 ( .A(n1455), .B(n1654), .Z(n1108) );
  NANDN U1546 ( .A(n1106), .B(n1105), .Z(n1107) );
  AND U1547 ( .A(n1108), .B(n1107), .Z(n1247) );
  AND U1548 ( .A(x[73]), .B(y[206]), .Z(n2075) );
  NAND U1549 ( .A(n1233), .B(n2075), .Z(n1112) );
  NANDN U1550 ( .A(n1110), .B(n1109), .Z(n1111) );
  NAND U1551 ( .A(n1112), .B(n1111), .Z(n1246) );
  XNOR U1552 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U1553 ( .A(y[204]), .B(x[69]), .Z(n1286) );
  NAND U1554 ( .A(x[72]), .B(y[201]), .Z(n1113) );
  XNOR U1555 ( .A(n1286), .B(n1113), .Z(n1226) );
  XOR U1556 ( .A(n1226), .B(n1225), .Z(n1240) );
  NAND U1557 ( .A(x[71]), .B(y[202]), .Z(n1241) );
  NAND U1558 ( .A(y[205]), .B(x[68]), .Z(n1114) );
  XNOR U1559 ( .A(n1115), .B(n1114), .Z(n1192) );
  NAND U1560 ( .A(x[75]), .B(y[198]), .Z(n1193) );
  XOR U1561 ( .A(n1192), .B(n1193), .Z(n1243) );
  XOR U1562 ( .A(n1242), .B(n1243), .Z(n1249) );
  XNOR U1563 ( .A(n1248), .B(n1249), .Z(n1252) );
  XOR U1564 ( .A(n1253), .B(n1252), .Z(n1255) );
  XOR U1565 ( .A(n1254), .B(n1255), .Z(n1175) );
  NANDN U1566 ( .A(n1117), .B(n1116), .Z(n1121) );
  NANDN U1567 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U1568 ( .A(n1121), .B(n1120), .Z(n1174) );
  NANDN U1569 ( .A(n1123), .B(n1122), .Z(n1127) );
  NANDN U1570 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1571 ( .A(n1127), .B(n1126), .Z(n1183) );
  NAND U1572 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U1573 ( .A(n1131), .B(n1130), .Z(n1132) );
  NAND U1574 ( .A(n1133), .B(n1132), .Z(n1261) );
  AND U1575 ( .A(y[203]), .B(x[77]), .Z(n2094) );
  AND U1576 ( .A(x[69]), .B(y[195]), .Z(n1134) );
  NAND U1577 ( .A(n2094), .B(n1134), .Z(n1137) );
  NANDN U1578 ( .A(n1135), .B(n1818), .Z(n1136) );
  NAND U1579 ( .A(n1137), .B(n1136), .Z(n1214) );
  AND U1580 ( .A(y[208]), .B(x[65]), .Z(n1139) );
  NAND U1581 ( .A(x[73]), .B(y[200]), .Z(n1138) );
  XNOR U1582 ( .A(n1139), .B(n1138), .Z(n1229) );
  NAND U1583 ( .A(n1140), .B(o[16]), .Z(n1230) );
  XNOR U1584 ( .A(n1229), .B(n1230), .Z(n1213) );
  AND U1585 ( .A(y[197]), .B(x[76]), .Z(n1142) );
  NAND U1586 ( .A(x[79]), .B(y[194]), .Z(n1141) );
  XNOR U1587 ( .A(n1142), .B(n1141), .Z(n1188) );
  AND U1588 ( .A(y[195]), .B(x[78]), .Z(n1187) );
  XOR U1589 ( .A(n1188), .B(n1187), .Z(n1212) );
  XOR U1590 ( .A(n1213), .B(n1212), .Z(n1215) );
  XOR U1591 ( .A(n1214), .B(n1215), .Z(n1259) );
  NAND U1592 ( .A(y[207]), .B(x[72]), .Z(n1910) );
  AND U1593 ( .A(y[200]), .B(x[65]), .Z(n1304) );
  XOR U1594 ( .A(n1220), .B(n1221), .Z(n1222) );
  AND U1595 ( .A(x[64]), .B(y[209]), .Z(n1202) );
  AND U1596 ( .A(x[81]), .B(y[192]), .Z(n1201) );
  XOR U1597 ( .A(n1202), .B(n1201), .Z(n1204) );
  AND U1598 ( .A(x[80]), .B(y[193]), .Z(n1198) );
  XOR U1599 ( .A(n1198), .B(o[17]), .Z(n1203) );
  XOR U1600 ( .A(n1204), .B(n1203), .Z(n1217) );
  AND U1601 ( .A(x[74]), .B(y[199]), .Z(n1153) );
  NAND U1602 ( .A(x[66]), .B(y[207]), .Z(n1152) );
  XNOR U1603 ( .A(n1153), .B(n1152), .Z(n1234) );
  NAND U1604 ( .A(y[206]), .B(x[67]), .Z(n1235) );
  XNOR U1605 ( .A(n1234), .B(n1235), .Z(n1216) );
  XOR U1606 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U1607 ( .A(n1219), .B(n1218), .Z(n1223) );
  XNOR U1608 ( .A(n1222), .B(n1223), .Z(n1258) );
  XOR U1609 ( .A(n1259), .B(n1258), .Z(n1260) );
  XNOR U1610 ( .A(n1261), .B(n1260), .Z(n1180) );
  NANDN U1611 ( .A(n1155), .B(n1154), .Z(n1159) );
  NANDN U1612 ( .A(n1157), .B(n1156), .Z(n1158) );
  AND U1613 ( .A(n1159), .B(n1158), .Z(n1181) );
  XOR U1614 ( .A(n1180), .B(n1181), .Z(n1182) );
  XOR U1615 ( .A(n1183), .B(n1182), .Z(n1265) );
  XOR U1616 ( .A(n1266), .B(n1265), .Z(n1267) );
  XOR U1617 ( .A(n1268), .B(n1267), .Z(n1264) );
  NANDN U1618 ( .A(n1161), .B(n1160), .Z(n1165) );
  NAND U1619 ( .A(n1163), .B(n1162), .Z(n1164) );
  NAND U1620 ( .A(n1165), .B(n1164), .Z(n1263) );
  NANDN U1621 ( .A(n1166), .B(n1167), .Z(n1172) );
  NOR U1622 ( .A(n1168), .B(n1167), .Z(n1170) );
  OR U1623 ( .A(n1170), .B(n1169), .Z(n1171) );
  AND U1624 ( .A(n1172), .B(n1171), .Z(n1262) );
  XOR U1625 ( .A(n1263), .B(n1262), .Z(n1173) );
  XNOR U1626 ( .A(n1264), .B(n1173), .Z(N50) );
  NANDN U1627 ( .A(n1175), .B(n1174), .Z(n1179) );
  NANDN U1628 ( .A(n1177), .B(n1176), .Z(n1178) );
  AND U1629 ( .A(n1179), .B(n1178), .Z(n1376) );
  NAND U1630 ( .A(n1181), .B(n1180), .Z(n1185) );
  NANDN U1631 ( .A(n1183), .B(n1182), .Z(n1184) );
  AND U1632 ( .A(n1185), .B(n1184), .Z(n1373) );
  AND U1633 ( .A(y[194]), .B(x[76]), .Z(n1507) );
  AND U1634 ( .A(x[79]), .B(y[197]), .Z(n1186) );
  NAND U1635 ( .A(n1507), .B(n1186), .Z(n1190) );
  NAND U1636 ( .A(n1188), .B(n1187), .Z(n1189) );
  NAND U1637 ( .A(n1190), .B(n1189), .Z(n1348) );
  NAND U1638 ( .A(n2426), .B(n1191), .Z(n1195) );
  NANDN U1639 ( .A(n1193), .B(n1192), .Z(n1194) );
  AND U1640 ( .A(n1195), .B(n1194), .Z(n1341) );
  AND U1641 ( .A(y[209]), .B(x[65]), .Z(n1197) );
  NAND U1642 ( .A(x[74]), .B(y[200]), .Z(n1196) );
  XNOR U1643 ( .A(n1197), .B(n1196), .Z(n1305) );
  NAND U1644 ( .A(n1198), .B(o[17]), .Z(n1306) );
  XNOR U1645 ( .A(n1305), .B(n1306), .Z(n1339) );
  AND U1646 ( .A(x[79]), .B(y[195]), .Z(n1200) );
  NAND U1647 ( .A(x[73]), .B(y[201]), .Z(n1199) );
  XNOR U1648 ( .A(n1200), .B(n1199), .Z(n1296) );
  NAND U1649 ( .A(x[78]), .B(y[196]), .Z(n1297) );
  XNOR U1650 ( .A(n1296), .B(n1297), .Z(n1338) );
  XOR U1651 ( .A(n1339), .B(n1338), .Z(n1340) );
  XNOR U1652 ( .A(n1341), .B(n1340), .Z(n1349) );
  XOR U1653 ( .A(n1348), .B(n1349), .Z(n1351) );
  NAND U1654 ( .A(n1202), .B(n1201), .Z(n1206) );
  NAND U1655 ( .A(n1204), .B(n1203), .Z(n1205) );
  NAND U1656 ( .A(n1206), .B(n1205), .Z(n1360) );
  AND U1657 ( .A(y[199]), .B(x[75]), .Z(n1208) );
  NAND U1658 ( .A(y[194]), .B(x[80]), .Z(n1207) );
  XNOR U1659 ( .A(n1208), .B(n1207), .Z(n1292) );
  NAND U1660 ( .A(x[66]), .B(y[208]), .Z(n1293) );
  XNOR U1661 ( .A(n1292), .B(n1293), .Z(n1361) );
  XOR U1662 ( .A(n1360), .B(n1361), .Z(n1363) );
  AND U1663 ( .A(x[70]), .B(y[204]), .Z(n1210) );
  NAND U1664 ( .A(y[205]), .B(x[69]), .Z(n1209) );
  XNOR U1665 ( .A(n1210), .B(n1209), .Z(n1287) );
  NAND U1666 ( .A(y[206]), .B(x[68]), .Z(n1211) );
  XNOR U1667 ( .A(n2080), .B(n1211), .Z(n1327) );
  NAND U1668 ( .A(x[71]), .B(y[203]), .Z(n1328) );
  XOR U1669 ( .A(n1327), .B(n1328), .Z(n1288) );
  XNOR U1670 ( .A(n1287), .B(n1288), .Z(n1362) );
  XOR U1671 ( .A(n1363), .B(n1362), .Z(n1350) );
  XOR U1672 ( .A(n1351), .B(n1350), .Z(n1277) );
  XOR U1673 ( .A(n1343), .B(n1342), .Z(n1345) );
  XOR U1674 ( .A(n1345), .B(n1344), .Z(n1276) );
  XNOR U1675 ( .A(n1277), .B(n1276), .Z(n1279) );
  AND U1676 ( .A(y[204]), .B(x[72]), .Z(n1553) );
  NAND U1677 ( .A(n1553), .B(n1224), .Z(n1228) );
  NAND U1678 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1679 ( .A(n1228), .B(n1227), .Z(n1355) );
  AND U1680 ( .A(x[73]), .B(y[208]), .Z(n2186) );
  NAND U1681 ( .A(n2186), .B(n1304), .Z(n1232) );
  NANDN U1682 ( .A(n1230), .B(n1229), .Z(n1231) );
  NAND U1683 ( .A(n1232), .B(n1231), .Z(n1354) );
  XOR U1684 ( .A(n1355), .B(n1354), .Z(n1357) );
  AND U1685 ( .A(y[207]), .B(x[74]), .Z(n2103) );
  IV U1686 ( .A(n2103), .Z(n2185) );
  NANDN U1687 ( .A(n2185), .B(n1233), .Z(n1237) );
  NANDN U1688 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1689 ( .A(n1237), .B(n1236), .Z(n1337) );
  AND U1690 ( .A(x[64]), .B(y[210]), .Z(n1309) );
  NAND U1691 ( .A(y[192]), .B(x[82]), .Z(n1310) );
  XNOR U1692 ( .A(n1309), .B(n1310), .Z(n1312) );
  NAND U1693 ( .A(x[81]), .B(y[193]), .Z(n1331) );
  XNOR U1694 ( .A(o[18]), .B(n1331), .Z(n1311) );
  XOR U1695 ( .A(n1312), .B(n1311), .Z(n1335) );
  AND U1696 ( .A(y[197]), .B(x[77]), .Z(n1239) );
  NAND U1697 ( .A(y[207]), .B(x[67]), .Z(n1238) );
  XNOR U1698 ( .A(n1239), .B(n1238), .Z(n1318) );
  NAND U1699 ( .A(x[76]), .B(y[198]), .Z(n1319) );
  XNOR U1700 ( .A(n1318), .B(n1319), .Z(n1334) );
  XOR U1701 ( .A(n1335), .B(n1334), .Z(n1336) );
  XNOR U1702 ( .A(n1337), .B(n1336), .Z(n1356) );
  XOR U1703 ( .A(n1357), .B(n1356), .Z(n1281) );
  NANDN U1704 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U1705 ( .A(n1243), .B(n1242), .Z(n1244) );
  AND U1706 ( .A(n1245), .B(n1244), .Z(n1280) );
  XNOR U1707 ( .A(n1281), .B(n1280), .Z(n1283) );
  NANDN U1708 ( .A(n1247), .B(n1246), .Z(n1251) );
  NANDN U1709 ( .A(n1249), .B(n1248), .Z(n1250) );
  AND U1710 ( .A(n1251), .B(n1250), .Z(n1282) );
  XOR U1711 ( .A(n1283), .B(n1282), .Z(n1278) );
  XOR U1712 ( .A(n1279), .B(n1278), .Z(n1275) );
  NANDN U1713 ( .A(n1253), .B(n1252), .Z(n1257) );
  OR U1714 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U1715 ( .A(n1257), .B(n1256), .Z(n1272) );
  XOR U1716 ( .A(n1272), .B(n1273), .Z(n1274) );
  XOR U1717 ( .A(n1275), .B(n1274), .Z(n1374) );
  XNOR U1718 ( .A(n1376), .B(n1375), .Z(n1369) );
  NAND U1719 ( .A(n1266), .B(n1265), .Z(n1270) );
  NANDN U1720 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1721 ( .A(n1270), .B(n1269), .Z(n1367) );
  IV U1722 ( .A(n1367), .Z(n1366) );
  XOR U1723 ( .A(n1368), .B(n1366), .Z(n1271) );
  XNOR U1724 ( .A(n1369), .B(n1271), .Z(N51) );
  NANDN U1725 ( .A(n1281), .B(n1280), .Z(n1285) );
  NAND U1726 ( .A(n1283), .B(n1282), .Z(n1284) );
  AND U1727 ( .A(n1285), .B(n1284), .Z(n1383) );
  AND U1728 ( .A(y[205]), .B(x[70]), .Z(n1333) );
  NAND U1729 ( .A(n1333), .B(n1286), .Z(n1290) );
  NANDN U1730 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U1731 ( .A(n1290), .B(n1289), .Z(n1388) );
  AND U1732 ( .A(x[80]), .B(y[199]), .Z(n1291) );
  NAND U1733 ( .A(n1291), .B(n1654), .Z(n1295) );
  NANDN U1734 ( .A(n1293), .B(n1292), .Z(n1294) );
  AND U1735 ( .A(n1295), .B(n1294), .Z(n1387) );
  AND U1736 ( .A(y[201]), .B(x[79]), .Z(n2106) );
  NAND U1737 ( .A(n2106), .B(n1416), .Z(n1299) );
  NANDN U1738 ( .A(n1297), .B(n1296), .Z(n1298) );
  AND U1739 ( .A(n1299), .B(n1298), .Z(n1407) );
  NAND U1740 ( .A(y[210]), .B(x[65]), .Z(n1300) );
  XNOR U1741 ( .A(n1301), .B(n1300), .Z(n1454) );
  AND U1742 ( .A(x[77]), .B(y[198]), .Z(n1303) );
  NAND U1743 ( .A(y[209]), .B(x[66]), .Z(n1302) );
  XNOR U1744 ( .A(n1303), .B(n1302), .Z(n1422) );
  XOR U1745 ( .A(n1405), .B(n1404), .Z(n1406) );
  XOR U1746 ( .A(n1387), .B(n1386), .Z(n1389) );
  XOR U1747 ( .A(n1388), .B(n1389), .Z(n1381) );
  AND U1748 ( .A(x[74]), .B(y[209]), .Z(n2595) );
  NAND U1749 ( .A(n2595), .B(n1304), .Z(n1308) );
  NANDN U1750 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U1751 ( .A(n1308), .B(n1307), .Z(n1466) );
  NANDN U1752 ( .A(n1310), .B(n1309), .Z(n1314) );
  NAND U1753 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U1754 ( .A(n1314), .B(n1313), .Z(n1464) );
  AND U1755 ( .A(x[73]), .B(y[202]), .Z(n1316) );
  NAND U1756 ( .A(y[195]), .B(x[80]), .Z(n1315) );
  XNOR U1757 ( .A(n1316), .B(n1315), .Z(n1417) );
  NAND U1758 ( .A(x[79]), .B(y[196]), .Z(n1418) );
  XNOR U1759 ( .A(n1417), .B(n1418), .Z(n1463) );
  XNOR U1760 ( .A(n1466), .B(n1465), .Z(n1394) );
  AND U1761 ( .A(y[207]), .B(x[77]), .Z(n2712) );
  NANDN U1762 ( .A(n1317), .B(n2712), .Z(n1321) );
  NANDN U1763 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U1764 ( .A(n1321), .B(n1320), .Z(n1472) );
  AND U1765 ( .A(x[81]), .B(y[194]), .Z(n1323) );
  NAND U1766 ( .A(x[74]), .B(y[201]), .Z(n1322) );
  XNOR U1767 ( .A(n1323), .B(n1322), .Z(n1460) );
  NAND U1768 ( .A(y[193]), .B(x[82]), .Z(n1436) );
  XNOR U1769 ( .A(o[19]), .B(n1436), .Z(n1459) );
  XOR U1770 ( .A(n1460), .B(n1459), .Z(n1470) );
  AND U1771 ( .A(y[208]), .B(x[67]), .Z(n1325) );
  NAND U1772 ( .A(x[75]), .B(y[200]), .Z(n1324) );
  XNOR U1773 ( .A(n1325), .B(n1324), .Z(n1430) );
  XOR U1774 ( .A(n1470), .B(n1469), .Z(n1471) );
  NAND U1775 ( .A(n1703), .B(n1326), .Z(n1330) );
  NANDN U1776 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U1777 ( .A(n1330), .B(n1329), .Z(n1413) );
  AND U1778 ( .A(x[64]), .B(y[211]), .Z(n1441) );
  NAND U1779 ( .A(y[192]), .B(x[83]), .Z(n1442) );
  XNOR U1780 ( .A(n1441), .B(n1442), .Z(n1444) );
  ANDN U1781 ( .B(o[18]), .A(n1331), .Z(n1443) );
  XOR U1782 ( .A(n1444), .B(n1443), .Z(n1411) );
  AND U1783 ( .A(x[68]), .B(y[207]), .Z(n1567) );
  NAND U1784 ( .A(y[206]), .B(x[69]), .Z(n1332) );
  XOR U1785 ( .A(n1333), .B(n1332), .Z(n1438) );
  XNOR U1786 ( .A(n1567), .B(n1438), .Z(n1410) );
  XOR U1787 ( .A(n1411), .B(n1410), .Z(n1412) );
  XNOR U1788 ( .A(n1413), .B(n1412), .Z(n1392) );
  XOR U1789 ( .A(n1393), .B(n1392), .Z(n1395) );
  XOR U1790 ( .A(n1394), .B(n1395), .Z(n1400) );
  XOR U1791 ( .A(n1399), .B(n1398), .Z(n1401) );
  XOR U1792 ( .A(n1400), .B(n1401), .Z(n1380) );
  XNOR U1793 ( .A(n1381), .B(n1380), .Z(n1382) );
  XOR U1794 ( .A(n1383), .B(n1382), .Z(n1483) );
  NAND U1795 ( .A(n1343), .B(n1342), .Z(n1347) );
  NAND U1796 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U1797 ( .A(n1347), .B(n1346), .Z(n1481) );
  NAND U1798 ( .A(n1349), .B(n1348), .Z(n1353) );
  NAND U1799 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1800 ( .A(n1353), .B(n1352), .Z(n1477) );
  NAND U1801 ( .A(n1355), .B(n1354), .Z(n1359) );
  NAND U1802 ( .A(n1357), .B(n1356), .Z(n1358) );
  NAND U1803 ( .A(n1359), .B(n1358), .Z(n1476) );
  NAND U1804 ( .A(n1361), .B(n1360), .Z(n1365) );
  NAND U1805 ( .A(n1363), .B(n1362), .Z(n1364) );
  NAND U1806 ( .A(n1365), .B(n1364), .Z(n1475) );
  XNOR U1807 ( .A(n1476), .B(n1475), .Z(n1478) );
  XOR U1808 ( .A(n1477), .B(n1478), .Z(n1482) );
  XNOR U1809 ( .A(n1481), .B(n1482), .Z(n1484) );
  XOR U1810 ( .A(n1483), .B(n1484), .Z(n1494) );
  XNOR U1811 ( .A(n1495), .B(n1494), .Z(n1497) );
  XOR U1812 ( .A(n1496), .B(n1497), .Z(n1490) );
  OR U1813 ( .A(n1368), .B(n1366), .Z(n1372) );
  ANDN U1814 ( .B(n1368), .A(n1367), .Z(n1370) );
  OR U1815 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1816 ( .A(n1372), .B(n1371), .Z(n1489) );
  NANDN U1817 ( .A(n1374), .B(n1373), .Z(n1378) );
  NAND U1818 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U1819 ( .A(n1378), .B(n1377), .Z(n1488) );
  IV U1820 ( .A(n1488), .Z(n1487) );
  XOR U1821 ( .A(n1489), .B(n1487), .Z(n1379) );
  XNOR U1822 ( .A(n1490), .B(n1379), .Z(N52) );
  NANDN U1823 ( .A(n1381), .B(n1380), .Z(n1385) );
  NANDN U1824 ( .A(n1383), .B(n1382), .Z(n1384) );
  AND U1825 ( .A(n1385), .B(n1384), .Z(n1604) );
  NANDN U1826 ( .A(n1387), .B(n1386), .Z(n1391) );
  OR U1827 ( .A(n1389), .B(n1388), .Z(n1390) );
  AND U1828 ( .A(n1391), .B(n1390), .Z(n1611) );
  NANDN U1829 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U1830 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U1831 ( .A(n1397), .B(n1396), .Z(n1609) );
  NANDN U1832 ( .A(n1399), .B(n1398), .Z(n1403) );
  NANDN U1833 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1834 ( .A(n1403), .B(n1402), .Z(n1608) );
  XNOR U1835 ( .A(n1609), .B(n1608), .Z(n1610) );
  XOR U1836 ( .A(n1611), .B(n1610), .Z(n1603) );
  NAND U1837 ( .A(n1405), .B(n1404), .Z(n1409) );
  NANDN U1838 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U1839 ( .A(n1409), .B(n1408), .Z(n1502) );
  NAND U1840 ( .A(n1411), .B(n1410), .Z(n1415) );
  NAND U1841 ( .A(n1413), .B(n1412), .Z(n1414) );
  NAND U1842 ( .A(n1415), .B(n1414), .Z(n1501) );
  AND U1843 ( .A(x[80]), .B(y[202]), .Z(n2338) );
  NAND U1844 ( .A(n2338), .B(n1416), .Z(n1420) );
  NANDN U1845 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U1846 ( .A(n1420), .B(n1419), .Z(n1542) );
  AND U1847 ( .A(x[77]), .B(y[209]), .Z(n2942) );
  NAND U1848 ( .A(n2942), .B(n1421), .Z(n1425) );
  NANDN U1849 ( .A(n1423), .B(n1422), .Z(n1424) );
  AND U1850 ( .A(n1425), .B(n1424), .Z(n1587) );
  NAND U1851 ( .A(y[196]), .B(x[80]), .Z(n1426) );
  XNOR U1852 ( .A(n1427), .B(n1426), .Z(n1548) );
  NAND U1853 ( .A(y[210]), .B(x[66]), .Z(n1549) );
  XNOR U1854 ( .A(n1548), .B(n1549), .Z(n1585) );
  NAND U1855 ( .A(y[197]), .B(x[79]), .Z(n1428) );
  XNOR U1856 ( .A(n1429), .B(n1428), .Z(n1518) );
  NAND U1857 ( .A(x[78]), .B(y[198]), .Z(n1519) );
  XNOR U1858 ( .A(n1518), .B(n1519), .Z(n1584) );
  XOR U1859 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U1860 ( .A(n1587), .B(n1586), .Z(n1541) );
  XNOR U1861 ( .A(n1542), .B(n1541), .Z(n1544) );
  AND U1862 ( .A(x[75]), .B(y[208]), .Z(n2598) );
  NANDN U1863 ( .A(n1682), .B(n2598), .Z(n1433) );
  NANDN U1864 ( .A(n1431), .B(n1430), .Z(n1432) );
  AND U1865 ( .A(n1433), .B(n1432), .Z(n1593) );
  AND U1866 ( .A(y[211]), .B(x[65]), .Z(n1435) );
  NAND U1867 ( .A(x[75]), .B(y[201]), .Z(n1434) );
  XNOR U1868 ( .A(n1435), .B(n1434), .Z(n1514) );
  NAND U1869 ( .A(y[193]), .B(x[83]), .Z(n1522) );
  XNOR U1870 ( .A(o[20]), .B(n1522), .Z(n1513) );
  XOR U1871 ( .A(n1514), .B(n1513), .Z(n1591) );
  AND U1872 ( .A(y[212]), .B(x[64]), .Z(n1572) );
  NAND U1873 ( .A(y[192]), .B(x[84]), .Z(n1573) );
  XNOR U1874 ( .A(n1572), .B(n1573), .Z(n1575) );
  ANDN U1875 ( .B(o[19]), .A(n1436), .Z(n1574) );
  XOR U1876 ( .A(n1575), .B(n1574), .Z(n1590) );
  XOR U1877 ( .A(n1591), .B(n1590), .Z(n1592) );
  XNOR U1878 ( .A(n1593), .B(n1592), .Z(n1543) );
  XOR U1879 ( .A(n1544), .B(n1543), .Z(n1503) );
  XOR U1880 ( .A(n1504), .B(n1503), .Z(n1599) );
  AND U1881 ( .A(y[206]), .B(x[70]), .Z(n1524) );
  AND U1882 ( .A(x[69]), .B(y[205]), .Z(n1437) );
  NAND U1883 ( .A(n1524), .B(n1437), .Z(n1440) );
  NANDN U1884 ( .A(n1438), .B(n1567), .Z(n1439) );
  AND U1885 ( .A(n1440), .B(n1439), .Z(n1532) );
  NANDN U1886 ( .A(n1442), .B(n1441), .Z(n1446) );
  NAND U1887 ( .A(n1444), .B(n1443), .Z(n1445) );
  AND U1888 ( .A(n1446), .B(n1445), .Z(n1530) );
  AND U1889 ( .A(x[76]), .B(y[200]), .Z(n1448) );
  NAND U1890 ( .A(x[82]), .B(y[194]), .Z(n1447) );
  XNOR U1891 ( .A(n1448), .B(n1447), .Z(n1508) );
  NAND U1892 ( .A(x[81]), .B(y[195]), .Z(n1509) );
  XNOR U1893 ( .A(n1508), .B(n1509), .Z(n1529) );
  XNOR U1894 ( .A(n1530), .B(n1529), .Z(n1531) );
  XOR U1895 ( .A(n1532), .B(n1531), .Z(n1536) );
  AND U1896 ( .A(x[77]), .B(y[199]), .Z(n1450) );
  NAND U1897 ( .A(y[209]), .B(x[67]), .Z(n1449) );
  XNOR U1898 ( .A(n1450), .B(n1449), .Z(n1554) );
  XOR U1899 ( .A(n1554), .B(n1553), .Z(n1526) );
  AND U1900 ( .A(y[207]), .B(x[69]), .Z(n1452) );
  NAND U1901 ( .A(y[208]), .B(x[68]), .Z(n1451) );
  XNOR U1902 ( .A(n1452), .B(n1451), .Z(n1569) );
  AND U1903 ( .A(y[205]), .B(x[71]), .Z(n1568) );
  XNOR U1904 ( .A(n1569), .B(n1568), .Z(n1523) );
  XNOR U1905 ( .A(n1524), .B(n1523), .Z(n1525) );
  XOR U1906 ( .A(n1526), .B(n1525), .Z(n1580) );
  AND U1907 ( .A(y[210]), .B(x[72]), .Z(n2659) );
  AND U1908 ( .A(x[65]), .B(y[203]), .Z(n1453) );
  NAND U1909 ( .A(n2659), .B(n1453), .Z(n1457) );
  NANDN U1910 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1911 ( .A(n1457), .B(n1456), .Z(n1579) );
  AND U1912 ( .A(y[201]), .B(x[81]), .Z(n2344) );
  NAND U1913 ( .A(n2344), .B(n1458), .Z(n1462) );
  NAND U1914 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1915 ( .A(n1462), .B(n1461), .Z(n1578) );
  XNOR U1916 ( .A(n1579), .B(n1578), .Z(n1581) );
  XNOR U1917 ( .A(n1580), .B(n1581), .Z(n1535) );
  XOR U1918 ( .A(n1536), .B(n1535), .Z(n1537) );
  NANDN U1919 ( .A(n1464), .B(n1463), .Z(n1468) );
  NAND U1920 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1921 ( .A(n1468), .B(n1467), .Z(n1538) );
  NAND U1922 ( .A(n1470), .B(n1469), .Z(n1474) );
  NANDN U1923 ( .A(n1472), .B(n1471), .Z(n1473) );
  NAND U1924 ( .A(n1474), .B(n1473), .Z(n1597) );
  XOR U1925 ( .A(n1599), .B(n1598), .Z(n1602) );
  XOR U1926 ( .A(n1603), .B(n1602), .Z(n1605) );
  XOR U1927 ( .A(n1604), .B(n1605), .Z(n1619) );
  NAND U1928 ( .A(n1476), .B(n1475), .Z(n1480) );
  NANDN U1929 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U1930 ( .A(n1480), .B(n1479), .Z(n1618) );
  NANDN U1931 ( .A(n1482), .B(n1481), .Z(n1486) );
  NAND U1932 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1933 ( .A(n1486), .B(n1485), .Z(n1617) );
  XOR U1934 ( .A(n1618), .B(n1617), .Z(n1620) );
  XNOR U1935 ( .A(n1619), .B(n1620), .Z(n1614) );
  OR U1936 ( .A(n1489), .B(n1487), .Z(n1493) );
  ANDN U1937 ( .B(n1489), .A(n1488), .Z(n1491) );
  OR U1938 ( .A(n1491), .B(n1490), .Z(n1492) );
  AND U1939 ( .A(n1493), .B(n1492), .Z(n1616) );
  NAND U1940 ( .A(n1495), .B(n1494), .Z(n1499) );
  NANDN U1941 ( .A(n1497), .B(n1496), .Z(n1498) );
  NAND U1942 ( .A(n1499), .B(n1498), .Z(n1615) );
  XOR U1943 ( .A(n1616), .B(n1615), .Z(n1500) );
  XNOR U1944 ( .A(n1614), .B(n1500), .Z(N53) );
  NANDN U1945 ( .A(n1502), .B(n1501), .Z(n1506) );
  NAND U1946 ( .A(n1504), .B(n1503), .Z(n1505) );
  AND U1947 ( .A(n1506), .B(n1505), .Z(n1633) );
  NAND U1948 ( .A(y[200]), .B(x[82]), .Z(n2347) );
  NANDN U1949 ( .A(n2347), .B(n1507), .Z(n1511) );
  NANDN U1950 ( .A(n1509), .B(n1508), .Z(n1510) );
  AND U1951 ( .A(n1511), .B(n1510), .Z(n1711) );
  AND U1952 ( .A(x[75]), .B(y[211]), .Z(n3148) );
  AND U1953 ( .A(y[201]), .B(x[65]), .Z(n1512) );
  NAND U1954 ( .A(n3148), .B(n1512), .Z(n1516) );
  NAND U1955 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U1956 ( .A(n1516), .B(n1515), .Z(n1710) );
  XNOR U1957 ( .A(n1711), .B(n1710), .Z(n1713) );
  AND U1958 ( .A(x[79]), .B(y[203]), .Z(n2333) );
  NAND U1959 ( .A(n2333), .B(n1517), .Z(n1521) );
  NANDN U1960 ( .A(n1519), .B(n1518), .Z(n1520) );
  NAND U1961 ( .A(n1521), .B(n1520), .Z(n1667) );
  AND U1962 ( .A(y[213]), .B(x[64]), .Z(n1688) );
  NAND U1963 ( .A(y[192]), .B(x[85]), .Z(n1689) );
  XNOR U1964 ( .A(n1688), .B(n1689), .Z(n1691) );
  ANDN U1965 ( .B(o[20]), .A(n1522), .Z(n1690) );
  XOR U1966 ( .A(n1691), .B(n1690), .Z(n1666) );
  AND U1967 ( .A(x[69]), .B(y[208]), .Z(n1672) );
  AND U1968 ( .A(x[80]), .B(y[197]), .Z(n1671) );
  XOR U1969 ( .A(n1672), .B(n1671), .Z(n1674) );
  AND U1970 ( .A(x[79]), .B(y[198]), .Z(n1673) );
  XOR U1971 ( .A(n1674), .B(n1673), .Z(n1665) );
  XOR U1972 ( .A(n1666), .B(n1665), .Z(n1668) );
  XOR U1973 ( .A(n1667), .B(n1668), .Z(n1712) );
  XOR U1974 ( .A(n1713), .B(n1712), .Z(n1705) );
  NANDN U1975 ( .A(n1524), .B(n1523), .Z(n1528) );
  NANDN U1976 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1977 ( .A(n1528), .B(n1527), .Z(n1704) );
  XNOR U1978 ( .A(n1705), .B(n1704), .Z(n1707) );
  NANDN U1979 ( .A(n1530), .B(n1529), .Z(n1534) );
  NANDN U1980 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1981 ( .A(n1534), .B(n1533), .Z(n1706) );
  XOR U1982 ( .A(n1707), .B(n1706), .Z(n1631) );
  NAND U1983 ( .A(n1536), .B(n1535), .Z(n1540) );
  NANDN U1984 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1985 ( .A(n1540), .B(n1539), .Z(n1630) );
  NANDN U1986 ( .A(n1542), .B(n1541), .Z(n1546) );
  NAND U1987 ( .A(n1544), .B(n1543), .Z(n1545) );
  AND U1988 ( .A(n1546), .B(n1545), .Z(n1731) );
  NAND U1989 ( .A(n2338), .B(n1547), .Z(n1551) );
  NANDN U1990 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U1991 ( .A(n1551), .B(n1550), .Z(n1637) );
  NAND U1992 ( .A(n2942), .B(n1552), .Z(n1556) );
  NAND U1993 ( .A(n1554), .B(n1553), .Z(n1555) );
  AND U1994 ( .A(n1556), .B(n1555), .Z(n1725) );
  AND U1995 ( .A(y[202]), .B(x[75]), .Z(n1558) );
  NAND U1996 ( .A(x[83]), .B(y[194]), .Z(n1557) );
  XNOR U1997 ( .A(n1558), .B(n1557), .Z(n1656) );
  AND U1998 ( .A(y[193]), .B(x[84]), .Z(n1687) );
  XOR U1999 ( .A(n1687), .B(o[21]), .Z(n1655) );
  XOR U2000 ( .A(n1656), .B(n1655), .Z(n1723) );
  NAND U2001 ( .A(x[82]), .B(y[195]), .Z(n1559) );
  XNOR U2002 ( .A(n1560), .B(n1559), .Z(n1695) );
  NAND U2003 ( .A(y[212]), .B(x[65]), .Z(n1696) );
  XNOR U2004 ( .A(n1695), .B(n1696), .Z(n1722) );
  XOR U2005 ( .A(n1723), .B(n1722), .Z(n1724) );
  XNOR U2006 ( .A(n1725), .B(n1724), .Z(n1636) );
  XNOR U2007 ( .A(n1637), .B(n1636), .Z(n1639) );
  AND U2008 ( .A(x[71]), .B(y[206]), .Z(n1908) );
  AND U2009 ( .A(x[70]), .B(y[207]), .Z(n1562) );
  NAND U2010 ( .A(y[199]), .B(x[78]), .Z(n1561) );
  XOR U2011 ( .A(n1562), .B(n1561), .Z(n1699) );
  XNOR U2012 ( .A(n1908), .B(n1699), .Z(n1645) );
  NAND U2013 ( .A(y[204]), .B(x[73]), .Z(n1643) );
  NAND U2014 ( .A(y[205]), .B(x[72]), .Z(n1642) );
  XOR U2015 ( .A(n1643), .B(n1642), .Z(n1644) );
  AND U2016 ( .A(y[196]), .B(x[81]), .Z(n1564) );
  NAND U2017 ( .A(x[76]), .B(y[201]), .Z(n1563) );
  XNOR U2018 ( .A(n1564), .B(n1563), .Z(n1648) );
  NAND U2019 ( .A(y[211]), .B(x[66]), .Z(n1649) );
  XNOR U2020 ( .A(n1648), .B(n1649), .Z(n1660) );
  AND U2021 ( .A(x[67]), .B(y[210]), .Z(n1566) );
  NAND U2022 ( .A(x[77]), .B(y[200]), .Z(n1565) );
  XNOR U2023 ( .A(n1566), .B(n1565), .Z(n1684) );
  AND U2024 ( .A(x[68]), .B(y[209]), .Z(n1683) );
  XOR U2025 ( .A(n1684), .B(n1683), .Z(n1659) );
  XOR U2026 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U2027 ( .A(n1672), .B(n1567), .Z(n1571) );
  NAND U2028 ( .A(n1569), .B(n1568), .Z(n1570) );
  AND U2029 ( .A(n1571), .B(n1570), .Z(n1717) );
  NANDN U2030 ( .A(n1573), .B(n1572), .Z(n1577) );
  NAND U2031 ( .A(n1575), .B(n1574), .Z(n1576) );
  NAND U2032 ( .A(n1577), .B(n1576), .Z(n1716) );
  XNOR U2033 ( .A(n1717), .B(n1716), .Z(n1718) );
  XOR U2034 ( .A(n1719), .B(n1718), .Z(n1638) );
  XOR U2035 ( .A(n1639), .B(n1638), .Z(n1729) );
  NANDN U2036 ( .A(n1579), .B(n1578), .Z(n1583) );
  NAND U2037 ( .A(n1581), .B(n1580), .Z(n1582) );
  NAND U2038 ( .A(n1583), .B(n1582), .Z(n1736) );
  NAND U2039 ( .A(n1585), .B(n1584), .Z(n1589) );
  NANDN U2040 ( .A(n1587), .B(n1586), .Z(n1588) );
  NAND U2041 ( .A(n1589), .B(n1588), .Z(n1735) );
  NAND U2042 ( .A(n1591), .B(n1590), .Z(n1595) );
  NANDN U2043 ( .A(n1593), .B(n1592), .Z(n1594) );
  NAND U2044 ( .A(n1595), .B(n1594), .Z(n1734) );
  XOR U2045 ( .A(n1735), .B(n1734), .Z(n1737) );
  XOR U2046 ( .A(n1736), .B(n1737), .Z(n1728) );
  XOR U2047 ( .A(n1729), .B(n1728), .Z(n1730) );
  XOR U2048 ( .A(n1731), .B(n1730), .Z(n1625) );
  NANDN U2049 ( .A(n1597), .B(n1596), .Z(n1601) );
  NANDN U2050 ( .A(n1599), .B(n1598), .Z(n1600) );
  NAND U2051 ( .A(n1601), .B(n1600), .Z(n1624) );
  XOR U2052 ( .A(n1625), .B(n1624), .Z(n1627) );
  XNOR U2053 ( .A(n1626), .B(n1627), .Z(n1742) );
  NANDN U2054 ( .A(n1603), .B(n1602), .Z(n1607) );
  NANDN U2055 ( .A(n1605), .B(n1604), .Z(n1606) );
  AND U2056 ( .A(n1607), .B(n1606), .Z(n1741) );
  NANDN U2057 ( .A(n1609), .B(n1608), .Z(n1613) );
  NAND U2058 ( .A(n1611), .B(n1610), .Z(n1612) );
  AND U2059 ( .A(n1613), .B(n1612), .Z(n1740) );
  XNOR U2060 ( .A(n1741), .B(n1740), .Z(n1743) );
  XOR U2061 ( .A(n1742), .B(n1743), .Z(n1746) );
  NAND U2062 ( .A(n1618), .B(n1617), .Z(n1622) );
  NAND U2063 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U2064 ( .A(n1622), .B(n1621), .Z(n1744) );
  XOR U2065 ( .A(n1745), .B(n1744), .Z(n1623) );
  XNOR U2066 ( .A(n1746), .B(n1623), .Z(N54) );
  NAND U2067 ( .A(n1625), .B(n1624), .Z(n1629) );
  NAND U2068 ( .A(n1627), .B(n1626), .Z(n1628) );
  AND U2069 ( .A(n1629), .B(n1628), .Z(n1751) );
  NANDN U2070 ( .A(n1631), .B(n1630), .Z(n1635) );
  NANDN U2071 ( .A(n1633), .B(n1632), .Z(n1634) );
  AND U2072 ( .A(n1635), .B(n1634), .Z(n1749) );
  NANDN U2073 ( .A(n1637), .B(n1636), .Z(n1641) );
  NAND U2074 ( .A(n1639), .B(n1638), .Z(n1640) );
  AND U2075 ( .A(n1641), .B(n1640), .Z(n1872) );
  NAND U2076 ( .A(n1643), .B(n1642), .Z(n1647) );
  NANDN U2077 ( .A(n1645), .B(n1644), .Z(n1646) );
  AND U2078 ( .A(n1647), .B(n1646), .Z(n1866) );
  NAND U2079 ( .A(n2344), .B(n1818), .Z(n1651) );
  NANDN U2080 ( .A(n1649), .B(n1648), .Z(n1650) );
  AND U2081 ( .A(n1651), .B(n1650), .Z(n1796) );
  AND U2082 ( .A(x[69]), .B(y[209]), .Z(n1840) );
  AND U2083 ( .A(x[81]), .B(y[197]), .Z(n1839) );
  XOR U2084 ( .A(n1840), .B(n1839), .Z(n1842) );
  AND U2085 ( .A(x[80]), .B(y[198]), .Z(n1841) );
  XOR U2086 ( .A(n1842), .B(n1841), .Z(n1794) );
  AND U2087 ( .A(y[196]), .B(x[82]), .Z(n1653) );
  NAND U2088 ( .A(y[202]), .B(x[76]), .Z(n1652) );
  XNOR U2089 ( .A(n1653), .B(n1652), .Z(n1820) );
  AND U2090 ( .A(x[68]), .B(y[210]), .Z(n1819) );
  XOR U2091 ( .A(n1820), .B(n1819), .Z(n1793) );
  XOR U2092 ( .A(n1794), .B(n1793), .Z(n1795) );
  XOR U2093 ( .A(n1796), .B(n1795), .Z(n1863) );
  AND U2094 ( .A(x[83]), .B(y[202]), .Z(n2837) );
  NAND U2095 ( .A(n2837), .B(n1654), .Z(n1658) );
  NAND U2096 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U2097 ( .A(n1658), .B(n1657), .Z(n1864) );
  XOR U2098 ( .A(n1863), .B(n1864), .Z(n1865) );
  XOR U2099 ( .A(n1866), .B(n1865), .Z(n1869) );
  NAND U2100 ( .A(n1660), .B(n1659), .Z(n1664) );
  NANDN U2101 ( .A(n1662), .B(n1661), .Z(n1663) );
  AND U2102 ( .A(n1664), .B(n1663), .Z(n1852) );
  NAND U2103 ( .A(n1666), .B(n1665), .Z(n1670) );
  NAND U2104 ( .A(n1668), .B(n1667), .Z(n1669) );
  NAND U2105 ( .A(n1670), .B(n1669), .Z(n1851) );
  XNOR U2106 ( .A(n1852), .B(n1851), .Z(n1854) );
  NAND U2107 ( .A(n1672), .B(n1671), .Z(n1676) );
  AND U2108 ( .A(n1674), .B(n1673), .Z(n1675) );
  ANDN U2109 ( .B(n1676), .A(n1675), .Z(n1815) );
  AND U2110 ( .A(x[84]), .B(y[194]), .Z(n1678) );
  NAND U2111 ( .A(x[77]), .B(y[201]), .Z(n1677) );
  XNOR U2112 ( .A(n1678), .B(n1677), .Z(n1836) );
  AND U2113 ( .A(y[212]), .B(x[66]), .Z(n1835) );
  XOR U2114 ( .A(n1836), .B(n1835), .Z(n1813) );
  AND U2115 ( .A(y[208]), .B(x[70]), .Z(n1680) );
  NAND U2116 ( .A(x[79]), .B(y[199]), .Z(n1679) );
  XNOR U2117 ( .A(n1680), .B(n1679), .Z(n1847) );
  XOR U2118 ( .A(n1847), .B(n1681), .Z(n1812) );
  XOR U2119 ( .A(n1813), .B(n1812), .Z(n1814) );
  XNOR U2120 ( .A(n1815), .B(n1814), .Z(n1858) );
  AND U2121 ( .A(y[210]), .B(x[77]), .Z(n3146) );
  NANDN U2122 ( .A(n1682), .B(n3146), .Z(n1686) );
  NAND U2123 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2124 ( .A(n1686), .B(n1685), .Z(n1784) );
  AND U2125 ( .A(y[213]), .B(x[65]), .Z(n1807) );
  XOR U2126 ( .A(n1808), .B(n1807), .Z(n1806) );
  NAND U2127 ( .A(n1687), .B(o[21]), .Z(n1805) );
  XNOR U2128 ( .A(n1806), .B(n1805), .Z(n1781) );
  AND U2129 ( .A(y[200]), .B(x[78]), .Z(n1799) );
  NAND U2130 ( .A(x[67]), .B(y[211]), .Z(n1800) );
  XNOR U2131 ( .A(n1799), .B(n1800), .Z(n1801) );
  NAND U2132 ( .A(y[195]), .B(x[83]), .Z(n1802) );
  XOR U2133 ( .A(n1801), .B(n1802), .Z(n1782) );
  XNOR U2134 ( .A(n1781), .B(n1782), .Z(n1783) );
  XNOR U2135 ( .A(n1784), .B(n1783), .Z(n1857) );
  XOR U2136 ( .A(n1858), .B(n1857), .Z(n1860) );
  NANDN U2137 ( .A(n1689), .B(n1688), .Z(n1693) );
  NAND U2138 ( .A(n1691), .B(n1690), .Z(n1692) );
  AND U2139 ( .A(n1693), .B(n1692), .Z(n1776) );
  AND U2140 ( .A(x[82]), .B(y[203]), .Z(n2839) );
  NAND U2141 ( .A(n2839), .B(n1694), .Z(n1698) );
  NANDN U2142 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U2143 ( .A(n1698), .B(n1697), .Z(n1775) );
  XNOR U2144 ( .A(n1776), .B(n1775), .Z(n1778) );
  AND U2145 ( .A(x[78]), .B(y[207]), .Z(n2849) );
  NAND U2146 ( .A(n1846), .B(n2849), .Z(n1701) );
  NANDN U2147 ( .A(n1699), .B(n1908), .Z(n1700) );
  NAND U2148 ( .A(n1701), .B(n1700), .Z(n1789) );
  AND U2149 ( .A(x[64]), .B(y[214]), .Z(n1824) );
  AND U2150 ( .A(x[86]), .B(y[192]), .Z(n1823) );
  XOR U2151 ( .A(n1824), .B(n1823), .Z(n1826) );
  AND U2152 ( .A(y[193]), .B(x[85]), .Z(n1845) );
  XOR U2153 ( .A(n1845), .B(o[22]), .Z(n1825) );
  XOR U2154 ( .A(n1826), .B(n1825), .Z(n1788) );
  NAND U2155 ( .A(y[207]), .B(x[71]), .Z(n1702) );
  XNOR U2156 ( .A(n1703), .B(n1702), .Z(n1830) );
  XOR U2157 ( .A(n1830), .B(n1829), .Z(n1787) );
  XOR U2158 ( .A(n1788), .B(n1787), .Z(n1790) );
  XOR U2159 ( .A(n1789), .B(n1790), .Z(n1777) );
  XOR U2160 ( .A(n1778), .B(n1777), .Z(n1859) );
  XOR U2161 ( .A(n1860), .B(n1859), .Z(n1853) );
  XOR U2162 ( .A(n1854), .B(n1853), .Z(n1870) );
  XOR U2163 ( .A(n1869), .B(n1870), .Z(n1871) );
  XOR U2164 ( .A(n1872), .B(n1871), .Z(n1765) );
  NANDN U2165 ( .A(n1705), .B(n1704), .Z(n1709) );
  NAND U2166 ( .A(n1707), .B(n1706), .Z(n1708) );
  AND U2167 ( .A(n1709), .B(n1708), .Z(n1764) );
  NANDN U2168 ( .A(n1711), .B(n1710), .Z(n1715) );
  NAND U2169 ( .A(n1713), .B(n1712), .Z(n1714) );
  AND U2170 ( .A(n1715), .B(n1714), .Z(n1772) );
  NANDN U2171 ( .A(n1717), .B(n1716), .Z(n1721) );
  NAND U2172 ( .A(n1719), .B(n1718), .Z(n1720) );
  AND U2173 ( .A(n1721), .B(n1720), .Z(n1770) );
  NAND U2174 ( .A(n1723), .B(n1722), .Z(n1727) );
  NANDN U2175 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U2176 ( .A(n1727), .B(n1726), .Z(n1769) );
  XNOR U2177 ( .A(n1770), .B(n1769), .Z(n1771) );
  XOR U2178 ( .A(n1772), .B(n1771), .Z(n1763) );
  XNOR U2179 ( .A(n1764), .B(n1763), .Z(n1766) );
  XNOR U2180 ( .A(n1765), .B(n1766), .Z(n1759) );
  NAND U2181 ( .A(n1729), .B(n1728), .Z(n1733) );
  NANDN U2182 ( .A(n1731), .B(n1730), .Z(n1732) );
  AND U2183 ( .A(n1733), .B(n1732), .Z(n1758) );
  NAND U2184 ( .A(n1735), .B(n1734), .Z(n1739) );
  NAND U2185 ( .A(n1737), .B(n1736), .Z(n1738) );
  NAND U2186 ( .A(n1739), .B(n1738), .Z(n1757) );
  XNOR U2187 ( .A(n1758), .B(n1757), .Z(n1760) );
  XOR U2188 ( .A(n1759), .B(n1760), .Z(n1748) );
  XNOR U2189 ( .A(n1751), .B(n1750), .Z(n1756) );
  XOR U2190 ( .A(n1754), .B(n1755), .Z(n1747) );
  XNOR U2191 ( .A(n1756), .B(n1747), .Z(N55) );
  NANDN U2192 ( .A(n1749), .B(n1748), .Z(n1753) );
  NAND U2193 ( .A(n1751), .B(n1750), .Z(n1752) );
  NAND U2194 ( .A(n1753), .B(n1752), .Z(n1883) );
  IV U2195 ( .A(n1883), .Z(n1882) );
  NANDN U2196 ( .A(n1758), .B(n1757), .Z(n1762) );
  NAND U2197 ( .A(n1760), .B(n1759), .Z(n1761) );
  AND U2198 ( .A(n1762), .B(n1761), .Z(n1879) );
  NANDN U2199 ( .A(n1764), .B(n1763), .Z(n1768) );
  NAND U2200 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U2201 ( .A(n1768), .B(n1767), .Z(n1877) );
  NANDN U2202 ( .A(n1770), .B(n1769), .Z(n1774) );
  NANDN U2203 ( .A(n1772), .B(n1771), .Z(n1773) );
  AND U2204 ( .A(n1774), .B(n1773), .Z(n2004) );
  NANDN U2205 ( .A(n1776), .B(n1775), .Z(n1780) );
  NAND U2206 ( .A(n1778), .B(n1777), .Z(n1779) );
  NAND U2207 ( .A(n1780), .B(n1779), .Z(n1997) );
  NANDN U2208 ( .A(n1782), .B(n1781), .Z(n1786) );
  NANDN U2209 ( .A(n1784), .B(n1783), .Z(n1785) );
  NAND U2210 ( .A(n1786), .B(n1785), .Z(n1996) );
  NAND U2211 ( .A(n1788), .B(n1787), .Z(n1792) );
  NAND U2212 ( .A(n1790), .B(n1789), .Z(n1791) );
  NAND U2213 ( .A(n1792), .B(n1791), .Z(n1995) );
  XOR U2214 ( .A(n1996), .B(n1995), .Z(n1998) );
  XOR U2215 ( .A(n1997), .B(n1998), .Z(n2015) );
  NAND U2216 ( .A(n1794), .B(n1793), .Z(n1798) );
  NANDN U2217 ( .A(n1796), .B(n1795), .Z(n1797) );
  NAND U2218 ( .A(n1798), .B(n1797), .Z(n2013) );
  NANDN U2219 ( .A(n1800), .B(n1799), .Z(n1804) );
  NANDN U2220 ( .A(n1802), .B(n1801), .Z(n1803) );
  AND U2221 ( .A(n1804), .B(n1803), .Z(n1942) );
  ANDN U2222 ( .B(n1806), .A(n1805), .Z(n1810) );
  NAND U2223 ( .A(n1808), .B(n1807), .Z(n1809) );
  NANDN U2224 ( .A(n1810), .B(n1809), .Z(n1941) );
  XNOR U2225 ( .A(n1942), .B(n1941), .Z(n1944) );
  NAND U2226 ( .A(y[208]), .B(x[71]), .Z(n1811) );
  XNOR U2227 ( .A(n2075), .B(n1811), .Z(n1909) );
  NAND U2228 ( .A(y[205]), .B(x[74]), .Z(n1948) );
  XNOR U2229 ( .A(n1947), .B(n1948), .Z(n1949) );
  AND U2230 ( .A(x[70]), .B(y[209]), .Z(n1900) );
  NAND U2231 ( .A(y[200]), .B(x[79]), .Z(n1901) );
  XNOR U2232 ( .A(n1900), .B(n1901), .Z(n1902) );
  NAND U2233 ( .A(y[204]), .B(x[75]), .Z(n1903) );
  XOR U2234 ( .A(n1902), .B(n1903), .Z(n1950) );
  XNOR U2235 ( .A(n1949), .B(n1950), .Z(n1943) );
  XOR U2236 ( .A(n1944), .B(n1943), .Z(n2014) );
  XNOR U2237 ( .A(n2013), .B(n2014), .Z(n2016) );
  NAND U2238 ( .A(n1813), .B(n1812), .Z(n1817) );
  NANDN U2239 ( .A(n1815), .B(n1814), .Z(n1816) );
  NAND U2240 ( .A(n1817), .B(n1816), .Z(n1935) );
  NAND U2241 ( .A(x[82]), .B(y[202]), .Z(n2678) );
  NANDN U2242 ( .A(n2678), .B(n1818), .Z(n1822) );
  NAND U2243 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2244 ( .A(n1822), .B(n1821), .Z(n1972) );
  NAND U2245 ( .A(n1824), .B(n1823), .Z(n1828) );
  NAND U2246 ( .A(n1826), .B(n1825), .Z(n1827) );
  NAND U2247 ( .A(n1828), .B(n1827), .Z(n1971) );
  XOR U2248 ( .A(n1972), .B(n1971), .Z(n1973) );
  NANDN U2249 ( .A(n1910), .B(n1908), .Z(n1832) );
  NAND U2250 ( .A(n1830), .B(n1829), .Z(n1831) );
  NAND U2251 ( .A(n1832), .B(n1831), .Z(n1985) );
  AND U2252 ( .A(x[64]), .B(y[215]), .Z(n1919) );
  NAND U2253 ( .A(x[87]), .B(y[192]), .Z(n1920) );
  XNOR U2254 ( .A(n1919), .B(n1920), .Z(n1921) );
  NAND U2255 ( .A(x[86]), .B(y[193]), .Z(n1899) );
  XOR U2256 ( .A(o[23]), .B(n1899), .Z(n1922) );
  XNOR U2257 ( .A(n1921), .B(n1922), .Z(n1984) );
  AND U2258 ( .A(x[84]), .B(y[195]), .Z(n2500) );
  NAND U2259 ( .A(y[199]), .B(x[80]), .Z(n1833) );
  XNOR U2260 ( .A(n2500), .B(n1833), .Z(n1895) );
  NAND U2261 ( .A(x[83]), .B(y[196]), .Z(n1896) );
  XNOR U2262 ( .A(n1895), .B(n1896), .Z(n1983) );
  XOR U2263 ( .A(n1984), .B(n1983), .Z(n1986) );
  XNOR U2264 ( .A(n1985), .B(n1986), .Z(n1974) );
  XOR U2265 ( .A(n1935), .B(n1936), .Z(n1938) );
  AND U2266 ( .A(y[201]), .B(x[84]), .Z(n2860) );
  AND U2267 ( .A(y[194]), .B(x[77]), .Z(n1834) );
  NAND U2268 ( .A(n2860), .B(n1834), .Z(n1838) );
  NAND U2269 ( .A(n1836), .B(n1835), .Z(n1837) );
  NAND U2270 ( .A(n1838), .B(n1837), .Z(n1929) );
  NAND U2271 ( .A(n1840), .B(n1839), .Z(n1844) );
  NAND U2272 ( .A(n1842), .B(n1841), .Z(n1843) );
  NAND U2273 ( .A(n1844), .B(n1843), .Z(n1991) );
  AND U2274 ( .A(y[202]), .B(x[77]), .Z(n1965) );
  NAND U2275 ( .A(y[213]), .B(x[66]), .Z(n1966) );
  XNOR U2276 ( .A(n1965), .B(n1966), .Z(n1967) );
  NAND U2277 ( .A(y[194]), .B(x[85]), .Z(n1968) );
  XNOR U2278 ( .A(n1967), .B(n1968), .Z(n1990) );
  AND U2279 ( .A(x[76]), .B(y[203]), .Z(n1913) );
  NAND U2280 ( .A(x[65]), .B(y[214]), .Z(n1914) );
  XNOR U2281 ( .A(n1913), .B(n1914), .Z(n1916) );
  AND U2282 ( .A(n1845), .B(o[22]), .Z(n1915) );
  XOR U2283 ( .A(n1916), .B(n1915), .Z(n1989) );
  XOR U2284 ( .A(n1990), .B(n1989), .Z(n1992) );
  XOR U2285 ( .A(n1991), .B(n1992), .Z(n1930) );
  XOR U2286 ( .A(n1929), .B(n1930), .Z(n1932) );
  AND U2287 ( .A(x[79]), .B(y[208]), .Z(n3096) );
  NAND U2288 ( .A(n3096), .B(n1846), .Z(n1850) );
  NANDN U2289 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U2290 ( .A(n1850), .B(n1849), .Z(n1979) );
  AND U2291 ( .A(y[201]), .B(x[78]), .Z(n1959) );
  NAND U2292 ( .A(y[212]), .B(x[67]), .Z(n1960) );
  XNOR U2293 ( .A(n1959), .B(n1960), .Z(n1961) );
  NAND U2294 ( .A(x[68]), .B(y[211]), .Z(n1962) );
  XNOR U2295 ( .A(n1961), .B(n1962), .Z(n1978) );
  AND U2296 ( .A(x[69]), .B(y[210]), .Z(n1953) );
  NAND U2297 ( .A(x[82]), .B(y[197]), .Z(n1954) );
  XNOR U2298 ( .A(n1953), .B(n1954), .Z(n1956) );
  AND U2299 ( .A(x[81]), .B(y[198]), .Z(n1955) );
  XOR U2300 ( .A(n1956), .B(n1955), .Z(n1977) );
  XOR U2301 ( .A(n1978), .B(n1977), .Z(n1980) );
  XOR U2302 ( .A(n1979), .B(n1980), .Z(n1931) );
  XOR U2303 ( .A(n1932), .B(n1931), .Z(n1937) );
  XOR U2304 ( .A(n1938), .B(n1937), .Z(n2001) );
  XOR U2305 ( .A(n2002), .B(n2001), .Z(n2003) );
  XOR U2306 ( .A(n2004), .B(n2003), .Z(n1891) );
  NANDN U2307 ( .A(n1852), .B(n1851), .Z(n1856) );
  NAND U2308 ( .A(n1854), .B(n1853), .Z(n1855) );
  AND U2309 ( .A(n1856), .B(n1855), .Z(n2010) );
  NAND U2310 ( .A(n1858), .B(n1857), .Z(n1862) );
  NAND U2311 ( .A(n1860), .B(n1859), .Z(n1861) );
  AND U2312 ( .A(n1862), .B(n1861), .Z(n2008) );
  NAND U2313 ( .A(n1864), .B(n1863), .Z(n1868) );
  NANDN U2314 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2315 ( .A(n1868), .B(n1867), .Z(n2007) );
  XNOR U2316 ( .A(n2008), .B(n2007), .Z(n2009) );
  XOR U2317 ( .A(n2010), .B(n2009), .Z(n1889) );
  NAND U2318 ( .A(n1870), .B(n1869), .Z(n1874) );
  NANDN U2319 ( .A(n1872), .B(n1871), .Z(n1873) );
  AND U2320 ( .A(n1874), .B(n1873), .Z(n1890) );
  XOR U2321 ( .A(n1889), .B(n1890), .Z(n1892) );
  XOR U2322 ( .A(n1891), .B(n1892), .Z(n1876) );
  XNOR U2323 ( .A(n1877), .B(n1876), .Z(n1878) );
  XOR U2324 ( .A(n1879), .B(n1878), .Z(n1885) );
  XNOR U2325 ( .A(n1884), .B(n1885), .Z(n1875) );
  XOR U2326 ( .A(n1882), .B(n1875), .Z(N56) );
  NANDN U2327 ( .A(n1877), .B(n1876), .Z(n1881) );
  NAND U2328 ( .A(n1879), .B(n1878), .Z(n1880) );
  NAND U2329 ( .A(n1881), .B(n1880), .Z(n2155) );
  IV U2330 ( .A(n2155), .Z(n2153) );
  OR U2331 ( .A(n1884), .B(n1882), .Z(n1888) );
  ANDN U2332 ( .B(n1884), .A(n1883), .Z(n1886) );
  OR U2333 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2334 ( .A(n1888), .B(n1887), .Z(n2154) );
  NAND U2335 ( .A(n1890), .B(n1889), .Z(n1894) );
  NAND U2336 ( .A(n1892), .B(n1891), .Z(n1893) );
  AND U2337 ( .A(n1894), .B(n1893), .Z(n2150) );
  AND U2338 ( .A(x[80]), .B(y[195]), .Z(n2048) );
  AND U2339 ( .A(y[199]), .B(x[84]), .Z(n2424) );
  NAND U2340 ( .A(n2048), .B(n2424), .Z(n1898) );
  NANDN U2341 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2342 ( .A(n1898), .B(n1897), .Z(n2068) );
  AND U2343 ( .A(y[194]), .B(x[86]), .Z(n2085) );
  XOR U2344 ( .A(n2086), .B(n2085), .Z(n2088) );
  AND U2345 ( .A(y[214]), .B(x[66]), .Z(n2087) );
  XOR U2346 ( .A(n2088), .B(n2087), .Z(n2066) );
  AND U2347 ( .A(x[65]), .B(y[215]), .Z(n2093) );
  XOR U2348 ( .A(n2094), .B(n2093), .Z(n2092) );
  ANDN U2349 ( .B(o[23]), .A(n1899), .Z(n2091) );
  XOR U2350 ( .A(n2092), .B(n2091), .Z(n2065) );
  XOR U2351 ( .A(n2066), .B(n2065), .Z(n2067) );
  XNOR U2352 ( .A(n2068), .B(n2067), .Z(n2123) );
  NANDN U2353 ( .A(n1901), .B(n1900), .Z(n1905) );
  NANDN U2354 ( .A(n1903), .B(n1902), .Z(n1904) );
  AND U2355 ( .A(n1905), .B(n1904), .Z(n2062) );
  AND U2356 ( .A(x[85]), .B(y[195]), .Z(n1907) );
  NAND U2357 ( .A(y[200]), .B(x[80]), .Z(n1906) );
  XNOR U2358 ( .A(n1907), .B(n1906), .Z(n2049) );
  NAND U2359 ( .A(x[69]), .B(y[211]), .Z(n2050) );
  XNOR U2360 ( .A(n2049), .B(n2050), .Z(n2059) );
  AND U2361 ( .A(y[196]), .B(x[84]), .Z(n2259) );
  NAND U2362 ( .A(y[210]), .B(x[70]), .Z(n2438) );
  XNOR U2363 ( .A(n2259), .B(n2438), .Z(n2055) );
  NAND U2364 ( .A(x[83]), .B(y[197]), .Z(n2056) );
  XOR U2365 ( .A(n2055), .B(n2056), .Z(n2060) );
  XNOR U2366 ( .A(n2059), .B(n2060), .Z(n2061) );
  XNOR U2367 ( .A(n2062), .B(n2061), .Z(n2040) );
  NAND U2368 ( .A(n2186), .B(n1908), .Z(n1912) );
  NANDN U2369 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2370 ( .A(n1912), .B(n1911), .Z(n2039) );
  NANDN U2371 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2372 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2373 ( .A(n1918), .B(n1917), .Z(n2038) );
  XOR U2374 ( .A(n2039), .B(n2038), .Z(n2041) );
  XOR U2375 ( .A(n2040), .B(n2041), .Z(n2124) );
  XNOR U2376 ( .A(n2123), .B(n2124), .Z(n2125) );
  NANDN U2377 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U2378 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2379 ( .A(n1924), .B(n1923), .Z(n2118) );
  AND U2380 ( .A(y[213]), .B(x[67]), .Z(n2105) );
  XOR U2381 ( .A(n2106), .B(n2105), .Z(n2108) );
  NAND U2382 ( .A(x[68]), .B(y[212]), .Z(n2107) );
  XNOR U2383 ( .A(n2108), .B(n2107), .Z(n2117) );
  XNOR U2384 ( .A(n2118), .B(n2117), .Z(n2119) );
  AND U2385 ( .A(x[73]), .B(y[207]), .Z(n1926) );
  NAND U2386 ( .A(x[74]), .B(y[206]), .Z(n1925) );
  XNOR U2387 ( .A(n1926), .B(n1925), .Z(n2076) );
  AND U2388 ( .A(x[72]), .B(y[208]), .Z(n1928) );
  NAND U2389 ( .A(y[202]), .B(x[78]), .Z(n1927) );
  XNOR U2390 ( .A(n1928), .B(n1927), .Z(n2081) );
  NAND U2391 ( .A(y[205]), .B(x[75]), .Z(n2082) );
  XOR U2392 ( .A(n2081), .B(n2082), .Z(n2077) );
  XOR U2393 ( .A(n2076), .B(n2077), .Z(n2120) );
  XOR U2394 ( .A(n2119), .B(n2120), .Z(n2126) );
  XOR U2395 ( .A(n2125), .B(n2126), .Z(n2135) );
  NAND U2396 ( .A(n1930), .B(n1929), .Z(n1934) );
  NAND U2397 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2398 ( .A(n1934), .B(n1933), .Z(n2136) );
  XOR U2399 ( .A(n2135), .B(n2136), .Z(n2138) );
  NAND U2400 ( .A(n1936), .B(n1935), .Z(n1940) );
  NAND U2401 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U2402 ( .A(n1940), .B(n1939), .Z(n2137) );
  XOR U2403 ( .A(n2138), .B(n2137), .Z(n2144) );
  NANDN U2404 ( .A(n1942), .B(n1941), .Z(n1946) );
  NAND U2405 ( .A(n1944), .B(n1943), .Z(n1945) );
  AND U2406 ( .A(n1946), .B(n1945), .Z(n2132) );
  NANDN U2407 ( .A(n1948), .B(n1947), .Z(n1952) );
  NANDN U2408 ( .A(n1950), .B(n1949), .Z(n1951) );
  AND U2409 ( .A(n1952), .B(n1951), .Z(n2130) );
  NANDN U2410 ( .A(n1954), .B(n1953), .Z(n1958) );
  NAND U2411 ( .A(n1956), .B(n1955), .Z(n1957) );
  AND U2412 ( .A(n1958), .B(n1957), .Z(n2047) );
  AND U2413 ( .A(x[64]), .B(y[216]), .Z(n2111) );
  NAND U2414 ( .A(x[88]), .B(y[192]), .Z(n2112) );
  XNOR U2415 ( .A(n2111), .B(n2112), .Z(n2113) );
  NAND U2416 ( .A(x[87]), .B(y[193]), .Z(n2104) );
  XOR U2417 ( .A(o[24]), .B(n2104), .Z(n2114) );
  XNOR U2418 ( .A(n2113), .B(n2114), .Z(n2045) );
  AND U2419 ( .A(x[71]), .B(y[209]), .Z(n2098) );
  AND U2420 ( .A(x[82]), .B(y[198]), .Z(n2097) );
  XOR U2421 ( .A(n2098), .B(n2097), .Z(n2100) );
  AND U2422 ( .A(x[81]), .B(y[199]), .Z(n2099) );
  XOR U2423 ( .A(n2100), .B(n2099), .Z(n2044) );
  XOR U2424 ( .A(n2045), .B(n2044), .Z(n2046) );
  XNOR U2425 ( .A(n2047), .B(n2046), .Z(n2034) );
  NANDN U2426 ( .A(n1960), .B(n1959), .Z(n1964) );
  NANDN U2427 ( .A(n1962), .B(n1961), .Z(n1963) );
  AND U2428 ( .A(n1964), .B(n1963), .Z(n2033) );
  NANDN U2429 ( .A(n1966), .B(n1965), .Z(n1970) );
  NANDN U2430 ( .A(n1968), .B(n1967), .Z(n1969) );
  NAND U2431 ( .A(n1970), .B(n1969), .Z(n2032) );
  XOR U2432 ( .A(n2033), .B(n2032), .Z(n2035) );
  XNOR U2433 ( .A(n2034), .B(n2035), .Z(n2129) );
  XNOR U2434 ( .A(n2130), .B(n2129), .Z(n2131) );
  XOR U2435 ( .A(n2132), .B(n2131), .Z(n2028) );
  NAND U2436 ( .A(n1972), .B(n1971), .Z(n1976) );
  NANDN U2437 ( .A(n1974), .B(n1973), .Z(n1975) );
  AND U2438 ( .A(n1976), .B(n1975), .Z(n2072) );
  NAND U2439 ( .A(n1978), .B(n1977), .Z(n1982) );
  NAND U2440 ( .A(n1980), .B(n1979), .Z(n1981) );
  AND U2441 ( .A(n1982), .B(n1981), .Z(n2070) );
  NAND U2442 ( .A(n1984), .B(n1983), .Z(n1988) );
  NAND U2443 ( .A(n1986), .B(n1985), .Z(n1987) );
  AND U2444 ( .A(n1988), .B(n1987), .Z(n2069) );
  XOR U2445 ( .A(n2070), .B(n2069), .Z(n2071) );
  XOR U2446 ( .A(n2072), .B(n2071), .Z(n2027) );
  NAND U2447 ( .A(n1990), .B(n1989), .Z(n1994) );
  NAND U2448 ( .A(n1992), .B(n1991), .Z(n1993) );
  AND U2449 ( .A(n1994), .B(n1993), .Z(n2026) );
  XOR U2450 ( .A(n2027), .B(n2026), .Z(n2029) );
  XOR U2451 ( .A(n2028), .B(n2029), .Z(n2142) );
  NAND U2452 ( .A(n1996), .B(n1995), .Z(n2000) );
  NAND U2453 ( .A(n1998), .B(n1997), .Z(n1999) );
  AND U2454 ( .A(n2000), .B(n1999), .Z(n2141) );
  XOR U2455 ( .A(n2142), .B(n2141), .Z(n2143) );
  XOR U2456 ( .A(n2144), .B(n2143), .Z(n2148) );
  NAND U2457 ( .A(n2002), .B(n2001), .Z(n2006) );
  NANDN U2458 ( .A(n2004), .B(n2003), .Z(n2005) );
  NAND U2459 ( .A(n2006), .B(n2005), .Z(n2022) );
  NANDN U2460 ( .A(n2008), .B(n2007), .Z(n2012) );
  NANDN U2461 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U2462 ( .A(n2012), .B(n2011), .Z(n2021) );
  NAND U2463 ( .A(n2014), .B(n2013), .Z(n2018) );
  NANDN U2464 ( .A(n2016), .B(n2015), .Z(n2017) );
  NAND U2465 ( .A(n2018), .B(n2017), .Z(n2020) );
  XOR U2466 ( .A(n2021), .B(n2020), .Z(n2023) );
  XOR U2467 ( .A(n2022), .B(n2023), .Z(n2147) );
  XNOR U2468 ( .A(n2148), .B(n2147), .Z(n2149) );
  XOR U2469 ( .A(n2150), .B(n2149), .Z(n2156) );
  XNOR U2470 ( .A(n2154), .B(n2156), .Z(n2019) );
  XOR U2471 ( .A(n2153), .B(n2019), .Z(N57) );
  NAND U2472 ( .A(n2021), .B(n2020), .Z(n2025) );
  NAND U2473 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2474 ( .A(n2025), .B(n2024), .Z(n2305) );
  NAND U2475 ( .A(n2027), .B(n2026), .Z(n2031) );
  NAND U2476 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U2477 ( .A(n2031), .B(n2030), .Z(n2169) );
  NANDN U2478 ( .A(n2033), .B(n2032), .Z(n2037) );
  NANDN U2479 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U2480 ( .A(n2037), .B(n2036), .Z(n2174) );
  NANDN U2481 ( .A(n2039), .B(n2038), .Z(n2043) );
  NANDN U2482 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2483 ( .A(n2043), .B(n2042), .Z(n2173) );
  XNOR U2484 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2485 ( .A(y[200]), .B(x[85]), .Z(n3156) );
  NAND U2486 ( .A(n3156), .B(n2048), .Z(n2052) );
  NANDN U2487 ( .A(n2050), .B(n2049), .Z(n2051) );
  AND U2488 ( .A(n2052), .B(n2051), .Z(n2279) );
  AND U2489 ( .A(x[86]), .B(y[195]), .Z(n2248) );
  AND U2490 ( .A(x[69]), .B(y[212]), .Z(n2247) );
  NAND U2491 ( .A(x[81]), .B(y[200]), .Z(n2246) );
  XOR U2492 ( .A(n2247), .B(n2246), .Z(n2249) );
  XOR U2493 ( .A(n2248), .B(n2249), .Z(n2277) );
  AND U2494 ( .A(x[84]), .B(y[197]), .Z(n2054) );
  NAND U2495 ( .A(x[85]), .B(y[196]), .Z(n2053) );
  XNOR U2496 ( .A(n2054), .B(n2053), .Z(n2261) );
  AND U2497 ( .A(x[83]), .B(y[198]), .Z(n2260) );
  XOR U2498 ( .A(n2261), .B(n2260), .Z(n2276) );
  XNOR U2499 ( .A(n2277), .B(n2276), .Z(n2278) );
  XOR U2500 ( .A(n2279), .B(n2278), .Z(n2204) );
  NANDN U2501 ( .A(n2438), .B(n2259), .Z(n2058) );
  NANDN U2502 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U2503 ( .A(n2058), .B(n2057), .Z(n2284) );
  AND U2504 ( .A(x[79]), .B(y[202]), .Z(n2266) );
  AND U2505 ( .A(y[199]), .B(x[82]), .Z(n2265) );
  NAND U2506 ( .A(x[70]), .B(y[211]), .Z(n2264) );
  XOR U2507 ( .A(n2265), .B(n2264), .Z(n2267) );
  XOR U2508 ( .A(n2266), .B(n2267), .Z(n2283) );
  AND U2509 ( .A(x[87]), .B(y[194]), .Z(n2242) );
  AND U2510 ( .A(x[68]), .B(y[213]), .Z(n2241) );
  NAND U2511 ( .A(x[80]), .B(y[201]), .Z(n2240) );
  XOR U2512 ( .A(n2241), .B(n2240), .Z(n2243) );
  XNOR U2513 ( .A(n2242), .B(n2243), .Z(n2282) );
  XOR U2514 ( .A(n2283), .B(n2282), .Z(n2285) );
  XNOR U2515 ( .A(n2284), .B(n2285), .Z(n2203) );
  XOR U2516 ( .A(n2204), .B(n2203), .Z(n2205) );
  XOR U2517 ( .A(n2206), .B(n2205), .Z(n2218) );
  NANDN U2518 ( .A(n2060), .B(n2059), .Z(n2064) );
  NANDN U2519 ( .A(n2062), .B(n2061), .Z(n2063) );
  AND U2520 ( .A(n2064), .B(n2063), .Z(n2216) );
  XNOR U2521 ( .A(n2216), .B(n2215), .Z(n2217) );
  XOR U2522 ( .A(n2218), .B(n2217), .Z(n2176) );
  XOR U2523 ( .A(n2175), .B(n2176), .Z(n2168) );
  NAND U2524 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U2525 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U2526 ( .A(n2074), .B(n2073), .Z(n2167) );
  XOR U2527 ( .A(n2168), .B(n2167), .Z(n2170) );
  XOR U2528 ( .A(n2169), .B(n2170), .Z(n2164) );
  NANDN U2529 ( .A(n2185), .B(n2075), .Z(n2079) );
  NANDN U2530 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U2531 ( .A(n2079), .B(n2078), .Z(n2210) );
  AND U2532 ( .A(x[78]), .B(y[208]), .Z(n3060) );
  NAND U2533 ( .A(n3060), .B(n2080), .Z(n2084) );
  NANDN U2534 ( .A(n2082), .B(n2081), .Z(n2083) );
  AND U2535 ( .A(n2084), .B(n2083), .Z(n2237) );
  AND U2536 ( .A(x[75]), .B(y[206]), .Z(n2255) );
  AND U2537 ( .A(x[76]), .B(y[205]), .Z(n2254) );
  NAND U2538 ( .A(x[71]), .B(y[210]), .Z(n2253) );
  XOR U2539 ( .A(n2254), .B(n2253), .Z(n2256) );
  XOR U2540 ( .A(n2255), .B(n2256), .Z(n2235) );
  NAND U2541 ( .A(x[88]), .B(y[193]), .Z(n2252) );
  XNOR U2542 ( .A(o[25]), .B(n2252), .Z(n2222) );
  NAND U2543 ( .A(x[65]), .B(y[216]), .Z(n2223) );
  XNOR U2544 ( .A(n2222), .B(n2223), .Z(n2224) );
  NAND U2545 ( .A(y[204]), .B(x[77]), .Z(n2225) );
  XNOR U2546 ( .A(n2224), .B(n2225), .Z(n2234) );
  XNOR U2547 ( .A(n2235), .B(n2234), .Z(n2236) );
  XNOR U2548 ( .A(n2237), .B(n2236), .Z(n2209) );
  XNOR U2549 ( .A(n2210), .B(n2209), .Z(n2212) );
  AND U2550 ( .A(n2086), .B(n2085), .Z(n2090) );
  NAND U2551 ( .A(n2088), .B(n2087), .Z(n2089) );
  NANDN U2552 ( .A(n2090), .B(n2089), .Z(n2198) );
  AND U2553 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U2554 ( .A(n2094), .B(n2093), .Z(n2095) );
  NANDN U2555 ( .A(n2096), .B(n2095), .Z(n2197) );
  XOR U2556 ( .A(n2198), .B(n2197), .Z(n2199) );
  NAND U2557 ( .A(n2098), .B(n2097), .Z(n2102) );
  NAND U2558 ( .A(n2100), .B(n2099), .Z(n2101) );
  NAND U2559 ( .A(n2102), .B(n2101), .Z(n2193) );
  AND U2560 ( .A(x[72]), .B(y[209]), .Z(n2188) );
  XOR U2561 ( .A(n2186), .B(n2103), .Z(n2187) );
  XOR U2562 ( .A(n2188), .B(n2187), .Z(n2192) );
  ANDN U2563 ( .B(o[24]), .A(n2104), .Z(n2182) );
  AND U2564 ( .A(x[89]), .B(y[192]), .Z(n2180) );
  NAND U2565 ( .A(y[217]), .B(x[64]), .Z(n2179) );
  XNOR U2566 ( .A(n2180), .B(n2179), .Z(n2181) );
  XOR U2567 ( .A(n2182), .B(n2181), .Z(n2191) );
  XNOR U2568 ( .A(n2192), .B(n2191), .Z(n2194) );
  XNOR U2569 ( .A(n2199), .B(n2200), .Z(n2211) );
  XOR U2570 ( .A(n2212), .B(n2211), .Z(n2291) );
  NAND U2571 ( .A(n2106), .B(n2105), .Z(n2110) );
  ANDN U2572 ( .B(n2108), .A(n2107), .Z(n2109) );
  ANDN U2573 ( .B(n2110), .A(n2109), .Z(n2272) );
  NANDN U2574 ( .A(n2112), .B(n2111), .Z(n2116) );
  NANDN U2575 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U2576 ( .A(n2116), .B(n2115), .Z(n2271) );
  AND U2577 ( .A(x[78]), .B(y[203]), .Z(n2229) );
  AND U2578 ( .A(y[215]), .B(x[66]), .Z(n2228) );
  XOR U2579 ( .A(n2229), .B(n2228), .Z(n2231) );
  AND U2580 ( .A(x[67]), .B(y[214]), .Z(n2230) );
  XOR U2581 ( .A(n2231), .B(n2230), .Z(n2270) );
  XOR U2582 ( .A(n2271), .B(n2270), .Z(n2273) );
  XOR U2583 ( .A(n2272), .B(n2273), .Z(n2289) );
  NANDN U2584 ( .A(n2118), .B(n2117), .Z(n2122) );
  NANDN U2585 ( .A(n2120), .B(n2119), .Z(n2121) );
  AND U2586 ( .A(n2122), .B(n2121), .Z(n2288) );
  XNOR U2587 ( .A(n2289), .B(n2288), .Z(n2290) );
  XNOR U2588 ( .A(n2291), .B(n2290), .Z(n2294) );
  NANDN U2589 ( .A(n2124), .B(n2123), .Z(n2128) );
  NANDN U2590 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U2591 ( .A(n2128), .B(n2127), .Z(n2295) );
  XNOR U2592 ( .A(n2294), .B(n2295), .Z(n2296) );
  NANDN U2593 ( .A(n2130), .B(n2129), .Z(n2134) );
  NANDN U2594 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U2595 ( .A(n2134), .B(n2133), .Z(n2297) );
  XOR U2596 ( .A(n2296), .B(n2297), .Z(n2161) );
  NAND U2597 ( .A(n2136), .B(n2135), .Z(n2140) );
  NAND U2598 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U2599 ( .A(n2140), .B(n2139), .Z(n2162) );
  XOR U2600 ( .A(n2161), .B(n2162), .Z(n2163) );
  NAND U2601 ( .A(n2142), .B(n2141), .Z(n2146) );
  NAND U2602 ( .A(n2144), .B(n2143), .Z(n2145) );
  NAND U2603 ( .A(n2146), .B(n2145), .Z(n2303) );
  XNOR U2604 ( .A(n2305), .B(n2306), .Z(n2302) );
  NANDN U2605 ( .A(n2148), .B(n2147), .Z(n2152) );
  NAND U2606 ( .A(n2150), .B(n2149), .Z(n2151) );
  NAND U2607 ( .A(n2152), .B(n2151), .Z(n2301) );
  NANDN U2608 ( .A(n2153), .B(n2154), .Z(n2159) );
  NOR U2609 ( .A(n2155), .B(n2154), .Z(n2157) );
  OR U2610 ( .A(n2157), .B(n2156), .Z(n2158) );
  AND U2611 ( .A(n2159), .B(n2158), .Z(n2300) );
  XOR U2612 ( .A(n2301), .B(n2300), .Z(n2160) );
  XNOR U2613 ( .A(n2302), .B(n2160), .Z(N58) );
  NAND U2614 ( .A(n2162), .B(n2161), .Z(n2166) );
  NANDN U2615 ( .A(n2164), .B(n2163), .Z(n2165) );
  NAND U2616 ( .A(n2166), .B(n2165), .Z(n2456) );
  NAND U2617 ( .A(n2168), .B(n2167), .Z(n2172) );
  NAND U2618 ( .A(n2170), .B(n2169), .Z(n2171) );
  AND U2619 ( .A(n2172), .B(n2171), .Z(n2457) );
  XOR U2620 ( .A(n2456), .B(n2457), .Z(n2459) );
  NANDN U2621 ( .A(n2174), .B(n2173), .Z(n2178) );
  NANDN U2622 ( .A(n2176), .B(n2175), .Z(n2177) );
  AND U2623 ( .A(n2178), .B(n2177), .Z(n2453) );
  AND U2624 ( .A(x[66]), .B(y[216]), .Z(n2332) );
  XOR U2625 ( .A(n2333), .B(n2332), .Z(n2335) );
  NAND U2626 ( .A(y[194]), .B(x[88]), .Z(n2334) );
  XNOR U2627 ( .A(n2335), .B(n2334), .Z(n2374) );
  NANDN U2628 ( .A(n2180), .B(n2179), .Z(n2184) );
  NANDN U2629 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U2630 ( .A(n2184), .B(n2183), .Z(n2375) );
  XNOR U2631 ( .A(n2374), .B(n2375), .Z(n2376) );
  NANDN U2632 ( .A(n2186), .B(n2185), .Z(n2190) );
  NANDN U2633 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U2634 ( .A(n2190), .B(n2189), .Z(n2377) );
  XOR U2635 ( .A(n2376), .B(n2377), .Z(n2405) );
  NAND U2636 ( .A(n2192), .B(n2191), .Z(n2196) );
  NANDN U2637 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U2638 ( .A(n2196), .B(n2195), .Z(n2406) );
  XOR U2639 ( .A(n2405), .B(n2406), .Z(n2408) );
  NAND U2640 ( .A(n2198), .B(n2197), .Z(n2202) );
  NANDN U2641 ( .A(n2200), .B(n2199), .Z(n2201) );
  AND U2642 ( .A(n2202), .B(n2201), .Z(n2407) );
  XOR U2643 ( .A(n2408), .B(n2407), .Z(n2402) );
  NAND U2644 ( .A(n2204), .B(n2203), .Z(n2208) );
  NAND U2645 ( .A(n2206), .B(n2205), .Z(n2207) );
  AND U2646 ( .A(n2208), .B(n2207), .Z(n2400) );
  NANDN U2647 ( .A(n2210), .B(n2209), .Z(n2214) );
  NAND U2648 ( .A(n2212), .B(n2211), .Z(n2213) );
  AND U2649 ( .A(n2214), .B(n2213), .Z(n2399) );
  XNOR U2650 ( .A(n2400), .B(n2399), .Z(n2401) );
  XOR U2651 ( .A(n2402), .B(n2401), .Z(n2451) );
  NANDN U2652 ( .A(n2216), .B(n2215), .Z(n2220) );
  NANDN U2653 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U2654 ( .A(n2220), .B(n2219), .Z(n2319) );
  AND U2655 ( .A(x[76]), .B(y[206]), .Z(n2572) );
  AND U2656 ( .A(y[213]), .B(x[69]), .Z(n2388) );
  XOR U2657 ( .A(n2572), .B(n2388), .Z(n2390) );
  NAND U2658 ( .A(x[74]), .B(y[208]), .Z(n2389) );
  XNOR U2659 ( .A(n2390), .B(n2389), .Z(n2414) );
  AND U2660 ( .A(x[71]), .B(y[211]), .Z(n2412) );
  NAND U2661 ( .A(x[70]), .B(y[212]), .Z(n2221) );
  XNOR U2662 ( .A(n2659), .B(n2221), .Z(n2439) );
  NAND U2663 ( .A(x[73]), .B(y[209]), .Z(n2440) );
  XNOR U2664 ( .A(n2439), .B(n2440), .Z(n2411) );
  XOR U2665 ( .A(n2412), .B(n2411), .Z(n2413) );
  XOR U2666 ( .A(n2414), .B(n2413), .Z(n2358) );
  NANDN U2667 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U2668 ( .A(n2225), .B(n2224), .Z(n2226) );
  NAND U2669 ( .A(n2227), .B(n2226), .Z(n2357) );
  NAND U2670 ( .A(n2229), .B(n2228), .Z(n2233) );
  NAND U2671 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U2672 ( .A(n2233), .B(n2232), .Z(n2356) );
  XNOR U2673 ( .A(n2357), .B(n2356), .Z(n2359) );
  NANDN U2674 ( .A(n2235), .B(n2234), .Z(n2239) );
  NANDN U2675 ( .A(n2237), .B(n2236), .Z(n2238) );
  AND U2676 ( .A(n2239), .B(n2238), .Z(n2362) );
  NANDN U2677 ( .A(n2241), .B(n2240), .Z(n2245) );
  OR U2678 ( .A(n2243), .B(n2242), .Z(n2244) );
  AND U2679 ( .A(n2245), .B(n2244), .Z(n2322) );
  NANDN U2680 ( .A(n2247), .B(n2246), .Z(n2251) );
  OR U2681 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2682 ( .A(n2251), .B(n2250), .Z(n2323) );
  XNOR U2683 ( .A(n2322), .B(n2323), .Z(n2324) );
  ANDN U2684 ( .B(o[25]), .A(n2252), .Z(n2431) );
  NAND U2685 ( .A(x[78]), .B(y[204]), .Z(n2432) );
  XNOR U2686 ( .A(n2431), .B(n2432), .Z(n2433) );
  NAND U2687 ( .A(x[65]), .B(y[217]), .Z(n2434) );
  XNOR U2688 ( .A(n2433), .B(n2434), .Z(n2380) );
  NAND U2689 ( .A(y[193]), .B(x[89]), .Z(n2443) );
  XNOR U2690 ( .A(o[26]), .B(n2443), .Z(n2393) );
  NAND U2691 ( .A(x[90]), .B(y[192]), .Z(n2394) );
  XNOR U2692 ( .A(n2393), .B(n2394), .Z(n2395) );
  NAND U2693 ( .A(x[64]), .B(y[218]), .Z(n2396) );
  XOR U2694 ( .A(n2395), .B(n2396), .Z(n2381) );
  XNOR U2695 ( .A(n2380), .B(n2381), .Z(n2382) );
  NANDN U2696 ( .A(n2254), .B(n2253), .Z(n2258) );
  OR U2697 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U2698 ( .A(n2258), .B(n2257), .Z(n2383) );
  XOR U2699 ( .A(n2382), .B(n2383), .Z(n2325) );
  XOR U2700 ( .A(n2324), .B(n2325), .Z(n2370) );
  AND U2701 ( .A(x[85]), .B(y[197]), .Z(n2425) );
  NAND U2702 ( .A(n2425), .B(n2259), .Z(n2263) );
  NAND U2703 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U2704 ( .A(n2263), .B(n2262), .Z(n2352) );
  XOR U2705 ( .A(n2426), .B(n2425), .Z(n2428) );
  NAND U2706 ( .A(y[198]), .B(x[84]), .Z(n2427) );
  XNOR U2707 ( .A(n2428), .B(n2427), .Z(n2351) );
  NAND U2708 ( .A(x[87]), .B(y[195]), .Z(n2339) );
  XNOR U2709 ( .A(n2338), .B(n2339), .Z(n2341) );
  AND U2710 ( .A(x[86]), .B(y[196]), .Z(n2340) );
  XOR U2711 ( .A(n2341), .B(n2340), .Z(n2350) );
  XOR U2712 ( .A(n2351), .B(n2350), .Z(n2353) );
  XOR U2713 ( .A(n2352), .B(n2353), .Z(n2369) );
  AND U2714 ( .A(x[67]), .B(y[215]), .Z(n2417) );
  NAND U2715 ( .A(x[75]), .B(y[207]), .Z(n2418) );
  XNOR U2716 ( .A(n2417), .B(n2418), .Z(n2419) );
  NAND U2717 ( .A(x[83]), .B(y[199]), .Z(n2420) );
  XNOR U2718 ( .A(n2419), .B(n2420), .Z(n2329) );
  NAND U2719 ( .A(x[68]), .B(y[214]), .Z(n2345) );
  XNOR U2720 ( .A(n2344), .B(n2345), .Z(n2346) );
  XOR U2721 ( .A(n2329), .B(n2328), .Z(n2331) );
  NANDN U2722 ( .A(n2265), .B(n2264), .Z(n2269) );
  OR U2723 ( .A(n2267), .B(n2266), .Z(n2268) );
  AND U2724 ( .A(n2269), .B(n2268), .Z(n2330) );
  XNOR U2725 ( .A(n2331), .B(n2330), .Z(n2368) );
  XOR U2726 ( .A(n2370), .B(n2371), .Z(n2364) );
  XOR U2727 ( .A(n2365), .B(n2364), .Z(n2317) );
  NANDN U2728 ( .A(n2271), .B(n2270), .Z(n2275) );
  OR U2729 ( .A(n2273), .B(n2272), .Z(n2274) );
  NAND U2730 ( .A(n2275), .B(n2274), .Z(n2446) );
  NANDN U2731 ( .A(n2277), .B(n2276), .Z(n2281) );
  NANDN U2732 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U2733 ( .A(n2281), .B(n2280), .Z(n2445) );
  NANDN U2734 ( .A(n2283), .B(n2282), .Z(n2287) );
  OR U2735 ( .A(n2285), .B(n2284), .Z(n2286) );
  NAND U2736 ( .A(n2287), .B(n2286), .Z(n2444) );
  XOR U2737 ( .A(n2445), .B(n2444), .Z(n2447) );
  XOR U2738 ( .A(n2446), .B(n2447), .Z(n2316) );
  XNOR U2739 ( .A(n2317), .B(n2316), .Z(n2318) );
  XNOR U2740 ( .A(n2319), .B(n2318), .Z(n2450) );
  XNOR U2741 ( .A(n2451), .B(n2450), .Z(n2452) );
  XNOR U2742 ( .A(n2453), .B(n2452), .Z(n2312) );
  NANDN U2743 ( .A(n2289), .B(n2288), .Z(n2293) );
  NANDN U2744 ( .A(n2291), .B(n2290), .Z(n2292) );
  AND U2745 ( .A(n2293), .B(n2292), .Z(n2310) );
  NANDN U2746 ( .A(n2295), .B(n2294), .Z(n2299) );
  NANDN U2747 ( .A(n2297), .B(n2296), .Z(n2298) );
  NAND U2748 ( .A(n2299), .B(n2298), .Z(n2311) );
  XOR U2749 ( .A(n2310), .B(n2311), .Z(n2313) );
  XNOR U2750 ( .A(n2312), .B(n2313), .Z(n2458) );
  XNOR U2751 ( .A(n2459), .B(n2458), .Z(n2465) );
  NANDN U2752 ( .A(n2304), .B(n2303), .Z(n2308) );
  NANDN U2753 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2754 ( .A(n2308), .B(n2307), .Z(n2463) );
  IV U2755 ( .A(n2463), .Z(n2462) );
  XOR U2756 ( .A(n2464), .B(n2462), .Z(n2309) );
  XNOR U2757 ( .A(n2465), .B(n2309), .Z(N59) );
  NANDN U2758 ( .A(n2311), .B(n2310), .Z(n2315) );
  NANDN U2759 ( .A(n2313), .B(n2312), .Z(n2314) );
  AND U2760 ( .A(n2315), .B(n2314), .Z(n2622) );
  NANDN U2761 ( .A(n2317), .B(n2316), .Z(n2321) );
  NANDN U2762 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2763 ( .A(n2321), .B(n2320), .Z(n2472) );
  NANDN U2764 ( .A(n2323), .B(n2322), .Z(n2327) );
  NANDN U2765 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2766 ( .A(n2327), .B(n2326), .Z(n2497) );
  NAND U2767 ( .A(n2333), .B(n2332), .Z(n2337) );
  ANDN U2768 ( .B(n2335), .A(n2334), .Z(n2336) );
  ANDN U2769 ( .B(n2337), .A(n2336), .Z(n2549) );
  NANDN U2770 ( .A(n2339), .B(n2338), .Z(n2343) );
  NAND U2771 ( .A(n2341), .B(n2340), .Z(n2342) );
  NAND U2772 ( .A(n2343), .B(n2342), .Z(n2548) );
  XNOR U2773 ( .A(n2549), .B(n2548), .Z(n2550) );
  NANDN U2774 ( .A(n2345), .B(n2344), .Z(n2349) );
  NANDN U2775 ( .A(n2347), .B(n2346), .Z(n2348) );
  AND U2776 ( .A(n2349), .B(n2348), .Z(n2563) );
  AND U2777 ( .A(x[64]), .B(y[219]), .Z(n2517) );
  NAND U2778 ( .A(y[192]), .B(x[91]), .Z(n2518) );
  XNOR U2779 ( .A(n2517), .B(n2518), .Z(n2519) );
  AND U2780 ( .A(y[193]), .B(x[90]), .Z(n2523) );
  XOR U2781 ( .A(o[27]), .B(n2523), .Z(n2520) );
  XOR U2782 ( .A(n2519), .B(n2520), .Z(n2560) );
  AND U2783 ( .A(y[210]), .B(x[73]), .Z(n2526) );
  NAND U2784 ( .A(x[85]), .B(y[198]), .Z(n2527) );
  XNOR U2785 ( .A(n2526), .B(n2527), .Z(n2528) );
  NAND U2786 ( .A(y[201]), .B(x[82]), .Z(n2529) );
  XOR U2787 ( .A(n2528), .B(n2529), .Z(n2561) );
  XNOR U2788 ( .A(n2560), .B(n2561), .Z(n2562) );
  XOR U2789 ( .A(n2563), .B(n2562), .Z(n2551) );
  XNOR U2790 ( .A(n2550), .B(n2551), .Z(n2494) );
  XNOR U2791 ( .A(n2495), .B(n2494), .Z(n2496) );
  XOR U2792 ( .A(n2497), .B(n2496), .Z(n2615) );
  NAND U2793 ( .A(n2351), .B(n2350), .Z(n2355) );
  NAND U2794 ( .A(n2353), .B(n2352), .Z(n2354) );
  AND U2795 ( .A(n2355), .B(n2354), .Z(n2614) );
  NAND U2796 ( .A(n2357), .B(n2356), .Z(n2361) );
  NANDN U2797 ( .A(n2359), .B(n2358), .Z(n2360) );
  AND U2798 ( .A(n2361), .B(n2360), .Z(n2613) );
  XOR U2799 ( .A(n2614), .B(n2613), .Z(n2616) );
  XOR U2800 ( .A(n2615), .B(n2616), .Z(n2471) );
  NANDN U2801 ( .A(n2363), .B(n2362), .Z(n2367) );
  NAND U2802 ( .A(n2365), .B(n2364), .Z(n2366) );
  AND U2803 ( .A(n2367), .B(n2366), .Z(n2604) );
  NANDN U2804 ( .A(n2369), .B(n2368), .Z(n2373) );
  NAND U2805 ( .A(n2371), .B(n2370), .Z(n2372) );
  AND U2806 ( .A(n2373), .B(n2372), .Z(n2602) );
  NANDN U2807 ( .A(n2375), .B(n2374), .Z(n2379) );
  NANDN U2808 ( .A(n2377), .B(n2376), .Z(n2378) );
  AND U2809 ( .A(n2379), .B(n2378), .Z(n2491) );
  NANDN U2810 ( .A(n2381), .B(n2380), .Z(n2385) );
  NANDN U2811 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U2812 ( .A(n2385), .B(n2384), .Z(n2489) );
  AND U2813 ( .A(y[200]), .B(x[83]), .Z(n2505) );
  NAND U2814 ( .A(y[194]), .B(x[89]), .Z(n2506) );
  XNOR U2815 ( .A(n2505), .B(n2506), .Z(n2507) );
  NAND U2816 ( .A(y[213]), .B(x[70]), .Z(n2508) );
  XNOR U2817 ( .A(n2507), .B(n2508), .Z(n2542) );
  AND U2818 ( .A(y[204]), .B(x[79]), .Z(n2583) );
  NAND U2819 ( .A(y[217]), .B(x[66]), .Z(n2584) );
  XNOR U2820 ( .A(n2583), .B(n2584), .Z(n2585) );
  NAND U2821 ( .A(x[67]), .B(y[216]), .Z(n2586) );
  XOR U2822 ( .A(n2585), .B(n2586), .Z(n2543) );
  XNOR U2823 ( .A(n2542), .B(n2543), .Z(n2544) );
  AND U2824 ( .A(x[80]), .B(y[203]), .Z(n2596) );
  XOR U2825 ( .A(n2596), .B(n2595), .Z(n2597) );
  XOR U2826 ( .A(n2598), .B(n2597), .Z(n2574) );
  AND U2827 ( .A(x[77]), .B(y[206]), .Z(n2387) );
  NAND U2828 ( .A(y[207]), .B(x[76]), .Z(n2386) );
  XNOR U2829 ( .A(n2387), .B(n2386), .Z(n2573) );
  XOR U2830 ( .A(n2574), .B(n2573), .Z(n2545) );
  XOR U2831 ( .A(n2544), .B(n2545), .Z(n2568) );
  NAND U2832 ( .A(n2572), .B(n2388), .Z(n2392) );
  ANDN U2833 ( .B(n2390), .A(n2389), .Z(n2391) );
  ANDN U2834 ( .B(n2392), .A(n2391), .Z(n2567) );
  NANDN U2835 ( .A(n2394), .B(n2393), .Z(n2398) );
  NANDN U2836 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U2837 ( .A(n2398), .B(n2397), .Z(n2566) );
  XOR U2838 ( .A(n2567), .B(n2566), .Z(n2569) );
  XNOR U2839 ( .A(n2568), .B(n2569), .Z(n2488) );
  XNOR U2840 ( .A(n2489), .B(n2488), .Z(n2490) );
  XNOR U2841 ( .A(n2491), .B(n2490), .Z(n2601) );
  XOR U2842 ( .A(n2602), .B(n2601), .Z(n2603) );
  XOR U2843 ( .A(n2604), .B(n2603), .Z(n2470) );
  XNOR U2844 ( .A(n2472), .B(n2473), .Z(n2478) );
  NANDN U2845 ( .A(n2400), .B(n2399), .Z(n2404) );
  NAND U2846 ( .A(n2402), .B(n2401), .Z(n2403) );
  NAND U2847 ( .A(n2404), .B(n2403), .Z(n2476) );
  NAND U2848 ( .A(n2406), .B(n2405), .Z(n2410) );
  NAND U2849 ( .A(n2408), .B(n2407), .Z(n2409) );
  NAND U2850 ( .A(n2410), .B(n2409), .Z(n2482) );
  NAND U2851 ( .A(n2412), .B(n2411), .Z(n2416) );
  NAND U2852 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U2853 ( .A(n2416), .B(n2415), .Z(n2609) );
  NANDN U2854 ( .A(n2418), .B(n2417), .Z(n2422) );
  NANDN U2855 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U2856 ( .A(n2422), .B(n2421), .Z(n2539) );
  NAND U2857 ( .A(x[88]), .B(y[195]), .Z(n2423) );
  XNOR U2858 ( .A(n2424), .B(n2423), .Z(n2501) );
  NAND U2859 ( .A(y[212]), .B(x[71]), .Z(n2502) );
  XNOR U2860 ( .A(n2501), .B(n2502), .Z(n2536) );
  AND U2861 ( .A(y[211]), .B(x[72]), .Z(n2589) );
  NAND U2862 ( .A(x[87]), .B(y[196]), .Z(n2590) );
  XNOR U2863 ( .A(n2589), .B(n2590), .Z(n2591) );
  NAND U2864 ( .A(x[86]), .B(y[197]), .Z(n2592) );
  XOR U2865 ( .A(n2591), .B(n2592), .Z(n2537) );
  XNOR U2866 ( .A(n2536), .B(n2537), .Z(n2538) );
  XOR U2867 ( .A(n2539), .B(n2538), .Z(n2607) );
  NAND U2868 ( .A(n2426), .B(n2425), .Z(n2430) );
  ANDN U2869 ( .B(n2428), .A(n2427), .Z(n2429) );
  ANDN U2870 ( .B(n2430), .A(n2429), .Z(n2533) );
  NANDN U2871 ( .A(n2432), .B(n2431), .Z(n2436) );
  NANDN U2872 ( .A(n2434), .B(n2433), .Z(n2435) );
  NAND U2873 ( .A(n2436), .B(n2435), .Z(n2532) );
  XNOR U2874 ( .A(n2533), .B(n2532), .Z(n2535) );
  AND U2875 ( .A(y[212]), .B(x[72]), .Z(n2437) );
  NANDN U2876 ( .A(n2438), .B(n2437), .Z(n2442) );
  NANDN U2877 ( .A(n2440), .B(n2439), .Z(n2441) );
  NAND U2878 ( .A(n2442), .B(n2441), .Z(n2556) );
  ANDN U2879 ( .B(o[26]), .A(n2443), .Z(n2579) );
  AND U2880 ( .A(x[78]), .B(y[205]), .Z(n2577) );
  NAND U2881 ( .A(x[65]), .B(y[218]), .Z(n2578) );
  XOR U2882 ( .A(n2577), .B(n2578), .Z(n2580) );
  XNOR U2883 ( .A(n2579), .B(n2580), .Z(n2555) );
  AND U2884 ( .A(x[81]), .B(y[202]), .Z(n2511) );
  NAND U2885 ( .A(x[68]), .B(y[215]), .Z(n2512) );
  XNOR U2886 ( .A(n2511), .B(n2512), .Z(n2514) );
  AND U2887 ( .A(x[69]), .B(y[214]), .Z(n2513) );
  XOR U2888 ( .A(n2514), .B(n2513), .Z(n2554) );
  XOR U2889 ( .A(n2555), .B(n2554), .Z(n2557) );
  XOR U2890 ( .A(n2556), .B(n2557), .Z(n2534) );
  XOR U2891 ( .A(n2535), .B(n2534), .Z(n2608) );
  XNOR U2892 ( .A(n2609), .B(n2610), .Z(n2483) );
  XOR U2893 ( .A(n2482), .B(n2483), .Z(n2485) );
  NAND U2894 ( .A(n2445), .B(n2444), .Z(n2449) );
  NAND U2895 ( .A(n2447), .B(n2446), .Z(n2448) );
  AND U2896 ( .A(n2449), .B(n2448), .Z(n2484) );
  XOR U2897 ( .A(n2485), .B(n2484), .Z(n2477) );
  XNOR U2898 ( .A(n2476), .B(n2477), .Z(n2479) );
  NANDN U2899 ( .A(n2451), .B(n2450), .Z(n2455) );
  NANDN U2900 ( .A(n2453), .B(n2452), .Z(n2454) );
  NAND U2901 ( .A(n2455), .B(n2454), .Z(n2619) );
  XOR U2902 ( .A(n2620), .B(n2619), .Z(n2621) );
  XNOR U2903 ( .A(n2622), .B(n2621), .Z(n2627) );
  NAND U2904 ( .A(n2457), .B(n2456), .Z(n2461) );
  NAND U2905 ( .A(n2459), .B(n2458), .Z(n2460) );
  AND U2906 ( .A(n2461), .B(n2460), .Z(n2626) );
  OR U2907 ( .A(n2464), .B(n2462), .Z(n2468) );
  ANDN U2908 ( .B(n2464), .A(n2463), .Z(n2466) );
  OR U2909 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2910 ( .A(n2468), .B(n2467), .Z(n2625) );
  XNOR U2911 ( .A(n2626), .B(n2625), .Z(n2469) );
  XNOR U2912 ( .A(n2627), .B(n2469), .Z(N60) );
  NANDN U2913 ( .A(n2471), .B(n2470), .Z(n2475) );
  NAND U2914 ( .A(n2473), .B(n2472), .Z(n2474) );
  NAND U2915 ( .A(n2475), .B(n2474), .Z(n2787) );
  NAND U2916 ( .A(n2477), .B(n2476), .Z(n2481) );
  NANDN U2917 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2918 ( .A(n2481), .B(n2480), .Z(n2788) );
  XOR U2919 ( .A(n2787), .B(n2788), .Z(n2790) );
  NAND U2920 ( .A(n2483), .B(n2482), .Z(n2487) );
  NAND U2921 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2922 ( .A(n2487), .B(n2486), .Z(n2630) );
  NANDN U2923 ( .A(n2489), .B(n2488), .Z(n2493) );
  NANDN U2924 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2925 ( .A(n2493), .B(n2492), .Z(n2776) );
  NANDN U2926 ( .A(n2495), .B(n2494), .Z(n2499) );
  NANDN U2927 ( .A(n2497), .B(n2496), .Z(n2498) );
  NAND U2928 ( .A(n2499), .B(n2498), .Z(n2775) );
  XNOR U2929 ( .A(n2776), .B(n2775), .Z(n2778) );
  AND U2930 ( .A(x[88]), .B(y[199]), .Z(n3162) );
  NAND U2931 ( .A(n2500), .B(n3162), .Z(n2504) );
  NANDN U2932 ( .A(n2502), .B(n2501), .Z(n2503) );
  AND U2933 ( .A(n2504), .B(n2503), .Z(n2759) );
  AND U2934 ( .A(y[195]), .B(x[89]), .Z(n2696) );
  XOR U2935 ( .A(n2697), .B(n2696), .Z(n2695) );
  NAND U2936 ( .A(x[65]), .B(y[219]), .Z(n2694) );
  XNOR U2937 ( .A(n2695), .B(n2694), .Z(n2757) );
  AND U2938 ( .A(x[80]), .B(y[204]), .Z(n2688) );
  NAND U2939 ( .A(x[88]), .B(y[196]), .Z(n2689) );
  XNOR U2940 ( .A(n2688), .B(n2689), .Z(n2690) );
  NAND U2941 ( .A(y[218]), .B(x[66]), .Z(n2691) );
  XOR U2942 ( .A(n2690), .B(n2691), .Z(n2758) );
  XOR U2943 ( .A(n2757), .B(n2758), .Z(n2760) );
  XOR U2944 ( .A(n2759), .B(n2760), .Z(n2742) );
  NANDN U2945 ( .A(n2506), .B(n2505), .Z(n2510) );
  NANDN U2946 ( .A(n2508), .B(n2507), .Z(n2509) );
  AND U2947 ( .A(n2510), .B(n2509), .Z(n2765) );
  NAND U2948 ( .A(y[217]), .B(x[67]), .Z(n2713) );
  XNOR U2949 ( .A(n2712), .B(n2713), .Z(n2714) );
  NAND U2950 ( .A(x[87]), .B(y[197]), .Z(n2715) );
  XNOR U2951 ( .A(n2714), .B(n2715), .Z(n2763) );
  AND U2952 ( .A(x[69]), .B(y[215]), .Z(n2681) );
  NAND U2953 ( .A(y[199]), .B(x[85]), .Z(n2682) );
  XNOR U2954 ( .A(n2681), .B(n2682), .Z(n2683) );
  NAND U2955 ( .A(y[200]), .B(x[84]), .Z(n2684) );
  XOR U2956 ( .A(n2683), .B(n2684), .Z(n2764) );
  XOR U2957 ( .A(n2763), .B(n2764), .Z(n2766) );
  XOR U2958 ( .A(n2765), .B(n2766), .Z(n2740) );
  NANDN U2959 ( .A(n2512), .B(n2511), .Z(n2516) );
  NAND U2960 ( .A(n2514), .B(n2513), .Z(n2515) );
  AND U2961 ( .A(n2516), .B(n2515), .Z(n2752) );
  NANDN U2962 ( .A(n2518), .B(n2517), .Z(n2522) );
  NAND U2963 ( .A(n2520), .B(n2519), .Z(n2521) );
  NAND U2964 ( .A(n2522), .B(n2521), .Z(n2751) );
  XNOR U2965 ( .A(n2752), .B(n2751), .Z(n2754) );
  AND U2966 ( .A(n2523), .B(o[27]), .Z(n2656) );
  AND U2967 ( .A(x[64]), .B(y[220]), .Z(n2654) );
  AND U2968 ( .A(y[192]), .B(x[92]), .Z(n2653) );
  XOR U2969 ( .A(n2654), .B(n2653), .Z(n2655) );
  XOR U2970 ( .A(n2656), .B(n2655), .Z(n2642) );
  AND U2971 ( .A(x[74]), .B(y[210]), .Z(n2525) );
  NAND U2972 ( .A(x[72]), .B(y[212]), .Z(n2524) );
  XNOR U2973 ( .A(n2525), .B(n2524), .Z(n2661) );
  AND U2974 ( .A(y[211]), .B(x[73]), .Z(n2660) );
  XOR U2975 ( .A(n2661), .B(n2660), .Z(n2641) );
  XOR U2976 ( .A(n2642), .B(n2641), .Z(n2644) );
  NANDN U2977 ( .A(n2527), .B(n2526), .Z(n2531) );
  NANDN U2978 ( .A(n2529), .B(n2528), .Z(n2530) );
  NAND U2979 ( .A(n2531), .B(n2530), .Z(n2643) );
  XOR U2980 ( .A(n2644), .B(n2643), .Z(n2753) );
  XNOR U2981 ( .A(n2754), .B(n2753), .Z(n2739) );
  XNOR U2982 ( .A(n2740), .B(n2739), .Z(n2741) );
  XOR U2983 ( .A(n2742), .B(n2741), .Z(n2781) );
  NANDN U2984 ( .A(n2537), .B(n2536), .Z(n2541) );
  NANDN U2985 ( .A(n2539), .B(n2538), .Z(n2540) );
  AND U2986 ( .A(n2541), .B(n2540), .Z(n2734) );
  NANDN U2987 ( .A(n2543), .B(n2542), .Z(n2547) );
  NAND U2988 ( .A(n2545), .B(n2544), .Z(n2546) );
  NAND U2989 ( .A(n2547), .B(n2546), .Z(n2733) );
  XNOR U2990 ( .A(n2734), .B(n2733), .Z(n2735) );
  XNOR U2991 ( .A(n2736), .B(n2735), .Z(n2782) );
  XOR U2992 ( .A(n2781), .B(n2782), .Z(n2784) );
  NANDN U2993 ( .A(n2549), .B(n2548), .Z(n2553) );
  NANDN U2994 ( .A(n2551), .B(n2550), .Z(n2552) );
  AND U2995 ( .A(n2553), .B(n2552), .Z(n2747) );
  NAND U2996 ( .A(n2555), .B(n2554), .Z(n2559) );
  NAND U2997 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U2998 ( .A(n2559), .B(n2558), .Z(n2746) );
  NANDN U2999 ( .A(n2561), .B(n2560), .Z(n2565) );
  NANDN U3000 ( .A(n2563), .B(n2562), .Z(n2564) );
  NAND U3001 ( .A(n2565), .B(n2564), .Z(n2745) );
  XOR U3002 ( .A(n2746), .B(n2745), .Z(n2748) );
  XOR U3003 ( .A(n2747), .B(n2748), .Z(n2728) );
  NANDN U3004 ( .A(n2567), .B(n2566), .Z(n2571) );
  NANDN U3005 ( .A(n2569), .B(n2568), .Z(n2570) );
  AND U3006 ( .A(n2571), .B(n2570), .Z(n2727) );
  XNOR U3007 ( .A(n2728), .B(n2727), .Z(n2729) );
  NAND U3008 ( .A(n2572), .B(n2712), .Z(n2576) );
  NAND U3009 ( .A(n2574), .B(n2573), .Z(n2575) );
  AND U3010 ( .A(n2576), .B(n2575), .Z(n2666) );
  NANDN U3011 ( .A(n2578), .B(n2577), .Z(n2582) );
  NANDN U3012 ( .A(n2580), .B(n2579), .Z(n2581) );
  AND U3013 ( .A(n2582), .B(n2581), .Z(n2665) );
  NANDN U3014 ( .A(n2584), .B(n2583), .Z(n2588) );
  NANDN U3015 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U3016 ( .A(n2588), .B(n2587), .Z(n2664) );
  XOR U3017 ( .A(n2665), .B(n2664), .Z(n2667) );
  XOR U3018 ( .A(n2666), .B(n2667), .Z(n2772) );
  AND U3019 ( .A(x[81]), .B(y[203]), .Z(n2648) );
  AND U3020 ( .A(x[86]), .B(y[198]), .Z(n2647) );
  XOR U3021 ( .A(n2648), .B(n2647), .Z(n2650) );
  AND U3022 ( .A(x[68]), .B(y[216]), .Z(n2649) );
  XOR U3023 ( .A(n2650), .B(n2649), .Z(n2670) );
  AND U3024 ( .A(y[214]), .B(x[70]), .Z(n2878) );
  NAND U3025 ( .A(y[201]), .B(x[83]), .Z(n2676) );
  XNOR U3026 ( .A(n2878), .B(n2676), .Z(n2677) );
  XOR U3027 ( .A(n2670), .B(n2671), .Z(n2673) );
  NANDN U3028 ( .A(n2590), .B(n2589), .Z(n2594) );
  NANDN U3029 ( .A(n2592), .B(n2591), .Z(n2593) );
  NAND U3030 ( .A(n2594), .B(n2593), .Z(n2672) );
  XOR U3031 ( .A(n2673), .B(n2672), .Z(n2770) );
  AND U3032 ( .A(y[213]), .B(x[71]), .Z(n2701) );
  AND U3033 ( .A(x[76]), .B(y[208]), .Z(n2700) );
  XOR U3034 ( .A(n2701), .B(n2700), .Z(n2703) );
  AND U3035 ( .A(x[75]), .B(y[209]), .Z(n2702) );
  XOR U3036 ( .A(n2703), .B(n2702), .Z(n2707) );
  AND U3037 ( .A(y[205]), .B(x[79]), .Z(n2721) );
  AND U3038 ( .A(y[193]), .B(x[91]), .Z(n2687) );
  XOR U3039 ( .A(o[28]), .B(n2687), .Z(n2719) );
  AND U3040 ( .A(y[194]), .B(x[90]), .Z(n2718) );
  XOR U3041 ( .A(n2719), .B(n2718), .Z(n2720) );
  XNOR U3042 ( .A(n2721), .B(n2720), .Z(n2706) );
  XNOR U3043 ( .A(n2707), .B(n2706), .Z(n2708) );
  OR U3044 ( .A(n2596), .B(n2595), .Z(n2600) );
  NANDN U3045 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U3046 ( .A(n2600), .B(n2599), .Z(n2709) );
  XNOR U3047 ( .A(n2708), .B(n2709), .Z(n2769) );
  XNOR U3048 ( .A(n2770), .B(n2769), .Z(n2771) );
  XOR U3049 ( .A(n2772), .B(n2771), .Z(n2730) );
  XOR U3050 ( .A(n2729), .B(n2730), .Z(n2783) );
  XOR U3051 ( .A(n2784), .B(n2783), .Z(n2777) );
  XOR U3052 ( .A(n2778), .B(n2777), .Z(n2629) );
  XOR U3053 ( .A(n2630), .B(n2629), .Z(n2631) );
  NAND U3054 ( .A(n2602), .B(n2601), .Z(n2606) );
  NAND U3055 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U3056 ( .A(n2606), .B(n2605), .Z(n2637) );
  NANDN U3057 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U3058 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U3059 ( .A(n2612), .B(n2611), .Z(n2636) );
  NAND U3060 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U3061 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U3062 ( .A(n2618), .B(n2617), .Z(n2635) );
  XOR U3063 ( .A(n2636), .B(n2635), .Z(n2638) );
  XNOR U3064 ( .A(n2637), .B(n2638), .Z(n2632) );
  XNOR U3065 ( .A(n2790), .B(n2789), .Z(n2795) );
  NAND U3066 ( .A(n2620), .B(n2619), .Z(n2624) );
  NANDN U3067 ( .A(n2622), .B(n2621), .Z(n2623) );
  NAND U3068 ( .A(n2624), .B(n2623), .Z(n2793) );
  XOR U3069 ( .A(n2793), .B(n2794), .Z(n2628) );
  XNOR U3070 ( .A(n2795), .B(n2628), .Z(N61) );
  NAND U3071 ( .A(n2630), .B(n2629), .Z(n2634) );
  NANDN U3072 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U3073 ( .A(n2634), .B(n2633), .Z(n2802) );
  NAND U3074 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U3075 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U3076 ( .A(n2640), .B(n2639), .Z(n2800) );
  NAND U3077 ( .A(n2642), .B(n2641), .Z(n2646) );
  NAND U3078 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U3079 ( .A(n2646), .B(n2645), .Z(n2909) );
  NAND U3080 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U3081 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U3082 ( .A(n2652), .B(n2651), .Z(n2946) );
  NAND U3083 ( .A(n2654), .B(n2653), .Z(n2658) );
  NAND U3084 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U3085 ( .A(n2658), .B(n2657), .Z(n2945) );
  XOR U3086 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U3087 ( .A(x[74]), .B(y[212]), .Z(n2944) );
  NAND U3088 ( .A(n2659), .B(n2944), .Z(n2663) );
  NAND U3089 ( .A(n2661), .B(n2660), .Z(n2662) );
  NAND U3090 ( .A(n2663), .B(n2662), .Z(n2917) );
  AND U3091 ( .A(x[86]), .B(y[199]), .Z(n2855) );
  AND U3092 ( .A(x[76]), .B(y[209]), .Z(n3145) );
  AND U3093 ( .A(x[65]), .B(y[220]), .Z(n2854) );
  XOR U3094 ( .A(n3145), .B(n2854), .Z(n2856) );
  XOR U3095 ( .A(n2855), .B(n2856), .Z(n2916) );
  NAND U3096 ( .A(y[206]), .B(x[79]), .Z(n2859) );
  XOR U3097 ( .A(n3156), .B(n2859), .Z(n2861) );
  XNOR U3098 ( .A(n2860), .B(n2861), .Z(n2915) );
  XOR U3099 ( .A(n2916), .B(n2915), .Z(n2918) );
  XNOR U3100 ( .A(n2917), .B(n2918), .Z(n2948) );
  NANDN U3101 ( .A(n2665), .B(n2664), .Z(n2669) );
  OR U3102 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U3103 ( .A(n2669), .B(n2668), .Z(n2911) );
  XOR U3104 ( .A(n2912), .B(n2911), .Z(n2906) );
  NAND U3105 ( .A(n2671), .B(n2670), .Z(n2675) );
  NAND U3106 ( .A(n2673), .B(n2672), .Z(n2674) );
  AND U3107 ( .A(n2675), .B(n2674), .Z(n2904) );
  NANDN U3108 ( .A(n2676), .B(n2878), .Z(n2680) );
  NANDN U3109 ( .A(n2678), .B(n2677), .Z(n2679) );
  NAND U3110 ( .A(n2680), .B(n2679), .Z(n2930) );
  AND U3111 ( .A(x[89]), .B(y[196]), .Z(n2851) );
  AND U3112 ( .A(y[195]), .B(x[90]), .Z(n2848) );
  XOR U3113 ( .A(n2849), .B(n2848), .Z(n2850) );
  XOR U3114 ( .A(n2851), .B(n2850), .Z(n2928) );
  AND U3115 ( .A(y[193]), .B(x[92]), .Z(n2864) );
  XOR U3116 ( .A(o[29]), .B(n2864), .Z(n2938) );
  AND U3117 ( .A(x[64]), .B(y[221]), .Z(n2936) );
  AND U3118 ( .A(y[192]), .B(x[93]), .Z(n2935) );
  XOR U3119 ( .A(n2936), .B(n2935), .Z(n2937) );
  XNOR U3120 ( .A(n2938), .B(n2937), .Z(n2927) );
  XOR U3121 ( .A(n2930), .B(n2929), .Z(n2897) );
  NANDN U3122 ( .A(n2682), .B(n2681), .Z(n2686) );
  NANDN U3123 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U3124 ( .A(n2686), .B(n2685), .Z(n2887) );
  AND U3125 ( .A(o[28]), .B(n2687), .Z(n2827) );
  AND U3126 ( .A(x[80]), .B(y[205]), .Z(n2825) );
  AND U3127 ( .A(y[194]), .B(x[91]), .Z(n2824) );
  XOR U3128 ( .A(n2825), .B(n2824), .Z(n2826) );
  XOR U3129 ( .A(n2827), .B(n2826), .Z(n2886) );
  AND U3130 ( .A(x[66]), .B(y[219]), .Z(n2836) );
  XOR U3131 ( .A(n2837), .B(n2836), .Z(n2838) );
  XOR U3132 ( .A(n2839), .B(n2838), .Z(n2885) );
  XOR U3133 ( .A(n2886), .B(n2885), .Z(n2888) );
  XOR U3134 ( .A(n2887), .B(n2888), .Z(n2898) );
  NANDN U3135 ( .A(n2689), .B(n2688), .Z(n2693) );
  NANDN U3136 ( .A(n2691), .B(n2690), .Z(n2692) );
  NAND U3137 ( .A(n2693), .B(n2692), .Z(n2922) );
  ANDN U3138 ( .B(n2695), .A(n2694), .Z(n2699) );
  NAND U3139 ( .A(n2697), .B(n2696), .Z(n2698) );
  NANDN U3140 ( .A(n2699), .B(n2698), .Z(n2921) );
  XOR U3141 ( .A(n2922), .B(n2921), .Z(n2923) );
  NAND U3142 ( .A(n2701), .B(n2700), .Z(n2705) );
  NAND U3143 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U3144 ( .A(n2705), .B(n2704), .Z(n2820) );
  AND U3145 ( .A(y[210]), .B(x[75]), .Z(n2875) );
  AND U3146 ( .A(y[218]), .B(x[67]), .Z(n2873) );
  AND U3147 ( .A(x[81]), .B(y[204]), .Z(n2872) );
  XOR U3148 ( .A(n2873), .B(n2872), .Z(n2874) );
  XOR U3149 ( .A(n2875), .B(n2874), .Z(n2819) );
  AND U3150 ( .A(x[87]), .B(y[198]), .Z(n3161) );
  AND U3151 ( .A(x[77]), .B(y[208]), .Z(n2868) );
  AND U3152 ( .A(x[88]), .B(y[197]), .Z(n2867) );
  XOR U3153 ( .A(n2868), .B(n2867), .Z(n2869) );
  XOR U3154 ( .A(n3161), .B(n2869), .Z(n2818) );
  XOR U3155 ( .A(n2819), .B(n2818), .Z(n2821) );
  XNOR U3156 ( .A(n2820), .B(n2821), .Z(n2924) );
  NANDN U3157 ( .A(n2707), .B(n2706), .Z(n2711) );
  NANDN U3158 ( .A(n2709), .B(n2708), .Z(n2710) );
  AND U3159 ( .A(n2711), .B(n2710), .Z(n2813) );
  NANDN U3160 ( .A(n2713), .B(n2712), .Z(n2717) );
  NANDN U3161 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3162 ( .A(n2717), .B(n2716), .Z(n2843) );
  NAND U3163 ( .A(n2719), .B(n2718), .Z(n2723) );
  NAND U3164 ( .A(n2721), .B(n2720), .Z(n2722) );
  NAND U3165 ( .A(n2723), .B(n2722), .Z(n2842) );
  XOR U3166 ( .A(n2843), .B(n2842), .Z(n2845) );
  AND U3167 ( .A(y[213]), .B(x[72]), .Z(n2880) );
  AND U3168 ( .A(x[70]), .B(y[215]), .Z(n2725) );
  NAND U3169 ( .A(y[214]), .B(x[71]), .Z(n2724) );
  XNOR U3170 ( .A(n2725), .B(n2724), .Z(n2879) );
  XNOR U3171 ( .A(n2880), .B(n2879), .Z(n2933) );
  NAND U3172 ( .A(y[212]), .B(x[73]), .Z(n3112) );
  AND U3173 ( .A(x[69]), .B(y[216]), .Z(n2833) );
  AND U3174 ( .A(x[68]), .B(y[217]), .Z(n2831) );
  AND U3175 ( .A(y[211]), .B(x[74]), .Z(n2830) );
  XOR U3176 ( .A(n2831), .B(n2830), .Z(n2832) );
  XNOR U3177 ( .A(n2833), .B(n2832), .Z(n2934) );
  XOR U3178 ( .A(n3112), .B(n2934), .Z(n2726) );
  XNOR U3179 ( .A(n2933), .B(n2726), .Z(n2844) );
  XNOR U3180 ( .A(n2845), .B(n2844), .Z(n2812) );
  XNOR U3181 ( .A(n2813), .B(n2812), .Z(n2814) );
  XNOR U3182 ( .A(n2815), .B(n2814), .Z(n2903) );
  XNOR U3183 ( .A(n2904), .B(n2903), .Z(n2905) );
  XNOR U3184 ( .A(n2906), .B(n2905), .Z(n2957) );
  NANDN U3185 ( .A(n2728), .B(n2727), .Z(n2732) );
  NANDN U3186 ( .A(n2730), .B(n2729), .Z(n2731) );
  NAND U3187 ( .A(n2732), .B(n2731), .Z(n2958) );
  XNOR U3188 ( .A(n2957), .B(n2958), .Z(n2959) );
  NANDN U3189 ( .A(n2734), .B(n2733), .Z(n2738) );
  NANDN U3190 ( .A(n2736), .B(n2735), .Z(n2737) );
  AND U3191 ( .A(n2738), .B(n2737), .Z(n2952) );
  NANDN U3192 ( .A(n2740), .B(n2739), .Z(n2744) );
  NANDN U3193 ( .A(n2742), .B(n2741), .Z(n2743) );
  AND U3194 ( .A(n2744), .B(n2743), .Z(n2951) );
  XNOR U3195 ( .A(n2952), .B(n2951), .Z(n2953) );
  NANDN U3196 ( .A(n2746), .B(n2745), .Z(n2750) );
  OR U3197 ( .A(n2748), .B(n2747), .Z(n2749) );
  NAND U3198 ( .A(n2750), .B(n2749), .Z(n2965) );
  NANDN U3199 ( .A(n2752), .B(n2751), .Z(n2756) );
  NAND U3200 ( .A(n2754), .B(n2753), .Z(n2755) );
  AND U3201 ( .A(n2756), .B(n2755), .Z(n2894) );
  NANDN U3202 ( .A(n2758), .B(n2757), .Z(n2762) );
  OR U3203 ( .A(n2760), .B(n2759), .Z(n2761) );
  AND U3204 ( .A(n2762), .B(n2761), .Z(n2892) );
  NANDN U3205 ( .A(n2764), .B(n2763), .Z(n2768) );
  OR U3206 ( .A(n2766), .B(n2765), .Z(n2767) );
  NAND U3207 ( .A(n2768), .B(n2767), .Z(n2891) );
  XNOR U3208 ( .A(n2892), .B(n2891), .Z(n2893) );
  XNOR U3209 ( .A(n2894), .B(n2893), .Z(n2964) );
  NANDN U3210 ( .A(n2770), .B(n2769), .Z(n2774) );
  NANDN U3211 ( .A(n2772), .B(n2771), .Z(n2773) );
  AND U3212 ( .A(n2774), .B(n2773), .Z(n2963) );
  XOR U3213 ( .A(n2964), .B(n2963), .Z(n2966) );
  XOR U3214 ( .A(n2965), .B(n2966), .Z(n2954) );
  XOR U3215 ( .A(n2953), .B(n2954), .Z(n2960) );
  XOR U3216 ( .A(n2959), .B(n2960), .Z(n2808) );
  NANDN U3217 ( .A(n2776), .B(n2775), .Z(n2780) );
  NAND U3218 ( .A(n2778), .B(n2777), .Z(n2779) );
  AND U3219 ( .A(n2780), .B(n2779), .Z(n2807) );
  NAND U3220 ( .A(n2782), .B(n2781), .Z(n2786) );
  NAND U3221 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U3222 ( .A(n2786), .B(n2785), .Z(n2806) );
  XOR U3223 ( .A(n2807), .B(n2806), .Z(n2809) );
  XNOR U3224 ( .A(n2808), .B(n2809), .Z(n2801) );
  XOR U3225 ( .A(n2800), .B(n2801), .Z(n2803) );
  XOR U3226 ( .A(n2802), .B(n2803), .Z(n2799) );
  NAND U3227 ( .A(n2788), .B(n2787), .Z(n2792) );
  NAND U3228 ( .A(n2790), .B(n2789), .Z(n2791) );
  AND U3229 ( .A(n2792), .B(n2791), .Z(n2798) );
  XNOR U3230 ( .A(n2798), .B(n2797), .Z(n2796) );
  XNOR U3231 ( .A(n2799), .B(n2796), .Z(N62) );
  NAND U3232 ( .A(n2801), .B(n2800), .Z(n2805) );
  NAND U3233 ( .A(n2803), .B(n2802), .Z(n2804) );
  NAND U3234 ( .A(n2805), .B(n2804), .Z(n3264) );
  NANDN U3235 ( .A(n2807), .B(n2806), .Z(n2811) );
  NANDN U3236 ( .A(n2809), .B(n2808), .Z(n2810) );
  AND U3237 ( .A(n2811), .B(n2810), .Z(n2970) );
  NANDN U3238 ( .A(n2813), .B(n2812), .Z(n2817) );
  NAND U3239 ( .A(n2815), .B(n2814), .Z(n2816) );
  AND U3240 ( .A(n2817), .B(n2816), .Z(n3243) );
  NAND U3241 ( .A(n2819), .B(n2818), .Z(n2823) );
  NAND U3242 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U3243 ( .A(n2823), .B(n2822), .Z(n3226) );
  NAND U3244 ( .A(n2825), .B(n2824), .Z(n2829) );
  NAND U3245 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3246 ( .A(n2829), .B(n2828), .Z(n3177) );
  NAND U3247 ( .A(n2831), .B(n2830), .Z(n2835) );
  NAND U3248 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U3249 ( .A(n2835), .B(n2834), .Z(n3180) );
  AND U3250 ( .A(x[70]), .B(y[216]), .Z(n3026) );
  AND U3251 ( .A(x[69]), .B(y[217]), .Z(n3028) );
  AND U3252 ( .A(x[83]), .B(y[203]), .Z(n3027) );
  XOR U3253 ( .A(n3028), .B(n3027), .Z(n3025) );
  XNOR U3254 ( .A(n3026), .B(n3025), .Z(n2987) );
  AND U3255 ( .A(x[68]), .B(y[218]), .Z(n3140) );
  AND U3256 ( .A(x[67]), .B(y[219]), .Z(n3142) );
  AND U3257 ( .A(y[204]), .B(x[82]), .Z(n3141) );
  XOR U3258 ( .A(n3142), .B(n3141), .Z(n3139) );
  XOR U3259 ( .A(n3140), .B(n3139), .Z(n2990) );
  NAND U3260 ( .A(n2837), .B(n2836), .Z(n2841) );
  NAND U3261 ( .A(n2839), .B(n2838), .Z(n2840) );
  AND U3262 ( .A(n2841), .B(n2840), .Z(n2989) );
  XOR U3263 ( .A(n2987), .B(n2988), .Z(n3179) );
  XOR U3264 ( .A(n3180), .B(n3179), .Z(n3178) );
  XOR U3265 ( .A(n3177), .B(n3178), .Z(n3225) );
  NAND U3266 ( .A(n2843), .B(n2842), .Z(n2847) );
  NAND U3267 ( .A(n2845), .B(n2844), .Z(n2846) );
  AND U3268 ( .A(n2847), .B(n2846), .Z(n3227) );
  XOR U3269 ( .A(n3228), .B(n3227), .Z(n3246) );
  AND U3270 ( .A(n2849), .B(n2848), .Z(n2853) );
  NAND U3271 ( .A(n2851), .B(n2850), .Z(n2852) );
  NANDN U3272 ( .A(n2853), .B(n2852), .Z(n3171) );
  AND U3273 ( .A(n3145), .B(n2854), .Z(n2858) );
  NAND U3274 ( .A(n2856), .B(n2855), .Z(n2857) );
  NANDN U3275 ( .A(n2858), .B(n2857), .Z(n3174) );
  NANDN U3276 ( .A(n2859), .B(n3156), .Z(n2863) );
  NANDN U3277 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U3278 ( .A(n2863), .B(n2862), .Z(n3000) );
  AND U3279 ( .A(n2864), .B(o[29]), .Z(n3064) );
  AND U3280 ( .A(y[194]), .B(x[92]), .Z(n3066) );
  AND U3281 ( .A(x[80]), .B(y[206]), .Z(n3065) );
  XOR U3282 ( .A(n3066), .B(n3065), .Z(n3063) );
  XOR U3283 ( .A(n3064), .B(n3063), .Z(n3002) );
  AND U3284 ( .A(x[89]), .B(y[197]), .Z(n3160) );
  AND U3285 ( .A(y[198]), .B(x[88]), .Z(n2866) );
  NAND U3286 ( .A(y[199]), .B(x[87]), .Z(n2865) );
  XNOR U3287 ( .A(n2866), .B(n2865), .Z(n3159) );
  XNOR U3288 ( .A(n3160), .B(n3159), .Z(n3001) );
  XNOR U3289 ( .A(n3000), .B(n2999), .Z(n3173) );
  XOR U3290 ( .A(n3174), .B(n3173), .Z(n3172) );
  XOR U3291 ( .A(n3171), .B(n3172), .Z(n3220) );
  NAND U3292 ( .A(n2868), .B(n2867), .Z(n2871) );
  NAND U3293 ( .A(n3161), .B(n2869), .Z(n2870) );
  NAND U3294 ( .A(n2871), .B(n2870), .Z(n3202) );
  NAND U3295 ( .A(n2873), .B(n2872), .Z(n2877) );
  NAND U3296 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U3297 ( .A(n2877), .B(n2876), .Z(n2994) );
  AND U3298 ( .A(x[64]), .B(y[222]), .Z(n3116) );
  AND U3299 ( .A(y[193]), .B(x[93]), .Z(n3095) );
  XOR U3300 ( .A(o[30]), .B(n3095), .Z(n3118) );
  AND U3301 ( .A(y[192]), .B(x[94]), .Z(n3117) );
  XOR U3302 ( .A(n3118), .B(n3117), .Z(n3115) );
  XOR U3303 ( .A(n3116), .B(n3115), .Z(n2996) );
  AND U3304 ( .A(y[202]), .B(x[84]), .Z(n3059) );
  XOR U3305 ( .A(n3060), .B(n3059), .Z(n3058) );
  AND U3306 ( .A(y[214]), .B(x[72]), .Z(n3057) );
  XNOR U3307 ( .A(n3058), .B(n3057), .Z(n2995) );
  XNOR U3308 ( .A(n2994), .B(n2993), .Z(n3201) );
  XOR U3309 ( .A(n3202), .B(n3201), .Z(n3199) );
  AND U3310 ( .A(x[71]), .B(y[215]), .Z(n3154) );
  NAND U3311 ( .A(n2878), .B(n3154), .Z(n2882) );
  NAND U3312 ( .A(n2880), .B(n2879), .Z(n2881) );
  AND U3313 ( .A(n2882), .B(n2881), .Z(n3007) );
  AND U3314 ( .A(y[200]), .B(x[86]), .Z(n2884) );
  AND U3315 ( .A(x[85]), .B(y[201]), .Z(n2883) );
  XOR U3316 ( .A(n2884), .B(n2883), .Z(n3153) );
  XOR U3317 ( .A(n3154), .B(n3153), .Z(n3010) );
  AND U3318 ( .A(x[81]), .B(y[205]), .Z(n3014) );
  AND U3319 ( .A(x[66]), .B(y[220]), .Z(n3016) );
  AND U3320 ( .A(x[90]), .B(y[196]), .Z(n3015) );
  XOR U3321 ( .A(n3016), .B(n3015), .Z(n3013) );
  XNOR U3322 ( .A(n3014), .B(n3013), .Z(n3009) );
  XNOR U3323 ( .A(n3007), .B(n3008), .Z(n3200) );
  NAND U3324 ( .A(n2886), .B(n2885), .Z(n2890) );
  NAND U3325 ( .A(n2888), .B(n2887), .Z(n2889) );
  NAND U3326 ( .A(n2890), .B(n2889), .Z(n3221) );
  XOR U3327 ( .A(n3222), .B(n3221), .Z(n3219) );
  XOR U3328 ( .A(n3220), .B(n3219), .Z(n3245) );
  XNOR U3329 ( .A(n3243), .B(n3244), .Z(n3240) );
  NANDN U3330 ( .A(n2892), .B(n2891), .Z(n2896) );
  NANDN U3331 ( .A(n2894), .B(n2893), .Z(n2895) );
  AND U3332 ( .A(n2896), .B(n2895), .Z(n3239) );
  NANDN U3333 ( .A(n2898), .B(n2897), .Z(n2902) );
  NANDN U3334 ( .A(n2900), .B(n2899), .Z(n2901) );
  NAND U3335 ( .A(n2902), .B(n2901), .Z(n3237) );
  XOR U3336 ( .A(n3238), .B(n3237), .Z(n3256) );
  NANDN U3337 ( .A(n2904), .B(n2903), .Z(n2908) );
  NANDN U3338 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U3339 ( .A(n2908), .B(n2907), .Z(n3257) );
  NANDN U3340 ( .A(n2910), .B(n2909), .Z(n2914) );
  NAND U3341 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U3342 ( .A(n2914), .B(n2913), .Z(n3211) );
  NAND U3343 ( .A(n2916), .B(n2915), .Z(n2920) );
  NAND U3344 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3345 ( .A(n2920), .B(n2919), .Z(n3195) );
  NAND U3346 ( .A(n2922), .B(n2921), .Z(n2926) );
  NANDN U3347 ( .A(n2924), .B(n2923), .Z(n2925) );
  NAND U3348 ( .A(n2926), .B(n2925), .Z(n3196) );
  XNOR U3349 ( .A(n3195), .B(n3196), .Z(n3194) );
  NANDN U3350 ( .A(n2928), .B(n2927), .Z(n2932) );
  OR U3351 ( .A(n2930), .B(n2929), .Z(n2931) );
  NAND U3352 ( .A(n2932), .B(n2931), .Z(n3193) );
  XOR U3353 ( .A(n3194), .B(n3193), .Z(n3214) );
  NAND U3354 ( .A(n2936), .B(n2935), .Z(n2940) );
  NAND U3355 ( .A(n2938), .B(n2937), .Z(n2939) );
  NAND U3356 ( .A(n2940), .B(n2939), .Z(n3051) );
  AND U3357 ( .A(y[210]), .B(x[76]), .Z(n2941) );
  XOR U3358 ( .A(n2942), .B(n2941), .Z(n3147) );
  XOR U3359 ( .A(n3148), .B(n3147), .Z(n3110) );
  AND U3360 ( .A(x[73]), .B(y[213]), .Z(n2943) );
  XOR U3361 ( .A(n2944), .B(n2943), .Z(n3109) );
  XOR U3362 ( .A(n3110), .B(n3109), .Z(n3054) );
  AND U3363 ( .A(y[195]), .B(x[91]), .Z(n3022) );
  AND U3364 ( .A(x[65]), .B(y[221]), .Z(n3021) );
  XOR U3365 ( .A(n3022), .B(n3021), .Z(n3019) );
  XOR U3366 ( .A(n3020), .B(n3019), .Z(n3053) );
  XOR U3367 ( .A(n3054), .B(n3053), .Z(n3052) );
  XOR U3368 ( .A(n3051), .B(n3052), .Z(n2984) );
  NAND U3369 ( .A(n2946), .B(n2945), .Z(n2950) );
  NANDN U3370 ( .A(n2948), .B(n2947), .Z(n2949) );
  AND U3371 ( .A(n2950), .B(n2949), .Z(n2981) );
  XNOR U3372 ( .A(n2982), .B(n2981), .Z(n3213) );
  XNOR U3373 ( .A(n3211), .B(n3212), .Z(n3258) );
  XOR U3374 ( .A(n3256), .B(n3255), .Z(n2971) );
  NANDN U3375 ( .A(n2952), .B(n2951), .Z(n2956) );
  NAND U3376 ( .A(n2954), .B(n2953), .Z(n2955) );
  AND U3377 ( .A(n2956), .B(n2955), .Z(n2978) );
  NANDN U3378 ( .A(n2958), .B(n2957), .Z(n2962) );
  NAND U3379 ( .A(n2960), .B(n2959), .Z(n2961) );
  AND U3380 ( .A(n2962), .B(n2961), .Z(n2977) );
  XOR U3381 ( .A(n2978), .B(n2977), .Z(n2976) );
  NAND U3382 ( .A(n2964), .B(n2963), .Z(n2968) );
  NAND U3383 ( .A(n2966), .B(n2965), .Z(n2967) );
  AND U3384 ( .A(n2968), .B(n2967), .Z(n2975) );
  XNOR U3385 ( .A(n2976), .B(n2975), .Z(n2972) );
  XOR U3386 ( .A(n2970), .B(n2969), .Z(n3261) );
  XNOR U3387 ( .A(n3262), .B(n3261), .Z(N63) );
  NANDN U3388 ( .A(n2970), .B(n2969), .Z(n2974) );
  ANDN U3389 ( .B(n2972), .A(n2971), .Z(n2973) );
  ANDN U3390 ( .B(n2974), .A(n2973), .Z(n3254) );
  NAND U3391 ( .A(n2976), .B(n2975), .Z(n2980) );
  AND U3392 ( .A(n2978), .B(n2977), .Z(n2979) );
  ANDN U3393 ( .B(n2980), .A(n2979), .Z(n3236) );
  NAND U3394 ( .A(n2982), .B(n2981), .Z(n2986) );
  NANDN U3395 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U3396 ( .A(n2986), .B(n2985), .Z(n3210) );
  NANDN U3397 ( .A(n2988), .B(n2987), .Z(n2992) );
  NANDN U3398 ( .A(n2990), .B(n2989), .Z(n2991) );
  AND U3399 ( .A(n2992), .B(n2991), .Z(n3192) );
  NAND U3400 ( .A(n2994), .B(n2993), .Z(n2998) );
  NANDN U3401 ( .A(n2996), .B(n2995), .Z(n2997) );
  AND U3402 ( .A(n2998), .B(n2997), .Z(n3006) );
  NAND U3403 ( .A(n3000), .B(n2999), .Z(n3004) );
  NANDN U3404 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U3405 ( .A(n3004), .B(n3003), .Z(n3005) );
  XNOR U3406 ( .A(n3006), .B(n3005), .Z(n3190) );
  NANDN U3407 ( .A(n3008), .B(n3007), .Z(n3012) );
  NANDN U3408 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U3409 ( .A(n3012), .B(n3011), .Z(n3188) );
  NAND U3410 ( .A(n3014), .B(n3013), .Z(n3018) );
  NAND U3411 ( .A(n3016), .B(n3015), .Z(n3017) );
  AND U3412 ( .A(n3018), .B(n3017), .Z(n3050) );
  NAND U3413 ( .A(n3020), .B(n3019), .Z(n3024) );
  NAND U3414 ( .A(n3022), .B(n3021), .Z(n3023) );
  AND U3415 ( .A(n3024), .B(n3023), .Z(n3032) );
  NAND U3416 ( .A(n3026), .B(n3025), .Z(n3030) );
  NAND U3417 ( .A(n3028), .B(n3027), .Z(n3029) );
  NAND U3418 ( .A(n3030), .B(n3029), .Z(n3031) );
  XNOR U3419 ( .A(n3032), .B(n3031), .Z(n3048) );
  AND U3420 ( .A(y[216]), .B(x[71]), .Z(n3034) );
  NAND U3421 ( .A(y[218]), .B(x[69]), .Z(n3033) );
  XNOR U3422 ( .A(n3034), .B(n3033), .Z(n3038) );
  AND U3423 ( .A(y[221]), .B(x[66]), .Z(n3036) );
  NAND U3424 ( .A(y[200]), .B(x[87]), .Z(n3035) );
  XNOR U3425 ( .A(n3036), .B(n3035), .Z(n3037) );
  XOR U3426 ( .A(n3038), .B(n3037), .Z(n3046) );
  AND U3427 ( .A(x[91]), .B(y[196]), .Z(n3040) );
  NAND U3428 ( .A(x[70]), .B(y[217]), .Z(n3039) );
  XNOR U3429 ( .A(n3040), .B(n3039), .Z(n3044) );
  AND U3430 ( .A(y[220]), .B(x[67]), .Z(n3042) );
  NAND U3431 ( .A(x[82]), .B(y[205]), .Z(n3041) );
  XNOR U3432 ( .A(n3042), .B(n3041), .Z(n3043) );
  XNOR U3433 ( .A(n3044), .B(n3043), .Z(n3045) );
  XNOR U3434 ( .A(n3046), .B(n3045), .Z(n3047) );
  XNOR U3435 ( .A(n3048), .B(n3047), .Z(n3049) );
  XNOR U3436 ( .A(n3050), .B(n3049), .Z(n3138) );
  NAND U3437 ( .A(n3052), .B(n3051), .Z(n3056) );
  NAND U3438 ( .A(n3054), .B(n3053), .Z(n3055) );
  AND U3439 ( .A(n3056), .B(n3055), .Z(n3136) );
  NAND U3440 ( .A(n3058), .B(n3057), .Z(n3062) );
  NAND U3441 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U3442 ( .A(n3062), .B(n3061), .Z(n3070) );
  NAND U3443 ( .A(n3064), .B(n3063), .Z(n3068) );
  NAND U3444 ( .A(n3066), .B(n3065), .Z(n3067) );
  NAND U3445 ( .A(n3068), .B(n3067), .Z(n3069) );
  XNOR U3446 ( .A(n3070), .B(n3069), .Z(n3134) );
  AND U3447 ( .A(y[223]), .B(x[64]), .Z(n3072) );
  NAND U3448 ( .A(y[207]), .B(x[80]), .Z(n3071) );
  XNOR U3449 ( .A(n3072), .B(n3071), .Z(n3076) );
  AND U3450 ( .A(x[84]), .B(y[203]), .Z(n3074) );
  NAND U3451 ( .A(x[93]), .B(y[194]), .Z(n3073) );
  XNOR U3452 ( .A(n3074), .B(n3073), .Z(n3075) );
  XOR U3453 ( .A(n3076), .B(n3075), .Z(n3078) );
  AND U3454 ( .A(y[201]), .B(x[86]), .Z(n3155) );
  AND U3455 ( .A(y[213]), .B(x[74]), .Z(n3111) );
  XNOR U3456 ( .A(n3155), .B(n3111), .Z(n3077) );
  XNOR U3457 ( .A(n3078), .B(n3077), .Z(n3094) );
  AND U3458 ( .A(x[73]), .B(y[214]), .Z(n3080) );
  NAND U3459 ( .A(y[198]), .B(x[89]), .Z(n3079) );
  XNOR U3460 ( .A(n3080), .B(n3079), .Z(n3084) );
  AND U3461 ( .A(y[209]), .B(x[78]), .Z(n3082) );
  NAND U3462 ( .A(y[206]), .B(x[81]), .Z(n3081) );
  XNOR U3463 ( .A(n3082), .B(n3081), .Z(n3083) );
  XOR U3464 ( .A(n3084), .B(n3083), .Z(n3092) );
  AND U3465 ( .A(x[94]), .B(y[193]), .Z(n3086) );
  NAND U3466 ( .A(x[75]), .B(y[212]), .Z(n3085) );
  XNOR U3467 ( .A(n3086), .B(n3085), .Z(n3090) );
  AND U3468 ( .A(y[211]), .B(x[76]), .Z(n3088) );
  NAND U3469 ( .A(y[197]), .B(x[90]), .Z(n3087) );
  XNOR U3470 ( .A(n3088), .B(n3087), .Z(n3089) );
  XNOR U3471 ( .A(n3090), .B(n3089), .Z(n3091) );
  XNOR U3472 ( .A(n3092), .B(n3091), .Z(n3093) );
  XOR U3473 ( .A(n3094), .B(n3093), .Z(n3108) );
  AND U3474 ( .A(x[85]), .B(y[202]), .Z(n3102) );
  AND U3475 ( .A(n3095), .B(o[30]), .Z(n3100) );
  XOR U3476 ( .A(n3146), .B(o[31]), .Z(n3098) );
  XNOR U3477 ( .A(n3162), .B(n3096), .Z(n3097) );
  XNOR U3478 ( .A(n3098), .B(n3097), .Z(n3099) );
  XNOR U3479 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U3480 ( .A(n3102), .B(n3101), .Z(n3106) );
  AND U3481 ( .A(y[222]), .B(x[65]), .Z(n3104) );
  NAND U3482 ( .A(x[92]), .B(y[195]), .Z(n3103) );
  XNOR U3483 ( .A(n3104), .B(n3103), .Z(n3105) );
  XNOR U3484 ( .A(n3106), .B(n3105), .Z(n3107) );
  XNOR U3485 ( .A(n3108), .B(n3107), .Z(n3124) );
  NAND U3486 ( .A(n3110), .B(n3109), .Z(n3114) );
  NANDN U3487 ( .A(n3112), .B(n3111), .Z(n3113) );
  AND U3488 ( .A(n3114), .B(n3113), .Z(n3122) );
  NAND U3489 ( .A(n3116), .B(n3115), .Z(n3120) );
  NAND U3490 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U3491 ( .A(n3120), .B(n3119), .Z(n3121) );
  XNOR U3492 ( .A(n3122), .B(n3121), .Z(n3123) );
  XOR U3493 ( .A(n3124), .B(n3123), .Z(n3132) );
  AND U3494 ( .A(x[72]), .B(y[215]), .Z(n3126) );
  NAND U3495 ( .A(x[83]), .B(y[204]), .Z(n3125) );
  XNOR U3496 ( .A(n3126), .B(n3125), .Z(n3130) );
  AND U3497 ( .A(x[95]), .B(y[192]), .Z(n3128) );
  NAND U3498 ( .A(y[219]), .B(x[68]), .Z(n3127) );
  XNOR U3499 ( .A(n3128), .B(n3127), .Z(n3129) );
  XNOR U3500 ( .A(n3130), .B(n3129), .Z(n3131) );
  XNOR U3501 ( .A(n3132), .B(n3131), .Z(n3133) );
  XNOR U3502 ( .A(n3134), .B(n3133), .Z(n3135) );
  XNOR U3503 ( .A(n3136), .B(n3135), .Z(n3137) );
  XOR U3504 ( .A(n3138), .B(n3137), .Z(n3170) );
  NAND U3505 ( .A(n3140), .B(n3139), .Z(n3144) );
  NAND U3506 ( .A(n3142), .B(n3141), .Z(n3143) );
  AND U3507 ( .A(n3144), .B(n3143), .Z(n3152) );
  NAND U3508 ( .A(n3146), .B(n3145), .Z(n3150) );
  NAND U3509 ( .A(n3148), .B(n3147), .Z(n3149) );
  AND U3510 ( .A(n3150), .B(n3149), .Z(n3151) );
  XNOR U3511 ( .A(n3152), .B(n3151), .Z(n3168) );
  NAND U3512 ( .A(n3154), .B(n3153), .Z(n3158) );
  NAND U3513 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3514 ( .A(n3158), .B(n3157), .Z(n3166) );
  NAND U3515 ( .A(n3160), .B(n3159), .Z(n3164) );
  NAND U3516 ( .A(n3162), .B(n3161), .Z(n3163) );
  NAND U3517 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U3518 ( .A(n3166), .B(n3165), .Z(n3167) );
  XOR U3519 ( .A(n3168), .B(n3167), .Z(n3169) );
  XNOR U3520 ( .A(n3170), .B(n3169), .Z(n3186) );
  NAND U3521 ( .A(n3172), .B(n3171), .Z(n3176) );
  NAND U3522 ( .A(n3174), .B(n3173), .Z(n3175) );
  AND U3523 ( .A(n3176), .B(n3175), .Z(n3184) );
  NAND U3524 ( .A(n3178), .B(n3177), .Z(n3182) );
  NAND U3525 ( .A(n3180), .B(n3179), .Z(n3181) );
  NAND U3526 ( .A(n3182), .B(n3181), .Z(n3183) );
  XNOR U3527 ( .A(n3184), .B(n3183), .Z(n3185) );
  XNOR U3528 ( .A(n3186), .B(n3185), .Z(n3187) );
  XNOR U3529 ( .A(n3188), .B(n3187), .Z(n3189) );
  XNOR U3530 ( .A(n3190), .B(n3189), .Z(n3191) );
  XNOR U3531 ( .A(n3192), .B(n3191), .Z(n3208) );
  NAND U3532 ( .A(n3194), .B(n3193), .Z(n3198) );
  NANDN U3533 ( .A(n3196), .B(n3195), .Z(n3197) );
  AND U3534 ( .A(n3198), .B(n3197), .Z(n3206) );
  NANDN U3535 ( .A(n3200), .B(n3199), .Z(n3204) );
  NAND U3536 ( .A(n3202), .B(n3201), .Z(n3203) );
  NAND U3537 ( .A(n3204), .B(n3203), .Z(n3205) );
  XNOR U3538 ( .A(n3206), .B(n3205), .Z(n3207) );
  XNOR U3539 ( .A(n3208), .B(n3207), .Z(n3209) );
  XNOR U3540 ( .A(n3210), .B(n3209), .Z(n3218) );
  NANDN U3541 ( .A(n3212), .B(n3211), .Z(n3216) );
  NANDN U3542 ( .A(n3214), .B(n3213), .Z(n3215) );
  NAND U3543 ( .A(n3216), .B(n3215), .Z(n3217) );
  XNOR U3544 ( .A(n3218), .B(n3217), .Z(n3234) );
  NAND U3545 ( .A(n3220), .B(n3219), .Z(n3224) );
  NAND U3546 ( .A(n3222), .B(n3221), .Z(n3223) );
  AND U3547 ( .A(n3224), .B(n3223), .Z(n3232) );
  ANDN U3548 ( .B(n3226), .A(n3225), .Z(n3230) );
  AND U3549 ( .A(n3228), .B(n3227), .Z(n3229) );
  OR U3550 ( .A(n3230), .B(n3229), .Z(n3231) );
  XNOR U3551 ( .A(n3232), .B(n3231), .Z(n3233) );
  XNOR U3552 ( .A(n3234), .B(n3233), .Z(n3235) );
  XNOR U3553 ( .A(n3236), .B(n3235), .Z(n3252) );
  NAND U3554 ( .A(n3238), .B(n3237), .Z(n3242) );
  NANDN U3555 ( .A(n3240), .B(n3239), .Z(n3241) );
  AND U3556 ( .A(n3242), .B(n3241), .Z(n3250) );
  NANDN U3557 ( .A(n3244), .B(n3243), .Z(n3248) );
  NANDN U3558 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U3559 ( .A(n3248), .B(n3247), .Z(n3249) );
  XNOR U3560 ( .A(n3250), .B(n3249), .Z(n3251) );
  XNOR U3561 ( .A(n3252), .B(n3251), .Z(n3253) );
  XNOR U3562 ( .A(n3254), .B(n3253), .Z(n3270) );
  NAND U3563 ( .A(n3256), .B(n3255), .Z(n3260) );
  NANDN U3564 ( .A(n3258), .B(n3257), .Z(n3259) );
  AND U3565 ( .A(n3260), .B(n3259), .Z(n3268) );
  NAND U3566 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U3567 ( .A(n3264), .B(n3263), .Z(n3265) );
  NAND U3568 ( .A(n3266), .B(n3265), .Z(n3267) );
  XNOR U3569 ( .A(n3268), .B(n3267), .Z(n3269) );
  XNOR U3570 ( .A(n3270), .B(n3269), .Z(N64) );
  AND U3571 ( .A(x[64]), .B(y[224]), .Z(n3902) );
  XOR U3572 ( .A(n3902), .B(o[32]), .Z(N97) );
  AND U3573 ( .A(x[65]), .B(y[224]), .Z(n3280) );
  AND U3574 ( .A(x[64]), .B(y[225]), .Z(n3271) );
  XNOR U3575 ( .A(n3271), .B(o[33]), .Z(n3274) );
  XNOR U3576 ( .A(n3280), .B(n3274), .Z(n3276) );
  NAND U3577 ( .A(n3902), .B(o[32]), .Z(n3275) );
  XNOR U3578 ( .A(n3276), .B(n3275), .Z(N98) );
  AND U3579 ( .A(n3271), .B(o[33]), .Z(n3282) );
  AND U3580 ( .A(x[66]), .B(y[224]), .Z(n3273) );
  AND U3581 ( .A(y[225]), .B(x[65]), .Z(n3272) );
  XOR U3582 ( .A(n3273), .B(n3272), .Z(n3281) );
  XOR U3583 ( .A(n3282), .B(n3281), .Z(n3287) );
  NANDN U3584 ( .A(n3280), .B(n3274), .Z(n3278) );
  NAND U3585 ( .A(n3276), .B(n3275), .Z(n3277) );
  NAND U3586 ( .A(n3278), .B(n3277), .Z(n3285) );
  NAND U3587 ( .A(x[64]), .B(y[226]), .Z(n3290) );
  XNOR U3588 ( .A(o[34]), .B(n3290), .Z(n3286) );
  XOR U3589 ( .A(n3285), .B(n3286), .Z(n3279) );
  XNOR U3590 ( .A(n3287), .B(n3279), .Z(N99) );
  NAND U3591 ( .A(x[66]), .B(y[225]), .Z(n3299) );
  NANDN U3592 ( .A(n3299), .B(n3280), .Z(n3284) );
  NAND U3593 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U3594 ( .A(n3284), .B(n3283), .Z(n3306) );
  AND U3595 ( .A(x[65]), .B(y[226]), .Z(n3397) );
  XOR U3596 ( .A(n3397), .B(n3301), .Z(n3303) );
  AND U3597 ( .A(y[224]), .B(x[67]), .Z(n3289) );
  NAND U3598 ( .A(y[227]), .B(x[64]), .Z(n3288) );
  XNOR U3599 ( .A(n3289), .B(n3288), .Z(n3294) );
  ANDN U3600 ( .B(o[34]), .A(n3290), .Z(n3293) );
  XOR U3601 ( .A(n3294), .B(n3293), .Z(n3302) );
  XOR U3602 ( .A(n3303), .B(n3302), .Z(n3308) );
  XNOR U3603 ( .A(n3307), .B(n3308), .Z(n3291) );
  XOR U3604 ( .A(n3306), .B(n3291), .Z(N100) );
  AND U3605 ( .A(x[67]), .B(y[227]), .Z(n3292) );
  NAND U3606 ( .A(n3902), .B(n3292), .Z(n3296) );
  NAND U3607 ( .A(n3294), .B(n3293), .Z(n3295) );
  AND U3608 ( .A(n3296), .B(n3295), .Z(n3330) );
  AND U3609 ( .A(y[228]), .B(x[64]), .Z(n3298) );
  NAND U3610 ( .A(y[224]), .B(x[68]), .Z(n3297) );
  XNOR U3611 ( .A(n3298), .B(n3297), .Z(n3321) );
  ANDN U3612 ( .B(o[35]), .A(n3299), .Z(n3320) );
  XOR U3613 ( .A(n3321), .B(n3320), .Z(n3328) );
  AND U3614 ( .A(x[66]), .B(y[226]), .Z(n3449) );
  NAND U3615 ( .A(y[227]), .B(x[65]), .Z(n3300) );
  XNOR U3616 ( .A(n3449), .B(n3300), .Z(n3316) );
  NAND U3617 ( .A(x[67]), .B(y[225]), .Z(n3314) );
  XOR U3618 ( .A(o[36]), .B(n3314), .Z(n3317) );
  XNOR U3619 ( .A(n3316), .B(n3317), .Z(n3327) );
  XOR U3620 ( .A(n3328), .B(n3327), .Z(n3329) );
  XOR U3621 ( .A(n3330), .B(n3329), .Z(n3326) );
  NAND U3622 ( .A(n3397), .B(n3301), .Z(n3305) );
  NAND U3623 ( .A(n3303), .B(n3302), .Z(n3304) );
  NAND U3624 ( .A(n3305), .B(n3304), .Z(n3325) );
  XOR U3625 ( .A(n3325), .B(n3324), .Z(n3309) );
  XNOR U3626 ( .A(n3326), .B(n3309), .Z(N101) );
  AND U3627 ( .A(y[226]), .B(x[67]), .Z(n3311) );
  NAND U3628 ( .A(y[228]), .B(x[65]), .Z(n3310) );
  XNOR U3629 ( .A(n3311), .B(n3310), .Z(n3335) );
  AND U3630 ( .A(x[68]), .B(y[225]), .Z(n3344) );
  XOR U3631 ( .A(n3344), .B(o[37]), .Z(n3334) );
  XNOR U3632 ( .A(n3335), .B(n3334), .Z(n3338) );
  NAND U3633 ( .A(x[66]), .B(y[227]), .Z(n3406) );
  AND U3634 ( .A(y[229]), .B(x[64]), .Z(n3313) );
  NAND U3635 ( .A(y[224]), .B(x[69]), .Z(n3312) );
  XNOR U3636 ( .A(n3313), .B(n3312), .Z(n3341) );
  ANDN U3637 ( .B(o[36]), .A(n3314), .Z(n3340) );
  XOR U3638 ( .A(n3341), .B(n3340), .Z(n3339) );
  XOR U3639 ( .A(n3406), .B(n3339), .Z(n3315) );
  XOR U3640 ( .A(n3338), .B(n3315), .Z(n3350) );
  NANDN U3641 ( .A(n3406), .B(n3397), .Z(n3319) );
  NANDN U3642 ( .A(n3317), .B(n3316), .Z(n3318) );
  AND U3643 ( .A(n3319), .B(n3318), .Z(n3348) );
  AND U3644 ( .A(x[68]), .B(y[228]), .Z(n4121) );
  NAND U3645 ( .A(n4121), .B(n3902), .Z(n3323) );
  NAND U3646 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U3647 ( .A(n3323), .B(n3322), .Z(n3347) );
  XNOR U3648 ( .A(n3348), .B(n3347), .Z(n3349) );
  XOR U3649 ( .A(n3350), .B(n3349), .Z(n3356) );
  NAND U3650 ( .A(n3328), .B(n3327), .Z(n3332) );
  NANDN U3651 ( .A(n3330), .B(n3329), .Z(n3331) );
  AND U3652 ( .A(n3332), .B(n3331), .Z(n3355) );
  IV U3653 ( .A(n3355), .Z(n3353) );
  XOR U3654 ( .A(n3354), .B(n3353), .Z(n3333) );
  XNOR U3655 ( .A(n3356), .B(n3333), .Z(N102) );
  AND U3656 ( .A(x[67]), .B(y[228]), .Z(n3407) );
  NAND U3657 ( .A(n3407), .B(n3397), .Z(n3337) );
  NAND U3658 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U3659 ( .A(n3337), .B(n3336), .Z(n3361) );
  XOR U3660 ( .A(n3361), .B(n3362), .Z(n3364) );
  AND U3661 ( .A(x[69]), .B(y[229]), .Z(n3568) );
  AND U3662 ( .A(y[224]), .B(x[70]), .Z(n3343) );
  NAND U3663 ( .A(y[230]), .B(x[64]), .Z(n3342) );
  XNOR U3664 ( .A(n3343), .B(n3342), .Z(n3375) );
  NAND U3665 ( .A(n3344), .B(o[37]), .Z(n3376) );
  XNOR U3666 ( .A(n3375), .B(n3376), .Z(n3370) );
  XNOR U3667 ( .A(n3371), .B(n3370), .Z(n3373) );
  AND U3668 ( .A(y[228]), .B(x[66]), .Z(n3855) );
  NAND U3669 ( .A(y[227]), .B(x[67]), .Z(n3345) );
  XNOR U3670 ( .A(n3855), .B(n3345), .Z(n3380) );
  AND U3671 ( .A(y[229]), .B(x[65]), .Z(n3598) );
  NAND U3672 ( .A(y[226]), .B(x[68]), .Z(n3346) );
  XNOR U3673 ( .A(n3598), .B(n3346), .Z(n3382) );
  NAND U3674 ( .A(x[69]), .B(y[225]), .Z(n3389) );
  XOR U3675 ( .A(n3382), .B(n3381), .Z(n3379) );
  XOR U3676 ( .A(n3380), .B(n3379), .Z(n3372) );
  XOR U3677 ( .A(n3373), .B(n3372), .Z(n3363) );
  XNOR U3678 ( .A(n3364), .B(n3363), .Z(n3369) );
  NANDN U3679 ( .A(n3348), .B(n3347), .Z(n3352) );
  NAND U3680 ( .A(n3350), .B(n3349), .Z(n3351) );
  NAND U3681 ( .A(n3352), .B(n3351), .Z(n3368) );
  NANDN U3682 ( .A(n3353), .B(n3354), .Z(n3359) );
  NOR U3683 ( .A(n3355), .B(n3354), .Z(n3357) );
  OR U3684 ( .A(n3357), .B(n3356), .Z(n3358) );
  AND U3685 ( .A(n3359), .B(n3358), .Z(n3367) );
  XOR U3686 ( .A(n3368), .B(n3367), .Z(n3360) );
  XNOR U3687 ( .A(n3369), .B(n3360), .Z(N103) );
  NAND U3688 ( .A(n3362), .B(n3361), .Z(n3366) );
  NAND U3689 ( .A(n3364), .B(n3363), .Z(n3365) );
  NAND U3690 ( .A(n3366), .B(n3365), .Z(n3427) );
  AND U3691 ( .A(y[230]), .B(x[65]), .Z(n3770) );
  NAND U3692 ( .A(y[226]), .B(x[69]), .Z(n3374) );
  XNOR U3693 ( .A(n3770), .B(n3374), .Z(n3400) );
  NAND U3694 ( .A(x[70]), .B(y[225]), .Z(n3403) );
  XNOR U3695 ( .A(o[39]), .B(n3403), .Z(n3399) );
  XOR U3696 ( .A(n3400), .B(n3399), .Z(n3418) );
  AND U3697 ( .A(x[70]), .B(y[230]), .Z(n3617) );
  NAND U3698 ( .A(n3902), .B(n3617), .Z(n3378) );
  NANDN U3699 ( .A(n3376), .B(n3375), .Z(n3377) );
  AND U3700 ( .A(n3378), .B(n3377), .Z(n3417) );
  XOR U3701 ( .A(n3420), .B(n3419), .Z(n3424) );
  AND U3702 ( .A(x[68]), .B(y[229]), .Z(n3907) );
  NAND U3703 ( .A(n3907), .B(n3397), .Z(n3384) );
  NAND U3704 ( .A(n3382), .B(n3381), .Z(n3383) );
  AND U3705 ( .A(n3384), .B(n3383), .Z(n3394) );
  AND U3706 ( .A(y[229]), .B(x[66]), .Z(n3386) );
  NAND U3707 ( .A(y[227]), .B(x[68]), .Z(n3385) );
  XNOR U3708 ( .A(n3386), .B(n3385), .Z(n3408) );
  XOR U3709 ( .A(n3408), .B(n3407), .Z(n3392) );
  AND U3710 ( .A(y[224]), .B(x[71]), .Z(n3388) );
  NAND U3711 ( .A(y[231]), .B(x[64]), .Z(n3387) );
  XNOR U3712 ( .A(n3388), .B(n3387), .Z(n3412) );
  ANDN U3713 ( .B(o[38]), .A(n3389), .Z(n3411) );
  XNOR U3714 ( .A(n3412), .B(n3411), .Z(n3391) );
  XOR U3715 ( .A(n3394), .B(n3393), .Z(n3423) );
  XOR U3716 ( .A(n3424), .B(n3423), .Z(n3425) );
  XOR U3717 ( .A(n3426), .B(n3425), .Z(n3429) );
  XNOR U3718 ( .A(n3428), .B(n3429), .Z(n3390) );
  XNOR U3719 ( .A(n3427), .B(n3390), .Z(N104) );
  NANDN U3720 ( .A(n3392), .B(n3391), .Z(n3396) );
  NAND U3721 ( .A(n3394), .B(n3393), .Z(n3395) );
  AND U3722 ( .A(n3396), .B(n3395), .Z(n3462) );
  AND U3723 ( .A(x[69]), .B(y[230]), .Z(n3398) );
  NAND U3724 ( .A(n3398), .B(n3397), .Z(n3402) );
  NAND U3725 ( .A(n3400), .B(n3399), .Z(n3401) );
  AND U3726 ( .A(n3402), .B(n3401), .Z(n3460) );
  ANDN U3727 ( .B(o[39]), .A(n3403), .Z(n3440) );
  AND U3728 ( .A(y[231]), .B(x[65]), .Z(n3897) );
  NAND U3729 ( .A(y[227]), .B(x[69]), .Z(n3404) );
  XNOR U3730 ( .A(n3897), .B(n3404), .Z(n3441) );
  XNOR U3731 ( .A(n3440), .B(n3441), .Z(n3445) );
  NAND U3732 ( .A(x[67]), .B(y[229]), .Z(n4226) );
  AND U3733 ( .A(y[230]), .B(x[66]), .Z(n4302) );
  AND U3734 ( .A(y[226]), .B(x[70]), .Z(n3405) );
  XOR U3735 ( .A(n4302), .B(n3405), .Z(n3450) );
  XOR U3736 ( .A(n4121), .B(n3450), .Z(n3444) );
  XOR U3737 ( .A(n3445), .B(n3446), .Z(n3459) );
  XNOR U3738 ( .A(n3462), .B(n3461), .Z(n3470) );
  NANDN U3739 ( .A(n3406), .B(n3907), .Z(n3410) );
  NAND U3740 ( .A(n3408), .B(n3407), .Z(n3409) );
  AND U3741 ( .A(n3410), .B(n3409), .Z(n3456) );
  AND U3742 ( .A(x[71]), .B(y[231]), .Z(n3791) );
  NAND U3743 ( .A(n3902), .B(n3791), .Z(n3414) );
  NAND U3744 ( .A(n3412), .B(n3411), .Z(n3413) );
  AND U3745 ( .A(n3414), .B(n3413), .Z(n3454) );
  AND U3746 ( .A(y[224]), .B(x[72]), .Z(n3416) );
  NAND U3747 ( .A(y[232]), .B(x[64]), .Z(n3415) );
  XNOR U3748 ( .A(n3416), .B(n3415), .Z(n3432) );
  NAND U3749 ( .A(x[71]), .B(y[225]), .Z(n3435) );
  XNOR U3750 ( .A(o[40]), .B(n3435), .Z(n3431) );
  XOR U3751 ( .A(n3432), .B(n3431), .Z(n3453) );
  NANDN U3752 ( .A(n3418), .B(n3417), .Z(n3422) );
  NAND U3753 ( .A(n3420), .B(n3419), .Z(n3421) );
  NAND U3754 ( .A(n3422), .B(n3421), .Z(n3468) );
  XOR U3755 ( .A(n3470), .B(n3471), .Z(n3467) );
  XOR U3756 ( .A(n3466), .B(n3465), .Z(n3430) );
  XNOR U3757 ( .A(n3467), .B(n3430), .Z(N105) );
  AND U3758 ( .A(x[72]), .B(y[232]), .Z(n3922) );
  NAND U3759 ( .A(n3922), .B(n3902), .Z(n3434) );
  NAND U3760 ( .A(n3432), .B(n3431), .Z(n3433) );
  AND U3761 ( .A(n3434), .B(n3433), .Z(n3510) );
  ANDN U3762 ( .B(o[40]), .A(n3435), .Z(n3484) );
  AND U3763 ( .A(y[226]), .B(x[71]), .Z(n3846) );
  NAND U3764 ( .A(y[228]), .B(x[69]), .Z(n3436) );
  XNOR U3765 ( .A(n3846), .B(n3436), .Z(n3483) );
  XOR U3766 ( .A(n3484), .B(n3483), .Z(n3508) );
  AND U3767 ( .A(y[224]), .B(x[73]), .Z(n3438) );
  NAND U3768 ( .A(y[233]), .B(x[64]), .Z(n3437) );
  XNOR U3769 ( .A(n3438), .B(n3437), .Z(n3490) );
  NAND U3770 ( .A(x[72]), .B(y[225]), .Z(n3499) );
  XNOR U3771 ( .A(o[41]), .B(n3499), .Z(n3489) );
  XNOR U3772 ( .A(n3490), .B(n3489), .Z(n3507) );
  XNOR U3773 ( .A(n3508), .B(n3507), .Z(n3509) );
  XNOR U3774 ( .A(n3510), .B(n3509), .Z(n3504) );
  AND U3775 ( .A(y[227]), .B(x[70]), .Z(n3859) );
  NAND U3776 ( .A(y[232]), .B(x[65]), .Z(n3439) );
  XNOR U3777 ( .A(n3859), .B(n3439), .Z(n3494) );
  XOR U3778 ( .A(n3907), .B(n3494), .Z(n3514) );
  AND U3779 ( .A(x[66]), .B(y[231]), .Z(n4101) );
  NAND U3780 ( .A(x[67]), .B(y[230]), .Z(n3869) );
  XNOR U3781 ( .A(n4101), .B(n3869), .Z(n3513) );
  XOR U3782 ( .A(n3514), .B(n3513), .Z(n3502) );
  NAND U3783 ( .A(x[69]), .B(y[231]), .Z(n3697) );
  AND U3784 ( .A(x[65]), .B(y[227]), .Z(n3493) );
  NANDN U3785 ( .A(n3697), .B(n3493), .Z(n3443) );
  NAND U3786 ( .A(n3441), .B(n3440), .Z(n3442) );
  NAND U3787 ( .A(n3443), .B(n3442), .Z(n3501) );
  XOR U3788 ( .A(n3502), .B(n3501), .Z(n3503) );
  XNOR U3789 ( .A(n3504), .B(n3503), .Z(n3477) );
  NANDN U3790 ( .A(n3444), .B(n4226), .Z(n3448) );
  NANDN U3791 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U3792 ( .A(n3448), .B(n3447), .Z(n3475) );
  NAND U3793 ( .A(n3617), .B(n3449), .Z(n3452) );
  NAND U3794 ( .A(n4121), .B(n3450), .Z(n3451) );
  AND U3795 ( .A(n3452), .B(n3451), .Z(n3476) );
  XNOR U3796 ( .A(n3475), .B(n3476), .Z(n3478) );
  NANDN U3797 ( .A(n3454), .B(n3453), .Z(n3458) );
  NANDN U3798 ( .A(n3456), .B(n3455), .Z(n3457) );
  AND U3799 ( .A(n3458), .B(n3457), .Z(n3518) );
  NANDN U3800 ( .A(n3460), .B(n3459), .Z(n3464) );
  NAND U3801 ( .A(n3462), .B(n3461), .Z(n3463) );
  NAND U3802 ( .A(n3464), .B(n3463), .Z(n3517) );
  XNOR U3803 ( .A(n3519), .B(n3520), .Z(n3525) );
  NANDN U3804 ( .A(n3469), .B(n3468), .Z(n3473) );
  NANDN U3805 ( .A(n3471), .B(n3470), .Z(n3472) );
  AND U3806 ( .A(n3473), .B(n3472), .Z(n3523) );
  XOR U3807 ( .A(n3524), .B(n3523), .Z(n3474) );
  XNOR U3808 ( .A(n3525), .B(n3474), .Z(N106) );
  NAND U3809 ( .A(n3476), .B(n3475), .Z(n3480) );
  NANDN U3810 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3811 ( .A(n3480), .B(n3479), .Z(n3583) );
  AND U3812 ( .A(x[71]), .B(y[228]), .Z(n3482) );
  AND U3813 ( .A(x[69]), .B(y[226]), .Z(n3481) );
  NAND U3814 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U3815 ( .A(n3484), .B(n3483), .Z(n3485) );
  AND U3816 ( .A(n3486), .B(n3485), .Z(n3575) );
  AND U3817 ( .A(y[227]), .B(x[71]), .Z(n3488) );
  NAND U3818 ( .A(y[230]), .B(x[68]), .Z(n3487) );
  XNOR U3819 ( .A(n3488), .B(n3487), .Z(n3547) );
  AND U3820 ( .A(x[70]), .B(y[228]), .Z(n3546) );
  XOR U3821 ( .A(n3547), .B(n3546), .Z(n3573) );
  AND U3822 ( .A(x[72]), .B(y[226]), .Z(n3766) );
  NAND U3823 ( .A(x[73]), .B(y[225]), .Z(n3556) );
  XNOR U3824 ( .A(o[42]), .B(n3556), .Z(n3567) );
  XOR U3825 ( .A(n3766), .B(n3567), .Z(n3569) );
  XNOR U3826 ( .A(n3569), .B(n3568), .Z(n3572) );
  XNOR U3827 ( .A(n3573), .B(n3572), .Z(n3574) );
  XOR U3828 ( .A(n3575), .B(n3574), .Z(n3536) );
  AND U3829 ( .A(x[73]), .B(y[233]), .Z(n4130) );
  NAND U3830 ( .A(n4130), .B(n3902), .Z(n3492) );
  NAND U3831 ( .A(n3490), .B(n3489), .Z(n3491) );
  AND U3832 ( .A(n3492), .B(n3491), .Z(n3534) );
  AND U3833 ( .A(x[70]), .B(y[232]), .Z(n3801) );
  NAND U3834 ( .A(n3801), .B(n3493), .Z(n3496) );
  NAND U3835 ( .A(n3907), .B(n3494), .Z(n3495) );
  AND U3836 ( .A(n3496), .B(n3495), .Z(n3542) );
  AND U3837 ( .A(y[224]), .B(x[74]), .Z(n3498) );
  NAND U3838 ( .A(y[234]), .B(x[64]), .Z(n3497) );
  XNOR U3839 ( .A(n3498), .B(n3497), .Z(n3551) );
  ANDN U3840 ( .B(o[41]), .A(n3499), .Z(n3550) );
  XOR U3841 ( .A(n3551), .B(n3550), .Z(n3540) );
  AND U3842 ( .A(y[231]), .B(x[67]), .Z(n4439) );
  NAND U3843 ( .A(y[233]), .B(x[65]), .Z(n3500) );
  XNOR U3844 ( .A(n4439), .B(n3500), .Z(n3563) );
  NAND U3845 ( .A(x[66]), .B(y[232]), .Z(n3564) );
  XNOR U3846 ( .A(n3563), .B(n3564), .Z(n3539) );
  XOR U3847 ( .A(n3540), .B(n3539), .Z(n3541) );
  XNOR U3848 ( .A(n3542), .B(n3541), .Z(n3533) );
  XNOR U3849 ( .A(n3534), .B(n3533), .Z(n3535) );
  XNOR U3850 ( .A(n3536), .B(n3535), .Z(n3582) );
  NAND U3851 ( .A(n3502), .B(n3501), .Z(n3506) );
  NAND U3852 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U3853 ( .A(n3506), .B(n3505), .Z(n3530) );
  NANDN U3854 ( .A(n3508), .B(n3507), .Z(n3512) );
  NAND U3855 ( .A(n3510), .B(n3509), .Z(n3511) );
  AND U3856 ( .A(n3512), .B(n3511), .Z(n3527) );
  ANDN U3857 ( .B(n3869), .A(n4101), .Z(n3516) );
  NANDN U3858 ( .A(n3514), .B(n3513), .Z(n3515) );
  NANDN U3859 ( .A(n3516), .B(n3515), .Z(n3528) );
  XNOR U3860 ( .A(n3527), .B(n3528), .Z(n3529) );
  XOR U3861 ( .A(n3530), .B(n3529), .Z(n3581) );
  XOR U3862 ( .A(n3583), .B(n3584), .Z(n3580) );
  NANDN U3863 ( .A(n3518), .B(n3517), .Z(n3522) );
  NAND U3864 ( .A(n3520), .B(n3519), .Z(n3521) );
  NAND U3865 ( .A(n3522), .B(n3521), .Z(n3578) );
  XOR U3866 ( .A(n3578), .B(n3579), .Z(n3526) );
  XNOR U3867 ( .A(n3580), .B(n3526), .Z(N107) );
  NANDN U3868 ( .A(n3528), .B(n3527), .Z(n3532) );
  NANDN U3869 ( .A(n3530), .B(n3529), .Z(n3531) );
  AND U3870 ( .A(n3532), .B(n3531), .Z(n3652) );
  NANDN U3871 ( .A(n3534), .B(n3533), .Z(n3538) );
  NANDN U3872 ( .A(n3536), .B(n3535), .Z(n3537) );
  AND U3873 ( .A(n3538), .B(n3537), .Z(n3650) );
  NAND U3874 ( .A(n3540), .B(n3539), .Z(n3544) );
  NANDN U3875 ( .A(n3542), .B(n3541), .Z(n3543) );
  AND U3876 ( .A(n3544), .B(n3543), .Z(n3639) );
  AND U3877 ( .A(x[71]), .B(y[230]), .Z(n3692) );
  AND U3878 ( .A(x[68]), .B(y[227]), .Z(n3545) );
  NAND U3879 ( .A(n3692), .B(n3545), .Z(n3549) );
  NAND U3880 ( .A(n3547), .B(n3546), .Z(n3548) );
  AND U3881 ( .A(n3549), .B(n3548), .Z(n3637) );
  AND U3882 ( .A(x[74]), .B(y[234]), .Z(n4308) );
  NAND U3883 ( .A(n4308), .B(n3902), .Z(n3553) );
  NAND U3884 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U3885 ( .A(n3553), .B(n3552), .Z(n3633) );
  AND U3886 ( .A(y[224]), .B(x[75]), .Z(n3555) );
  NAND U3887 ( .A(y[235]), .B(x[64]), .Z(n3554) );
  XNOR U3888 ( .A(n3555), .B(n3554), .Z(n3609) );
  ANDN U3889 ( .B(o[42]), .A(n3556), .Z(n3608) );
  XOR U3890 ( .A(n3609), .B(n3608), .Z(n3631) );
  AND U3891 ( .A(y[229]), .B(x[70]), .Z(n3558) );
  NAND U3892 ( .A(y[234]), .B(x[65]), .Z(n3557) );
  XNOR U3893 ( .A(n3558), .B(n3557), .Z(n3600) );
  NAND U3894 ( .A(x[74]), .B(y[225]), .Z(n3618) );
  XNOR U3895 ( .A(o[43]), .B(n3618), .Z(n3599) );
  XOR U3896 ( .A(n3600), .B(n3599), .Z(n3630) );
  XOR U3897 ( .A(n3631), .B(n3630), .Z(n3632) );
  XNOR U3898 ( .A(n3633), .B(n3632), .Z(n3636) );
  XNOR U3899 ( .A(n3637), .B(n3636), .Z(n3638) );
  XOR U3900 ( .A(n3639), .B(n3638), .Z(n3621) );
  AND U3901 ( .A(x[67]), .B(y[232]), .Z(n4575) );
  AND U3902 ( .A(y[233]), .B(x[66]), .Z(n3560) );
  NAND U3903 ( .A(y[230]), .B(x[69]), .Z(n3559) );
  XNOR U3904 ( .A(n3560), .B(n3559), .Z(n3595) );
  AND U3905 ( .A(x[68]), .B(y[231]), .Z(n3594) );
  XNOR U3906 ( .A(n3595), .B(n3594), .Z(n3625) );
  XNOR U3907 ( .A(n4575), .B(n3625), .Z(n3627) );
  AND U3908 ( .A(y[226]), .B(x[73]), .Z(n3562) );
  NAND U3909 ( .A(y[228]), .B(x[71]), .Z(n3561) );
  XNOR U3910 ( .A(n3562), .B(n3561), .Z(n3613) );
  AND U3911 ( .A(x[72]), .B(y[227]), .Z(n3612) );
  XNOR U3912 ( .A(n3613), .B(n3612), .Z(n3626) );
  XOR U3913 ( .A(n3627), .B(n3626), .Z(n3591) );
  NAND U3914 ( .A(x[67]), .B(y[233]), .Z(n3688) );
  NANDN U3915 ( .A(n3688), .B(n3897), .Z(n3566) );
  NANDN U3916 ( .A(n3564), .B(n3563), .Z(n3565) );
  AND U3917 ( .A(n3566), .B(n3565), .Z(n3589) );
  NAND U3918 ( .A(n3766), .B(n3567), .Z(n3571) );
  NAND U3919 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U3920 ( .A(n3571), .B(n3570), .Z(n3588) );
  XNOR U3921 ( .A(n3589), .B(n3588), .Z(n3590) );
  XOR U3922 ( .A(n3591), .B(n3590), .Z(n3620) );
  NANDN U3923 ( .A(n3573), .B(n3572), .Z(n3577) );
  NAND U3924 ( .A(n3575), .B(n3574), .Z(n3576) );
  NAND U3925 ( .A(n3577), .B(n3576), .Z(n3619) );
  XOR U3926 ( .A(n3620), .B(n3619), .Z(n3622) );
  XNOR U3927 ( .A(n3621), .B(n3622), .Z(n3649) );
  XNOR U3928 ( .A(n3650), .B(n3649), .Z(n3651) );
  XOR U3929 ( .A(n3652), .B(n3651), .Z(n3645) );
  NANDN U3930 ( .A(n3582), .B(n3581), .Z(n3586) );
  NAND U3931 ( .A(n3584), .B(n3583), .Z(n3585) );
  AND U3932 ( .A(n3586), .B(n3585), .Z(n3643) );
  IV U3933 ( .A(n3643), .Z(n3642) );
  XOR U3934 ( .A(n3644), .B(n3642), .Z(n3587) );
  XNOR U3935 ( .A(n3645), .B(n3587), .Z(N108) );
  NANDN U3936 ( .A(n3589), .B(n3588), .Z(n3593) );
  NANDN U3937 ( .A(n3591), .B(n3590), .Z(n3592) );
  AND U3938 ( .A(n3593), .B(n3592), .Z(n3729) );
  AND U3939 ( .A(x[69]), .B(y[233]), .Z(n4094) );
  NAND U3940 ( .A(n4302), .B(n4094), .Z(n3597) );
  NAND U3941 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U3942 ( .A(n3597), .B(n3596), .Z(n3676) );
  AND U3943 ( .A(x[70]), .B(y[234]), .Z(n3913) );
  NAND U3944 ( .A(n3913), .B(n3598), .Z(n3602) );
  NAND U3945 ( .A(n3600), .B(n3599), .Z(n3601) );
  NAND U3946 ( .A(n3602), .B(n3601), .Z(n3675) );
  XOR U3947 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U3948 ( .A(x[73]), .B(y[227]), .Z(n4297) );
  AND U3949 ( .A(y[226]), .B(x[74]), .Z(n4339) );
  NAND U3950 ( .A(y[232]), .B(x[68]), .Z(n3603) );
  XOR U3951 ( .A(n4339), .B(n3603), .Z(n3719) );
  XNOR U3952 ( .A(n4297), .B(n3719), .Z(n3698) );
  NAND U3953 ( .A(x[71]), .B(y[229]), .Z(n3696) );
  XOR U3954 ( .A(n3697), .B(n3696), .Z(n3699) );
  AND U3955 ( .A(y[224]), .B(x[76]), .Z(n3605) );
  NAND U3956 ( .A(y[236]), .B(x[64]), .Z(n3604) );
  XNOR U3957 ( .A(n3605), .B(n3604), .Z(n3713) );
  NAND U3958 ( .A(x[75]), .B(y[225]), .Z(n3693) );
  XNOR U3959 ( .A(o[44]), .B(n3693), .Z(n3712) );
  XOR U3960 ( .A(n3713), .B(n3712), .Z(n3682) );
  AND U3961 ( .A(y[228]), .B(x[72]), .Z(n3607) );
  NAND U3962 ( .A(y[234]), .B(x[66]), .Z(n3606) );
  XNOR U3963 ( .A(n3607), .B(n3606), .Z(n3687) );
  XOR U3964 ( .A(n3682), .B(n3681), .Z(n3683) );
  XNOR U3965 ( .A(n3677), .B(n3678), .Z(n3727) );
  AND U3966 ( .A(x[75]), .B(y[235]), .Z(n4685) );
  NAND U3967 ( .A(n4685), .B(n3902), .Z(n3611) );
  NAND U3968 ( .A(n3609), .B(n3608), .Z(n3610) );
  AND U3969 ( .A(n3611), .B(n3610), .Z(n3705) );
  AND U3970 ( .A(x[73]), .B(y[228]), .Z(n3695) );
  NAND U3971 ( .A(n3846), .B(n3695), .Z(n3615) );
  NAND U3972 ( .A(n3613), .B(n3612), .Z(n3614) );
  AND U3973 ( .A(n3615), .B(n3614), .Z(n3703) );
  NAND U3974 ( .A(y[235]), .B(x[65]), .Z(n3616) );
  XNOR U3975 ( .A(n3617), .B(n3616), .Z(n3709) );
  ANDN U3976 ( .B(o[43]), .A(n3618), .Z(n3708) );
  XOR U3977 ( .A(n3709), .B(n3708), .Z(n3702) );
  XNOR U3978 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR U3979 ( .A(n3705), .B(n3704), .Z(n3726) );
  XOR U3980 ( .A(n3727), .B(n3726), .Z(n3728) );
  XOR U3981 ( .A(n3729), .B(n3728), .Z(n3657) );
  NAND U3982 ( .A(n3620), .B(n3619), .Z(n3624) );
  NAND U3983 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U3984 ( .A(n3624), .B(n3623), .Z(n3656) );
  XOR U3985 ( .A(n3657), .B(n3656), .Z(n3659) );
  NANDN U3986 ( .A(n4575), .B(n3625), .Z(n3629) );
  NAND U3987 ( .A(n3627), .B(n3626), .Z(n3628) );
  AND U3988 ( .A(n3629), .B(n3628), .Z(n3670) );
  NAND U3989 ( .A(n3631), .B(n3630), .Z(n3635) );
  NANDN U3990 ( .A(n3633), .B(n3632), .Z(n3634) );
  AND U3991 ( .A(n3635), .B(n3634), .Z(n3669) );
  XNOR U3992 ( .A(n3670), .B(n3669), .Z(n3671) );
  NANDN U3993 ( .A(n3637), .B(n3636), .Z(n3641) );
  NANDN U3994 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U3995 ( .A(n3641), .B(n3640), .Z(n3672) );
  XNOR U3996 ( .A(n3671), .B(n3672), .Z(n3658) );
  XNOR U3997 ( .A(n3659), .B(n3658), .Z(n3665) );
  OR U3998 ( .A(n3644), .B(n3642), .Z(n3648) );
  ANDN U3999 ( .B(n3644), .A(n3643), .Z(n3646) );
  OR U4000 ( .A(n3646), .B(n3645), .Z(n3647) );
  AND U4001 ( .A(n3648), .B(n3647), .Z(n3663) );
  NANDN U4002 ( .A(n3650), .B(n3649), .Z(n3654) );
  NANDN U4003 ( .A(n3652), .B(n3651), .Z(n3653) );
  AND U4004 ( .A(n3654), .B(n3653), .Z(n3664) );
  IV U4005 ( .A(n3664), .Z(n3662) );
  XOR U4006 ( .A(n3663), .B(n3662), .Z(n3655) );
  XNOR U4007 ( .A(n3665), .B(n3655), .Z(N109) );
  NAND U4008 ( .A(n3657), .B(n3656), .Z(n3661) );
  NAND U4009 ( .A(n3659), .B(n3658), .Z(n3660) );
  AND U4010 ( .A(n3661), .B(n3660), .Z(n3740) );
  NANDN U4011 ( .A(n3662), .B(n3663), .Z(n3668) );
  NOR U4012 ( .A(n3664), .B(n3663), .Z(n3666) );
  OR U4013 ( .A(n3666), .B(n3665), .Z(n3667) );
  AND U4014 ( .A(n3668), .B(n3667), .Z(n3739) );
  NANDN U4015 ( .A(n3670), .B(n3669), .Z(n3674) );
  NANDN U4016 ( .A(n3672), .B(n3671), .Z(n3673) );
  AND U4017 ( .A(n3674), .B(n3673), .Z(n3736) );
  NAND U4018 ( .A(n3676), .B(n3675), .Z(n3680) );
  NANDN U4019 ( .A(n3678), .B(n3677), .Z(n3679) );
  NAND U4020 ( .A(n3680), .B(n3679), .Z(n3742) );
  NAND U4021 ( .A(n3682), .B(n3681), .Z(n3686) );
  NANDN U4022 ( .A(n3684), .B(n3683), .Z(n3685) );
  NAND U4023 ( .A(n3686), .B(n3685), .Z(n3750) );
  AND U4024 ( .A(y[234]), .B(x[72]), .Z(n4925) );
  NAND U4025 ( .A(n4925), .B(n3855), .Z(n3690) );
  NANDN U4026 ( .A(n3688), .B(n3687), .Z(n3689) );
  AND U4027 ( .A(n3690), .B(n3689), .Z(n3781) );
  NAND U4028 ( .A(y[236]), .B(x[65]), .Z(n3691) );
  XNOR U4029 ( .A(n3692), .B(n3691), .Z(n3772) );
  ANDN U4030 ( .B(o[44]), .A(n3693), .Z(n3771) );
  XOR U4031 ( .A(n3772), .B(n3771), .Z(n3779) );
  AND U4032 ( .A(x[70]), .B(y[231]), .Z(n4723) );
  NAND U4033 ( .A(y[235]), .B(x[66]), .Z(n3694) );
  XOR U4034 ( .A(n3695), .B(n3694), .Z(n3784) );
  XNOR U4035 ( .A(n4723), .B(n3784), .Z(n3778) );
  XOR U4036 ( .A(n3779), .B(n3778), .Z(n3780) );
  XNOR U4037 ( .A(n3781), .B(n3780), .Z(n3749) );
  NAND U4038 ( .A(n3697), .B(n3696), .Z(n3701) );
  ANDN U4039 ( .B(n3699), .A(n3698), .Z(n3700) );
  ANDN U4040 ( .B(n3701), .A(n3700), .Z(n3748) );
  XOR U4041 ( .A(n3749), .B(n3748), .Z(n3751) );
  XOR U4042 ( .A(n3750), .B(n3751), .Z(n3743) );
  XOR U4043 ( .A(n3742), .B(n3743), .Z(n3745) );
  NANDN U4044 ( .A(n3703), .B(n3702), .Z(n3707) );
  NANDN U4045 ( .A(n3705), .B(n3704), .Z(n3706) );
  AND U4046 ( .A(n3707), .B(n3706), .Z(n3757) );
  NAND U4047 ( .A(x[70]), .B(y[235]), .Z(n4096) );
  NANDN U4048 ( .A(n4096), .B(n3770), .Z(n3711) );
  NAND U4049 ( .A(n3709), .B(n3708), .Z(n3710) );
  AND U4050 ( .A(n3711), .B(n3710), .Z(n3763) );
  AND U4051 ( .A(x[76]), .B(y[236]), .Z(n4931) );
  NAND U4052 ( .A(n4931), .B(n3902), .Z(n3715) );
  NAND U4053 ( .A(n3713), .B(n3712), .Z(n3714) );
  AND U4054 ( .A(n3715), .B(n3714), .Z(n3761) );
  AND U4055 ( .A(x[74]), .B(y[227]), .Z(n4587) );
  AND U4056 ( .A(y[229]), .B(x[72]), .Z(n3717) );
  NAND U4057 ( .A(y[226]), .B(x[75]), .Z(n3716) );
  XOR U4058 ( .A(n3717), .B(n3716), .Z(n3767) );
  XNOR U4059 ( .A(n4587), .B(n3767), .Z(n3760) );
  XNOR U4060 ( .A(n3761), .B(n3760), .Z(n3762) );
  XNOR U4061 ( .A(n3763), .B(n3762), .Z(n3755) );
  AND U4062 ( .A(x[74]), .B(y[232]), .Z(n4127) );
  AND U4063 ( .A(x[68]), .B(y[226]), .Z(n3718) );
  NAND U4064 ( .A(n4127), .B(n3718), .Z(n3721) );
  NANDN U4065 ( .A(n3719), .B(n4297), .Z(n3720) );
  AND U4066 ( .A(n3721), .B(n3720), .Z(n3805) );
  AND U4067 ( .A(y[224]), .B(x[77]), .Z(n3723) );
  NAND U4068 ( .A(y[237]), .B(x[64]), .Z(n3722) );
  XNOR U4069 ( .A(n3723), .B(n3722), .Z(n3797) );
  NAND U4070 ( .A(x[76]), .B(y[225]), .Z(n3789) );
  XNOR U4071 ( .A(o[45]), .B(n3789), .Z(n3796) );
  XOR U4072 ( .A(n3797), .B(n3796), .Z(n3803) );
  AND U4073 ( .A(y[234]), .B(x[67]), .Z(n3725) );
  NAND U4074 ( .A(y[232]), .B(x[69]), .Z(n3724) );
  XNOR U4075 ( .A(n3725), .B(n3724), .Z(n3792) );
  NAND U4076 ( .A(x[68]), .B(y[233]), .Z(n3793) );
  XNOR U4077 ( .A(n3792), .B(n3793), .Z(n3802) );
  XOR U4078 ( .A(n3803), .B(n3802), .Z(n3804) );
  XNOR U4079 ( .A(n3805), .B(n3804), .Z(n3754) );
  XOR U4080 ( .A(n3755), .B(n3754), .Z(n3756) );
  XNOR U4081 ( .A(n3757), .B(n3756), .Z(n3744) );
  XOR U4082 ( .A(n3745), .B(n3744), .Z(n3734) );
  NAND U4083 ( .A(n3727), .B(n3726), .Z(n3731) );
  NANDN U4084 ( .A(n3729), .B(n3728), .Z(n3730) );
  AND U4085 ( .A(n3731), .B(n3730), .Z(n3733) );
  XNOR U4086 ( .A(n3734), .B(n3733), .Z(n3735) );
  XNOR U4087 ( .A(n3736), .B(n3735), .Z(n3741) );
  XNOR U4088 ( .A(n3739), .B(n3741), .Z(n3732) );
  XOR U4089 ( .A(n3740), .B(n3732), .Z(N110) );
  NANDN U4090 ( .A(n3734), .B(n3733), .Z(n3738) );
  NANDN U4091 ( .A(n3736), .B(n3735), .Z(n3737) );
  NAND U4092 ( .A(n3738), .B(n3737), .Z(n3817) );
  IV U4093 ( .A(n3817), .Z(n3815) );
  NAND U4094 ( .A(n3743), .B(n3742), .Z(n3747) );
  NAND U4095 ( .A(n3745), .B(n3744), .Z(n3746) );
  NAND U4096 ( .A(n3747), .B(n3746), .Z(n3810) );
  NAND U4097 ( .A(n3749), .B(n3748), .Z(n3753) );
  NAND U4098 ( .A(n3751), .B(n3750), .Z(n3752) );
  NAND U4099 ( .A(n3753), .B(n3752), .Z(n3809) );
  XOR U4100 ( .A(n3810), .B(n3809), .Z(n3811) );
  NAND U4101 ( .A(n3755), .B(n3754), .Z(n3759) );
  NANDN U4102 ( .A(n3757), .B(n3756), .Z(n3758) );
  AND U4103 ( .A(n3759), .B(n3758), .Z(n3825) );
  NANDN U4104 ( .A(n3761), .B(n3760), .Z(n3765) );
  NANDN U4105 ( .A(n3763), .B(n3762), .Z(n3764) );
  AND U4106 ( .A(n3765), .B(n3764), .Z(n3831) );
  AND U4107 ( .A(x[75]), .B(y[229]), .Z(n3925) );
  NAND U4108 ( .A(n3925), .B(n3766), .Z(n3769) );
  NANDN U4109 ( .A(n3767), .B(n4587), .Z(n3768) );
  AND U4110 ( .A(n3769), .B(n3768), .Z(n3885) );
  NAND U4111 ( .A(x[71]), .B(y[236]), .Z(n4312) );
  NANDN U4112 ( .A(n4312), .B(n3770), .Z(n3774) );
  NAND U4113 ( .A(n3772), .B(n3771), .Z(n3773) );
  NAND U4114 ( .A(n3774), .B(n3773), .Z(n3884) );
  XNOR U4115 ( .A(n3885), .B(n3884), .Z(n3887) );
  AND U4116 ( .A(x[68]), .B(y[234]), .Z(n4235) );
  AND U4117 ( .A(y[230]), .B(x[72]), .Z(n3776) );
  NAND U4118 ( .A(y[235]), .B(x[67]), .Z(n3775) );
  XOR U4119 ( .A(n3776), .B(n3775), .Z(n3870) );
  XNOR U4120 ( .A(n4094), .B(n3870), .Z(n3879) );
  XOR U4121 ( .A(n4235), .B(n3879), .Z(n3881) );
  AND U4122 ( .A(x[73]), .B(y[229]), .Z(n4404) );
  AND U4123 ( .A(y[228]), .B(x[74]), .Z(n4434) );
  AND U4124 ( .A(y[236]), .B(x[66]), .Z(n3777) );
  XOR U4125 ( .A(n4434), .B(n3777), .Z(n3856) );
  XOR U4126 ( .A(n4404), .B(n3856), .Z(n3880) );
  XOR U4127 ( .A(n3881), .B(n3880), .Z(n3886) );
  XOR U4128 ( .A(n3887), .B(n3886), .Z(n3829) );
  NAND U4129 ( .A(n3779), .B(n3778), .Z(n3783) );
  NANDN U4130 ( .A(n3781), .B(n3780), .Z(n3782) );
  AND U4131 ( .A(n3783), .B(n3782), .Z(n3828) );
  XNOR U4132 ( .A(n3829), .B(n3828), .Z(n3830) );
  XOR U4133 ( .A(n3831), .B(n3830), .Z(n3823) );
  AND U4134 ( .A(x[73]), .B(y[235]), .Z(n4310) );
  NAND U4135 ( .A(n4310), .B(n3855), .Z(n3786) );
  NANDN U4136 ( .A(n3784), .B(n4723), .Z(n3785) );
  AND U4137 ( .A(n3786), .B(n3785), .Z(n3843) );
  AND U4138 ( .A(y[238]), .B(x[64]), .Z(n3788) );
  NAND U4139 ( .A(y[224]), .B(x[78]), .Z(n3787) );
  XNOR U4140 ( .A(n3788), .B(n3787), .Z(n3866) );
  ANDN U4141 ( .B(o[45]), .A(n3789), .Z(n3865) );
  XOR U4142 ( .A(n3866), .B(n3865), .Z(n3841) );
  NAND U4143 ( .A(y[226]), .B(x[76]), .Z(n3790) );
  XNOR U4144 ( .A(n3791), .B(n3790), .Z(n3848) );
  NAND U4145 ( .A(x[77]), .B(y[225]), .Z(n3854) );
  XNOR U4146 ( .A(o[46]), .B(n3854), .Z(n3847) );
  XOR U4147 ( .A(n3848), .B(n3847), .Z(n3840) );
  XOR U4148 ( .A(n3841), .B(n3840), .Z(n3842) );
  XOR U4149 ( .A(n3843), .B(n3842), .Z(n3891) );
  NAND U4150 ( .A(x[69]), .B(y[234]), .Z(n3914) );
  NANDN U4151 ( .A(n3914), .B(n4575), .Z(n3795) );
  NANDN U4152 ( .A(n3793), .B(n3792), .Z(n3794) );
  AND U4153 ( .A(n3795), .B(n3794), .Z(n3837) );
  AND U4154 ( .A(x[77]), .B(y[237]), .Z(n5295) );
  NAND U4155 ( .A(n5295), .B(n3902), .Z(n3799) );
  NAND U4156 ( .A(n3797), .B(n3796), .Z(n3798) );
  AND U4157 ( .A(n3799), .B(n3798), .Z(n3835) );
  NAND U4158 ( .A(y[227]), .B(x[75]), .Z(n3800) );
  XNOR U4159 ( .A(n3801), .B(n3800), .Z(n3861) );
  NAND U4160 ( .A(x[65]), .B(y[237]), .Z(n3862) );
  XNOR U4161 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U4162 ( .A(n3837), .B(n3836), .Z(n3890) );
  XOR U4163 ( .A(n3891), .B(n3890), .Z(n3893) );
  NAND U4164 ( .A(n3803), .B(n3802), .Z(n3807) );
  NANDN U4165 ( .A(n3805), .B(n3804), .Z(n3806) );
  AND U4166 ( .A(n3807), .B(n3806), .Z(n3892) );
  XNOR U4167 ( .A(n3893), .B(n3892), .Z(n3822) );
  XNOR U4168 ( .A(n3823), .B(n3822), .Z(n3824) );
  XOR U4169 ( .A(n3825), .B(n3824), .Z(n3812) );
  XNOR U4170 ( .A(n3811), .B(n3812), .Z(n3818) );
  XNOR U4171 ( .A(n3816), .B(n3818), .Z(n3808) );
  XOR U4172 ( .A(n3815), .B(n3808), .Z(N111) );
  NAND U4173 ( .A(n3810), .B(n3809), .Z(n3814) );
  NANDN U4174 ( .A(n3812), .B(n3811), .Z(n3813) );
  AND U4175 ( .A(n3814), .B(n3813), .Z(n3982) );
  NANDN U4176 ( .A(n3815), .B(n3816), .Z(n3821) );
  NOR U4177 ( .A(n3817), .B(n3816), .Z(n3819) );
  OR U4178 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U4179 ( .A(n3821), .B(n3820), .Z(n3983) );
  NANDN U4180 ( .A(n3823), .B(n3822), .Z(n3827) );
  NANDN U4181 ( .A(n3825), .B(n3824), .Z(n3826) );
  AND U4182 ( .A(n3827), .B(n3826), .Z(n3979) );
  NANDN U4183 ( .A(n3829), .B(n3828), .Z(n3833) );
  NAND U4184 ( .A(n3831), .B(n3830), .Z(n3832) );
  NAND U4185 ( .A(n3833), .B(n3832), .Z(n3954) );
  NANDN U4186 ( .A(n3835), .B(n3834), .Z(n3839) );
  NANDN U4187 ( .A(n3837), .B(n3836), .Z(n3838) );
  AND U4188 ( .A(n3839), .B(n3838), .Z(n3961) );
  NAND U4189 ( .A(n3841), .B(n3840), .Z(n3845) );
  NANDN U4190 ( .A(n3843), .B(n3842), .Z(n3844) );
  AND U4191 ( .A(n3845), .B(n3844), .Z(n3959) );
  NAND U4192 ( .A(x[76]), .B(y[231]), .Z(n4304) );
  NANDN U4193 ( .A(n4304), .B(n3846), .Z(n3850) );
  NAND U4194 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4195 ( .A(n3850), .B(n3849), .Z(n3935) );
  AND U4196 ( .A(y[226]), .B(x[77]), .Z(n4711) );
  NAND U4197 ( .A(y[228]), .B(x[75]), .Z(n3851) );
  XNOR U4198 ( .A(n4711), .B(n3851), .Z(n3939) );
  AND U4199 ( .A(x[76]), .B(y[227]), .Z(n3938) );
  XOR U4200 ( .A(n3939), .B(n3938), .Z(n3933) );
  AND U4201 ( .A(y[224]), .B(x[79]), .Z(n3853) );
  NAND U4202 ( .A(y[239]), .B(x[64]), .Z(n3852) );
  XNOR U4203 ( .A(n3853), .B(n3852), .Z(n3904) );
  ANDN U4204 ( .B(o[46]), .A(n3854), .Z(n3903) );
  XNOR U4205 ( .A(n3904), .B(n3903), .Z(n3932) );
  XNOR U4206 ( .A(n3933), .B(n3932), .Z(n3934) );
  XOR U4207 ( .A(n3935), .B(n3934), .Z(n3967) );
  AND U4208 ( .A(x[74]), .B(y[236]), .Z(n4724) );
  NAND U4209 ( .A(n4724), .B(n3855), .Z(n3858) );
  NAND U4210 ( .A(n4404), .B(n3856), .Z(n3857) );
  AND U4211 ( .A(n3858), .B(n3857), .Z(n3965) );
  AND U4212 ( .A(x[75]), .B(y[232]), .Z(n3860) );
  NAND U4213 ( .A(n3860), .B(n3859), .Z(n3864) );
  NANDN U4214 ( .A(n3862), .B(n3861), .Z(n3863) );
  NAND U4215 ( .A(n3864), .B(n3863), .Z(n3964) );
  AND U4216 ( .A(x[78]), .B(y[238]), .Z(n5557) );
  NAND U4217 ( .A(n3902), .B(n5557), .Z(n3868) );
  NAND U4218 ( .A(n3866), .B(n3865), .Z(n3867) );
  AND U4219 ( .A(n3868), .B(n3867), .Z(n3927) );
  AND U4220 ( .A(x[72]), .B(y[235]), .Z(n4210) );
  NANDN U4221 ( .A(n3869), .B(n4210), .Z(n3872) );
  NANDN U4222 ( .A(n3870), .B(n4094), .Z(n3871) );
  NAND U4223 ( .A(n3872), .B(n3871), .Z(n3926) );
  XNOR U4224 ( .A(n3927), .B(n3926), .Z(n3929) );
  AND U4225 ( .A(y[229]), .B(x[74]), .Z(n3874) );
  NAND U4226 ( .A(y[235]), .B(x[68]), .Z(n3873) );
  XNOR U4227 ( .A(n3874), .B(n3873), .Z(n3909) );
  AND U4228 ( .A(x[71]), .B(y[232]), .Z(n3908) );
  XOR U4229 ( .A(n3909), .B(n3908), .Z(n3916) );
  NAND U4230 ( .A(x[70]), .B(y[233]), .Z(n4013) );
  XOR U4231 ( .A(n4013), .B(n3914), .Z(n3915) );
  XNOR U4232 ( .A(n3916), .B(n3915), .Z(n3949) );
  AND U4233 ( .A(y[230]), .B(x[73]), .Z(n3876) );
  NAND U4234 ( .A(y[237]), .B(x[66]), .Z(n3875) );
  XNOR U4235 ( .A(n3876), .B(n3875), .Z(n3917) );
  NAND U4236 ( .A(x[67]), .B(y[236]), .Z(n3918) );
  XNOR U4237 ( .A(n3917), .B(n3918), .Z(n3947) );
  AND U4238 ( .A(y[231]), .B(x[72]), .Z(n3878) );
  NAND U4239 ( .A(y[238]), .B(x[65]), .Z(n3877) );
  XNOR U4240 ( .A(n3878), .B(n3877), .Z(n3899) );
  NAND U4241 ( .A(x[78]), .B(y[225]), .Z(n3923) );
  XNOR U4242 ( .A(o[47]), .B(n3923), .Z(n3898) );
  XOR U4243 ( .A(n3899), .B(n3898), .Z(n3946) );
  XOR U4244 ( .A(n3947), .B(n3946), .Z(n3948) );
  XNOR U4245 ( .A(n3949), .B(n3948), .Z(n3928) );
  XOR U4246 ( .A(n3929), .B(n3928), .Z(n3971) );
  NAND U4247 ( .A(n4235), .B(n3879), .Z(n3883) );
  NAND U4248 ( .A(n3881), .B(n3880), .Z(n3882) );
  AND U4249 ( .A(n3883), .B(n3882), .Z(n3970) );
  NANDN U4250 ( .A(n3885), .B(n3884), .Z(n3889) );
  NAND U4251 ( .A(n3887), .B(n3886), .Z(n3888) );
  AND U4252 ( .A(n3889), .B(n3888), .Z(n3972) );
  XOR U4253 ( .A(n3973), .B(n3972), .Z(n3952) );
  XOR U4254 ( .A(n3953), .B(n3952), .Z(n3955) );
  XOR U4255 ( .A(n3954), .B(n3955), .Z(n3976) );
  NAND U4256 ( .A(n3891), .B(n3890), .Z(n3895) );
  NAND U4257 ( .A(n3893), .B(n3892), .Z(n3894) );
  AND U4258 ( .A(n3895), .B(n3894), .Z(n3977) );
  XOR U4259 ( .A(n3976), .B(n3977), .Z(n3978) );
  XNOR U4260 ( .A(n3979), .B(n3978), .Z(n3984) );
  XNOR U4261 ( .A(n3983), .B(n3984), .Z(n3896) );
  XOR U4262 ( .A(n3982), .B(n3896), .Z(N112) );
  AND U4263 ( .A(x[72]), .B(y[238]), .Z(n4596) );
  NAND U4264 ( .A(n4596), .B(n3897), .Z(n3901) );
  NAND U4265 ( .A(n3899), .B(n3898), .Z(n3900) );
  AND U4266 ( .A(n3901), .B(n3900), .Z(n4043) );
  AND U4267 ( .A(x[79]), .B(y[239]), .Z(n6012) );
  NAND U4268 ( .A(n6012), .B(n3902), .Z(n3906) );
  NAND U4269 ( .A(n3904), .B(n3903), .Z(n3905) );
  NAND U4270 ( .A(n3906), .B(n3905), .Z(n4042) );
  XNOR U4271 ( .A(n4043), .B(n4042), .Z(n4045) );
  AND U4272 ( .A(x[74]), .B(y[235]), .Z(n4447) );
  NAND U4273 ( .A(n4447), .B(n3907), .Z(n3911) );
  NAND U4274 ( .A(n3909), .B(n3908), .Z(n3910) );
  NAND U4275 ( .A(n3911), .B(n3910), .Z(n4000) );
  AND U4276 ( .A(x[64]), .B(y[240]), .Z(n4022) );
  NAND U4277 ( .A(x[80]), .B(y[224]), .Z(n4023) );
  XNOR U4278 ( .A(n4022), .B(n4023), .Z(n4024) );
  NAND U4279 ( .A(x[79]), .B(y[225]), .Z(n4010) );
  XOR U4280 ( .A(o[48]), .B(n4010), .Z(n4025) );
  XNOR U4281 ( .A(n4024), .B(n4025), .Z(n3999) );
  NAND U4282 ( .A(y[233]), .B(x[71]), .Z(n3912) );
  XNOR U4283 ( .A(n3913), .B(n3912), .Z(n4015) );
  AND U4284 ( .A(x[74]), .B(y[230]), .Z(n4014) );
  XOR U4285 ( .A(n4015), .B(n4014), .Z(n3998) );
  XOR U4286 ( .A(n3999), .B(n3998), .Z(n4001) );
  XOR U4287 ( .A(n4000), .B(n4001), .Z(n4044) );
  XOR U4288 ( .A(n4045), .B(n4044), .Z(n3995) );
  AND U4289 ( .A(x[73]), .B(y[237]), .Z(n4706) );
  NAND U4290 ( .A(n4706), .B(n4302), .Z(n3920) );
  NANDN U4291 ( .A(n3918), .B(n3917), .Z(n3919) );
  NAND U4292 ( .A(n3920), .B(n3919), .Z(n4032) );
  NAND U4293 ( .A(y[239]), .B(x[65]), .Z(n3921) );
  XNOR U4294 ( .A(n3922), .B(n3921), .Z(n4019) );
  ANDN U4295 ( .B(o[47]), .A(n3923), .Z(n4018) );
  XOR U4296 ( .A(n4019), .B(n4018), .Z(n4031) );
  NAND U4297 ( .A(y[226]), .B(x[78]), .Z(n3924) );
  XNOR U4298 ( .A(n3925), .B(n3924), .Z(n4054) );
  NAND U4299 ( .A(x[68]), .B(y[236]), .Z(n4055) );
  XNOR U4300 ( .A(n4054), .B(n4055), .Z(n4030) );
  XOR U4301 ( .A(n4031), .B(n4030), .Z(n4033) );
  XNOR U4302 ( .A(n4032), .B(n4033), .Z(n3992) );
  XNOR U4303 ( .A(n3993), .B(n3992), .Z(n3994) );
  XNOR U4304 ( .A(n3995), .B(n3994), .Z(n4036) );
  NANDN U4305 ( .A(n3927), .B(n3926), .Z(n3931) );
  NAND U4306 ( .A(n3929), .B(n3928), .Z(n3930) );
  NAND U4307 ( .A(n3931), .B(n3930), .Z(n4037) );
  XNOR U4308 ( .A(n4036), .B(n4037), .Z(n4039) );
  NANDN U4309 ( .A(n3933), .B(n3932), .Z(n3937) );
  NAND U4310 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U4311 ( .A(n3937), .B(n3936), .Z(n4068) );
  AND U4312 ( .A(x[75]), .B(y[226]), .Z(n4548) );
  AND U4313 ( .A(x[77]), .B(y[228]), .Z(n4065) );
  NAND U4314 ( .A(n4548), .B(n4065), .Z(n3941) );
  NAND U4315 ( .A(n3939), .B(n3938), .Z(n3940) );
  AND U4316 ( .A(n3941), .B(n3940), .Z(n4051) );
  AND U4317 ( .A(y[231]), .B(x[73]), .Z(n3943) );
  NAND U4318 ( .A(y[238]), .B(x[66]), .Z(n3942) );
  XNOR U4319 ( .A(n3943), .B(n3942), .Z(n4058) );
  NAND U4320 ( .A(x[67]), .B(y[237]), .Z(n4059) );
  XNOR U4321 ( .A(n4058), .B(n4059), .Z(n4049) );
  AND U4322 ( .A(x[76]), .B(y[228]), .Z(n4695) );
  AND U4323 ( .A(y[227]), .B(x[77]), .Z(n3945) );
  NAND U4324 ( .A(y[235]), .B(x[69]), .Z(n3944) );
  XOR U4325 ( .A(n3945), .B(n3944), .Z(n4005) );
  XNOR U4326 ( .A(n4695), .B(n4005), .Z(n4048) );
  XOR U4327 ( .A(n4049), .B(n4048), .Z(n4050) );
  XNOR U4328 ( .A(n4051), .B(n4050), .Z(n4067) );
  NAND U4329 ( .A(n3947), .B(n3946), .Z(n3951) );
  NANDN U4330 ( .A(n3949), .B(n3948), .Z(n3950) );
  AND U4331 ( .A(n3951), .B(n3950), .Z(n4066) );
  XNOR U4332 ( .A(n4067), .B(n4066), .Z(n4069) );
  XOR U4333 ( .A(n4068), .B(n4069), .Z(n4038) );
  XOR U4334 ( .A(n4039), .B(n4038), .Z(n4076) );
  NANDN U4335 ( .A(n3953), .B(n3952), .Z(n3957) );
  NANDN U4336 ( .A(n3955), .B(n3954), .Z(n3956) );
  AND U4337 ( .A(n3957), .B(n3956), .Z(n4075) );
  XNOR U4338 ( .A(n4076), .B(n4075), .Z(n4078) );
  NANDN U4339 ( .A(n3959), .B(n3958), .Z(n3963) );
  NANDN U4340 ( .A(n3961), .B(n3960), .Z(n3962) );
  AND U4341 ( .A(n3963), .B(n3962), .Z(n3989) );
  NANDN U4342 ( .A(n3965), .B(n3964), .Z(n3969) );
  NANDN U4343 ( .A(n3967), .B(n3966), .Z(n3968) );
  AND U4344 ( .A(n3969), .B(n3968), .Z(n3987) );
  NANDN U4345 ( .A(n3971), .B(n3970), .Z(n3975) );
  NAND U4346 ( .A(n3973), .B(n3972), .Z(n3974) );
  AND U4347 ( .A(n3975), .B(n3974), .Z(n3986) );
  XNOR U4348 ( .A(n4078), .B(n4077), .Z(n4074) );
  NAND U4349 ( .A(n3977), .B(n3976), .Z(n3981) );
  NANDN U4350 ( .A(n3979), .B(n3978), .Z(n3980) );
  NAND U4351 ( .A(n3981), .B(n3980), .Z(n4073) );
  XOR U4352 ( .A(n4073), .B(n4072), .Z(n3985) );
  XNOR U4353 ( .A(n4074), .B(n3985), .Z(N113) );
  NANDN U4354 ( .A(n3987), .B(n3986), .Z(n3991) );
  NANDN U4355 ( .A(n3989), .B(n3988), .Z(n3990) );
  AND U4356 ( .A(n3991), .B(n3990), .Z(n4175) );
  NANDN U4357 ( .A(n3993), .B(n3992), .Z(n3997) );
  NANDN U4358 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U4359 ( .A(n3997), .B(n3996), .Z(n4090) );
  NAND U4360 ( .A(n3999), .B(n3998), .Z(n4003) );
  NAND U4361 ( .A(n4001), .B(n4000), .Z(n4002) );
  AND U4362 ( .A(n4003), .B(n4002), .Z(n4169) );
  AND U4363 ( .A(x[77]), .B(y[235]), .Z(n4939) );
  AND U4364 ( .A(x[69]), .B(y[227]), .Z(n4004) );
  NAND U4365 ( .A(n4939), .B(n4004), .Z(n4007) );
  NANDN U4366 ( .A(n4005), .B(n4695), .Z(n4006) );
  AND U4367 ( .A(n4007), .B(n4006), .Z(n4145) );
  AND U4368 ( .A(y[232]), .B(x[73]), .Z(n4009) );
  NAND U4369 ( .A(y[240]), .B(x[65]), .Z(n4008) );
  XNOR U4370 ( .A(n4009), .B(n4008), .Z(n4100) );
  ANDN U4371 ( .B(o[48]), .A(n4010), .Z(n4099) );
  XOR U4372 ( .A(n4100), .B(n4099), .Z(n4143) );
  AND U4373 ( .A(y[226]), .B(x[79]), .Z(n4012) );
  NAND U4374 ( .A(y[229]), .B(x[76]), .Z(n4011) );
  XNOR U4375 ( .A(n4012), .B(n4011), .Z(n4118) );
  AND U4376 ( .A(x[78]), .B(y[227]), .Z(n4117) );
  XOR U4377 ( .A(n4118), .B(n4117), .Z(n4142) );
  XOR U4378 ( .A(n4143), .B(n4142), .Z(n4144) );
  XNOR U4379 ( .A(n4145), .B(n4144), .Z(n4167) );
  AND U4380 ( .A(x[71]), .B(y[234]), .Z(n4107) );
  NANDN U4381 ( .A(n4013), .B(n4107), .Z(n4017) );
  NAND U4382 ( .A(n4015), .B(n4014), .Z(n4016) );
  AND U4383 ( .A(n4017), .B(n4016), .Z(n4155) );
  AND U4384 ( .A(x[72]), .B(y[239]), .Z(n4851) );
  AND U4385 ( .A(x[65]), .B(y[232]), .Z(n4213) );
  NAND U4386 ( .A(n4851), .B(n4213), .Z(n4021) );
  NAND U4387 ( .A(n4019), .B(n4018), .Z(n4020) );
  NAND U4388 ( .A(n4021), .B(n4020), .Z(n4154) );
  XNOR U4389 ( .A(n4155), .B(n4154), .Z(n4157) );
  NANDN U4390 ( .A(n4023), .B(n4022), .Z(n4027) );
  NANDN U4391 ( .A(n4025), .B(n4024), .Z(n4026) );
  AND U4392 ( .A(n4027), .B(n4026), .Z(n4151) );
  AND U4393 ( .A(x[64]), .B(y[241]), .Z(n4132) );
  AND U4394 ( .A(x[81]), .B(y[224]), .Z(n4131) );
  XOR U4395 ( .A(n4132), .B(n4131), .Z(n4134) );
  AND U4396 ( .A(x[80]), .B(y[225]), .Z(n4128) );
  XOR U4397 ( .A(n4128), .B(o[49]), .Z(n4133) );
  XOR U4398 ( .A(n4134), .B(n4133), .Z(n4149) );
  AND U4399 ( .A(y[231]), .B(x[74]), .Z(n4029) );
  NAND U4400 ( .A(y[239]), .B(x[66]), .Z(n4028) );
  XNOR U4401 ( .A(n4029), .B(n4028), .Z(n4103) );
  AND U4402 ( .A(x[67]), .B(y[238]), .Z(n4102) );
  XOR U4403 ( .A(n4103), .B(n4102), .Z(n4148) );
  XOR U4404 ( .A(n4149), .B(n4148), .Z(n4150) );
  XNOR U4405 ( .A(n4151), .B(n4150), .Z(n4156) );
  XOR U4406 ( .A(n4157), .B(n4156), .Z(n4166) );
  XOR U4407 ( .A(n4167), .B(n4166), .Z(n4168) );
  XNOR U4408 ( .A(n4169), .B(n4168), .Z(n4089) );
  NAND U4409 ( .A(n4031), .B(n4030), .Z(n4035) );
  NAND U4410 ( .A(n4033), .B(n4032), .Z(n4034) );
  AND U4411 ( .A(n4035), .B(n4034), .Z(n4088) );
  XOR U4412 ( .A(n4089), .B(n4088), .Z(n4091) );
  XOR U4413 ( .A(n4090), .B(n4091), .Z(n4173) );
  NANDN U4414 ( .A(n4037), .B(n4036), .Z(n4041) );
  NAND U4415 ( .A(n4039), .B(n4038), .Z(n4040) );
  NAND U4416 ( .A(n4041), .B(n4040), .Z(n4084) );
  NANDN U4417 ( .A(n4043), .B(n4042), .Z(n4047) );
  NAND U4418 ( .A(n4045), .B(n4044), .Z(n4046) );
  AND U4419 ( .A(n4047), .B(n4046), .Z(n4163) );
  NAND U4420 ( .A(n4049), .B(n4048), .Z(n4053) );
  NANDN U4421 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U4422 ( .A(n4053), .B(n4052), .Z(n4161) );
  NAND U4423 ( .A(x[78]), .B(y[229]), .Z(n4336) );
  NANDN U4424 ( .A(n4336), .B(n4548), .Z(n4057) );
  NANDN U4425 ( .A(n4055), .B(n4054), .Z(n4056) );
  AND U4426 ( .A(n4057), .B(n4056), .Z(n4111) );
  AND U4427 ( .A(y[238]), .B(x[73]), .Z(n4920) );
  NAND U4428 ( .A(n4101), .B(n4920), .Z(n4061) );
  NANDN U4429 ( .A(n4059), .B(n4058), .Z(n4060) );
  NAND U4430 ( .A(n4061), .B(n4060), .Z(n4110) );
  XNOR U4431 ( .A(n4111), .B(n4110), .Z(n4112) );
  AND U4432 ( .A(y[233]), .B(x[72]), .Z(n4063) );
  NAND U4433 ( .A(y[236]), .B(x[69]), .Z(n4062) );
  XNOR U4434 ( .A(n4063), .B(n4062), .Z(n4095) );
  XOR U4435 ( .A(n4107), .B(n4106), .Z(n4108) );
  NAND U4436 ( .A(y[237]), .B(x[68]), .Z(n4064) );
  XNOR U4437 ( .A(n4065), .B(n4064), .Z(n4122) );
  NAND U4438 ( .A(x[75]), .B(y[230]), .Z(n4123) );
  XOR U4439 ( .A(n4122), .B(n4123), .Z(n4109) );
  XOR U4440 ( .A(n4108), .B(n4109), .Z(n4113) );
  XNOR U4441 ( .A(n4112), .B(n4113), .Z(n4160) );
  XNOR U4442 ( .A(n4161), .B(n4160), .Z(n4162) );
  XNOR U4443 ( .A(n4163), .B(n4162), .Z(n4083) );
  NANDN U4444 ( .A(n4067), .B(n4066), .Z(n4071) );
  NAND U4445 ( .A(n4069), .B(n4068), .Z(n4070) );
  NAND U4446 ( .A(n4071), .B(n4070), .Z(n4082) );
  XOR U4447 ( .A(n4083), .B(n4082), .Z(n4085) );
  XOR U4448 ( .A(n4084), .B(n4085), .Z(n4172) );
  XOR U4449 ( .A(n4173), .B(n4172), .Z(n4174) );
  XOR U4450 ( .A(n4175), .B(n4174), .Z(n4180) );
  NANDN U4451 ( .A(n4076), .B(n4075), .Z(n4080) );
  NAND U4452 ( .A(n4078), .B(n4077), .Z(n4079) );
  NAND U4453 ( .A(n4080), .B(n4079), .Z(n4178) );
  XNOR U4454 ( .A(n4179), .B(n4178), .Z(n4081) );
  XNOR U4455 ( .A(n4180), .B(n4081), .Z(N114) );
  NANDN U4456 ( .A(n4083), .B(n4082), .Z(n4087) );
  NANDN U4457 ( .A(n4085), .B(n4084), .Z(n4086) );
  AND U4458 ( .A(n4087), .B(n4086), .Z(n4281) );
  NANDN U4459 ( .A(n4089), .B(n4088), .Z(n4093) );
  NANDN U4460 ( .A(n4091), .B(n4090), .Z(n4092) );
  AND U4461 ( .A(n4093), .B(n4092), .Z(n4278) );
  AND U4462 ( .A(x[72]), .B(y[236]), .Z(n4440) );
  NAND U4463 ( .A(n4440), .B(n4094), .Z(n4098) );
  NANDN U4464 ( .A(n4096), .B(n4095), .Z(n4097) );
  NAND U4465 ( .A(n4098), .B(n4097), .Z(n4264) );
  AND U4466 ( .A(x[73]), .B(y[240]), .Z(n5093) );
  XOR U4467 ( .A(n4264), .B(n4263), .Z(n4265) );
  AND U4468 ( .A(x[74]), .B(y[239]), .Z(n4948) );
  IV U4469 ( .A(n4948), .Z(n5092) );
  AND U4470 ( .A(x[64]), .B(y[242]), .Z(n4218) );
  NAND U4471 ( .A(x[82]), .B(y[224]), .Z(n4219) );
  XNOR U4472 ( .A(n4218), .B(n4219), .Z(n4220) );
  NAND U4473 ( .A(x[81]), .B(y[225]), .Z(n4240) );
  XOR U4474 ( .A(o[50]), .B(n4240), .Z(n4221) );
  XNOR U4475 ( .A(n4220), .B(n4221), .Z(n4244) );
  AND U4476 ( .A(y[229]), .B(x[77]), .Z(n4105) );
  NAND U4477 ( .A(y[239]), .B(x[67]), .Z(n4104) );
  XNOR U4478 ( .A(n4105), .B(n4104), .Z(n4227) );
  NAND U4479 ( .A(x[76]), .B(y[230]), .Z(n4228) );
  XNOR U4480 ( .A(n4227), .B(n4228), .Z(n4243) );
  XOR U4481 ( .A(n4244), .B(n4243), .Z(n4245) );
  XNOR U4482 ( .A(n4246), .B(n4245), .Z(n4266) );
  XNOR U4483 ( .A(n4265), .B(n4266), .Z(n4195) );
  XNOR U4484 ( .A(n4195), .B(n4194), .Z(n4197) );
  NANDN U4485 ( .A(n4111), .B(n4110), .Z(n4115) );
  NANDN U4486 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U4487 ( .A(n4115), .B(n4114), .Z(n4196) );
  XOR U4488 ( .A(n4197), .B(n4196), .Z(n4191) );
  AND U4489 ( .A(x[79]), .B(y[229]), .Z(n4116) );
  AND U4490 ( .A(x[76]), .B(y[226]), .Z(n4394) );
  NAND U4491 ( .A(n4116), .B(n4394), .Z(n4120) );
  NAND U4492 ( .A(n4118), .B(n4117), .Z(n4119) );
  NAND U4493 ( .A(n4120), .B(n4119), .Z(n4257) );
  NAND U4494 ( .A(n5295), .B(n4121), .Z(n4125) );
  NANDN U4495 ( .A(n4123), .B(n4122), .Z(n4124) );
  NAND U4496 ( .A(n4125), .B(n4124), .Z(n4249) );
  NAND U4497 ( .A(y[241]), .B(x[65]), .Z(n4126) );
  XNOR U4498 ( .A(n4127), .B(n4126), .Z(n4214) );
  NAND U4499 ( .A(n4128), .B(o[49]), .Z(n4215) );
  XNOR U4500 ( .A(n4214), .B(n4215), .Z(n4248) );
  NAND U4501 ( .A(y[227]), .B(x[79]), .Z(n4129) );
  XNOR U4502 ( .A(n4130), .B(n4129), .Z(n4206) );
  AND U4503 ( .A(x[78]), .B(y[228]), .Z(n4205) );
  XOR U4504 ( .A(n4206), .B(n4205), .Z(n4247) );
  XOR U4505 ( .A(n4248), .B(n4247), .Z(n4250) );
  XOR U4506 ( .A(n4249), .B(n4250), .Z(n4258) );
  XOR U4507 ( .A(n4257), .B(n4258), .Z(n4260) );
  NAND U4508 ( .A(n4132), .B(n4131), .Z(n4136) );
  NAND U4509 ( .A(n4134), .B(n4133), .Z(n4135) );
  NAND U4510 ( .A(n4136), .B(n4135), .Z(n4269) );
  AND U4511 ( .A(y[231]), .B(x[75]), .Z(n4138) );
  NAND U4512 ( .A(y[226]), .B(x[80]), .Z(n4137) );
  XNOR U4513 ( .A(n4138), .B(n4137), .Z(n4204) );
  AND U4514 ( .A(x[66]), .B(y[240]), .Z(n4203) );
  XOR U4515 ( .A(n4204), .B(n4203), .Z(n4270) );
  XOR U4516 ( .A(n4269), .B(n4270), .Z(n4272) );
  AND U4517 ( .A(y[236]), .B(x[70]), .Z(n4140) );
  NAND U4518 ( .A(y[237]), .B(x[69]), .Z(n4139) );
  XNOR U4519 ( .A(n4140), .B(n4139), .Z(n4200) );
  NAND U4520 ( .A(y[238]), .B(x[68]), .Z(n4141) );
  XNOR U4521 ( .A(n4925), .B(n4141), .Z(n4236) );
  NAND U4522 ( .A(x[71]), .B(y[235]), .Z(n4237) );
  XNOR U4523 ( .A(n4236), .B(n4237), .Z(n4199) );
  XOR U4524 ( .A(n4200), .B(n4199), .Z(n4271) );
  XOR U4525 ( .A(n4272), .B(n4271), .Z(n4259) );
  XOR U4526 ( .A(n4260), .B(n4259), .Z(n4189) );
  NAND U4527 ( .A(n4143), .B(n4142), .Z(n4147) );
  NANDN U4528 ( .A(n4145), .B(n4144), .Z(n4146) );
  AND U4529 ( .A(n4147), .B(n4146), .Z(n4252) );
  NAND U4530 ( .A(n4149), .B(n4148), .Z(n4153) );
  NANDN U4531 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U4532 ( .A(n4153), .B(n4152), .Z(n4251) );
  XOR U4533 ( .A(n4252), .B(n4251), .Z(n4254) );
  NANDN U4534 ( .A(n4155), .B(n4154), .Z(n4159) );
  NAND U4535 ( .A(n4157), .B(n4156), .Z(n4158) );
  AND U4536 ( .A(n4159), .B(n4158), .Z(n4253) );
  XOR U4537 ( .A(n4254), .B(n4253), .Z(n4188) );
  XOR U4538 ( .A(n4191), .B(n4190), .Z(n4185) );
  NANDN U4539 ( .A(n4161), .B(n4160), .Z(n4165) );
  NANDN U4540 ( .A(n4163), .B(n4162), .Z(n4164) );
  AND U4541 ( .A(n4165), .B(n4164), .Z(n4183) );
  NAND U4542 ( .A(n4167), .B(n4166), .Z(n4171) );
  NANDN U4543 ( .A(n4169), .B(n4168), .Z(n4170) );
  NAND U4544 ( .A(n4171), .B(n4170), .Z(n4182) );
  XNOR U4545 ( .A(n4278), .B(n4279), .Z(n4280) );
  XNOR U4546 ( .A(n4281), .B(n4280), .Z(n4277) );
  NAND U4547 ( .A(n4173), .B(n4172), .Z(n4177) );
  NANDN U4548 ( .A(n4175), .B(n4174), .Z(n4176) );
  NAND U4549 ( .A(n4177), .B(n4176), .Z(n4275) );
  XOR U4550 ( .A(n4275), .B(n4276), .Z(n4181) );
  XNOR U4551 ( .A(n4277), .B(n4181), .Z(N115) );
  NANDN U4552 ( .A(n4183), .B(n4182), .Z(n4187) );
  NANDN U4553 ( .A(n4185), .B(n4184), .Z(n4186) );
  AND U4554 ( .A(n4187), .B(n4186), .Z(n4381) );
  NANDN U4555 ( .A(n4189), .B(n4188), .Z(n4193) );
  NAND U4556 ( .A(n4191), .B(n4190), .Z(n4192) );
  AND U4557 ( .A(n4193), .B(n4192), .Z(n4379) );
  AND U4558 ( .A(x[70]), .B(y[237]), .Z(n4242) );
  AND U4559 ( .A(x[69]), .B(y[236]), .Z(n4198) );
  NAND U4560 ( .A(n4242), .B(n4198), .Z(n4202) );
  NAND U4561 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U4562 ( .A(n4202), .B(n4201), .Z(n4356) );
  AND U4563 ( .A(x[79]), .B(y[233]), .Z(n4951) );
  NAND U4564 ( .A(n4951), .B(n4297), .Z(n4208) );
  NAND U4565 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U4566 ( .A(n4208), .B(n4207), .Z(n4292) );
  NAND U4567 ( .A(y[242]), .B(x[65]), .Z(n4209) );
  XNOR U4568 ( .A(n4210), .B(n4209), .Z(n4335) );
  AND U4569 ( .A(y[230]), .B(x[77]), .Z(n4212) );
  NAND U4570 ( .A(y[241]), .B(x[66]), .Z(n4211) );
  XNOR U4571 ( .A(n4212), .B(n4211), .Z(n4303) );
  XOR U4572 ( .A(n4290), .B(n4289), .Z(n4291) );
  XNOR U4573 ( .A(n4292), .B(n4291), .Z(n4355) );
  XOR U4574 ( .A(n4354), .B(n4355), .Z(n4357) );
  XOR U4575 ( .A(n4356), .B(n4357), .Z(n4286) );
  NAND U4576 ( .A(x[74]), .B(y[241]), .Z(n5392) );
  NANDN U4577 ( .A(n5392), .B(n4213), .Z(n4217) );
  NANDN U4578 ( .A(n4215), .B(n4214), .Z(n4216) );
  AND U4579 ( .A(n4217), .B(n4216), .Z(n4347) );
  NANDN U4580 ( .A(n4219), .B(n4218), .Z(n4223) );
  NANDN U4581 ( .A(n4221), .B(n4220), .Z(n4222) );
  AND U4582 ( .A(n4223), .B(n4222), .Z(n4345) );
  AND U4583 ( .A(y[234]), .B(x[73]), .Z(n4225) );
  NAND U4584 ( .A(y[227]), .B(x[80]), .Z(n4224) );
  XNOR U4585 ( .A(n4225), .B(n4224), .Z(n4298) );
  NAND U4586 ( .A(x[79]), .B(y[228]), .Z(n4299) );
  XNOR U4587 ( .A(n4298), .B(n4299), .Z(n4344) );
  XNOR U4588 ( .A(n4345), .B(n4344), .Z(n4346) );
  XOR U4589 ( .A(n4347), .B(n4346), .Z(n4360) );
  AND U4590 ( .A(x[77]), .B(y[239]), .Z(n5587) );
  NANDN U4591 ( .A(n4226), .B(n5587), .Z(n4230) );
  NANDN U4592 ( .A(n4228), .B(n4227), .Z(n4229) );
  AND U4593 ( .A(n4230), .B(n4229), .Z(n4353) );
  AND U4594 ( .A(y[233]), .B(x[74]), .Z(n4232) );
  NAND U4595 ( .A(y[226]), .B(x[81]), .Z(n4231) );
  XNOR U4596 ( .A(n4232), .B(n4231), .Z(n4340) );
  NAND U4597 ( .A(x[82]), .B(y[225]), .Z(n4317) );
  XOR U4598 ( .A(o[51]), .B(n4317), .Z(n4341) );
  XNOR U4599 ( .A(n4340), .B(n4341), .Z(n4351) );
  AND U4600 ( .A(y[240]), .B(x[67]), .Z(n4234) );
  NAND U4601 ( .A(y[232]), .B(x[75]), .Z(n4233) );
  XNOR U4602 ( .A(n4234), .B(n4233), .Z(n4311) );
  XOR U4603 ( .A(n4351), .B(n4350), .Z(n4352) );
  XOR U4604 ( .A(n4353), .B(n4352), .Z(n4358) );
  NAND U4605 ( .A(n4596), .B(n4235), .Z(n4239) );
  NANDN U4606 ( .A(n4237), .B(n4236), .Z(n4238) );
  AND U4607 ( .A(n4239), .B(n4238), .Z(n4296) );
  AND U4608 ( .A(x[64]), .B(y[243]), .Z(n4322) );
  NAND U4609 ( .A(x[83]), .B(y[224]), .Z(n4323) );
  XNOR U4610 ( .A(n4322), .B(n4323), .Z(n4325) );
  ANDN U4611 ( .B(o[50]), .A(n4240), .Z(n4324) );
  XOR U4612 ( .A(n4325), .B(n4324), .Z(n4294) );
  AND U4613 ( .A(x[68]), .B(y[239]), .Z(n4454) );
  NAND U4614 ( .A(y[238]), .B(x[69]), .Z(n4241) );
  XOR U4615 ( .A(n4242), .B(n4241), .Z(n4319) );
  XNOR U4616 ( .A(n4454), .B(n4319), .Z(n4293) );
  XOR U4617 ( .A(n4294), .B(n4293), .Z(n4295) );
  XOR U4618 ( .A(n4296), .B(n4295), .Z(n4359) );
  XOR U4619 ( .A(n4358), .B(n4359), .Z(n4361) );
  XOR U4620 ( .A(n4360), .B(n4361), .Z(n4364) );
  XNOR U4621 ( .A(n4362), .B(n4363), .Z(n4365) );
  XNOR U4622 ( .A(n4364), .B(n4365), .Z(n4285) );
  XNOR U4623 ( .A(n4286), .B(n4285), .Z(n4288) );
  XOR U4624 ( .A(n4287), .B(n4288), .Z(n4375) );
  NAND U4625 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U4626 ( .A(n4254), .B(n4253), .Z(n4255) );
  AND U4627 ( .A(n4256), .B(n4255), .Z(n4372) );
  NAND U4628 ( .A(n4258), .B(n4257), .Z(n4262) );
  NAND U4629 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U4630 ( .A(n4262), .B(n4261), .Z(n4368) );
  NAND U4631 ( .A(n4264), .B(n4263), .Z(n4268) );
  NANDN U4632 ( .A(n4266), .B(n4265), .Z(n4267) );
  NAND U4633 ( .A(n4268), .B(n4267), .Z(n4367) );
  NAND U4634 ( .A(n4270), .B(n4269), .Z(n4274) );
  NAND U4635 ( .A(n4272), .B(n4271), .Z(n4273) );
  NAND U4636 ( .A(n4274), .B(n4273), .Z(n4366) );
  XNOR U4637 ( .A(n4367), .B(n4366), .Z(n4369) );
  XOR U4638 ( .A(n4368), .B(n4369), .Z(n4373) );
  XNOR U4639 ( .A(n4372), .B(n4373), .Z(n4374) );
  XNOR U4640 ( .A(n4375), .B(n4374), .Z(n4378) );
  XOR U4641 ( .A(n4379), .B(n4378), .Z(n4380) );
  XOR U4642 ( .A(n4381), .B(n4380), .Z(n4386) );
  NANDN U4643 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U4644 ( .A(n4281), .B(n4280), .Z(n4282) );
  NAND U4645 ( .A(n4283), .B(n4282), .Z(n4384) );
  XNOR U4646 ( .A(n4385), .B(n4384), .Z(n4284) );
  XNOR U4647 ( .A(n4386), .B(n4284), .Z(N116) );
  XNOR U4648 ( .A(n4389), .B(n4388), .Z(n4391) );
  AND U4649 ( .A(x[80]), .B(y[234]), .Z(n5214) );
  NAND U4650 ( .A(n5214), .B(n4297), .Z(n4301) );
  NANDN U4651 ( .A(n4299), .B(n4298), .Z(n4300) );
  AND U4652 ( .A(n4301), .B(n4300), .Z(n4429) );
  AND U4653 ( .A(x[77]), .B(y[241]), .Z(n5820) );
  NAND U4654 ( .A(n5820), .B(n4302), .Z(n4306) );
  NANDN U4655 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4656 ( .A(n4306), .B(n4305), .Z(n4474) );
  NAND U4657 ( .A(y[228]), .B(x[80]), .Z(n4307) );
  XNOR U4658 ( .A(n4308), .B(n4307), .Z(n4435) );
  NAND U4659 ( .A(x[66]), .B(y[242]), .Z(n4436) );
  XNOR U4660 ( .A(n4435), .B(n4436), .Z(n4472) );
  NAND U4661 ( .A(y[229]), .B(x[79]), .Z(n4309) );
  XNOR U4662 ( .A(n4310), .B(n4309), .Z(n4405) );
  NAND U4663 ( .A(x[78]), .B(y[230]), .Z(n4406) );
  XNOR U4664 ( .A(n4405), .B(n4406), .Z(n4471) );
  XOR U4665 ( .A(n4472), .B(n4471), .Z(n4473) );
  XNOR U4666 ( .A(n4474), .B(n4473), .Z(n4428) );
  XNOR U4667 ( .A(n4429), .B(n4428), .Z(n4431) );
  NAND U4668 ( .A(x[75]), .B(y[240]), .Z(n5394) );
  NANDN U4669 ( .A(n5394), .B(n4575), .Z(n4314) );
  NANDN U4670 ( .A(n4312), .B(n4311), .Z(n4313) );
  AND U4671 ( .A(n4314), .B(n4313), .Z(n4480) );
  AND U4672 ( .A(y[233]), .B(x[75]), .Z(n4316) );
  NAND U4673 ( .A(y[243]), .B(x[65]), .Z(n4315) );
  XNOR U4674 ( .A(n4316), .B(n4315), .Z(n4401) );
  NAND U4675 ( .A(x[83]), .B(y[225]), .Z(n4409) );
  XNOR U4676 ( .A(o[52]), .B(n4409), .Z(n4400) );
  XOR U4677 ( .A(n4401), .B(n4400), .Z(n4478) );
  AND U4678 ( .A(x[64]), .B(y[244]), .Z(n4459) );
  NAND U4679 ( .A(x[84]), .B(y[224]), .Z(n4460) );
  XNOR U4680 ( .A(n4459), .B(n4460), .Z(n4462) );
  ANDN U4681 ( .B(o[51]), .A(n4317), .Z(n4461) );
  XOR U4682 ( .A(n4462), .B(n4461), .Z(n4477) );
  XOR U4683 ( .A(n4478), .B(n4477), .Z(n4479) );
  XNOR U4684 ( .A(n4480), .B(n4479), .Z(n4430) );
  XOR U4685 ( .A(n4431), .B(n4430), .Z(n4390) );
  XOR U4686 ( .A(n4391), .B(n4390), .Z(n4486) );
  AND U4687 ( .A(x[70]), .B(y[238]), .Z(n4411) );
  AND U4688 ( .A(x[69]), .B(y[237]), .Z(n4318) );
  NAND U4689 ( .A(n4411), .B(n4318), .Z(n4321) );
  NANDN U4690 ( .A(n4319), .B(n4454), .Z(n4320) );
  AND U4691 ( .A(n4321), .B(n4320), .Z(n4419) );
  NANDN U4692 ( .A(n4323), .B(n4322), .Z(n4327) );
  NAND U4693 ( .A(n4325), .B(n4324), .Z(n4326) );
  AND U4694 ( .A(n4327), .B(n4326), .Z(n4417) );
  AND U4695 ( .A(y[226]), .B(x[82]), .Z(n4329) );
  NAND U4696 ( .A(y[232]), .B(x[76]), .Z(n4328) );
  XNOR U4697 ( .A(n4329), .B(n4328), .Z(n4395) );
  NAND U4698 ( .A(x[81]), .B(y[227]), .Z(n4396) );
  XNOR U4699 ( .A(n4395), .B(n4396), .Z(n4416) );
  XNOR U4700 ( .A(n4417), .B(n4416), .Z(n4418) );
  XOR U4701 ( .A(n4419), .B(n4418), .Z(n4423) );
  AND U4702 ( .A(y[231]), .B(x[77]), .Z(n4331) );
  NAND U4703 ( .A(y[241]), .B(x[67]), .Z(n4330) );
  XNOR U4704 ( .A(n4331), .B(n4330), .Z(n4441) );
  XOR U4705 ( .A(n4441), .B(n4440), .Z(n4413) );
  AND U4706 ( .A(y[239]), .B(x[69]), .Z(n4333) );
  NAND U4707 ( .A(y[240]), .B(x[68]), .Z(n4332) );
  XNOR U4708 ( .A(n4333), .B(n4332), .Z(n4456) );
  AND U4709 ( .A(x[71]), .B(y[237]), .Z(n4455) );
  XNOR U4710 ( .A(n4456), .B(n4455), .Z(n4410) );
  XNOR U4711 ( .A(n4411), .B(n4410), .Z(n4412) );
  XOR U4712 ( .A(n4413), .B(n4412), .Z(n4467) );
  AND U4713 ( .A(x[72]), .B(y[242]), .Z(n5537) );
  AND U4714 ( .A(x[65]), .B(y[235]), .Z(n4334) );
  NAND U4715 ( .A(n5537), .B(n4334), .Z(n4338) );
  NANDN U4716 ( .A(n4336), .B(n4335), .Z(n4337) );
  AND U4717 ( .A(n4338), .B(n4337), .Z(n4466) );
  AND U4718 ( .A(x[81]), .B(y[233]), .Z(n5220) );
  NAND U4719 ( .A(n5220), .B(n4339), .Z(n4343) );
  NANDN U4720 ( .A(n4341), .B(n4340), .Z(n4342) );
  NAND U4721 ( .A(n4343), .B(n4342), .Z(n4465) );
  XNOR U4722 ( .A(n4466), .B(n4465), .Z(n4468) );
  XNOR U4723 ( .A(n4467), .B(n4468), .Z(n4422) );
  XOR U4724 ( .A(n4423), .B(n4422), .Z(n4424) );
  NANDN U4725 ( .A(n4345), .B(n4344), .Z(n4349) );
  NANDN U4726 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U4727 ( .A(n4349), .B(n4348), .Z(n4425) );
  XNOR U4728 ( .A(n4424), .B(n4425), .Z(n4483) );
  XNOR U4729 ( .A(n4483), .B(n4484), .Z(n4485) );
  XNOR U4730 ( .A(n4486), .B(n4485), .Z(n4490) );
  XOR U4731 ( .A(n4493), .B(n4494), .Z(n4495) );
  XOR U4732 ( .A(n4496), .B(n4495), .Z(n4489) );
  XOR U4733 ( .A(n4490), .B(n4489), .Z(n4492) );
  XOR U4734 ( .A(n4491), .B(n4492), .Z(n4502) );
  NAND U4735 ( .A(n4367), .B(n4366), .Z(n4371) );
  NANDN U4736 ( .A(n4369), .B(n4368), .Z(n4370) );
  AND U4737 ( .A(n4371), .B(n4370), .Z(n4500) );
  NANDN U4738 ( .A(n4373), .B(n4372), .Z(n4377) );
  NANDN U4739 ( .A(n4375), .B(n4374), .Z(n4376) );
  AND U4740 ( .A(n4377), .B(n4376), .Z(n4499) );
  XOR U4741 ( .A(n4500), .B(n4499), .Z(n4501) );
  XOR U4742 ( .A(n4502), .B(n4501), .Z(n4507) );
  NAND U4743 ( .A(n4379), .B(n4378), .Z(n4383) );
  NANDN U4744 ( .A(n4381), .B(n4380), .Z(n4382) );
  NAND U4745 ( .A(n4383), .B(n4382), .Z(n4505) );
  XOR U4746 ( .A(n4505), .B(n4506), .Z(n4387) );
  XNOR U4747 ( .A(n4507), .B(n4387), .Z(N117) );
  NANDN U4748 ( .A(n4389), .B(n4388), .Z(n4393) );
  NAND U4749 ( .A(n4391), .B(n4390), .Z(n4392) );
  AND U4750 ( .A(n4393), .B(n4392), .Z(n4527) );
  AND U4751 ( .A(x[82]), .B(y[232]), .Z(n5222) );
  NAND U4752 ( .A(n5222), .B(n4394), .Z(n4398) );
  NANDN U4753 ( .A(n4396), .B(n4395), .Z(n4397) );
  AND U4754 ( .A(n4398), .B(n4397), .Z(n4604) );
  AND U4755 ( .A(x[75]), .B(y[243]), .Z(n6018) );
  AND U4756 ( .A(x[65]), .B(y[233]), .Z(n4399) );
  NAND U4757 ( .A(n6018), .B(n4399), .Z(n4403) );
  NAND U4758 ( .A(n4401), .B(n4400), .Z(n4402) );
  NAND U4759 ( .A(n4403), .B(n4402), .Z(n4603) );
  XNOR U4760 ( .A(n4604), .B(n4603), .Z(n4606) );
  AND U4761 ( .A(x[79]), .B(y[235]), .Z(n5209) );
  NAND U4762 ( .A(n5209), .B(n4404), .Z(n4408) );
  NANDN U4763 ( .A(n4406), .B(n4405), .Z(n4407) );
  AND U4764 ( .A(n4408), .B(n4407), .Z(n4562) );
  AND U4765 ( .A(x[64]), .B(y[245]), .Z(n4581) );
  NAND U4766 ( .A(x[85]), .B(y[224]), .Z(n4582) );
  XNOR U4767 ( .A(n4581), .B(n4582), .Z(n4584) );
  ANDN U4768 ( .B(o[52]), .A(n4409), .Z(n4583) );
  XOR U4769 ( .A(n4584), .B(n4583), .Z(n4560) );
  AND U4770 ( .A(x[69]), .B(y[240]), .Z(n4566) );
  AND U4771 ( .A(x[80]), .B(y[229]), .Z(n4565) );
  XOR U4772 ( .A(n4566), .B(n4565), .Z(n4568) );
  NAND U4773 ( .A(x[79]), .B(y[230]), .Z(n4567) );
  XNOR U4774 ( .A(n4568), .B(n4567), .Z(n4559) );
  XOR U4775 ( .A(n4560), .B(n4559), .Z(n4561) );
  XNOR U4776 ( .A(n4562), .B(n4561), .Z(n4605) );
  XOR U4777 ( .A(n4606), .B(n4605), .Z(n4598) );
  NANDN U4778 ( .A(n4411), .B(n4410), .Z(n4415) );
  NANDN U4779 ( .A(n4413), .B(n4412), .Z(n4414) );
  NAND U4780 ( .A(n4415), .B(n4414), .Z(n4597) );
  XNOR U4781 ( .A(n4598), .B(n4597), .Z(n4600) );
  NANDN U4782 ( .A(n4417), .B(n4416), .Z(n4421) );
  NANDN U4783 ( .A(n4419), .B(n4418), .Z(n4420) );
  AND U4784 ( .A(n4421), .B(n4420), .Z(n4599) );
  XOR U4785 ( .A(n4600), .B(n4599), .Z(n4525) );
  NAND U4786 ( .A(n4423), .B(n4422), .Z(n4427) );
  NANDN U4787 ( .A(n4425), .B(n4424), .Z(n4426) );
  AND U4788 ( .A(n4427), .B(n4426), .Z(n4524) );
  XNOR U4789 ( .A(n4525), .B(n4524), .Z(n4526) );
  XOR U4790 ( .A(n4527), .B(n4526), .Z(n4520) );
  NANDN U4791 ( .A(n4429), .B(n4428), .Z(n4433) );
  NAND U4792 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U4793 ( .A(n4433), .B(n4432), .Z(n4624) );
  NAND U4794 ( .A(n5214), .B(n4434), .Z(n4438) );
  NANDN U4795 ( .A(n4436), .B(n4435), .Z(n4437) );
  AND U4796 ( .A(n4438), .B(n4437), .Z(n4531) );
  NAND U4797 ( .A(n5820), .B(n4439), .Z(n4443) );
  NAND U4798 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U4799 ( .A(n4443), .B(n4442), .Z(n4618) );
  AND U4800 ( .A(y[226]), .B(x[83]), .Z(n4445) );
  NAND U4801 ( .A(y[234]), .B(x[75]), .Z(n4444) );
  XNOR U4802 ( .A(n4445), .B(n4444), .Z(n4550) );
  NAND U4803 ( .A(x[84]), .B(y[225]), .Z(n4580) );
  XNOR U4804 ( .A(o[53]), .B(n4580), .Z(n4549) );
  XOR U4805 ( .A(n4550), .B(n4549), .Z(n4616) );
  NAND U4806 ( .A(y[227]), .B(x[82]), .Z(n4446) );
  XNOR U4807 ( .A(n4447), .B(n4446), .Z(n4588) );
  NAND U4808 ( .A(x[65]), .B(y[244]), .Z(n4589) );
  XNOR U4809 ( .A(n4588), .B(n4589), .Z(n4615) );
  XOR U4810 ( .A(n4616), .B(n4615), .Z(n4617) );
  XNOR U4811 ( .A(n4618), .B(n4617), .Z(n4530) );
  XNOR U4812 ( .A(n4531), .B(n4530), .Z(n4533) );
  AND U4813 ( .A(x[71]), .B(y[238]), .Z(n4850) );
  AND U4814 ( .A(y[239]), .B(x[70]), .Z(n4449) );
  NAND U4815 ( .A(y[231]), .B(x[78]), .Z(n4448) );
  XNOR U4816 ( .A(n4449), .B(n4448), .Z(n4592) );
  XOR U4817 ( .A(n4850), .B(n4592), .Z(n4539) );
  AND U4818 ( .A(x[73]), .B(y[236]), .Z(n4537) );
  NAND U4819 ( .A(x[72]), .B(y[237]), .Z(n4536) );
  XNOR U4820 ( .A(n4537), .B(n4536), .Z(n4538) );
  XOR U4821 ( .A(n4539), .B(n4538), .Z(n4555) );
  AND U4822 ( .A(y[233]), .B(x[76]), .Z(n4451) );
  NAND U4823 ( .A(y[228]), .B(x[81]), .Z(n4450) );
  XNOR U4824 ( .A(n4451), .B(n4450), .Z(n4542) );
  NAND U4825 ( .A(x[66]), .B(y[243]), .Z(n4543) );
  XNOR U4826 ( .A(n4542), .B(n4543), .Z(n4554) );
  AND U4827 ( .A(y[232]), .B(x[77]), .Z(n4453) );
  NAND U4828 ( .A(y[242]), .B(x[67]), .Z(n4452) );
  XNOR U4829 ( .A(n4453), .B(n4452), .Z(n4576) );
  NAND U4830 ( .A(x[68]), .B(y[241]), .Z(n4577) );
  XNOR U4831 ( .A(n4576), .B(n4577), .Z(n4553) );
  XOR U4832 ( .A(n4554), .B(n4553), .Z(n4556) );
  XOR U4833 ( .A(n4555), .B(n4556), .Z(n4612) );
  NAND U4834 ( .A(n4566), .B(n4454), .Z(n4458) );
  NAND U4835 ( .A(n4456), .B(n4455), .Z(n4457) );
  AND U4836 ( .A(n4458), .B(n4457), .Z(n4610) );
  NANDN U4837 ( .A(n4460), .B(n4459), .Z(n4464) );
  NAND U4838 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U4839 ( .A(n4464), .B(n4463), .Z(n4609) );
  XNOR U4840 ( .A(n4610), .B(n4609), .Z(n4611) );
  XOR U4841 ( .A(n4612), .B(n4611), .Z(n4532) );
  XOR U4842 ( .A(n4533), .B(n4532), .Z(n4622) );
  NANDN U4843 ( .A(n4466), .B(n4465), .Z(n4470) );
  NAND U4844 ( .A(n4468), .B(n4467), .Z(n4469) );
  NAND U4845 ( .A(n4470), .B(n4469), .Z(n4629) );
  NAND U4846 ( .A(n4472), .B(n4471), .Z(n4476) );
  NANDN U4847 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U4848 ( .A(n4476), .B(n4475), .Z(n4628) );
  NAND U4849 ( .A(n4478), .B(n4477), .Z(n4482) );
  NANDN U4850 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U4851 ( .A(n4482), .B(n4481), .Z(n4627) );
  XOR U4852 ( .A(n4628), .B(n4627), .Z(n4630) );
  XOR U4853 ( .A(n4629), .B(n4630), .Z(n4621) );
  XOR U4854 ( .A(n4622), .B(n4621), .Z(n4623) );
  XOR U4855 ( .A(n4624), .B(n4623), .Z(n4519) );
  NANDN U4856 ( .A(n4484), .B(n4483), .Z(n4488) );
  NANDN U4857 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U4858 ( .A(n4488), .B(n4487), .Z(n4518) );
  XOR U4859 ( .A(n4519), .B(n4518), .Z(n4521) );
  XOR U4860 ( .A(n4520), .B(n4521), .Z(n4512) );
  NAND U4861 ( .A(n4494), .B(n4493), .Z(n4498) );
  NAND U4862 ( .A(n4496), .B(n4495), .Z(n4497) );
  AND U4863 ( .A(n4498), .B(n4497), .Z(n4509) );
  XOR U4864 ( .A(n4510), .B(n4509), .Z(n4511) );
  XOR U4865 ( .A(n4512), .B(n4511), .Z(n4517) );
  NAND U4866 ( .A(n4500), .B(n4499), .Z(n4504) );
  NAND U4867 ( .A(n4502), .B(n4501), .Z(n4503) );
  AND U4868 ( .A(n4504), .B(n4503), .Z(n4515) );
  XNOR U4869 ( .A(n4515), .B(n4516), .Z(n4508) );
  XNOR U4870 ( .A(n4517), .B(n4508), .Z(N118) );
  NAND U4871 ( .A(n4510), .B(n4509), .Z(n4514) );
  NANDN U4872 ( .A(n4512), .B(n4511), .Z(n4513) );
  AND U4873 ( .A(n4514), .B(n4513), .Z(n4759) );
  NAND U4874 ( .A(n4519), .B(n4518), .Z(n4523) );
  NAND U4875 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U4876 ( .A(n4523), .B(n4522), .Z(n4755) );
  NANDN U4877 ( .A(n4525), .B(n4524), .Z(n4529) );
  NANDN U4878 ( .A(n4527), .B(n4526), .Z(n4528) );
  AND U4879 ( .A(n4529), .B(n4528), .Z(n4753) );
  NANDN U4880 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U4881 ( .A(n4533), .B(n4532), .Z(n4534) );
  AND U4882 ( .A(n4535), .B(n4534), .Z(n4749) );
  NANDN U4883 ( .A(n4537), .B(n4536), .Z(n4541) );
  NANDN U4884 ( .A(n4539), .B(n4538), .Z(n4540) );
  AND U4885 ( .A(n4541), .B(n4540), .Z(n4743) );
  NAND U4886 ( .A(n5220), .B(n4695), .Z(n4545) );
  NANDN U4887 ( .A(n4543), .B(n4542), .Z(n4544) );
  NAND U4888 ( .A(n4545), .B(n4544), .Z(n4672) );
  AND U4889 ( .A(x[69]), .B(y[241]), .Z(n4716) );
  NAND U4890 ( .A(x[81]), .B(y[229]), .Z(n4717) );
  XNOR U4891 ( .A(n4716), .B(n4717), .Z(n4718) );
  NAND U4892 ( .A(x[80]), .B(y[230]), .Z(n4719) );
  XNOR U4893 ( .A(n4718), .B(n4719), .Z(n4671) );
  AND U4894 ( .A(y[228]), .B(x[82]), .Z(n4547) );
  NAND U4895 ( .A(y[234]), .B(x[76]), .Z(n4546) );
  XNOR U4896 ( .A(n4547), .B(n4546), .Z(n4696) );
  NAND U4897 ( .A(x[68]), .B(y[242]), .Z(n4697) );
  XNOR U4898 ( .A(n4696), .B(n4697), .Z(n4670) );
  XOR U4899 ( .A(n4671), .B(n4670), .Z(n4673) );
  XNOR U4900 ( .A(n4672), .B(n4673), .Z(n4740) );
  AND U4901 ( .A(x[83]), .B(y[234]), .Z(n5717) );
  NAND U4902 ( .A(n5717), .B(n4548), .Z(n4552) );
  NAND U4903 ( .A(n4550), .B(n4549), .Z(n4551) );
  AND U4904 ( .A(n4552), .B(n4551), .Z(n4741) );
  XOR U4905 ( .A(n4740), .B(n4741), .Z(n4742) );
  XOR U4906 ( .A(n4743), .B(n4742), .Z(n4746) );
  NAND U4907 ( .A(n4554), .B(n4553), .Z(n4558) );
  NAND U4908 ( .A(n4556), .B(n4555), .Z(n4557) );
  AND U4909 ( .A(n4558), .B(n4557), .Z(n4729) );
  NAND U4910 ( .A(n4560), .B(n4559), .Z(n4564) );
  NANDN U4911 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U4912 ( .A(n4564), .B(n4563), .Z(n4728) );
  XNOR U4913 ( .A(n4729), .B(n4728), .Z(n4731) );
  NAND U4914 ( .A(n4566), .B(n4565), .Z(n4570) );
  ANDN U4915 ( .B(n4568), .A(n4567), .Z(n4569) );
  ANDN U4916 ( .B(n4570), .A(n4569), .Z(n4692) );
  AND U4917 ( .A(y[226]), .B(x[84]), .Z(n4572) );
  NAND U4918 ( .A(y[233]), .B(x[77]), .Z(n4571) );
  XNOR U4919 ( .A(n4572), .B(n4571), .Z(n4712) );
  NAND U4920 ( .A(x[66]), .B(y[244]), .Z(n4713) );
  XNOR U4921 ( .A(n4712), .B(n4713), .Z(n4690) );
  AND U4922 ( .A(y[231]), .B(x[79]), .Z(n4574) );
  NAND U4923 ( .A(y[240]), .B(x[70]), .Z(n4573) );
  XOR U4924 ( .A(n4574), .B(n4573), .Z(n4725) );
  XNOR U4925 ( .A(n4724), .B(n4725), .Z(n4689) );
  XOR U4926 ( .A(n4690), .B(n4689), .Z(n4691) );
  XNOR U4927 ( .A(n4692), .B(n4691), .Z(n4735) );
  AND U4928 ( .A(x[77]), .B(y[242]), .Z(n6020) );
  NAND U4929 ( .A(n4575), .B(n6020), .Z(n4579) );
  NANDN U4930 ( .A(n4577), .B(n4576), .Z(n4578) );
  AND U4931 ( .A(n4579), .B(n4578), .Z(n4661) );
  AND U4932 ( .A(x[65]), .B(y[245]), .Z(n4684) );
  XOR U4933 ( .A(n4685), .B(n4684), .Z(n4683) );
  ANDN U4934 ( .B(o[53]), .A(n4580), .Z(n4682) );
  XOR U4935 ( .A(n4683), .B(n4682), .Z(n4659) );
  AND U4936 ( .A(x[78]), .B(y[232]), .Z(n4676) );
  NAND U4937 ( .A(x[67]), .B(y[243]), .Z(n4677) );
  XNOR U4938 ( .A(n4676), .B(n4677), .Z(n4678) );
  NAND U4939 ( .A(x[83]), .B(y[227]), .Z(n4679) );
  XNOR U4940 ( .A(n4678), .B(n4679), .Z(n4658) );
  XOR U4941 ( .A(n4659), .B(n4658), .Z(n4660) );
  XNOR U4942 ( .A(n4661), .B(n4660), .Z(n4734) );
  XOR U4943 ( .A(n4735), .B(n4734), .Z(n4737) );
  NANDN U4944 ( .A(n4582), .B(n4581), .Z(n4586) );
  NAND U4945 ( .A(n4584), .B(n4583), .Z(n4585) );
  AND U4946 ( .A(n4586), .B(n4585), .Z(n4653) );
  AND U4947 ( .A(x[82]), .B(y[235]), .Z(n5719) );
  NAND U4948 ( .A(n5719), .B(n4587), .Z(n4591) );
  NANDN U4949 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U4950 ( .A(n4591), .B(n4590), .Z(n4652) );
  XNOR U4951 ( .A(n4653), .B(n4652), .Z(n4655) );
  AND U4952 ( .A(x[78]), .B(y[239]), .Z(n5729) );
  NAND U4953 ( .A(n4723), .B(n5729), .Z(n4594) );
  NAND U4954 ( .A(n4850), .B(n4592), .Z(n4593) );
  AND U4955 ( .A(n4594), .B(n4593), .Z(n4667) );
  AND U4956 ( .A(x[64]), .B(y[246]), .Z(n4700) );
  NAND U4957 ( .A(x[86]), .B(y[224]), .Z(n4701) );
  XNOR U4958 ( .A(n4700), .B(n4701), .Z(n4703) );
  NAND U4959 ( .A(x[85]), .B(y[225]), .Z(n4722) );
  XNOR U4960 ( .A(o[54]), .B(n4722), .Z(n4702) );
  XOR U4961 ( .A(n4703), .B(n4702), .Z(n4665) );
  NAND U4962 ( .A(y[239]), .B(x[71]), .Z(n4595) );
  XOR U4963 ( .A(n4596), .B(n4595), .Z(n4707) );
  XNOR U4964 ( .A(n4706), .B(n4707), .Z(n4664) );
  XOR U4965 ( .A(n4665), .B(n4664), .Z(n4666) );
  XNOR U4966 ( .A(n4667), .B(n4666), .Z(n4654) );
  XOR U4967 ( .A(n4655), .B(n4654), .Z(n4736) );
  XOR U4968 ( .A(n4737), .B(n4736), .Z(n4730) );
  XOR U4969 ( .A(n4731), .B(n4730), .Z(n4747) );
  XOR U4970 ( .A(n4746), .B(n4747), .Z(n4748) );
  XOR U4971 ( .A(n4749), .B(n4748), .Z(n4642) );
  NANDN U4972 ( .A(n4598), .B(n4597), .Z(n4602) );
  NAND U4973 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U4974 ( .A(n4602), .B(n4601), .Z(n4641) );
  NANDN U4975 ( .A(n4604), .B(n4603), .Z(n4608) );
  NAND U4976 ( .A(n4606), .B(n4605), .Z(n4607) );
  AND U4977 ( .A(n4608), .B(n4607), .Z(n4649) );
  NANDN U4978 ( .A(n4610), .B(n4609), .Z(n4614) );
  NAND U4979 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U4980 ( .A(n4614), .B(n4613), .Z(n4647) );
  NAND U4981 ( .A(n4616), .B(n4615), .Z(n4620) );
  NANDN U4982 ( .A(n4618), .B(n4617), .Z(n4619) );
  NAND U4983 ( .A(n4620), .B(n4619), .Z(n4646) );
  XNOR U4984 ( .A(n4647), .B(n4646), .Z(n4648) );
  XOR U4985 ( .A(n4649), .B(n4648), .Z(n4640) );
  XNOR U4986 ( .A(n4641), .B(n4640), .Z(n4643) );
  XNOR U4987 ( .A(n4642), .B(n4643), .Z(n4636) );
  NAND U4988 ( .A(n4622), .B(n4621), .Z(n4626) );
  NANDN U4989 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U4990 ( .A(n4626), .B(n4625), .Z(n4635) );
  NAND U4991 ( .A(n4628), .B(n4627), .Z(n4632) );
  NAND U4992 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U4993 ( .A(n4632), .B(n4631), .Z(n4634) );
  XNOR U4994 ( .A(n4635), .B(n4634), .Z(n4637) );
  XOR U4995 ( .A(n4636), .B(n4637), .Z(n4752) );
  XNOR U4996 ( .A(n4753), .B(n4752), .Z(n4754) );
  XOR U4997 ( .A(n4755), .B(n4754), .Z(n4760) );
  XOR U4998 ( .A(n4758), .B(n4760), .Z(n4633) );
  XOR U4999 ( .A(n4759), .B(n4633), .Z(N119) );
  NANDN U5000 ( .A(n4635), .B(n4634), .Z(n4639) );
  NAND U5001 ( .A(n4637), .B(n4636), .Z(n4638) );
  AND U5002 ( .A(n4639), .B(n4638), .Z(n4765) );
  NANDN U5003 ( .A(n4641), .B(n4640), .Z(n4645) );
  NAND U5004 ( .A(n4643), .B(n4642), .Z(n4644) );
  AND U5005 ( .A(n4645), .B(n4644), .Z(n4763) );
  NANDN U5006 ( .A(n4647), .B(n4646), .Z(n4651) );
  NANDN U5007 ( .A(n4649), .B(n4648), .Z(n4650) );
  AND U5008 ( .A(n4651), .B(n4650), .Z(n4886) );
  NANDN U5009 ( .A(n4653), .B(n4652), .Z(n4657) );
  NAND U5010 ( .A(n4655), .B(n4654), .Z(n4656) );
  AND U5011 ( .A(n4657), .B(n4656), .Z(n4834) );
  NAND U5012 ( .A(n4659), .B(n4658), .Z(n4663) );
  NANDN U5013 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U5014 ( .A(n4663), .B(n4662), .Z(n4832) );
  NAND U5015 ( .A(n4665), .B(n4664), .Z(n4669) );
  NANDN U5016 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U5017 ( .A(n4669), .B(n4668), .Z(n4831) );
  XNOR U5018 ( .A(n4832), .B(n4831), .Z(n4833) );
  XNOR U5019 ( .A(n4834), .B(n4833), .Z(n4898) );
  NAND U5020 ( .A(n4671), .B(n4670), .Z(n4675) );
  NAND U5021 ( .A(n4673), .B(n4672), .Z(n4674) );
  AND U5022 ( .A(n4675), .B(n4674), .Z(n4896) );
  NANDN U5023 ( .A(n4677), .B(n4676), .Z(n4681) );
  NANDN U5024 ( .A(n4679), .B(n4678), .Z(n4680) );
  AND U5025 ( .A(n4681), .B(n4680), .Z(n4778) );
  AND U5026 ( .A(n4683), .B(n4682), .Z(n4687) );
  NAND U5027 ( .A(n4685), .B(n4684), .Z(n4686) );
  NANDN U5028 ( .A(n4687), .B(n4686), .Z(n4777) );
  XNOR U5029 ( .A(n4778), .B(n4777), .Z(n4780) );
  NAND U5030 ( .A(y[240]), .B(x[71]), .Z(n4688) );
  XOR U5031 ( .A(n4920), .B(n4688), .Z(n4852) );
  XNOR U5032 ( .A(n4851), .B(n4852), .Z(n4783) );
  NAND U5033 ( .A(x[74]), .B(y[237]), .Z(n4784) );
  XNOR U5034 ( .A(n4783), .B(n4784), .Z(n4786) );
  AND U5035 ( .A(x[70]), .B(y[241]), .Z(n4842) );
  NAND U5036 ( .A(x[79]), .B(y[232]), .Z(n4843) );
  XNOR U5037 ( .A(n4842), .B(n4843), .Z(n4844) );
  NAND U5038 ( .A(x[75]), .B(y[236]), .Z(n4845) );
  XNOR U5039 ( .A(n4844), .B(n4845), .Z(n4785) );
  XOR U5040 ( .A(n4786), .B(n4785), .Z(n4779) );
  XOR U5041 ( .A(n4780), .B(n4779), .Z(n4895) );
  XNOR U5042 ( .A(n4896), .B(n4895), .Z(n4897) );
  XOR U5043 ( .A(n4898), .B(n4897), .Z(n4884) );
  NAND U5044 ( .A(n4690), .B(n4689), .Z(n4694) );
  NANDN U5045 ( .A(n4692), .B(n4691), .Z(n4693) );
  AND U5046 ( .A(n4694), .B(n4693), .Z(n4878) );
  AND U5047 ( .A(x[82]), .B(y[234]), .Z(n5575) );
  NAND U5048 ( .A(n5575), .B(n4695), .Z(n4699) );
  NANDN U5049 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U5050 ( .A(n4699), .B(n4698), .Z(n4820) );
  NANDN U5051 ( .A(n4701), .B(n4700), .Z(n4705) );
  NAND U5052 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U5053 ( .A(n4705), .B(n4704), .Z(n4819) );
  XOR U5054 ( .A(n4820), .B(n4819), .Z(n4821) );
  NAND U5055 ( .A(n4850), .B(n4851), .Z(n4709) );
  NANDN U5056 ( .A(n4707), .B(n4706), .Z(n4708) );
  NAND U5057 ( .A(n4709), .B(n4708), .Z(n4815) );
  AND U5058 ( .A(x[64]), .B(y[247]), .Z(n4861) );
  NAND U5059 ( .A(x[87]), .B(y[224]), .Z(n4862) );
  XNOR U5060 ( .A(n4861), .B(n4862), .Z(n4864) );
  NAND U5061 ( .A(x[86]), .B(y[225]), .Z(n4841) );
  XNOR U5062 ( .A(o[55]), .B(n4841), .Z(n4863) );
  XOR U5063 ( .A(n4864), .B(n4863), .Z(n4814) );
  AND U5064 ( .A(y[227]), .B(x[84]), .Z(n5433) );
  NAND U5065 ( .A(y[231]), .B(x[80]), .Z(n4710) );
  XNOR U5066 ( .A(n5433), .B(n4710), .Z(n4837) );
  NAND U5067 ( .A(x[83]), .B(y[228]), .Z(n4838) );
  XNOR U5068 ( .A(n4837), .B(n4838), .Z(n4813) );
  XOR U5069 ( .A(n4814), .B(n4813), .Z(n4816) );
  XNOR U5070 ( .A(n4815), .B(n4816), .Z(n4822) );
  XNOR U5071 ( .A(n4821), .B(n4822), .Z(n4877) );
  XNOR U5072 ( .A(n4878), .B(n4877), .Z(n4880) );
  AND U5073 ( .A(x[84]), .B(y[233]), .Z(n5741) );
  NAND U5074 ( .A(n5741), .B(n4711), .Z(n4715) );
  NANDN U5075 ( .A(n4713), .B(n4712), .Z(n4714) );
  AND U5076 ( .A(n4715), .B(n4714), .Z(n4872) );
  NANDN U5077 ( .A(n4717), .B(n4716), .Z(n4721) );
  NANDN U5078 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U5079 ( .A(n4721), .B(n4720), .Z(n4827) );
  AND U5080 ( .A(x[77]), .B(y[234]), .Z(n4801) );
  NAND U5081 ( .A(x[66]), .B(y[245]), .Z(n4802) );
  XNOR U5082 ( .A(n4801), .B(n4802), .Z(n4803) );
  NAND U5083 ( .A(x[85]), .B(y[226]), .Z(n4804) );
  XNOR U5084 ( .A(n4803), .B(n4804), .Z(n4826) );
  AND U5085 ( .A(x[76]), .B(y[235]), .Z(n4855) );
  NAND U5086 ( .A(x[65]), .B(y[246]), .Z(n4856) );
  XNOR U5087 ( .A(n4855), .B(n4856), .Z(n4858) );
  ANDN U5088 ( .B(o[54]), .A(n4722), .Z(n4857) );
  XOR U5089 ( .A(n4858), .B(n4857), .Z(n4825) );
  XOR U5090 ( .A(n4826), .B(n4825), .Z(n4828) );
  XOR U5091 ( .A(n4827), .B(n4828), .Z(n4871) );
  XNOR U5092 ( .A(n4872), .B(n4871), .Z(n4874) );
  AND U5093 ( .A(x[79]), .B(y[240]), .Z(n5953) );
  NAND U5094 ( .A(n5953), .B(n4723), .Z(n4727) );
  NANDN U5095 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U5096 ( .A(n4727), .B(n4726), .Z(n4809) );
  AND U5097 ( .A(x[78]), .B(y[233]), .Z(n4795) );
  NAND U5098 ( .A(x[67]), .B(y[244]), .Z(n4796) );
  XNOR U5099 ( .A(n4795), .B(n4796), .Z(n4797) );
  NAND U5100 ( .A(x[68]), .B(y[243]), .Z(n4798) );
  XNOR U5101 ( .A(n4797), .B(n4798), .Z(n4808) );
  AND U5102 ( .A(x[69]), .B(y[242]), .Z(n4789) );
  NAND U5103 ( .A(x[82]), .B(y[229]), .Z(n4790) );
  XNOR U5104 ( .A(n4789), .B(n4790), .Z(n4792) );
  AND U5105 ( .A(x[81]), .B(y[230]), .Z(n4791) );
  XOR U5106 ( .A(n4792), .B(n4791), .Z(n4807) );
  XOR U5107 ( .A(n4808), .B(n4807), .Z(n4810) );
  XOR U5108 ( .A(n4809), .B(n4810), .Z(n4873) );
  XOR U5109 ( .A(n4874), .B(n4873), .Z(n4879) );
  XOR U5110 ( .A(n4880), .B(n4879), .Z(n4883) );
  XOR U5111 ( .A(n4884), .B(n4883), .Z(n4885) );
  XOR U5112 ( .A(n4886), .B(n4885), .Z(n4773) );
  NANDN U5113 ( .A(n4729), .B(n4728), .Z(n4733) );
  NAND U5114 ( .A(n4731), .B(n4730), .Z(n4732) );
  AND U5115 ( .A(n4733), .B(n4732), .Z(n4892) );
  NAND U5116 ( .A(n4735), .B(n4734), .Z(n4739) );
  NAND U5117 ( .A(n4737), .B(n4736), .Z(n4738) );
  AND U5118 ( .A(n4739), .B(n4738), .Z(n4890) );
  NAND U5119 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U5120 ( .A(n4743), .B(n4742), .Z(n4744) );
  AND U5121 ( .A(n4745), .B(n4744), .Z(n4889) );
  XNOR U5122 ( .A(n4890), .B(n4889), .Z(n4891) );
  XOR U5123 ( .A(n4892), .B(n4891), .Z(n4771) );
  NAND U5124 ( .A(n4747), .B(n4746), .Z(n4751) );
  NANDN U5125 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U5126 ( .A(n4751), .B(n4750), .Z(n4772) );
  XOR U5127 ( .A(n4771), .B(n4772), .Z(n4774) );
  XOR U5128 ( .A(n4773), .B(n4774), .Z(n4762) );
  XNOR U5129 ( .A(n4763), .B(n4762), .Z(n4764) );
  XOR U5130 ( .A(n4765), .B(n4764), .Z(n4770) );
  NANDN U5131 ( .A(n4753), .B(n4752), .Z(n4757) );
  NAND U5132 ( .A(n4755), .B(n4754), .Z(n4756) );
  NAND U5133 ( .A(n4757), .B(n4756), .Z(n4769) );
  XOR U5134 ( .A(n4769), .B(n4768), .Z(n4761) );
  XNOR U5135 ( .A(n4770), .B(n4761), .Z(N120) );
  NANDN U5136 ( .A(n4763), .B(n4762), .Z(n4767) );
  NAND U5137 ( .A(n4765), .B(n4764), .Z(n4766) );
  NAND U5138 ( .A(n4767), .B(n4766), .Z(n5041) );
  IV U5139 ( .A(n5041), .Z(n5039) );
  NAND U5140 ( .A(n4772), .B(n4771), .Z(n4776) );
  NAND U5141 ( .A(n4774), .B(n4773), .Z(n4775) );
  AND U5142 ( .A(n4776), .B(n4775), .Z(n5036) );
  NANDN U5143 ( .A(n4778), .B(n4777), .Z(n4782) );
  NAND U5144 ( .A(n4780), .B(n4779), .Z(n4781) );
  AND U5145 ( .A(n4782), .B(n4781), .Z(n4977) );
  NANDN U5146 ( .A(n4784), .B(n4783), .Z(n4788) );
  NAND U5147 ( .A(n4786), .B(n4785), .Z(n4787) );
  AND U5148 ( .A(n4788), .B(n4787), .Z(n4975) );
  NANDN U5149 ( .A(n4790), .B(n4789), .Z(n4794) );
  NAND U5150 ( .A(n4792), .B(n4791), .Z(n4793) );
  AND U5151 ( .A(n4794), .B(n4793), .Z(n5001) );
  AND U5152 ( .A(x[64]), .B(y[248]), .Z(n4957) );
  AND U5153 ( .A(x[88]), .B(y[224]), .Z(n4956) );
  XOR U5154 ( .A(n4957), .B(n4956), .Z(n4959) );
  AND U5155 ( .A(x[87]), .B(y[225]), .Z(n4949) );
  XOR U5156 ( .A(n4949), .B(o[56]), .Z(n4958) );
  XOR U5157 ( .A(n4959), .B(n4958), .Z(n4999) );
  AND U5158 ( .A(x[71]), .B(y[241]), .Z(n4943) );
  AND U5159 ( .A(x[82]), .B(y[230]), .Z(n4942) );
  XOR U5160 ( .A(n4943), .B(n4942), .Z(n4945) );
  AND U5161 ( .A(x[81]), .B(y[231]), .Z(n4944) );
  XOR U5162 ( .A(n4945), .B(n4944), .Z(n4998) );
  XOR U5163 ( .A(n4999), .B(n4998), .Z(n5000) );
  XNOR U5164 ( .A(n5001), .B(n5000), .Z(n4989) );
  NANDN U5165 ( .A(n4796), .B(n4795), .Z(n4800) );
  NANDN U5166 ( .A(n4798), .B(n4797), .Z(n4799) );
  AND U5167 ( .A(n4800), .B(n4799), .Z(n4987) );
  NANDN U5168 ( .A(n4802), .B(n4801), .Z(n4806) );
  NANDN U5169 ( .A(n4804), .B(n4803), .Z(n4805) );
  NAND U5170 ( .A(n4806), .B(n4805), .Z(n4986) );
  XNOR U5171 ( .A(n4987), .B(n4986), .Z(n4988) );
  XOR U5172 ( .A(n4989), .B(n4988), .Z(n4974) );
  XNOR U5173 ( .A(n4975), .B(n4974), .Z(n4976) );
  XOR U5174 ( .A(n4977), .B(n4976), .Z(n4982) );
  NAND U5175 ( .A(n4808), .B(n4807), .Z(n4812) );
  NAND U5176 ( .A(n4810), .B(n4809), .Z(n4811) );
  AND U5177 ( .A(n4812), .B(n4811), .Z(n5028) );
  NAND U5178 ( .A(n4814), .B(n4813), .Z(n4818) );
  NAND U5179 ( .A(n4816), .B(n4815), .Z(n4817) );
  AND U5180 ( .A(n4818), .B(n4817), .Z(n5027) );
  XOR U5181 ( .A(n5028), .B(n5027), .Z(n5030) );
  NAND U5182 ( .A(n4820), .B(n4819), .Z(n4824) );
  NANDN U5183 ( .A(n4822), .B(n4821), .Z(n4823) );
  AND U5184 ( .A(n4824), .B(n4823), .Z(n5029) );
  XOR U5185 ( .A(n5030), .B(n5029), .Z(n4980) );
  NAND U5186 ( .A(n4826), .B(n4825), .Z(n4830) );
  NAND U5187 ( .A(n4828), .B(n4827), .Z(n4829) );
  NAND U5188 ( .A(n4830), .B(n4829), .Z(n4981) );
  XNOR U5189 ( .A(n4980), .B(n4981), .Z(n4983) );
  XOR U5190 ( .A(n4982), .B(n4983), .Z(n4908) );
  NANDN U5191 ( .A(n4832), .B(n4831), .Z(n4836) );
  NANDN U5192 ( .A(n4834), .B(n4833), .Z(n4835) );
  NAND U5193 ( .A(n4836), .B(n4835), .Z(n4909) );
  XNOR U5194 ( .A(n4908), .B(n4909), .Z(n4911) );
  AND U5195 ( .A(x[80]), .B(y[227]), .Z(n5004) );
  AND U5196 ( .A(x[84]), .B(y[231]), .Z(n5320) );
  NAND U5197 ( .A(n5004), .B(n5320), .Z(n4840) );
  NANDN U5198 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U5199 ( .A(n4840), .B(n4839), .Z(n5024) );
  AND U5200 ( .A(x[86]), .B(y[226]), .Z(n4930) );
  XOR U5201 ( .A(n4931), .B(n4930), .Z(n4933) );
  AND U5202 ( .A(x[66]), .B(y[246]), .Z(n4932) );
  XOR U5203 ( .A(n4933), .B(n4932), .Z(n5022) );
  AND U5204 ( .A(x[65]), .B(y[247]), .Z(n4938) );
  XOR U5205 ( .A(n4939), .B(n4938), .Z(n4937) );
  ANDN U5206 ( .B(o[55]), .A(n4841), .Z(n4936) );
  XOR U5207 ( .A(n4937), .B(n4936), .Z(n5021) );
  XOR U5208 ( .A(n5022), .B(n5021), .Z(n5023) );
  XNOR U5209 ( .A(n5024), .B(n5023), .Z(n4969) );
  NANDN U5210 ( .A(n4843), .B(n4842), .Z(n4847) );
  NANDN U5211 ( .A(n4845), .B(n4844), .Z(n4846) );
  AND U5212 ( .A(n4847), .B(n4846), .Z(n5018) );
  AND U5213 ( .A(y[227]), .B(x[85]), .Z(n4849) );
  NAND U5214 ( .A(y[232]), .B(x[80]), .Z(n4848) );
  XNOR U5215 ( .A(n4849), .B(n4848), .Z(n5006) );
  AND U5216 ( .A(x[69]), .B(y[243]), .Z(n5005) );
  XOR U5217 ( .A(n5006), .B(n5005), .Z(n5016) );
  AND U5218 ( .A(x[84]), .B(y[228]), .Z(n5160) );
  NAND U5219 ( .A(x[70]), .B(y[242]), .Z(n5307) );
  XNOR U5220 ( .A(n5160), .B(n5307), .Z(n5012) );
  AND U5221 ( .A(x[83]), .B(y[229]), .Z(n5011) );
  XOR U5222 ( .A(n5012), .B(n5011), .Z(n5015) );
  XOR U5223 ( .A(n5016), .B(n5015), .Z(n5017) );
  XNOR U5224 ( .A(n5018), .B(n5017), .Z(n4995) );
  NAND U5225 ( .A(n5093), .B(n4850), .Z(n4854) );
  NANDN U5226 ( .A(n4852), .B(n4851), .Z(n4853) );
  AND U5227 ( .A(n4854), .B(n4853), .Z(n4993) );
  NANDN U5228 ( .A(n4856), .B(n4855), .Z(n4860) );
  NAND U5229 ( .A(n4858), .B(n4857), .Z(n4859) );
  NAND U5230 ( .A(n4860), .B(n4859), .Z(n4992) );
  XNOR U5231 ( .A(n4993), .B(n4992), .Z(n4994) );
  XOR U5232 ( .A(n4995), .B(n4994), .Z(n4968) );
  XOR U5233 ( .A(n4969), .B(n4968), .Z(n4971) );
  NANDN U5234 ( .A(n4862), .B(n4861), .Z(n4866) );
  NAND U5235 ( .A(n4864), .B(n4863), .Z(n4865) );
  AND U5236 ( .A(n4866), .B(n4865), .Z(n4963) );
  AND U5237 ( .A(x[67]), .B(y[245]), .Z(n4950) );
  XOR U5238 ( .A(n4951), .B(n4950), .Z(n4953) );
  NAND U5239 ( .A(x[68]), .B(y[244]), .Z(n4952) );
  XNOR U5240 ( .A(n4953), .B(n4952), .Z(n4962) );
  AND U5241 ( .A(y[238]), .B(x[74]), .Z(n4868) );
  NAND U5242 ( .A(y[239]), .B(x[73]), .Z(n4867) );
  XNOR U5243 ( .A(n4868), .B(n4867), .Z(n4922) );
  AND U5244 ( .A(y[240]), .B(x[72]), .Z(n4870) );
  NAND U5245 ( .A(y[234]), .B(x[78]), .Z(n4869) );
  XNOR U5246 ( .A(n4870), .B(n4869), .Z(n4926) );
  NAND U5247 ( .A(x[75]), .B(y[237]), .Z(n4927) );
  XOR U5248 ( .A(n4922), .B(n4921), .Z(n4964) );
  XOR U5249 ( .A(n4965), .B(n4964), .Z(n4970) );
  XOR U5250 ( .A(n4971), .B(n4970), .Z(n4915) );
  NANDN U5251 ( .A(n4872), .B(n4871), .Z(n4876) );
  NAND U5252 ( .A(n4874), .B(n4873), .Z(n4875) );
  AND U5253 ( .A(n4876), .B(n4875), .Z(n4914) );
  XNOR U5254 ( .A(n4915), .B(n4914), .Z(n4916) );
  NANDN U5255 ( .A(n4878), .B(n4877), .Z(n4882) );
  NAND U5256 ( .A(n4880), .B(n4879), .Z(n4881) );
  NAND U5257 ( .A(n4882), .B(n4881), .Z(n4917) );
  XNOR U5258 ( .A(n4916), .B(n4917), .Z(n4910) );
  XOR U5259 ( .A(n4911), .B(n4910), .Z(n5034) );
  NAND U5260 ( .A(n4884), .B(n4883), .Z(n4888) );
  NANDN U5261 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5262 ( .A(n4888), .B(n4887), .Z(n4905) );
  NANDN U5263 ( .A(n4890), .B(n4889), .Z(n4894) );
  NANDN U5264 ( .A(n4892), .B(n4891), .Z(n4893) );
  AND U5265 ( .A(n4894), .B(n4893), .Z(n4903) );
  NANDN U5266 ( .A(n4896), .B(n4895), .Z(n4900) );
  NAND U5267 ( .A(n4898), .B(n4897), .Z(n4899) );
  NAND U5268 ( .A(n4900), .B(n4899), .Z(n4902) );
  XNOR U5269 ( .A(n4903), .B(n4902), .Z(n4904) );
  XNOR U5270 ( .A(n4905), .B(n4904), .Z(n5033) );
  XNOR U5271 ( .A(n5034), .B(n5033), .Z(n5035) );
  XOR U5272 ( .A(n5036), .B(n5035), .Z(n5042) );
  XNOR U5273 ( .A(n5040), .B(n5042), .Z(n4901) );
  XOR U5274 ( .A(n5039), .B(n4901), .Z(N121) );
  NANDN U5275 ( .A(n4903), .B(n4902), .Z(n4907) );
  NANDN U5276 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U5277 ( .A(n4907), .B(n4906), .Z(n5050) );
  NANDN U5278 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U5279 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U5280 ( .A(n4913), .B(n4912), .Z(n5048) );
  NANDN U5281 ( .A(n4915), .B(n4914), .Z(n4919) );
  NANDN U5282 ( .A(n4917), .B(n4916), .Z(n4918) );
  AND U5283 ( .A(n4919), .B(n4918), .Z(n5057) );
  NANDN U5284 ( .A(n5092), .B(n4920), .Z(n4924) );
  NAND U5285 ( .A(n4922), .B(n4921), .Z(n4923) );
  AND U5286 ( .A(n4924), .B(n4923), .Z(n5117) );
  AND U5287 ( .A(x[78]), .B(y[240]), .Z(n6000) );
  NAND U5288 ( .A(n6000), .B(n4925), .Z(n4929) );
  NANDN U5289 ( .A(n4927), .B(n4926), .Z(n4928) );
  AND U5290 ( .A(n4929), .B(n4928), .Z(n5144) );
  NAND U5291 ( .A(x[75]), .B(y[238]), .Z(n5158) );
  NAND U5292 ( .A(x[76]), .B(y[237]), .Z(n5156) );
  NAND U5293 ( .A(x[71]), .B(y[242]), .Z(n5157) );
  XNOR U5294 ( .A(n5156), .B(n5157), .Z(n5159) );
  XOR U5295 ( .A(n5158), .B(n5159), .Z(n5141) );
  NAND U5296 ( .A(x[88]), .B(y[225]), .Z(n5155) );
  XNOR U5297 ( .A(o[57]), .B(n5155), .Z(n5129) );
  NAND U5298 ( .A(x[65]), .B(y[248]), .Z(n5130) );
  NAND U5299 ( .A(x[77]), .B(y[236]), .Z(n5132) );
  XOR U5300 ( .A(n5141), .B(n5142), .Z(n5143) );
  XNOR U5301 ( .A(n5117), .B(n5116), .Z(n5119) );
  NAND U5302 ( .A(n4931), .B(n4930), .Z(n4935) );
  AND U5303 ( .A(n4933), .B(n4932), .Z(n4934) );
  ANDN U5304 ( .B(n4935), .A(n4934), .Z(n5105) );
  AND U5305 ( .A(n4937), .B(n4936), .Z(n4941) );
  NAND U5306 ( .A(n4939), .B(n4938), .Z(n4940) );
  NANDN U5307 ( .A(n4941), .B(n4940), .Z(n5104) );
  XNOR U5308 ( .A(n5105), .B(n5104), .Z(n5107) );
  NAND U5309 ( .A(n4943), .B(n4942), .Z(n4947) );
  NAND U5310 ( .A(n4945), .B(n4944), .Z(n4946) );
  AND U5311 ( .A(n4947), .B(n4946), .Z(n5101) );
  AND U5312 ( .A(x[72]), .B(y[241]), .Z(n5095) );
  XOR U5313 ( .A(n5093), .B(n4948), .Z(n5094) );
  XOR U5314 ( .A(n5095), .B(n5094), .Z(n5099) );
  AND U5315 ( .A(n4949), .B(o[56]), .Z(n5088) );
  AND U5316 ( .A(x[89]), .B(y[224]), .Z(n5087) );
  NAND U5317 ( .A(x[64]), .B(y[249]), .Z(n5086) );
  XOR U5318 ( .A(n5087), .B(n5086), .Z(n5089) );
  XNOR U5319 ( .A(n5088), .B(n5089), .Z(n5098) );
  XOR U5320 ( .A(n5099), .B(n5098), .Z(n5100) );
  XNOR U5321 ( .A(n5101), .B(n5100), .Z(n5106) );
  XOR U5322 ( .A(n5107), .B(n5106), .Z(n5118) );
  XOR U5323 ( .A(n5119), .B(n5118), .Z(n5071) );
  NAND U5324 ( .A(n4951), .B(n4950), .Z(n4955) );
  ANDN U5325 ( .B(n4953), .A(n4952), .Z(n4954) );
  ANDN U5326 ( .B(n4955), .A(n4954), .Z(n5172) );
  NAND U5327 ( .A(n4957), .B(n4956), .Z(n4961) );
  NAND U5328 ( .A(n4959), .B(n4958), .Z(n4960) );
  AND U5329 ( .A(n4961), .B(n4960), .Z(n5170) );
  AND U5330 ( .A(x[78]), .B(y[235]), .Z(n5135) );
  NAND U5331 ( .A(x[66]), .B(y[247]), .Z(n5136) );
  XNOR U5332 ( .A(n5135), .B(n5136), .Z(n5137) );
  NAND U5333 ( .A(x[67]), .B(y[246]), .Z(n5138) );
  XNOR U5334 ( .A(n5137), .B(n5138), .Z(n5169) );
  XNOR U5335 ( .A(n5170), .B(n5169), .Z(n5171) );
  XOR U5336 ( .A(n5172), .B(n5171), .Z(n5068) );
  NANDN U5337 ( .A(n4963), .B(n4962), .Z(n4967) );
  NAND U5338 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U5339 ( .A(n4967), .B(n4966), .Z(n5069) );
  XOR U5340 ( .A(n5068), .B(n5069), .Z(n5070) );
  NAND U5341 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U5342 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U5343 ( .A(n4973), .B(n4972), .Z(n5075) );
  XNOR U5344 ( .A(n5074), .B(n5075), .Z(n5076) );
  NANDN U5345 ( .A(n4975), .B(n4974), .Z(n4979) );
  NANDN U5346 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5347 ( .A(n4979), .B(n4978), .Z(n5077) );
  XNOR U5348 ( .A(n5076), .B(n5077), .Z(n5056) );
  XNOR U5349 ( .A(n5057), .B(n5056), .Z(n5059) );
  NANDN U5350 ( .A(n4981), .B(n4980), .Z(n4985) );
  NAND U5351 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5352 ( .A(n4985), .B(n4984), .Z(n5064) );
  NANDN U5353 ( .A(n4987), .B(n4986), .Z(n4991) );
  NAND U5354 ( .A(n4989), .B(n4988), .Z(n4990) );
  AND U5355 ( .A(n4991), .B(n4990), .Z(n5081) );
  NANDN U5356 ( .A(n4993), .B(n4992), .Z(n4997) );
  NAND U5357 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5358 ( .A(n4997), .B(n4996), .Z(n5080) );
  XNOR U5359 ( .A(n5081), .B(n5080), .Z(n5083) );
  NAND U5360 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U5361 ( .A(n5001), .B(n5000), .Z(n5002) );
  AND U5362 ( .A(n5003), .B(n5002), .Z(n5113) );
  AND U5363 ( .A(x[85]), .B(y[232]), .Z(n5879) );
  NAND U5364 ( .A(n5879), .B(n5004), .Z(n5008) );
  NAND U5365 ( .A(n5006), .B(n5005), .Z(n5007) );
  NAND U5366 ( .A(n5008), .B(n5007), .Z(n5177) );
  NAND U5367 ( .A(x[86]), .B(y[227]), .Z(n5153) );
  NAND U5368 ( .A(x[69]), .B(y[244]), .Z(n5151) );
  NAND U5369 ( .A(x[81]), .B(y[232]), .Z(n5152) );
  XOR U5370 ( .A(n5151), .B(n5152), .Z(n5154) );
  XOR U5371 ( .A(n5153), .B(n5154), .Z(n5176) );
  AND U5372 ( .A(y[229]), .B(x[84]), .Z(n5010) );
  NAND U5373 ( .A(y[228]), .B(x[85]), .Z(n5009) );
  XNOR U5374 ( .A(n5010), .B(n5009), .Z(n5162) );
  AND U5375 ( .A(x[83]), .B(y[230]), .Z(n5161) );
  XOR U5376 ( .A(n5162), .B(n5161), .Z(n5175) );
  XOR U5377 ( .A(n5177), .B(n5178), .Z(n5111) );
  NANDN U5378 ( .A(n5307), .B(n5160), .Z(n5014) );
  NAND U5379 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U5380 ( .A(n5014), .B(n5013), .Z(n5183) );
  NAND U5381 ( .A(x[79]), .B(y[234]), .Z(n5167) );
  NAND U5382 ( .A(x[82]), .B(y[231]), .Z(n5165) );
  NAND U5383 ( .A(x[70]), .B(y[243]), .Z(n5166) );
  XOR U5384 ( .A(n5165), .B(n5166), .Z(n5168) );
  XOR U5385 ( .A(n5167), .B(n5168), .Z(n5182) );
  NAND U5386 ( .A(x[87]), .B(y[226]), .Z(n5150) );
  NAND U5387 ( .A(x[68]), .B(y[245]), .Z(n5147) );
  NAND U5388 ( .A(x[80]), .B(y[233]), .Z(n5148) );
  XOR U5389 ( .A(n5147), .B(n5148), .Z(n5149) );
  XNOR U5390 ( .A(n5150), .B(n5149), .Z(n5181) );
  XOR U5391 ( .A(n5183), .B(n5184), .Z(n5110) );
  XNOR U5392 ( .A(n5111), .B(n5110), .Z(n5112) );
  XOR U5393 ( .A(n5113), .B(n5112), .Z(n5125) );
  NAND U5394 ( .A(n5016), .B(n5015), .Z(n5020) );
  NANDN U5395 ( .A(n5018), .B(n5017), .Z(n5019) );
  AND U5396 ( .A(n5020), .B(n5019), .Z(n5123) );
  NAND U5397 ( .A(n5022), .B(n5021), .Z(n5026) );
  NANDN U5398 ( .A(n5024), .B(n5023), .Z(n5025) );
  NAND U5399 ( .A(n5026), .B(n5025), .Z(n5122) );
  XNOR U5400 ( .A(n5123), .B(n5122), .Z(n5124) );
  XNOR U5401 ( .A(n5125), .B(n5124), .Z(n5082) );
  XOR U5402 ( .A(n5083), .B(n5082), .Z(n5063) );
  NAND U5403 ( .A(n5028), .B(n5027), .Z(n5032) );
  NAND U5404 ( .A(n5030), .B(n5029), .Z(n5031) );
  NAND U5405 ( .A(n5032), .B(n5031), .Z(n5062) );
  XNOR U5406 ( .A(n5063), .B(n5062), .Z(n5065) );
  XOR U5407 ( .A(n5064), .B(n5065), .Z(n5058) );
  XOR U5408 ( .A(n5059), .B(n5058), .Z(n5047) );
  XNOR U5409 ( .A(n5048), .B(n5047), .Z(n5049) );
  XOR U5410 ( .A(n5050), .B(n5049), .Z(n5055) );
  NANDN U5411 ( .A(n5034), .B(n5033), .Z(n5038) );
  NAND U5412 ( .A(n5036), .B(n5035), .Z(n5037) );
  NAND U5413 ( .A(n5038), .B(n5037), .Z(n5054) );
  NANDN U5414 ( .A(n5039), .B(n5040), .Z(n5045) );
  NOR U5415 ( .A(n5041), .B(n5040), .Z(n5043) );
  OR U5416 ( .A(n5043), .B(n5042), .Z(n5044) );
  AND U5417 ( .A(n5045), .B(n5044), .Z(n5053) );
  XOR U5418 ( .A(n5054), .B(n5053), .Z(n5046) );
  XNOR U5419 ( .A(n5055), .B(n5046), .Z(N122) );
  NANDN U5420 ( .A(n5048), .B(n5047), .Z(n5052) );
  NAND U5421 ( .A(n5050), .B(n5049), .Z(n5051) );
  NAND U5422 ( .A(n5052), .B(n5051), .Z(n5335) );
  IV U5423 ( .A(n5335), .Z(n5333) );
  NANDN U5424 ( .A(n5057), .B(n5056), .Z(n5061) );
  NAND U5425 ( .A(n5059), .B(n5058), .Z(n5060) );
  AND U5426 ( .A(n5061), .B(n5060), .Z(n5327) );
  NANDN U5427 ( .A(n5063), .B(n5062), .Z(n5067) );
  NAND U5428 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5429 ( .A(n5067), .B(n5066), .Z(n5328) );
  XNOR U5430 ( .A(n5327), .B(n5328), .Z(n5330) );
  NAND U5431 ( .A(n5069), .B(n5068), .Z(n5073) );
  NANDN U5432 ( .A(n5071), .B(n5070), .Z(n5072) );
  AND U5433 ( .A(n5073), .B(n5072), .Z(n5188) );
  NANDN U5434 ( .A(n5075), .B(n5074), .Z(n5079) );
  NANDN U5435 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5436 ( .A(n5079), .B(n5078), .Z(n5189) );
  XNOR U5437 ( .A(n5188), .B(n5189), .Z(n5191) );
  NANDN U5438 ( .A(n5081), .B(n5080), .Z(n5085) );
  NAND U5439 ( .A(n5083), .B(n5082), .Z(n5084) );
  AND U5440 ( .A(n5085), .B(n5084), .Z(n5197) );
  AND U5441 ( .A(x[66]), .B(y[248]), .Z(n5208) );
  XOR U5442 ( .A(n5209), .B(n5208), .Z(n5211) );
  NAND U5443 ( .A(x[88]), .B(y[226]), .Z(n5210) );
  XNOR U5444 ( .A(n5211), .B(n5210), .Z(n5251) );
  NANDN U5445 ( .A(n5087), .B(n5086), .Z(n5091) );
  OR U5446 ( .A(n5089), .B(n5088), .Z(n5090) );
  AND U5447 ( .A(n5091), .B(n5090), .Z(n5250) );
  XOR U5448 ( .A(n5251), .B(n5250), .Z(n5253) );
  NANDN U5449 ( .A(n5093), .B(n5092), .Z(n5097) );
  NANDN U5450 ( .A(n5095), .B(n5094), .Z(n5096) );
  AND U5451 ( .A(n5097), .B(n5096), .Z(n5252) );
  XOR U5452 ( .A(n5253), .B(n5252), .Z(n5284) );
  NAND U5453 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U5454 ( .A(n5101), .B(n5100), .Z(n5102) );
  AND U5455 ( .A(n5103), .B(n5102), .Z(n5283) );
  NANDN U5456 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U5457 ( .A(n5107), .B(n5106), .Z(n5108) );
  AND U5458 ( .A(n5109), .B(n5108), .Z(n5285) );
  XOR U5459 ( .A(n5286), .B(n5285), .Z(n5280) );
  NANDN U5460 ( .A(n5111), .B(n5110), .Z(n5115) );
  NAND U5461 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5462 ( .A(n5115), .B(n5114), .Z(n5277) );
  NANDN U5463 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U5464 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U5465 ( .A(n5121), .B(n5120), .Z(n5278) );
  XOR U5466 ( .A(n5277), .B(n5278), .Z(n5279) );
  XOR U5467 ( .A(n5280), .B(n5279), .Z(n5195) );
  NANDN U5468 ( .A(n5123), .B(n5122), .Z(n5127) );
  NANDN U5469 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U5470 ( .A(n5127), .B(n5126), .Z(n5273) );
  AND U5471 ( .A(x[76]), .B(y[238]), .Z(n5402) );
  AND U5472 ( .A(x[69]), .B(y[245]), .Z(n5260) );
  XOR U5473 ( .A(n5402), .B(n5260), .Z(n5262) );
  NAND U5474 ( .A(x[74]), .B(y[240]), .Z(n5261) );
  XNOR U5475 ( .A(n5262), .B(n5261), .Z(n5292) );
  AND U5476 ( .A(x[71]), .B(y[243]), .Z(n5290) );
  NAND U5477 ( .A(y[244]), .B(x[70]), .Z(n5128) );
  XNOR U5478 ( .A(n5537), .B(n5128), .Z(n5308) );
  NAND U5479 ( .A(x[73]), .B(y[241]), .Z(n5309) );
  XNOR U5480 ( .A(n5308), .B(n5309), .Z(n5289) );
  XOR U5481 ( .A(n5290), .B(n5289), .Z(n5291) );
  XOR U5482 ( .A(n5292), .B(n5291), .Z(n5234) );
  NANDN U5483 ( .A(n5130), .B(n5129), .Z(n5134) );
  NANDN U5484 ( .A(n5132), .B(n5131), .Z(n5133) );
  NAND U5485 ( .A(n5134), .B(n5133), .Z(n5233) );
  NANDN U5486 ( .A(n5136), .B(n5135), .Z(n5140) );
  NANDN U5487 ( .A(n5138), .B(n5137), .Z(n5139) );
  NAND U5488 ( .A(n5140), .B(n5139), .Z(n5232) );
  XNOR U5489 ( .A(n5233), .B(n5232), .Z(n5235) );
  NAND U5490 ( .A(n5142), .B(n5141), .Z(n5146) );
  NANDN U5491 ( .A(n5144), .B(n5143), .Z(n5145) );
  AND U5492 ( .A(n5146), .B(n5145), .Z(n5238) );
  XOR U5493 ( .A(n5201), .B(n5200), .Z(n5202) );
  ANDN U5494 ( .B(o[57]), .A(n5155), .Z(n5301) );
  NAND U5495 ( .A(x[78]), .B(y[236]), .Z(n5302) );
  XNOR U5496 ( .A(n5301), .B(n5302), .Z(n5303) );
  NAND U5497 ( .A(x[65]), .B(y[249]), .Z(n5304) );
  XNOR U5498 ( .A(n5303), .B(n5304), .Z(n5255) );
  NAND U5499 ( .A(x[89]), .B(y[225]), .Z(n5312) );
  XNOR U5500 ( .A(o[58]), .B(n5312), .Z(n5265) );
  NAND U5501 ( .A(x[90]), .B(y[224]), .Z(n5266) );
  XNOR U5502 ( .A(n5265), .B(n5266), .Z(n5268) );
  AND U5503 ( .A(x[64]), .B(y[250]), .Z(n5267) );
  XOR U5504 ( .A(n5268), .B(n5267), .Z(n5254) );
  XOR U5505 ( .A(n5255), .B(n5254), .Z(n5257) );
  XOR U5506 ( .A(n5257), .B(n5256), .Z(n5203) );
  XNOR U5507 ( .A(n5202), .B(n5203), .Z(n5246) );
  AND U5508 ( .A(x[85]), .B(y[229]), .Z(n5296) );
  NAND U5509 ( .A(n5296), .B(n5160), .Z(n5164) );
  NAND U5510 ( .A(n5162), .B(n5161), .Z(n5163) );
  NAND U5511 ( .A(n5164), .B(n5163), .Z(n5228) );
  XOR U5512 ( .A(n5296), .B(n5295), .Z(n5298) );
  NAND U5513 ( .A(x[84]), .B(y[230]), .Z(n5297) );
  XNOR U5514 ( .A(n5298), .B(n5297), .Z(n5227) );
  NAND U5515 ( .A(x[87]), .B(y[227]), .Z(n5215) );
  XNOR U5516 ( .A(n5214), .B(n5215), .Z(n5217) );
  AND U5517 ( .A(x[86]), .B(y[228]), .Z(n5216) );
  XOR U5518 ( .A(n5217), .B(n5216), .Z(n5226) );
  XOR U5519 ( .A(n5227), .B(n5226), .Z(n5229) );
  XOR U5520 ( .A(n5228), .B(n5229), .Z(n5245) );
  AND U5521 ( .A(x[75]), .B(y[239]), .Z(n5313) );
  NAND U5522 ( .A(x[83]), .B(y[231]), .Z(n5314) );
  XNOR U5523 ( .A(n5313), .B(n5314), .Z(n5315) );
  NAND U5524 ( .A(x[67]), .B(y[247]), .Z(n5316) );
  XNOR U5525 ( .A(n5315), .B(n5316), .Z(n5205) );
  NAND U5526 ( .A(x[68]), .B(y[246]), .Z(n5221) );
  XNOR U5527 ( .A(n5220), .B(n5221), .Z(n5223) );
  XOR U5528 ( .A(n5223), .B(n5222), .Z(n5204) );
  XOR U5529 ( .A(n5205), .B(n5204), .Z(n5206) );
  XNOR U5530 ( .A(n5206), .B(n5207), .Z(n5244) );
  XOR U5531 ( .A(n5246), .B(n5247), .Z(n5241) );
  XNOR U5532 ( .A(n5240), .B(n5241), .Z(n5272) );
  NANDN U5533 ( .A(n5170), .B(n5169), .Z(n5174) );
  NANDN U5534 ( .A(n5172), .B(n5171), .Z(n5173) );
  NAND U5535 ( .A(n5174), .B(n5173), .Z(n5323) );
  NANDN U5536 ( .A(n5176), .B(n5175), .Z(n5180) );
  NAND U5537 ( .A(n5178), .B(n5177), .Z(n5179) );
  NAND U5538 ( .A(n5180), .B(n5179), .Z(n5322) );
  NANDN U5539 ( .A(n5182), .B(n5181), .Z(n5186) );
  NANDN U5540 ( .A(n5184), .B(n5183), .Z(n5185) );
  NAND U5541 ( .A(n5186), .B(n5185), .Z(n5321) );
  XOR U5542 ( .A(n5322), .B(n5321), .Z(n5324) );
  XOR U5543 ( .A(n5323), .B(n5324), .Z(n5271) );
  XOR U5544 ( .A(n5273), .B(n5274), .Z(n5194) );
  XNOR U5545 ( .A(n5195), .B(n5194), .Z(n5196) );
  XNOR U5546 ( .A(n5197), .B(n5196), .Z(n5190) );
  XOR U5547 ( .A(n5191), .B(n5190), .Z(n5329) );
  XOR U5548 ( .A(n5330), .B(n5329), .Z(n5336) );
  XNOR U5549 ( .A(n5334), .B(n5336), .Z(n5187) );
  XOR U5550 ( .A(n5333), .B(n5187), .Z(N123) );
  NANDN U5551 ( .A(n5189), .B(n5188), .Z(n5193) );
  NAND U5552 ( .A(n5191), .B(n5190), .Z(n5192) );
  AND U5553 ( .A(n5193), .B(n5192), .Z(n5344) );
  NANDN U5554 ( .A(n5195), .B(n5194), .Z(n5199) );
  NANDN U5555 ( .A(n5197), .B(n5196), .Z(n5198) );
  AND U5556 ( .A(n5199), .B(n5198), .Z(n5342) );
  NAND U5557 ( .A(n5209), .B(n5208), .Z(n5213) );
  ANDN U5558 ( .B(n5211), .A(n5210), .Z(n5212) );
  ANDN U5559 ( .B(n5213), .A(n5212), .Z(n5375) );
  NANDN U5560 ( .A(n5215), .B(n5214), .Z(n5219) );
  NAND U5561 ( .A(n5217), .B(n5216), .Z(n5218) );
  NAND U5562 ( .A(n5219), .B(n5218), .Z(n5374) );
  XNOR U5563 ( .A(n5375), .B(n5374), .Z(n5376) );
  NANDN U5564 ( .A(n5221), .B(n5220), .Z(n5225) );
  NAND U5565 ( .A(n5223), .B(n5222), .Z(n5224) );
  AND U5566 ( .A(n5225), .B(n5224), .Z(n5389) );
  AND U5567 ( .A(x[64]), .B(y[251]), .Z(n5459) );
  NAND U5568 ( .A(x[91]), .B(y[224]), .Z(n5460) );
  XNOR U5569 ( .A(n5459), .B(n5460), .Z(n5462) );
  NAND U5570 ( .A(x[90]), .B(y[225]), .Z(n5450) );
  XNOR U5571 ( .A(o[59]), .B(n5450), .Z(n5461) );
  XOR U5572 ( .A(n5462), .B(n5461), .Z(n5386) );
  AND U5573 ( .A(x[73]), .B(y[242]), .Z(n5444) );
  NAND U5574 ( .A(x[85]), .B(y[230]), .Z(n5445) );
  XNOR U5575 ( .A(n5444), .B(n5445), .Z(n5446) );
  NAND U5576 ( .A(x[82]), .B(y[233]), .Z(n5447) );
  XOR U5577 ( .A(n5446), .B(n5447), .Z(n5387) );
  XNOR U5578 ( .A(n5386), .B(n5387), .Z(n5388) );
  XOR U5579 ( .A(n5389), .B(n5388), .Z(n5377) );
  XNOR U5580 ( .A(n5376), .B(n5377), .Z(n5468) );
  XOR U5581 ( .A(n5467), .B(n5468), .Z(n5470) );
  XOR U5582 ( .A(n5469), .B(n5470), .Z(n5486) );
  NAND U5583 ( .A(n5227), .B(n5226), .Z(n5231) );
  NAND U5584 ( .A(n5229), .B(n5228), .Z(n5230) );
  AND U5585 ( .A(n5231), .B(n5230), .Z(n5484) );
  NAND U5586 ( .A(n5233), .B(n5232), .Z(n5237) );
  NANDN U5587 ( .A(n5235), .B(n5234), .Z(n5236) );
  AND U5588 ( .A(n5237), .B(n5236), .Z(n5483) );
  XOR U5589 ( .A(n5484), .B(n5483), .Z(n5485) );
  NANDN U5590 ( .A(n5239), .B(n5238), .Z(n5243) );
  NANDN U5591 ( .A(n5241), .B(n5240), .Z(n5242) );
  AND U5592 ( .A(n5243), .B(n5242), .Z(n5474) );
  NANDN U5593 ( .A(n5245), .B(n5244), .Z(n5249) );
  NANDN U5594 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U5595 ( .A(n5249), .B(n5248), .Z(n5472) );
  AND U5596 ( .A(x[79]), .B(y[236]), .Z(n5407) );
  AND U5597 ( .A(x[66]), .B(y[249]), .Z(n5408) );
  XOR U5598 ( .A(n5407), .B(n5408), .Z(n5409) );
  AND U5599 ( .A(x[67]), .B(y[248]), .Z(n5410) );
  XOR U5600 ( .A(n5409), .B(n5410), .Z(n5427) );
  AND U5601 ( .A(x[83]), .B(y[232]), .Z(n5438) );
  NAND U5602 ( .A(x[89]), .B(y[226]), .Z(n5439) );
  XNOR U5603 ( .A(n5438), .B(n5439), .Z(n5440) );
  NAND U5604 ( .A(x[70]), .B(y[245]), .Z(n5441) );
  XOR U5605 ( .A(n5440), .B(n5441), .Z(n5428) );
  XNOR U5606 ( .A(n5427), .B(n5428), .Z(n5429) );
  NAND U5607 ( .A(x[80]), .B(y[235]), .Z(n5393) );
  XOR U5608 ( .A(n5393), .B(n5392), .Z(n5395) );
  XOR U5609 ( .A(n5394), .B(n5395), .Z(n5404) );
  AND U5610 ( .A(y[238]), .B(x[77]), .Z(n5259) );
  NAND U5611 ( .A(y[239]), .B(x[76]), .Z(n5258) );
  XNOR U5612 ( .A(n5259), .B(n5258), .Z(n5403) );
  XOR U5613 ( .A(n5404), .B(n5403), .Z(n5430) );
  XNOR U5614 ( .A(n5429), .B(n5430), .Z(n5370) );
  NAND U5615 ( .A(n5402), .B(n5260), .Z(n5264) );
  ANDN U5616 ( .B(n5262), .A(n5261), .Z(n5263) );
  ANDN U5617 ( .B(n5264), .A(n5263), .Z(n5369) );
  NANDN U5618 ( .A(n5266), .B(n5265), .Z(n5270) );
  NAND U5619 ( .A(n5268), .B(n5267), .Z(n5269) );
  NAND U5620 ( .A(n5270), .B(n5269), .Z(n5368) );
  XOR U5621 ( .A(n5369), .B(n5368), .Z(n5371) );
  XNOR U5622 ( .A(n5370), .B(n5371), .Z(n5464) );
  XOR U5623 ( .A(n5463), .B(n5464), .Z(n5466) );
  XOR U5624 ( .A(n5465), .B(n5466), .Z(n5471) );
  XOR U5625 ( .A(n5472), .B(n5471), .Z(n5473) );
  XOR U5626 ( .A(n5474), .B(n5473), .Z(n5350) );
  NANDN U5627 ( .A(n5272), .B(n5271), .Z(n5276) );
  NAND U5628 ( .A(n5274), .B(n5273), .Z(n5275) );
  NAND U5629 ( .A(n5276), .B(n5275), .Z(n5352) );
  XOR U5630 ( .A(n5353), .B(n5352), .Z(n5359) );
  NAND U5631 ( .A(n5278), .B(n5277), .Z(n5282) );
  NAND U5632 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U5633 ( .A(n5282), .B(n5281), .Z(n5356) );
  NANDN U5634 ( .A(n5284), .B(n5283), .Z(n5288) );
  NAND U5635 ( .A(n5286), .B(n5285), .Z(n5287) );
  NAND U5636 ( .A(n5288), .B(n5287), .Z(n5363) );
  NAND U5637 ( .A(n5290), .B(n5289), .Z(n5294) );
  NAND U5638 ( .A(n5292), .B(n5291), .Z(n5293) );
  NAND U5639 ( .A(n5294), .B(n5293), .Z(n5479) );
  NAND U5640 ( .A(n5296), .B(n5295), .Z(n5300) );
  ANDN U5641 ( .B(n5298), .A(n5297), .Z(n5299) );
  ANDN U5642 ( .B(n5300), .A(n5299), .Z(n5420) );
  NANDN U5643 ( .A(n5302), .B(n5301), .Z(n5306) );
  NANDN U5644 ( .A(n5304), .B(n5303), .Z(n5305) );
  NAND U5645 ( .A(n5306), .B(n5305), .Z(n5419) );
  XNOR U5646 ( .A(n5420), .B(n5419), .Z(n5422) );
  AND U5647 ( .A(y[244]), .B(x[72]), .Z(n5452) );
  NANDN U5648 ( .A(n5307), .B(n5452), .Z(n5311) );
  NANDN U5649 ( .A(n5309), .B(n5308), .Z(n5310) );
  NAND U5650 ( .A(n5311), .B(n5310), .Z(n5383) );
  ANDN U5651 ( .B(o[58]), .A(n5312), .Z(n5415) );
  AND U5652 ( .A(x[78]), .B(y[237]), .Z(n5414) );
  AND U5653 ( .A(x[65]), .B(y[250]), .Z(n5413) );
  XOR U5654 ( .A(n5414), .B(n5413), .Z(n5416) );
  XOR U5655 ( .A(n5415), .B(n5416), .Z(n5380) );
  AND U5656 ( .A(x[81]), .B(y[234]), .Z(n5453) );
  NAND U5657 ( .A(x[68]), .B(y[247]), .Z(n5454) );
  XNOR U5658 ( .A(n5453), .B(n5454), .Z(n5456) );
  AND U5659 ( .A(x[69]), .B(y[246]), .Z(n5455) );
  XOR U5660 ( .A(n5456), .B(n5455), .Z(n5381) );
  XOR U5661 ( .A(n5380), .B(n5381), .Z(n5382) );
  XOR U5662 ( .A(n5383), .B(n5382), .Z(n5421) );
  XOR U5663 ( .A(n5422), .B(n5421), .Z(n5478) );
  NANDN U5664 ( .A(n5314), .B(n5313), .Z(n5318) );
  NANDN U5665 ( .A(n5316), .B(n5315), .Z(n5317) );
  AND U5666 ( .A(n5318), .B(n5317), .Z(n5426) );
  NAND U5667 ( .A(y[227]), .B(x[88]), .Z(n5319) );
  XNOR U5668 ( .A(n5320), .B(n5319), .Z(n5434) );
  NAND U5669 ( .A(x[71]), .B(y[244]), .Z(n5435) );
  XNOR U5670 ( .A(n5434), .B(n5435), .Z(n5424) );
  AND U5671 ( .A(x[72]), .B(y[243]), .Z(n5396) );
  AND U5672 ( .A(x[87]), .B(y[228]), .Z(n5397) );
  XOR U5673 ( .A(n5396), .B(n5397), .Z(n5398) );
  AND U5674 ( .A(x[86]), .B(y[229]), .Z(n5399) );
  XOR U5675 ( .A(n5398), .B(n5399), .Z(n5423) );
  XOR U5676 ( .A(n5424), .B(n5423), .Z(n5425) );
  XNOR U5677 ( .A(n5426), .B(n5425), .Z(n5477) );
  XOR U5678 ( .A(n5478), .B(n5477), .Z(n5480) );
  XNOR U5679 ( .A(n5479), .B(n5480), .Z(n5362) );
  XOR U5680 ( .A(n5363), .B(n5362), .Z(n5365) );
  NAND U5681 ( .A(n5322), .B(n5321), .Z(n5326) );
  NAND U5682 ( .A(n5324), .B(n5323), .Z(n5325) );
  AND U5683 ( .A(n5326), .B(n5325), .Z(n5364) );
  XOR U5684 ( .A(n5365), .B(n5364), .Z(n5357) );
  XOR U5685 ( .A(n5356), .B(n5357), .Z(n5358) );
  XOR U5686 ( .A(n5342), .B(n5341), .Z(n5343) );
  XOR U5687 ( .A(n5344), .B(n5343), .Z(n5349) );
  NANDN U5688 ( .A(n5328), .B(n5327), .Z(n5332) );
  NAND U5689 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5690 ( .A(n5332), .B(n5331), .Z(n5348) );
  NANDN U5691 ( .A(n5333), .B(n5334), .Z(n5339) );
  NOR U5692 ( .A(n5335), .B(n5334), .Z(n5337) );
  OR U5693 ( .A(n5337), .B(n5336), .Z(n5338) );
  AND U5694 ( .A(n5339), .B(n5338), .Z(n5347) );
  XOR U5695 ( .A(n5348), .B(n5347), .Z(n5340) );
  XNOR U5696 ( .A(n5349), .B(n5340), .Z(N124) );
  NAND U5697 ( .A(n5342), .B(n5341), .Z(n5346) );
  NAND U5698 ( .A(n5344), .B(n5343), .Z(n5345) );
  NAND U5699 ( .A(n5346), .B(n5345), .Z(n5498) );
  IV U5700 ( .A(n5498), .Z(n5496) );
  NANDN U5701 ( .A(n5351), .B(n5350), .Z(n5355) );
  NAND U5702 ( .A(n5353), .B(n5352), .Z(n5354) );
  NAND U5703 ( .A(n5355), .B(n5354), .Z(n5490) );
  NAND U5704 ( .A(n5357), .B(n5356), .Z(n5361) );
  NANDN U5705 ( .A(n5359), .B(n5358), .Z(n5360) );
  AND U5706 ( .A(n5361), .B(n5360), .Z(n5491) );
  XOR U5707 ( .A(n5490), .B(n5491), .Z(n5493) );
  NAND U5708 ( .A(n5363), .B(n5362), .Z(n5367) );
  NAND U5709 ( .A(n5365), .B(n5364), .Z(n5366) );
  AND U5710 ( .A(n5367), .B(n5366), .Z(n5503) );
  NANDN U5711 ( .A(n5369), .B(n5368), .Z(n5373) );
  NANDN U5712 ( .A(n5371), .B(n5370), .Z(n5372) );
  AND U5713 ( .A(n5373), .B(n5372), .Z(n5516) );
  NANDN U5714 ( .A(n5375), .B(n5374), .Z(n5379) );
  NANDN U5715 ( .A(n5377), .B(n5376), .Z(n5378) );
  AND U5716 ( .A(n5379), .B(n5378), .Z(n5619) );
  NAND U5717 ( .A(n5381), .B(n5380), .Z(n5385) );
  NAND U5718 ( .A(n5383), .B(n5382), .Z(n5384) );
  AND U5719 ( .A(n5385), .B(n5384), .Z(n5617) );
  NANDN U5720 ( .A(n5387), .B(n5386), .Z(n5391) );
  NANDN U5721 ( .A(n5389), .B(n5388), .Z(n5390) );
  NAND U5722 ( .A(n5391), .B(n5390), .Z(n5616) );
  XNOR U5723 ( .A(n5617), .B(n5616), .Z(n5618) );
  XNOR U5724 ( .A(n5619), .B(n5618), .Z(n5515) );
  XNOR U5725 ( .A(n5516), .B(n5515), .Z(n5518) );
  AND U5726 ( .A(x[71]), .B(y[245]), .Z(n5561) );
  AND U5727 ( .A(x[76]), .B(y[240]), .Z(n5560) );
  XOR U5728 ( .A(n5561), .B(n5560), .Z(n5563) );
  AND U5729 ( .A(x[75]), .B(y[241]), .Z(n5562) );
  XOR U5730 ( .A(n5563), .B(n5562), .Z(n5593) );
  AND U5731 ( .A(x[91]), .B(y[225]), .Z(n5572) );
  XOR U5732 ( .A(o[60]), .B(n5572), .Z(n5581) );
  AND U5733 ( .A(x[90]), .B(y[226]), .Z(n5580) );
  XOR U5734 ( .A(n5581), .B(n5580), .Z(n5583) );
  AND U5735 ( .A(x[79]), .B(y[237]), .Z(n5582) );
  XNOR U5736 ( .A(n5583), .B(n5582), .Z(n5592) );
  XOR U5737 ( .A(n5594), .B(n5595), .Z(n5623) );
  NAND U5738 ( .A(n5397), .B(n5396), .Z(n5401) );
  NAND U5739 ( .A(n5399), .B(n5398), .Z(n5400) );
  NAND U5740 ( .A(n5401), .B(n5400), .Z(n5600) );
  AND U5741 ( .A(x[81]), .B(y[235]), .Z(n5526) );
  AND U5742 ( .A(x[86]), .B(y[230]), .Z(n5525) );
  XOR U5743 ( .A(n5526), .B(n5525), .Z(n5528) );
  AND U5744 ( .A(x[68]), .B(y[248]), .Z(n5527) );
  XOR U5745 ( .A(n5528), .B(n5527), .Z(n5599) );
  AND U5746 ( .A(x[70]), .B(y[246]), .Z(n5758) );
  AND U5747 ( .A(x[83]), .B(y[233]), .Z(n5573) );
  XOR U5748 ( .A(n5758), .B(n5573), .Z(n5574) );
  XOR U5749 ( .A(n5575), .B(n5574), .Z(n5598) );
  XOR U5750 ( .A(n5599), .B(n5598), .Z(n5601) );
  XOR U5751 ( .A(n5600), .B(n5601), .Z(n5622) );
  XOR U5752 ( .A(n5623), .B(n5622), .Z(n5625) );
  NAND U5753 ( .A(n5402), .B(n5587), .Z(n5406) );
  NANDN U5754 ( .A(n5404), .B(n5403), .Z(n5405) );
  NAND U5755 ( .A(n5406), .B(n5405), .Z(n5521) );
  NAND U5756 ( .A(n5408), .B(n5407), .Z(n5412) );
  NAND U5757 ( .A(n5410), .B(n5409), .Z(n5411) );
  NAND U5758 ( .A(n5412), .B(n5411), .Z(n5520) );
  NAND U5759 ( .A(n5414), .B(n5413), .Z(n5418) );
  NAND U5760 ( .A(n5416), .B(n5415), .Z(n5417) );
  NAND U5761 ( .A(n5418), .B(n5417), .Z(n5519) );
  XOR U5762 ( .A(n5520), .B(n5519), .Z(n5522) );
  XOR U5763 ( .A(n5521), .B(n5522), .Z(n5624) );
  XOR U5764 ( .A(n5625), .B(n5624), .Z(n5517) );
  XOR U5765 ( .A(n5518), .B(n5517), .Z(n5651) );
  NANDN U5766 ( .A(n5428), .B(n5427), .Z(n5432) );
  NANDN U5767 ( .A(n5430), .B(n5429), .Z(n5431) );
  NAND U5768 ( .A(n5432), .B(n5431), .Z(n5604) );
  XNOR U5769 ( .A(n5605), .B(n5604), .Z(n5606) );
  XOR U5770 ( .A(n5607), .B(n5606), .Z(n5648) );
  AND U5771 ( .A(x[88]), .B(y[231]), .Z(n5954) );
  NAND U5772 ( .A(n5433), .B(n5954), .Z(n5437) );
  NANDN U5773 ( .A(n5435), .B(n5434), .Z(n5436) );
  NAND U5774 ( .A(n5437), .B(n5436), .Z(n5640) );
  AND U5775 ( .A(x[89]), .B(y[227]), .Z(n5556) );
  XOR U5776 ( .A(n5557), .B(n5556), .Z(n5555) );
  AND U5777 ( .A(x[65]), .B(y[251]), .Z(n5554) );
  XOR U5778 ( .A(n5555), .B(n5554), .Z(n5639) );
  AND U5779 ( .A(x[80]), .B(y[236]), .Z(n5549) );
  AND U5780 ( .A(x[88]), .B(y[228]), .Z(n5548) );
  XOR U5781 ( .A(n5549), .B(n5548), .Z(n5551) );
  AND U5782 ( .A(x[66]), .B(y[250]), .Z(n5550) );
  XOR U5783 ( .A(n5551), .B(n5550), .Z(n5638) );
  XOR U5784 ( .A(n5639), .B(n5638), .Z(n5641) );
  XNOR U5785 ( .A(n5640), .B(n5641), .Z(n5613) );
  NANDN U5786 ( .A(n5439), .B(n5438), .Z(n5443) );
  NANDN U5787 ( .A(n5441), .B(n5440), .Z(n5442) );
  NAND U5788 ( .A(n5443), .B(n5442), .Z(n5634) );
  AND U5789 ( .A(x[67]), .B(y[249]), .Z(n5586) );
  XOR U5790 ( .A(n5587), .B(n5586), .Z(n5589) );
  AND U5791 ( .A(x[87]), .B(y[229]), .Z(n5588) );
  XOR U5792 ( .A(n5589), .B(n5588), .Z(n5633) );
  AND U5793 ( .A(x[69]), .B(y[247]), .Z(n5567) );
  AND U5794 ( .A(x[85]), .B(y[231]), .Z(n5566) );
  XOR U5795 ( .A(n5567), .B(n5566), .Z(n5569) );
  AND U5796 ( .A(x[84]), .B(y[232]), .Z(n5568) );
  XOR U5797 ( .A(n5569), .B(n5568), .Z(n5632) );
  XOR U5798 ( .A(n5633), .B(n5632), .Z(n5635) );
  XNOR U5799 ( .A(n5634), .B(n5635), .Z(n5611) );
  NANDN U5800 ( .A(n5445), .B(n5444), .Z(n5449) );
  NANDN U5801 ( .A(n5447), .B(n5446), .Z(n5448) );
  NAND U5802 ( .A(n5449), .B(n5448), .Z(n5544) );
  ANDN U5803 ( .B(o[59]), .A(n5450), .Z(n5534) );
  AND U5804 ( .A(x[64]), .B(y[252]), .Z(n5532) );
  AND U5805 ( .A(x[92]), .B(y[224]), .Z(n5531) );
  XOR U5806 ( .A(n5532), .B(n5531), .Z(n5533) );
  XOR U5807 ( .A(n5534), .B(n5533), .Z(n5543) );
  NAND U5808 ( .A(y[242]), .B(x[74]), .Z(n5451) );
  XNOR U5809 ( .A(n5452), .B(n5451), .Z(n5539) );
  AND U5810 ( .A(x[73]), .B(y[243]), .Z(n5538) );
  XOR U5811 ( .A(n5539), .B(n5538), .Z(n5542) );
  XOR U5812 ( .A(n5543), .B(n5542), .Z(n5545) );
  XOR U5813 ( .A(n5544), .B(n5545), .Z(n5629) );
  NANDN U5814 ( .A(n5454), .B(n5453), .Z(n5458) );
  NAND U5815 ( .A(n5456), .B(n5455), .Z(n5457) );
  NAND U5816 ( .A(n5458), .B(n5457), .Z(n5627) );
  XOR U5817 ( .A(n5627), .B(n5626), .Z(n5628) );
  XNOR U5818 ( .A(n5629), .B(n5628), .Z(n5610) );
  XOR U5819 ( .A(n5611), .B(n5610), .Z(n5612) );
  XOR U5820 ( .A(n5613), .B(n5612), .Z(n5649) );
  XOR U5821 ( .A(n5648), .B(n5649), .Z(n5650) );
  XOR U5822 ( .A(n5651), .B(n5650), .Z(n5646) );
  XNOR U5823 ( .A(n5644), .B(n5645), .Z(n5647) );
  XOR U5824 ( .A(n5646), .B(n5647), .Z(n5504) );
  NAND U5825 ( .A(n5472), .B(n5471), .Z(n5476) );
  NAND U5826 ( .A(n5474), .B(n5473), .Z(n5475) );
  NAND U5827 ( .A(n5476), .B(n5475), .Z(n5511) );
  NAND U5828 ( .A(n5478), .B(n5477), .Z(n5482) );
  NAND U5829 ( .A(n5480), .B(n5479), .Z(n5481) );
  NAND U5830 ( .A(n5482), .B(n5481), .Z(n5509) );
  NAND U5831 ( .A(n5484), .B(n5483), .Z(n5488) );
  NANDN U5832 ( .A(n5486), .B(n5485), .Z(n5487) );
  AND U5833 ( .A(n5488), .B(n5487), .Z(n5510) );
  XOR U5834 ( .A(n5509), .B(n5510), .Z(n5512) );
  XOR U5835 ( .A(n5511), .B(n5512), .Z(n5505) );
  XOR U5836 ( .A(n5506), .B(n5505), .Z(n5492) );
  XOR U5837 ( .A(n5493), .B(n5492), .Z(n5499) );
  XNOR U5838 ( .A(n5497), .B(n5499), .Z(n5489) );
  XOR U5839 ( .A(n5496), .B(n5489), .Z(N125) );
  NAND U5840 ( .A(n5491), .B(n5490), .Z(n5495) );
  NAND U5841 ( .A(n5493), .B(n5492), .Z(n5494) );
  AND U5842 ( .A(n5495), .B(n5494), .Z(n5653) );
  NANDN U5843 ( .A(n5496), .B(n5497), .Z(n5502) );
  NOR U5844 ( .A(n5498), .B(n5497), .Z(n5500) );
  OR U5845 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U5846 ( .A(n5502), .B(n5501), .Z(n5654) );
  NANDN U5847 ( .A(n5504), .B(n5503), .Z(n5508) );
  NAND U5848 ( .A(n5506), .B(n5505), .Z(n5507) );
  NAND U5849 ( .A(n5508), .B(n5507), .Z(n5658) );
  NAND U5850 ( .A(n5510), .B(n5509), .Z(n5514) );
  NAND U5851 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5852 ( .A(n5514), .B(n5513), .Z(n5656) );
  NAND U5853 ( .A(n5520), .B(n5519), .Z(n5524) );
  NAND U5854 ( .A(n5522), .B(n5521), .Z(n5523) );
  AND U5855 ( .A(n5524), .B(n5523), .Z(n5786) );
  NAND U5856 ( .A(n5526), .B(n5525), .Z(n5530) );
  NAND U5857 ( .A(n5528), .B(n5527), .Z(n5529) );
  NAND U5858 ( .A(n5530), .B(n5529), .Z(n5824) );
  NAND U5859 ( .A(n5532), .B(n5531), .Z(n5536) );
  NAND U5860 ( .A(n5534), .B(n5533), .Z(n5535) );
  NAND U5861 ( .A(n5536), .B(n5535), .Z(n5823) );
  XOR U5862 ( .A(n5824), .B(n5823), .Z(n5825) );
  AND U5863 ( .A(x[74]), .B(y[244]), .Z(n5822) );
  NAND U5864 ( .A(n5537), .B(n5822), .Z(n5541) );
  NAND U5865 ( .A(n5539), .B(n5538), .Z(n5540) );
  NAND U5866 ( .A(n5541), .B(n5540), .Z(n5792) );
  AND U5867 ( .A(x[76]), .B(y[241]), .Z(n6019) );
  AND U5868 ( .A(x[65]), .B(y[252]), .Z(n5734) );
  XOR U5869 ( .A(n6019), .B(n5734), .Z(n5736) );
  AND U5870 ( .A(x[86]), .B(y[231]), .Z(n5735) );
  XOR U5871 ( .A(n5736), .B(n5735), .Z(n5791) );
  AND U5872 ( .A(x[79]), .B(y[238]), .Z(n5739) );
  XOR U5873 ( .A(n5879), .B(n5739), .Z(n5740) );
  XOR U5874 ( .A(n5741), .B(n5740), .Z(n5790) );
  XOR U5875 ( .A(n5791), .B(n5790), .Z(n5793) );
  XNOR U5876 ( .A(n5792), .B(n5793), .Z(n5826) );
  NAND U5877 ( .A(n5543), .B(n5542), .Z(n5547) );
  NAND U5878 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U5879 ( .A(n5547), .B(n5546), .Z(n5784) );
  XNOR U5880 ( .A(n5786), .B(n5787), .Z(n5781) );
  NAND U5881 ( .A(n5549), .B(n5548), .Z(n5553) );
  NAND U5882 ( .A(n5551), .B(n5550), .Z(n5552) );
  NAND U5883 ( .A(n5553), .B(n5552), .Z(n5797) );
  AND U5884 ( .A(n5555), .B(n5554), .Z(n5559) );
  NAND U5885 ( .A(n5557), .B(n5556), .Z(n5558) );
  NANDN U5886 ( .A(n5559), .B(n5558), .Z(n5796) );
  XOR U5887 ( .A(n5797), .B(n5796), .Z(n5798) );
  NAND U5888 ( .A(n5561), .B(n5560), .Z(n5565) );
  NAND U5889 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U5890 ( .A(n5565), .B(n5564), .Z(n5700) );
  AND U5891 ( .A(x[75]), .B(y[242]), .Z(n5755) );
  AND U5892 ( .A(x[67]), .B(y[250]), .Z(n5753) );
  AND U5893 ( .A(x[81]), .B(y[236]), .Z(n5752) );
  XOR U5894 ( .A(n5753), .B(n5752), .Z(n5754) );
  XOR U5895 ( .A(n5755), .B(n5754), .Z(n5699) );
  AND U5896 ( .A(x[87]), .B(y[230]), .Z(n5922) );
  AND U5897 ( .A(x[77]), .B(y[240]), .Z(n5748) );
  AND U5898 ( .A(x[88]), .B(y[229]), .Z(n5747) );
  XOR U5899 ( .A(n5748), .B(n5747), .Z(n5749) );
  XOR U5900 ( .A(n5922), .B(n5749), .Z(n5698) );
  XOR U5901 ( .A(n5699), .B(n5698), .Z(n5701) );
  XNOR U5902 ( .A(n5700), .B(n5701), .Z(n5799) );
  NAND U5903 ( .A(n5567), .B(n5566), .Z(n5571) );
  NAND U5904 ( .A(n5569), .B(n5568), .Z(n5570) );
  NAND U5905 ( .A(n5571), .B(n5570), .Z(n5767) );
  AND U5906 ( .A(n5572), .B(o[60]), .Z(n5707) );
  AND U5907 ( .A(x[80]), .B(y[237]), .Z(n5705) );
  AND U5908 ( .A(x[91]), .B(y[226]), .Z(n5704) );
  XOR U5909 ( .A(n5705), .B(n5704), .Z(n5706) );
  XOR U5910 ( .A(n5707), .B(n5706), .Z(n5766) );
  AND U5911 ( .A(x[66]), .B(y[251]), .Z(n5716) );
  XOR U5912 ( .A(n5717), .B(n5716), .Z(n5718) );
  XOR U5913 ( .A(n5719), .B(n5718), .Z(n5765) );
  XOR U5914 ( .A(n5766), .B(n5765), .Z(n5768) );
  XOR U5915 ( .A(n5767), .B(n5768), .Z(n5687) );
  NAND U5916 ( .A(n5758), .B(n5573), .Z(n5577) );
  NAND U5917 ( .A(n5575), .B(n5574), .Z(n5576) );
  AND U5918 ( .A(n5577), .B(n5576), .Z(n5804) );
  AND U5919 ( .A(x[92]), .B(y[225]), .Z(n5744) );
  XOR U5920 ( .A(o[61]), .B(n5744), .Z(n5816) );
  AND U5921 ( .A(x[64]), .B(y[253]), .Z(n5814) );
  AND U5922 ( .A(x[93]), .B(y[224]), .Z(n5813) );
  XOR U5923 ( .A(n5814), .B(n5813), .Z(n5815) );
  XOR U5924 ( .A(n5816), .B(n5815), .Z(n5803) );
  AND U5925 ( .A(x[89]), .B(y[228]), .Z(n5731) );
  AND U5926 ( .A(x[90]), .B(y[227]), .Z(n5728) );
  XOR U5927 ( .A(n5729), .B(n5728), .Z(n5730) );
  XNOR U5928 ( .A(n5731), .B(n5730), .Z(n5802) );
  XNOR U5929 ( .A(n5804), .B(n5805), .Z(n5686) );
  AND U5930 ( .A(y[247]), .B(x[70]), .Z(n5579) );
  NAND U5931 ( .A(y[246]), .B(x[71]), .Z(n5578) );
  XNOR U5932 ( .A(n5579), .B(n5578), .Z(n5760) );
  AND U5933 ( .A(x[72]), .B(y[245]), .Z(n5759) );
  XOR U5934 ( .A(n5760), .B(n5759), .Z(n5808) );
  AND U5935 ( .A(x[73]), .B(y[244]), .Z(n5970) );
  XOR U5936 ( .A(n5808), .B(n5970), .Z(n5810) );
  AND U5937 ( .A(x[68]), .B(y[249]), .Z(n5711) );
  AND U5938 ( .A(x[74]), .B(y[243]), .Z(n5710) );
  XOR U5939 ( .A(n5711), .B(n5710), .Z(n5713) );
  AND U5940 ( .A(x[69]), .B(y[248]), .Z(n5712) );
  XOR U5941 ( .A(n5713), .B(n5712), .Z(n5809) );
  XOR U5942 ( .A(n5810), .B(n5809), .Z(n5724) );
  NAND U5943 ( .A(n5581), .B(n5580), .Z(n5585) );
  NAND U5944 ( .A(n5583), .B(n5582), .Z(n5584) );
  NAND U5945 ( .A(n5585), .B(n5584), .Z(n5723) );
  NAND U5946 ( .A(n5587), .B(n5586), .Z(n5591) );
  NAND U5947 ( .A(n5589), .B(n5588), .Z(n5590) );
  NAND U5948 ( .A(n5591), .B(n5590), .Z(n5722) );
  XNOR U5949 ( .A(n5723), .B(n5722), .Z(n5725) );
  NANDN U5950 ( .A(n5593), .B(n5592), .Z(n5597) );
  NANDN U5951 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U5952 ( .A(n5597), .B(n5596), .Z(n5692) );
  XNOR U5953 ( .A(n5694), .B(n5695), .Z(n5779) );
  NAND U5954 ( .A(n5599), .B(n5598), .Z(n5603) );
  NAND U5955 ( .A(n5601), .B(n5600), .Z(n5602) );
  NAND U5956 ( .A(n5603), .B(n5602), .Z(n5778) );
  XNOR U5957 ( .A(n5680), .B(n5679), .Z(n5682) );
  NANDN U5958 ( .A(n5605), .B(n5604), .Z(n5609) );
  NANDN U5959 ( .A(n5607), .B(n5606), .Z(n5608) );
  AND U5960 ( .A(n5609), .B(n5608), .Z(n5673) );
  NAND U5961 ( .A(n5611), .B(n5610), .Z(n5615) );
  NAND U5962 ( .A(n5613), .B(n5612), .Z(n5614) );
  AND U5963 ( .A(n5615), .B(n5614), .Z(n5672) );
  XNOR U5964 ( .A(n5673), .B(n5672), .Z(n5675) );
  NANDN U5965 ( .A(n5617), .B(n5616), .Z(n5621) );
  NANDN U5966 ( .A(n5619), .B(n5618), .Z(n5620) );
  NAND U5967 ( .A(n5621), .B(n5620), .Z(n5669) );
  NAND U5968 ( .A(n5627), .B(n5626), .Z(n5631) );
  NAND U5969 ( .A(n5629), .B(n5628), .Z(n5630) );
  NAND U5970 ( .A(n5631), .B(n5630), .Z(n5773) );
  NAND U5971 ( .A(n5633), .B(n5632), .Z(n5637) );
  NAND U5972 ( .A(n5635), .B(n5634), .Z(n5636) );
  NAND U5973 ( .A(n5637), .B(n5636), .Z(n5772) );
  NAND U5974 ( .A(n5639), .B(n5638), .Z(n5643) );
  NAND U5975 ( .A(n5641), .B(n5640), .Z(n5642) );
  NAND U5976 ( .A(n5643), .B(n5642), .Z(n5771) );
  XOR U5977 ( .A(n5772), .B(n5771), .Z(n5774) );
  XOR U5978 ( .A(n5773), .B(n5774), .Z(n5666) );
  XOR U5979 ( .A(n5667), .B(n5666), .Z(n5668) );
  XOR U5980 ( .A(n5669), .B(n5668), .Z(n5674) );
  XOR U5981 ( .A(n5675), .B(n5674), .Z(n5681) );
  XOR U5982 ( .A(n5682), .B(n5681), .Z(n5664) );
  XNOR U5983 ( .A(n5663), .B(n5662), .Z(n5665) );
  XNOR U5984 ( .A(n5664), .B(n5665), .Z(n5657) );
  XOR U5985 ( .A(n5656), .B(n5657), .Z(n5659) );
  XOR U5986 ( .A(n5658), .B(n5659), .Z(n5655) );
  XNOR U5987 ( .A(n5654), .B(n5655), .Z(n5652) );
  XOR U5988 ( .A(n5653), .B(n5652), .Z(N126) );
  NAND U5989 ( .A(n5657), .B(n5656), .Z(n5661) );
  NAND U5990 ( .A(n5659), .B(n5658), .Z(n5660) );
  AND U5991 ( .A(n5661), .B(n5660), .Z(n6109) );
  XNOR U5992 ( .A(n6110), .B(n6109), .Z(n6112) );
  NAND U5993 ( .A(n5667), .B(n5666), .Z(n5671) );
  NAND U5994 ( .A(n5669), .B(n5668), .Z(n5670) );
  AND U5995 ( .A(n5671), .B(n5670), .Z(n5830) );
  NANDN U5996 ( .A(n5673), .B(n5672), .Z(n5678) );
  IV U5997 ( .A(n5674), .Z(n5676) );
  NANDN U5998 ( .A(n5676), .B(n5675), .Z(n5677) );
  AND U5999 ( .A(n5678), .B(n5677), .Z(n5831) );
  NANDN U6000 ( .A(n5680), .B(n5679), .Z(n5685) );
  IV U6001 ( .A(n5681), .Z(n5683) );
  NANDN U6002 ( .A(n5683), .B(n5682), .Z(n5684) );
  NAND U6003 ( .A(n5685), .B(n5684), .Z(n5832) );
  XOR U6004 ( .A(n5830), .B(n5829), .Z(n6105) );
  NANDN U6005 ( .A(n5687), .B(n5686), .Z(n5691) );
  NANDN U6006 ( .A(n5689), .B(n5688), .Z(n5690) );
  AND U6007 ( .A(n5691), .B(n5690), .Z(n6100) );
  NANDN U6008 ( .A(n5693), .B(n5692), .Z(n5697) );
  NANDN U6009 ( .A(n5695), .B(n5694), .Z(n5696) );
  AND U6010 ( .A(n5697), .B(n5696), .Z(n6091) );
  NAND U6011 ( .A(n5699), .B(n5698), .Z(n5703) );
  NAND U6012 ( .A(n5701), .B(n5700), .Z(n5702) );
  AND U6013 ( .A(n5703), .B(n5702), .Z(n6078) );
  NAND U6014 ( .A(n5705), .B(n5704), .Z(n5709) );
  NAND U6015 ( .A(n5707), .B(n5706), .Z(n5708) );
  AND U6016 ( .A(n5709), .B(n5708), .Z(n6036) );
  NAND U6017 ( .A(n5711), .B(n5710), .Z(n5715) );
  NAND U6018 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U6019 ( .A(n5715), .B(n5714), .Z(n6038) );
  AND U6020 ( .A(x[70]), .B(y[248]), .Z(n6004) );
  AND U6021 ( .A(x[69]), .B(y[249]), .Z(n6005) );
  NAND U6022 ( .A(x[83]), .B(y[235]), .Z(n6006) );
  XOR U6023 ( .A(n6004), .B(n6003), .Z(n5909) );
  AND U6024 ( .A(x[68]), .B(y[250]), .Z(n5883) );
  AND U6025 ( .A(x[67]), .B(y[251]), .Z(n5884) );
  NAND U6026 ( .A(x[82]), .B(y[236]), .Z(n5885) );
  XOR U6027 ( .A(n5883), .B(n5882), .Z(n5911) );
  NAND U6028 ( .A(n5717), .B(n5716), .Z(n5721) );
  NAND U6029 ( .A(n5719), .B(n5718), .Z(n5720) );
  AND U6030 ( .A(n5721), .B(n5720), .Z(n5910) );
  XOR U6031 ( .A(n5909), .B(n5908), .Z(n6037) );
  XOR U6032 ( .A(n6036), .B(n6035), .Z(n6077) );
  XOR U6033 ( .A(n6078), .B(n6077), .Z(n6075) );
  NAND U6034 ( .A(n5723), .B(n5722), .Z(n5727) );
  NANDN U6035 ( .A(n5725), .B(n5724), .Z(n5726) );
  NAND U6036 ( .A(n5727), .B(n5726), .Z(n6076) );
  XOR U6037 ( .A(n6075), .B(n6076), .Z(n6093) );
  NAND U6038 ( .A(n5729), .B(n5728), .Z(n5733) );
  AND U6039 ( .A(n5731), .B(n5730), .Z(n5732) );
  ANDN U6040 ( .B(n5733), .A(n5732), .Z(n6030) );
  NAND U6041 ( .A(n6019), .B(n5734), .Z(n5738) );
  AND U6042 ( .A(n5736), .B(n5735), .Z(n5737) );
  ANDN U6043 ( .B(n5738), .A(n5737), .Z(n6032) );
  NAND U6044 ( .A(n5879), .B(n5739), .Z(n5743) );
  NAND U6045 ( .A(n5741), .B(n5740), .Z(n5742) );
  AND U6046 ( .A(n5743), .B(n5742), .Z(n5846) );
  AND U6047 ( .A(n5744), .B(o[61]), .Z(n5872) );
  AND U6048 ( .A(x[92]), .B(y[226]), .Z(n5874) );
  AND U6049 ( .A(x[80]), .B(y[238]), .Z(n5873) );
  XOR U6050 ( .A(n5874), .B(n5873), .Z(n5871) );
  XOR U6051 ( .A(n5872), .B(n5871), .Z(n5848) );
  AND U6052 ( .A(x[89]), .B(y[229]), .Z(n5921) );
  AND U6053 ( .A(y[230]), .B(x[88]), .Z(n5746) );
  NAND U6054 ( .A(y[231]), .B(x[87]), .Z(n5745) );
  XNOR U6055 ( .A(n5746), .B(n5745), .Z(n5920) );
  XNOR U6056 ( .A(n5921), .B(n5920), .Z(n5847) );
  XNOR U6057 ( .A(n5846), .B(n5845), .Z(n6031) );
  XNOR U6058 ( .A(n6030), .B(n6029), .Z(n6070) );
  NAND U6059 ( .A(n5748), .B(n5747), .Z(n5751) );
  NAND U6060 ( .A(n5922), .B(n5749), .Z(n5750) );
  AND U6061 ( .A(n5751), .B(n5750), .Z(n6060) );
  NAND U6062 ( .A(n5753), .B(n5752), .Z(n5757) );
  NAND U6063 ( .A(n5755), .B(n5754), .Z(n5756) );
  AND U6064 ( .A(n5757), .B(n5756), .Z(n5858) );
  AND U6065 ( .A(x[64]), .B(y[254]), .Z(n5974) );
  AND U6066 ( .A(x[93]), .B(y[225]), .Z(n5952) );
  XOR U6067 ( .A(o[62]), .B(n5952), .Z(n5976) );
  AND U6068 ( .A(x[94]), .B(y[224]), .Z(n5975) );
  XOR U6069 ( .A(n5976), .B(n5975), .Z(n5973) );
  XOR U6070 ( .A(n5974), .B(n5973), .Z(n5860) );
  AND U6071 ( .A(x[84]), .B(y[234]), .Z(n5999) );
  XOR U6072 ( .A(n6000), .B(n5999), .Z(n5998) );
  AND U6073 ( .A(x[72]), .B(y[246]), .Z(n5997) );
  XNOR U6074 ( .A(n5998), .B(n5997), .Z(n5859) );
  XNOR U6075 ( .A(n5858), .B(n5857), .Z(n6059) );
  AND U6076 ( .A(x[71]), .B(y[247]), .Z(n5878) );
  NAND U6077 ( .A(n5758), .B(n5878), .Z(n5762) );
  NAND U6078 ( .A(n5760), .B(n5759), .Z(n5761) );
  AND U6079 ( .A(n5762), .B(n5761), .Z(n5852) );
  AND U6080 ( .A(y[233]), .B(x[85]), .Z(n5764) );
  NAND U6081 ( .A(y[232]), .B(x[86]), .Z(n5763) );
  XNOR U6082 ( .A(n5764), .B(n5763), .Z(n5877) );
  XOR U6083 ( .A(n5878), .B(n5877), .Z(n5854) );
  AND U6084 ( .A(x[81]), .B(y[237]), .Z(n5915) );
  AND U6085 ( .A(x[66]), .B(y[252]), .Z(n5917) );
  AND U6086 ( .A(x[90]), .B(y[228]), .Z(n5916) );
  XOR U6087 ( .A(n5917), .B(n5916), .Z(n5914) );
  XNOR U6088 ( .A(n5915), .B(n5914), .Z(n5853) );
  XOR U6089 ( .A(n5852), .B(n5851), .Z(n6058) );
  XNOR U6090 ( .A(n6057), .B(n6058), .Z(n6071) );
  NAND U6091 ( .A(n5766), .B(n5765), .Z(n5770) );
  NAND U6092 ( .A(n5768), .B(n5767), .Z(n5769) );
  AND U6093 ( .A(n5770), .B(n5769), .Z(n6072) );
  XOR U6094 ( .A(n6070), .B(n6069), .Z(n6094) );
  XNOR U6095 ( .A(n6093), .B(n6094), .Z(n6092) );
  NAND U6096 ( .A(n5772), .B(n5771), .Z(n5776) );
  NAND U6097 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U6098 ( .A(n5776), .B(n5775), .Z(n6099) );
  XOR U6099 ( .A(n6102), .B(n6099), .Z(n5777) );
  XOR U6100 ( .A(n6100), .B(n5777), .Z(n6086) );
  NANDN U6101 ( .A(n5779), .B(n5778), .Z(n5783) );
  NANDN U6102 ( .A(n5781), .B(n5780), .Z(n5782) );
  AND U6103 ( .A(n5783), .B(n5782), .Z(n6088) );
  NANDN U6104 ( .A(n5785), .B(n5784), .Z(n5789) );
  NANDN U6105 ( .A(n5787), .B(n5786), .Z(n5788) );
  AND U6106 ( .A(n5789), .B(n5788), .Z(n5834) );
  NAND U6107 ( .A(n5791), .B(n5790), .Z(n5795) );
  NAND U6108 ( .A(n5793), .B(n5792), .Z(n5794) );
  AND U6109 ( .A(n5795), .B(n5794), .Z(n6053) );
  NAND U6110 ( .A(n5797), .B(n5796), .Z(n5801) );
  NANDN U6111 ( .A(n5799), .B(n5798), .Z(n5800) );
  NAND U6112 ( .A(n5801), .B(n5800), .Z(n6054) );
  XNOR U6113 ( .A(n6053), .B(n6054), .Z(n6052) );
  NANDN U6114 ( .A(n5803), .B(n5802), .Z(n5807) );
  NANDN U6115 ( .A(n5805), .B(n5804), .Z(n5806) );
  NAND U6116 ( .A(n5807), .B(n5806), .Z(n6051) );
  XOR U6117 ( .A(n6052), .B(n6051), .Z(n5836) );
  NAND U6118 ( .A(n5808), .B(n5970), .Z(n5812) );
  NAND U6119 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6120 ( .A(n5812), .B(n5811), .Z(n5841) );
  NAND U6121 ( .A(n5814), .B(n5813), .Z(n5818) );
  NAND U6122 ( .A(n5816), .B(n5815), .Z(n5817) );
  NAND U6123 ( .A(n5818), .B(n5817), .Z(n5865) );
  AND U6124 ( .A(y[242]), .B(x[76]), .Z(n5819) );
  XOR U6125 ( .A(n5820), .B(n5819), .Z(n6017) );
  XOR U6126 ( .A(n6018), .B(n6017), .Z(n5968) );
  AND U6127 ( .A(y[245]), .B(x[73]), .Z(n5821) );
  XOR U6128 ( .A(n5822), .B(n5821), .Z(n5967) );
  XOR U6129 ( .A(n5968), .B(n5967), .Z(n5868) );
  AND U6130 ( .A(x[91]), .B(y[227]), .Z(n6014) );
  AND U6131 ( .A(x[65]), .B(y[253]), .Z(n6013) );
  XOR U6132 ( .A(n6014), .B(n6013), .Z(n6011) );
  XOR U6133 ( .A(n6012), .B(n6011), .Z(n5867) );
  XOR U6134 ( .A(n5868), .B(n5867), .Z(n5866) );
  XOR U6135 ( .A(n5865), .B(n5866), .Z(n5842) );
  NAND U6136 ( .A(n5824), .B(n5823), .Z(n5828) );
  NANDN U6137 ( .A(n5826), .B(n5825), .Z(n5827) );
  AND U6138 ( .A(n5828), .B(n5827), .Z(n5839) );
  XNOR U6139 ( .A(n5840), .B(n5839), .Z(n5835) );
  XOR U6140 ( .A(n5834), .B(n5833), .Z(n6087) );
  XOR U6141 ( .A(n6086), .B(n6085), .Z(n6106) );
  XOR U6142 ( .A(n6105), .B(n6106), .Z(n6107) );
  XOR U6143 ( .A(n6108), .B(n6107), .Z(n6111) );
  XNOR U6144 ( .A(n6112), .B(n6111), .Z(N127) );
  NANDN U6145 ( .A(n5836), .B(n5835), .Z(n5837) );
  NAND U6146 ( .A(n5840), .B(n5839), .Z(n5844) );
  NANDN U6147 ( .A(n5842), .B(n5841), .Z(n5843) );
  AND U6148 ( .A(n5844), .B(n5843), .Z(n6068) );
  NAND U6149 ( .A(n5846), .B(n5845), .Z(n5850) );
  NANDN U6150 ( .A(n5848), .B(n5847), .Z(n5849) );
  AND U6151 ( .A(n5850), .B(n5849), .Z(n6050) );
  NAND U6152 ( .A(n5852), .B(n5851), .Z(n5856) );
  NANDN U6153 ( .A(n5854), .B(n5853), .Z(n5855) );
  AND U6154 ( .A(n5856), .B(n5855), .Z(n5864) );
  NAND U6155 ( .A(n5858), .B(n5857), .Z(n5862) );
  NANDN U6156 ( .A(n5860), .B(n5859), .Z(n5861) );
  NAND U6157 ( .A(n5862), .B(n5861), .Z(n5863) );
  XNOR U6158 ( .A(n5864), .B(n5863), .Z(n6048) );
  NAND U6159 ( .A(n5866), .B(n5865), .Z(n5870) );
  NAND U6160 ( .A(n5868), .B(n5867), .Z(n5869) );
  AND U6161 ( .A(n5870), .B(n5869), .Z(n6046) );
  NAND U6162 ( .A(n5872), .B(n5871), .Z(n5876) );
  NAND U6163 ( .A(n5874), .B(n5873), .Z(n5875) );
  AND U6164 ( .A(n5876), .B(n5875), .Z(n5907) );
  NAND U6165 ( .A(n5878), .B(n5877), .Z(n5881) );
  AND U6166 ( .A(x[86]), .B(y[233]), .Z(n5933) );
  NAND U6167 ( .A(n5879), .B(n5933), .Z(n5880) );
  AND U6168 ( .A(n5881), .B(n5880), .Z(n5889) );
  NAND U6169 ( .A(n5883), .B(n5882), .Z(n5887) );
  NANDN U6170 ( .A(n5885), .B(n5884), .Z(n5886) );
  NAND U6171 ( .A(n5887), .B(n5886), .Z(n5888) );
  XNOR U6172 ( .A(n5889), .B(n5888), .Z(n5905) );
  AND U6173 ( .A(y[237]), .B(x[82]), .Z(n5891) );
  NAND U6174 ( .A(y[252]), .B(x[67]), .Z(n5890) );
  XNOR U6175 ( .A(n5891), .B(n5890), .Z(n5895) );
  AND U6176 ( .A(y[247]), .B(x[72]), .Z(n5893) );
  NAND U6177 ( .A(y[253]), .B(x[66]), .Z(n5892) );
  XNOR U6178 ( .A(n5893), .B(n5892), .Z(n5894) );
  XOR U6179 ( .A(n5895), .B(n5894), .Z(n5903) );
  AND U6180 ( .A(y[224]), .B(x[95]), .Z(n5897) );
  NAND U6181 ( .A(y[251]), .B(x[68]), .Z(n5896) );
  XNOR U6182 ( .A(n5897), .B(n5896), .Z(n5901) );
  AND U6183 ( .A(y[248]), .B(x[71]), .Z(n5899) );
  NAND U6184 ( .A(y[250]), .B(x[69]), .Z(n5898) );
  XNOR U6185 ( .A(n5899), .B(n5898), .Z(n5900) );
  XNOR U6186 ( .A(n5901), .B(n5900), .Z(n5902) );
  XNOR U6187 ( .A(n5903), .B(n5902), .Z(n5904) );
  XNOR U6188 ( .A(n5905), .B(n5904), .Z(n5906) );
  XNOR U6189 ( .A(n5907), .B(n5906), .Z(n5996) );
  NANDN U6190 ( .A(n5909), .B(n5908), .Z(n5913) );
  NANDN U6191 ( .A(n5911), .B(n5910), .Z(n5912) );
  AND U6192 ( .A(n5913), .B(n5912), .Z(n5994) );
  NAND U6193 ( .A(n5915), .B(n5914), .Z(n5919) );
  NAND U6194 ( .A(n5917), .B(n5916), .Z(n5918) );
  AND U6195 ( .A(n5919), .B(n5918), .Z(n5926) );
  NAND U6196 ( .A(n5921), .B(n5920), .Z(n5924) );
  NAND U6197 ( .A(n5954), .B(n5922), .Z(n5923) );
  NAND U6198 ( .A(n5924), .B(n5923), .Z(n5925) );
  XNOR U6199 ( .A(n5926), .B(n5925), .Z(n5992) );
  AND U6200 ( .A(y[227]), .B(x[92]), .Z(n5928) );
  NAND U6201 ( .A(y[243]), .B(x[76]), .Z(n5927) );
  XNOR U6202 ( .A(n5928), .B(n5927), .Z(n5932) );
  AND U6203 ( .A(y[255]), .B(x[64]), .Z(n5930) );
  NAND U6204 ( .A(y[254]), .B(x[65]), .Z(n5929) );
  XNOR U6205 ( .A(n5930), .B(n5929), .Z(n5931) );
  XOR U6206 ( .A(n5932), .B(n5931), .Z(n5935) );
  AND U6207 ( .A(x[74]), .B(y[245]), .Z(n5969) );
  XNOR U6208 ( .A(n5933), .B(n5969), .Z(n5934) );
  XNOR U6209 ( .A(n5935), .B(n5934), .Z(n5951) );
  AND U6210 ( .A(y[226]), .B(x[93]), .Z(n5937) );
  NAND U6211 ( .A(y[235]), .B(x[84]), .Z(n5936) );
  XNOR U6212 ( .A(n5937), .B(n5936), .Z(n5941) );
  AND U6213 ( .A(y[225]), .B(x[94]), .Z(n5939) );
  NAND U6214 ( .A(y[236]), .B(x[83]), .Z(n5938) );
  XNOR U6215 ( .A(n5939), .B(n5938), .Z(n5940) );
  XOR U6216 ( .A(n5941), .B(n5940), .Z(n5949) );
  AND U6217 ( .A(y[246]), .B(x[73]), .Z(n5943) );
  NAND U6218 ( .A(y[230]), .B(x[89]), .Z(n5942) );
  XNOR U6219 ( .A(n5943), .B(n5942), .Z(n5947) );
  AND U6220 ( .A(y[241]), .B(x[78]), .Z(n5945) );
  NAND U6221 ( .A(y[239]), .B(x[80]), .Z(n5944) );
  XNOR U6222 ( .A(n5945), .B(n5944), .Z(n5946) );
  XNOR U6223 ( .A(n5947), .B(n5946), .Z(n5948) );
  XNOR U6224 ( .A(n5949), .B(n5948), .Z(n5950) );
  XOR U6225 ( .A(n5951), .B(n5950), .Z(n5966) );
  AND U6226 ( .A(y[232]), .B(x[87]), .Z(n5960) );
  AND U6227 ( .A(n5952), .B(o[62]), .Z(n5958) );
  XOR U6228 ( .A(n6020), .B(o[63]), .Z(n5956) );
  XNOR U6229 ( .A(n5954), .B(n5953), .Z(n5955) );
  XNOR U6230 ( .A(n5956), .B(n5955), .Z(n5957) );
  XNOR U6231 ( .A(n5958), .B(n5957), .Z(n5959) );
  XNOR U6232 ( .A(n5960), .B(n5959), .Z(n5964) );
  AND U6233 ( .A(y[244]), .B(x[75]), .Z(n5962) );
  NAND U6234 ( .A(y[229]), .B(x[90]), .Z(n5961) );
  XNOR U6235 ( .A(n5962), .B(n5961), .Z(n5963) );
  XNOR U6236 ( .A(n5964), .B(n5963), .Z(n5965) );
  XNOR U6237 ( .A(n5966), .B(n5965), .Z(n5982) );
  NAND U6238 ( .A(n5968), .B(n5967), .Z(n5972) );
  NAND U6239 ( .A(n5970), .B(n5969), .Z(n5971) );
  AND U6240 ( .A(n5972), .B(n5971), .Z(n5980) );
  NAND U6241 ( .A(n5974), .B(n5973), .Z(n5978) );
  NAND U6242 ( .A(n5976), .B(n5975), .Z(n5977) );
  NAND U6243 ( .A(n5978), .B(n5977), .Z(n5979) );
  XNOR U6244 ( .A(n5980), .B(n5979), .Z(n5981) );
  XOR U6245 ( .A(n5982), .B(n5981), .Z(n5990) );
  AND U6246 ( .A(y[228]), .B(x[91]), .Z(n5984) );
  NAND U6247 ( .A(y[238]), .B(x[81]), .Z(n5983) );
  XNOR U6248 ( .A(n5984), .B(n5983), .Z(n5988) );
  AND U6249 ( .A(y[234]), .B(x[85]), .Z(n5986) );
  NAND U6250 ( .A(y[249]), .B(x[70]), .Z(n5985) );
  XNOR U6251 ( .A(n5986), .B(n5985), .Z(n5987) );
  XNOR U6252 ( .A(n5988), .B(n5987), .Z(n5989) );
  XNOR U6253 ( .A(n5990), .B(n5989), .Z(n5991) );
  XNOR U6254 ( .A(n5992), .B(n5991), .Z(n5993) );
  XNOR U6255 ( .A(n5994), .B(n5993), .Z(n5995) );
  XOR U6256 ( .A(n5996), .B(n5995), .Z(n6028) );
  NAND U6257 ( .A(n5998), .B(n5997), .Z(n6002) );
  NAND U6258 ( .A(n6000), .B(n5999), .Z(n6001) );
  AND U6259 ( .A(n6002), .B(n6001), .Z(n6010) );
  NAND U6260 ( .A(n6004), .B(n6003), .Z(n6008) );
  NANDN U6261 ( .A(n6006), .B(n6005), .Z(n6007) );
  NAND U6262 ( .A(n6008), .B(n6007), .Z(n6009) );
  XNOR U6263 ( .A(n6010), .B(n6009), .Z(n6026) );
  NAND U6264 ( .A(n6012), .B(n6011), .Z(n6016) );
  NAND U6265 ( .A(n6014), .B(n6013), .Z(n6015) );
  AND U6266 ( .A(n6016), .B(n6015), .Z(n6024) );
  NAND U6267 ( .A(n6018), .B(n6017), .Z(n6022) );
  NAND U6268 ( .A(n6020), .B(n6019), .Z(n6021) );
  NAND U6269 ( .A(n6022), .B(n6021), .Z(n6023) );
  XNOR U6270 ( .A(n6024), .B(n6023), .Z(n6025) );
  XNOR U6271 ( .A(n6026), .B(n6025), .Z(n6027) );
  XNOR U6272 ( .A(n6028), .B(n6027), .Z(n6044) );
  NANDN U6273 ( .A(n6030), .B(n6029), .Z(n6034) );
  NANDN U6274 ( .A(n6032), .B(n6031), .Z(n6033) );
  AND U6275 ( .A(n6034), .B(n6033), .Z(n6042) );
  NANDN U6276 ( .A(n6036), .B(n6035), .Z(n6040) );
  NANDN U6277 ( .A(n6038), .B(n6037), .Z(n6039) );
  NAND U6278 ( .A(n6040), .B(n6039), .Z(n6041) );
  XNOR U6279 ( .A(n6042), .B(n6041), .Z(n6043) );
  XNOR U6280 ( .A(n6044), .B(n6043), .Z(n6045) );
  XNOR U6281 ( .A(n6046), .B(n6045), .Z(n6047) );
  XNOR U6282 ( .A(n6048), .B(n6047), .Z(n6049) );
  XNOR U6283 ( .A(n6050), .B(n6049), .Z(n6066) );
  NAND U6284 ( .A(n6052), .B(n6051), .Z(n6056) );
  NANDN U6285 ( .A(n6054), .B(n6053), .Z(n6055) );
  AND U6286 ( .A(n6056), .B(n6055), .Z(n6064) );
  NANDN U6287 ( .A(n6058), .B(n6057), .Z(n6062) );
  NANDN U6288 ( .A(n6060), .B(n6059), .Z(n6061) );
  NAND U6289 ( .A(n6062), .B(n6061), .Z(n6063) );
  XNOR U6290 ( .A(n6064), .B(n6063), .Z(n6065) );
  XNOR U6291 ( .A(n6066), .B(n6065), .Z(n6067) );
  XNOR U6292 ( .A(n6068), .B(n6067), .Z(n6084) );
  NAND U6293 ( .A(n6070), .B(n6069), .Z(n6074) );
  NANDN U6294 ( .A(n6072), .B(n6071), .Z(n6073) );
  AND U6295 ( .A(n6074), .B(n6073), .Z(n6082) );
  NANDN U6296 ( .A(n6076), .B(n6075), .Z(n6080) );
  NAND U6297 ( .A(n6078), .B(n6077), .Z(n6079) );
  NAND U6298 ( .A(n6080), .B(n6079), .Z(n6081) );
  XNOR U6299 ( .A(n6082), .B(n6081), .Z(n6083) );
  NAND U6300 ( .A(n6086), .B(n6085), .Z(n6090) );
  NANDN U6301 ( .A(n6088), .B(n6087), .Z(n6089) );
  AND U6302 ( .A(n6090), .B(n6089), .Z(n6098) );
  NANDN U6303 ( .A(n6092), .B(n6091), .Z(n6096) );
  NAND U6304 ( .A(n6094), .B(n6093), .Z(n6095) );
  NAND U6305 ( .A(n6096), .B(n6095), .Z(n6097) );
  OR U6306 ( .A(n6099), .B(n6100), .Z(n6104) );
  AND U6307 ( .A(n6100), .B(n6099), .Z(n6101) );
  OR U6308 ( .A(n6102), .B(n6101), .Z(n6103) );
  AND U6309 ( .A(x[64]), .B(y[256]), .Z(n6771) );
  XOR U6310 ( .A(n6771), .B(o[64]), .Z(N161) );
  NAND U6311 ( .A(x[65]), .B(y[256]), .Z(n6116) );
  AND U6312 ( .A(x[64]), .B(y[257]), .Z(n6115) );
  XNOR U6313 ( .A(n6115), .B(o[65]), .Z(n6117) );
  XOR U6314 ( .A(n6116), .B(n6117), .Z(n6119) );
  NAND U6315 ( .A(n6771), .B(o[64]), .Z(n6118) );
  XNOR U6316 ( .A(n6119), .B(n6118), .Z(N162) );
  AND U6317 ( .A(y[256]), .B(x[66]), .Z(n6114) );
  NAND U6318 ( .A(y[257]), .B(x[65]), .Z(n6113) );
  XNOR U6319 ( .A(n6114), .B(n6113), .Z(n6131) );
  AND U6320 ( .A(n6115), .B(o[65]), .Z(n6130) );
  XNOR U6321 ( .A(n6131), .B(n6130), .Z(n6128) );
  AND U6322 ( .A(x[64]), .B(y[258]), .Z(n6125) );
  XOR U6323 ( .A(n6125), .B(o[66]), .Z(n6126) );
  IV U6324 ( .A(n6116), .Z(n6129) );
  NANDN U6325 ( .A(n6129), .B(n6117), .Z(n6121) );
  NAND U6326 ( .A(n6119), .B(n6118), .Z(n6120) );
  AND U6327 ( .A(n6121), .B(n6120), .Z(n6127) );
  XOR U6328 ( .A(n6126), .B(n6127), .Z(n6122) );
  XNOR U6329 ( .A(n6128), .B(n6122), .Z(N163) );
  AND U6330 ( .A(x[65]), .B(y[258]), .Z(n6258) );
  NAND U6331 ( .A(x[66]), .B(y[257]), .Z(n6142) );
  XOR U6332 ( .A(n6258), .B(n6151), .Z(n6153) );
  AND U6333 ( .A(y[256]), .B(x[67]), .Z(n6124) );
  NAND U6334 ( .A(y[259]), .B(x[64]), .Z(n6123) );
  XNOR U6335 ( .A(n6124), .B(n6123), .Z(n6136) );
  NAND U6336 ( .A(n6125), .B(o[66]), .Z(n6137) );
  XNOR U6337 ( .A(n6153), .B(n6152), .Z(n6147) );
  NANDN U6338 ( .A(n6142), .B(n6129), .Z(n6133) );
  NAND U6339 ( .A(n6131), .B(n6130), .Z(n6132) );
  NAND U6340 ( .A(n6133), .B(n6132), .Z(n6145) );
  IV U6341 ( .A(n6145), .Z(n6144) );
  XOR U6342 ( .A(n6146), .B(n6144), .Z(n6134) );
  XNOR U6343 ( .A(n6147), .B(n6134), .Z(N164) );
  AND U6344 ( .A(x[67]), .B(y[259]), .Z(n6135) );
  NAND U6345 ( .A(n6771), .B(n6135), .Z(n6139) );
  NANDN U6346 ( .A(n6137), .B(n6136), .Z(n6138) );
  AND U6347 ( .A(n6139), .B(n6138), .Z(n6181) );
  AND U6348 ( .A(y[260]), .B(x[64]), .Z(n6141) );
  NAND U6349 ( .A(y[256]), .B(x[68]), .Z(n6140) );
  XNOR U6350 ( .A(n6141), .B(n6140), .Z(n6168) );
  ANDN U6351 ( .B(o[67]), .A(n6142), .Z(n6167) );
  XOR U6352 ( .A(n6168), .B(n6167), .Z(n6179) );
  AND U6353 ( .A(y[258]), .B(x[66]), .Z(n6314) );
  NAND U6354 ( .A(y[259]), .B(x[65]), .Z(n6143) );
  XNOR U6355 ( .A(n6314), .B(n6143), .Z(n6164) );
  NAND U6356 ( .A(x[67]), .B(y[257]), .Z(n6161) );
  XNOR U6357 ( .A(o[68]), .B(n6161), .Z(n6163) );
  XOR U6358 ( .A(n6164), .B(n6163), .Z(n6178) );
  XOR U6359 ( .A(n6179), .B(n6178), .Z(n6180) );
  XOR U6360 ( .A(n6181), .B(n6180), .Z(n6174) );
  OR U6361 ( .A(n6146), .B(n6144), .Z(n6150) );
  ANDN U6362 ( .B(n6146), .A(n6145), .Z(n6148) );
  OR U6363 ( .A(n6148), .B(n6147), .Z(n6149) );
  AND U6364 ( .A(n6150), .B(n6149), .Z(n6173) );
  NAND U6365 ( .A(n6258), .B(n6151), .Z(n6155) );
  NAND U6366 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6367 ( .A(n6155), .B(n6154), .Z(n6172) );
  IV U6368 ( .A(n6172), .Z(n6171) );
  XOR U6369 ( .A(n6173), .B(n6171), .Z(n6156) );
  XNOR U6370 ( .A(n6174), .B(n6156), .Z(N165) );
  AND U6371 ( .A(y[258]), .B(x[67]), .Z(n6158) );
  NAND U6372 ( .A(y[260]), .B(x[65]), .Z(n6157) );
  XNOR U6373 ( .A(n6158), .B(n6157), .Z(n6186) );
  AND U6374 ( .A(x[68]), .B(y[257]), .Z(n6197) );
  XOR U6375 ( .A(n6197), .B(o[69]), .Z(n6185) );
  XNOR U6376 ( .A(n6186), .B(n6185), .Z(n6189) );
  NAND U6377 ( .A(x[66]), .B(y[259]), .Z(n6267) );
  AND U6378 ( .A(y[261]), .B(x[64]), .Z(n6160) );
  NAND U6379 ( .A(y[256]), .B(x[69]), .Z(n6159) );
  XNOR U6380 ( .A(n6160), .B(n6159), .Z(n6192) );
  ANDN U6381 ( .B(o[68]), .A(n6161), .Z(n6191) );
  XOR U6382 ( .A(n6192), .B(n6191), .Z(n6190) );
  XOR U6383 ( .A(n6267), .B(n6190), .Z(n6162) );
  XOR U6384 ( .A(n6189), .B(n6162), .Z(n6210) );
  NANDN U6385 ( .A(n6267), .B(n6258), .Z(n6166) );
  NAND U6386 ( .A(n6164), .B(n6163), .Z(n6165) );
  AND U6387 ( .A(n6166), .B(n6165), .Z(n6208) );
  AND U6388 ( .A(x[68]), .B(y[260]), .Z(n6979) );
  NAND U6389 ( .A(n6979), .B(n6771), .Z(n6170) );
  NAND U6390 ( .A(n6168), .B(n6167), .Z(n6169) );
  NAND U6391 ( .A(n6170), .B(n6169), .Z(n6207) );
  XNOR U6392 ( .A(n6210), .B(n6209), .Z(n6204) );
  OR U6393 ( .A(n6173), .B(n6171), .Z(n6177) );
  ANDN U6394 ( .B(n6173), .A(n6172), .Z(n6175) );
  OR U6395 ( .A(n6175), .B(n6174), .Z(n6176) );
  AND U6396 ( .A(n6177), .B(n6176), .Z(n6202) );
  NAND U6397 ( .A(n6179), .B(n6178), .Z(n6183) );
  NANDN U6398 ( .A(n6181), .B(n6180), .Z(n6182) );
  NAND U6399 ( .A(n6183), .B(n6182), .Z(n6201) );
  IV U6400 ( .A(n6201), .Z(n6200) );
  XOR U6401 ( .A(n6202), .B(n6200), .Z(n6184) );
  XNOR U6402 ( .A(n6204), .B(n6184), .Z(N166) );
  AND U6403 ( .A(x[67]), .B(y[260]), .Z(n6269) );
  NAND U6404 ( .A(n6258), .B(n6269), .Z(n6188) );
  NAND U6405 ( .A(n6186), .B(n6185), .Z(n6187) );
  AND U6406 ( .A(n6188), .B(n6187), .Z(n6246) );
  XNOR U6407 ( .A(n6246), .B(n6245), .Z(n6248) );
  AND U6408 ( .A(x[69]), .B(y[261]), .Z(n6433) );
  NAND U6409 ( .A(n6771), .B(n6433), .Z(n6194) );
  NAND U6410 ( .A(n6192), .B(n6191), .Z(n6193) );
  AND U6411 ( .A(n6194), .B(n6193), .Z(n6215) );
  AND U6412 ( .A(y[256]), .B(x[70]), .Z(n6196) );
  NAND U6413 ( .A(y[262]), .B(x[64]), .Z(n6195) );
  XNOR U6414 ( .A(n6196), .B(n6195), .Z(n6221) );
  NAND U6415 ( .A(n6197), .B(o[69]), .Z(n6222) );
  XNOR U6416 ( .A(n6221), .B(n6222), .Z(n6214) );
  AND U6417 ( .A(y[260]), .B(x[66]), .Z(n6711) );
  NAND U6418 ( .A(y[259]), .B(x[67]), .Z(n6198) );
  XNOR U6419 ( .A(n6711), .B(n6198), .Z(n6226) );
  AND U6420 ( .A(x[65]), .B(y[261]), .Z(n6493) );
  NAND U6421 ( .A(y[258]), .B(x[68]), .Z(n6199) );
  XNOR U6422 ( .A(n6493), .B(n6199), .Z(n6230) );
  NAND U6423 ( .A(x[69]), .B(y[257]), .Z(n6235) );
  XNOR U6424 ( .A(o[70]), .B(n6235), .Z(n6229) );
  XOR U6425 ( .A(n6230), .B(n6229), .Z(n6225) );
  XOR U6426 ( .A(n6226), .B(n6225), .Z(n6216) );
  XOR U6427 ( .A(n6217), .B(n6216), .Z(n6247) );
  XNOR U6428 ( .A(n6248), .B(n6247), .Z(n6241) );
  OR U6429 ( .A(n6202), .B(n6200), .Z(n6206) );
  ANDN U6430 ( .B(n6202), .A(n6201), .Z(n6203) );
  OR U6431 ( .A(n6204), .B(n6203), .Z(n6205) );
  AND U6432 ( .A(n6206), .B(n6205), .Z(n6240) );
  NANDN U6433 ( .A(n6208), .B(n6207), .Z(n6212) );
  NAND U6434 ( .A(n6210), .B(n6209), .Z(n6211) );
  NAND U6435 ( .A(n6212), .B(n6211), .Z(n6239) );
  IV U6436 ( .A(n6239), .Z(n6238) );
  XOR U6437 ( .A(n6240), .B(n6238), .Z(n6213) );
  XNOR U6438 ( .A(n6241), .B(n6213), .Z(N167) );
  NANDN U6439 ( .A(n6215), .B(n6214), .Z(n6219) );
  NAND U6440 ( .A(n6217), .B(n6216), .Z(n6218) );
  AND U6441 ( .A(n6219), .B(n6218), .Z(n6287) );
  AND U6442 ( .A(y[262]), .B(x[65]), .Z(n6626) );
  NAND U6443 ( .A(y[258]), .B(x[69]), .Z(n6220) );
  XNOR U6444 ( .A(n6626), .B(n6220), .Z(n6261) );
  NAND U6445 ( .A(x[70]), .B(y[257]), .Z(n6265) );
  XNOR U6446 ( .A(o[71]), .B(n6265), .Z(n6260) );
  XOR U6447 ( .A(n6261), .B(n6260), .Z(n6279) );
  AND U6448 ( .A(x[70]), .B(y[262]), .Z(n6513) );
  NAND U6449 ( .A(n6771), .B(n6513), .Z(n6224) );
  NANDN U6450 ( .A(n6222), .B(n6221), .Z(n6223) );
  AND U6451 ( .A(n6224), .B(n6223), .Z(n6278) );
  XNOR U6452 ( .A(n6279), .B(n6278), .Z(n6280) );
  NANDN U6453 ( .A(n6267), .B(n6269), .Z(n6228) );
  NAND U6454 ( .A(n6226), .B(n6225), .Z(n6227) );
  NAND U6455 ( .A(n6228), .B(n6227), .Z(n6281) );
  XNOR U6456 ( .A(n6280), .B(n6281), .Z(n6285) );
  AND U6457 ( .A(x[68]), .B(y[261]), .Z(n6776) );
  NAND U6458 ( .A(n6776), .B(n6258), .Z(n6232) );
  NAND U6459 ( .A(n6230), .B(n6229), .Z(n6231) );
  AND U6460 ( .A(n6232), .B(n6231), .Z(n6255) );
  AND U6461 ( .A(y[261]), .B(x[66]), .Z(n6234) );
  NAND U6462 ( .A(y[259]), .B(x[68]), .Z(n6233) );
  XNOR U6463 ( .A(n6234), .B(n6233), .Z(n6268) );
  XOR U6464 ( .A(n6269), .B(n6268), .Z(n6253) );
  ANDN U6465 ( .B(o[70]), .A(n6235), .Z(n6273) );
  AND U6466 ( .A(y[256]), .B(x[71]), .Z(n6237) );
  NAND U6467 ( .A(y[263]), .B(x[64]), .Z(n6236) );
  XNOR U6468 ( .A(n6237), .B(n6236), .Z(n6272) );
  XNOR U6469 ( .A(n6273), .B(n6272), .Z(n6252) );
  XNOR U6470 ( .A(n6253), .B(n6252), .Z(n6254) );
  XOR U6471 ( .A(n6255), .B(n6254), .Z(n6284) );
  XOR U6472 ( .A(n6285), .B(n6284), .Z(n6286) );
  XNOR U6473 ( .A(n6287), .B(n6286), .Z(n6293) );
  OR U6474 ( .A(n6240), .B(n6238), .Z(n6244) );
  ANDN U6475 ( .B(n6240), .A(n6239), .Z(n6242) );
  OR U6476 ( .A(n6242), .B(n6241), .Z(n6243) );
  AND U6477 ( .A(n6244), .B(n6243), .Z(n6291) );
  NANDN U6478 ( .A(n6246), .B(n6245), .Z(n6250) );
  NAND U6479 ( .A(n6248), .B(n6247), .Z(n6249) );
  AND U6480 ( .A(n6250), .B(n6249), .Z(n6292) );
  IV U6481 ( .A(n6292), .Z(n6290) );
  XOR U6482 ( .A(n6291), .B(n6290), .Z(n6251) );
  XNOR U6483 ( .A(n6293), .B(n6251), .Z(N168) );
  NANDN U6484 ( .A(n6253), .B(n6252), .Z(n6257) );
  NAND U6485 ( .A(n6255), .B(n6254), .Z(n6256) );
  AND U6486 ( .A(n6257), .B(n6256), .Z(n6327) );
  AND U6487 ( .A(x[69]), .B(y[262]), .Z(n6259) );
  NAND U6488 ( .A(n6259), .B(n6258), .Z(n6263) );
  NAND U6489 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U6490 ( .A(n6263), .B(n6262), .Z(n6325) );
  AND U6491 ( .A(y[263]), .B(x[65]), .Z(n6766) );
  NAND U6492 ( .A(y[259]), .B(x[69]), .Z(n6264) );
  XNOR U6493 ( .A(n6766), .B(n6264), .Z(n6308) );
  ANDN U6494 ( .B(o[71]), .A(n6265), .Z(n6307) );
  XOR U6495 ( .A(n6308), .B(n6307), .Z(n6313) );
  NAND U6496 ( .A(x[67]), .B(y[261]), .Z(n7117) );
  AND U6497 ( .A(y[262]), .B(x[66]), .Z(n7242) );
  NAND U6498 ( .A(y[258]), .B(x[70]), .Z(n6266) );
  XNOR U6499 ( .A(n7242), .B(n6266), .Z(n6315) );
  XNOR U6500 ( .A(n6979), .B(n6315), .Z(n6311) );
  XOR U6501 ( .A(n7117), .B(n6311), .Z(n6312) );
  XOR U6502 ( .A(n6313), .B(n6312), .Z(n6324) );
  XNOR U6503 ( .A(n6325), .B(n6324), .Z(n6326) );
  XOR U6504 ( .A(n6327), .B(n6326), .Z(n6336) );
  NANDN U6505 ( .A(n6267), .B(n6776), .Z(n6271) );
  NAND U6506 ( .A(n6269), .B(n6268), .Z(n6270) );
  AND U6507 ( .A(n6271), .B(n6270), .Z(n6321) );
  AND U6508 ( .A(x[71]), .B(y[263]), .Z(n6647) );
  NAND U6509 ( .A(n6771), .B(n6647), .Z(n6275) );
  NAND U6510 ( .A(n6273), .B(n6272), .Z(n6274) );
  AND U6511 ( .A(n6275), .B(n6274), .Z(n6319) );
  AND U6512 ( .A(y[256]), .B(x[72]), .Z(n6277) );
  NAND U6513 ( .A(y[264]), .B(x[64]), .Z(n6276) );
  XNOR U6514 ( .A(n6277), .B(n6276), .Z(n6299) );
  NAND U6515 ( .A(x[71]), .B(y[257]), .Z(n6303) );
  XNOR U6516 ( .A(o[72]), .B(n6303), .Z(n6298) );
  XOR U6517 ( .A(n6299), .B(n6298), .Z(n6318) );
  XNOR U6518 ( .A(n6319), .B(n6318), .Z(n6320) );
  XOR U6519 ( .A(n6321), .B(n6320), .Z(n6334) );
  NANDN U6520 ( .A(n6279), .B(n6278), .Z(n6283) );
  NANDN U6521 ( .A(n6281), .B(n6280), .Z(n6282) );
  NAND U6522 ( .A(n6283), .B(n6282), .Z(n6333) );
  XOR U6523 ( .A(n6334), .B(n6333), .Z(n6335) );
  XOR U6524 ( .A(n6336), .B(n6335), .Z(n6332) );
  NAND U6525 ( .A(n6285), .B(n6284), .Z(n6289) );
  NAND U6526 ( .A(n6287), .B(n6286), .Z(n6288) );
  NAND U6527 ( .A(n6289), .B(n6288), .Z(n6330) );
  NANDN U6528 ( .A(n6290), .B(n6291), .Z(n6296) );
  NOR U6529 ( .A(n6292), .B(n6291), .Z(n6294) );
  OR U6530 ( .A(n6294), .B(n6293), .Z(n6295) );
  AND U6531 ( .A(n6296), .B(n6295), .Z(n6331) );
  XOR U6532 ( .A(n6330), .B(n6331), .Z(n6297) );
  XNOR U6533 ( .A(n6332), .B(n6297), .Z(N169) );
  AND U6534 ( .A(x[72]), .B(y[264]), .Z(n6793) );
  NAND U6535 ( .A(n6793), .B(n6771), .Z(n6301) );
  NAND U6536 ( .A(n6299), .B(n6298), .Z(n6300) );
  AND U6537 ( .A(n6301), .B(n6300), .Z(n6375) );
  AND U6538 ( .A(y[258]), .B(x[71]), .Z(n6702) );
  NAND U6539 ( .A(y[260]), .B(x[69]), .Z(n6302) );
  XNOR U6540 ( .A(n6702), .B(n6302), .Z(n6349) );
  ANDN U6541 ( .B(o[72]), .A(n6303), .Z(n6348) );
  XOR U6542 ( .A(n6349), .B(n6348), .Z(n6373) );
  AND U6543 ( .A(y[256]), .B(x[73]), .Z(n6305) );
  NAND U6544 ( .A(y[265]), .B(x[64]), .Z(n6304) );
  XNOR U6545 ( .A(n6305), .B(n6304), .Z(n6355) );
  NAND U6546 ( .A(x[72]), .B(y[257]), .Z(n6362) );
  XNOR U6547 ( .A(n6355), .B(n6354), .Z(n6372) );
  XOR U6548 ( .A(n6375), .B(n6374), .Z(n6369) );
  AND U6549 ( .A(y[259]), .B(x[70]), .Z(n6715) );
  NAND U6550 ( .A(y[264]), .B(x[65]), .Z(n6306) );
  XNOR U6551 ( .A(n6715), .B(n6306), .Z(n6359) );
  XOR U6552 ( .A(n6776), .B(n6359), .Z(n6379) );
  NAND U6553 ( .A(x[66]), .B(y[263]), .Z(n7027) );
  NAND U6554 ( .A(x[67]), .B(y[262]), .Z(n6725) );
  XOR U6555 ( .A(n7027), .B(n6725), .Z(n6378) );
  NAND U6556 ( .A(x[69]), .B(y[263]), .Z(n6549) );
  AND U6557 ( .A(x[65]), .B(y[259]), .Z(n6358) );
  NANDN U6558 ( .A(n6549), .B(n6358), .Z(n6310) );
  NAND U6559 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U6560 ( .A(n6310), .B(n6309), .Z(n6366) );
  XOR U6561 ( .A(n6367), .B(n6366), .Z(n6368) );
  XOR U6562 ( .A(n6369), .B(n6368), .Z(n6342) );
  NAND U6563 ( .A(n6513), .B(n6314), .Z(n6317) );
  NAND U6564 ( .A(n6979), .B(n6315), .Z(n6316) );
  AND U6565 ( .A(n6317), .B(n6316), .Z(n6340) );
  XNOR U6566 ( .A(n6341), .B(n6340), .Z(n6343) );
  XNOR U6567 ( .A(n6342), .B(n6343), .Z(n6387) );
  NANDN U6568 ( .A(n6319), .B(n6318), .Z(n6323) );
  NANDN U6569 ( .A(n6321), .B(n6320), .Z(n6322) );
  AND U6570 ( .A(n6323), .B(n6322), .Z(n6386) );
  NANDN U6571 ( .A(n6325), .B(n6324), .Z(n6329) );
  NAND U6572 ( .A(n6327), .B(n6326), .Z(n6328) );
  NAND U6573 ( .A(n6329), .B(n6328), .Z(n6385) );
  XNOR U6574 ( .A(n6386), .B(n6385), .Z(n6388) );
  XNOR U6575 ( .A(n6387), .B(n6388), .Z(n6384) );
  NAND U6576 ( .A(n6334), .B(n6333), .Z(n6338) );
  NANDN U6577 ( .A(n6336), .B(n6335), .Z(n6337) );
  AND U6578 ( .A(n6338), .B(n6337), .Z(n6383) );
  XOR U6579 ( .A(n6382), .B(n6383), .Z(n6339) );
  XNOR U6580 ( .A(n6384), .B(n6339), .Z(N170) );
  NANDN U6581 ( .A(n6341), .B(n6340), .Z(n6345) );
  NAND U6582 ( .A(n6343), .B(n6342), .Z(n6344) );
  AND U6583 ( .A(n6345), .B(n6344), .Z(n6453) );
  AND U6584 ( .A(x[71]), .B(y[260]), .Z(n6347) );
  AND U6585 ( .A(x[69]), .B(y[258]), .Z(n6346) );
  NAND U6586 ( .A(n6347), .B(n6346), .Z(n6351) );
  NAND U6587 ( .A(n6349), .B(n6348), .Z(n6350) );
  AND U6588 ( .A(n6351), .B(n6350), .Z(n6440) );
  AND U6589 ( .A(y[259]), .B(x[71]), .Z(n6353) );
  NAND U6590 ( .A(y[262]), .B(x[68]), .Z(n6352) );
  XNOR U6591 ( .A(n6353), .B(n6352), .Z(n6412) );
  AND U6592 ( .A(x[70]), .B(y[260]), .Z(n6411) );
  XOR U6593 ( .A(n6412), .B(n6411), .Z(n6438) );
  AND U6594 ( .A(x[72]), .B(y[258]), .Z(n6622) );
  AND U6595 ( .A(x[73]), .B(y[257]), .Z(n6421) );
  XOR U6596 ( .A(n6421), .B(o[74]), .Z(n6432) );
  XOR U6597 ( .A(n6622), .B(n6432), .Z(n6434) );
  XNOR U6598 ( .A(n6434), .B(n6433), .Z(n6437) );
  XOR U6599 ( .A(n6440), .B(n6439), .Z(n6401) );
  AND U6600 ( .A(x[73]), .B(y[265]), .Z(n6988) );
  NAND U6601 ( .A(n6988), .B(n6771), .Z(n6357) );
  NAND U6602 ( .A(n6355), .B(n6354), .Z(n6356) );
  AND U6603 ( .A(n6357), .B(n6356), .Z(n6399) );
  AND U6604 ( .A(x[70]), .B(y[264]), .Z(n6657) );
  NAND U6605 ( .A(n6657), .B(n6358), .Z(n6361) );
  NAND U6606 ( .A(n6776), .B(n6359), .Z(n6360) );
  NAND U6607 ( .A(n6361), .B(n6360), .Z(n6406) );
  ANDN U6608 ( .B(o[73]), .A(n6362), .Z(n6416) );
  AND U6609 ( .A(x[74]), .B(y[256]), .Z(n6364) );
  AND U6610 ( .A(y[266]), .B(x[64]), .Z(n6363) );
  XOR U6611 ( .A(n6364), .B(n6363), .Z(n6415) );
  XOR U6612 ( .A(n6416), .B(n6415), .Z(n6405) );
  AND U6613 ( .A(y[263]), .B(x[67]), .Z(n7365) );
  NAND U6614 ( .A(y[265]), .B(x[65]), .Z(n6365) );
  XNOR U6615 ( .A(n7365), .B(n6365), .Z(n6429) );
  AND U6616 ( .A(x[66]), .B(y[264]), .Z(n6428) );
  XOR U6617 ( .A(n6429), .B(n6428), .Z(n6404) );
  XOR U6618 ( .A(n6405), .B(n6404), .Z(n6407) );
  XOR U6619 ( .A(n6406), .B(n6407), .Z(n6398) );
  NAND U6620 ( .A(n6367), .B(n6366), .Z(n6371) );
  NANDN U6621 ( .A(n6369), .B(n6368), .Z(n6370) );
  AND U6622 ( .A(n6371), .B(n6370), .Z(n6395) );
  NANDN U6623 ( .A(n6373), .B(n6372), .Z(n6377) );
  NAND U6624 ( .A(n6375), .B(n6374), .Z(n6376) );
  AND U6625 ( .A(n6377), .B(n6376), .Z(n6392) );
  AND U6626 ( .A(n7027), .B(n6725), .Z(n6381) );
  NANDN U6627 ( .A(n6379), .B(n6378), .Z(n6380) );
  NANDN U6628 ( .A(n6381), .B(n6380), .Z(n6393) );
  XOR U6629 ( .A(n6395), .B(n6394), .Z(n6450) );
  XOR U6630 ( .A(n6451), .B(n6450), .Z(n6452) );
  XOR U6631 ( .A(n6453), .B(n6452), .Z(n6446) );
  NANDN U6632 ( .A(n6386), .B(n6385), .Z(n6390) );
  NAND U6633 ( .A(n6388), .B(n6387), .Z(n6389) );
  AND U6634 ( .A(n6390), .B(n6389), .Z(n6445) );
  IV U6635 ( .A(n6445), .Z(n6443) );
  XOR U6636 ( .A(n6444), .B(n6443), .Z(n6391) );
  XNOR U6637 ( .A(n6446), .B(n6391), .Z(N171) );
  NANDN U6638 ( .A(n6393), .B(n6392), .Z(n6397) );
  NANDN U6639 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U6640 ( .A(n6397), .B(n6396), .Z(n6460) );
  NANDN U6641 ( .A(n6399), .B(n6398), .Z(n6403) );
  NANDN U6642 ( .A(n6401), .B(n6400), .Z(n6402) );
  AND U6643 ( .A(n6403), .B(n6402), .Z(n6458) );
  NAND U6644 ( .A(n6405), .B(n6404), .Z(n6409) );
  NAND U6645 ( .A(n6407), .B(n6406), .Z(n6408) );
  NAND U6646 ( .A(n6409), .B(n6408), .Z(n6479) );
  AND U6647 ( .A(x[71]), .B(y[262]), .Z(n6544) );
  AND U6648 ( .A(x[68]), .B(y[259]), .Z(n6410) );
  NAND U6649 ( .A(n6544), .B(n6410), .Z(n6414) );
  NAND U6650 ( .A(n6412), .B(n6411), .Z(n6413) );
  NAND U6651 ( .A(n6414), .B(n6413), .Z(n6477) );
  AND U6652 ( .A(x[74]), .B(y[266]), .Z(n7248) );
  NAND U6653 ( .A(n7248), .B(n6771), .Z(n6418) );
  NAND U6654 ( .A(n6416), .B(n6415), .Z(n6417) );
  NAND U6655 ( .A(n6418), .B(n6417), .Z(n6473) );
  AND U6656 ( .A(y[256]), .B(x[75]), .Z(n6420) );
  NAND U6657 ( .A(y[267]), .B(x[64]), .Z(n6419) );
  XNOR U6658 ( .A(n6420), .B(n6419), .Z(n6503) );
  NAND U6659 ( .A(n6421), .B(o[74]), .Z(n6504) );
  XNOR U6660 ( .A(n6503), .B(n6504), .Z(n6472) );
  AND U6661 ( .A(y[261]), .B(x[70]), .Z(n6423) );
  NAND U6662 ( .A(y[266]), .B(x[65]), .Z(n6422) );
  XNOR U6663 ( .A(n6423), .B(n6422), .Z(n6495) );
  NAND U6664 ( .A(x[74]), .B(y[257]), .Z(n6511) );
  XNOR U6665 ( .A(o[75]), .B(n6511), .Z(n6494) );
  XOR U6666 ( .A(n6495), .B(n6494), .Z(n6471) );
  XOR U6667 ( .A(n6472), .B(n6471), .Z(n6474) );
  XOR U6668 ( .A(n6473), .B(n6474), .Z(n6478) );
  XOR U6669 ( .A(n6477), .B(n6478), .Z(n6480) );
  XNOR U6670 ( .A(n6479), .B(n6480), .Z(n6516) );
  AND U6671 ( .A(x[67]), .B(y[264]), .Z(n7497) );
  AND U6672 ( .A(y[265]), .B(x[66]), .Z(n6425) );
  NAND U6673 ( .A(y[262]), .B(x[69]), .Z(n6424) );
  XNOR U6674 ( .A(n6425), .B(n6424), .Z(n6490) );
  AND U6675 ( .A(x[68]), .B(y[263]), .Z(n6489) );
  XNOR U6676 ( .A(n6490), .B(n6489), .Z(n6466) );
  XNOR U6677 ( .A(n7497), .B(n6466), .Z(n6467) );
  AND U6678 ( .A(y[258]), .B(x[73]), .Z(n6427) );
  NAND U6679 ( .A(y[260]), .B(x[71]), .Z(n6426) );
  XNOR U6680 ( .A(n6427), .B(n6426), .Z(n6507) );
  NAND U6681 ( .A(x[72]), .B(y[259]), .Z(n6508) );
  XNOR U6682 ( .A(n6507), .B(n6508), .Z(n6468) );
  NAND U6683 ( .A(x[67]), .B(y[265]), .Z(n6540) );
  NANDN U6684 ( .A(n6540), .B(n6766), .Z(n6431) );
  NAND U6685 ( .A(n6429), .B(n6428), .Z(n6430) );
  NAND U6686 ( .A(n6431), .B(n6430), .Z(n6484) );
  NAND U6687 ( .A(n6622), .B(n6432), .Z(n6436) );
  NAND U6688 ( .A(n6434), .B(n6433), .Z(n6435) );
  NAND U6689 ( .A(n6436), .B(n6435), .Z(n6483) );
  XOR U6690 ( .A(n6484), .B(n6483), .Z(n6485) );
  NANDN U6691 ( .A(n6438), .B(n6437), .Z(n6442) );
  NAND U6692 ( .A(n6440), .B(n6439), .Z(n6441) );
  NAND U6693 ( .A(n6442), .B(n6441), .Z(n6514) );
  XOR U6694 ( .A(n6516), .B(n6517), .Z(n6457) );
  XOR U6695 ( .A(n6460), .B(n6459), .Z(n6465) );
  NANDN U6696 ( .A(n6443), .B(n6444), .Z(n6449) );
  NOR U6697 ( .A(n6445), .B(n6444), .Z(n6447) );
  OR U6698 ( .A(n6447), .B(n6446), .Z(n6448) );
  AND U6699 ( .A(n6449), .B(n6448), .Z(n6463) );
  NAND U6700 ( .A(n6451), .B(n6450), .Z(n6455) );
  NANDN U6701 ( .A(n6453), .B(n6452), .Z(n6454) );
  AND U6702 ( .A(n6455), .B(n6454), .Z(n6464) );
  XOR U6703 ( .A(n6463), .B(n6464), .Z(n6456) );
  XNOR U6704 ( .A(n6465), .B(n6456), .Z(N172) );
  NANDN U6705 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6706 ( .A(n6460), .B(n6459), .Z(n6461) );
  NAND U6707 ( .A(n6462), .B(n6461), .Z(n6585) );
  IV U6708 ( .A(n6585), .Z(n6584) );
  NANDN U6709 ( .A(n7497), .B(n6466), .Z(n6470) );
  NANDN U6710 ( .A(n6468), .B(n6467), .Z(n6469) );
  NAND U6711 ( .A(n6470), .B(n6469), .Z(n6521) );
  NAND U6712 ( .A(n6472), .B(n6471), .Z(n6476) );
  NAND U6713 ( .A(n6474), .B(n6473), .Z(n6475) );
  AND U6714 ( .A(n6476), .B(n6475), .Z(n6522) );
  XOR U6715 ( .A(n6521), .B(n6522), .Z(n6524) );
  NAND U6716 ( .A(n6478), .B(n6477), .Z(n6482) );
  NAND U6717 ( .A(n6480), .B(n6479), .Z(n6481) );
  AND U6718 ( .A(n6482), .B(n6481), .Z(n6523) );
  XOR U6719 ( .A(n6524), .B(n6523), .Z(n6593) );
  NAND U6720 ( .A(n6484), .B(n6483), .Z(n6488) );
  NANDN U6721 ( .A(n6486), .B(n6485), .Z(n6487) );
  NAND U6722 ( .A(n6488), .B(n6487), .Z(n6580) );
  AND U6723 ( .A(x[69]), .B(y[265]), .Z(n7018) );
  NAND U6724 ( .A(n7242), .B(n7018), .Z(n6492) );
  NAND U6725 ( .A(n6490), .B(n6489), .Z(n6491) );
  AND U6726 ( .A(n6492), .B(n6491), .Z(n6528) );
  AND U6727 ( .A(x[70]), .B(y[266]), .Z(n6782) );
  NAND U6728 ( .A(n6782), .B(n6493), .Z(n6497) );
  NAND U6729 ( .A(n6495), .B(n6494), .Z(n6496) );
  NAND U6730 ( .A(n6497), .B(n6496), .Z(n6527) );
  AND U6731 ( .A(x[73]), .B(y[259]), .Z(n7237) );
  AND U6732 ( .A(y[258]), .B(x[74]), .Z(n7232) );
  NAND U6733 ( .A(y[264]), .B(x[68]), .Z(n6498) );
  XOR U6734 ( .A(n7232), .B(n6498), .Z(n6571) );
  XNOR U6735 ( .A(n7237), .B(n6571), .Z(n6550) );
  NAND U6736 ( .A(x[71]), .B(y[261]), .Z(n6548) );
  XOR U6737 ( .A(n6549), .B(n6548), .Z(n6551) );
  AND U6738 ( .A(y[256]), .B(x[76]), .Z(n6500) );
  NAND U6739 ( .A(y[268]), .B(x[64]), .Z(n6499) );
  XNOR U6740 ( .A(n6500), .B(n6499), .Z(n6565) );
  NAND U6741 ( .A(x[75]), .B(y[257]), .Z(n6545) );
  XNOR U6742 ( .A(o[76]), .B(n6545), .Z(n6564) );
  XOR U6743 ( .A(n6565), .B(n6564), .Z(n6534) );
  AND U6744 ( .A(y[260]), .B(x[72]), .Z(n6502) );
  NAND U6745 ( .A(y[266]), .B(x[66]), .Z(n6501) );
  XNOR U6746 ( .A(n6502), .B(n6501), .Z(n6539) );
  XNOR U6747 ( .A(n6539), .B(n6540), .Z(n6533) );
  XOR U6748 ( .A(n6534), .B(n6533), .Z(n6536) );
  XOR U6749 ( .A(n6535), .B(n6536), .Z(n6529) );
  XOR U6750 ( .A(n6530), .B(n6529), .Z(n6578) );
  AND U6751 ( .A(x[75]), .B(y[267]), .Z(n7602) );
  NAND U6752 ( .A(n7602), .B(n6771), .Z(n6506) );
  NANDN U6753 ( .A(n6504), .B(n6503), .Z(n6505) );
  AND U6754 ( .A(n6506), .B(n6505), .Z(n6557) );
  AND U6755 ( .A(x[73]), .B(y[260]), .Z(n6547) );
  NAND U6756 ( .A(n6702), .B(n6547), .Z(n6510) );
  NANDN U6757 ( .A(n6508), .B(n6507), .Z(n6509) );
  AND U6758 ( .A(n6510), .B(n6509), .Z(n6555) );
  ANDN U6759 ( .B(o[75]), .A(n6511), .Z(n6560) );
  NAND U6760 ( .A(y[267]), .B(x[65]), .Z(n6512) );
  XOR U6761 ( .A(n6513), .B(n6512), .Z(n6561) );
  XNOR U6762 ( .A(n6560), .B(n6561), .Z(n6554) );
  XNOR U6763 ( .A(n6555), .B(n6554), .Z(n6556) );
  XOR U6764 ( .A(n6557), .B(n6556), .Z(n6579) );
  XNOR U6765 ( .A(n6578), .B(n6579), .Z(n6581) );
  XOR U6766 ( .A(n6580), .B(n6581), .Z(n6592) );
  NANDN U6767 ( .A(n6515), .B(n6514), .Z(n6519) );
  NANDN U6768 ( .A(n6517), .B(n6516), .Z(n6518) );
  NAND U6769 ( .A(n6519), .B(n6518), .Z(n6591) );
  XNOR U6770 ( .A(n6593), .B(n6594), .Z(n6587) );
  XNOR U6771 ( .A(n6586), .B(n6587), .Z(n6520) );
  XOR U6772 ( .A(n6584), .B(n6520), .Z(N173) );
  NAND U6773 ( .A(n6522), .B(n6521), .Z(n6526) );
  NAND U6774 ( .A(n6524), .B(n6523), .Z(n6525) );
  NAND U6775 ( .A(n6526), .B(n6525), .Z(n6673) );
  NANDN U6776 ( .A(n6528), .B(n6527), .Z(n6532) );
  NAND U6777 ( .A(n6530), .B(n6529), .Z(n6531) );
  AND U6778 ( .A(n6532), .B(n6531), .Z(n6599) );
  NAND U6779 ( .A(n6534), .B(n6533), .Z(n6538) );
  NAND U6780 ( .A(n6536), .B(n6535), .Z(n6537) );
  NAND U6781 ( .A(n6538), .B(n6537), .Z(n6606) );
  AND U6782 ( .A(y[266]), .B(x[72]), .Z(n7893) );
  NAND U6783 ( .A(n7893), .B(n6711), .Z(n6542) );
  NANDN U6784 ( .A(n6540), .B(n6539), .Z(n6541) );
  AND U6785 ( .A(n6542), .B(n6541), .Z(n6637) );
  NAND U6786 ( .A(y[268]), .B(x[65]), .Z(n6543) );
  XNOR U6787 ( .A(n6544), .B(n6543), .Z(n6628) );
  ANDN U6788 ( .B(o[76]), .A(n6545), .Z(n6627) );
  XOR U6789 ( .A(n6628), .B(n6627), .Z(n6635) );
  AND U6790 ( .A(x[70]), .B(y[263]), .Z(n7640) );
  NAND U6791 ( .A(y[267]), .B(x[66]), .Z(n6546) );
  XOR U6792 ( .A(n6547), .B(n6546), .Z(n6640) );
  XNOR U6793 ( .A(n7640), .B(n6640), .Z(n6634) );
  XOR U6794 ( .A(n6635), .B(n6634), .Z(n6636) );
  XNOR U6795 ( .A(n6637), .B(n6636), .Z(n6605) );
  NAND U6796 ( .A(n6549), .B(n6548), .Z(n6553) );
  ANDN U6797 ( .B(n6551), .A(n6550), .Z(n6552) );
  ANDN U6798 ( .B(n6553), .A(n6552), .Z(n6604) );
  XOR U6799 ( .A(n6605), .B(n6604), .Z(n6607) );
  XOR U6800 ( .A(n6606), .B(n6607), .Z(n6598) );
  NANDN U6801 ( .A(n6555), .B(n6554), .Z(n6559) );
  NANDN U6802 ( .A(n6557), .B(n6556), .Z(n6558) );
  AND U6803 ( .A(n6559), .B(n6558), .Z(n6613) );
  AND U6804 ( .A(x[70]), .B(y[267]), .Z(n6908) );
  IV U6805 ( .A(n6908), .Z(n7020) );
  NANDN U6806 ( .A(n7020), .B(n6626), .Z(n6563) );
  NANDN U6807 ( .A(n6561), .B(n6560), .Z(n6562) );
  AND U6808 ( .A(n6563), .B(n6562), .Z(n6619) );
  AND U6809 ( .A(x[76]), .B(y[268]), .Z(n7899) );
  NAND U6810 ( .A(n7899), .B(n6771), .Z(n6567) );
  NAND U6811 ( .A(n6565), .B(n6564), .Z(n6566) );
  AND U6812 ( .A(n6567), .B(n6566), .Z(n6617) );
  AND U6813 ( .A(x[74]), .B(y[259]), .Z(n7509) );
  AND U6814 ( .A(y[261]), .B(x[72]), .Z(n6569) );
  NAND U6815 ( .A(y[258]), .B(x[75]), .Z(n6568) );
  XOR U6816 ( .A(n6569), .B(n6568), .Z(n6623) );
  XNOR U6817 ( .A(n7509), .B(n6623), .Z(n6616) );
  XNOR U6818 ( .A(n6617), .B(n6616), .Z(n6618) );
  XNOR U6819 ( .A(n6619), .B(n6618), .Z(n6611) );
  AND U6820 ( .A(x[74]), .B(y[264]), .Z(n6985) );
  AND U6821 ( .A(x[68]), .B(y[258]), .Z(n6570) );
  NAND U6822 ( .A(n6985), .B(n6570), .Z(n6573) );
  NANDN U6823 ( .A(n6571), .B(n7237), .Z(n6572) );
  AND U6824 ( .A(n6573), .B(n6572), .Z(n6661) );
  AND U6825 ( .A(y[256]), .B(x[77]), .Z(n6575) );
  NAND U6826 ( .A(y[269]), .B(x[64]), .Z(n6574) );
  XNOR U6827 ( .A(n6575), .B(n6574), .Z(n6653) );
  NAND U6828 ( .A(x[76]), .B(y[257]), .Z(n6645) );
  XNOR U6829 ( .A(o[77]), .B(n6645), .Z(n6652) );
  XOR U6830 ( .A(n6653), .B(n6652), .Z(n6659) );
  AND U6831 ( .A(y[266]), .B(x[67]), .Z(n6577) );
  NAND U6832 ( .A(y[264]), .B(x[69]), .Z(n6576) );
  XNOR U6833 ( .A(n6577), .B(n6576), .Z(n6648) );
  NAND U6834 ( .A(x[68]), .B(y[265]), .Z(n6649) );
  XNOR U6835 ( .A(n6648), .B(n6649), .Z(n6658) );
  XOR U6836 ( .A(n6659), .B(n6658), .Z(n6660) );
  XNOR U6837 ( .A(n6661), .B(n6660), .Z(n6610) );
  XOR U6838 ( .A(n6611), .B(n6610), .Z(n6612) );
  XNOR U6839 ( .A(n6613), .B(n6612), .Z(n6600) );
  XOR U6840 ( .A(n6601), .B(n6600), .Z(n6672) );
  NANDN U6841 ( .A(n6579), .B(n6578), .Z(n6583) );
  NAND U6842 ( .A(n6581), .B(n6580), .Z(n6582) );
  AND U6843 ( .A(n6583), .B(n6582), .Z(n6671) );
  XOR U6844 ( .A(n6673), .B(n6674), .Z(n6667) );
  OR U6845 ( .A(n6586), .B(n6584), .Z(n6590) );
  ANDN U6846 ( .B(n6586), .A(n6585), .Z(n6588) );
  OR U6847 ( .A(n6588), .B(n6587), .Z(n6589) );
  AND U6848 ( .A(n6590), .B(n6589), .Z(n6666) );
  NANDN U6849 ( .A(n6592), .B(n6591), .Z(n6596) );
  NANDN U6850 ( .A(n6594), .B(n6593), .Z(n6595) );
  AND U6851 ( .A(n6596), .B(n6595), .Z(n6665) );
  IV U6852 ( .A(n6665), .Z(n6664) );
  XOR U6853 ( .A(n6666), .B(n6664), .Z(n6597) );
  XNOR U6854 ( .A(n6667), .B(n6597), .Z(N174) );
  NANDN U6855 ( .A(n6599), .B(n6598), .Z(n6603) );
  NAND U6856 ( .A(n6601), .B(n6600), .Z(n6602) );
  AND U6857 ( .A(n6603), .B(n6602), .Z(n6760) );
  NAND U6858 ( .A(n6605), .B(n6604), .Z(n6609) );
  NAND U6859 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND U6860 ( .A(n6609), .B(n6608), .Z(n6759) );
  NAND U6861 ( .A(n6611), .B(n6610), .Z(n6615) );
  NANDN U6862 ( .A(n6613), .B(n6612), .Z(n6614) );
  AND U6863 ( .A(n6615), .B(n6614), .Z(n6681) );
  NANDN U6864 ( .A(n6617), .B(n6616), .Z(n6621) );
  NANDN U6865 ( .A(n6619), .B(n6618), .Z(n6620) );
  AND U6866 ( .A(n6621), .B(n6620), .Z(n6687) );
  AND U6867 ( .A(x[75]), .B(y[261]), .Z(n6796) );
  NAND U6868 ( .A(n6796), .B(n6622), .Z(n6625) );
  NANDN U6869 ( .A(n6623), .B(n7509), .Z(n6624) );
  AND U6870 ( .A(n6625), .B(n6624), .Z(n6741) );
  NAND U6871 ( .A(x[71]), .B(y[268]), .Z(n7252) );
  NANDN U6872 ( .A(n7252), .B(n6626), .Z(n6630) );
  NAND U6873 ( .A(n6628), .B(n6627), .Z(n6629) );
  NAND U6874 ( .A(n6630), .B(n6629), .Z(n6740) );
  XNOR U6875 ( .A(n6741), .B(n6740), .Z(n6743) );
  AND U6876 ( .A(x[68]), .B(y[266]), .Z(n7126) );
  AND U6877 ( .A(y[262]), .B(x[72]), .Z(n6632) );
  NAND U6878 ( .A(y[267]), .B(x[67]), .Z(n6631) );
  XOR U6879 ( .A(n6632), .B(n6631), .Z(n6726) );
  XNOR U6880 ( .A(n7018), .B(n6726), .Z(n6735) );
  XOR U6881 ( .A(n7126), .B(n6735), .Z(n6737) );
  AND U6882 ( .A(x[73]), .B(y[261]), .Z(n7330) );
  AND U6883 ( .A(y[260]), .B(x[74]), .Z(n7360) );
  AND U6884 ( .A(y[268]), .B(x[66]), .Z(n6633) );
  XOR U6885 ( .A(n7360), .B(n6633), .Z(n6712) );
  XOR U6886 ( .A(n7330), .B(n6712), .Z(n6736) );
  XOR U6887 ( .A(n6737), .B(n6736), .Z(n6742) );
  XOR U6888 ( .A(n6743), .B(n6742), .Z(n6685) );
  NAND U6889 ( .A(n6635), .B(n6634), .Z(n6639) );
  NANDN U6890 ( .A(n6637), .B(n6636), .Z(n6638) );
  AND U6891 ( .A(n6639), .B(n6638), .Z(n6684) );
  XNOR U6892 ( .A(n6685), .B(n6684), .Z(n6686) );
  XOR U6893 ( .A(n6687), .B(n6686), .Z(n6679) );
  AND U6894 ( .A(x[73]), .B(y[267]), .Z(n7250) );
  NAND U6895 ( .A(n7250), .B(n6711), .Z(n6642) );
  NANDN U6896 ( .A(n6640), .B(n7640), .Z(n6641) );
  AND U6897 ( .A(n6642), .B(n6641), .Z(n6699) );
  AND U6898 ( .A(y[270]), .B(x[64]), .Z(n6644) );
  NAND U6899 ( .A(y[256]), .B(x[78]), .Z(n6643) );
  XNOR U6900 ( .A(n6644), .B(n6643), .Z(n6722) );
  ANDN U6901 ( .B(o[77]), .A(n6645), .Z(n6721) );
  XOR U6902 ( .A(n6722), .B(n6721), .Z(n6697) );
  NAND U6903 ( .A(y[258]), .B(x[76]), .Z(n6646) );
  XNOR U6904 ( .A(n6647), .B(n6646), .Z(n6704) );
  NAND U6905 ( .A(x[77]), .B(y[257]), .Z(n6710) );
  XNOR U6906 ( .A(o[78]), .B(n6710), .Z(n6703) );
  XOR U6907 ( .A(n6704), .B(n6703), .Z(n6696) );
  XOR U6908 ( .A(n6697), .B(n6696), .Z(n6698) );
  XOR U6909 ( .A(n6699), .B(n6698), .Z(n6747) );
  AND U6910 ( .A(x[69]), .B(y[266]), .Z(n6783) );
  NAND U6911 ( .A(n7497), .B(n6783), .Z(n6651) );
  NANDN U6912 ( .A(n6649), .B(n6648), .Z(n6650) );
  AND U6913 ( .A(n6651), .B(n6650), .Z(n6693) );
  AND U6914 ( .A(x[77]), .B(y[269]), .Z(n8225) );
  NAND U6915 ( .A(n8225), .B(n6771), .Z(n6655) );
  NAND U6916 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U6917 ( .A(n6655), .B(n6654), .Z(n6691) );
  NAND U6918 ( .A(y[259]), .B(x[75]), .Z(n6656) );
  XNOR U6919 ( .A(n6657), .B(n6656), .Z(n6717) );
  NAND U6920 ( .A(x[65]), .B(y[269]), .Z(n6718) );
  XNOR U6921 ( .A(n6717), .B(n6718), .Z(n6690) );
  XNOR U6922 ( .A(n6691), .B(n6690), .Z(n6692) );
  XOR U6923 ( .A(n6693), .B(n6692), .Z(n6746) );
  XOR U6924 ( .A(n6747), .B(n6746), .Z(n6749) );
  NAND U6925 ( .A(n6659), .B(n6658), .Z(n6663) );
  NANDN U6926 ( .A(n6661), .B(n6660), .Z(n6662) );
  AND U6927 ( .A(n6663), .B(n6662), .Z(n6748) );
  XNOR U6928 ( .A(n6749), .B(n6748), .Z(n6678) );
  XNOR U6929 ( .A(n6679), .B(n6678), .Z(n6680) );
  XNOR U6930 ( .A(n6681), .B(n6680), .Z(n6761) );
  XNOR U6931 ( .A(n6762), .B(n6761), .Z(n6755) );
  OR U6932 ( .A(n6666), .B(n6664), .Z(n6670) );
  ANDN U6933 ( .B(n6666), .A(n6665), .Z(n6668) );
  OR U6934 ( .A(n6668), .B(n6667), .Z(n6669) );
  AND U6935 ( .A(n6670), .B(n6669), .Z(n6754) );
  NANDN U6936 ( .A(n6672), .B(n6671), .Z(n6676) );
  NAND U6937 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U6938 ( .A(n6676), .B(n6675), .Z(n6753) );
  IV U6939 ( .A(n6753), .Z(n6752) );
  XOR U6940 ( .A(n6754), .B(n6752), .Z(n6677) );
  XNOR U6941 ( .A(n6755), .B(n6677), .Z(N175) );
  NANDN U6942 ( .A(n6679), .B(n6678), .Z(n6683) );
  NANDN U6943 ( .A(n6681), .B(n6680), .Z(n6682) );
  AND U6944 ( .A(n6683), .B(n6682), .Z(n6857) );
  NANDN U6945 ( .A(n6685), .B(n6684), .Z(n6689) );
  NAND U6946 ( .A(n6687), .B(n6686), .Z(n6688) );
  NAND U6947 ( .A(n6689), .B(n6688), .Z(n6825) );
  NANDN U6948 ( .A(n6691), .B(n6690), .Z(n6695) );
  NANDN U6949 ( .A(n6693), .B(n6692), .Z(n6694) );
  AND U6950 ( .A(n6695), .B(n6694), .Z(n6832) );
  NAND U6951 ( .A(n6697), .B(n6696), .Z(n6701) );
  NANDN U6952 ( .A(n6699), .B(n6698), .Z(n6700) );
  AND U6953 ( .A(n6701), .B(n6700), .Z(n6830) );
  NAND U6954 ( .A(x[76]), .B(y[263]), .Z(n7244) );
  NANDN U6955 ( .A(n7244), .B(n6702), .Z(n6706) );
  NAND U6956 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U6957 ( .A(n6706), .B(n6705), .Z(n6806) );
  AND U6958 ( .A(y[258]), .B(x[77]), .Z(n7628) );
  NAND U6959 ( .A(y[260]), .B(x[75]), .Z(n6707) );
  XNOR U6960 ( .A(n7628), .B(n6707), .Z(n6810) );
  AND U6961 ( .A(x[76]), .B(y[259]), .Z(n6809) );
  XOR U6962 ( .A(n6810), .B(n6809), .Z(n6804) );
  AND U6963 ( .A(y[256]), .B(x[79]), .Z(n6709) );
  NAND U6964 ( .A(y[271]), .B(x[64]), .Z(n6708) );
  XNOR U6965 ( .A(n6709), .B(n6708), .Z(n6773) );
  ANDN U6966 ( .B(o[78]), .A(n6710), .Z(n6772) );
  XNOR U6967 ( .A(n6773), .B(n6772), .Z(n6803) );
  XNOR U6968 ( .A(n6804), .B(n6803), .Z(n6805) );
  XOR U6969 ( .A(n6806), .B(n6805), .Z(n6838) );
  NAND U6970 ( .A(x[74]), .B(y[268]), .Z(n7642) );
  NANDN U6971 ( .A(n7642), .B(n6711), .Z(n6714) );
  NAND U6972 ( .A(n7330), .B(n6712), .Z(n6713) );
  AND U6973 ( .A(n6714), .B(n6713), .Z(n6836) );
  AND U6974 ( .A(x[75]), .B(y[264]), .Z(n6716) );
  NAND U6975 ( .A(n6716), .B(n6715), .Z(n6720) );
  NANDN U6976 ( .A(n6718), .B(n6717), .Z(n6719) );
  NAND U6977 ( .A(n6720), .B(n6719), .Z(n6835) );
  XNOR U6978 ( .A(n6836), .B(n6835), .Z(n6837) );
  XNOR U6979 ( .A(n6838), .B(n6837), .Z(n6829) );
  XNOR U6980 ( .A(n6830), .B(n6829), .Z(n6831) );
  XNOR U6981 ( .A(n6832), .B(n6831), .Z(n6824) );
  AND U6982 ( .A(x[78]), .B(y[270]), .Z(n8460) );
  NAND U6983 ( .A(n8460), .B(n6771), .Z(n6724) );
  NAND U6984 ( .A(n6722), .B(n6721), .Z(n6723) );
  AND U6985 ( .A(n6724), .B(n6723), .Z(n6798) );
  AND U6986 ( .A(x[72]), .B(y[267]), .Z(n7101) );
  NANDN U6987 ( .A(n6725), .B(n7101), .Z(n6728) );
  NANDN U6988 ( .A(n6726), .B(n7018), .Z(n6727) );
  NAND U6989 ( .A(n6728), .B(n6727), .Z(n6797) );
  XNOR U6990 ( .A(n6798), .B(n6797), .Z(n6800) );
  AND U6991 ( .A(y[261]), .B(x[74]), .Z(n6730) );
  NAND U6992 ( .A(y[267]), .B(x[68]), .Z(n6729) );
  XNOR U6993 ( .A(n6730), .B(n6729), .Z(n6778) );
  AND U6994 ( .A(x[71]), .B(y[264]), .Z(n6777) );
  XOR U6995 ( .A(n6778), .B(n6777), .Z(n6785) );
  NAND U6996 ( .A(x[70]), .B(y[265]), .Z(n6938) );
  XNOR U6997 ( .A(n6938), .B(n6783), .Z(n6784) );
  AND U6998 ( .A(y[262]), .B(x[73]), .Z(n6732) );
  NAND U6999 ( .A(y[269]), .B(x[66]), .Z(n6731) );
  XNOR U7000 ( .A(n6732), .B(n6731), .Z(n6788) );
  NAND U7001 ( .A(x[67]), .B(y[268]), .Z(n6789) );
  AND U7002 ( .A(y[263]), .B(x[72]), .Z(n6734) );
  NAND U7003 ( .A(y[270]), .B(x[65]), .Z(n6733) );
  XNOR U7004 ( .A(n6734), .B(n6733), .Z(n6768) );
  NAND U7005 ( .A(x[78]), .B(y[257]), .Z(n6794) );
  XNOR U7006 ( .A(o[79]), .B(n6794), .Z(n6767) );
  XOR U7007 ( .A(n6768), .B(n6767), .Z(n6817) );
  XOR U7008 ( .A(n6818), .B(n6817), .Z(n6820) );
  XOR U7009 ( .A(n6819), .B(n6820), .Z(n6799) );
  XOR U7010 ( .A(n6800), .B(n6799), .Z(n6842) );
  NAND U7011 ( .A(n7126), .B(n6735), .Z(n6739) );
  NAND U7012 ( .A(n6737), .B(n6736), .Z(n6738) );
  AND U7013 ( .A(n6739), .B(n6738), .Z(n6841) );
  XNOR U7014 ( .A(n6842), .B(n6841), .Z(n6844) );
  NANDN U7015 ( .A(n6741), .B(n6740), .Z(n6745) );
  NAND U7016 ( .A(n6743), .B(n6742), .Z(n6744) );
  AND U7017 ( .A(n6745), .B(n6744), .Z(n6843) );
  XOR U7018 ( .A(n6844), .B(n6843), .Z(n6823) );
  XOR U7019 ( .A(n6825), .B(n6826), .Z(n6854) );
  NAND U7020 ( .A(n6747), .B(n6746), .Z(n6751) );
  NAND U7021 ( .A(n6749), .B(n6748), .Z(n6750) );
  AND U7022 ( .A(n6751), .B(n6750), .Z(n6855) );
  XOR U7023 ( .A(n6854), .B(n6855), .Z(n6856) );
  XOR U7024 ( .A(n6857), .B(n6856), .Z(n6850) );
  OR U7025 ( .A(n6754), .B(n6752), .Z(n6758) );
  ANDN U7026 ( .B(n6754), .A(n6753), .Z(n6756) );
  OR U7027 ( .A(n6756), .B(n6755), .Z(n6757) );
  AND U7028 ( .A(n6758), .B(n6757), .Z(n6849) );
  NANDN U7029 ( .A(n6760), .B(n6759), .Z(n6764) );
  NAND U7030 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U7031 ( .A(n6764), .B(n6763), .Z(n6848) );
  IV U7032 ( .A(n6848), .Z(n6847) );
  XOR U7033 ( .A(n6849), .B(n6847), .Z(n6765) );
  XNOR U7034 ( .A(n6850), .B(n6765), .Z(N176) );
  AND U7035 ( .A(x[72]), .B(y[270]), .Z(n7518) );
  NAND U7036 ( .A(n7518), .B(n6766), .Z(n6770) );
  NAND U7037 ( .A(n6768), .B(n6767), .Z(n6769) );
  AND U7038 ( .A(n6770), .B(n6769), .Z(n6887) );
  AND U7039 ( .A(x[79]), .B(y[271]), .Z(n8840) );
  NAND U7040 ( .A(n8840), .B(n6771), .Z(n6775) );
  NAND U7041 ( .A(n6773), .B(n6772), .Z(n6774) );
  NAND U7042 ( .A(n6775), .B(n6774), .Z(n6886) );
  AND U7043 ( .A(x[74]), .B(y[267]), .Z(n7373) );
  NAND U7044 ( .A(n7373), .B(n6776), .Z(n6780) );
  NAND U7045 ( .A(n6778), .B(n6777), .Z(n6779) );
  NAND U7046 ( .A(n6780), .B(n6779), .Z(n6925) );
  AND U7047 ( .A(x[64]), .B(y[272]), .Z(n6947) );
  NAND U7048 ( .A(x[80]), .B(y[256]), .Z(n6948) );
  XNOR U7049 ( .A(n6947), .B(n6948), .Z(n6950) );
  NAND U7050 ( .A(x[79]), .B(y[257]), .Z(n6935) );
  XNOR U7051 ( .A(o[80]), .B(n6935), .Z(n6949) );
  XOR U7052 ( .A(n6950), .B(n6949), .Z(n6924) );
  NAND U7053 ( .A(y[265]), .B(x[71]), .Z(n6781) );
  XNOR U7054 ( .A(n6782), .B(n6781), .Z(n6940) );
  AND U7055 ( .A(x[74]), .B(y[262]), .Z(n6939) );
  XOR U7056 ( .A(n6940), .B(n6939), .Z(n6923) );
  XOR U7057 ( .A(n6924), .B(n6923), .Z(n6926) );
  XOR U7058 ( .A(n6925), .B(n6926), .Z(n6888) );
  XOR U7059 ( .A(n6889), .B(n6888), .Z(n6920) );
  NANDN U7060 ( .A(n6783), .B(n6938), .Z(n6787) );
  NANDN U7061 ( .A(n6785), .B(n6784), .Z(n6786) );
  AND U7062 ( .A(n6787), .B(n6786), .Z(n6918) );
  NAND U7063 ( .A(x[73]), .B(y[269]), .Z(n7624) );
  NANDN U7064 ( .A(n7624), .B(n7242), .Z(n6791) );
  NANDN U7065 ( .A(n6789), .B(n6788), .Z(n6790) );
  AND U7066 ( .A(n6791), .B(n6790), .Z(n6958) );
  NAND U7067 ( .A(y[271]), .B(x[65]), .Z(n6792) );
  XNOR U7068 ( .A(n6793), .B(n6792), .Z(n6944) );
  ANDN U7069 ( .B(o[79]), .A(n6794), .Z(n6943) );
  XOR U7070 ( .A(n6944), .B(n6943), .Z(n6956) );
  NAND U7071 ( .A(y[258]), .B(x[78]), .Z(n6795) );
  XNOR U7072 ( .A(n6796), .B(n6795), .Z(n6898) );
  NAND U7073 ( .A(x[68]), .B(y[268]), .Z(n6899) );
  XNOR U7074 ( .A(n6898), .B(n6899), .Z(n6955) );
  XOR U7075 ( .A(n6956), .B(n6955), .Z(n6957) );
  XOR U7076 ( .A(n6958), .B(n6957), .Z(n6917) );
  NANDN U7077 ( .A(n6798), .B(n6797), .Z(n6802) );
  NAND U7078 ( .A(n6800), .B(n6799), .Z(n6801) );
  NAND U7079 ( .A(n6802), .B(n6801), .Z(n6881) );
  XNOR U7080 ( .A(n6880), .B(n6881), .Z(n6883) );
  NANDN U7081 ( .A(n6804), .B(n6803), .Z(n6808) );
  NAND U7082 ( .A(n6806), .B(n6805), .Z(n6807) );
  AND U7083 ( .A(n6808), .B(n6807), .Z(n6914) );
  AND U7084 ( .A(x[77]), .B(y[260]), .Z(n6910) );
  AND U7085 ( .A(x[75]), .B(y[258]), .Z(n7470) );
  NAND U7086 ( .A(n6910), .B(n7470), .Z(n6812) );
  NAND U7087 ( .A(n6810), .B(n6809), .Z(n6811) );
  AND U7088 ( .A(n6812), .B(n6811), .Z(n6895) );
  AND U7089 ( .A(y[263]), .B(x[73]), .Z(n6814) );
  NAND U7090 ( .A(y[270]), .B(x[66]), .Z(n6813) );
  XNOR U7091 ( .A(n6814), .B(n6813), .Z(n6902) );
  NAND U7092 ( .A(x[67]), .B(y[269]), .Z(n6903) );
  XNOR U7093 ( .A(n6902), .B(n6903), .Z(n6893) );
  AND U7094 ( .A(x[76]), .B(y[260]), .Z(n7612) );
  AND U7095 ( .A(y[259]), .B(x[77]), .Z(n6816) );
  NAND U7096 ( .A(y[267]), .B(x[69]), .Z(n6815) );
  XOR U7097 ( .A(n6816), .B(n6815), .Z(n6930) );
  XNOR U7098 ( .A(n7612), .B(n6930), .Z(n6892) );
  XOR U7099 ( .A(n6893), .B(n6892), .Z(n6894) );
  NAND U7100 ( .A(n6818), .B(n6817), .Z(n6822) );
  NAND U7101 ( .A(n6820), .B(n6819), .Z(n6821) );
  AND U7102 ( .A(n6822), .B(n6821), .Z(n6912) );
  XOR U7103 ( .A(n6911), .B(n6912), .Z(n6913) );
  XOR U7104 ( .A(n6883), .B(n6882), .Z(n6862) );
  NANDN U7105 ( .A(n6824), .B(n6823), .Z(n6828) );
  NANDN U7106 ( .A(n6826), .B(n6825), .Z(n6827) );
  AND U7107 ( .A(n6828), .B(n6827), .Z(n6861) );
  NANDN U7108 ( .A(n6830), .B(n6829), .Z(n6834) );
  NANDN U7109 ( .A(n6832), .B(n6831), .Z(n6833) );
  AND U7110 ( .A(n6834), .B(n6833), .Z(n6877) );
  NANDN U7111 ( .A(n6836), .B(n6835), .Z(n6840) );
  NANDN U7112 ( .A(n6838), .B(n6837), .Z(n6839) );
  AND U7113 ( .A(n6840), .B(n6839), .Z(n6875) );
  NANDN U7114 ( .A(n6842), .B(n6841), .Z(n6846) );
  NAND U7115 ( .A(n6844), .B(n6843), .Z(n6845) );
  AND U7116 ( .A(n6846), .B(n6845), .Z(n6874) );
  XNOR U7117 ( .A(n6875), .B(n6874), .Z(n6876) );
  XOR U7118 ( .A(n6877), .B(n6876), .Z(n6864) );
  XNOR U7119 ( .A(n6863), .B(n6864), .Z(n6870) );
  OR U7120 ( .A(n6849), .B(n6847), .Z(n6853) );
  ANDN U7121 ( .B(n6849), .A(n6848), .Z(n6851) );
  OR U7122 ( .A(n6851), .B(n6850), .Z(n6852) );
  AND U7123 ( .A(n6853), .B(n6852), .Z(n6868) );
  NAND U7124 ( .A(n6855), .B(n6854), .Z(n6859) );
  NANDN U7125 ( .A(n6857), .B(n6856), .Z(n6858) );
  AND U7126 ( .A(n6859), .B(n6858), .Z(n6869) );
  IV U7127 ( .A(n6869), .Z(n6867) );
  XOR U7128 ( .A(n6868), .B(n6867), .Z(n6860) );
  XNOR U7129 ( .A(n6870), .B(n6860), .Z(N177) );
  NANDN U7130 ( .A(n6862), .B(n6861), .Z(n6866) );
  NANDN U7131 ( .A(n6864), .B(n6863), .Z(n6865) );
  AND U7132 ( .A(n6866), .B(n6865), .Z(n7064) );
  NANDN U7133 ( .A(n6867), .B(n6868), .Z(n6873) );
  NOR U7134 ( .A(n6869), .B(n6868), .Z(n6871) );
  OR U7135 ( .A(n6871), .B(n6870), .Z(n6872) );
  AND U7136 ( .A(n6873), .B(n6872), .Z(n7065) );
  NANDN U7137 ( .A(n6875), .B(n6874), .Z(n6879) );
  NANDN U7138 ( .A(n6877), .B(n6876), .Z(n6878) );
  AND U7139 ( .A(n6879), .B(n6878), .Z(n7061) );
  NANDN U7140 ( .A(n6881), .B(n6880), .Z(n6885) );
  NAND U7141 ( .A(n6883), .B(n6882), .Z(n6884) );
  AND U7142 ( .A(n6885), .B(n6884), .Z(n6965) );
  NANDN U7143 ( .A(n6887), .B(n6886), .Z(n6891) );
  NAND U7144 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U7145 ( .A(n6891), .B(n6890), .Z(n7049) );
  NAND U7146 ( .A(n6893), .B(n6892), .Z(n6897) );
  NANDN U7147 ( .A(n6895), .B(n6894), .Z(n6896) );
  AND U7148 ( .A(n6897), .B(n6896), .Z(n7047) );
  NAND U7149 ( .A(x[78]), .B(y[261]), .Z(n7229) );
  NANDN U7150 ( .A(n7229), .B(n7470), .Z(n6901) );
  NANDN U7151 ( .A(n6899), .B(n6898), .Z(n6900) );
  AND U7152 ( .A(n6901), .B(n6900), .Z(n7041) );
  AND U7153 ( .A(y[270]), .B(x[73]), .Z(n7888) );
  NANDN U7154 ( .A(n7027), .B(n7888), .Z(n6905) );
  NANDN U7155 ( .A(n6903), .B(n6902), .Z(n6904) );
  NAND U7156 ( .A(n6905), .B(n6904), .Z(n7040) );
  XNOR U7157 ( .A(n7041), .B(n7040), .Z(n7043) );
  AND U7158 ( .A(x[71]), .B(y[266]), .Z(n7035) );
  AND U7159 ( .A(y[265]), .B(x[72]), .Z(n6907) );
  NAND U7160 ( .A(y[268]), .B(x[69]), .Z(n6906) );
  XNOR U7161 ( .A(n6907), .B(n6906), .Z(n7019) );
  XOR U7162 ( .A(n7019), .B(n6908), .Z(n7034) );
  XOR U7163 ( .A(n7035), .B(n7034), .Z(n7037) );
  NAND U7164 ( .A(y[269]), .B(x[68]), .Z(n6909) );
  XNOR U7165 ( .A(n6910), .B(n6909), .Z(n6980) );
  NAND U7166 ( .A(x[75]), .B(y[262]), .Z(n6981) );
  XNOR U7167 ( .A(n6980), .B(n6981), .Z(n7036) );
  XOR U7168 ( .A(n7037), .B(n7036), .Z(n7042) );
  XOR U7169 ( .A(n7043), .B(n7042), .Z(n7046) );
  NAND U7170 ( .A(n6912), .B(n6911), .Z(n6916) );
  NANDN U7171 ( .A(n6914), .B(n6913), .Z(n6915) );
  NAND U7172 ( .A(n6916), .B(n6915), .Z(n6962) );
  XOR U7173 ( .A(n6963), .B(n6962), .Z(n6964) );
  NANDN U7174 ( .A(n6918), .B(n6917), .Z(n6922) );
  NANDN U7175 ( .A(n6920), .B(n6919), .Z(n6921) );
  AND U7176 ( .A(n6922), .B(n6921), .Z(n6971) );
  NAND U7177 ( .A(n6924), .B(n6923), .Z(n6928) );
  NAND U7178 ( .A(n6926), .B(n6925), .Z(n6927) );
  AND U7179 ( .A(n6928), .B(n6927), .Z(n7055) );
  AND U7180 ( .A(x[77]), .B(y[267]), .Z(n7907) );
  AND U7181 ( .A(x[69]), .B(y[259]), .Z(n6929) );
  NAND U7182 ( .A(n7907), .B(n6929), .Z(n6932) );
  NANDN U7183 ( .A(n6930), .B(n7612), .Z(n6931) );
  AND U7184 ( .A(n6932), .B(n6931), .Z(n7003) );
  AND U7185 ( .A(y[264]), .B(x[73]), .Z(n6934) );
  NAND U7186 ( .A(y[272]), .B(x[65]), .Z(n6933) );
  XNOR U7187 ( .A(n6934), .B(n6933), .Z(n7024) );
  ANDN U7188 ( .B(o[80]), .A(n6935), .Z(n7023) );
  XOR U7189 ( .A(n7024), .B(n7023), .Z(n7001) );
  AND U7190 ( .A(y[258]), .B(x[79]), .Z(n6937) );
  NAND U7191 ( .A(y[261]), .B(x[76]), .Z(n6936) );
  XNOR U7192 ( .A(n6937), .B(n6936), .Z(n6975) );
  NAND U7193 ( .A(x[78]), .B(y[259]), .Z(n6976) );
  XOR U7194 ( .A(n7001), .B(n7000), .Z(n7002) );
  XNOR U7195 ( .A(n7003), .B(n7002), .Z(n7053) );
  NANDN U7196 ( .A(n6938), .B(n7035), .Z(n6942) );
  NAND U7197 ( .A(n6940), .B(n6939), .Z(n6941) );
  AND U7198 ( .A(n6942), .B(n6941), .Z(n7013) );
  NAND U7199 ( .A(x[72]), .B(y[271]), .Z(n7706) );
  AND U7200 ( .A(x[65]), .B(y[264]), .Z(n7104) );
  NANDN U7201 ( .A(n7706), .B(n7104), .Z(n6946) );
  NAND U7202 ( .A(n6944), .B(n6943), .Z(n6945) );
  NAND U7203 ( .A(n6946), .B(n6945), .Z(n7012) );
  XNOR U7204 ( .A(n7013), .B(n7012), .Z(n7015) );
  NANDN U7205 ( .A(n6948), .B(n6947), .Z(n6952) );
  NAND U7206 ( .A(n6950), .B(n6949), .Z(n6951) );
  AND U7207 ( .A(n6952), .B(n6951), .Z(n7009) );
  AND U7208 ( .A(x[64]), .B(y[273]), .Z(n6989) );
  NAND U7209 ( .A(x[81]), .B(y[256]), .Z(n6990) );
  NAND U7210 ( .A(x[80]), .B(y[257]), .Z(n6986) );
  XNOR U7211 ( .A(o[81]), .B(n6986), .Z(n6991) );
  XOR U7212 ( .A(n6992), .B(n6991), .Z(n7007) );
  AND U7213 ( .A(y[263]), .B(x[74]), .Z(n6954) );
  NAND U7214 ( .A(y[271]), .B(x[66]), .Z(n6953) );
  XNOR U7215 ( .A(n6954), .B(n6953), .Z(n7028) );
  NAND U7216 ( .A(x[67]), .B(y[270]), .Z(n7029) );
  XNOR U7217 ( .A(n7028), .B(n7029), .Z(n7006) );
  XOR U7218 ( .A(n7007), .B(n7006), .Z(n7008) );
  XNOR U7219 ( .A(n7009), .B(n7008), .Z(n7014) );
  XOR U7220 ( .A(n7015), .B(n7014), .Z(n7052) );
  XOR U7221 ( .A(n7053), .B(n7052), .Z(n7054) );
  NAND U7222 ( .A(n6956), .B(n6955), .Z(n6960) );
  NANDN U7223 ( .A(n6958), .B(n6957), .Z(n6959) );
  AND U7224 ( .A(n6960), .B(n6959), .Z(n6969) );
  XOR U7225 ( .A(n6968), .B(n6969), .Z(n6970) );
  XOR U7226 ( .A(n6971), .B(n6970), .Z(n7058) );
  XOR U7227 ( .A(n7059), .B(n7058), .Z(n7060) );
  XNOR U7228 ( .A(n7061), .B(n7060), .Z(n7066) );
  XNOR U7229 ( .A(n7065), .B(n7066), .Z(n6961) );
  XOR U7230 ( .A(n7064), .B(n6961), .Z(N178) );
  NAND U7231 ( .A(n6963), .B(n6962), .Z(n6967) );
  NANDN U7232 ( .A(n6965), .B(n6964), .Z(n6966) );
  AND U7233 ( .A(n6967), .B(n6966), .Z(n7176) );
  NAND U7234 ( .A(n6969), .B(n6968), .Z(n6973) );
  NANDN U7235 ( .A(n6971), .B(n6970), .Z(n6972) );
  AND U7236 ( .A(n6973), .B(n6972), .Z(n7174) );
  AND U7237 ( .A(x[76]), .B(y[258]), .Z(n7320) );
  AND U7238 ( .A(x[79]), .B(y[261]), .Z(n6974) );
  NAND U7239 ( .A(n7320), .B(n6974), .Z(n6978) );
  NANDN U7240 ( .A(n6976), .B(n6975), .Z(n6977) );
  AND U7241 ( .A(n6978), .B(n6977), .Z(n7153) );
  NAND U7242 ( .A(n8225), .B(n6979), .Z(n6983) );
  NANDN U7243 ( .A(n6981), .B(n6980), .Z(n6982) );
  AND U7244 ( .A(n6983), .B(n6982), .Z(n7143) );
  NAND U7245 ( .A(y[273]), .B(x[65]), .Z(n6984) );
  XNOR U7246 ( .A(n6985), .B(n6984), .Z(n7106) );
  ANDN U7247 ( .B(o[81]), .A(n6986), .Z(n7105) );
  XOR U7248 ( .A(n7106), .B(n7105), .Z(n7141) );
  NAND U7249 ( .A(y[259]), .B(x[79]), .Z(n6987) );
  XNOR U7250 ( .A(n6988), .B(n6987), .Z(n7096) );
  NAND U7251 ( .A(x[78]), .B(y[260]), .Z(n7097) );
  XNOR U7252 ( .A(n7096), .B(n7097), .Z(n7140) );
  XOR U7253 ( .A(n7141), .B(n7140), .Z(n7142) );
  XNOR U7254 ( .A(n7143), .B(n7142), .Z(n7152) );
  XNOR U7255 ( .A(n7153), .B(n7152), .Z(n7155) );
  NANDN U7256 ( .A(n6990), .B(n6989), .Z(n6994) );
  NAND U7257 ( .A(n6992), .B(n6991), .Z(n6993) );
  AND U7258 ( .A(n6994), .B(n6993), .Z(n7165) );
  AND U7259 ( .A(y[263]), .B(x[75]), .Z(n6996) );
  NAND U7260 ( .A(y[258]), .B(x[80]), .Z(n6995) );
  XNOR U7261 ( .A(n6996), .B(n6995), .Z(n7092) );
  NAND U7262 ( .A(x[66]), .B(y[272]), .Z(n7093) );
  XNOR U7263 ( .A(n7092), .B(n7093), .Z(n7164) );
  AND U7264 ( .A(y[268]), .B(x[70]), .Z(n6998) );
  NAND U7265 ( .A(y[269]), .B(x[69]), .Z(n6997) );
  XNOR U7266 ( .A(n6998), .B(n6997), .Z(n7088) );
  NAND U7267 ( .A(y[270]), .B(x[68]), .Z(n6999) );
  XNOR U7268 ( .A(n7893), .B(n6999), .Z(n7127) );
  NAND U7269 ( .A(x[71]), .B(y[267]), .Z(n7128) );
  XNOR U7270 ( .A(n7127), .B(n7128), .Z(n7087) );
  XOR U7271 ( .A(n7088), .B(n7087), .Z(n7166) );
  XOR U7272 ( .A(n7167), .B(n7166), .Z(n7154) );
  XOR U7273 ( .A(n7155), .B(n7154), .Z(n7075) );
  NAND U7274 ( .A(n7001), .B(n7000), .Z(n7005) );
  NANDN U7275 ( .A(n7003), .B(n7002), .Z(n7004) );
  AND U7276 ( .A(n7005), .B(n7004), .Z(n7146) );
  NAND U7277 ( .A(n7007), .B(n7006), .Z(n7011) );
  NANDN U7278 ( .A(n7009), .B(n7008), .Z(n7010) );
  NAND U7279 ( .A(n7011), .B(n7010), .Z(n7147) );
  XNOR U7280 ( .A(n7146), .B(n7147), .Z(n7148) );
  NANDN U7281 ( .A(n7013), .B(n7012), .Z(n7017) );
  NAND U7282 ( .A(n7015), .B(n7014), .Z(n7016) );
  NAND U7283 ( .A(n7017), .B(n7016), .Z(n7149) );
  XNOR U7284 ( .A(n7148), .B(n7149), .Z(n7074) );
  AND U7285 ( .A(x[72]), .B(y[268]), .Z(n7366) );
  NAND U7286 ( .A(n7366), .B(n7018), .Z(n7022) );
  NANDN U7287 ( .A(n7020), .B(n7019), .Z(n7021) );
  NAND U7288 ( .A(n7022), .B(n7021), .Z(n7159) );
  NAND U7289 ( .A(x[73]), .B(y[272]), .Z(n7991) );
  NANDN U7290 ( .A(n7991), .B(n7104), .Z(n7026) );
  NAND U7291 ( .A(n7024), .B(n7023), .Z(n7025) );
  NAND U7292 ( .A(n7026), .B(n7025), .Z(n7158) );
  XOR U7293 ( .A(n7159), .B(n7158), .Z(n7161) );
  NAND U7294 ( .A(x[74]), .B(y[271]), .Z(n7992) );
  OR U7295 ( .A(n7027), .B(n7992), .Z(n7031) );
  NANDN U7296 ( .A(n7029), .B(n7028), .Z(n7030) );
  AND U7297 ( .A(n7031), .B(n7030), .Z(n7137) );
  AND U7298 ( .A(x[64]), .B(y[274]), .Z(n7109) );
  NAND U7299 ( .A(x[82]), .B(y[256]), .Z(n7110) );
  XNOR U7300 ( .A(n7109), .B(n7110), .Z(n7112) );
  NAND U7301 ( .A(x[81]), .B(y[257]), .Z(n7131) );
  XNOR U7302 ( .A(o[82]), .B(n7131), .Z(n7111) );
  XOR U7303 ( .A(n7112), .B(n7111), .Z(n7135) );
  AND U7304 ( .A(y[261]), .B(x[77]), .Z(n7033) );
  NAND U7305 ( .A(y[271]), .B(x[67]), .Z(n7032) );
  XNOR U7306 ( .A(n7033), .B(n7032), .Z(n7118) );
  NAND U7307 ( .A(x[76]), .B(y[262]), .Z(n7119) );
  XNOR U7308 ( .A(n7118), .B(n7119), .Z(n7134) );
  XOR U7309 ( .A(n7135), .B(n7134), .Z(n7136) );
  XNOR U7310 ( .A(n7137), .B(n7136), .Z(n7160) );
  XOR U7311 ( .A(n7161), .B(n7160), .Z(n7081) );
  NAND U7312 ( .A(n7035), .B(n7034), .Z(n7039) );
  NAND U7313 ( .A(n7037), .B(n7036), .Z(n7038) );
  AND U7314 ( .A(n7039), .B(n7038), .Z(n7080) );
  XNOR U7315 ( .A(n7081), .B(n7080), .Z(n7082) );
  NANDN U7316 ( .A(n7041), .B(n7040), .Z(n7045) );
  NAND U7317 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7318 ( .A(n7045), .B(n7044), .Z(n7083) );
  XNOR U7319 ( .A(n7082), .B(n7083), .Z(n7076) );
  XOR U7320 ( .A(n7077), .B(n7076), .Z(n7071) );
  NANDN U7321 ( .A(n7047), .B(n7046), .Z(n7051) );
  NANDN U7322 ( .A(n7049), .B(n7048), .Z(n7050) );
  AND U7323 ( .A(n7051), .B(n7050), .Z(n7069) );
  NAND U7324 ( .A(n7053), .B(n7052), .Z(n7057) );
  NANDN U7325 ( .A(n7055), .B(n7054), .Z(n7056) );
  NAND U7326 ( .A(n7057), .B(n7056), .Z(n7068) );
  XOR U7327 ( .A(n7174), .B(n7173), .Z(n7175) );
  XNOR U7328 ( .A(n7176), .B(n7175), .Z(n7172) );
  NAND U7329 ( .A(n7059), .B(n7058), .Z(n7063) );
  NANDN U7330 ( .A(n7061), .B(n7060), .Z(n7062) );
  NAND U7331 ( .A(n7063), .B(n7062), .Z(n7171) );
  XOR U7332 ( .A(n7171), .B(n7170), .Z(n7067) );
  XNOR U7333 ( .A(n7172), .B(n7067), .Z(N179) );
  NANDN U7334 ( .A(n7069), .B(n7068), .Z(n7073) );
  NANDN U7335 ( .A(n7071), .B(n7070), .Z(n7072) );
  AND U7336 ( .A(n7073), .B(n7072), .Z(n7183) );
  NANDN U7337 ( .A(n7075), .B(n7074), .Z(n7079) );
  NAND U7338 ( .A(n7077), .B(n7076), .Z(n7078) );
  AND U7339 ( .A(n7079), .B(n7078), .Z(n7181) );
  NANDN U7340 ( .A(n7081), .B(n7080), .Z(n7085) );
  NANDN U7341 ( .A(n7083), .B(n7082), .Z(n7084) );
  AND U7342 ( .A(n7085), .B(n7084), .Z(n7196) );
  AND U7343 ( .A(x[70]), .B(y[269]), .Z(n7133) );
  AND U7344 ( .A(x[69]), .B(y[268]), .Z(n7086) );
  NAND U7345 ( .A(n7133), .B(n7086), .Z(n7090) );
  NAND U7346 ( .A(n7088), .B(n7087), .Z(n7089) );
  AND U7347 ( .A(n7090), .B(n7089), .Z(n7285) );
  AND U7348 ( .A(x[80]), .B(y[263]), .Z(n7091) );
  NAND U7349 ( .A(n7091), .B(n7470), .Z(n7095) );
  NANDN U7350 ( .A(n7093), .B(n7092), .Z(n7094) );
  AND U7351 ( .A(n7095), .B(n7094), .Z(n7283) );
  AND U7352 ( .A(x[79]), .B(y[265]), .Z(n7918) );
  NAND U7353 ( .A(n7918), .B(n7237), .Z(n7099) );
  NANDN U7354 ( .A(n7097), .B(n7096), .Z(n7098) );
  AND U7355 ( .A(n7099), .B(n7098), .Z(n7261) );
  NAND U7356 ( .A(y[274]), .B(x[65]), .Z(n7100) );
  XNOR U7357 ( .A(n7101), .B(n7100), .Z(n7228) );
  AND U7358 ( .A(y[262]), .B(x[77]), .Z(n7103) );
  NAND U7359 ( .A(y[273]), .B(x[66]), .Z(n7102) );
  XNOR U7360 ( .A(n7103), .B(n7102), .Z(n7243) );
  XOR U7361 ( .A(n7259), .B(n7258), .Z(n7260) );
  XNOR U7362 ( .A(n7261), .B(n7260), .Z(n7282) );
  XNOR U7363 ( .A(n7283), .B(n7282), .Z(n7284) );
  XOR U7364 ( .A(n7285), .B(n7284), .Z(n7194) );
  NAND U7365 ( .A(x[74]), .B(y[273]), .Z(n8315) );
  NANDN U7366 ( .A(n8315), .B(n7104), .Z(n7108) );
  NAND U7367 ( .A(n7106), .B(n7105), .Z(n7107) );
  AND U7368 ( .A(n7108), .B(n7107), .Z(n7208) );
  NANDN U7369 ( .A(n7110), .B(n7109), .Z(n7114) );
  NAND U7370 ( .A(n7112), .B(n7111), .Z(n7113) );
  AND U7371 ( .A(n7114), .B(n7113), .Z(n7206) );
  AND U7372 ( .A(y[266]), .B(x[73]), .Z(n7116) );
  NAND U7373 ( .A(y[259]), .B(x[80]), .Z(n7115) );
  XNOR U7374 ( .A(n7116), .B(n7115), .Z(n7238) );
  NAND U7375 ( .A(x[79]), .B(y[260]), .Z(n7239) );
  XNOR U7376 ( .A(n7238), .B(n7239), .Z(n7205) );
  XNOR U7377 ( .A(n7206), .B(n7205), .Z(n7207) );
  XOR U7378 ( .A(n7208), .B(n7207), .Z(n7278) );
  AND U7379 ( .A(x[77]), .B(y[271]), .Z(n8482) );
  NANDN U7380 ( .A(n7117), .B(n8482), .Z(n7121) );
  NANDN U7381 ( .A(n7119), .B(n7118), .Z(n7120) );
  AND U7382 ( .A(n7121), .B(n7120), .Z(n7202) );
  AND U7383 ( .A(y[265]), .B(x[74]), .Z(n7123) );
  NAND U7384 ( .A(y[258]), .B(x[81]), .Z(n7122) );
  XNOR U7385 ( .A(n7123), .B(n7122), .Z(n7234) );
  NAND U7386 ( .A(x[82]), .B(y[257]), .Z(n7257) );
  XNOR U7387 ( .A(o[83]), .B(n7257), .Z(n7233) );
  XOR U7388 ( .A(n7234), .B(n7233), .Z(n7200) );
  AND U7389 ( .A(y[272]), .B(x[67]), .Z(n7125) );
  NAND U7390 ( .A(y[264]), .B(x[75]), .Z(n7124) );
  XNOR U7391 ( .A(n7125), .B(n7124), .Z(n7251) );
  XOR U7392 ( .A(n7200), .B(n7199), .Z(n7201) );
  XOR U7393 ( .A(n7202), .B(n7201), .Z(n7277) );
  NAND U7394 ( .A(n7518), .B(n7126), .Z(n7130) );
  NANDN U7395 ( .A(n7128), .B(n7127), .Z(n7129) );
  AND U7396 ( .A(n7130), .B(n7129), .Z(n7267) );
  ANDN U7397 ( .B(o[82]), .A(n7131), .Z(n7218) );
  AND U7398 ( .A(x[64]), .B(y[275]), .Z(n7215) );
  NAND U7399 ( .A(x[83]), .B(y[256]), .Z(n7216) );
  XNOR U7400 ( .A(n7215), .B(n7216), .Z(n7217) );
  XOR U7401 ( .A(n7218), .B(n7217), .Z(n7265) );
  AND U7402 ( .A(x[68]), .B(y[271]), .Z(n7386) );
  NAND U7403 ( .A(y[270]), .B(x[69]), .Z(n7132) );
  XOR U7404 ( .A(n7133), .B(n7132), .Z(n7212) );
  XNOR U7405 ( .A(n7386), .B(n7212), .Z(n7264) );
  XOR U7406 ( .A(n7265), .B(n7264), .Z(n7266) );
  XOR U7407 ( .A(n7267), .B(n7266), .Z(n7276) );
  XOR U7408 ( .A(n7277), .B(n7276), .Z(n7279) );
  XNOR U7409 ( .A(n7278), .B(n7279), .Z(n7272) );
  NAND U7410 ( .A(n7135), .B(n7134), .Z(n7139) );
  NANDN U7411 ( .A(n7137), .B(n7136), .Z(n7138) );
  AND U7412 ( .A(n7139), .B(n7138), .Z(n7271) );
  NAND U7413 ( .A(n7141), .B(n7140), .Z(n7145) );
  NANDN U7414 ( .A(n7143), .B(n7142), .Z(n7144) );
  NAND U7415 ( .A(n7145), .B(n7144), .Z(n7270) );
  XNOR U7416 ( .A(n7271), .B(n7270), .Z(n7273) );
  XNOR U7417 ( .A(n7272), .B(n7273), .Z(n7193) );
  XOR U7418 ( .A(n7194), .B(n7193), .Z(n7195) );
  XOR U7419 ( .A(n7196), .B(n7195), .Z(n7296) );
  NANDN U7420 ( .A(n7147), .B(n7146), .Z(n7151) );
  NANDN U7421 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U7422 ( .A(n7151), .B(n7150), .Z(n7295) );
  NANDN U7423 ( .A(n7153), .B(n7152), .Z(n7157) );
  NAND U7424 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7425 ( .A(n7157), .B(n7156), .Z(n7291) );
  NAND U7426 ( .A(n7159), .B(n7158), .Z(n7163) );
  NAND U7427 ( .A(n7161), .B(n7160), .Z(n7162) );
  AND U7428 ( .A(n7163), .B(n7162), .Z(n7289) );
  NANDN U7429 ( .A(n7165), .B(n7164), .Z(n7169) );
  NAND U7430 ( .A(n7167), .B(n7166), .Z(n7168) );
  NAND U7431 ( .A(n7169), .B(n7168), .Z(n7288) );
  XOR U7432 ( .A(n7295), .B(n7294), .Z(n7297) );
  XOR U7433 ( .A(n7296), .B(n7297), .Z(n7180) );
  XOR U7434 ( .A(n7181), .B(n7180), .Z(n7182) );
  XOR U7435 ( .A(n7183), .B(n7182), .Z(n7189) );
  NAND U7436 ( .A(n7174), .B(n7173), .Z(n7178) );
  NAND U7437 ( .A(n7176), .B(n7175), .Z(n7177) );
  NAND U7438 ( .A(n7178), .B(n7177), .Z(n7187) );
  IV U7439 ( .A(n7187), .Z(n7186) );
  XOR U7440 ( .A(n7188), .B(n7186), .Z(n7179) );
  XNOR U7441 ( .A(n7189), .B(n7179), .Z(N180) );
  NAND U7442 ( .A(n7181), .B(n7180), .Z(n7185) );
  NANDN U7443 ( .A(n7183), .B(n7182), .Z(n7184) );
  NAND U7444 ( .A(n7185), .B(n7184), .Z(n7308) );
  IV U7445 ( .A(n7308), .Z(n7307) );
  OR U7446 ( .A(n7188), .B(n7186), .Z(n7192) );
  ANDN U7447 ( .B(n7188), .A(n7187), .Z(n7190) );
  OR U7448 ( .A(n7190), .B(n7189), .Z(n7191) );
  AND U7449 ( .A(n7192), .B(n7191), .Z(n7309) );
  NAND U7450 ( .A(n7194), .B(n7193), .Z(n7198) );
  NANDN U7451 ( .A(n7196), .B(n7195), .Z(n7197) );
  AND U7452 ( .A(n7198), .B(n7197), .Z(n7418) );
  NAND U7453 ( .A(n7200), .B(n7199), .Z(n7204) );
  NANDN U7454 ( .A(n7202), .B(n7201), .Z(n7203) );
  AND U7455 ( .A(n7204), .B(n7203), .Z(n7410) );
  NANDN U7456 ( .A(n7206), .B(n7205), .Z(n7210) );
  NANDN U7457 ( .A(n7208), .B(n7207), .Z(n7209) );
  AND U7458 ( .A(n7210), .B(n7209), .Z(n7351) );
  AND U7459 ( .A(x[70]), .B(y[270]), .Z(n7337) );
  AND U7460 ( .A(x[69]), .B(y[269]), .Z(n7211) );
  NAND U7461 ( .A(n7337), .B(n7211), .Z(n7214) );
  NANDN U7462 ( .A(n7212), .B(n7386), .Z(n7213) );
  AND U7463 ( .A(n7214), .B(n7213), .Z(n7345) );
  NANDN U7464 ( .A(n7216), .B(n7215), .Z(n7220) );
  NAND U7465 ( .A(n7218), .B(n7217), .Z(n7219) );
  AND U7466 ( .A(n7220), .B(n7219), .Z(n7343) );
  AND U7467 ( .A(y[258]), .B(x[82]), .Z(n7222) );
  NAND U7468 ( .A(y[264]), .B(x[76]), .Z(n7221) );
  XNOR U7469 ( .A(n7222), .B(n7221), .Z(n7321) );
  NAND U7470 ( .A(x[81]), .B(y[259]), .Z(n7322) );
  XNOR U7471 ( .A(n7321), .B(n7322), .Z(n7342) );
  XNOR U7472 ( .A(n7343), .B(n7342), .Z(n7344) );
  XOR U7473 ( .A(n7345), .B(n7344), .Z(n7349) );
  AND U7474 ( .A(y[263]), .B(x[77]), .Z(n7224) );
  NAND U7475 ( .A(y[273]), .B(x[67]), .Z(n7223) );
  XNOR U7476 ( .A(n7224), .B(n7223), .Z(n7367) );
  XOR U7477 ( .A(n7367), .B(n7366), .Z(n7339) );
  AND U7478 ( .A(y[271]), .B(x[69]), .Z(n7226) );
  NAND U7479 ( .A(y[272]), .B(x[68]), .Z(n7225) );
  XNOR U7480 ( .A(n7226), .B(n7225), .Z(n7388) );
  AND U7481 ( .A(x[71]), .B(y[269]), .Z(n7387) );
  XNOR U7482 ( .A(n7388), .B(n7387), .Z(n7336) );
  XNOR U7483 ( .A(n7337), .B(n7336), .Z(n7338) );
  XOR U7484 ( .A(n7339), .B(n7338), .Z(n7393) );
  AND U7485 ( .A(x[72]), .B(y[274]), .Z(n8440) );
  AND U7486 ( .A(x[65]), .B(y[267]), .Z(n7227) );
  NAND U7487 ( .A(n8440), .B(n7227), .Z(n7231) );
  NANDN U7488 ( .A(n7229), .B(n7228), .Z(n7230) );
  AND U7489 ( .A(n7231), .B(n7230), .Z(n7392) );
  AND U7490 ( .A(x[81]), .B(y[265]), .Z(n8147) );
  NAND U7491 ( .A(n8147), .B(n7232), .Z(n7236) );
  NAND U7492 ( .A(n7234), .B(n7233), .Z(n7235) );
  NAND U7493 ( .A(n7236), .B(n7235), .Z(n7391) );
  XNOR U7494 ( .A(n7392), .B(n7391), .Z(n7394) );
  XNOR U7495 ( .A(n7393), .B(n7394), .Z(n7348) );
  XOR U7496 ( .A(n7349), .B(n7348), .Z(n7350) );
  XOR U7497 ( .A(n7351), .B(n7350), .Z(n7409) );
  XOR U7498 ( .A(n7410), .B(n7409), .Z(n7412) );
  AND U7499 ( .A(x[80]), .B(y[266]), .Z(n8141) );
  NAND U7500 ( .A(n8141), .B(n7237), .Z(n7241) );
  NANDN U7501 ( .A(n7239), .B(n7238), .Z(n7240) );
  AND U7502 ( .A(n7241), .B(n7240), .Z(n7355) );
  AND U7503 ( .A(x[77]), .B(y[273]), .Z(n8711) );
  NAND U7504 ( .A(n8711), .B(n7242), .Z(n7246) );
  NANDN U7505 ( .A(n7244), .B(n7243), .Z(n7245) );
  AND U7506 ( .A(n7246), .B(n7245), .Z(n7400) );
  NAND U7507 ( .A(y[260]), .B(x[80]), .Z(n7247) );
  XNOR U7508 ( .A(n7248), .B(n7247), .Z(n7361) );
  NAND U7509 ( .A(x[66]), .B(y[274]), .Z(n7362) );
  XNOR U7510 ( .A(n7361), .B(n7362), .Z(n7398) );
  NAND U7511 ( .A(y[261]), .B(x[79]), .Z(n7249) );
  XNOR U7512 ( .A(n7250), .B(n7249), .Z(n7331) );
  NAND U7513 ( .A(x[78]), .B(y[262]), .Z(n7332) );
  XNOR U7514 ( .A(n7331), .B(n7332), .Z(n7397) );
  XOR U7515 ( .A(n7398), .B(n7397), .Z(n7399) );
  XNOR U7516 ( .A(n7400), .B(n7399), .Z(n7354) );
  XNOR U7517 ( .A(n7355), .B(n7354), .Z(n7357) );
  NAND U7518 ( .A(x[75]), .B(y[272]), .Z(n8316) );
  NANDN U7519 ( .A(n8316), .B(n7497), .Z(n7254) );
  NANDN U7520 ( .A(n7252), .B(n7251), .Z(n7253) );
  AND U7521 ( .A(n7254), .B(n7253), .Z(n7406) );
  AND U7522 ( .A(y[265]), .B(x[75]), .Z(n7256) );
  NAND U7523 ( .A(y[275]), .B(x[65]), .Z(n7255) );
  XNOR U7524 ( .A(n7256), .B(n7255), .Z(n7327) );
  NAND U7525 ( .A(x[83]), .B(y[257]), .Z(n7335) );
  XNOR U7526 ( .A(o[84]), .B(n7335), .Z(n7326) );
  XOR U7527 ( .A(n7327), .B(n7326), .Z(n7404) );
  ANDN U7528 ( .B(o[83]), .A(n7257), .Z(n7383) );
  AND U7529 ( .A(x[64]), .B(y[276]), .Z(n7380) );
  NAND U7530 ( .A(x[84]), .B(y[256]), .Z(n7381) );
  XNOR U7531 ( .A(n7380), .B(n7381), .Z(n7382) );
  XOR U7532 ( .A(n7383), .B(n7382), .Z(n7403) );
  XOR U7533 ( .A(n7404), .B(n7403), .Z(n7405) );
  XNOR U7534 ( .A(n7406), .B(n7405), .Z(n7356) );
  XOR U7535 ( .A(n7357), .B(n7356), .Z(n7317) );
  NAND U7536 ( .A(n7259), .B(n7258), .Z(n7263) );
  NANDN U7537 ( .A(n7261), .B(n7260), .Z(n7262) );
  AND U7538 ( .A(n7263), .B(n7262), .Z(n7314) );
  NAND U7539 ( .A(n7265), .B(n7264), .Z(n7269) );
  NANDN U7540 ( .A(n7267), .B(n7266), .Z(n7268) );
  NAND U7541 ( .A(n7269), .B(n7268), .Z(n7315) );
  XNOR U7542 ( .A(n7314), .B(n7315), .Z(n7316) );
  XNOR U7543 ( .A(n7317), .B(n7316), .Z(n7411) );
  XOR U7544 ( .A(n7412), .B(n7411), .Z(n7416) );
  NANDN U7545 ( .A(n7271), .B(n7270), .Z(n7275) );
  NAND U7546 ( .A(n7273), .B(n7272), .Z(n7274) );
  AND U7547 ( .A(n7275), .B(n7274), .Z(n7424) );
  NAND U7548 ( .A(n7277), .B(n7276), .Z(n7281) );
  NAND U7549 ( .A(n7279), .B(n7278), .Z(n7280) );
  AND U7550 ( .A(n7281), .B(n7280), .Z(n7422) );
  NANDN U7551 ( .A(n7283), .B(n7282), .Z(n7287) );
  NANDN U7552 ( .A(n7285), .B(n7284), .Z(n7286) );
  AND U7553 ( .A(n7287), .B(n7286), .Z(n7421) );
  XNOR U7554 ( .A(n7424), .B(n7423), .Z(n7415) );
  XNOR U7555 ( .A(n7416), .B(n7415), .Z(n7417) );
  XOR U7556 ( .A(n7418), .B(n7417), .Z(n7304) );
  NANDN U7557 ( .A(n7289), .B(n7288), .Z(n7293) );
  NANDN U7558 ( .A(n7291), .B(n7290), .Z(n7292) );
  AND U7559 ( .A(n7293), .B(n7292), .Z(n7301) );
  NAND U7560 ( .A(n7295), .B(n7294), .Z(n7299) );
  NAND U7561 ( .A(n7297), .B(n7296), .Z(n7298) );
  NAND U7562 ( .A(n7299), .B(n7298), .Z(n7302) );
  XNOR U7563 ( .A(n7301), .B(n7302), .Z(n7303) );
  XNOR U7564 ( .A(n7304), .B(n7303), .Z(n7310) );
  XNOR U7565 ( .A(n7309), .B(n7310), .Z(n7300) );
  XOR U7566 ( .A(n7307), .B(n7300), .Z(N181) );
  NANDN U7567 ( .A(n7302), .B(n7301), .Z(n7306) );
  NANDN U7568 ( .A(n7304), .B(n7303), .Z(n7305) );
  NAND U7569 ( .A(n7306), .B(n7305), .Z(n7551) );
  IV U7570 ( .A(n7551), .Z(n7549) );
  OR U7571 ( .A(n7309), .B(n7307), .Z(n7313) );
  ANDN U7572 ( .B(n7309), .A(n7308), .Z(n7311) );
  OR U7573 ( .A(n7311), .B(n7310), .Z(n7312) );
  AND U7574 ( .A(n7313), .B(n7312), .Z(n7550) );
  NANDN U7575 ( .A(n7315), .B(n7314), .Z(n7319) );
  NANDN U7576 ( .A(n7317), .B(n7316), .Z(n7318) );
  AND U7577 ( .A(n7319), .B(n7318), .Z(n7437) );
  NAND U7578 ( .A(x[82]), .B(y[264]), .Z(n8150) );
  NANDN U7579 ( .A(n8150), .B(n7320), .Z(n7324) );
  NANDN U7580 ( .A(n7322), .B(n7321), .Z(n7323) );
  AND U7581 ( .A(n7324), .B(n7323), .Z(n7526) );
  AND U7582 ( .A(x[75]), .B(y[275]), .Z(n8924) );
  AND U7583 ( .A(x[65]), .B(y[265]), .Z(n7325) );
  NAND U7584 ( .A(n8924), .B(n7325), .Z(n7329) );
  NAND U7585 ( .A(n7327), .B(n7326), .Z(n7328) );
  NAND U7586 ( .A(n7329), .B(n7328), .Z(n7525) );
  XNOR U7587 ( .A(n7526), .B(n7525), .Z(n7528) );
  AND U7588 ( .A(x[79]), .B(y[267]), .Z(n8136) );
  NAND U7589 ( .A(n8136), .B(n7330), .Z(n7334) );
  NANDN U7590 ( .A(n7332), .B(n7331), .Z(n7333) );
  AND U7591 ( .A(n7334), .B(n7333), .Z(n7484) );
  ANDN U7592 ( .B(o[84]), .A(n7335), .Z(n7506) );
  AND U7593 ( .A(x[64]), .B(y[277]), .Z(n7503) );
  NAND U7594 ( .A(x[85]), .B(y[256]), .Z(n7504) );
  XNOR U7595 ( .A(n7503), .B(n7504), .Z(n7505) );
  XOR U7596 ( .A(n7506), .B(n7505), .Z(n7482) );
  AND U7597 ( .A(x[69]), .B(y[272]), .Z(n7488) );
  AND U7598 ( .A(x[80]), .B(y[261]), .Z(n7487) );
  XOR U7599 ( .A(n7488), .B(n7487), .Z(n7490) );
  NAND U7600 ( .A(x[79]), .B(y[262]), .Z(n7489) );
  XNOR U7601 ( .A(n7490), .B(n7489), .Z(n7481) );
  XOR U7602 ( .A(n7482), .B(n7481), .Z(n7483) );
  XNOR U7603 ( .A(n7484), .B(n7483), .Z(n7527) );
  XOR U7604 ( .A(n7528), .B(n7527), .Z(n7520) );
  NANDN U7605 ( .A(n7337), .B(n7336), .Z(n7341) );
  NANDN U7606 ( .A(n7339), .B(n7338), .Z(n7340) );
  NAND U7607 ( .A(n7341), .B(n7340), .Z(n7519) );
  XNOR U7608 ( .A(n7520), .B(n7519), .Z(n7522) );
  NANDN U7609 ( .A(n7343), .B(n7342), .Z(n7347) );
  NANDN U7610 ( .A(n7345), .B(n7344), .Z(n7346) );
  AND U7611 ( .A(n7347), .B(n7346), .Z(n7521) );
  XOR U7612 ( .A(n7522), .B(n7521), .Z(n7435) );
  NAND U7613 ( .A(n7349), .B(n7348), .Z(n7353) );
  NAND U7614 ( .A(n7351), .B(n7350), .Z(n7352) );
  AND U7615 ( .A(n7353), .B(n7352), .Z(n7434) );
  XNOR U7616 ( .A(n7435), .B(n7434), .Z(n7436) );
  XOR U7617 ( .A(n7437), .B(n7436), .Z(n7431) );
  NANDN U7618 ( .A(n7355), .B(n7354), .Z(n7359) );
  NAND U7619 ( .A(n7357), .B(n7356), .Z(n7358) );
  AND U7620 ( .A(n7359), .B(n7358), .Z(n7443) );
  NAND U7621 ( .A(n8141), .B(n7360), .Z(n7364) );
  NANDN U7622 ( .A(n7362), .B(n7361), .Z(n7363) );
  AND U7623 ( .A(n7364), .B(n7363), .Z(n7453) );
  NAND U7624 ( .A(n7365), .B(n8711), .Z(n7369) );
  NAND U7625 ( .A(n7367), .B(n7366), .Z(n7368) );
  AND U7626 ( .A(n7369), .B(n7368), .Z(n7540) );
  AND U7627 ( .A(y[258]), .B(x[83]), .Z(n7371) );
  NAND U7628 ( .A(y[266]), .B(x[75]), .Z(n7370) );
  XNOR U7629 ( .A(n7371), .B(n7370), .Z(n7472) );
  NAND U7630 ( .A(x[84]), .B(y[257]), .Z(n7502) );
  XNOR U7631 ( .A(o[85]), .B(n7502), .Z(n7471) );
  XOR U7632 ( .A(n7472), .B(n7471), .Z(n7538) );
  NAND U7633 ( .A(y[259]), .B(x[82]), .Z(n7372) );
  XNOR U7634 ( .A(n7373), .B(n7372), .Z(n7510) );
  NAND U7635 ( .A(x[65]), .B(y[276]), .Z(n7511) );
  XNOR U7636 ( .A(n7510), .B(n7511), .Z(n7537) );
  XOR U7637 ( .A(n7538), .B(n7537), .Z(n7539) );
  XNOR U7638 ( .A(n7540), .B(n7539), .Z(n7452) );
  XNOR U7639 ( .A(n7453), .B(n7452), .Z(n7455) );
  AND U7640 ( .A(x[71]), .B(y[270]), .Z(n7704) );
  AND U7641 ( .A(y[271]), .B(x[70]), .Z(n7375) );
  NAND U7642 ( .A(y[263]), .B(x[78]), .Z(n7374) );
  XNOR U7643 ( .A(n7375), .B(n7374), .Z(n7514) );
  XOR U7644 ( .A(n7704), .B(n7514), .Z(n7461) );
  AND U7645 ( .A(x[73]), .B(y[268]), .Z(n7459) );
  NAND U7646 ( .A(x[72]), .B(y[269]), .Z(n7458) );
  XNOR U7647 ( .A(n7459), .B(n7458), .Z(n7460) );
  XOR U7648 ( .A(n7461), .B(n7460), .Z(n7477) );
  AND U7649 ( .A(y[265]), .B(x[76]), .Z(n7377) );
  NAND U7650 ( .A(y[260]), .B(x[81]), .Z(n7376) );
  XNOR U7651 ( .A(n7377), .B(n7376), .Z(n7464) );
  NAND U7652 ( .A(x[66]), .B(y[275]), .Z(n7465) );
  XNOR U7653 ( .A(n7464), .B(n7465), .Z(n7476) );
  AND U7654 ( .A(y[264]), .B(x[77]), .Z(n7379) );
  NAND U7655 ( .A(y[274]), .B(x[67]), .Z(n7378) );
  XNOR U7656 ( .A(n7379), .B(n7378), .Z(n7498) );
  NAND U7657 ( .A(x[68]), .B(y[273]), .Z(n7499) );
  XNOR U7658 ( .A(n7498), .B(n7499), .Z(n7475) );
  XOR U7659 ( .A(n7476), .B(n7475), .Z(n7478) );
  XOR U7660 ( .A(n7477), .B(n7478), .Z(n7534) );
  NANDN U7661 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U7662 ( .A(n7383), .B(n7382), .Z(n7384) );
  AND U7663 ( .A(n7385), .B(n7384), .Z(n7532) );
  NAND U7664 ( .A(n7488), .B(n7386), .Z(n7390) );
  NAND U7665 ( .A(n7388), .B(n7387), .Z(n7389) );
  NAND U7666 ( .A(n7390), .B(n7389), .Z(n7531) );
  XNOR U7667 ( .A(n7532), .B(n7531), .Z(n7533) );
  XOR U7668 ( .A(n7534), .B(n7533), .Z(n7454) );
  XOR U7669 ( .A(n7455), .B(n7454), .Z(n7441) );
  NANDN U7670 ( .A(n7392), .B(n7391), .Z(n7396) );
  NAND U7671 ( .A(n7394), .B(n7393), .Z(n7395) );
  NAND U7672 ( .A(n7396), .B(n7395), .Z(n7448) );
  NAND U7673 ( .A(n7398), .B(n7397), .Z(n7402) );
  NANDN U7674 ( .A(n7400), .B(n7399), .Z(n7401) );
  NAND U7675 ( .A(n7402), .B(n7401), .Z(n7447) );
  NAND U7676 ( .A(n7404), .B(n7403), .Z(n7408) );
  NANDN U7677 ( .A(n7406), .B(n7405), .Z(n7407) );
  NAND U7678 ( .A(n7408), .B(n7407), .Z(n7446) );
  XOR U7679 ( .A(n7447), .B(n7446), .Z(n7449) );
  XOR U7680 ( .A(n7448), .B(n7449), .Z(n7440) );
  XOR U7681 ( .A(n7441), .B(n7440), .Z(n7442) );
  XOR U7682 ( .A(n7443), .B(n7442), .Z(n7429) );
  NAND U7683 ( .A(n7410), .B(n7409), .Z(n7414) );
  NAND U7684 ( .A(n7412), .B(n7411), .Z(n7413) );
  NAND U7685 ( .A(n7414), .B(n7413), .Z(n7428) );
  XOR U7686 ( .A(n7429), .B(n7428), .Z(n7430) );
  XOR U7687 ( .A(n7431), .B(n7430), .Z(n7545) );
  NANDN U7688 ( .A(n7416), .B(n7415), .Z(n7420) );
  NAND U7689 ( .A(n7418), .B(n7417), .Z(n7419) );
  AND U7690 ( .A(n7420), .B(n7419), .Z(n7544) );
  NANDN U7691 ( .A(n7422), .B(n7421), .Z(n7426) );
  NAND U7692 ( .A(n7424), .B(n7423), .Z(n7425) );
  AND U7693 ( .A(n7426), .B(n7425), .Z(n7543) );
  XNOR U7694 ( .A(n7544), .B(n7543), .Z(n7546) );
  XOR U7695 ( .A(n7545), .B(n7546), .Z(n7552) );
  XNOR U7696 ( .A(n7550), .B(n7552), .Z(n7427) );
  XOR U7697 ( .A(n7549), .B(n7427), .Z(N182) );
  NAND U7698 ( .A(n7429), .B(n7428), .Z(n7433) );
  NANDN U7699 ( .A(n7431), .B(n7430), .Z(n7432) );
  AND U7700 ( .A(n7433), .B(n7432), .Z(n7681) );
  NANDN U7701 ( .A(n7435), .B(n7434), .Z(n7439) );
  NAND U7702 ( .A(n7437), .B(n7436), .Z(n7438) );
  AND U7703 ( .A(n7439), .B(n7438), .Z(n7679) );
  NAND U7704 ( .A(n7441), .B(n7440), .Z(n7445) );
  NANDN U7705 ( .A(n7443), .B(n7442), .Z(n7444) );
  AND U7706 ( .A(n7445), .B(n7444), .Z(n7558) );
  NAND U7707 ( .A(n7447), .B(n7446), .Z(n7451) );
  NAND U7708 ( .A(n7449), .B(n7448), .Z(n7450) );
  NAND U7709 ( .A(n7451), .B(n7450), .Z(n7557) );
  XNOR U7710 ( .A(n7558), .B(n7557), .Z(n7560) );
  NANDN U7711 ( .A(n7453), .B(n7452), .Z(n7457) );
  NAND U7712 ( .A(n7455), .B(n7454), .Z(n7456) );
  AND U7713 ( .A(n7457), .B(n7456), .Z(n7666) );
  NANDN U7714 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U7715 ( .A(n7461), .B(n7460), .Z(n7462) );
  AND U7716 ( .A(n7463), .B(n7462), .Z(n7660) );
  NAND U7717 ( .A(n8147), .B(n7612), .Z(n7467) );
  NANDN U7718 ( .A(n7465), .B(n7464), .Z(n7466) );
  NAND U7719 ( .A(n7467), .B(n7466), .Z(n7589) );
  AND U7720 ( .A(x[69]), .B(y[273]), .Z(n7633) );
  NAND U7721 ( .A(x[81]), .B(y[261]), .Z(n7634) );
  XNOR U7722 ( .A(n7633), .B(n7634), .Z(n7635) );
  NAND U7723 ( .A(x[80]), .B(y[262]), .Z(n7636) );
  XNOR U7724 ( .A(n7635), .B(n7636), .Z(n7588) );
  AND U7725 ( .A(y[260]), .B(x[82]), .Z(n7469) );
  NAND U7726 ( .A(y[266]), .B(x[76]), .Z(n7468) );
  XNOR U7727 ( .A(n7469), .B(n7468), .Z(n7613) );
  NAND U7728 ( .A(x[68]), .B(y[274]), .Z(n7614) );
  XNOR U7729 ( .A(n7613), .B(n7614), .Z(n7587) );
  XOR U7730 ( .A(n7588), .B(n7587), .Z(n7590) );
  XNOR U7731 ( .A(n7589), .B(n7590), .Z(n7657) );
  AND U7732 ( .A(x[83]), .B(y[266]), .Z(n8609) );
  NAND U7733 ( .A(n7470), .B(n8609), .Z(n7474) );
  NAND U7734 ( .A(n7472), .B(n7471), .Z(n7473) );
  AND U7735 ( .A(n7474), .B(n7473), .Z(n7658) );
  XOR U7736 ( .A(n7657), .B(n7658), .Z(n7659) );
  XOR U7737 ( .A(n7660), .B(n7659), .Z(n7663) );
  NAND U7738 ( .A(n7476), .B(n7475), .Z(n7480) );
  NAND U7739 ( .A(n7478), .B(n7477), .Z(n7479) );
  AND U7740 ( .A(n7480), .B(n7479), .Z(n7646) );
  NAND U7741 ( .A(n7482), .B(n7481), .Z(n7486) );
  NANDN U7742 ( .A(n7484), .B(n7483), .Z(n7485) );
  NAND U7743 ( .A(n7486), .B(n7485), .Z(n7645) );
  XNOR U7744 ( .A(n7646), .B(n7645), .Z(n7648) );
  NAND U7745 ( .A(n7488), .B(n7487), .Z(n7492) );
  ANDN U7746 ( .B(n7490), .A(n7489), .Z(n7491) );
  ANDN U7747 ( .B(n7492), .A(n7491), .Z(n7609) );
  AND U7748 ( .A(y[258]), .B(x[84]), .Z(n7494) );
  NAND U7749 ( .A(y[265]), .B(x[77]), .Z(n7493) );
  XNOR U7750 ( .A(n7494), .B(n7493), .Z(n7629) );
  NAND U7751 ( .A(x[66]), .B(y[276]), .Z(n7630) );
  XNOR U7752 ( .A(n7629), .B(n7630), .Z(n7607) );
  AND U7753 ( .A(y[263]), .B(x[79]), .Z(n7496) );
  NAND U7754 ( .A(y[272]), .B(x[70]), .Z(n7495) );
  XNOR U7755 ( .A(n7496), .B(n7495), .Z(n7641) );
  XOR U7756 ( .A(n7607), .B(n7606), .Z(n7608) );
  XNOR U7757 ( .A(n7609), .B(n7608), .Z(n7652) );
  AND U7758 ( .A(x[77]), .B(y[274]), .Z(n8922) );
  NAND U7759 ( .A(n7497), .B(n8922), .Z(n7501) );
  NANDN U7760 ( .A(n7499), .B(n7498), .Z(n7500) );
  AND U7761 ( .A(n7501), .B(n7500), .Z(n7578) );
  AND U7762 ( .A(x[65]), .B(y[277]), .Z(n7601) );
  XOR U7763 ( .A(n7602), .B(n7601), .Z(n7600) );
  ANDN U7764 ( .B(o[85]), .A(n7502), .Z(n7599) );
  XOR U7765 ( .A(n7600), .B(n7599), .Z(n7576) );
  AND U7766 ( .A(x[78]), .B(y[264]), .Z(n7593) );
  NAND U7767 ( .A(x[67]), .B(y[275]), .Z(n7594) );
  XNOR U7768 ( .A(n7593), .B(n7594), .Z(n7595) );
  NAND U7769 ( .A(x[83]), .B(y[259]), .Z(n7596) );
  XNOR U7770 ( .A(n7595), .B(n7596), .Z(n7575) );
  XOR U7771 ( .A(n7576), .B(n7575), .Z(n7577) );
  XNOR U7772 ( .A(n7578), .B(n7577), .Z(n7651) );
  XOR U7773 ( .A(n7652), .B(n7651), .Z(n7654) );
  NANDN U7774 ( .A(n7504), .B(n7503), .Z(n7508) );
  NAND U7775 ( .A(n7506), .B(n7505), .Z(n7507) );
  AND U7776 ( .A(n7508), .B(n7507), .Z(n7570) );
  AND U7777 ( .A(x[82]), .B(y[267]), .Z(n8611) );
  NAND U7778 ( .A(n8611), .B(n7509), .Z(n7513) );
  NANDN U7779 ( .A(n7511), .B(n7510), .Z(n7512) );
  NAND U7780 ( .A(n7513), .B(n7512), .Z(n7569) );
  XNOR U7781 ( .A(n7570), .B(n7569), .Z(n7572) );
  AND U7782 ( .A(x[78]), .B(y[271]), .Z(n8621) );
  NAND U7783 ( .A(n7640), .B(n8621), .Z(n7516) );
  NAND U7784 ( .A(n7704), .B(n7514), .Z(n7515) );
  AND U7785 ( .A(n7516), .B(n7515), .Z(n7584) );
  AND U7786 ( .A(x[64]), .B(y[278]), .Z(n7617) );
  NAND U7787 ( .A(x[86]), .B(y[256]), .Z(n7618) );
  XNOR U7788 ( .A(n7617), .B(n7618), .Z(n7620) );
  NAND U7789 ( .A(x[85]), .B(y[257]), .Z(n7639) );
  XNOR U7790 ( .A(o[86]), .B(n7639), .Z(n7619) );
  XOR U7791 ( .A(n7620), .B(n7619), .Z(n7582) );
  NAND U7792 ( .A(y[271]), .B(x[71]), .Z(n7517) );
  XNOR U7793 ( .A(n7518), .B(n7517), .Z(n7623) );
  XOR U7794 ( .A(n7582), .B(n7581), .Z(n7583) );
  XNOR U7795 ( .A(n7584), .B(n7583), .Z(n7571) );
  XOR U7796 ( .A(n7572), .B(n7571), .Z(n7653) );
  XOR U7797 ( .A(n7654), .B(n7653), .Z(n7647) );
  XOR U7798 ( .A(n7648), .B(n7647), .Z(n7664) );
  XOR U7799 ( .A(n7663), .B(n7664), .Z(n7665) );
  XNOR U7800 ( .A(n7666), .B(n7665), .Z(n7672) );
  NANDN U7801 ( .A(n7520), .B(n7519), .Z(n7524) );
  NAND U7802 ( .A(n7522), .B(n7521), .Z(n7523) );
  AND U7803 ( .A(n7524), .B(n7523), .Z(n7670) );
  NANDN U7804 ( .A(n7526), .B(n7525), .Z(n7530) );
  NAND U7805 ( .A(n7528), .B(n7527), .Z(n7529) );
  AND U7806 ( .A(n7530), .B(n7529), .Z(n7566) );
  NANDN U7807 ( .A(n7532), .B(n7531), .Z(n7536) );
  NAND U7808 ( .A(n7534), .B(n7533), .Z(n7535) );
  AND U7809 ( .A(n7536), .B(n7535), .Z(n7564) );
  NAND U7810 ( .A(n7538), .B(n7537), .Z(n7542) );
  NANDN U7811 ( .A(n7540), .B(n7539), .Z(n7541) );
  NAND U7812 ( .A(n7542), .B(n7541), .Z(n7563) );
  XNOR U7813 ( .A(n7564), .B(n7563), .Z(n7565) );
  XNOR U7814 ( .A(n7566), .B(n7565), .Z(n7669) );
  XOR U7815 ( .A(n7670), .B(n7669), .Z(n7671) );
  XOR U7816 ( .A(n7672), .B(n7671), .Z(n7559) );
  XOR U7817 ( .A(n7560), .B(n7559), .Z(n7678) );
  XNOR U7818 ( .A(n7679), .B(n7678), .Z(n7680) );
  XNOR U7819 ( .A(n7681), .B(n7680), .Z(n7677) );
  NANDN U7820 ( .A(n7544), .B(n7543), .Z(n7548) );
  NAND U7821 ( .A(n7546), .B(n7545), .Z(n7547) );
  NAND U7822 ( .A(n7548), .B(n7547), .Z(n7676) );
  NANDN U7823 ( .A(n7549), .B(n7550), .Z(n7555) );
  NOR U7824 ( .A(n7551), .B(n7550), .Z(n7553) );
  OR U7825 ( .A(n7553), .B(n7552), .Z(n7554) );
  AND U7826 ( .A(n7555), .B(n7554), .Z(n7675) );
  XOR U7827 ( .A(n7676), .B(n7675), .Z(n7556) );
  XNOR U7828 ( .A(n7677), .B(n7556), .Z(N183) );
  NANDN U7829 ( .A(n7558), .B(n7557), .Z(n7562) );
  NAND U7830 ( .A(n7560), .B(n7559), .Z(n7561) );
  AND U7831 ( .A(n7562), .B(n7561), .Z(n7825) );
  NANDN U7832 ( .A(n7564), .B(n7563), .Z(n7568) );
  NANDN U7833 ( .A(n7566), .B(n7565), .Z(n7567) );
  AND U7834 ( .A(n7568), .B(n7567), .Z(n7800) );
  NANDN U7835 ( .A(n7570), .B(n7569), .Z(n7574) );
  NAND U7836 ( .A(n7572), .B(n7571), .Z(n7573) );
  AND U7837 ( .A(n7574), .B(n7573), .Z(n7794) );
  NAND U7838 ( .A(n7576), .B(n7575), .Z(n7580) );
  NANDN U7839 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U7840 ( .A(n7580), .B(n7579), .Z(n7792) );
  NAND U7841 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U7842 ( .A(n7584), .B(n7583), .Z(n7585) );
  NAND U7843 ( .A(n7586), .B(n7585), .Z(n7791) );
  XNOR U7844 ( .A(n7792), .B(n7791), .Z(n7793) );
  XNOR U7845 ( .A(n7794), .B(n7793), .Z(n7812) );
  NAND U7846 ( .A(n7588), .B(n7587), .Z(n7592) );
  NAND U7847 ( .A(n7590), .B(n7589), .Z(n7591) );
  AND U7848 ( .A(n7592), .B(n7591), .Z(n7810) );
  NANDN U7849 ( .A(n7594), .B(n7593), .Z(n7598) );
  NANDN U7850 ( .A(n7596), .B(n7595), .Z(n7597) );
  AND U7851 ( .A(n7598), .B(n7597), .Z(n7738) );
  AND U7852 ( .A(n7600), .B(n7599), .Z(n7604) );
  NAND U7853 ( .A(n7602), .B(n7601), .Z(n7603) );
  NANDN U7854 ( .A(n7604), .B(n7603), .Z(n7737) );
  XNOR U7855 ( .A(n7738), .B(n7737), .Z(n7740) );
  NAND U7856 ( .A(y[272]), .B(x[71]), .Z(n7605) );
  XNOR U7857 ( .A(n7888), .B(n7605), .Z(n7705) );
  NAND U7858 ( .A(x[74]), .B(y[269]), .Z(n7744) );
  XNOR U7859 ( .A(n7743), .B(n7744), .Z(n7746) );
  AND U7860 ( .A(x[70]), .B(y[273]), .Z(n7696) );
  NAND U7861 ( .A(x[79]), .B(y[264]), .Z(n7697) );
  XNOR U7862 ( .A(n7696), .B(n7697), .Z(n7698) );
  NAND U7863 ( .A(x[75]), .B(y[268]), .Z(n7699) );
  XNOR U7864 ( .A(n7698), .B(n7699), .Z(n7745) );
  XOR U7865 ( .A(n7746), .B(n7745), .Z(n7739) );
  XOR U7866 ( .A(n7740), .B(n7739), .Z(n7809) );
  XNOR U7867 ( .A(n7810), .B(n7809), .Z(n7811) );
  XOR U7868 ( .A(n7812), .B(n7811), .Z(n7798) );
  NAND U7869 ( .A(n7607), .B(n7606), .Z(n7611) );
  NANDN U7870 ( .A(n7609), .B(n7608), .Z(n7610) );
  AND U7871 ( .A(n7611), .B(n7610), .Z(n7732) );
  AND U7872 ( .A(x[82]), .B(y[266]), .Z(n8470) );
  NAND U7873 ( .A(n8470), .B(n7612), .Z(n7616) );
  NANDN U7874 ( .A(n7614), .B(n7613), .Z(n7615) );
  AND U7875 ( .A(n7616), .B(n7615), .Z(n7768) );
  NANDN U7876 ( .A(n7618), .B(n7617), .Z(n7622) );
  NAND U7877 ( .A(n7620), .B(n7619), .Z(n7621) );
  NAND U7878 ( .A(n7622), .B(n7621), .Z(n7767) );
  XNOR U7879 ( .A(n7768), .B(n7767), .Z(n7770) );
  NANDN U7880 ( .A(n7706), .B(n7704), .Z(n7626) );
  NANDN U7881 ( .A(n7624), .B(n7623), .Z(n7625) );
  AND U7882 ( .A(n7626), .B(n7625), .Z(n7782) );
  AND U7883 ( .A(x[64]), .B(y[279]), .Z(n7715) );
  NAND U7884 ( .A(x[87]), .B(y[256]), .Z(n7716) );
  XNOR U7885 ( .A(n7715), .B(n7716), .Z(n7718) );
  NAND U7886 ( .A(x[86]), .B(y[257]), .Z(n7695) );
  XNOR U7887 ( .A(o[87]), .B(n7695), .Z(n7717) );
  XOR U7888 ( .A(n7718), .B(n7717), .Z(n7780) );
  AND U7889 ( .A(y[259]), .B(x[84]), .Z(n8349) );
  NAND U7890 ( .A(y[263]), .B(x[80]), .Z(n7627) );
  XNOR U7891 ( .A(n8349), .B(n7627), .Z(n7691) );
  NAND U7892 ( .A(x[83]), .B(y[260]), .Z(n7692) );
  XNOR U7893 ( .A(n7691), .B(n7692), .Z(n7779) );
  XOR U7894 ( .A(n7780), .B(n7779), .Z(n7781) );
  XOR U7895 ( .A(n7770), .B(n7769), .Z(n7731) );
  XNOR U7896 ( .A(n7732), .B(n7731), .Z(n7734) );
  AND U7897 ( .A(x[84]), .B(y[265]), .Z(n8633) );
  NAND U7898 ( .A(n8633), .B(n7628), .Z(n7632) );
  NANDN U7899 ( .A(n7630), .B(n7629), .Z(n7631) );
  AND U7900 ( .A(n7632), .B(n7631), .Z(n7726) );
  NANDN U7901 ( .A(n7634), .B(n7633), .Z(n7638) );
  NANDN U7902 ( .A(n7636), .B(n7635), .Z(n7637) );
  AND U7903 ( .A(n7638), .B(n7637), .Z(n7788) );
  AND U7904 ( .A(x[77]), .B(y[266]), .Z(n7761) );
  NAND U7905 ( .A(x[66]), .B(y[277]), .Z(n7762) );
  XNOR U7906 ( .A(n7761), .B(n7762), .Z(n7763) );
  NAND U7907 ( .A(x[85]), .B(y[258]), .Z(n7764) );
  XNOR U7908 ( .A(n7763), .B(n7764), .Z(n7786) );
  AND U7909 ( .A(x[76]), .B(y[267]), .Z(n7709) );
  NAND U7910 ( .A(x[65]), .B(y[278]), .Z(n7710) );
  XNOR U7911 ( .A(n7709), .B(n7710), .Z(n7712) );
  ANDN U7912 ( .B(o[86]), .A(n7639), .Z(n7711) );
  XOR U7913 ( .A(n7712), .B(n7711), .Z(n7785) );
  XOR U7914 ( .A(n7786), .B(n7785), .Z(n7787) );
  XNOR U7915 ( .A(n7788), .B(n7787), .Z(n7725) );
  XNOR U7916 ( .A(n7726), .B(n7725), .Z(n7728) );
  AND U7917 ( .A(x[79]), .B(y[272]), .Z(n8871) );
  NAND U7918 ( .A(n8871), .B(n7640), .Z(n7644) );
  NANDN U7919 ( .A(n7642), .B(n7641), .Z(n7643) );
  AND U7920 ( .A(n7644), .B(n7643), .Z(n7776) );
  AND U7921 ( .A(x[78]), .B(y[265]), .Z(n7755) );
  NAND U7922 ( .A(x[67]), .B(y[276]), .Z(n7756) );
  XNOR U7923 ( .A(n7755), .B(n7756), .Z(n7757) );
  NAND U7924 ( .A(x[68]), .B(y[275]), .Z(n7758) );
  XNOR U7925 ( .A(n7757), .B(n7758), .Z(n7774) );
  AND U7926 ( .A(x[69]), .B(y[274]), .Z(n7749) );
  NAND U7927 ( .A(x[82]), .B(y[261]), .Z(n7750) );
  XNOR U7928 ( .A(n7749), .B(n7750), .Z(n7751) );
  NAND U7929 ( .A(x[81]), .B(y[262]), .Z(n7752) );
  XNOR U7930 ( .A(n7751), .B(n7752), .Z(n7773) );
  XOR U7931 ( .A(n7774), .B(n7773), .Z(n7775) );
  XNOR U7932 ( .A(n7776), .B(n7775), .Z(n7727) );
  XOR U7933 ( .A(n7728), .B(n7727), .Z(n7733) );
  XOR U7934 ( .A(n7734), .B(n7733), .Z(n7797) );
  XOR U7935 ( .A(n7798), .B(n7797), .Z(n7799) );
  XOR U7936 ( .A(n7800), .B(n7799), .Z(n7687) );
  NANDN U7937 ( .A(n7646), .B(n7645), .Z(n7650) );
  NAND U7938 ( .A(n7648), .B(n7647), .Z(n7649) );
  AND U7939 ( .A(n7650), .B(n7649), .Z(n7806) );
  NAND U7940 ( .A(n7652), .B(n7651), .Z(n7656) );
  NAND U7941 ( .A(n7654), .B(n7653), .Z(n7655) );
  AND U7942 ( .A(n7656), .B(n7655), .Z(n7804) );
  NAND U7943 ( .A(n7658), .B(n7657), .Z(n7662) );
  NANDN U7944 ( .A(n7660), .B(n7659), .Z(n7661) );
  AND U7945 ( .A(n7662), .B(n7661), .Z(n7803) );
  XNOR U7946 ( .A(n7804), .B(n7803), .Z(n7805) );
  XOR U7947 ( .A(n7806), .B(n7805), .Z(n7685) );
  NAND U7948 ( .A(n7664), .B(n7663), .Z(n7668) );
  NANDN U7949 ( .A(n7666), .B(n7665), .Z(n7667) );
  AND U7950 ( .A(n7668), .B(n7667), .Z(n7686) );
  XOR U7951 ( .A(n7685), .B(n7686), .Z(n7688) );
  XOR U7952 ( .A(n7687), .B(n7688), .Z(n7822) );
  NAND U7953 ( .A(n7670), .B(n7669), .Z(n7674) );
  NAND U7954 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U7955 ( .A(n7674), .B(n7673), .Z(n7823) );
  XNOR U7956 ( .A(n7822), .B(n7823), .Z(n7824) );
  XNOR U7957 ( .A(n7825), .B(n7824), .Z(n7818) );
  NANDN U7958 ( .A(n7679), .B(n7678), .Z(n7683) );
  NAND U7959 ( .A(n7681), .B(n7680), .Z(n7682) );
  AND U7960 ( .A(n7683), .B(n7682), .Z(n7817) );
  IV U7961 ( .A(n7817), .Z(n7815) );
  XOR U7962 ( .A(n7816), .B(n7815), .Z(n7684) );
  XNOR U7963 ( .A(n7818), .B(n7684), .Z(N184) );
  NAND U7964 ( .A(n7686), .B(n7685), .Z(n7690) );
  NAND U7965 ( .A(n7688), .B(n7687), .Z(n7689) );
  AND U7966 ( .A(n7690), .B(n7689), .Z(n7965) );
  AND U7967 ( .A(x[84]), .B(y[263]), .Z(n8223) );
  AND U7968 ( .A(x[80]), .B(y[259]), .Z(n7853) );
  NAND U7969 ( .A(n8223), .B(n7853), .Z(n7694) );
  NANDN U7970 ( .A(n7692), .B(n7691), .Z(n7693) );
  AND U7971 ( .A(n7694), .B(n7693), .Z(n7879) );
  AND U7972 ( .A(x[86]), .B(y[258]), .Z(n7898) );
  XOR U7973 ( .A(n7899), .B(n7898), .Z(n7900) );
  NAND U7974 ( .A(x[66]), .B(y[278]), .Z(n7901) );
  XNOR U7975 ( .A(n7900), .B(n7901), .Z(n7877) );
  AND U7976 ( .A(x[65]), .B(y[279]), .Z(n7906) );
  XOR U7977 ( .A(n7907), .B(n7906), .Z(n7905) );
  ANDN U7978 ( .B(o[87]), .A(n7695), .Z(n7904) );
  XOR U7979 ( .A(n7905), .B(n7904), .Z(n7876) );
  XOR U7980 ( .A(n7877), .B(n7876), .Z(n7878) );
  XNOR U7981 ( .A(n7879), .B(n7878), .Z(n7936) );
  NANDN U7982 ( .A(n7697), .B(n7696), .Z(n7701) );
  NANDN U7983 ( .A(n7699), .B(n7698), .Z(n7700) );
  AND U7984 ( .A(n7701), .B(n7700), .Z(n7873) );
  AND U7985 ( .A(y[259]), .B(x[85]), .Z(n7703) );
  NAND U7986 ( .A(y[264]), .B(x[80]), .Z(n7702) );
  XNOR U7987 ( .A(n7703), .B(n7702), .Z(n7854) );
  NAND U7988 ( .A(x[69]), .B(y[275]), .Z(n7855) );
  XNOR U7989 ( .A(n7854), .B(n7855), .Z(n7871) );
  AND U7990 ( .A(x[70]), .B(y[274]), .Z(n8236) );
  NAND U7991 ( .A(x[84]), .B(y[260]), .Z(n8057) );
  NAND U7992 ( .A(x[83]), .B(y[261]), .Z(n7861) );
  XNOR U7993 ( .A(n7860), .B(n7861), .Z(n7870) );
  XOR U7994 ( .A(n7871), .B(n7870), .Z(n7872) );
  XNOR U7995 ( .A(n7873), .B(n7872), .Z(n7850) );
  NANDN U7996 ( .A(n7991), .B(n7704), .Z(n7708) );
  NANDN U7997 ( .A(n7706), .B(n7705), .Z(n7707) );
  AND U7998 ( .A(n7708), .B(n7707), .Z(n7848) );
  NANDN U7999 ( .A(n7710), .B(n7709), .Z(n7714) );
  NAND U8000 ( .A(n7712), .B(n7711), .Z(n7713) );
  NAND U8001 ( .A(n7714), .B(n7713), .Z(n7847) );
  XNOR U8002 ( .A(n7848), .B(n7847), .Z(n7849) );
  XOR U8003 ( .A(n7850), .B(n7849), .Z(n7935) );
  XOR U8004 ( .A(n7936), .B(n7935), .Z(n7938) );
  NANDN U8005 ( .A(n7716), .B(n7715), .Z(n7720) );
  NAND U8006 ( .A(n7718), .B(n7717), .Z(n7719) );
  AND U8007 ( .A(n7720), .B(n7719), .Z(n7930) );
  AND U8008 ( .A(x[67]), .B(y[277]), .Z(n7917) );
  XOR U8009 ( .A(n7918), .B(n7917), .Z(n7920) );
  NAND U8010 ( .A(x[68]), .B(y[276]), .Z(n7919) );
  XNOR U8011 ( .A(n7920), .B(n7919), .Z(n7929) );
  XNOR U8012 ( .A(n7930), .B(n7929), .Z(n7932) );
  AND U8013 ( .A(y[270]), .B(x[74]), .Z(n7722) );
  NAND U8014 ( .A(y[271]), .B(x[73]), .Z(n7721) );
  XNOR U8015 ( .A(n7722), .B(n7721), .Z(n7890) );
  AND U8016 ( .A(y[272]), .B(x[72]), .Z(n7724) );
  NAND U8017 ( .A(y[266]), .B(x[78]), .Z(n7723) );
  XNOR U8018 ( .A(n7724), .B(n7723), .Z(n7894) );
  NAND U8019 ( .A(x[75]), .B(y[269]), .Z(n7895) );
  XOR U8020 ( .A(n7890), .B(n7889), .Z(n7931) );
  XOR U8021 ( .A(n7932), .B(n7931), .Z(n7937) );
  XOR U8022 ( .A(n7938), .B(n7937), .Z(n7948) );
  NANDN U8023 ( .A(n7726), .B(n7725), .Z(n7730) );
  NAND U8024 ( .A(n7728), .B(n7727), .Z(n7729) );
  AND U8025 ( .A(n7730), .B(n7729), .Z(n7947) );
  XNOR U8026 ( .A(n7948), .B(n7947), .Z(n7949) );
  NANDN U8027 ( .A(n7732), .B(n7731), .Z(n7736) );
  NAND U8028 ( .A(n7734), .B(n7733), .Z(n7735) );
  NAND U8029 ( .A(n7736), .B(n7735), .Z(n7950) );
  XNOR U8030 ( .A(n7949), .B(n7950), .Z(n7956) );
  NANDN U8031 ( .A(n7738), .B(n7737), .Z(n7742) );
  NAND U8032 ( .A(n7740), .B(n7739), .Z(n7741) );
  AND U8033 ( .A(n7742), .B(n7741), .Z(n7944) );
  NANDN U8034 ( .A(n7744), .B(n7743), .Z(n7748) );
  NAND U8035 ( .A(n7746), .B(n7745), .Z(n7747) );
  AND U8036 ( .A(n7748), .B(n7747), .Z(n7942) );
  NANDN U8037 ( .A(n7750), .B(n7749), .Z(n7754) );
  NANDN U8038 ( .A(n7752), .B(n7751), .Z(n7753) );
  AND U8039 ( .A(n7754), .B(n7753), .Z(n7867) );
  AND U8040 ( .A(x[64]), .B(y[280]), .Z(n7924) );
  AND U8041 ( .A(x[88]), .B(y[256]), .Z(n7923) );
  XOR U8042 ( .A(n7924), .B(n7923), .Z(n7926) );
  AND U8043 ( .A(x[87]), .B(y[257]), .Z(n7916) );
  XOR U8044 ( .A(n7916), .B(o[88]), .Z(n7925) );
  XOR U8045 ( .A(n7926), .B(n7925), .Z(n7865) );
  AND U8046 ( .A(x[71]), .B(y[273]), .Z(n7910) );
  NAND U8047 ( .A(x[82]), .B(y[262]), .Z(n7911) );
  XNOR U8048 ( .A(n7910), .B(n7911), .Z(n7912) );
  NAND U8049 ( .A(x[81]), .B(y[263]), .Z(n7913) );
  XNOR U8050 ( .A(n7912), .B(n7913), .Z(n7864) );
  XOR U8051 ( .A(n7865), .B(n7864), .Z(n7866) );
  XNOR U8052 ( .A(n7867), .B(n7866), .Z(n7844) );
  NANDN U8053 ( .A(n7756), .B(n7755), .Z(n7760) );
  NANDN U8054 ( .A(n7758), .B(n7757), .Z(n7759) );
  AND U8055 ( .A(n7760), .B(n7759), .Z(n7842) );
  NANDN U8056 ( .A(n7762), .B(n7761), .Z(n7766) );
  NANDN U8057 ( .A(n7764), .B(n7763), .Z(n7765) );
  NAND U8058 ( .A(n7766), .B(n7765), .Z(n7841) );
  XNOR U8059 ( .A(n7842), .B(n7841), .Z(n7843) );
  XOR U8060 ( .A(n7844), .B(n7843), .Z(n7941) );
  XNOR U8061 ( .A(n7942), .B(n7941), .Z(n7943) );
  XOR U8062 ( .A(n7944), .B(n7943), .Z(n7837) );
  NANDN U8063 ( .A(n7768), .B(n7767), .Z(n7772) );
  NAND U8064 ( .A(n7770), .B(n7769), .Z(n7771) );
  AND U8065 ( .A(n7772), .B(n7771), .Z(n7885) );
  NAND U8066 ( .A(n7774), .B(n7773), .Z(n7778) );
  NANDN U8067 ( .A(n7776), .B(n7775), .Z(n7777) );
  AND U8068 ( .A(n7778), .B(n7777), .Z(n7882) );
  NAND U8069 ( .A(n7780), .B(n7779), .Z(n7784) );
  NANDN U8070 ( .A(n7782), .B(n7781), .Z(n7783) );
  NAND U8071 ( .A(n7784), .B(n7783), .Z(n7883) );
  XOR U8072 ( .A(n7885), .B(n7884), .Z(n7835) );
  NAND U8073 ( .A(n7786), .B(n7785), .Z(n7790) );
  NANDN U8074 ( .A(n7788), .B(n7787), .Z(n7789) );
  NAND U8075 ( .A(n7790), .B(n7789), .Z(n7836) );
  XNOR U8076 ( .A(n7835), .B(n7836), .Z(n7838) );
  XOR U8077 ( .A(n7837), .B(n7838), .Z(n7953) );
  NANDN U8078 ( .A(n7792), .B(n7791), .Z(n7796) );
  NANDN U8079 ( .A(n7794), .B(n7793), .Z(n7795) );
  NAND U8080 ( .A(n7796), .B(n7795), .Z(n7954) );
  XNOR U8081 ( .A(n7953), .B(n7954), .Z(n7955) );
  XOR U8082 ( .A(n7956), .B(n7955), .Z(n7963) );
  NAND U8083 ( .A(n7798), .B(n7797), .Z(n7802) );
  NANDN U8084 ( .A(n7800), .B(n7799), .Z(n7801) );
  AND U8085 ( .A(n7802), .B(n7801), .Z(n7832) );
  NANDN U8086 ( .A(n7804), .B(n7803), .Z(n7808) );
  NANDN U8087 ( .A(n7806), .B(n7805), .Z(n7807) );
  AND U8088 ( .A(n7808), .B(n7807), .Z(n7830) );
  NANDN U8089 ( .A(n7810), .B(n7809), .Z(n7814) );
  NAND U8090 ( .A(n7812), .B(n7811), .Z(n7813) );
  NAND U8091 ( .A(n7814), .B(n7813), .Z(n7829) );
  XNOR U8092 ( .A(n7830), .B(n7829), .Z(n7831) );
  XNOR U8093 ( .A(n7832), .B(n7831), .Z(n7962) );
  XNOR U8094 ( .A(n7963), .B(n7962), .Z(n7964) );
  XNOR U8095 ( .A(n7965), .B(n7964), .Z(n7961) );
  NANDN U8096 ( .A(n7815), .B(n7816), .Z(n7821) );
  NOR U8097 ( .A(n7817), .B(n7816), .Z(n7819) );
  OR U8098 ( .A(n7819), .B(n7818), .Z(n7820) );
  AND U8099 ( .A(n7821), .B(n7820), .Z(n7959) );
  NANDN U8100 ( .A(n7823), .B(n7822), .Z(n7827) );
  NAND U8101 ( .A(n7825), .B(n7824), .Z(n7826) );
  AND U8102 ( .A(n7827), .B(n7826), .Z(n7960) );
  XOR U8103 ( .A(n7959), .B(n7960), .Z(n7828) );
  XNOR U8104 ( .A(n7961), .B(n7828), .Z(N185) );
  NANDN U8105 ( .A(n7830), .B(n7829), .Z(n7834) );
  NANDN U8106 ( .A(n7832), .B(n7831), .Z(n7833) );
  AND U8107 ( .A(n7834), .B(n7833), .Z(n8106) );
  NANDN U8108 ( .A(n7836), .B(n7835), .Z(n7840) );
  NAND U8109 ( .A(n7838), .B(n7837), .Z(n7839) );
  AND U8110 ( .A(n7840), .B(n7839), .Z(n7978) );
  NANDN U8111 ( .A(n7842), .B(n7841), .Z(n7846) );
  NAND U8112 ( .A(n7844), .B(n7843), .Z(n7845) );
  AND U8113 ( .A(n7846), .B(n7845), .Z(n7982) );
  NANDN U8114 ( .A(n7848), .B(n7847), .Z(n7852) );
  NAND U8115 ( .A(n7850), .B(n7849), .Z(n7851) );
  NAND U8116 ( .A(n7852), .B(n7851), .Z(n7981) );
  XNOR U8117 ( .A(n7982), .B(n7981), .Z(n7984) );
  AND U8118 ( .A(x[85]), .B(y[264]), .Z(n8791) );
  NAND U8119 ( .A(n8791), .B(n7853), .Z(n7857) );
  NANDN U8120 ( .A(n7855), .B(n7854), .Z(n7856) );
  NAND U8121 ( .A(n7857), .B(n7856), .Z(n8074) );
  NAND U8122 ( .A(x[86]), .B(y[259]), .Z(n8050) );
  NAND U8123 ( .A(x[69]), .B(y[276]), .Z(n8048) );
  NAND U8124 ( .A(x[81]), .B(y[264]), .Z(n8049) );
  XOR U8125 ( .A(n8048), .B(n8049), .Z(n8051) );
  XOR U8126 ( .A(n8050), .B(n8051), .Z(n8073) );
  AND U8127 ( .A(y[261]), .B(x[84]), .Z(n7859) );
  NAND U8128 ( .A(y[260]), .B(x[85]), .Z(n7858) );
  XNOR U8129 ( .A(n7859), .B(n7858), .Z(n8059) );
  AND U8130 ( .A(x[83]), .B(y[262]), .Z(n8058) );
  XOR U8131 ( .A(n8059), .B(n8058), .Z(n8072) );
  XOR U8132 ( .A(n8073), .B(n8072), .Z(n8075) );
  XOR U8133 ( .A(n8074), .B(n8075), .Z(n8008) );
  NANDN U8134 ( .A(n8057), .B(n8236), .Z(n7863) );
  NANDN U8135 ( .A(n7861), .B(n7860), .Z(n7862) );
  NAND U8136 ( .A(n7863), .B(n7862), .Z(n8080) );
  NAND U8137 ( .A(x[79]), .B(y[266]), .Z(n8064) );
  NAND U8138 ( .A(x[82]), .B(y[263]), .Z(n8062) );
  NAND U8139 ( .A(x[70]), .B(y[275]), .Z(n8063) );
  XOR U8140 ( .A(n8062), .B(n8063), .Z(n8065) );
  XOR U8141 ( .A(n8064), .B(n8065), .Z(n8079) );
  NAND U8142 ( .A(x[87]), .B(y[258]), .Z(n8047) );
  NAND U8143 ( .A(x[68]), .B(y[277]), .Z(n8044) );
  NAND U8144 ( .A(x[80]), .B(y[265]), .Z(n8045) );
  XOR U8145 ( .A(n8044), .B(n8045), .Z(n8046) );
  XNOR U8146 ( .A(n8047), .B(n8046), .Z(n8078) );
  XOR U8147 ( .A(n8079), .B(n8078), .Z(n8081) );
  XOR U8148 ( .A(n8080), .B(n8081), .Z(n8007) );
  XOR U8149 ( .A(n8008), .B(n8007), .Z(n8010) );
  NAND U8150 ( .A(n7865), .B(n7864), .Z(n7869) );
  NANDN U8151 ( .A(n7867), .B(n7866), .Z(n7868) );
  AND U8152 ( .A(n7869), .B(n7868), .Z(n8009) );
  XOR U8153 ( .A(n8010), .B(n8009), .Z(n8022) );
  NAND U8154 ( .A(n7871), .B(n7870), .Z(n7875) );
  NANDN U8155 ( .A(n7873), .B(n7872), .Z(n7874) );
  AND U8156 ( .A(n7875), .B(n7874), .Z(n8020) );
  NAND U8157 ( .A(n7877), .B(n7876), .Z(n7881) );
  NANDN U8158 ( .A(n7879), .B(n7878), .Z(n7880) );
  NAND U8159 ( .A(n7881), .B(n7880), .Z(n8019) );
  XNOR U8160 ( .A(n8020), .B(n8019), .Z(n8021) );
  XNOR U8161 ( .A(n8022), .B(n8021), .Z(n7983) );
  XOR U8162 ( .A(n7984), .B(n7983), .Z(n7976) );
  NANDN U8163 ( .A(n7883), .B(n7882), .Z(n7887) );
  NAND U8164 ( .A(n7885), .B(n7884), .Z(n7886) );
  NAND U8165 ( .A(n7887), .B(n7886), .Z(n7975) );
  NANDN U8166 ( .A(n7992), .B(n7888), .Z(n7892) );
  NAND U8167 ( .A(n7890), .B(n7889), .Z(n7891) );
  AND U8168 ( .A(n7892), .B(n7891), .Z(n8014) );
  AND U8169 ( .A(x[78]), .B(y[272]), .Z(n8931) );
  NAND U8170 ( .A(n8931), .B(n7893), .Z(n7897) );
  NANDN U8171 ( .A(n7895), .B(n7894), .Z(n7896) );
  NAND U8172 ( .A(n7897), .B(n7896), .Z(n8040) );
  NAND U8173 ( .A(x[75]), .B(y[270]), .Z(n8055) );
  NAND U8174 ( .A(x[76]), .B(y[269]), .Z(n8053) );
  NAND U8175 ( .A(x[71]), .B(y[274]), .Z(n8054) );
  XOR U8176 ( .A(n8053), .B(n8054), .Z(n8056) );
  XOR U8177 ( .A(n8055), .B(n8056), .Z(n8039) );
  NAND U8178 ( .A(x[88]), .B(y[257]), .Z(n8052) );
  XNOR U8179 ( .A(o[89]), .B(n8052), .Z(n8027) );
  AND U8180 ( .A(x[65]), .B(y[280]), .Z(n8026) );
  XOR U8181 ( .A(n8027), .B(n8026), .Z(n8029) );
  AND U8182 ( .A(x[77]), .B(y[268]), .Z(n8028) );
  XOR U8183 ( .A(n8029), .B(n8028), .Z(n8038) );
  XOR U8184 ( .A(n8040), .B(n8041), .Z(n8013) );
  XNOR U8185 ( .A(n8014), .B(n8013), .Z(n8016) );
  AND U8186 ( .A(n7899), .B(n7898), .Z(n7903) );
  NANDN U8187 ( .A(n7901), .B(n7900), .Z(n7902) );
  NANDN U8188 ( .A(n7903), .B(n7902), .Z(n8002) );
  AND U8189 ( .A(n7905), .B(n7904), .Z(n7909) );
  NAND U8190 ( .A(n7907), .B(n7906), .Z(n7908) );
  NANDN U8191 ( .A(n7909), .B(n7908), .Z(n8001) );
  XOR U8192 ( .A(n8002), .B(n8001), .Z(n8003) );
  NANDN U8193 ( .A(n7911), .B(n7910), .Z(n7915) );
  NANDN U8194 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND U8195 ( .A(n7915), .B(n7914), .Z(n7997) );
  NAND U8196 ( .A(x[72]), .B(y[273]), .Z(n7993) );
  XOR U8197 ( .A(n7991), .B(n7992), .Z(n7994) );
  XOR U8198 ( .A(n7993), .B(n7994), .Z(n7996) );
  NAND U8199 ( .A(n7916), .B(o[88]), .Z(n7990) );
  NAND U8200 ( .A(x[89]), .B(y[256]), .Z(n7987) );
  NAND U8201 ( .A(x[64]), .B(y[281]), .Z(n7988) );
  XOR U8202 ( .A(n7987), .B(n7988), .Z(n7989) );
  XNOR U8203 ( .A(n7990), .B(n7989), .Z(n7995) );
  XOR U8204 ( .A(n7996), .B(n7995), .Z(n7998) );
  XOR U8205 ( .A(n7997), .B(n7998), .Z(n8004) );
  XNOR U8206 ( .A(n8003), .B(n8004), .Z(n8015) );
  XOR U8207 ( .A(n8016), .B(n8015), .Z(n8093) );
  NAND U8208 ( .A(n7918), .B(n7917), .Z(n7922) );
  ANDN U8209 ( .B(n7920), .A(n7919), .Z(n7921) );
  ANDN U8210 ( .B(n7922), .A(n7921), .Z(n8069) );
  NAND U8211 ( .A(n7924), .B(n7923), .Z(n7928) );
  NAND U8212 ( .A(n7926), .B(n7925), .Z(n7927) );
  AND U8213 ( .A(n7928), .B(n7927), .Z(n8067) );
  AND U8214 ( .A(x[78]), .B(y[267]), .Z(n8033) );
  AND U8215 ( .A(x[66]), .B(y[279]), .Z(n8032) );
  XOR U8216 ( .A(n8033), .B(n8032), .Z(n8035) );
  AND U8217 ( .A(x[67]), .B(y[278]), .Z(n8034) );
  XOR U8218 ( .A(n8035), .B(n8034), .Z(n8066) );
  XNOR U8219 ( .A(n8067), .B(n8066), .Z(n8068) );
  XNOR U8220 ( .A(n8069), .B(n8068), .Z(n8091) );
  NANDN U8221 ( .A(n7930), .B(n7929), .Z(n7934) );
  NAND U8222 ( .A(n7932), .B(n7931), .Z(n7933) );
  AND U8223 ( .A(n7934), .B(n7933), .Z(n8090) );
  XNOR U8224 ( .A(n8091), .B(n8090), .Z(n8092) );
  XNOR U8225 ( .A(n8093), .B(n8092), .Z(n8084) );
  NAND U8226 ( .A(n7936), .B(n7935), .Z(n7940) );
  NAND U8227 ( .A(n7938), .B(n7937), .Z(n7939) );
  NAND U8228 ( .A(n7940), .B(n7939), .Z(n8085) );
  XNOR U8229 ( .A(n8084), .B(n8085), .Z(n8087) );
  NANDN U8230 ( .A(n7942), .B(n7941), .Z(n7946) );
  NANDN U8231 ( .A(n7944), .B(n7943), .Z(n7945) );
  AND U8232 ( .A(n7946), .B(n7945), .Z(n8086) );
  XOR U8233 ( .A(n8087), .B(n8086), .Z(n7970) );
  NANDN U8234 ( .A(n7948), .B(n7947), .Z(n7952) );
  NANDN U8235 ( .A(n7950), .B(n7949), .Z(n7951) );
  AND U8236 ( .A(n7952), .B(n7951), .Z(n7969) );
  XNOR U8237 ( .A(n7971), .B(n7972), .Z(n8104) );
  NANDN U8238 ( .A(n7954), .B(n7953), .Z(n7958) );
  NAND U8239 ( .A(n7956), .B(n7955), .Z(n7957) );
  NAND U8240 ( .A(n7958), .B(n7957), .Z(n8103) );
  XOR U8241 ( .A(n8104), .B(n8103), .Z(n8105) );
  XNOR U8242 ( .A(n8106), .B(n8105), .Z(n8099) );
  NANDN U8243 ( .A(n7963), .B(n7962), .Z(n7967) );
  NAND U8244 ( .A(n7965), .B(n7964), .Z(n7966) );
  AND U8245 ( .A(n7967), .B(n7966), .Z(n8098) );
  IV U8246 ( .A(n8098), .Z(n8096) );
  XOR U8247 ( .A(n8097), .B(n8096), .Z(n7968) );
  XNOR U8248 ( .A(n8099), .B(n7968), .Z(N186) );
  NANDN U8249 ( .A(n7970), .B(n7969), .Z(n7974) );
  NAND U8250 ( .A(n7972), .B(n7971), .Z(n7973) );
  AND U8251 ( .A(n7974), .B(n7973), .Z(n8111) );
  NANDN U8252 ( .A(n7976), .B(n7975), .Z(n7980) );
  NANDN U8253 ( .A(n7978), .B(n7977), .Z(n7979) );
  AND U8254 ( .A(n7980), .B(n7979), .Z(n8110) );
  NANDN U8255 ( .A(n7982), .B(n7981), .Z(n7986) );
  NAND U8256 ( .A(n7984), .B(n7983), .Z(n7985) );
  AND U8257 ( .A(n7986), .B(n7985), .Z(n8257) );
  AND U8258 ( .A(x[66]), .B(y[280]), .Z(n8135) );
  XOR U8259 ( .A(n8136), .B(n8135), .Z(n8138) );
  NAND U8260 ( .A(x[88]), .B(y[258]), .Z(n8137) );
  XNOR U8261 ( .A(n8138), .B(n8137), .Z(n8172) );
  XOR U8262 ( .A(n8172), .B(n8171), .Z(n8174) );
  XOR U8263 ( .A(n8174), .B(n8173), .Z(n8205) );
  NANDN U8264 ( .A(n7996), .B(n7995), .Z(n8000) );
  NANDN U8265 ( .A(n7998), .B(n7997), .Z(n7999) );
  AND U8266 ( .A(n8000), .B(n7999), .Z(n8204) );
  XNOR U8267 ( .A(n8205), .B(n8204), .Z(n8207) );
  NAND U8268 ( .A(n8002), .B(n8001), .Z(n8006) );
  NANDN U8269 ( .A(n8004), .B(n8003), .Z(n8005) );
  AND U8270 ( .A(n8006), .B(n8005), .Z(n8206) );
  XOR U8271 ( .A(n8207), .B(n8206), .Z(n8251) );
  NAND U8272 ( .A(n8008), .B(n8007), .Z(n8012) );
  NAND U8273 ( .A(n8010), .B(n8009), .Z(n8011) );
  AND U8274 ( .A(n8012), .B(n8011), .Z(n8249) );
  NANDN U8275 ( .A(n8014), .B(n8013), .Z(n8018) );
  NAND U8276 ( .A(n8016), .B(n8015), .Z(n8017) );
  AND U8277 ( .A(n8018), .B(n8017), .Z(n8248) );
  XNOR U8278 ( .A(n8249), .B(n8248), .Z(n8250) );
  XOR U8279 ( .A(n8251), .B(n8250), .Z(n8255) );
  NANDN U8280 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U8281 ( .A(n8022), .B(n8021), .Z(n8023) );
  AND U8282 ( .A(n8024), .B(n8023), .Z(n8201) );
  NAND U8283 ( .A(y[276]), .B(x[70]), .Z(n8025) );
  XNOR U8284 ( .A(n8440), .B(n8025), .Z(n8237) );
  NAND U8285 ( .A(x[73]), .B(y[273]), .Z(n8238) );
  XNOR U8286 ( .A(n8237), .B(n8238), .Z(n8210) );
  NAND U8287 ( .A(x[71]), .B(y[275]), .Z(n8211) );
  XNOR U8288 ( .A(n8210), .B(n8211), .Z(n8212) );
  AND U8289 ( .A(x[76]), .B(y[270]), .Z(n8322) );
  AND U8290 ( .A(x[69]), .B(y[277]), .Z(n8181) );
  XOR U8291 ( .A(n8322), .B(n8181), .Z(n8183) );
  NAND U8292 ( .A(x[74]), .B(y[272]), .Z(n8182) );
  XOR U8293 ( .A(n8183), .B(n8182), .Z(n8213) );
  XNOR U8294 ( .A(n8212), .B(n8213), .Z(n8162) );
  NAND U8295 ( .A(n8027), .B(n8026), .Z(n8031) );
  NAND U8296 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U8297 ( .A(n8031), .B(n8030), .Z(n8160) );
  NAND U8298 ( .A(n8033), .B(n8032), .Z(n8037) );
  NAND U8299 ( .A(n8035), .B(n8034), .Z(n8036) );
  NAND U8300 ( .A(n8037), .B(n8036), .Z(n8159) );
  XNOR U8301 ( .A(n8160), .B(n8159), .Z(n8161) );
  XOR U8302 ( .A(n8162), .B(n8161), .Z(n8193) );
  NANDN U8303 ( .A(n8039), .B(n8038), .Z(n8043) );
  NAND U8304 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U8305 ( .A(n8043), .B(n8042), .Z(n8192) );
  XNOR U8306 ( .A(n8193), .B(n8192), .Z(n8195) );
  XNOR U8307 ( .A(n8125), .B(n8126), .Z(n8128) );
  ANDN U8308 ( .B(o[89]), .A(n8052), .Z(n8230) );
  NAND U8309 ( .A(x[78]), .B(y[268]), .Z(n8231) );
  XNOR U8310 ( .A(n8230), .B(n8231), .Z(n8232) );
  NAND U8311 ( .A(x[65]), .B(y[281]), .Z(n8233) );
  XNOR U8312 ( .A(n8232), .B(n8233), .Z(n8176) );
  NAND U8313 ( .A(x[89]), .B(y[257]), .Z(n8241) );
  XNOR U8314 ( .A(o[90]), .B(n8241), .Z(n8186) );
  NAND U8315 ( .A(x[90]), .B(y[256]), .Z(n8187) );
  XNOR U8316 ( .A(n8186), .B(n8187), .Z(n8189) );
  AND U8317 ( .A(x[64]), .B(y[282]), .Z(n8188) );
  XOR U8318 ( .A(n8189), .B(n8188), .Z(n8175) );
  XOR U8319 ( .A(n8176), .B(n8175), .Z(n8178) );
  XOR U8320 ( .A(n8178), .B(n8177), .Z(n8127) );
  XOR U8321 ( .A(n8128), .B(n8127), .Z(n8168) );
  AND U8322 ( .A(x[85]), .B(y[261]), .Z(n8224) );
  NANDN U8323 ( .A(n8057), .B(n8224), .Z(n8061) );
  NAND U8324 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U8325 ( .A(n8061), .B(n8060), .Z(n8156) );
  XOR U8326 ( .A(n8225), .B(n8224), .Z(n8227) );
  NAND U8327 ( .A(x[84]), .B(y[262]), .Z(n8226) );
  XNOR U8328 ( .A(n8227), .B(n8226), .Z(n8153) );
  NAND U8329 ( .A(x[87]), .B(y[259]), .Z(n8142) );
  XNOR U8330 ( .A(n8141), .B(n8142), .Z(n8143) );
  NAND U8331 ( .A(x[86]), .B(y[260]), .Z(n8144) );
  XOR U8332 ( .A(n8143), .B(n8144), .Z(n8154) );
  XNOR U8333 ( .A(n8153), .B(n8154), .Z(n8155) );
  XOR U8334 ( .A(n8156), .B(n8155), .Z(n8166) );
  AND U8335 ( .A(x[83]), .B(y[263]), .Z(n8216) );
  NAND U8336 ( .A(x[75]), .B(y[271]), .Z(n8217) );
  XNOR U8337 ( .A(n8216), .B(n8217), .Z(n8218) );
  NAND U8338 ( .A(x[67]), .B(y[279]), .Z(n8219) );
  XNOR U8339 ( .A(n8218), .B(n8219), .Z(n8132) );
  NAND U8340 ( .A(x[68]), .B(y[278]), .Z(n8148) );
  XNOR U8341 ( .A(n8147), .B(n8148), .Z(n8149) );
  XOR U8342 ( .A(n8132), .B(n8131), .Z(n8134) );
  XNOR U8343 ( .A(n8134), .B(n8133), .Z(n8165) );
  XOR U8344 ( .A(n8166), .B(n8165), .Z(n8167) );
  XNOR U8345 ( .A(n8168), .B(n8167), .Z(n8194) );
  XOR U8346 ( .A(n8195), .B(n8194), .Z(n8199) );
  NANDN U8347 ( .A(n8067), .B(n8066), .Z(n8071) );
  NANDN U8348 ( .A(n8069), .B(n8068), .Z(n8070) );
  AND U8349 ( .A(n8071), .B(n8070), .Z(n8245) );
  NANDN U8350 ( .A(n8073), .B(n8072), .Z(n8077) );
  NANDN U8351 ( .A(n8075), .B(n8074), .Z(n8076) );
  AND U8352 ( .A(n8077), .B(n8076), .Z(n8243) );
  NANDN U8353 ( .A(n8079), .B(n8078), .Z(n8083) );
  NANDN U8354 ( .A(n8081), .B(n8080), .Z(n8082) );
  NAND U8355 ( .A(n8083), .B(n8082), .Z(n8242) );
  XNOR U8356 ( .A(n8243), .B(n8242), .Z(n8244) );
  XNOR U8357 ( .A(n8245), .B(n8244), .Z(n8198) );
  XNOR U8358 ( .A(n8199), .B(n8198), .Z(n8200) );
  XNOR U8359 ( .A(n8201), .B(n8200), .Z(n8254) );
  XNOR U8360 ( .A(n8255), .B(n8254), .Z(n8256) );
  XNOR U8361 ( .A(n8257), .B(n8256), .Z(n8122) );
  NANDN U8362 ( .A(n8085), .B(n8084), .Z(n8089) );
  NAND U8363 ( .A(n8087), .B(n8086), .Z(n8088) );
  AND U8364 ( .A(n8089), .B(n8088), .Z(n8119) );
  NANDN U8365 ( .A(n8091), .B(n8090), .Z(n8095) );
  NANDN U8366 ( .A(n8093), .B(n8092), .Z(n8094) );
  NAND U8367 ( .A(n8095), .B(n8094), .Z(n8120) );
  XNOR U8368 ( .A(n8119), .B(n8120), .Z(n8121) );
  XOR U8369 ( .A(n8122), .B(n8121), .Z(n8112) );
  XNOR U8370 ( .A(n8113), .B(n8112), .Z(n8118) );
  NANDN U8371 ( .A(n8096), .B(n8097), .Z(n8102) );
  NOR U8372 ( .A(n8098), .B(n8097), .Z(n8100) );
  OR U8373 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8374 ( .A(n8102), .B(n8101), .Z(n8116) );
  NAND U8375 ( .A(n8104), .B(n8103), .Z(n8108) );
  NAND U8376 ( .A(n8106), .B(n8105), .Z(n8107) );
  AND U8377 ( .A(n8108), .B(n8107), .Z(n8117) );
  XOR U8378 ( .A(n8116), .B(n8117), .Z(n8109) );
  XNOR U8379 ( .A(n8118), .B(n8109), .Z(N187) );
  NANDN U8380 ( .A(n8111), .B(n8110), .Z(n8115) );
  NAND U8381 ( .A(n8113), .B(n8112), .Z(n8114) );
  NAND U8382 ( .A(n8115), .B(n8114), .Z(n8268) );
  IV U8383 ( .A(n8268), .Z(n8267) );
  NANDN U8384 ( .A(n8120), .B(n8119), .Z(n8124) );
  NAND U8385 ( .A(n8122), .B(n8121), .Z(n8123) );
  AND U8386 ( .A(n8124), .B(n8123), .Z(n8264) );
  NANDN U8387 ( .A(n8126), .B(n8125), .Z(n8130) );
  NAND U8388 ( .A(n8128), .B(n8127), .Z(n8129) );
  NAND U8389 ( .A(n8130), .B(n8129), .Z(n8385) );
  NAND U8390 ( .A(n8136), .B(n8135), .Z(n8140) );
  ANDN U8391 ( .B(n8138), .A(n8137), .Z(n8139) );
  ANDN U8392 ( .B(n8140), .A(n8139), .Z(n8299) );
  NANDN U8393 ( .A(n8142), .B(n8141), .Z(n8146) );
  NANDN U8394 ( .A(n8144), .B(n8143), .Z(n8145) );
  NAND U8395 ( .A(n8146), .B(n8145), .Z(n8298) );
  XNOR U8396 ( .A(n8299), .B(n8298), .Z(n8300) );
  NANDN U8397 ( .A(n8148), .B(n8147), .Z(n8152) );
  NANDN U8398 ( .A(n8150), .B(n8149), .Z(n8151) );
  AND U8399 ( .A(n8152), .B(n8151), .Z(n8311) );
  AND U8400 ( .A(x[64]), .B(y[283]), .Z(n8375) );
  NAND U8401 ( .A(x[91]), .B(y[256]), .Z(n8376) );
  XNOR U8402 ( .A(n8375), .B(n8376), .Z(n8378) );
  NAND U8403 ( .A(x[90]), .B(y[257]), .Z(n8366) );
  XOR U8404 ( .A(n8378), .B(n8377), .Z(n8308) );
  AND U8405 ( .A(x[73]), .B(y[274]), .Z(n8360) );
  NAND U8406 ( .A(x[85]), .B(y[262]), .Z(n8361) );
  XNOR U8407 ( .A(n8360), .B(n8361), .Z(n8362) );
  NAND U8408 ( .A(x[82]), .B(y[265]), .Z(n8363) );
  XOR U8409 ( .A(n8362), .B(n8363), .Z(n8309) );
  XNOR U8410 ( .A(n8308), .B(n8309), .Z(n8310) );
  XOR U8411 ( .A(n8311), .B(n8310), .Z(n8301) );
  XNOR U8412 ( .A(n8300), .B(n8301), .Z(n8384) );
  XOR U8413 ( .A(n8383), .B(n8384), .Z(n8386) );
  XOR U8414 ( .A(n8385), .B(n8386), .Z(n8402) );
  NANDN U8415 ( .A(n8154), .B(n8153), .Z(n8158) );
  NANDN U8416 ( .A(n8156), .B(n8155), .Z(n8157) );
  AND U8417 ( .A(n8158), .B(n8157), .Z(n8400) );
  NANDN U8418 ( .A(n8160), .B(n8159), .Z(n8164) );
  NAND U8419 ( .A(n8162), .B(n8161), .Z(n8163) );
  AND U8420 ( .A(n8164), .B(n8163), .Z(n8399) );
  XOR U8421 ( .A(n8400), .B(n8399), .Z(n8401) );
  NAND U8422 ( .A(n8166), .B(n8165), .Z(n8170) );
  NANDN U8423 ( .A(n8168), .B(n8167), .Z(n8169) );
  AND U8424 ( .A(n8170), .B(n8169), .Z(n8387) );
  AND U8425 ( .A(x[79]), .B(y[268]), .Z(n8328) );
  AND U8426 ( .A(x[66]), .B(y[281]), .Z(n8327) );
  XOR U8427 ( .A(n8328), .B(n8327), .Z(n8330) );
  AND U8428 ( .A(x[67]), .B(y[280]), .Z(n8329) );
  XOR U8429 ( .A(n8330), .B(n8329), .Z(n8343) );
  AND U8430 ( .A(x[83]), .B(y[264]), .Z(n8354) );
  NAND U8431 ( .A(x[89]), .B(y[258]), .Z(n8355) );
  XNOR U8432 ( .A(n8354), .B(n8355), .Z(n8356) );
  NAND U8433 ( .A(x[70]), .B(y[277]), .Z(n8357) );
  XOR U8434 ( .A(n8356), .B(n8357), .Z(n8344) );
  XNOR U8435 ( .A(n8343), .B(n8344), .Z(n8345) );
  NAND U8436 ( .A(x[80]), .B(y[267]), .Z(n8314) );
  XOR U8437 ( .A(n8314), .B(n8315), .Z(n8317) );
  XOR U8438 ( .A(n8316), .B(n8317), .Z(n8324) );
  AND U8439 ( .A(y[270]), .B(x[77]), .Z(n8180) );
  NAND U8440 ( .A(y[271]), .B(x[76]), .Z(n8179) );
  XNOR U8441 ( .A(n8180), .B(n8179), .Z(n8323) );
  XOR U8442 ( .A(n8324), .B(n8323), .Z(n8346) );
  XNOR U8443 ( .A(n8345), .B(n8346), .Z(n8295) );
  NAND U8444 ( .A(n8322), .B(n8181), .Z(n8185) );
  ANDN U8445 ( .B(n8183), .A(n8182), .Z(n8184) );
  ANDN U8446 ( .B(n8185), .A(n8184), .Z(n8293) );
  NANDN U8447 ( .A(n8187), .B(n8186), .Z(n8191) );
  NAND U8448 ( .A(n8189), .B(n8188), .Z(n8190) );
  NAND U8449 ( .A(n8191), .B(n8190), .Z(n8292) );
  XNOR U8450 ( .A(n8293), .B(n8292), .Z(n8294) );
  XOR U8451 ( .A(n8295), .B(n8294), .Z(n8379) );
  XNOR U8452 ( .A(n8380), .B(n8379), .Z(n8382) );
  XOR U8453 ( .A(n8381), .B(n8382), .Z(n8388) );
  NANDN U8454 ( .A(n8193), .B(n8192), .Z(n8197) );
  NAND U8455 ( .A(n8195), .B(n8194), .Z(n8196) );
  AND U8456 ( .A(n8197), .B(n8196), .Z(n8389) );
  XOR U8457 ( .A(n8390), .B(n8389), .Z(n8280) );
  NANDN U8458 ( .A(n8199), .B(n8198), .Z(n8203) );
  NANDN U8459 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND U8460 ( .A(n8203), .B(n8202), .Z(n8282) );
  XOR U8461 ( .A(n8283), .B(n8282), .Z(n8277) );
  NANDN U8462 ( .A(n8205), .B(n8204), .Z(n8209) );
  NAND U8463 ( .A(n8207), .B(n8206), .Z(n8208) );
  NAND U8464 ( .A(n8209), .B(n8208), .Z(n8286) );
  NANDN U8465 ( .A(n8211), .B(n8210), .Z(n8215) );
  NANDN U8466 ( .A(n8213), .B(n8212), .Z(n8214) );
  AND U8467 ( .A(n8215), .B(n8214), .Z(n8395) );
  NANDN U8468 ( .A(n8217), .B(n8216), .Z(n8221) );
  NANDN U8469 ( .A(n8219), .B(n8218), .Z(n8220) );
  AND U8470 ( .A(n8221), .B(n8220), .Z(n8342) );
  NAND U8471 ( .A(y[259]), .B(x[88]), .Z(n8222) );
  XNOR U8472 ( .A(n8223), .B(n8222), .Z(n8350) );
  NAND U8473 ( .A(x[71]), .B(y[276]), .Z(n8351) );
  XNOR U8474 ( .A(n8350), .B(n8351), .Z(n8340) );
  AND U8475 ( .A(x[72]), .B(y[275]), .Z(n8319) );
  AND U8476 ( .A(x[87]), .B(y[260]), .Z(n8318) );
  XOR U8477 ( .A(n8319), .B(n8318), .Z(n8321) );
  AND U8478 ( .A(x[86]), .B(y[261]), .Z(n8320) );
  XOR U8479 ( .A(n8321), .B(n8320), .Z(n8339) );
  XOR U8480 ( .A(n8340), .B(n8339), .Z(n8341) );
  XOR U8481 ( .A(n8342), .B(n8341), .Z(n8393) );
  NAND U8482 ( .A(n8225), .B(n8224), .Z(n8229) );
  ANDN U8483 ( .B(n8227), .A(n8226), .Z(n8228) );
  ANDN U8484 ( .B(n8229), .A(n8228), .Z(n8336) );
  NANDN U8485 ( .A(n8231), .B(n8230), .Z(n8235) );
  NANDN U8486 ( .A(n8233), .B(n8232), .Z(n8234) );
  NAND U8487 ( .A(n8235), .B(n8234), .Z(n8335) );
  XNOR U8488 ( .A(n8336), .B(n8335), .Z(n8338) );
  AND U8489 ( .A(x[72]), .B(y[276]), .Z(n8368) );
  NAND U8490 ( .A(n8236), .B(n8368), .Z(n8240) );
  NANDN U8491 ( .A(n8238), .B(n8237), .Z(n8239) );
  NAND U8492 ( .A(n8240), .B(n8239), .Z(n8306) );
  AND U8493 ( .A(x[78]), .B(y[269]), .Z(n8332) );
  AND U8494 ( .A(x[65]), .B(y[282]), .Z(n8331) );
  XOR U8495 ( .A(n8332), .B(n8331), .Z(n8334) );
  ANDN U8496 ( .B(o[90]), .A(n8241), .Z(n8333) );
  XOR U8497 ( .A(n8334), .B(n8333), .Z(n8305) );
  AND U8498 ( .A(x[81]), .B(y[266]), .Z(n8369) );
  NAND U8499 ( .A(x[68]), .B(y[279]), .Z(n8370) );
  XNOR U8500 ( .A(n8369), .B(n8370), .Z(n8372) );
  AND U8501 ( .A(x[69]), .B(y[278]), .Z(n8371) );
  XOR U8502 ( .A(n8372), .B(n8371), .Z(n8304) );
  XOR U8503 ( .A(n8305), .B(n8304), .Z(n8307) );
  XOR U8504 ( .A(n8306), .B(n8307), .Z(n8337) );
  XOR U8505 ( .A(n8338), .B(n8337), .Z(n8394) );
  XNOR U8506 ( .A(n8395), .B(n8396), .Z(n8287) );
  XOR U8507 ( .A(n8286), .B(n8287), .Z(n8289) );
  NANDN U8508 ( .A(n8243), .B(n8242), .Z(n8247) );
  NANDN U8509 ( .A(n8245), .B(n8244), .Z(n8246) );
  AND U8510 ( .A(n8247), .B(n8246), .Z(n8288) );
  XOR U8511 ( .A(n8289), .B(n8288), .Z(n8275) );
  NANDN U8512 ( .A(n8249), .B(n8248), .Z(n8253) );
  NAND U8513 ( .A(n8251), .B(n8250), .Z(n8252) );
  AND U8514 ( .A(n8253), .B(n8252), .Z(n8274) );
  XNOR U8515 ( .A(n8275), .B(n8274), .Z(n8276) );
  XOR U8516 ( .A(n8277), .B(n8276), .Z(n8262) );
  NANDN U8517 ( .A(n8255), .B(n8254), .Z(n8259) );
  NANDN U8518 ( .A(n8257), .B(n8256), .Z(n8258) );
  AND U8519 ( .A(n8259), .B(n8258), .Z(n8261) );
  XNOR U8520 ( .A(n8262), .B(n8261), .Z(n8263) );
  XOR U8521 ( .A(n8264), .B(n8263), .Z(n8270) );
  XNOR U8522 ( .A(n8269), .B(n8270), .Z(n8260) );
  XOR U8523 ( .A(n8267), .B(n8260), .Z(N188) );
  NANDN U8524 ( .A(n8262), .B(n8261), .Z(n8266) );
  NAND U8525 ( .A(n8264), .B(n8263), .Z(n8265) );
  NAND U8526 ( .A(n8266), .B(n8265), .Z(n8559) );
  IV U8527 ( .A(n8559), .Z(n8557) );
  OR U8528 ( .A(n8269), .B(n8267), .Z(n8273) );
  ANDN U8529 ( .B(n8269), .A(n8268), .Z(n8271) );
  OR U8530 ( .A(n8271), .B(n8270), .Z(n8272) );
  AND U8531 ( .A(n8273), .B(n8272), .Z(n8558) );
  NANDN U8532 ( .A(n8275), .B(n8274), .Z(n8279) );
  NAND U8533 ( .A(n8277), .B(n8276), .Z(n8278) );
  AND U8534 ( .A(n8279), .B(n8278), .Z(n8552) );
  NANDN U8535 ( .A(n8281), .B(n8280), .Z(n8285) );
  NAND U8536 ( .A(n8283), .B(n8282), .Z(n8284) );
  NAND U8537 ( .A(n8285), .B(n8284), .Z(n8551) );
  XNOR U8538 ( .A(n8552), .B(n8551), .Z(n8554) );
  NAND U8539 ( .A(n8287), .B(n8286), .Z(n8291) );
  NAND U8540 ( .A(n8289), .B(n8288), .Z(n8290) );
  AND U8541 ( .A(n8291), .B(n8290), .Z(n8407) );
  NANDN U8542 ( .A(n8293), .B(n8292), .Z(n8297) );
  NAND U8543 ( .A(n8295), .B(n8294), .Z(n8296) );
  AND U8544 ( .A(n8297), .B(n8296), .Z(n8419) );
  NANDN U8545 ( .A(n8299), .B(n8298), .Z(n8303) );
  NANDN U8546 ( .A(n8301), .B(n8300), .Z(n8302) );
  AND U8547 ( .A(n8303), .B(n8302), .Z(n8522) );
  NANDN U8548 ( .A(n8309), .B(n8308), .Z(n8313) );
  NANDN U8549 ( .A(n8311), .B(n8310), .Z(n8312) );
  NAND U8550 ( .A(n8313), .B(n8312), .Z(n8519) );
  XNOR U8551 ( .A(n8520), .B(n8519), .Z(n8521) );
  XNOR U8552 ( .A(n8522), .B(n8521), .Z(n8418) );
  XNOR U8553 ( .A(n8419), .B(n8418), .Z(n8421) );
  AND U8554 ( .A(x[71]), .B(y[277]), .Z(n8464) );
  AND U8555 ( .A(x[76]), .B(y[272]), .Z(n8463) );
  XOR U8556 ( .A(n8464), .B(n8463), .Z(n8466) );
  AND U8557 ( .A(x[75]), .B(y[273]), .Z(n8465) );
  XOR U8558 ( .A(n8466), .B(n8465), .Z(n8496) );
  AND U8559 ( .A(x[91]), .B(y[257]), .Z(n8480) );
  XOR U8560 ( .A(o[92]), .B(n8480), .Z(n8488) );
  AND U8561 ( .A(x[90]), .B(y[258]), .Z(n8487) );
  XOR U8562 ( .A(n8488), .B(n8487), .Z(n8490) );
  AND U8563 ( .A(x[79]), .B(y[269]), .Z(n8489) );
  XNOR U8564 ( .A(n8490), .B(n8489), .Z(n8495) );
  XOR U8565 ( .A(n8497), .B(n8498), .Z(n8538) );
  AND U8566 ( .A(x[81]), .B(y[267]), .Z(n8429) );
  AND U8567 ( .A(x[86]), .B(y[262]), .Z(n8428) );
  XOR U8568 ( .A(n8429), .B(n8428), .Z(n8431) );
  AND U8569 ( .A(x[68]), .B(y[280]), .Z(n8430) );
  XOR U8570 ( .A(n8431), .B(n8430), .Z(n8502) );
  AND U8571 ( .A(x[70]), .B(y[278]), .Z(n8650) );
  AND U8572 ( .A(x[83]), .B(y[265]), .Z(n8469) );
  XOR U8573 ( .A(n8650), .B(n8469), .Z(n8471) );
  XOR U8574 ( .A(n8471), .B(n8470), .Z(n8501) );
  XOR U8575 ( .A(n8502), .B(n8501), .Z(n8504) );
  XOR U8576 ( .A(n8503), .B(n8504), .Z(n8537) );
  XOR U8577 ( .A(n8538), .B(n8537), .Z(n8540) );
  NAND U8578 ( .A(n8322), .B(n8482), .Z(n8326) );
  NANDN U8579 ( .A(n8324), .B(n8323), .Z(n8325) );
  NAND U8580 ( .A(n8326), .B(n8325), .Z(n8424) );
  XOR U8581 ( .A(n8423), .B(n8422), .Z(n8425) );
  XOR U8582 ( .A(n8424), .B(n8425), .Z(n8539) );
  XOR U8583 ( .A(n8540), .B(n8539), .Z(n8420) );
  XOR U8584 ( .A(n8421), .B(n8420), .Z(n8548) );
  NANDN U8585 ( .A(n8344), .B(n8343), .Z(n8348) );
  NANDN U8586 ( .A(n8346), .B(n8345), .Z(n8347) );
  NAND U8587 ( .A(n8348), .B(n8347), .Z(n8507) );
  XNOR U8588 ( .A(n8508), .B(n8507), .Z(n8509) );
  XOR U8589 ( .A(n8510), .B(n8509), .Z(n8545) );
  AND U8590 ( .A(x[88]), .B(y[263]), .Z(n8872) );
  NAND U8591 ( .A(n8872), .B(n8349), .Z(n8353) );
  NANDN U8592 ( .A(n8351), .B(n8350), .Z(n8352) );
  NAND U8593 ( .A(n8353), .B(n8352), .Z(n8536) );
  AND U8594 ( .A(x[89]), .B(y[259]), .Z(n8459) );
  XOR U8595 ( .A(n8460), .B(n8459), .Z(n8458) );
  AND U8596 ( .A(x[65]), .B(y[283]), .Z(n8457) );
  XOR U8597 ( .A(n8458), .B(n8457), .Z(n8534) );
  AND U8598 ( .A(x[80]), .B(y[268]), .Z(n8452) );
  AND U8599 ( .A(x[88]), .B(y[260]), .Z(n8451) );
  XOR U8600 ( .A(n8452), .B(n8451), .Z(n8454) );
  AND U8601 ( .A(x[66]), .B(y[282]), .Z(n8453) );
  XOR U8602 ( .A(n8454), .B(n8453), .Z(n8533) );
  XOR U8603 ( .A(n8534), .B(n8533), .Z(n8535) );
  XNOR U8604 ( .A(n8536), .B(n8535), .Z(n8516) );
  NANDN U8605 ( .A(n8355), .B(n8354), .Z(n8359) );
  NANDN U8606 ( .A(n8357), .B(n8356), .Z(n8358) );
  NAND U8607 ( .A(n8359), .B(n8358), .Z(n8532) );
  AND U8608 ( .A(x[67]), .B(y[281]), .Z(n8481) );
  XOR U8609 ( .A(n8482), .B(n8481), .Z(n8484) );
  AND U8610 ( .A(x[87]), .B(y[261]), .Z(n8483) );
  XOR U8611 ( .A(n8484), .B(n8483), .Z(n8530) );
  AND U8612 ( .A(x[69]), .B(y[279]), .Z(n8475) );
  AND U8613 ( .A(x[85]), .B(y[263]), .Z(n8474) );
  XOR U8614 ( .A(n8475), .B(n8474), .Z(n8477) );
  AND U8615 ( .A(x[84]), .B(y[264]), .Z(n8476) );
  XOR U8616 ( .A(n8477), .B(n8476), .Z(n8529) );
  XOR U8617 ( .A(n8530), .B(n8529), .Z(n8531) );
  XNOR U8618 ( .A(n8532), .B(n8531), .Z(n8514) );
  NANDN U8619 ( .A(n8361), .B(n8360), .Z(n8365) );
  NANDN U8620 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U8621 ( .A(n8365), .B(n8364), .Z(n8447) );
  ANDN U8622 ( .B(o[91]), .A(n8366), .Z(n8437) );
  AND U8623 ( .A(x[64]), .B(y[284]), .Z(n8435) );
  AND U8624 ( .A(x[92]), .B(y[256]), .Z(n8434) );
  XOR U8625 ( .A(n8435), .B(n8434), .Z(n8436) );
  XOR U8626 ( .A(n8437), .B(n8436), .Z(n8446) );
  NAND U8627 ( .A(y[274]), .B(x[74]), .Z(n8367) );
  XNOR U8628 ( .A(n8368), .B(n8367), .Z(n8442) );
  AND U8629 ( .A(x[73]), .B(y[275]), .Z(n8441) );
  XOR U8630 ( .A(n8442), .B(n8441), .Z(n8445) );
  XOR U8631 ( .A(n8446), .B(n8445), .Z(n8448) );
  XOR U8632 ( .A(n8447), .B(n8448), .Z(n8528) );
  NANDN U8633 ( .A(n8370), .B(n8369), .Z(n8374) );
  NAND U8634 ( .A(n8372), .B(n8371), .Z(n8373) );
  NAND U8635 ( .A(n8374), .B(n8373), .Z(n8525) );
  XOR U8636 ( .A(n8525), .B(n8526), .Z(n8527) );
  XNOR U8637 ( .A(n8528), .B(n8527), .Z(n8513) );
  XOR U8638 ( .A(n8514), .B(n8513), .Z(n8515) );
  XOR U8639 ( .A(n8516), .B(n8515), .Z(n8546) );
  XOR U8640 ( .A(n8545), .B(n8546), .Z(n8547) );
  XNOR U8641 ( .A(n8548), .B(n8547), .Z(n8543) );
  XNOR U8642 ( .A(n8541), .B(n8542), .Z(n8544) );
  XOR U8643 ( .A(n8543), .B(n8544), .Z(n8406) );
  XOR U8644 ( .A(n8407), .B(n8406), .Z(n8408) );
  NANDN U8645 ( .A(n8388), .B(n8387), .Z(n8392) );
  NAND U8646 ( .A(n8390), .B(n8389), .Z(n8391) );
  NAND U8647 ( .A(n8392), .B(n8391), .Z(n8414) );
  NANDN U8648 ( .A(n8394), .B(n8393), .Z(n8398) );
  NANDN U8649 ( .A(n8396), .B(n8395), .Z(n8397) );
  AND U8650 ( .A(n8398), .B(n8397), .Z(n8413) );
  NAND U8651 ( .A(n8400), .B(n8399), .Z(n8404) );
  NANDN U8652 ( .A(n8402), .B(n8401), .Z(n8403) );
  AND U8653 ( .A(n8404), .B(n8403), .Z(n8412) );
  XOR U8654 ( .A(n8413), .B(n8412), .Z(n8415) );
  XNOR U8655 ( .A(n8414), .B(n8415), .Z(n8409) );
  XOR U8656 ( .A(n8554), .B(n8553), .Z(n8560) );
  XNOR U8657 ( .A(n8558), .B(n8560), .Z(n8405) );
  XOR U8658 ( .A(n8557), .B(n8405), .Z(N189) );
  NAND U8659 ( .A(n8407), .B(n8406), .Z(n8411) );
  NANDN U8660 ( .A(n8409), .B(n8408), .Z(n8410) );
  NAND U8661 ( .A(n8411), .B(n8410), .Z(n8570) );
  NAND U8662 ( .A(n8413), .B(n8412), .Z(n8417) );
  NAND U8663 ( .A(n8415), .B(n8414), .Z(n8416) );
  NAND U8664 ( .A(n8417), .B(n8416), .Z(n8569) );
  NAND U8665 ( .A(n8423), .B(n8422), .Z(n8427) );
  NAND U8666 ( .A(n8425), .B(n8424), .Z(n8426) );
  AND U8667 ( .A(n8427), .B(n8426), .Z(n8677) );
  NAND U8668 ( .A(n8429), .B(n8428), .Z(n8433) );
  NAND U8669 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U8670 ( .A(n8433), .B(n8432), .Z(n8715) );
  NAND U8671 ( .A(n8435), .B(n8434), .Z(n8439) );
  NAND U8672 ( .A(n8437), .B(n8436), .Z(n8438) );
  NAND U8673 ( .A(n8439), .B(n8438), .Z(n8714) );
  XOR U8674 ( .A(n8715), .B(n8714), .Z(n8716) );
  AND U8675 ( .A(x[74]), .B(y[276]), .Z(n8713) );
  NAND U8676 ( .A(n8440), .B(n8713), .Z(n8444) );
  NAND U8677 ( .A(n8442), .B(n8441), .Z(n8443) );
  NAND U8678 ( .A(n8444), .B(n8443), .Z(n8683) );
  AND U8679 ( .A(x[86]), .B(y[263]), .Z(n8628) );
  AND U8680 ( .A(x[65]), .B(y[284]), .Z(n8626) );
  AND U8681 ( .A(x[76]), .B(y[273]), .Z(n8921) );
  XOR U8682 ( .A(n8626), .B(n8921), .Z(n8627) );
  XOR U8683 ( .A(n8628), .B(n8627), .Z(n8682) );
  AND U8684 ( .A(x[79]), .B(y[270]), .Z(n8631) );
  XOR U8685 ( .A(n8791), .B(n8631), .Z(n8632) );
  XOR U8686 ( .A(n8633), .B(n8632), .Z(n8681) );
  XOR U8687 ( .A(n8682), .B(n8681), .Z(n8684) );
  XNOR U8688 ( .A(n8683), .B(n8684), .Z(n8717) );
  NAND U8689 ( .A(n8446), .B(n8445), .Z(n8450) );
  NAND U8690 ( .A(n8448), .B(n8447), .Z(n8449) );
  AND U8691 ( .A(n8450), .B(n8449), .Z(n8675) );
  XNOR U8692 ( .A(n8677), .B(n8678), .Z(n8672) );
  NAND U8693 ( .A(n8452), .B(n8451), .Z(n8456) );
  NAND U8694 ( .A(n8454), .B(n8453), .Z(n8455) );
  NAND U8695 ( .A(n8456), .B(n8455), .Z(n8688) );
  AND U8696 ( .A(n8458), .B(n8457), .Z(n8462) );
  NAND U8697 ( .A(n8460), .B(n8459), .Z(n8461) );
  NANDN U8698 ( .A(n8462), .B(n8461), .Z(n8687) );
  XOR U8699 ( .A(n8688), .B(n8687), .Z(n8689) );
  NAND U8700 ( .A(n8464), .B(n8463), .Z(n8468) );
  NAND U8701 ( .A(n8466), .B(n8465), .Z(n8467) );
  NAND U8702 ( .A(n8468), .B(n8467), .Z(n8592) );
  AND U8703 ( .A(x[75]), .B(y[274]), .Z(n8647) );
  AND U8704 ( .A(x[67]), .B(y[282]), .Z(n8645) );
  AND U8705 ( .A(x[81]), .B(y[268]), .Z(n8644) );
  XOR U8706 ( .A(n8645), .B(n8644), .Z(n8646) );
  XOR U8707 ( .A(n8647), .B(n8646), .Z(n8591) );
  AND U8708 ( .A(x[87]), .B(y[262]), .Z(n8834) );
  AND U8709 ( .A(x[77]), .B(y[272]), .Z(n8640) );
  AND U8710 ( .A(x[88]), .B(y[261]), .Z(n8639) );
  XOR U8711 ( .A(n8640), .B(n8639), .Z(n8641) );
  XOR U8712 ( .A(n8834), .B(n8641), .Z(n8590) );
  XOR U8713 ( .A(n8591), .B(n8590), .Z(n8593) );
  XNOR U8714 ( .A(n8592), .B(n8593), .Z(n8690) );
  NAND U8715 ( .A(n8650), .B(n8469), .Z(n8473) );
  NAND U8716 ( .A(n8471), .B(n8470), .Z(n8472) );
  AND U8717 ( .A(n8473), .B(n8472), .Z(n8695) );
  AND U8718 ( .A(x[89]), .B(y[260]), .Z(n8623) );
  AND U8719 ( .A(x[90]), .B(y[259]), .Z(n8620) );
  XOR U8720 ( .A(n8621), .B(n8620), .Z(n8622) );
  XOR U8721 ( .A(n8623), .B(n8622), .Z(n8694) );
  AND U8722 ( .A(x[92]), .B(y[257]), .Z(n8636) );
  XOR U8723 ( .A(o[93]), .B(n8636), .Z(n8707) );
  AND U8724 ( .A(x[64]), .B(y[285]), .Z(n8705) );
  AND U8725 ( .A(x[93]), .B(y[256]), .Z(n8704) );
  XOR U8726 ( .A(n8705), .B(n8704), .Z(n8706) );
  XNOR U8727 ( .A(n8707), .B(n8706), .Z(n8693) );
  XNOR U8728 ( .A(n8695), .B(n8696), .Z(n8578) );
  NAND U8729 ( .A(n8475), .B(n8474), .Z(n8479) );
  NAND U8730 ( .A(n8477), .B(n8476), .Z(n8478) );
  NAND U8731 ( .A(n8479), .B(n8478), .Z(n8659) );
  AND U8732 ( .A(o[92]), .B(n8480), .Z(n8599) );
  AND U8733 ( .A(x[80]), .B(y[269]), .Z(n8597) );
  AND U8734 ( .A(x[91]), .B(y[258]), .Z(n8596) );
  XOR U8735 ( .A(n8597), .B(n8596), .Z(n8598) );
  XOR U8736 ( .A(n8599), .B(n8598), .Z(n8658) );
  AND U8737 ( .A(x[66]), .B(y[283]), .Z(n8608) );
  XOR U8738 ( .A(n8609), .B(n8608), .Z(n8610) );
  XOR U8739 ( .A(n8611), .B(n8610), .Z(n8657) );
  XOR U8740 ( .A(n8658), .B(n8657), .Z(n8660) );
  XOR U8741 ( .A(n8659), .B(n8660), .Z(n8579) );
  NAND U8742 ( .A(n8482), .B(n8481), .Z(n8486) );
  NAND U8743 ( .A(n8484), .B(n8483), .Z(n8485) );
  NAND U8744 ( .A(n8486), .B(n8485), .Z(n8615) );
  NAND U8745 ( .A(n8488), .B(n8487), .Z(n8492) );
  NAND U8746 ( .A(n8490), .B(n8489), .Z(n8491) );
  NAND U8747 ( .A(n8492), .B(n8491), .Z(n8614) );
  XOR U8748 ( .A(n8615), .B(n8614), .Z(n8617) );
  AND U8749 ( .A(x[73]), .B(y[276]), .Z(n8888) );
  AND U8750 ( .A(x[72]), .B(y[277]), .Z(n8652) );
  AND U8751 ( .A(y[279]), .B(x[70]), .Z(n8494) );
  NAND U8752 ( .A(y[278]), .B(x[71]), .Z(n8493) );
  XNOR U8753 ( .A(n8494), .B(n8493), .Z(n8651) );
  XOR U8754 ( .A(n8652), .B(n8651), .Z(n8699) );
  XOR U8755 ( .A(n8888), .B(n8699), .Z(n8701) );
  AND U8756 ( .A(x[69]), .B(y[280]), .Z(n8605) );
  AND U8757 ( .A(x[68]), .B(y[281]), .Z(n8603) );
  AND U8758 ( .A(x[74]), .B(y[275]), .Z(n8602) );
  XOR U8759 ( .A(n8603), .B(n8602), .Z(n8604) );
  XOR U8760 ( .A(n8605), .B(n8604), .Z(n8700) );
  XOR U8761 ( .A(n8701), .B(n8700), .Z(n8616) );
  XOR U8762 ( .A(n8617), .B(n8616), .Z(n8585) );
  NANDN U8763 ( .A(n8496), .B(n8495), .Z(n8500) );
  NANDN U8764 ( .A(n8498), .B(n8497), .Z(n8499) );
  NAND U8765 ( .A(n8500), .B(n8499), .Z(n8584) );
  XNOR U8766 ( .A(n8586), .B(n8587), .Z(n8670) );
  NAND U8767 ( .A(n8502), .B(n8501), .Z(n8506) );
  NAND U8768 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U8769 ( .A(n8506), .B(n8505), .Z(n8669) );
  XNOR U8770 ( .A(n8736), .B(n8735), .Z(n8738) );
  NANDN U8771 ( .A(n8508), .B(n8507), .Z(n8512) );
  NANDN U8772 ( .A(n8510), .B(n8509), .Z(n8511) );
  AND U8773 ( .A(n8512), .B(n8511), .Z(n8729) );
  NAND U8774 ( .A(n8514), .B(n8513), .Z(n8518) );
  NAND U8775 ( .A(n8516), .B(n8515), .Z(n8517) );
  AND U8776 ( .A(n8518), .B(n8517), .Z(n8728) );
  XNOR U8777 ( .A(n8729), .B(n8728), .Z(n8731) );
  NANDN U8778 ( .A(n8520), .B(n8519), .Z(n8524) );
  NANDN U8779 ( .A(n8522), .B(n8521), .Z(n8523) );
  NAND U8780 ( .A(n8524), .B(n8523), .Z(n8723) );
  XOR U8781 ( .A(n8664), .B(n8663), .Z(n8666) );
  XOR U8782 ( .A(n8665), .B(n8666), .Z(n8721) );
  XOR U8783 ( .A(n8721), .B(n8720), .Z(n8724) );
  XOR U8784 ( .A(n8723), .B(n8724), .Z(n8730) );
  XOR U8785 ( .A(n8731), .B(n8730), .Z(n8737) );
  XOR U8786 ( .A(n8738), .B(n8737), .Z(n8577) );
  NAND U8787 ( .A(n8546), .B(n8545), .Z(n8550) );
  NANDN U8788 ( .A(n8548), .B(n8547), .Z(n8549) );
  NAND U8789 ( .A(n8550), .B(n8549), .Z(n8574) );
  XOR U8790 ( .A(n8575), .B(n8574), .Z(n8576) );
  XOR U8791 ( .A(n8577), .B(n8576), .Z(n8568) );
  XNOR U8792 ( .A(n8569), .B(n8568), .Z(n8571) );
  XOR U8793 ( .A(n8570), .B(n8571), .Z(n8567) );
  NANDN U8794 ( .A(n8552), .B(n8551), .Z(n8556) );
  NAND U8795 ( .A(n8554), .B(n8553), .Z(n8555) );
  NAND U8796 ( .A(n8556), .B(n8555), .Z(n8566) );
  NANDN U8797 ( .A(n8557), .B(n8558), .Z(n8563) );
  NOR U8798 ( .A(n8559), .B(n8558), .Z(n8561) );
  OR U8799 ( .A(n8561), .B(n8560), .Z(n8562) );
  AND U8800 ( .A(n8563), .B(n8562), .Z(n8565) );
  XOR U8801 ( .A(n8566), .B(n8565), .Z(n8564) );
  XNOR U8802 ( .A(n8567), .B(n8564), .Z(N190) );
  NAND U8803 ( .A(n8569), .B(n8568), .Z(n8573) );
  NANDN U8804 ( .A(n8571), .B(n8570), .Z(n8572) );
  NAND U8805 ( .A(n8573), .B(n8572), .Z(n9032) );
  NANDN U8806 ( .A(n8579), .B(n8578), .Z(n8583) );
  NANDN U8807 ( .A(n8581), .B(n8580), .Z(n8582) );
  AND U8808 ( .A(n8583), .B(n8582), .Z(n9011) );
  NANDN U8809 ( .A(n8585), .B(n8584), .Z(n8589) );
  NANDN U8810 ( .A(n8587), .B(n8586), .Z(n8588) );
  AND U8811 ( .A(n8589), .B(n8588), .Z(n9004) );
  NAND U8812 ( .A(n8591), .B(n8590), .Z(n8595) );
  NAND U8813 ( .A(n8593), .B(n8592), .Z(n8594) );
  AND U8814 ( .A(n8595), .B(n8594), .Z(n8994) );
  NAND U8815 ( .A(n8597), .B(n8596), .Z(n8601) );
  NAND U8816 ( .A(n8599), .B(n8598), .Z(n8600) );
  AND U8817 ( .A(n8601), .B(n8600), .Z(n8954) );
  NAND U8818 ( .A(n8603), .B(n8602), .Z(n8607) );
  NAND U8819 ( .A(n8605), .B(n8604), .Z(n8606) );
  AND U8820 ( .A(n8607), .B(n8606), .Z(n8956) );
  AND U8821 ( .A(x[70]), .B(y[280]), .Z(n8801) );
  AND U8822 ( .A(x[69]), .B(y[281]), .Z(n8803) );
  AND U8823 ( .A(x[83]), .B(y[267]), .Z(n8802) );
  XOR U8824 ( .A(n8803), .B(n8802), .Z(n8800) );
  XOR U8825 ( .A(n8801), .B(n8800), .Z(n8784) );
  AND U8826 ( .A(x[68]), .B(y[282]), .Z(n8916) );
  AND U8827 ( .A(x[67]), .B(y[283]), .Z(n8918) );
  AND U8828 ( .A(x[82]), .B(y[268]), .Z(n8917) );
  XOR U8829 ( .A(n8918), .B(n8917), .Z(n8915) );
  XOR U8830 ( .A(n8916), .B(n8915), .Z(n8786) );
  NAND U8831 ( .A(n8609), .B(n8608), .Z(n8613) );
  NAND U8832 ( .A(n8611), .B(n8610), .Z(n8612) );
  AND U8833 ( .A(n8613), .B(n8612), .Z(n8785) );
  XOR U8834 ( .A(n8784), .B(n8783), .Z(n8955) );
  XOR U8835 ( .A(n8954), .B(n8953), .Z(n8993) );
  XOR U8836 ( .A(n8994), .B(n8993), .Z(n8991) );
  NAND U8837 ( .A(n8615), .B(n8614), .Z(n8619) );
  NAND U8838 ( .A(n8617), .B(n8616), .Z(n8618) );
  NAND U8839 ( .A(n8619), .B(n8618), .Z(n8992) );
  XOR U8840 ( .A(n8991), .B(n8992), .Z(n9005) );
  NAND U8841 ( .A(n8621), .B(n8620), .Z(n8625) );
  AND U8842 ( .A(n8623), .B(n8622), .Z(n8624) );
  ANDN U8843 ( .B(n8625), .A(n8624), .Z(n8948) );
  NAND U8844 ( .A(n8626), .B(n8921), .Z(n8630) );
  NAND U8845 ( .A(n8628), .B(n8627), .Z(n8629) );
  AND U8846 ( .A(n8630), .B(n8629), .Z(n8950) );
  NAND U8847 ( .A(n8791), .B(n8631), .Z(n8635) );
  NAND U8848 ( .A(n8633), .B(n8632), .Z(n8634) );
  AND U8849 ( .A(n8635), .B(n8634), .Z(n8764) );
  AND U8850 ( .A(n8636), .B(o[93]), .Z(n8936) );
  AND U8851 ( .A(x[92]), .B(y[258]), .Z(n8938) );
  AND U8852 ( .A(x[80]), .B(y[270]), .Z(n8937) );
  XOR U8853 ( .A(n8938), .B(n8937), .Z(n8935) );
  XOR U8854 ( .A(n8936), .B(n8935), .Z(n8766) );
  AND U8855 ( .A(x[89]), .B(y[261]), .Z(n8833) );
  AND U8856 ( .A(y[262]), .B(x[88]), .Z(n8638) );
  NAND U8857 ( .A(y[263]), .B(x[87]), .Z(n8637) );
  XNOR U8858 ( .A(n8638), .B(n8637), .Z(n8832) );
  XNOR U8859 ( .A(n8833), .B(n8832), .Z(n8765) );
  XNOR U8860 ( .A(n8764), .B(n8763), .Z(n8949) );
  XNOR U8861 ( .A(n8948), .B(n8947), .Z(n8988) );
  NAND U8862 ( .A(n8640), .B(n8639), .Z(n8643) );
  NAND U8863 ( .A(n8834), .B(n8641), .Z(n8642) );
  AND U8864 ( .A(n8643), .B(n8642), .Z(n8978) );
  NAND U8865 ( .A(n8645), .B(n8644), .Z(n8649) );
  NAND U8866 ( .A(n8647), .B(n8646), .Z(n8648) );
  AND U8867 ( .A(n8649), .B(n8648), .Z(n8829) );
  AND U8868 ( .A(x[64]), .B(y[286]), .Z(n8892) );
  NAND U8869 ( .A(x[93]), .B(y[257]), .Z(n8870) );
  NAND U8870 ( .A(x[94]), .B(y[256]), .Z(n8894) );
  XOR U8871 ( .A(n8892), .B(n8891), .Z(n8826) );
  NAND U8872 ( .A(x[84]), .B(y[266]), .Z(n8932) );
  AND U8873 ( .A(x[72]), .B(y[278]), .Z(n8929) );
  XNOR U8874 ( .A(n8930), .B(n8929), .Z(n8827) );
  XNOR U8875 ( .A(n8826), .B(n8827), .Z(n8828) );
  XNOR U8876 ( .A(n8829), .B(n8828), .Z(n8977) );
  AND U8877 ( .A(x[71]), .B(y[279]), .Z(n8790) );
  NAND U8878 ( .A(n8650), .B(n8790), .Z(n8654) );
  NAND U8879 ( .A(n8652), .B(n8651), .Z(n8653) );
  AND U8880 ( .A(n8654), .B(n8653), .Z(n8776) );
  AND U8881 ( .A(y[265]), .B(x[85]), .Z(n8656) );
  NAND U8882 ( .A(y[264]), .B(x[86]), .Z(n8655) );
  XNOR U8883 ( .A(n8656), .B(n8655), .Z(n8789) );
  XOR U8884 ( .A(n8790), .B(n8789), .Z(n8778) );
  AND U8885 ( .A(x[81]), .B(y[269]), .Z(n8795) );
  AND U8886 ( .A(x[66]), .B(y[284]), .Z(n8797) );
  AND U8887 ( .A(x[90]), .B(y[260]), .Z(n8796) );
  XOR U8888 ( .A(n8797), .B(n8796), .Z(n8794) );
  XNOR U8889 ( .A(n8795), .B(n8794), .Z(n8777) );
  XOR U8890 ( .A(n8776), .B(n8775), .Z(n8976) );
  XNOR U8891 ( .A(n8975), .B(n8976), .Z(n8989) );
  NAND U8892 ( .A(n8658), .B(n8657), .Z(n8662) );
  NAND U8893 ( .A(n8660), .B(n8659), .Z(n8661) );
  AND U8894 ( .A(n8662), .B(n8661), .Z(n8990) );
  XOR U8895 ( .A(n8988), .B(n8987), .Z(n9006) );
  XOR U8896 ( .A(n9005), .B(n9006), .Z(n9003) );
  XOR U8897 ( .A(n9004), .B(n9003), .Z(n9013) );
  NAND U8898 ( .A(n8664), .B(n8663), .Z(n8668) );
  NAND U8899 ( .A(n8666), .B(n8665), .Z(n8667) );
  AND U8900 ( .A(n8668), .B(n8667), .Z(n9012) );
  NANDN U8901 ( .A(n8670), .B(n8669), .Z(n8674) );
  NANDN U8902 ( .A(n8672), .B(n8671), .Z(n8673) );
  AND U8903 ( .A(n8674), .B(n8673), .Z(n9002) );
  NANDN U8904 ( .A(n8676), .B(n8675), .Z(n8680) );
  NANDN U8905 ( .A(n8678), .B(n8677), .Z(n8679) );
  AND U8906 ( .A(n8680), .B(n8679), .Z(n8751) );
  NAND U8907 ( .A(n8682), .B(n8681), .Z(n8686) );
  NAND U8908 ( .A(n8684), .B(n8683), .Z(n8685) );
  AND U8909 ( .A(n8686), .B(n8685), .Z(n8759) );
  NAND U8910 ( .A(n8688), .B(n8687), .Z(n8692) );
  NANDN U8911 ( .A(n8690), .B(n8689), .Z(n8691) );
  NAND U8912 ( .A(n8692), .B(n8691), .Z(n8760) );
  XNOR U8913 ( .A(n8759), .B(n8760), .Z(n8758) );
  NANDN U8914 ( .A(n8694), .B(n8693), .Z(n8698) );
  NANDN U8915 ( .A(n8696), .B(n8695), .Z(n8697) );
  NAND U8916 ( .A(n8698), .B(n8697), .Z(n8757) );
  XOR U8917 ( .A(n8758), .B(n8757), .Z(n8754) );
  NAND U8918 ( .A(n8888), .B(n8699), .Z(n8703) );
  NAND U8919 ( .A(n8701), .B(n8700), .Z(n8702) );
  AND U8920 ( .A(n8703), .B(n8702), .Z(n8971) );
  NAND U8921 ( .A(n8705), .B(n8704), .Z(n8709) );
  NAND U8922 ( .A(n8707), .B(n8706), .Z(n8708) );
  NAND U8923 ( .A(n8709), .B(n8708), .Z(n8769) );
  AND U8924 ( .A(y[274]), .B(x[76]), .Z(n8710) );
  XOR U8925 ( .A(n8711), .B(n8710), .Z(n8923) );
  XOR U8926 ( .A(n8924), .B(n8923), .Z(n8886) );
  AND U8927 ( .A(y[277]), .B(x[73]), .Z(n8712) );
  XOR U8928 ( .A(n8713), .B(n8712), .Z(n8885) );
  XOR U8929 ( .A(n8886), .B(n8885), .Z(n8772) );
  AND U8930 ( .A(x[91]), .B(y[259]), .Z(n8838) );
  AND U8931 ( .A(x[65]), .B(y[285]), .Z(n8837) );
  XOR U8932 ( .A(n8838), .B(n8837), .Z(n8839) );
  XOR U8933 ( .A(n8840), .B(n8839), .Z(n8771) );
  XOR U8934 ( .A(n8772), .B(n8771), .Z(n8770) );
  XOR U8935 ( .A(n8769), .B(n8770), .Z(n8972) );
  NAND U8936 ( .A(n8715), .B(n8714), .Z(n8719) );
  NANDN U8937 ( .A(n8717), .B(n8716), .Z(n8718) );
  AND U8938 ( .A(n8719), .B(n8718), .Z(n8969) );
  XNOR U8939 ( .A(n8970), .B(n8969), .Z(n8753) );
  XOR U8940 ( .A(n8751), .B(n8750), .Z(n9001) );
  XOR U8941 ( .A(n9000), .B(n8999), .Z(n9025) );
  IV U8942 ( .A(n8720), .Z(n8722) );
  NANDN U8943 ( .A(n8722), .B(n8721), .Z(n8727) );
  IV U8944 ( .A(n8723), .Z(n8725) );
  NANDN U8945 ( .A(n8725), .B(n8724), .Z(n8726) );
  AND U8946 ( .A(n8727), .B(n8726), .Z(n8745) );
  NANDN U8947 ( .A(n8729), .B(n8728), .Z(n8734) );
  IV U8948 ( .A(n8730), .Z(n8732) );
  NANDN U8949 ( .A(n8732), .B(n8731), .Z(n8733) );
  AND U8950 ( .A(n8734), .B(n8733), .Z(n8746) );
  NANDN U8951 ( .A(n8736), .B(n8735), .Z(n8741) );
  IV U8952 ( .A(n8737), .Z(n8739) );
  NANDN U8953 ( .A(n8739), .B(n8738), .Z(n8740) );
  NAND U8954 ( .A(n8741), .B(n8740), .Z(n8747) );
  IV U8955 ( .A(n8747), .Z(n8742) );
  XOR U8956 ( .A(n8746), .B(n8742), .Z(n8744) );
  XOR U8957 ( .A(n8745), .B(n8744), .Z(n9026) );
  IV U8958 ( .A(n9026), .Z(n8743) );
  XOR U8959 ( .A(n9025), .B(n8743), .Z(n9023) );
  XNOR U8960 ( .A(n9024), .B(n9023), .Z(n9029) );
  XNOR U8961 ( .A(n9030), .B(n9029), .Z(N191) );
  NAND U8962 ( .A(n8745), .B(n8744), .Z(n8749) );
  NANDN U8963 ( .A(n8747), .B(n8746), .Z(n8748) );
  AND U8964 ( .A(n8749), .B(n8748), .Z(n9022) );
  IV U8965 ( .A(n8750), .Z(n8752) );
  NANDN U8966 ( .A(n8752), .B(n8751), .Z(n8756) );
  NANDN U8967 ( .A(n8754), .B(n8753), .Z(n8755) );
  AND U8968 ( .A(n8756), .B(n8755), .Z(n8998) );
  NAND U8969 ( .A(n8758), .B(n8757), .Z(n8762) );
  NANDN U8970 ( .A(n8760), .B(n8759), .Z(n8761) );
  AND U8971 ( .A(n8762), .B(n8761), .Z(n8986) );
  NAND U8972 ( .A(n8764), .B(n8763), .Z(n8768) );
  NANDN U8973 ( .A(n8766), .B(n8765), .Z(n8767) );
  AND U8974 ( .A(n8768), .B(n8767), .Z(n8968) );
  NAND U8975 ( .A(n8770), .B(n8769), .Z(n8774) );
  NAND U8976 ( .A(n8772), .B(n8771), .Z(n8773) );
  AND U8977 ( .A(n8774), .B(n8773), .Z(n8782) );
  NAND U8978 ( .A(n8776), .B(n8775), .Z(n8780) );
  NANDN U8979 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U8980 ( .A(n8780), .B(n8779), .Z(n8781) );
  XNOR U8981 ( .A(n8782), .B(n8781), .Z(n8966) );
  NANDN U8982 ( .A(n8784), .B(n8783), .Z(n8788) );
  NANDN U8983 ( .A(n8786), .B(n8785), .Z(n8787) );
  AND U8984 ( .A(n8788), .B(n8787), .Z(n8964) );
  NAND U8985 ( .A(n8790), .B(n8789), .Z(n8793) );
  AND U8986 ( .A(x[86]), .B(y[265]), .Z(n8851) );
  NAND U8987 ( .A(n8791), .B(n8851), .Z(n8792) );
  AND U8988 ( .A(n8793), .B(n8792), .Z(n8825) );
  NAND U8989 ( .A(n8795), .B(n8794), .Z(n8799) );
  NAND U8990 ( .A(n8797), .B(n8796), .Z(n8798) );
  AND U8991 ( .A(n8799), .B(n8798), .Z(n8807) );
  NAND U8992 ( .A(n8801), .B(n8800), .Z(n8805) );
  NAND U8993 ( .A(n8803), .B(n8802), .Z(n8804) );
  NAND U8994 ( .A(n8805), .B(n8804), .Z(n8806) );
  XNOR U8995 ( .A(n8807), .B(n8806), .Z(n8823) );
  AND U8996 ( .A(y[275]), .B(x[76]), .Z(n8809) );
  NAND U8997 ( .A(y[287]), .B(x[64]), .Z(n8808) );
  XNOR U8998 ( .A(n8809), .B(n8808), .Z(n8813) );
  AND U8999 ( .A(y[276]), .B(x[75]), .Z(n8811) );
  NAND U9000 ( .A(y[261]), .B(x[90]), .Z(n8810) );
  XNOR U9001 ( .A(n8811), .B(n8810), .Z(n8812) );
  XOR U9002 ( .A(n8813), .B(n8812), .Z(n8821) );
  AND U9003 ( .A(y[259]), .B(x[92]), .Z(n8815) );
  NAND U9004 ( .A(y[286]), .B(x[65]), .Z(n8814) );
  XNOR U9005 ( .A(n8815), .B(n8814), .Z(n8819) );
  AND U9006 ( .A(y[256]), .B(x[95]), .Z(n8817) );
  NAND U9007 ( .A(y[283]), .B(x[68]), .Z(n8816) );
  XNOR U9008 ( .A(n8817), .B(n8816), .Z(n8818) );
  XNOR U9009 ( .A(n8819), .B(n8818), .Z(n8820) );
  XNOR U9010 ( .A(n8821), .B(n8820), .Z(n8822) );
  XNOR U9011 ( .A(n8823), .B(n8822), .Z(n8824) );
  XNOR U9012 ( .A(n8825), .B(n8824), .Z(n8914) );
  ANDN U9013 ( .B(n8827), .A(n8826), .Z(n8831) );
  AND U9014 ( .A(n8829), .B(n8828), .Z(n8830) );
  NOR U9015 ( .A(n8831), .B(n8830), .Z(n8912) );
  NAND U9016 ( .A(n8833), .B(n8832), .Z(n8836) );
  NAND U9017 ( .A(n8872), .B(n8834), .Z(n8835) );
  AND U9018 ( .A(n8836), .B(n8835), .Z(n8844) );
  NAND U9019 ( .A(n8838), .B(n8837), .Z(n8842) );
  NAND U9020 ( .A(n8840), .B(n8839), .Z(n8841) );
  AND U9021 ( .A(n8842), .B(n8841), .Z(n8843) );
  XNOR U9022 ( .A(n8844), .B(n8843), .Z(n8910) );
  AND U9023 ( .A(y[280]), .B(x[71]), .Z(n8846) );
  NAND U9024 ( .A(y[264]), .B(x[87]), .Z(n8845) );
  XNOR U9025 ( .A(n8846), .B(n8845), .Z(n8850) );
  AND U9026 ( .A(y[260]), .B(x[91]), .Z(n8848) );
  NAND U9027 ( .A(y[285]), .B(x[66]), .Z(n8847) );
  XNOR U9028 ( .A(n8848), .B(n8847), .Z(n8849) );
  XOR U9029 ( .A(n8850), .B(n8849), .Z(n8853) );
  AND U9030 ( .A(x[74]), .B(y[277]), .Z(n8887) );
  XNOR U9031 ( .A(n8851), .B(n8887), .Z(n8852) );
  XNOR U9032 ( .A(n8853), .B(n8852), .Z(n8869) );
  AND U9033 ( .A(y[267]), .B(x[84]), .Z(n8855) );
  NAND U9034 ( .A(y[278]), .B(x[73]), .Z(n8854) );
  XNOR U9035 ( .A(n8855), .B(n8854), .Z(n8859) );
  AND U9036 ( .A(y[262]), .B(x[89]), .Z(n8857) );
  NAND U9037 ( .A(y[273]), .B(x[78]), .Z(n8856) );
  XNOR U9038 ( .A(n8857), .B(n8856), .Z(n8858) );
  XOR U9039 ( .A(n8859), .B(n8858), .Z(n8867) );
  AND U9040 ( .A(y[258]), .B(x[93]), .Z(n8861) );
  NAND U9041 ( .A(y[270]), .B(x[81]), .Z(n8860) );
  XNOR U9042 ( .A(n8861), .B(n8860), .Z(n8865) );
  AND U9043 ( .A(y[257]), .B(x[94]), .Z(n8863) );
  NAND U9044 ( .A(y[271]), .B(x[80]), .Z(n8862) );
  XNOR U9045 ( .A(n8863), .B(n8862), .Z(n8864) );
  XNOR U9046 ( .A(n8865), .B(n8864), .Z(n8866) );
  XNOR U9047 ( .A(n8867), .B(n8866), .Z(n8868) );
  XOR U9048 ( .A(n8869), .B(n8868), .Z(n8884) );
  AND U9049 ( .A(y[266]), .B(x[85]), .Z(n8878) );
  ANDN U9050 ( .B(o[94]), .A(n8870), .Z(n8876) );
  XOR U9051 ( .A(n8922), .B(o[95]), .Z(n8874) );
  XNOR U9052 ( .A(n8872), .B(n8871), .Z(n8873) );
  XNOR U9053 ( .A(n8874), .B(n8873), .Z(n8875) );
  XNOR U9054 ( .A(n8876), .B(n8875), .Z(n8877) );
  XNOR U9055 ( .A(n8878), .B(n8877), .Z(n8882) );
  AND U9056 ( .A(y[281]), .B(x[70]), .Z(n8880) );
  NAND U9057 ( .A(y[282]), .B(x[69]), .Z(n8879) );
  XNOR U9058 ( .A(n8880), .B(n8879), .Z(n8881) );
  XNOR U9059 ( .A(n8882), .B(n8881), .Z(n8883) );
  XNOR U9060 ( .A(n8884), .B(n8883), .Z(n8900) );
  NAND U9061 ( .A(n8886), .B(n8885), .Z(n8890) );
  NAND U9062 ( .A(n8888), .B(n8887), .Z(n8889) );
  AND U9063 ( .A(n8890), .B(n8889), .Z(n8898) );
  NAND U9064 ( .A(n8892), .B(n8891), .Z(n8896) );
  NANDN U9065 ( .A(n8894), .B(n8893), .Z(n8895) );
  NAND U9066 ( .A(n8896), .B(n8895), .Z(n8897) );
  XNOR U9067 ( .A(n8898), .B(n8897), .Z(n8899) );
  XOR U9068 ( .A(n8900), .B(n8899), .Z(n8908) );
  AND U9069 ( .A(y[279]), .B(x[72]), .Z(n8902) );
  NAND U9070 ( .A(y[268]), .B(x[83]), .Z(n8901) );
  XNOR U9071 ( .A(n8902), .B(n8901), .Z(n8906) );
  AND U9072 ( .A(y[269]), .B(x[82]), .Z(n8904) );
  NAND U9073 ( .A(y[284]), .B(x[67]), .Z(n8903) );
  XNOR U9074 ( .A(n8904), .B(n8903), .Z(n8905) );
  XNOR U9075 ( .A(n8906), .B(n8905), .Z(n8907) );
  XNOR U9076 ( .A(n8908), .B(n8907), .Z(n8909) );
  XOR U9077 ( .A(n8910), .B(n8909), .Z(n8911) );
  XNOR U9078 ( .A(n8912), .B(n8911), .Z(n8913) );
  XOR U9079 ( .A(n8914), .B(n8913), .Z(n8946) );
  NAND U9080 ( .A(n8916), .B(n8915), .Z(n8920) );
  NAND U9081 ( .A(n8918), .B(n8917), .Z(n8919) );
  AND U9082 ( .A(n8920), .B(n8919), .Z(n8928) );
  NAND U9083 ( .A(n8922), .B(n8921), .Z(n8926) );
  NAND U9084 ( .A(n8924), .B(n8923), .Z(n8925) );
  AND U9085 ( .A(n8926), .B(n8925), .Z(n8927) );
  XNOR U9086 ( .A(n8928), .B(n8927), .Z(n8944) );
  NAND U9087 ( .A(n8930), .B(n8929), .Z(n8934) );
  NANDN U9088 ( .A(n8932), .B(n8931), .Z(n8933) );
  AND U9089 ( .A(n8934), .B(n8933), .Z(n8942) );
  NAND U9090 ( .A(n8936), .B(n8935), .Z(n8940) );
  NAND U9091 ( .A(n8938), .B(n8937), .Z(n8939) );
  NAND U9092 ( .A(n8940), .B(n8939), .Z(n8941) );
  XNOR U9093 ( .A(n8942), .B(n8941), .Z(n8943) );
  XOR U9094 ( .A(n8944), .B(n8943), .Z(n8945) );
  XNOR U9095 ( .A(n8946), .B(n8945), .Z(n8962) );
  NANDN U9096 ( .A(n8948), .B(n8947), .Z(n8952) );
  NANDN U9097 ( .A(n8950), .B(n8949), .Z(n8951) );
  AND U9098 ( .A(n8952), .B(n8951), .Z(n8960) );
  NANDN U9099 ( .A(n8954), .B(n8953), .Z(n8958) );
  NANDN U9100 ( .A(n8956), .B(n8955), .Z(n8957) );
  NAND U9101 ( .A(n8958), .B(n8957), .Z(n8959) );
  XNOR U9102 ( .A(n8960), .B(n8959), .Z(n8961) );
  XNOR U9103 ( .A(n8962), .B(n8961), .Z(n8963) );
  XNOR U9104 ( .A(n8964), .B(n8963), .Z(n8965) );
  XNOR U9105 ( .A(n8966), .B(n8965), .Z(n8967) );
  XNOR U9106 ( .A(n8968), .B(n8967), .Z(n8984) );
  NAND U9107 ( .A(n8970), .B(n8969), .Z(n8974) );
  NANDN U9108 ( .A(n8972), .B(n8971), .Z(n8973) );
  AND U9109 ( .A(n8974), .B(n8973), .Z(n8982) );
  NANDN U9110 ( .A(n8976), .B(n8975), .Z(n8980) );
  NANDN U9111 ( .A(n8978), .B(n8977), .Z(n8979) );
  NAND U9112 ( .A(n8980), .B(n8979), .Z(n8981) );
  XNOR U9113 ( .A(n8982), .B(n8981), .Z(n8983) );
  XNOR U9114 ( .A(n8984), .B(n8983), .Z(n8985) );
  XNOR U9115 ( .A(n8986), .B(n8985), .Z(n8996) );
  XNOR U9116 ( .A(n8996), .B(n8995), .Z(n8997) );
  XNOR U9117 ( .A(n8998), .B(n8997), .Z(n9020) );
  NAND U9118 ( .A(n9004), .B(n9003), .Z(n9008) );
  NAND U9119 ( .A(n9006), .B(n9005), .Z(n9007) );
  NAND U9120 ( .A(n9008), .B(n9007), .Z(n9009) );
  XNOR U9121 ( .A(n9010), .B(n9009), .Z(n9018) );
  NANDN U9122 ( .A(n9012), .B(n9011), .Z(n9016) );
  ANDN U9123 ( .B(n9012), .A(n9011), .Z(n9014) );
  NANDN U9124 ( .A(n9014), .B(n9013), .Z(n9015) );
  NAND U9125 ( .A(n9016), .B(n9015), .Z(n9017) );
  XNOR U9126 ( .A(n9018), .B(n9017), .Z(n9019) );
  XNOR U9127 ( .A(n9020), .B(n9019), .Z(n9021) );
  XNOR U9128 ( .A(n9022), .B(n9021), .Z(n9038) );
  NAND U9129 ( .A(n9024), .B(n9023), .Z(n9028) );
  NANDN U9130 ( .A(n9026), .B(n9025), .Z(n9027) );
  AND U9131 ( .A(n9028), .B(n9027), .Z(n9036) );
  NAND U9132 ( .A(n9030), .B(n9029), .Z(n9034) );
  NANDN U9133 ( .A(n9032), .B(n9031), .Z(n9033) );
  NAND U9134 ( .A(n9034), .B(n9033), .Z(n9035) );
  XNOR U9135 ( .A(n9036), .B(n9035), .Z(n9037) );
  XNOR U9136 ( .A(n9038), .B(n9037), .Z(N192) );
endmodule

