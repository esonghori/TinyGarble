
module sum_N1024_CC4 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, \ADD_/c[255] , \ADD_/c[254] , \ADD_/c[253] ,
         \ADD_/c[252] , \ADD_/c[251] , \ADD_/c[250] , \ADD_/c[249] ,
         \ADD_/c[248] , \ADD_/c[247] , \ADD_/c[246] , \ADD_/c[245] ,
         \ADD_/c[244] , \ADD_/c[243] , \ADD_/c[242] , \ADD_/c[241] ,
         \ADD_/c[240] , \ADD_/c[239] , \ADD_/c[238] , \ADD_/c[237] ,
         \ADD_/c[236] , \ADD_/c[235] , \ADD_/c[234] , \ADD_/c[233] ,
         \ADD_/c[232] , \ADD_/c[231] , \ADD_/c[230] , \ADD_/c[229] ,
         \ADD_/c[228] , \ADD_/c[227] , \ADD_/c[226] , \ADD_/c[225] ,
         \ADD_/c[224] , \ADD_/c[223] , \ADD_/c[222] , \ADD_/c[221] ,
         \ADD_/c[220] , \ADD_/c[219] , \ADD_/c[218] , \ADD_/c[217] ,
         \ADD_/c[216] , \ADD_/c[215] , \ADD_/c[214] , \ADD_/c[213] ,
         \ADD_/c[212] , \ADD_/c[211] , \ADD_/c[210] , \ADD_/c[209] ,
         \ADD_/c[208] , \ADD_/c[207] , \ADD_/c[206] , \ADD_/c[205] ,
         \ADD_/c[204] , \ADD_/c[203] , \ADD_/c[202] , \ADD_/c[201] ,
         \ADD_/c[200] , \ADD_/c[199] , \ADD_/c[198] , \ADD_/c[197] ,
         \ADD_/c[196] , \ADD_/c[195] , \ADD_/c[194] , \ADD_/c[193] ,
         \ADD_/c[192] , \ADD_/c[191] , \ADD_/c[190] , \ADD_/c[189] ,
         \ADD_/c[188] , \ADD_/c[187] , \ADD_/c[186] , \ADD_/c[185] ,
         \ADD_/c[184] , \ADD_/c[183] , \ADD_/c[182] , \ADD_/c[181] ,
         \ADD_/c[180] , \ADD_/c[179] , \ADD_/c[178] , \ADD_/c[177] ,
         \ADD_/c[176] , \ADD_/c[175] , \ADD_/c[174] , \ADD_/c[173] ,
         \ADD_/c[172] , \ADD_/c[171] , \ADD_/c[170] , \ADD_/c[169] ,
         \ADD_/c[168] , \ADD_/c[167] , \ADD_/c[166] , \ADD_/c[165] ,
         \ADD_/c[164] , \ADD_/c[163] , \ADD_/c[162] , \ADD_/c[161] ,
         \ADD_/c[160] , \ADD_/c[159] , \ADD_/c[158] , \ADD_/c[157] ,
         \ADD_/c[156] , \ADD_/c[155] , \ADD_/c[154] , \ADD_/c[153] ,
         \ADD_/c[152] , \ADD_/c[151] , \ADD_/c[150] , \ADD_/c[149] ,
         \ADD_/c[148] , \ADD_/c[147] , \ADD_/c[146] , \ADD_/c[145] ,
         \ADD_/c[144] , \ADD_/c[143] , \ADD_/c[142] , \ADD_/c[141] ,
         \ADD_/c[140] , \ADD_/c[139] , \ADD_/c[138] , \ADD_/c[137] ,
         \ADD_/c[136] , \ADD_/c[135] , \ADD_/c[134] , \ADD_/c[133] ,
         \ADD_/c[132] , \ADD_/c[131] , \ADD_/c[130] , \ADD_/c[129] ,
         \ADD_/c[128] , \ADD_/c[127] , \ADD_/c[126] , \ADD_/c[125] ,
         \ADD_/c[124] , \ADD_/c[123] , \ADD_/c[122] , \ADD_/c[121] ,
         \ADD_/c[120] , \ADD_/c[119] , \ADD_/c[118] , \ADD_/c[117] ,
         \ADD_/c[116] , \ADD_/c[115] , \ADD_/c[114] , \ADD_/c[113] ,
         \ADD_/c[112] , \ADD_/c[111] , \ADD_/c[110] , \ADD_/c[109] ,
         \ADD_/c[108] , \ADD_/c[107] , \ADD_/c[106] , \ADD_/c[105] ,
         \ADD_/c[104] , \ADD_/c[103] , \ADD_/c[102] , \ADD_/c[101] ,
         \ADD_/c[100] , \ADD_/c[99] , \ADD_/c[98] , \ADD_/c[97] , \ADD_/c[96] ,
         \ADD_/c[95] , \ADD_/c[94] , \ADD_/c[93] , \ADD_/c[92] , \ADD_/c[91] ,
         \ADD_/c[90] , \ADD_/c[89] , \ADD_/c[88] , \ADD_/c[87] , \ADD_/c[86] ,
         \ADD_/c[85] , \ADD_/c[84] , \ADD_/c[83] , \ADD_/c[82] , \ADD_/c[81] ,
         \ADD_/c[80] , \ADD_/c[79] , \ADD_/c[78] , \ADD_/c[77] , \ADD_/c[76] ,
         \ADD_/c[75] , \ADD_/c[74] , \ADD_/c[73] , \ADD_/c[72] , \ADD_/c[71] ,
         \ADD_/c[70] , \ADD_/c[69] , \ADD_/c[68] , \ADD_/c[67] , \ADD_/c[66] ,
         \ADD_/c[65] , \ADD_/c[64] , \ADD_/c[63] , \ADD_/c[62] , \ADD_/c[61] ,
         \ADD_/c[60] , \ADD_/c[59] , \ADD_/c[58] , \ADD_/c[57] , \ADD_/c[56] ,
         \ADD_/c[55] , \ADD_/c[54] , \ADD_/c[53] , \ADD_/c[52] , \ADD_/c[51] ,
         \ADD_/c[50] , \ADD_/c[49] , \ADD_/c[48] , \ADD_/c[47] , \ADD_/c[46] ,
         \ADD_/c[45] , \ADD_/c[44] , \ADD_/c[43] , \ADD_/c[42] , \ADD_/c[41] ,
         \ADD_/c[40] , \ADD_/c[39] , \ADD_/c[38] , \ADD_/c[37] , \ADD_/c[36] ,
         \ADD_/c[35] , \ADD_/c[34] , \ADD_/c[33] , \ADD_/c[32] , \ADD_/c[31] ,
         \ADD_/c[30] , \ADD_/c[29] , \ADD_/c[28] , \ADD_/c[27] , \ADD_/c[26] ,
         \ADD_/c[25] , \ADD_/c[24] , \ADD_/c[23] , \ADD_/c[22] , \ADD_/c[21] ,
         \ADD_/c[20] , \ADD_/c[19] , \ADD_/c[18] , \ADD_/c[17] , \ADD_/c[16] ,
         \ADD_/c[15] , \ADD_/c[14] , \ADD_/c[13] , \ADD_/c[12] , \ADD_/c[11] ,
         \ADD_/c[10] , \ADD_/c[9] , \ADD_/c[8] , \ADD_/c[7] , \ADD_/c[6] ,
         \ADD_/c[5] , \ADD_/c[4] , \ADD_/c[3] , \ADD_/c[2] , \ADD_/c[1] ,
         \ADD_/FAINST[0].FA_/n3 , \ADD_/FAINST[0].FA_/n2 ,
         \ADD_/FAINST[0].FA_/n1 , \ADD_/FAINST[255].FA_/n3 ,
         \ADD_/FAINST[255].FA_/n2 , \ADD_/FAINST[255].FA_/n1 ,
         \ADD_/FAINST[254].FA_/n3 , \ADD_/FAINST[254].FA_/n2 ,
         \ADD_/FAINST[254].FA_/n1 , \ADD_/FAINST[253].FA_/n3 ,
         \ADD_/FAINST[253].FA_/n2 , \ADD_/FAINST[253].FA_/n1 ,
         \ADD_/FAINST[252].FA_/n3 , \ADD_/FAINST[252].FA_/n2 ,
         \ADD_/FAINST[252].FA_/n1 , \ADD_/FAINST[251].FA_/n3 ,
         \ADD_/FAINST[251].FA_/n2 , \ADD_/FAINST[251].FA_/n1 ,
         \ADD_/FAINST[250].FA_/n3 , \ADD_/FAINST[250].FA_/n2 ,
         \ADD_/FAINST[250].FA_/n1 , \ADD_/FAINST[249].FA_/n3 ,
         \ADD_/FAINST[249].FA_/n2 , \ADD_/FAINST[249].FA_/n1 ,
         \ADD_/FAINST[248].FA_/n3 , \ADD_/FAINST[248].FA_/n2 ,
         \ADD_/FAINST[248].FA_/n1 , \ADD_/FAINST[247].FA_/n3 ,
         \ADD_/FAINST[247].FA_/n2 , \ADD_/FAINST[247].FA_/n1 ,
         \ADD_/FAINST[246].FA_/n3 , \ADD_/FAINST[246].FA_/n2 ,
         \ADD_/FAINST[246].FA_/n1 , \ADD_/FAINST[245].FA_/n3 ,
         \ADD_/FAINST[245].FA_/n2 , \ADD_/FAINST[245].FA_/n1 ,
         \ADD_/FAINST[244].FA_/n3 , \ADD_/FAINST[244].FA_/n2 ,
         \ADD_/FAINST[244].FA_/n1 , \ADD_/FAINST[243].FA_/n3 ,
         \ADD_/FAINST[243].FA_/n2 , \ADD_/FAINST[243].FA_/n1 ,
         \ADD_/FAINST[242].FA_/n3 , \ADD_/FAINST[242].FA_/n2 ,
         \ADD_/FAINST[242].FA_/n1 , \ADD_/FAINST[241].FA_/n3 ,
         \ADD_/FAINST[241].FA_/n2 , \ADD_/FAINST[241].FA_/n1 ,
         \ADD_/FAINST[240].FA_/n3 , \ADD_/FAINST[240].FA_/n2 ,
         \ADD_/FAINST[240].FA_/n1 , \ADD_/FAINST[239].FA_/n3 ,
         \ADD_/FAINST[239].FA_/n2 , \ADD_/FAINST[239].FA_/n1 ,
         \ADD_/FAINST[238].FA_/n3 , \ADD_/FAINST[238].FA_/n2 ,
         \ADD_/FAINST[238].FA_/n1 , \ADD_/FAINST[237].FA_/n3 ,
         \ADD_/FAINST[237].FA_/n2 , \ADD_/FAINST[237].FA_/n1 ,
         \ADD_/FAINST[236].FA_/n3 , \ADD_/FAINST[236].FA_/n2 ,
         \ADD_/FAINST[236].FA_/n1 , \ADD_/FAINST[235].FA_/n3 ,
         \ADD_/FAINST[235].FA_/n2 , \ADD_/FAINST[235].FA_/n1 ,
         \ADD_/FAINST[234].FA_/n3 , \ADD_/FAINST[234].FA_/n2 ,
         \ADD_/FAINST[234].FA_/n1 , \ADD_/FAINST[233].FA_/n3 ,
         \ADD_/FAINST[233].FA_/n2 , \ADD_/FAINST[233].FA_/n1 ,
         \ADD_/FAINST[232].FA_/n3 , \ADD_/FAINST[232].FA_/n2 ,
         \ADD_/FAINST[232].FA_/n1 , \ADD_/FAINST[231].FA_/n3 ,
         \ADD_/FAINST[231].FA_/n2 , \ADD_/FAINST[231].FA_/n1 ,
         \ADD_/FAINST[230].FA_/n3 , \ADD_/FAINST[230].FA_/n2 ,
         \ADD_/FAINST[230].FA_/n1 , \ADD_/FAINST[229].FA_/n3 ,
         \ADD_/FAINST[229].FA_/n2 , \ADD_/FAINST[229].FA_/n1 ,
         \ADD_/FAINST[228].FA_/n3 , \ADD_/FAINST[228].FA_/n2 ,
         \ADD_/FAINST[228].FA_/n1 , \ADD_/FAINST[227].FA_/n3 ,
         \ADD_/FAINST[227].FA_/n2 , \ADD_/FAINST[227].FA_/n1 ,
         \ADD_/FAINST[226].FA_/n3 , \ADD_/FAINST[226].FA_/n2 ,
         \ADD_/FAINST[226].FA_/n1 , \ADD_/FAINST[225].FA_/n3 ,
         \ADD_/FAINST[225].FA_/n2 , \ADD_/FAINST[225].FA_/n1 ,
         \ADD_/FAINST[224].FA_/n3 , \ADD_/FAINST[224].FA_/n2 ,
         \ADD_/FAINST[224].FA_/n1 , \ADD_/FAINST[223].FA_/n3 ,
         \ADD_/FAINST[223].FA_/n2 , \ADD_/FAINST[223].FA_/n1 ,
         \ADD_/FAINST[222].FA_/n3 , \ADD_/FAINST[222].FA_/n2 ,
         \ADD_/FAINST[222].FA_/n1 , \ADD_/FAINST[221].FA_/n3 ,
         \ADD_/FAINST[221].FA_/n2 , \ADD_/FAINST[221].FA_/n1 ,
         \ADD_/FAINST[220].FA_/n3 , \ADD_/FAINST[220].FA_/n2 ,
         \ADD_/FAINST[220].FA_/n1 , \ADD_/FAINST[219].FA_/n3 ,
         \ADD_/FAINST[219].FA_/n2 , \ADD_/FAINST[219].FA_/n1 ,
         \ADD_/FAINST[218].FA_/n3 , \ADD_/FAINST[218].FA_/n2 ,
         \ADD_/FAINST[218].FA_/n1 , \ADD_/FAINST[217].FA_/n3 ,
         \ADD_/FAINST[217].FA_/n2 , \ADD_/FAINST[217].FA_/n1 ,
         \ADD_/FAINST[216].FA_/n3 , \ADD_/FAINST[216].FA_/n2 ,
         \ADD_/FAINST[216].FA_/n1 , \ADD_/FAINST[215].FA_/n3 ,
         \ADD_/FAINST[215].FA_/n2 , \ADD_/FAINST[215].FA_/n1 ,
         \ADD_/FAINST[214].FA_/n3 , \ADD_/FAINST[214].FA_/n2 ,
         \ADD_/FAINST[214].FA_/n1 , \ADD_/FAINST[213].FA_/n3 ,
         \ADD_/FAINST[213].FA_/n2 , \ADD_/FAINST[213].FA_/n1 ,
         \ADD_/FAINST[212].FA_/n3 , \ADD_/FAINST[212].FA_/n2 ,
         \ADD_/FAINST[212].FA_/n1 , \ADD_/FAINST[211].FA_/n3 ,
         \ADD_/FAINST[211].FA_/n2 , \ADD_/FAINST[211].FA_/n1 ,
         \ADD_/FAINST[210].FA_/n3 , \ADD_/FAINST[210].FA_/n2 ,
         \ADD_/FAINST[210].FA_/n1 , \ADD_/FAINST[209].FA_/n3 ,
         \ADD_/FAINST[209].FA_/n2 , \ADD_/FAINST[209].FA_/n1 ,
         \ADD_/FAINST[208].FA_/n3 , \ADD_/FAINST[208].FA_/n2 ,
         \ADD_/FAINST[208].FA_/n1 , \ADD_/FAINST[207].FA_/n3 ,
         \ADD_/FAINST[207].FA_/n2 , \ADD_/FAINST[207].FA_/n1 ,
         \ADD_/FAINST[206].FA_/n3 , \ADD_/FAINST[206].FA_/n2 ,
         \ADD_/FAINST[206].FA_/n1 , \ADD_/FAINST[205].FA_/n3 ,
         \ADD_/FAINST[205].FA_/n2 , \ADD_/FAINST[205].FA_/n1 ,
         \ADD_/FAINST[204].FA_/n3 , \ADD_/FAINST[204].FA_/n2 ,
         \ADD_/FAINST[204].FA_/n1 , \ADD_/FAINST[203].FA_/n3 ,
         \ADD_/FAINST[203].FA_/n2 , \ADD_/FAINST[203].FA_/n1 ,
         \ADD_/FAINST[202].FA_/n3 , \ADD_/FAINST[202].FA_/n2 ,
         \ADD_/FAINST[202].FA_/n1 , \ADD_/FAINST[201].FA_/n3 ,
         \ADD_/FAINST[201].FA_/n2 , \ADD_/FAINST[201].FA_/n1 ,
         \ADD_/FAINST[200].FA_/n3 , \ADD_/FAINST[200].FA_/n2 ,
         \ADD_/FAINST[200].FA_/n1 , \ADD_/FAINST[199].FA_/n3 ,
         \ADD_/FAINST[199].FA_/n2 , \ADD_/FAINST[199].FA_/n1 ,
         \ADD_/FAINST[198].FA_/n3 , \ADD_/FAINST[198].FA_/n2 ,
         \ADD_/FAINST[198].FA_/n1 , \ADD_/FAINST[197].FA_/n3 ,
         \ADD_/FAINST[197].FA_/n2 , \ADD_/FAINST[197].FA_/n1 ,
         \ADD_/FAINST[196].FA_/n3 , \ADD_/FAINST[196].FA_/n2 ,
         \ADD_/FAINST[196].FA_/n1 , \ADD_/FAINST[195].FA_/n3 ,
         \ADD_/FAINST[195].FA_/n2 , \ADD_/FAINST[195].FA_/n1 ,
         \ADD_/FAINST[194].FA_/n3 , \ADD_/FAINST[194].FA_/n2 ,
         \ADD_/FAINST[194].FA_/n1 , \ADD_/FAINST[193].FA_/n3 ,
         \ADD_/FAINST[193].FA_/n2 , \ADD_/FAINST[193].FA_/n1 ,
         \ADD_/FAINST[192].FA_/n3 , \ADD_/FAINST[192].FA_/n2 ,
         \ADD_/FAINST[192].FA_/n1 , \ADD_/FAINST[191].FA_/n3 ,
         \ADD_/FAINST[191].FA_/n2 , \ADD_/FAINST[191].FA_/n1 ,
         \ADD_/FAINST[190].FA_/n3 , \ADD_/FAINST[190].FA_/n2 ,
         \ADD_/FAINST[190].FA_/n1 , \ADD_/FAINST[189].FA_/n3 ,
         \ADD_/FAINST[189].FA_/n2 , \ADD_/FAINST[189].FA_/n1 ,
         \ADD_/FAINST[188].FA_/n3 , \ADD_/FAINST[188].FA_/n2 ,
         \ADD_/FAINST[188].FA_/n1 , \ADD_/FAINST[187].FA_/n3 ,
         \ADD_/FAINST[187].FA_/n2 , \ADD_/FAINST[187].FA_/n1 ,
         \ADD_/FAINST[186].FA_/n3 , \ADD_/FAINST[186].FA_/n2 ,
         \ADD_/FAINST[186].FA_/n1 , \ADD_/FAINST[185].FA_/n3 ,
         \ADD_/FAINST[185].FA_/n2 , \ADD_/FAINST[185].FA_/n1 ,
         \ADD_/FAINST[184].FA_/n3 , \ADD_/FAINST[184].FA_/n2 ,
         \ADD_/FAINST[184].FA_/n1 , \ADD_/FAINST[183].FA_/n3 ,
         \ADD_/FAINST[183].FA_/n2 , \ADD_/FAINST[183].FA_/n1 ,
         \ADD_/FAINST[182].FA_/n3 , \ADD_/FAINST[182].FA_/n2 ,
         \ADD_/FAINST[182].FA_/n1 , \ADD_/FAINST[181].FA_/n3 ,
         \ADD_/FAINST[181].FA_/n2 , \ADD_/FAINST[181].FA_/n1 ,
         \ADD_/FAINST[180].FA_/n3 , \ADD_/FAINST[180].FA_/n2 ,
         \ADD_/FAINST[180].FA_/n1 , \ADD_/FAINST[179].FA_/n3 ,
         \ADD_/FAINST[179].FA_/n2 , \ADD_/FAINST[179].FA_/n1 ,
         \ADD_/FAINST[178].FA_/n3 , \ADD_/FAINST[178].FA_/n2 ,
         \ADD_/FAINST[178].FA_/n1 , \ADD_/FAINST[177].FA_/n3 ,
         \ADD_/FAINST[177].FA_/n2 , \ADD_/FAINST[177].FA_/n1 ,
         \ADD_/FAINST[176].FA_/n3 , \ADD_/FAINST[176].FA_/n2 ,
         \ADD_/FAINST[176].FA_/n1 , \ADD_/FAINST[175].FA_/n3 ,
         \ADD_/FAINST[175].FA_/n2 , \ADD_/FAINST[175].FA_/n1 ,
         \ADD_/FAINST[174].FA_/n3 , \ADD_/FAINST[174].FA_/n2 ,
         \ADD_/FAINST[174].FA_/n1 , \ADD_/FAINST[173].FA_/n3 ,
         \ADD_/FAINST[173].FA_/n2 , \ADD_/FAINST[173].FA_/n1 ,
         \ADD_/FAINST[172].FA_/n3 , \ADD_/FAINST[172].FA_/n2 ,
         \ADD_/FAINST[172].FA_/n1 , \ADD_/FAINST[171].FA_/n3 ,
         \ADD_/FAINST[171].FA_/n2 , \ADD_/FAINST[171].FA_/n1 ,
         \ADD_/FAINST[170].FA_/n3 , \ADD_/FAINST[170].FA_/n2 ,
         \ADD_/FAINST[170].FA_/n1 , \ADD_/FAINST[169].FA_/n3 ,
         \ADD_/FAINST[169].FA_/n2 , \ADD_/FAINST[169].FA_/n1 ,
         \ADD_/FAINST[168].FA_/n3 , \ADD_/FAINST[168].FA_/n2 ,
         \ADD_/FAINST[168].FA_/n1 , \ADD_/FAINST[167].FA_/n3 ,
         \ADD_/FAINST[167].FA_/n2 , \ADD_/FAINST[167].FA_/n1 ,
         \ADD_/FAINST[166].FA_/n3 , \ADD_/FAINST[166].FA_/n2 ,
         \ADD_/FAINST[166].FA_/n1 , \ADD_/FAINST[165].FA_/n3 ,
         \ADD_/FAINST[165].FA_/n2 , \ADD_/FAINST[165].FA_/n1 ,
         \ADD_/FAINST[164].FA_/n3 , \ADD_/FAINST[164].FA_/n2 ,
         \ADD_/FAINST[164].FA_/n1 , \ADD_/FAINST[163].FA_/n3 ,
         \ADD_/FAINST[163].FA_/n2 , \ADD_/FAINST[163].FA_/n1 ,
         \ADD_/FAINST[162].FA_/n3 , \ADD_/FAINST[162].FA_/n2 ,
         \ADD_/FAINST[162].FA_/n1 , \ADD_/FAINST[161].FA_/n3 ,
         \ADD_/FAINST[161].FA_/n2 , \ADD_/FAINST[161].FA_/n1 ,
         \ADD_/FAINST[160].FA_/n3 , \ADD_/FAINST[160].FA_/n2 ,
         \ADD_/FAINST[160].FA_/n1 , \ADD_/FAINST[159].FA_/n3 ,
         \ADD_/FAINST[159].FA_/n2 , \ADD_/FAINST[159].FA_/n1 ,
         \ADD_/FAINST[158].FA_/n3 , \ADD_/FAINST[158].FA_/n2 ,
         \ADD_/FAINST[158].FA_/n1 , \ADD_/FAINST[157].FA_/n3 ,
         \ADD_/FAINST[157].FA_/n2 , \ADD_/FAINST[157].FA_/n1 ,
         \ADD_/FAINST[156].FA_/n3 , \ADD_/FAINST[156].FA_/n2 ,
         \ADD_/FAINST[156].FA_/n1 , \ADD_/FAINST[155].FA_/n3 ,
         \ADD_/FAINST[155].FA_/n2 , \ADD_/FAINST[155].FA_/n1 ,
         \ADD_/FAINST[154].FA_/n3 , \ADD_/FAINST[154].FA_/n2 ,
         \ADD_/FAINST[154].FA_/n1 , \ADD_/FAINST[153].FA_/n3 ,
         \ADD_/FAINST[153].FA_/n2 , \ADD_/FAINST[153].FA_/n1 ,
         \ADD_/FAINST[152].FA_/n3 , \ADD_/FAINST[152].FA_/n2 ,
         \ADD_/FAINST[152].FA_/n1 , \ADD_/FAINST[151].FA_/n3 ,
         \ADD_/FAINST[151].FA_/n2 , \ADD_/FAINST[151].FA_/n1 ,
         \ADD_/FAINST[150].FA_/n3 , \ADD_/FAINST[150].FA_/n2 ,
         \ADD_/FAINST[150].FA_/n1 , \ADD_/FAINST[149].FA_/n3 ,
         \ADD_/FAINST[149].FA_/n2 , \ADD_/FAINST[149].FA_/n1 ,
         \ADD_/FAINST[148].FA_/n3 , \ADD_/FAINST[148].FA_/n2 ,
         \ADD_/FAINST[148].FA_/n1 , \ADD_/FAINST[147].FA_/n3 ,
         \ADD_/FAINST[147].FA_/n2 , \ADD_/FAINST[147].FA_/n1 ,
         \ADD_/FAINST[146].FA_/n3 , \ADD_/FAINST[146].FA_/n2 ,
         \ADD_/FAINST[146].FA_/n1 , \ADD_/FAINST[145].FA_/n3 ,
         \ADD_/FAINST[145].FA_/n2 , \ADD_/FAINST[145].FA_/n1 ,
         \ADD_/FAINST[144].FA_/n3 , \ADD_/FAINST[144].FA_/n2 ,
         \ADD_/FAINST[144].FA_/n1 , \ADD_/FAINST[143].FA_/n3 ,
         \ADD_/FAINST[143].FA_/n2 , \ADD_/FAINST[143].FA_/n1 ,
         \ADD_/FAINST[142].FA_/n3 , \ADD_/FAINST[142].FA_/n2 ,
         \ADD_/FAINST[142].FA_/n1 , \ADD_/FAINST[141].FA_/n3 ,
         \ADD_/FAINST[141].FA_/n2 , \ADD_/FAINST[141].FA_/n1 ,
         \ADD_/FAINST[140].FA_/n3 , \ADD_/FAINST[140].FA_/n2 ,
         \ADD_/FAINST[140].FA_/n1 , \ADD_/FAINST[139].FA_/n3 ,
         \ADD_/FAINST[139].FA_/n2 , \ADD_/FAINST[139].FA_/n1 ,
         \ADD_/FAINST[138].FA_/n3 , \ADD_/FAINST[138].FA_/n2 ,
         \ADD_/FAINST[138].FA_/n1 , \ADD_/FAINST[137].FA_/n3 ,
         \ADD_/FAINST[137].FA_/n2 , \ADD_/FAINST[137].FA_/n1 ,
         \ADD_/FAINST[136].FA_/n3 , \ADD_/FAINST[136].FA_/n2 ,
         \ADD_/FAINST[136].FA_/n1 , \ADD_/FAINST[135].FA_/n3 ,
         \ADD_/FAINST[135].FA_/n2 , \ADD_/FAINST[135].FA_/n1 ,
         \ADD_/FAINST[134].FA_/n3 , \ADD_/FAINST[134].FA_/n2 ,
         \ADD_/FAINST[134].FA_/n1 , \ADD_/FAINST[133].FA_/n3 ,
         \ADD_/FAINST[133].FA_/n2 , \ADD_/FAINST[133].FA_/n1 ,
         \ADD_/FAINST[132].FA_/n3 , \ADD_/FAINST[132].FA_/n2 ,
         \ADD_/FAINST[132].FA_/n1 , \ADD_/FAINST[131].FA_/n3 ,
         \ADD_/FAINST[131].FA_/n2 , \ADD_/FAINST[131].FA_/n1 ,
         \ADD_/FAINST[130].FA_/n3 , \ADD_/FAINST[130].FA_/n2 ,
         \ADD_/FAINST[130].FA_/n1 , \ADD_/FAINST[129].FA_/n3 ,
         \ADD_/FAINST[129].FA_/n2 , \ADD_/FAINST[129].FA_/n1 ,
         \ADD_/FAINST[128].FA_/n3 , \ADD_/FAINST[128].FA_/n2 ,
         \ADD_/FAINST[128].FA_/n1 , \ADD_/FAINST[127].FA_/n3 ,
         \ADD_/FAINST[127].FA_/n2 , \ADD_/FAINST[127].FA_/n1 ,
         \ADD_/FAINST[126].FA_/n3 , \ADD_/FAINST[126].FA_/n2 ,
         \ADD_/FAINST[126].FA_/n1 , \ADD_/FAINST[125].FA_/n3 ,
         \ADD_/FAINST[125].FA_/n2 , \ADD_/FAINST[125].FA_/n1 ,
         \ADD_/FAINST[124].FA_/n3 , \ADD_/FAINST[124].FA_/n2 ,
         \ADD_/FAINST[124].FA_/n1 , \ADD_/FAINST[123].FA_/n3 ,
         \ADD_/FAINST[123].FA_/n2 , \ADD_/FAINST[123].FA_/n1 ,
         \ADD_/FAINST[122].FA_/n3 , \ADD_/FAINST[122].FA_/n2 ,
         \ADD_/FAINST[122].FA_/n1 , \ADD_/FAINST[121].FA_/n3 ,
         \ADD_/FAINST[121].FA_/n2 , \ADD_/FAINST[121].FA_/n1 ,
         \ADD_/FAINST[120].FA_/n3 , \ADD_/FAINST[120].FA_/n2 ,
         \ADD_/FAINST[120].FA_/n1 , \ADD_/FAINST[119].FA_/n3 ,
         \ADD_/FAINST[119].FA_/n2 , \ADD_/FAINST[119].FA_/n1 ,
         \ADD_/FAINST[118].FA_/n3 , \ADD_/FAINST[118].FA_/n2 ,
         \ADD_/FAINST[118].FA_/n1 , \ADD_/FAINST[117].FA_/n3 ,
         \ADD_/FAINST[117].FA_/n2 , \ADD_/FAINST[117].FA_/n1 ,
         \ADD_/FAINST[116].FA_/n3 , \ADD_/FAINST[116].FA_/n2 ,
         \ADD_/FAINST[116].FA_/n1 , \ADD_/FAINST[115].FA_/n3 ,
         \ADD_/FAINST[115].FA_/n2 , \ADD_/FAINST[115].FA_/n1 ,
         \ADD_/FAINST[114].FA_/n3 , \ADD_/FAINST[114].FA_/n2 ,
         \ADD_/FAINST[114].FA_/n1 , \ADD_/FAINST[113].FA_/n3 ,
         \ADD_/FAINST[113].FA_/n2 , \ADD_/FAINST[113].FA_/n1 ,
         \ADD_/FAINST[112].FA_/n3 , \ADD_/FAINST[112].FA_/n2 ,
         \ADD_/FAINST[112].FA_/n1 , \ADD_/FAINST[111].FA_/n3 ,
         \ADD_/FAINST[111].FA_/n2 , \ADD_/FAINST[111].FA_/n1 ,
         \ADD_/FAINST[110].FA_/n3 , \ADD_/FAINST[110].FA_/n2 ,
         \ADD_/FAINST[110].FA_/n1 , \ADD_/FAINST[109].FA_/n3 ,
         \ADD_/FAINST[109].FA_/n2 , \ADD_/FAINST[109].FA_/n1 ,
         \ADD_/FAINST[108].FA_/n3 , \ADD_/FAINST[108].FA_/n2 ,
         \ADD_/FAINST[108].FA_/n1 , \ADD_/FAINST[107].FA_/n3 ,
         \ADD_/FAINST[107].FA_/n2 , \ADD_/FAINST[107].FA_/n1 ,
         \ADD_/FAINST[106].FA_/n3 , \ADD_/FAINST[106].FA_/n2 ,
         \ADD_/FAINST[106].FA_/n1 , \ADD_/FAINST[105].FA_/n3 ,
         \ADD_/FAINST[105].FA_/n2 , \ADD_/FAINST[105].FA_/n1 ,
         \ADD_/FAINST[104].FA_/n3 , \ADD_/FAINST[104].FA_/n2 ,
         \ADD_/FAINST[104].FA_/n1 , \ADD_/FAINST[103].FA_/n3 ,
         \ADD_/FAINST[103].FA_/n2 , \ADD_/FAINST[103].FA_/n1 ,
         \ADD_/FAINST[102].FA_/n3 , \ADD_/FAINST[102].FA_/n2 ,
         \ADD_/FAINST[102].FA_/n1 , \ADD_/FAINST[101].FA_/n3 ,
         \ADD_/FAINST[101].FA_/n2 , \ADD_/FAINST[101].FA_/n1 ,
         \ADD_/FAINST[100].FA_/n3 , \ADD_/FAINST[100].FA_/n2 ,
         \ADD_/FAINST[100].FA_/n1 , \ADD_/FAINST[99].FA_/n3 ,
         \ADD_/FAINST[99].FA_/n2 , \ADD_/FAINST[99].FA_/n1 ,
         \ADD_/FAINST[98].FA_/n3 , \ADD_/FAINST[98].FA_/n2 ,
         \ADD_/FAINST[98].FA_/n1 , \ADD_/FAINST[97].FA_/n3 ,
         \ADD_/FAINST[97].FA_/n2 , \ADD_/FAINST[97].FA_/n1 ,
         \ADD_/FAINST[96].FA_/n3 , \ADD_/FAINST[96].FA_/n2 ,
         \ADD_/FAINST[96].FA_/n1 , \ADD_/FAINST[95].FA_/n3 ,
         \ADD_/FAINST[95].FA_/n2 , \ADD_/FAINST[95].FA_/n1 ,
         \ADD_/FAINST[94].FA_/n3 , \ADD_/FAINST[94].FA_/n2 ,
         \ADD_/FAINST[94].FA_/n1 , \ADD_/FAINST[93].FA_/n3 ,
         \ADD_/FAINST[93].FA_/n2 , \ADD_/FAINST[93].FA_/n1 ,
         \ADD_/FAINST[92].FA_/n3 , \ADD_/FAINST[92].FA_/n2 ,
         \ADD_/FAINST[92].FA_/n1 , \ADD_/FAINST[91].FA_/n3 ,
         \ADD_/FAINST[91].FA_/n2 , \ADD_/FAINST[91].FA_/n1 ,
         \ADD_/FAINST[90].FA_/n3 , \ADD_/FAINST[90].FA_/n2 ,
         \ADD_/FAINST[90].FA_/n1 , \ADD_/FAINST[89].FA_/n3 ,
         \ADD_/FAINST[89].FA_/n2 , \ADD_/FAINST[89].FA_/n1 ,
         \ADD_/FAINST[88].FA_/n3 , \ADD_/FAINST[88].FA_/n2 ,
         \ADD_/FAINST[88].FA_/n1 , \ADD_/FAINST[87].FA_/n3 ,
         \ADD_/FAINST[87].FA_/n2 , \ADD_/FAINST[87].FA_/n1 ,
         \ADD_/FAINST[86].FA_/n3 , \ADD_/FAINST[86].FA_/n2 ,
         \ADD_/FAINST[86].FA_/n1 , \ADD_/FAINST[85].FA_/n3 ,
         \ADD_/FAINST[85].FA_/n2 , \ADD_/FAINST[85].FA_/n1 ,
         \ADD_/FAINST[84].FA_/n3 , \ADD_/FAINST[84].FA_/n2 ,
         \ADD_/FAINST[84].FA_/n1 , \ADD_/FAINST[83].FA_/n3 ,
         \ADD_/FAINST[83].FA_/n2 , \ADD_/FAINST[83].FA_/n1 ,
         \ADD_/FAINST[82].FA_/n3 , \ADD_/FAINST[82].FA_/n2 ,
         \ADD_/FAINST[82].FA_/n1 , \ADD_/FAINST[81].FA_/n3 ,
         \ADD_/FAINST[81].FA_/n2 , \ADD_/FAINST[81].FA_/n1 ,
         \ADD_/FAINST[80].FA_/n3 , \ADD_/FAINST[80].FA_/n2 ,
         \ADD_/FAINST[80].FA_/n1 , \ADD_/FAINST[79].FA_/n3 ,
         \ADD_/FAINST[79].FA_/n2 , \ADD_/FAINST[79].FA_/n1 ,
         \ADD_/FAINST[78].FA_/n3 , \ADD_/FAINST[78].FA_/n2 ,
         \ADD_/FAINST[78].FA_/n1 , \ADD_/FAINST[77].FA_/n3 ,
         \ADD_/FAINST[77].FA_/n2 , \ADD_/FAINST[77].FA_/n1 ,
         \ADD_/FAINST[76].FA_/n3 , \ADD_/FAINST[76].FA_/n2 ,
         \ADD_/FAINST[76].FA_/n1 , \ADD_/FAINST[75].FA_/n3 ,
         \ADD_/FAINST[75].FA_/n2 , \ADD_/FAINST[75].FA_/n1 ,
         \ADD_/FAINST[74].FA_/n3 , \ADD_/FAINST[74].FA_/n2 ,
         \ADD_/FAINST[74].FA_/n1 , \ADD_/FAINST[73].FA_/n3 ,
         \ADD_/FAINST[73].FA_/n2 , \ADD_/FAINST[73].FA_/n1 ,
         \ADD_/FAINST[72].FA_/n3 , \ADD_/FAINST[72].FA_/n2 ,
         \ADD_/FAINST[72].FA_/n1 , \ADD_/FAINST[71].FA_/n3 ,
         \ADD_/FAINST[71].FA_/n2 , \ADD_/FAINST[71].FA_/n1 ,
         \ADD_/FAINST[70].FA_/n3 , \ADD_/FAINST[70].FA_/n2 ,
         \ADD_/FAINST[70].FA_/n1 , \ADD_/FAINST[69].FA_/n3 ,
         \ADD_/FAINST[69].FA_/n2 , \ADD_/FAINST[69].FA_/n1 ,
         \ADD_/FAINST[68].FA_/n3 , \ADD_/FAINST[68].FA_/n2 ,
         \ADD_/FAINST[68].FA_/n1 , \ADD_/FAINST[67].FA_/n3 ,
         \ADD_/FAINST[67].FA_/n2 , \ADD_/FAINST[67].FA_/n1 ,
         \ADD_/FAINST[66].FA_/n3 , \ADD_/FAINST[66].FA_/n2 ,
         \ADD_/FAINST[66].FA_/n1 , \ADD_/FAINST[65].FA_/n3 ,
         \ADD_/FAINST[65].FA_/n2 , \ADD_/FAINST[65].FA_/n1 ,
         \ADD_/FAINST[64].FA_/n3 , \ADD_/FAINST[64].FA_/n2 ,
         \ADD_/FAINST[64].FA_/n1 , \ADD_/FAINST[63].FA_/n3 ,
         \ADD_/FAINST[63].FA_/n2 , \ADD_/FAINST[63].FA_/n1 ,
         \ADD_/FAINST[62].FA_/n3 , \ADD_/FAINST[62].FA_/n2 ,
         \ADD_/FAINST[62].FA_/n1 , \ADD_/FAINST[61].FA_/n3 ,
         \ADD_/FAINST[61].FA_/n2 , \ADD_/FAINST[61].FA_/n1 ,
         \ADD_/FAINST[60].FA_/n3 , \ADD_/FAINST[60].FA_/n2 ,
         \ADD_/FAINST[60].FA_/n1 , \ADD_/FAINST[59].FA_/n3 ,
         \ADD_/FAINST[59].FA_/n2 , \ADD_/FAINST[59].FA_/n1 ,
         \ADD_/FAINST[58].FA_/n3 , \ADD_/FAINST[58].FA_/n2 ,
         \ADD_/FAINST[58].FA_/n1 , \ADD_/FAINST[57].FA_/n3 ,
         \ADD_/FAINST[57].FA_/n2 , \ADD_/FAINST[57].FA_/n1 ,
         \ADD_/FAINST[56].FA_/n3 , \ADD_/FAINST[56].FA_/n2 ,
         \ADD_/FAINST[56].FA_/n1 , \ADD_/FAINST[55].FA_/n3 ,
         \ADD_/FAINST[55].FA_/n2 , \ADD_/FAINST[55].FA_/n1 ,
         \ADD_/FAINST[54].FA_/n3 , \ADD_/FAINST[54].FA_/n2 ,
         \ADD_/FAINST[54].FA_/n1 , \ADD_/FAINST[53].FA_/n3 ,
         \ADD_/FAINST[53].FA_/n2 , \ADD_/FAINST[53].FA_/n1 ,
         \ADD_/FAINST[52].FA_/n3 , \ADD_/FAINST[52].FA_/n2 ,
         \ADD_/FAINST[52].FA_/n1 , \ADD_/FAINST[51].FA_/n3 ,
         \ADD_/FAINST[51].FA_/n2 , \ADD_/FAINST[51].FA_/n1 ,
         \ADD_/FAINST[50].FA_/n3 , \ADD_/FAINST[50].FA_/n2 ,
         \ADD_/FAINST[50].FA_/n1 , \ADD_/FAINST[49].FA_/n3 ,
         \ADD_/FAINST[49].FA_/n2 , \ADD_/FAINST[49].FA_/n1 ,
         \ADD_/FAINST[48].FA_/n3 , \ADD_/FAINST[48].FA_/n2 ,
         \ADD_/FAINST[48].FA_/n1 , \ADD_/FAINST[47].FA_/n3 ,
         \ADD_/FAINST[47].FA_/n2 , \ADD_/FAINST[47].FA_/n1 ,
         \ADD_/FAINST[46].FA_/n3 , \ADD_/FAINST[46].FA_/n2 ,
         \ADD_/FAINST[46].FA_/n1 , \ADD_/FAINST[45].FA_/n3 ,
         \ADD_/FAINST[45].FA_/n2 , \ADD_/FAINST[45].FA_/n1 ,
         \ADD_/FAINST[44].FA_/n3 , \ADD_/FAINST[44].FA_/n2 ,
         \ADD_/FAINST[44].FA_/n1 , \ADD_/FAINST[43].FA_/n3 ,
         \ADD_/FAINST[43].FA_/n2 , \ADD_/FAINST[43].FA_/n1 ,
         \ADD_/FAINST[42].FA_/n3 , \ADD_/FAINST[42].FA_/n2 ,
         \ADD_/FAINST[42].FA_/n1 , \ADD_/FAINST[41].FA_/n3 ,
         \ADD_/FAINST[41].FA_/n2 , \ADD_/FAINST[41].FA_/n1 ,
         \ADD_/FAINST[40].FA_/n3 , \ADD_/FAINST[40].FA_/n2 ,
         \ADD_/FAINST[40].FA_/n1 , \ADD_/FAINST[39].FA_/n3 ,
         \ADD_/FAINST[39].FA_/n2 , \ADD_/FAINST[39].FA_/n1 ,
         \ADD_/FAINST[38].FA_/n3 , \ADD_/FAINST[38].FA_/n2 ,
         \ADD_/FAINST[38].FA_/n1 , \ADD_/FAINST[37].FA_/n3 ,
         \ADD_/FAINST[37].FA_/n2 , \ADD_/FAINST[37].FA_/n1 ,
         \ADD_/FAINST[36].FA_/n3 , \ADD_/FAINST[36].FA_/n2 ,
         \ADD_/FAINST[36].FA_/n1 , \ADD_/FAINST[35].FA_/n3 ,
         \ADD_/FAINST[35].FA_/n2 , \ADD_/FAINST[35].FA_/n1 ,
         \ADD_/FAINST[34].FA_/n3 , \ADD_/FAINST[34].FA_/n2 ,
         \ADD_/FAINST[34].FA_/n1 , \ADD_/FAINST[33].FA_/n3 ,
         \ADD_/FAINST[33].FA_/n2 , \ADD_/FAINST[33].FA_/n1 ,
         \ADD_/FAINST[32].FA_/n3 , \ADD_/FAINST[32].FA_/n2 ,
         \ADD_/FAINST[32].FA_/n1 , \ADD_/FAINST[31].FA_/n3 ,
         \ADD_/FAINST[31].FA_/n2 , \ADD_/FAINST[31].FA_/n1 ,
         \ADD_/FAINST[30].FA_/n3 , \ADD_/FAINST[30].FA_/n2 ,
         \ADD_/FAINST[30].FA_/n1 , \ADD_/FAINST[29].FA_/n3 ,
         \ADD_/FAINST[29].FA_/n2 , \ADD_/FAINST[29].FA_/n1 ,
         \ADD_/FAINST[28].FA_/n3 , \ADD_/FAINST[28].FA_/n2 ,
         \ADD_/FAINST[28].FA_/n1 , \ADD_/FAINST[27].FA_/n3 ,
         \ADD_/FAINST[27].FA_/n2 , \ADD_/FAINST[27].FA_/n1 ,
         \ADD_/FAINST[26].FA_/n3 , \ADD_/FAINST[26].FA_/n2 ,
         \ADD_/FAINST[26].FA_/n1 , \ADD_/FAINST[25].FA_/n3 ,
         \ADD_/FAINST[25].FA_/n2 , \ADD_/FAINST[25].FA_/n1 ,
         \ADD_/FAINST[24].FA_/n3 , \ADD_/FAINST[24].FA_/n2 ,
         \ADD_/FAINST[24].FA_/n1 , \ADD_/FAINST[23].FA_/n3 ,
         \ADD_/FAINST[23].FA_/n2 , \ADD_/FAINST[23].FA_/n1 ,
         \ADD_/FAINST[22].FA_/n3 , \ADD_/FAINST[22].FA_/n2 ,
         \ADD_/FAINST[22].FA_/n1 , \ADD_/FAINST[21].FA_/n3 ,
         \ADD_/FAINST[21].FA_/n2 , \ADD_/FAINST[21].FA_/n1 ,
         \ADD_/FAINST[20].FA_/n3 , \ADD_/FAINST[20].FA_/n2 ,
         \ADD_/FAINST[20].FA_/n1 , \ADD_/FAINST[19].FA_/n3 ,
         \ADD_/FAINST[19].FA_/n2 , \ADD_/FAINST[19].FA_/n1 ,
         \ADD_/FAINST[18].FA_/n3 , \ADD_/FAINST[18].FA_/n2 ,
         \ADD_/FAINST[18].FA_/n1 , \ADD_/FAINST[17].FA_/n3 ,
         \ADD_/FAINST[17].FA_/n2 , \ADD_/FAINST[17].FA_/n1 ,
         \ADD_/FAINST[16].FA_/n3 , \ADD_/FAINST[16].FA_/n2 ,
         \ADD_/FAINST[16].FA_/n1 , \ADD_/FAINST[15].FA_/n3 ,
         \ADD_/FAINST[15].FA_/n2 , \ADD_/FAINST[15].FA_/n1 ,
         \ADD_/FAINST[14].FA_/n3 , \ADD_/FAINST[14].FA_/n2 ,
         \ADD_/FAINST[14].FA_/n1 , \ADD_/FAINST[13].FA_/n3 ,
         \ADD_/FAINST[13].FA_/n2 , \ADD_/FAINST[13].FA_/n1 ,
         \ADD_/FAINST[12].FA_/n3 , \ADD_/FAINST[12].FA_/n2 ,
         \ADD_/FAINST[12].FA_/n1 , \ADD_/FAINST[11].FA_/n3 ,
         \ADD_/FAINST[11].FA_/n2 , \ADD_/FAINST[11].FA_/n1 ,
         \ADD_/FAINST[10].FA_/n3 , \ADD_/FAINST[10].FA_/n2 ,
         \ADD_/FAINST[10].FA_/n1 , \ADD_/FAINST[9].FA_/n3 ,
         \ADD_/FAINST[9].FA_/n2 , \ADD_/FAINST[9].FA_/n1 ,
         \ADD_/FAINST[8].FA_/n3 , \ADD_/FAINST[8].FA_/n2 ,
         \ADD_/FAINST[8].FA_/n1 , \ADD_/FAINST[7].FA_/n3 ,
         \ADD_/FAINST[7].FA_/n2 , \ADD_/FAINST[7].FA_/n1 ,
         \ADD_/FAINST[6].FA_/n3 , \ADD_/FAINST[6].FA_/n2 ,
         \ADD_/FAINST[6].FA_/n1 , \ADD_/FAINST[5].FA_/n3 ,
         \ADD_/FAINST[5].FA_/n2 , \ADD_/FAINST[5].FA_/n1 ,
         \ADD_/FAINST[4].FA_/n3 , \ADD_/FAINST[4].FA_/n2 ,
         \ADD_/FAINST[4].FA_/n1 , \ADD_/FAINST[3].FA_/n3 ,
         \ADD_/FAINST[3].FA_/n2 , \ADD_/FAINST[3].FA_/n1 ,
         \ADD_/FAINST[2].FA_/n3 , \ADD_/FAINST[2].FA_/n2 ,
         \ADD_/FAINST[2].FA_/n1 , \ADD_/FAINST[1].FA_/n3 ,
         \ADD_/FAINST[1].FA_/n2 , \ADD_/FAINST[1].FA_/n1 ;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR \ADD_/FAINST[0].FA_/U5  ( .A(\ADD_/FAINST[0].FA_/n3 ), .B(carry_on), .Z(
        \ADD_/c[1] ) );
  XOR \ADD_/FAINST[0].FA_/U4  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(b[0]), .Z(c[0]) );
  AND \ADD_/FAINST[0].FA_/U3  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(
        \ADD_/FAINST[0].FA_/n2 ), .Z(\ADD_/FAINST[0].FA_/n3 ) );
  XOR \ADD_/FAINST[0].FA_/U2  ( .A(b[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n2 ) );
  XOR \ADD_/FAINST[0].FA_/U1  ( .A(a[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n1 ) );
  XOR \ADD_/FAINST[255].FA_/U5  ( .A(\ADD_/FAINST[255].FA_/n3 ), .B(
        \ADD_/c[255] ), .Z(carry_on_d) );
  XOR \ADD_/FAINST[255].FA_/U4  ( .A(\ADD_/FAINST[255].FA_/n1 ), .B(b[255]), 
        .Z(c[255]) );
  AND \ADD_/FAINST[255].FA_/U3  ( .A(\ADD_/FAINST[255].FA_/n1 ), .B(
        \ADD_/FAINST[255].FA_/n2 ), .Z(\ADD_/FAINST[255].FA_/n3 ) );
  XOR \ADD_/FAINST[255].FA_/U2  ( .A(b[255]), .B(\ADD_/c[255] ), .Z(
        \ADD_/FAINST[255].FA_/n2 ) );
  XOR \ADD_/FAINST[255].FA_/U1  ( .A(a[255]), .B(\ADD_/c[255] ), .Z(
        \ADD_/FAINST[255].FA_/n1 ) );
  XOR \ADD_/FAINST[254].FA_/U5  ( .A(\ADD_/FAINST[254].FA_/n3 ), .B(
        \ADD_/c[254] ), .Z(\ADD_/c[255] ) );
  XOR \ADD_/FAINST[254].FA_/U4  ( .A(\ADD_/FAINST[254].FA_/n1 ), .B(b[254]), 
        .Z(c[254]) );
  AND \ADD_/FAINST[254].FA_/U3  ( .A(\ADD_/FAINST[254].FA_/n1 ), .B(
        \ADD_/FAINST[254].FA_/n2 ), .Z(\ADD_/FAINST[254].FA_/n3 ) );
  XOR \ADD_/FAINST[254].FA_/U2  ( .A(b[254]), .B(\ADD_/c[254] ), .Z(
        \ADD_/FAINST[254].FA_/n2 ) );
  XOR \ADD_/FAINST[254].FA_/U1  ( .A(a[254]), .B(\ADD_/c[254] ), .Z(
        \ADD_/FAINST[254].FA_/n1 ) );
  XOR \ADD_/FAINST[253].FA_/U5  ( .A(\ADD_/FAINST[253].FA_/n3 ), .B(
        \ADD_/c[253] ), .Z(\ADD_/c[254] ) );
  XOR \ADD_/FAINST[253].FA_/U4  ( .A(\ADD_/FAINST[253].FA_/n1 ), .B(b[253]), 
        .Z(c[253]) );
  AND \ADD_/FAINST[253].FA_/U3  ( .A(\ADD_/FAINST[253].FA_/n1 ), .B(
        \ADD_/FAINST[253].FA_/n2 ), .Z(\ADD_/FAINST[253].FA_/n3 ) );
  XOR \ADD_/FAINST[253].FA_/U2  ( .A(b[253]), .B(\ADD_/c[253] ), .Z(
        \ADD_/FAINST[253].FA_/n2 ) );
  XOR \ADD_/FAINST[253].FA_/U1  ( .A(a[253]), .B(\ADD_/c[253] ), .Z(
        \ADD_/FAINST[253].FA_/n1 ) );
  XOR \ADD_/FAINST[252].FA_/U5  ( .A(\ADD_/FAINST[252].FA_/n3 ), .B(
        \ADD_/c[252] ), .Z(\ADD_/c[253] ) );
  XOR \ADD_/FAINST[252].FA_/U4  ( .A(\ADD_/FAINST[252].FA_/n1 ), .B(b[252]), 
        .Z(c[252]) );
  AND \ADD_/FAINST[252].FA_/U3  ( .A(\ADD_/FAINST[252].FA_/n1 ), .B(
        \ADD_/FAINST[252].FA_/n2 ), .Z(\ADD_/FAINST[252].FA_/n3 ) );
  XOR \ADD_/FAINST[252].FA_/U2  ( .A(b[252]), .B(\ADD_/c[252] ), .Z(
        \ADD_/FAINST[252].FA_/n2 ) );
  XOR \ADD_/FAINST[252].FA_/U1  ( .A(a[252]), .B(\ADD_/c[252] ), .Z(
        \ADD_/FAINST[252].FA_/n1 ) );
  XOR \ADD_/FAINST[251].FA_/U5  ( .A(\ADD_/FAINST[251].FA_/n3 ), .B(
        \ADD_/c[251] ), .Z(\ADD_/c[252] ) );
  XOR \ADD_/FAINST[251].FA_/U4  ( .A(\ADD_/FAINST[251].FA_/n1 ), .B(b[251]), 
        .Z(c[251]) );
  AND \ADD_/FAINST[251].FA_/U3  ( .A(\ADD_/FAINST[251].FA_/n1 ), .B(
        \ADD_/FAINST[251].FA_/n2 ), .Z(\ADD_/FAINST[251].FA_/n3 ) );
  XOR \ADD_/FAINST[251].FA_/U2  ( .A(b[251]), .B(\ADD_/c[251] ), .Z(
        \ADD_/FAINST[251].FA_/n2 ) );
  XOR \ADD_/FAINST[251].FA_/U1  ( .A(a[251]), .B(\ADD_/c[251] ), .Z(
        \ADD_/FAINST[251].FA_/n1 ) );
  XOR \ADD_/FAINST[250].FA_/U5  ( .A(\ADD_/FAINST[250].FA_/n3 ), .B(
        \ADD_/c[250] ), .Z(\ADD_/c[251] ) );
  XOR \ADD_/FAINST[250].FA_/U4  ( .A(\ADD_/FAINST[250].FA_/n1 ), .B(b[250]), 
        .Z(c[250]) );
  AND \ADD_/FAINST[250].FA_/U3  ( .A(\ADD_/FAINST[250].FA_/n1 ), .B(
        \ADD_/FAINST[250].FA_/n2 ), .Z(\ADD_/FAINST[250].FA_/n3 ) );
  XOR \ADD_/FAINST[250].FA_/U2  ( .A(b[250]), .B(\ADD_/c[250] ), .Z(
        \ADD_/FAINST[250].FA_/n2 ) );
  XOR \ADD_/FAINST[250].FA_/U1  ( .A(a[250]), .B(\ADD_/c[250] ), .Z(
        \ADD_/FAINST[250].FA_/n1 ) );
  XOR \ADD_/FAINST[249].FA_/U5  ( .A(\ADD_/FAINST[249].FA_/n3 ), .B(
        \ADD_/c[249] ), .Z(\ADD_/c[250] ) );
  XOR \ADD_/FAINST[249].FA_/U4  ( .A(\ADD_/FAINST[249].FA_/n1 ), .B(b[249]), 
        .Z(c[249]) );
  AND \ADD_/FAINST[249].FA_/U3  ( .A(\ADD_/FAINST[249].FA_/n1 ), .B(
        \ADD_/FAINST[249].FA_/n2 ), .Z(\ADD_/FAINST[249].FA_/n3 ) );
  XOR \ADD_/FAINST[249].FA_/U2  ( .A(b[249]), .B(\ADD_/c[249] ), .Z(
        \ADD_/FAINST[249].FA_/n2 ) );
  XOR \ADD_/FAINST[249].FA_/U1  ( .A(a[249]), .B(\ADD_/c[249] ), .Z(
        \ADD_/FAINST[249].FA_/n1 ) );
  XOR \ADD_/FAINST[248].FA_/U5  ( .A(\ADD_/FAINST[248].FA_/n3 ), .B(
        \ADD_/c[248] ), .Z(\ADD_/c[249] ) );
  XOR \ADD_/FAINST[248].FA_/U4  ( .A(\ADD_/FAINST[248].FA_/n1 ), .B(b[248]), 
        .Z(c[248]) );
  AND \ADD_/FAINST[248].FA_/U3  ( .A(\ADD_/FAINST[248].FA_/n1 ), .B(
        \ADD_/FAINST[248].FA_/n2 ), .Z(\ADD_/FAINST[248].FA_/n3 ) );
  XOR \ADD_/FAINST[248].FA_/U2  ( .A(b[248]), .B(\ADD_/c[248] ), .Z(
        \ADD_/FAINST[248].FA_/n2 ) );
  XOR \ADD_/FAINST[248].FA_/U1  ( .A(a[248]), .B(\ADD_/c[248] ), .Z(
        \ADD_/FAINST[248].FA_/n1 ) );
  XOR \ADD_/FAINST[247].FA_/U5  ( .A(\ADD_/FAINST[247].FA_/n3 ), .B(
        \ADD_/c[247] ), .Z(\ADD_/c[248] ) );
  XOR \ADD_/FAINST[247].FA_/U4  ( .A(\ADD_/FAINST[247].FA_/n1 ), .B(b[247]), 
        .Z(c[247]) );
  AND \ADD_/FAINST[247].FA_/U3  ( .A(\ADD_/FAINST[247].FA_/n1 ), .B(
        \ADD_/FAINST[247].FA_/n2 ), .Z(\ADD_/FAINST[247].FA_/n3 ) );
  XOR \ADD_/FAINST[247].FA_/U2  ( .A(b[247]), .B(\ADD_/c[247] ), .Z(
        \ADD_/FAINST[247].FA_/n2 ) );
  XOR \ADD_/FAINST[247].FA_/U1  ( .A(a[247]), .B(\ADD_/c[247] ), .Z(
        \ADD_/FAINST[247].FA_/n1 ) );
  XOR \ADD_/FAINST[246].FA_/U5  ( .A(\ADD_/FAINST[246].FA_/n3 ), .B(
        \ADD_/c[246] ), .Z(\ADD_/c[247] ) );
  XOR \ADD_/FAINST[246].FA_/U4  ( .A(\ADD_/FAINST[246].FA_/n1 ), .B(b[246]), 
        .Z(c[246]) );
  AND \ADD_/FAINST[246].FA_/U3  ( .A(\ADD_/FAINST[246].FA_/n1 ), .B(
        \ADD_/FAINST[246].FA_/n2 ), .Z(\ADD_/FAINST[246].FA_/n3 ) );
  XOR \ADD_/FAINST[246].FA_/U2  ( .A(b[246]), .B(\ADD_/c[246] ), .Z(
        \ADD_/FAINST[246].FA_/n2 ) );
  XOR \ADD_/FAINST[246].FA_/U1  ( .A(a[246]), .B(\ADD_/c[246] ), .Z(
        \ADD_/FAINST[246].FA_/n1 ) );
  XOR \ADD_/FAINST[245].FA_/U5  ( .A(\ADD_/FAINST[245].FA_/n3 ), .B(
        \ADD_/c[245] ), .Z(\ADD_/c[246] ) );
  XOR \ADD_/FAINST[245].FA_/U4  ( .A(\ADD_/FAINST[245].FA_/n1 ), .B(b[245]), 
        .Z(c[245]) );
  AND \ADD_/FAINST[245].FA_/U3  ( .A(\ADD_/FAINST[245].FA_/n1 ), .B(
        \ADD_/FAINST[245].FA_/n2 ), .Z(\ADD_/FAINST[245].FA_/n3 ) );
  XOR \ADD_/FAINST[245].FA_/U2  ( .A(b[245]), .B(\ADD_/c[245] ), .Z(
        \ADD_/FAINST[245].FA_/n2 ) );
  XOR \ADD_/FAINST[245].FA_/U1  ( .A(a[245]), .B(\ADD_/c[245] ), .Z(
        \ADD_/FAINST[245].FA_/n1 ) );
  XOR \ADD_/FAINST[244].FA_/U5  ( .A(\ADD_/FAINST[244].FA_/n3 ), .B(
        \ADD_/c[244] ), .Z(\ADD_/c[245] ) );
  XOR \ADD_/FAINST[244].FA_/U4  ( .A(\ADD_/FAINST[244].FA_/n1 ), .B(b[244]), 
        .Z(c[244]) );
  AND \ADD_/FAINST[244].FA_/U3  ( .A(\ADD_/FAINST[244].FA_/n1 ), .B(
        \ADD_/FAINST[244].FA_/n2 ), .Z(\ADD_/FAINST[244].FA_/n3 ) );
  XOR \ADD_/FAINST[244].FA_/U2  ( .A(b[244]), .B(\ADD_/c[244] ), .Z(
        \ADD_/FAINST[244].FA_/n2 ) );
  XOR \ADD_/FAINST[244].FA_/U1  ( .A(a[244]), .B(\ADD_/c[244] ), .Z(
        \ADD_/FAINST[244].FA_/n1 ) );
  XOR \ADD_/FAINST[243].FA_/U5  ( .A(\ADD_/FAINST[243].FA_/n3 ), .B(
        \ADD_/c[243] ), .Z(\ADD_/c[244] ) );
  XOR \ADD_/FAINST[243].FA_/U4  ( .A(\ADD_/FAINST[243].FA_/n1 ), .B(b[243]), 
        .Z(c[243]) );
  AND \ADD_/FAINST[243].FA_/U3  ( .A(\ADD_/FAINST[243].FA_/n1 ), .B(
        \ADD_/FAINST[243].FA_/n2 ), .Z(\ADD_/FAINST[243].FA_/n3 ) );
  XOR \ADD_/FAINST[243].FA_/U2  ( .A(b[243]), .B(\ADD_/c[243] ), .Z(
        \ADD_/FAINST[243].FA_/n2 ) );
  XOR \ADD_/FAINST[243].FA_/U1  ( .A(a[243]), .B(\ADD_/c[243] ), .Z(
        \ADD_/FAINST[243].FA_/n1 ) );
  XOR \ADD_/FAINST[242].FA_/U5  ( .A(\ADD_/FAINST[242].FA_/n3 ), .B(
        \ADD_/c[242] ), .Z(\ADD_/c[243] ) );
  XOR \ADD_/FAINST[242].FA_/U4  ( .A(\ADD_/FAINST[242].FA_/n1 ), .B(b[242]), 
        .Z(c[242]) );
  AND \ADD_/FAINST[242].FA_/U3  ( .A(\ADD_/FAINST[242].FA_/n1 ), .B(
        \ADD_/FAINST[242].FA_/n2 ), .Z(\ADD_/FAINST[242].FA_/n3 ) );
  XOR \ADD_/FAINST[242].FA_/U2  ( .A(b[242]), .B(\ADD_/c[242] ), .Z(
        \ADD_/FAINST[242].FA_/n2 ) );
  XOR \ADD_/FAINST[242].FA_/U1  ( .A(a[242]), .B(\ADD_/c[242] ), .Z(
        \ADD_/FAINST[242].FA_/n1 ) );
  XOR \ADD_/FAINST[241].FA_/U5  ( .A(\ADD_/FAINST[241].FA_/n3 ), .B(
        \ADD_/c[241] ), .Z(\ADD_/c[242] ) );
  XOR \ADD_/FAINST[241].FA_/U4  ( .A(\ADD_/FAINST[241].FA_/n1 ), .B(b[241]), 
        .Z(c[241]) );
  AND \ADD_/FAINST[241].FA_/U3  ( .A(\ADD_/FAINST[241].FA_/n1 ), .B(
        \ADD_/FAINST[241].FA_/n2 ), .Z(\ADD_/FAINST[241].FA_/n3 ) );
  XOR \ADD_/FAINST[241].FA_/U2  ( .A(b[241]), .B(\ADD_/c[241] ), .Z(
        \ADD_/FAINST[241].FA_/n2 ) );
  XOR \ADD_/FAINST[241].FA_/U1  ( .A(a[241]), .B(\ADD_/c[241] ), .Z(
        \ADD_/FAINST[241].FA_/n1 ) );
  XOR \ADD_/FAINST[240].FA_/U5  ( .A(\ADD_/FAINST[240].FA_/n3 ), .B(
        \ADD_/c[240] ), .Z(\ADD_/c[241] ) );
  XOR \ADD_/FAINST[240].FA_/U4  ( .A(\ADD_/FAINST[240].FA_/n1 ), .B(b[240]), 
        .Z(c[240]) );
  AND \ADD_/FAINST[240].FA_/U3  ( .A(\ADD_/FAINST[240].FA_/n1 ), .B(
        \ADD_/FAINST[240].FA_/n2 ), .Z(\ADD_/FAINST[240].FA_/n3 ) );
  XOR \ADD_/FAINST[240].FA_/U2  ( .A(b[240]), .B(\ADD_/c[240] ), .Z(
        \ADD_/FAINST[240].FA_/n2 ) );
  XOR \ADD_/FAINST[240].FA_/U1  ( .A(a[240]), .B(\ADD_/c[240] ), .Z(
        \ADD_/FAINST[240].FA_/n1 ) );
  XOR \ADD_/FAINST[239].FA_/U5  ( .A(\ADD_/FAINST[239].FA_/n3 ), .B(
        \ADD_/c[239] ), .Z(\ADD_/c[240] ) );
  XOR \ADD_/FAINST[239].FA_/U4  ( .A(\ADD_/FAINST[239].FA_/n1 ), .B(b[239]), 
        .Z(c[239]) );
  AND \ADD_/FAINST[239].FA_/U3  ( .A(\ADD_/FAINST[239].FA_/n1 ), .B(
        \ADD_/FAINST[239].FA_/n2 ), .Z(\ADD_/FAINST[239].FA_/n3 ) );
  XOR \ADD_/FAINST[239].FA_/U2  ( .A(b[239]), .B(\ADD_/c[239] ), .Z(
        \ADD_/FAINST[239].FA_/n2 ) );
  XOR \ADD_/FAINST[239].FA_/U1  ( .A(a[239]), .B(\ADD_/c[239] ), .Z(
        \ADD_/FAINST[239].FA_/n1 ) );
  XOR \ADD_/FAINST[238].FA_/U5  ( .A(\ADD_/FAINST[238].FA_/n3 ), .B(
        \ADD_/c[238] ), .Z(\ADD_/c[239] ) );
  XOR \ADD_/FAINST[238].FA_/U4  ( .A(\ADD_/FAINST[238].FA_/n1 ), .B(b[238]), 
        .Z(c[238]) );
  AND \ADD_/FAINST[238].FA_/U3  ( .A(\ADD_/FAINST[238].FA_/n1 ), .B(
        \ADD_/FAINST[238].FA_/n2 ), .Z(\ADD_/FAINST[238].FA_/n3 ) );
  XOR \ADD_/FAINST[238].FA_/U2  ( .A(b[238]), .B(\ADD_/c[238] ), .Z(
        \ADD_/FAINST[238].FA_/n2 ) );
  XOR \ADD_/FAINST[238].FA_/U1  ( .A(a[238]), .B(\ADD_/c[238] ), .Z(
        \ADD_/FAINST[238].FA_/n1 ) );
  XOR \ADD_/FAINST[237].FA_/U5  ( .A(\ADD_/FAINST[237].FA_/n3 ), .B(
        \ADD_/c[237] ), .Z(\ADD_/c[238] ) );
  XOR \ADD_/FAINST[237].FA_/U4  ( .A(\ADD_/FAINST[237].FA_/n1 ), .B(b[237]), 
        .Z(c[237]) );
  AND \ADD_/FAINST[237].FA_/U3  ( .A(\ADD_/FAINST[237].FA_/n1 ), .B(
        \ADD_/FAINST[237].FA_/n2 ), .Z(\ADD_/FAINST[237].FA_/n3 ) );
  XOR \ADD_/FAINST[237].FA_/U2  ( .A(b[237]), .B(\ADD_/c[237] ), .Z(
        \ADD_/FAINST[237].FA_/n2 ) );
  XOR \ADD_/FAINST[237].FA_/U1  ( .A(a[237]), .B(\ADD_/c[237] ), .Z(
        \ADD_/FAINST[237].FA_/n1 ) );
  XOR \ADD_/FAINST[236].FA_/U5  ( .A(\ADD_/FAINST[236].FA_/n3 ), .B(
        \ADD_/c[236] ), .Z(\ADD_/c[237] ) );
  XOR \ADD_/FAINST[236].FA_/U4  ( .A(\ADD_/FAINST[236].FA_/n1 ), .B(b[236]), 
        .Z(c[236]) );
  AND \ADD_/FAINST[236].FA_/U3  ( .A(\ADD_/FAINST[236].FA_/n1 ), .B(
        \ADD_/FAINST[236].FA_/n2 ), .Z(\ADD_/FAINST[236].FA_/n3 ) );
  XOR \ADD_/FAINST[236].FA_/U2  ( .A(b[236]), .B(\ADD_/c[236] ), .Z(
        \ADD_/FAINST[236].FA_/n2 ) );
  XOR \ADD_/FAINST[236].FA_/U1  ( .A(a[236]), .B(\ADD_/c[236] ), .Z(
        \ADD_/FAINST[236].FA_/n1 ) );
  XOR \ADD_/FAINST[235].FA_/U5  ( .A(\ADD_/FAINST[235].FA_/n3 ), .B(
        \ADD_/c[235] ), .Z(\ADD_/c[236] ) );
  XOR \ADD_/FAINST[235].FA_/U4  ( .A(\ADD_/FAINST[235].FA_/n1 ), .B(b[235]), 
        .Z(c[235]) );
  AND \ADD_/FAINST[235].FA_/U3  ( .A(\ADD_/FAINST[235].FA_/n1 ), .B(
        \ADD_/FAINST[235].FA_/n2 ), .Z(\ADD_/FAINST[235].FA_/n3 ) );
  XOR \ADD_/FAINST[235].FA_/U2  ( .A(b[235]), .B(\ADD_/c[235] ), .Z(
        \ADD_/FAINST[235].FA_/n2 ) );
  XOR \ADD_/FAINST[235].FA_/U1  ( .A(a[235]), .B(\ADD_/c[235] ), .Z(
        \ADD_/FAINST[235].FA_/n1 ) );
  XOR \ADD_/FAINST[234].FA_/U5  ( .A(\ADD_/FAINST[234].FA_/n3 ), .B(
        \ADD_/c[234] ), .Z(\ADD_/c[235] ) );
  XOR \ADD_/FAINST[234].FA_/U4  ( .A(\ADD_/FAINST[234].FA_/n1 ), .B(b[234]), 
        .Z(c[234]) );
  AND \ADD_/FAINST[234].FA_/U3  ( .A(\ADD_/FAINST[234].FA_/n1 ), .B(
        \ADD_/FAINST[234].FA_/n2 ), .Z(\ADD_/FAINST[234].FA_/n3 ) );
  XOR \ADD_/FAINST[234].FA_/U2  ( .A(b[234]), .B(\ADD_/c[234] ), .Z(
        \ADD_/FAINST[234].FA_/n2 ) );
  XOR \ADD_/FAINST[234].FA_/U1  ( .A(a[234]), .B(\ADD_/c[234] ), .Z(
        \ADD_/FAINST[234].FA_/n1 ) );
  XOR \ADD_/FAINST[233].FA_/U5  ( .A(\ADD_/FAINST[233].FA_/n3 ), .B(
        \ADD_/c[233] ), .Z(\ADD_/c[234] ) );
  XOR \ADD_/FAINST[233].FA_/U4  ( .A(\ADD_/FAINST[233].FA_/n1 ), .B(b[233]), 
        .Z(c[233]) );
  AND \ADD_/FAINST[233].FA_/U3  ( .A(\ADD_/FAINST[233].FA_/n1 ), .B(
        \ADD_/FAINST[233].FA_/n2 ), .Z(\ADD_/FAINST[233].FA_/n3 ) );
  XOR \ADD_/FAINST[233].FA_/U2  ( .A(b[233]), .B(\ADD_/c[233] ), .Z(
        \ADD_/FAINST[233].FA_/n2 ) );
  XOR \ADD_/FAINST[233].FA_/U1  ( .A(a[233]), .B(\ADD_/c[233] ), .Z(
        \ADD_/FAINST[233].FA_/n1 ) );
  XOR \ADD_/FAINST[232].FA_/U5  ( .A(\ADD_/FAINST[232].FA_/n3 ), .B(
        \ADD_/c[232] ), .Z(\ADD_/c[233] ) );
  XOR \ADD_/FAINST[232].FA_/U4  ( .A(\ADD_/FAINST[232].FA_/n1 ), .B(b[232]), 
        .Z(c[232]) );
  AND \ADD_/FAINST[232].FA_/U3  ( .A(\ADD_/FAINST[232].FA_/n1 ), .B(
        \ADD_/FAINST[232].FA_/n2 ), .Z(\ADD_/FAINST[232].FA_/n3 ) );
  XOR \ADD_/FAINST[232].FA_/U2  ( .A(b[232]), .B(\ADD_/c[232] ), .Z(
        \ADD_/FAINST[232].FA_/n2 ) );
  XOR \ADD_/FAINST[232].FA_/U1  ( .A(a[232]), .B(\ADD_/c[232] ), .Z(
        \ADD_/FAINST[232].FA_/n1 ) );
  XOR \ADD_/FAINST[231].FA_/U5  ( .A(\ADD_/FAINST[231].FA_/n3 ), .B(
        \ADD_/c[231] ), .Z(\ADD_/c[232] ) );
  XOR \ADD_/FAINST[231].FA_/U4  ( .A(\ADD_/FAINST[231].FA_/n1 ), .B(b[231]), 
        .Z(c[231]) );
  AND \ADD_/FAINST[231].FA_/U3  ( .A(\ADD_/FAINST[231].FA_/n1 ), .B(
        \ADD_/FAINST[231].FA_/n2 ), .Z(\ADD_/FAINST[231].FA_/n3 ) );
  XOR \ADD_/FAINST[231].FA_/U2  ( .A(b[231]), .B(\ADD_/c[231] ), .Z(
        \ADD_/FAINST[231].FA_/n2 ) );
  XOR \ADD_/FAINST[231].FA_/U1  ( .A(a[231]), .B(\ADD_/c[231] ), .Z(
        \ADD_/FAINST[231].FA_/n1 ) );
  XOR \ADD_/FAINST[230].FA_/U5  ( .A(\ADD_/FAINST[230].FA_/n3 ), .B(
        \ADD_/c[230] ), .Z(\ADD_/c[231] ) );
  XOR \ADD_/FAINST[230].FA_/U4  ( .A(\ADD_/FAINST[230].FA_/n1 ), .B(b[230]), 
        .Z(c[230]) );
  AND \ADD_/FAINST[230].FA_/U3  ( .A(\ADD_/FAINST[230].FA_/n1 ), .B(
        \ADD_/FAINST[230].FA_/n2 ), .Z(\ADD_/FAINST[230].FA_/n3 ) );
  XOR \ADD_/FAINST[230].FA_/U2  ( .A(b[230]), .B(\ADD_/c[230] ), .Z(
        \ADD_/FAINST[230].FA_/n2 ) );
  XOR \ADD_/FAINST[230].FA_/U1  ( .A(a[230]), .B(\ADD_/c[230] ), .Z(
        \ADD_/FAINST[230].FA_/n1 ) );
  XOR \ADD_/FAINST[229].FA_/U5  ( .A(\ADD_/FAINST[229].FA_/n3 ), .B(
        \ADD_/c[229] ), .Z(\ADD_/c[230] ) );
  XOR \ADD_/FAINST[229].FA_/U4  ( .A(\ADD_/FAINST[229].FA_/n1 ), .B(b[229]), 
        .Z(c[229]) );
  AND \ADD_/FAINST[229].FA_/U3  ( .A(\ADD_/FAINST[229].FA_/n1 ), .B(
        \ADD_/FAINST[229].FA_/n2 ), .Z(\ADD_/FAINST[229].FA_/n3 ) );
  XOR \ADD_/FAINST[229].FA_/U2  ( .A(b[229]), .B(\ADD_/c[229] ), .Z(
        \ADD_/FAINST[229].FA_/n2 ) );
  XOR \ADD_/FAINST[229].FA_/U1  ( .A(a[229]), .B(\ADD_/c[229] ), .Z(
        \ADD_/FAINST[229].FA_/n1 ) );
  XOR \ADD_/FAINST[228].FA_/U5  ( .A(\ADD_/FAINST[228].FA_/n3 ), .B(
        \ADD_/c[228] ), .Z(\ADD_/c[229] ) );
  XOR \ADD_/FAINST[228].FA_/U4  ( .A(\ADD_/FAINST[228].FA_/n1 ), .B(b[228]), 
        .Z(c[228]) );
  AND \ADD_/FAINST[228].FA_/U3  ( .A(\ADD_/FAINST[228].FA_/n1 ), .B(
        \ADD_/FAINST[228].FA_/n2 ), .Z(\ADD_/FAINST[228].FA_/n3 ) );
  XOR \ADD_/FAINST[228].FA_/U2  ( .A(b[228]), .B(\ADD_/c[228] ), .Z(
        \ADD_/FAINST[228].FA_/n2 ) );
  XOR \ADD_/FAINST[228].FA_/U1  ( .A(a[228]), .B(\ADD_/c[228] ), .Z(
        \ADD_/FAINST[228].FA_/n1 ) );
  XOR \ADD_/FAINST[227].FA_/U5  ( .A(\ADD_/FAINST[227].FA_/n3 ), .B(
        \ADD_/c[227] ), .Z(\ADD_/c[228] ) );
  XOR \ADD_/FAINST[227].FA_/U4  ( .A(\ADD_/FAINST[227].FA_/n1 ), .B(b[227]), 
        .Z(c[227]) );
  AND \ADD_/FAINST[227].FA_/U3  ( .A(\ADD_/FAINST[227].FA_/n1 ), .B(
        \ADD_/FAINST[227].FA_/n2 ), .Z(\ADD_/FAINST[227].FA_/n3 ) );
  XOR \ADD_/FAINST[227].FA_/U2  ( .A(b[227]), .B(\ADD_/c[227] ), .Z(
        \ADD_/FAINST[227].FA_/n2 ) );
  XOR \ADD_/FAINST[227].FA_/U1  ( .A(a[227]), .B(\ADD_/c[227] ), .Z(
        \ADD_/FAINST[227].FA_/n1 ) );
  XOR \ADD_/FAINST[226].FA_/U5  ( .A(\ADD_/FAINST[226].FA_/n3 ), .B(
        \ADD_/c[226] ), .Z(\ADD_/c[227] ) );
  XOR \ADD_/FAINST[226].FA_/U4  ( .A(\ADD_/FAINST[226].FA_/n1 ), .B(b[226]), 
        .Z(c[226]) );
  AND \ADD_/FAINST[226].FA_/U3  ( .A(\ADD_/FAINST[226].FA_/n1 ), .B(
        \ADD_/FAINST[226].FA_/n2 ), .Z(\ADD_/FAINST[226].FA_/n3 ) );
  XOR \ADD_/FAINST[226].FA_/U2  ( .A(b[226]), .B(\ADD_/c[226] ), .Z(
        \ADD_/FAINST[226].FA_/n2 ) );
  XOR \ADD_/FAINST[226].FA_/U1  ( .A(a[226]), .B(\ADD_/c[226] ), .Z(
        \ADD_/FAINST[226].FA_/n1 ) );
  XOR \ADD_/FAINST[225].FA_/U5  ( .A(\ADD_/FAINST[225].FA_/n3 ), .B(
        \ADD_/c[225] ), .Z(\ADD_/c[226] ) );
  XOR \ADD_/FAINST[225].FA_/U4  ( .A(\ADD_/FAINST[225].FA_/n1 ), .B(b[225]), 
        .Z(c[225]) );
  AND \ADD_/FAINST[225].FA_/U3  ( .A(\ADD_/FAINST[225].FA_/n1 ), .B(
        \ADD_/FAINST[225].FA_/n2 ), .Z(\ADD_/FAINST[225].FA_/n3 ) );
  XOR \ADD_/FAINST[225].FA_/U2  ( .A(b[225]), .B(\ADD_/c[225] ), .Z(
        \ADD_/FAINST[225].FA_/n2 ) );
  XOR \ADD_/FAINST[225].FA_/U1  ( .A(a[225]), .B(\ADD_/c[225] ), .Z(
        \ADD_/FAINST[225].FA_/n1 ) );
  XOR \ADD_/FAINST[224].FA_/U5  ( .A(\ADD_/FAINST[224].FA_/n3 ), .B(
        \ADD_/c[224] ), .Z(\ADD_/c[225] ) );
  XOR \ADD_/FAINST[224].FA_/U4  ( .A(\ADD_/FAINST[224].FA_/n1 ), .B(b[224]), 
        .Z(c[224]) );
  AND \ADD_/FAINST[224].FA_/U3  ( .A(\ADD_/FAINST[224].FA_/n1 ), .B(
        \ADD_/FAINST[224].FA_/n2 ), .Z(\ADD_/FAINST[224].FA_/n3 ) );
  XOR \ADD_/FAINST[224].FA_/U2  ( .A(b[224]), .B(\ADD_/c[224] ), .Z(
        \ADD_/FAINST[224].FA_/n2 ) );
  XOR \ADD_/FAINST[224].FA_/U1  ( .A(a[224]), .B(\ADD_/c[224] ), .Z(
        \ADD_/FAINST[224].FA_/n1 ) );
  XOR \ADD_/FAINST[223].FA_/U5  ( .A(\ADD_/FAINST[223].FA_/n3 ), .B(
        \ADD_/c[223] ), .Z(\ADD_/c[224] ) );
  XOR \ADD_/FAINST[223].FA_/U4  ( .A(\ADD_/FAINST[223].FA_/n1 ), .B(b[223]), 
        .Z(c[223]) );
  AND \ADD_/FAINST[223].FA_/U3  ( .A(\ADD_/FAINST[223].FA_/n1 ), .B(
        \ADD_/FAINST[223].FA_/n2 ), .Z(\ADD_/FAINST[223].FA_/n3 ) );
  XOR \ADD_/FAINST[223].FA_/U2  ( .A(b[223]), .B(\ADD_/c[223] ), .Z(
        \ADD_/FAINST[223].FA_/n2 ) );
  XOR \ADD_/FAINST[223].FA_/U1  ( .A(a[223]), .B(\ADD_/c[223] ), .Z(
        \ADD_/FAINST[223].FA_/n1 ) );
  XOR \ADD_/FAINST[222].FA_/U5  ( .A(\ADD_/FAINST[222].FA_/n3 ), .B(
        \ADD_/c[222] ), .Z(\ADD_/c[223] ) );
  XOR \ADD_/FAINST[222].FA_/U4  ( .A(\ADD_/FAINST[222].FA_/n1 ), .B(b[222]), 
        .Z(c[222]) );
  AND \ADD_/FAINST[222].FA_/U3  ( .A(\ADD_/FAINST[222].FA_/n1 ), .B(
        \ADD_/FAINST[222].FA_/n2 ), .Z(\ADD_/FAINST[222].FA_/n3 ) );
  XOR \ADD_/FAINST[222].FA_/U2  ( .A(b[222]), .B(\ADD_/c[222] ), .Z(
        \ADD_/FAINST[222].FA_/n2 ) );
  XOR \ADD_/FAINST[222].FA_/U1  ( .A(a[222]), .B(\ADD_/c[222] ), .Z(
        \ADD_/FAINST[222].FA_/n1 ) );
  XOR \ADD_/FAINST[221].FA_/U5  ( .A(\ADD_/FAINST[221].FA_/n3 ), .B(
        \ADD_/c[221] ), .Z(\ADD_/c[222] ) );
  XOR \ADD_/FAINST[221].FA_/U4  ( .A(\ADD_/FAINST[221].FA_/n1 ), .B(b[221]), 
        .Z(c[221]) );
  AND \ADD_/FAINST[221].FA_/U3  ( .A(\ADD_/FAINST[221].FA_/n1 ), .B(
        \ADD_/FAINST[221].FA_/n2 ), .Z(\ADD_/FAINST[221].FA_/n3 ) );
  XOR \ADD_/FAINST[221].FA_/U2  ( .A(b[221]), .B(\ADD_/c[221] ), .Z(
        \ADD_/FAINST[221].FA_/n2 ) );
  XOR \ADD_/FAINST[221].FA_/U1  ( .A(a[221]), .B(\ADD_/c[221] ), .Z(
        \ADD_/FAINST[221].FA_/n1 ) );
  XOR \ADD_/FAINST[220].FA_/U5  ( .A(\ADD_/FAINST[220].FA_/n3 ), .B(
        \ADD_/c[220] ), .Z(\ADD_/c[221] ) );
  XOR \ADD_/FAINST[220].FA_/U4  ( .A(\ADD_/FAINST[220].FA_/n1 ), .B(b[220]), 
        .Z(c[220]) );
  AND \ADD_/FAINST[220].FA_/U3  ( .A(\ADD_/FAINST[220].FA_/n1 ), .B(
        \ADD_/FAINST[220].FA_/n2 ), .Z(\ADD_/FAINST[220].FA_/n3 ) );
  XOR \ADD_/FAINST[220].FA_/U2  ( .A(b[220]), .B(\ADD_/c[220] ), .Z(
        \ADD_/FAINST[220].FA_/n2 ) );
  XOR \ADD_/FAINST[220].FA_/U1  ( .A(a[220]), .B(\ADD_/c[220] ), .Z(
        \ADD_/FAINST[220].FA_/n1 ) );
  XOR \ADD_/FAINST[219].FA_/U5  ( .A(\ADD_/FAINST[219].FA_/n3 ), .B(
        \ADD_/c[219] ), .Z(\ADD_/c[220] ) );
  XOR \ADD_/FAINST[219].FA_/U4  ( .A(\ADD_/FAINST[219].FA_/n1 ), .B(b[219]), 
        .Z(c[219]) );
  AND \ADD_/FAINST[219].FA_/U3  ( .A(\ADD_/FAINST[219].FA_/n1 ), .B(
        \ADD_/FAINST[219].FA_/n2 ), .Z(\ADD_/FAINST[219].FA_/n3 ) );
  XOR \ADD_/FAINST[219].FA_/U2  ( .A(b[219]), .B(\ADD_/c[219] ), .Z(
        \ADD_/FAINST[219].FA_/n2 ) );
  XOR \ADD_/FAINST[219].FA_/U1  ( .A(a[219]), .B(\ADD_/c[219] ), .Z(
        \ADD_/FAINST[219].FA_/n1 ) );
  XOR \ADD_/FAINST[218].FA_/U5  ( .A(\ADD_/FAINST[218].FA_/n3 ), .B(
        \ADD_/c[218] ), .Z(\ADD_/c[219] ) );
  XOR \ADD_/FAINST[218].FA_/U4  ( .A(\ADD_/FAINST[218].FA_/n1 ), .B(b[218]), 
        .Z(c[218]) );
  AND \ADD_/FAINST[218].FA_/U3  ( .A(\ADD_/FAINST[218].FA_/n1 ), .B(
        \ADD_/FAINST[218].FA_/n2 ), .Z(\ADD_/FAINST[218].FA_/n3 ) );
  XOR \ADD_/FAINST[218].FA_/U2  ( .A(b[218]), .B(\ADD_/c[218] ), .Z(
        \ADD_/FAINST[218].FA_/n2 ) );
  XOR \ADD_/FAINST[218].FA_/U1  ( .A(a[218]), .B(\ADD_/c[218] ), .Z(
        \ADD_/FAINST[218].FA_/n1 ) );
  XOR \ADD_/FAINST[217].FA_/U5  ( .A(\ADD_/FAINST[217].FA_/n3 ), .B(
        \ADD_/c[217] ), .Z(\ADD_/c[218] ) );
  XOR \ADD_/FAINST[217].FA_/U4  ( .A(\ADD_/FAINST[217].FA_/n1 ), .B(b[217]), 
        .Z(c[217]) );
  AND \ADD_/FAINST[217].FA_/U3  ( .A(\ADD_/FAINST[217].FA_/n1 ), .B(
        \ADD_/FAINST[217].FA_/n2 ), .Z(\ADD_/FAINST[217].FA_/n3 ) );
  XOR \ADD_/FAINST[217].FA_/U2  ( .A(b[217]), .B(\ADD_/c[217] ), .Z(
        \ADD_/FAINST[217].FA_/n2 ) );
  XOR \ADD_/FAINST[217].FA_/U1  ( .A(a[217]), .B(\ADD_/c[217] ), .Z(
        \ADD_/FAINST[217].FA_/n1 ) );
  XOR \ADD_/FAINST[216].FA_/U5  ( .A(\ADD_/FAINST[216].FA_/n3 ), .B(
        \ADD_/c[216] ), .Z(\ADD_/c[217] ) );
  XOR \ADD_/FAINST[216].FA_/U4  ( .A(\ADD_/FAINST[216].FA_/n1 ), .B(b[216]), 
        .Z(c[216]) );
  AND \ADD_/FAINST[216].FA_/U3  ( .A(\ADD_/FAINST[216].FA_/n1 ), .B(
        \ADD_/FAINST[216].FA_/n2 ), .Z(\ADD_/FAINST[216].FA_/n3 ) );
  XOR \ADD_/FAINST[216].FA_/U2  ( .A(b[216]), .B(\ADD_/c[216] ), .Z(
        \ADD_/FAINST[216].FA_/n2 ) );
  XOR \ADD_/FAINST[216].FA_/U1  ( .A(a[216]), .B(\ADD_/c[216] ), .Z(
        \ADD_/FAINST[216].FA_/n1 ) );
  XOR \ADD_/FAINST[215].FA_/U5  ( .A(\ADD_/FAINST[215].FA_/n3 ), .B(
        \ADD_/c[215] ), .Z(\ADD_/c[216] ) );
  XOR \ADD_/FAINST[215].FA_/U4  ( .A(\ADD_/FAINST[215].FA_/n1 ), .B(b[215]), 
        .Z(c[215]) );
  AND \ADD_/FAINST[215].FA_/U3  ( .A(\ADD_/FAINST[215].FA_/n1 ), .B(
        \ADD_/FAINST[215].FA_/n2 ), .Z(\ADD_/FAINST[215].FA_/n3 ) );
  XOR \ADD_/FAINST[215].FA_/U2  ( .A(b[215]), .B(\ADD_/c[215] ), .Z(
        \ADD_/FAINST[215].FA_/n2 ) );
  XOR \ADD_/FAINST[215].FA_/U1  ( .A(a[215]), .B(\ADD_/c[215] ), .Z(
        \ADD_/FAINST[215].FA_/n1 ) );
  XOR \ADD_/FAINST[214].FA_/U5  ( .A(\ADD_/FAINST[214].FA_/n3 ), .B(
        \ADD_/c[214] ), .Z(\ADD_/c[215] ) );
  XOR \ADD_/FAINST[214].FA_/U4  ( .A(\ADD_/FAINST[214].FA_/n1 ), .B(b[214]), 
        .Z(c[214]) );
  AND \ADD_/FAINST[214].FA_/U3  ( .A(\ADD_/FAINST[214].FA_/n1 ), .B(
        \ADD_/FAINST[214].FA_/n2 ), .Z(\ADD_/FAINST[214].FA_/n3 ) );
  XOR \ADD_/FAINST[214].FA_/U2  ( .A(b[214]), .B(\ADD_/c[214] ), .Z(
        \ADD_/FAINST[214].FA_/n2 ) );
  XOR \ADD_/FAINST[214].FA_/U1  ( .A(a[214]), .B(\ADD_/c[214] ), .Z(
        \ADD_/FAINST[214].FA_/n1 ) );
  XOR \ADD_/FAINST[213].FA_/U5  ( .A(\ADD_/FAINST[213].FA_/n3 ), .B(
        \ADD_/c[213] ), .Z(\ADD_/c[214] ) );
  XOR \ADD_/FAINST[213].FA_/U4  ( .A(\ADD_/FAINST[213].FA_/n1 ), .B(b[213]), 
        .Z(c[213]) );
  AND \ADD_/FAINST[213].FA_/U3  ( .A(\ADD_/FAINST[213].FA_/n1 ), .B(
        \ADD_/FAINST[213].FA_/n2 ), .Z(\ADD_/FAINST[213].FA_/n3 ) );
  XOR \ADD_/FAINST[213].FA_/U2  ( .A(b[213]), .B(\ADD_/c[213] ), .Z(
        \ADD_/FAINST[213].FA_/n2 ) );
  XOR \ADD_/FAINST[213].FA_/U1  ( .A(a[213]), .B(\ADD_/c[213] ), .Z(
        \ADD_/FAINST[213].FA_/n1 ) );
  XOR \ADD_/FAINST[212].FA_/U5  ( .A(\ADD_/FAINST[212].FA_/n3 ), .B(
        \ADD_/c[212] ), .Z(\ADD_/c[213] ) );
  XOR \ADD_/FAINST[212].FA_/U4  ( .A(\ADD_/FAINST[212].FA_/n1 ), .B(b[212]), 
        .Z(c[212]) );
  AND \ADD_/FAINST[212].FA_/U3  ( .A(\ADD_/FAINST[212].FA_/n1 ), .B(
        \ADD_/FAINST[212].FA_/n2 ), .Z(\ADD_/FAINST[212].FA_/n3 ) );
  XOR \ADD_/FAINST[212].FA_/U2  ( .A(b[212]), .B(\ADD_/c[212] ), .Z(
        \ADD_/FAINST[212].FA_/n2 ) );
  XOR \ADD_/FAINST[212].FA_/U1  ( .A(a[212]), .B(\ADD_/c[212] ), .Z(
        \ADD_/FAINST[212].FA_/n1 ) );
  XOR \ADD_/FAINST[211].FA_/U5  ( .A(\ADD_/FAINST[211].FA_/n3 ), .B(
        \ADD_/c[211] ), .Z(\ADD_/c[212] ) );
  XOR \ADD_/FAINST[211].FA_/U4  ( .A(\ADD_/FAINST[211].FA_/n1 ), .B(b[211]), 
        .Z(c[211]) );
  AND \ADD_/FAINST[211].FA_/U3  ( .A(\ADD_/FAINST[211].FA_/n1 ), .B(
        \ADD_/FAINST[211].FA_/n2 ), .Z(\ADD_/FAINST[211].FA_/n3 ) );
  XOR \ADD_/FAINST[211].FA_/U2  ( .A(b[211]), .B(\ADD_/c[211] ), .Z(
        \ADD_/FAINST[211].FA_/n2 ) );
  XOR \ADD_/FAINST[211].FA_/U1  ( .A(a[211]), .B(\ADD_/c[211] ), .Z(
        \ADD_/FAINST[211].FA_/n1 ) );
  XOR \ADD_/FAINST[210].FA_/U5  ( .A(\ADD_/FAINST[210].FA_/n3 ), .B(
        \ADD_/c[210] ), .Z(\ADD_/c[211] ) );
  XOR \ADD_/FAINST[210].FA_/U4  ( .A(\ADD_/FAINST[210].FA_/n1 ), .B(b[210]), 
        .Z(c[210]) );
  AND \ADD_/FAINST[210].FA_/U3  ( .A(\ADD_/FAINST[210].FA_/n1 ), .B(
        \ADD_/FAINST[210].FA_/n2 ), .Z(\ADD_/FAINST[210].FA_/n3 ) );
  XOR \ADD_/FAINST[210].FA_/U2  ( .A(b[210]), .B(\ADD_/c[210] ), .Z(
        \ADD_/FAINST[210].FA_/n2 ) );
  XOR \ADD_/FAINST[210].FA_/U1  ( .A(a[210]), .B(\ADD_/c[210] ), .Z(
        \ADD_/FAINST[210].FA_/n1 ) );
  XOR \ADD_/FAINST[209].FA_/U5  ( .A(\ADD_/FAINST[209].FA_/n3 ), .B(
        \ADD_/c[209] ), .Z(\ADD_/c[210] ) );
  XOR \ADD_/FAINST[209].FA_/U4  ( .A(\ADD_/FAINST[209].FA_/n1 ), .B(b[209]), 
        .Z(c[209]) );
  AND \ADD_/FAINST[209].FA_/U3  ( .A(\ADD_/FAINST[209].FA_/n1 ), .B(
        \ADD_/FAINST[209].FA_/n2 ), .Z(\ADD_/FAINST[209].FA_/n3 ) );
  XOR \ADD_/FAINST[209].FA_/U2  ( .A(b[209]), .B(\ADD_/c[209] ), .Z(
        \ADD_/FAINST[209].FA_/n2 ) );
  XOR \ADD_/FAINST[209].FA_/U1  ( .A(a[209]), .B(\ADD_/c[209] ), .Z(
        \ADD_/FAINST[209].FA_/n1 ) );
  XOR \ADD_/FAINST[208].FA_/U5  ( .A(\ADD_/FAINST[208].FA_/n3 ), .B(
        \ADD_/c[208] ), .Z(\ADD_/c[209] ) );
  XOR \ADD_/FAINST[208].FA_/U4  ( .A(\ADD_/FAINST[208].FA_/n1 ), .B(b[208]), 
        .Z(c[208]) );
  AND \ADD_/FAINST[208].FA_/U3  ( .A(\ADD_/FAINST[208].FA_/n1 ), .B(
        \ADD_/FAINST[208].FA_/n2 ), .Z(\ADD_/FAINST[208].FA_/n3 ) );
  XOR \ADD_/FAINST[208].FA_/U2  ( .A(b[208]), .B(\ADD_/c[208] ), .Z(
        \ADD_/FAINST[208].FA_/n2 ) );
  XOR \ADD_/FAINST[208].FA_/U1  ( .A(a[208]), .B(\ADD_/c[208] ), .Z(
        \ADD_/FAINST[208].FA_/n1 ) );
  XOR \ADD_/FAINST[207].FA_/U5  ( .A(\ADD_/FAINST[207].FA_/n3 ), .B(
        \ADD_/c[207] ), .Z(\ADD_/c[208] ) );
  XOR \ADD_/FAINST[207].FA_/U4  ( .A(\ADD_/FAINST[207].FA_/n1 ), .B(b[207]), 
        .Z(c[207]) );
  AND \ADD_/FAINST[207].FA_/U3  ( .A(\ADD_/FAINST[207].FA_/n1 ), .B(
        \ADD_/FAINST[207].FA_/n2 ), .Z(\ADD_/FAINST[207].FA_/n3 ) );
  XOR \ADD_/FAINST[207].FA_/U2  ( .A(b[207]), .B(\ADD_/c[207] ), .Z(
        \ADD_/FAINST[207].FA_/n2 ) );
  XOR \ADD_/FAINST[207].FA_/U1  ( .A(a[207]), .B(\ADD_/c[207] ), .Z(
        \ADD_/FAINST[207].FA_/n1 ) );
  XOR \ADD_/FAINST[206].FA_/U5  ( .A(\ADD_/FAINST[206].FA_/n3 ), .B(
        \ADD_/c[206] ), .Z(\ADD_/c[207] ) );
  XOR \ADD_/FAINST[206].FA_/U4  ( .A(\ADD_/FAINST[206].FA_/n1 ), .B(b[206]), 
        .Z(c[206]) );
  AND \ADD_/FAINST[206].FA_/U3  ( .A(\ADD_/FAINST[206].FA_/n1 ), .B(
        \ADD_/FAINST[206].FA_/n2 ), .Z(\ADD_/FAINST[206].FA_/n3 ) );
  XOR \ADD_/FAINST[206].FA_/U2  ( .A(b[206]), .B(\ADD_/c[206] ), .Z(
        \ADD_/FAINST[206].FA_/n2 ) );
  XOR \ADD_/FAINST[206].FA_/U1  ( .A(a[206]), .B(\ADD_/c[206] ), .Z(
        \ADD_/FAINST[206].FA_/n1 ) );
  XOR \ADD_/FAINST[205].FA_/U5  ( .A(\ADD_/FAINST[205].FA_/n3 ), .B(
        \ADD_/c[205] ), .Z(\ADD_/c[206] ) );
  XOR \ADD_/FAINST[205].FA_/U4  ( .A(\ADD_/FAINST[205].FA_/n1 ), .B(b[205]), 
        .Z(c[205]) );
  AND \ADD_/FAINST[205].FA_/U3  ( .A(\ADD_/FAINST[205].FA_/n1 ), .B(
        \ADD_/FAINST[205].FA_/n2 ), .Z(\ADD_/FAINST[205].FA_/n3 ) );
  XOR \ADD_/FAINST[205].FA_/U2  ( .A(b[205]), .B(\ADD_/c[205] ), .Z(
        \ADD_/FAINST[205].FA_/n2 ) );
  XOR \ADD_/FAINST[205].FA_/U1  ( .A(a[205]), .B(\ADD_/c[205] ), .Z(
        \ADD_/FAINST[205].FA_/n1 ) );
  XOR \ADD_/FAINST[204].FA_/U5  ( .A(\ADD_/FAINST[204].FA_/n3 ), .B(
        \ADD_/c[204] ), .Z(\ADD_/c[205] ) );
  XOR \ADD_/FAINST[204].FA_/U4  ( .A(\ADD_/FAINST[204].FA_/n1 ), .B(b[204]), 
        .Z(c[204]) );
  AND \ADD_/FAINST[204].FA_/U3  ( .A(\ADD_/FAINST[204].FA_/n1 ), .B(
        \ADD_/FAINST[204].FA_/n2 ), .Z(\ADD_/FAINST[204].FA_/n3 ) );
  XOR \ADD_/FAINST[204].FA_/U2  ( .A(b[204]), .B(\ADD_/c[204] ), .Z(
        \ADD_/FAINST[204].FA_/n2 ) );
  XOR \ADD_/FAINST[204].FA_/U1  ( .A(a[204]), .B(\ADD_/c[204] ), .Z(
        \ADD_/FAINST[204].FA_/n1 ) );
  XOR \ADD_/FAINST[203].FA_/U5  ( .A(\ADD_/FAINST[203].FA_/n3 ), .B(
        \ADD_/c[203] ), .Z(\ADD_/c[204] ) );
  XOR \ADD_/FAINST[203].FA_/U4  ( .A(\ADD_/FAINST[203].FA_/n1 ), .B(b[203]), 
        .Z(c[203]) );
  AND \ADD_/FAINST[203].FA_/U3  ( .A(\ADD_/FAINST[203].FA_/n1 ), .B(
        \ADD_/FAINST[203].FA_/n2 ), .Z(\ADD_/FAINST[203].FA_/n3 ) );
  XOR \ADD_/FAINST[203].FA_/U2  ( .A(b[203]), .B(\ADD_/c[203] ), .Z(
        \ADD_/FAINST[203].FA_/n2 ) );
  XOR \ADD_/FAINST[203].FA_/U1  ( .A(a[203]), .B(\ADD_/c[203] ), .Z(
        \ADD_/FAINST[203].FA_/n1 ) );
  XOR \ADD_/FAINST[202].FA_/U5  ( .A(\ADD_/FAINST[202].FA_/n3 ), .B(
        \ADD_/c[202] ), .Z(\ADD_/c[203] ) );
  XOR \ADD_/FAINST[202].FA_/U4  ( .A(\ADD_/FAINST[202].FA_/n1 ), .B(b[202]), 
        .Z(c[202]) );
  AND \ADD_/FAINST[202].FA_/U3  ( .A(\ADD_/FAINST[202].FA_/n1 ), .B(
        \ADD_/FAINST[202].FA_/n2 ), .Z(\ADD_/FAINST[202].FA_/n3 ) );
  XOR \ADD_/FAINST[202].FA_/U2  ( .A(b[202]), .B(\ADD_/c[202] ), .Z(
        \ADD_/FAINST[202].FA_/n2 ) );
  XOR \ADD_/FAINST[202].FA_/U1  ( .A(a[202]), .B(\ADD_/c[202] ), .Z(
        \ADD_/FAINST[202].FA_/n1 ) );
  XOR \ADD_/FAINST[201].FA_/U5  ( .A(\ADD_/FAINST[201].FA_/n3 ), .B(
        \ADD_/c[201] ), .Z(\ADD_/c[202] ) );
  XOR \ADD_/FAINST[201].FA_/U4  ( .A(\ADD_/FAINST[201].FA_/n1 ), .B(b[201]), 
        .Z(c[201]) );
  AND \ADD_/FAINST[201].FA_/U3  ( .A(\ADD_/FAINST[201].FA_/n1 ), .B(
        \ADD_/FAINST[201].FA_/n2 ), .Z(\ADD_/FAINST[201].FA_/n3 ) );
  XOR \ADD_/FAINST[201].FA_/U2  ( .A(b[201]), .B(\ADD_/c[201] ), .Z(
        \ADD_/FAINST[201].FA_/n2 ) );
  XOR \ADD_/FAINST[201].FA_/U1  ( .A(a[201]), .B(\ADD_/c[201] ), .Z(
        \ADD_/FAINST[201].FA_/n1 ) );
  XOR \ADD_/FAINST[200].FA_/U5  ( .A(\ADD_/FAINST[200].FA_/n3 ), .B(
        \ADD_/c[200] ), .Z(\ADD_/c[201] ) );
  XOR \ADD_/FAINST[200].FA_/U4  ( .A(\ADD_/FAINST[200].FA_/n1 ), .B(b[200]), 
        .Z(c[200]) );
  AND \ADD_/FAINST[200].FA_/U3  ( .A(\ADD_/FAINST[200].FA_/n1 ), .B(
        \ADD_/FAINST[200].FA_/n2 ), .Z(\ADD_/FAINST[200].FA_/n3 ) );
  XOR \ADD_/FAINST[200].FA_/U2  ( .A(b[200]), .B(\ADD_/c[200] ), .Z(
        \ADD_/FAINST[200].FA_/n2 ) );
  XOR \ADD_/FAINST[200].FA_/U1  ( .A(a[200]), .B(\ADD_/c[200] ), .Z(
        \ADD_/FAINST[200].FA_/n1 ) );
  XOR \ADD_/FAINST[199].FA_/U5  ( .A(\ADD_/FAINST[199].FA_/n3 ), .B(
        \ADD_/c[199] ), .Z(\ADD_/c[200] ) );
  XOR \ADD_/FAINST[199].FA_/U4  ( .A(\ADD_/FAINST[199].FA_/n1 ), .B(b[199]), 
        .Z(c[199]) );
  AND \ADD_/FAINST[199].FA_/U3  ( .A(\ADD_/FAINST[199].FA_/n1 ), .B(
        \ADD_/FAINST[199].FA_/n2 ), .Z(\ADD_/FAINST[199].FA_/n3 ) );
  XOR \ADD_/FAINST[199].FA_/U2  ( .A(b[199]), .B(\ADD_/c[199] ), .Z(
        \ADD_/FAINST[199].FA_/n2 ) );
  XOR \ADD_/FAINST[199].FA_/U1  ( .A(a[199]), .B(\ADD_/c[199] ), .Z(
        \ADD_/FAINST[199].FA_/n1 ) );
  XOR \ADD_/FAINST[198].FA_/U5  ( .A(\ADD_/FAINST[198].FA_/n3 ), .B(
        \ADD_/c[198] ), .Z(\ADD_/c[199] ) );
  XOR \ADD_/FAINST[198].FA_/U4  ( .A(\ADD_/FAINST[198].FA_/n1 ), .B(b[198]), 
        .Z(c[198]) );
  AND \ADD_/FAINST[198].FA_/U3  ( .A(\ADD_/FAINST[198].FA_/n1 ), .B(
        \ADD_/FAINST[198].FA_/n2 ), .Z(\ADD_/FAINST[198].FA_/n3 ) );
  XOR \ADD_/FAINST[198].FA_/U2  ( .A(b[198]), .B(\ADD_/c[198] ), .Z(
        \ADD_/FAINST[198].FA_/n2 ) );
  XOR \ADD_/FAINST[198].FA_/U1  ( .A(a[198]), .B(\ADD_/c[198] ), .Z(
        \ADD_/FAINST[198].FA_/n1 ) );
  XOR \ADD_/FAINST[197].FA_/U5  ( .A(\ADD_/FAINST[197].FA_/n3 ), .B(
        \ADD_/c[197] ), .Z(\ADD_/c[198] ) );
  XOR \ADD_/FAINST[197].FA_/U4  ( .A(\ADD_/FAINST[197].FA_/n1 ), .B(b[197]), 
        .Z(c[197]) );
  AND \ADD_/FAINST[197].FA_/U3  ( .A(\ADD_/FAINST[197].FA_/n1 ), .B(
        \ADD_/FAINST[197].FA_/n2 ), .Z(\ADD_/FAINST[197].FA_/n3 ) );
  XOR \ADD_/FAINST[197].FA_/U2  ( .A(b[197]), .B(\ADD_/c[197] ), .Z(
        \ADD_/FAINST[197].FA_/n2 ) );
  XOR \ADD_/FAINST[197].FA_/U1  ( .A(a[197]), .B(\ADD_/c[197] ), .Z(
        \ADD_/FAINST[197].FA_/n1 ) );
  XOR \ADD_/FAINST[196].FA_/U5  ( .A(\ADD_/FAINST[196].FA_/n3 ), .B(
        \ADD_/c[196] ), .Z(\ADD_/c[197] ) );
  XOR \ADD_/FAINST[196].FA_/U4  ( .A(\ADD_/FAINST[196].FA_/n1 ), .B(b[196]), 
        .Z(c[196]) );
  AND \ADD_/FAINST[196].FA_/U3  ( .A(\ADD_/FAINST[196].FA_/n1 ), .B(
        \ADD_/FAINST[196].FA_/n2 ), .Z(\ADD_/FAINST[196].FA_/n3 ) );
  XOR \ADD_/FAINST[196].FA_/U2  ( .A(b[196]), .B(\ADD_/c[196] ), .Z(
        \ADD_/FAINST[196].FA_/n2 ) );
  XOR \ADD_/FAINST[196].FA_/U1  ( .A(a[196]), .B(\ADD_/c[196] ), .Z(
        \ADD_/FAINST[196].FA_/n1 ) );
  XOR \ADD_/FAINST[195].FA_/U5  ( .A(\ADD_/FAINST[195].FA_/n3 ), .B(
        \ADD_/c[195] ), .Z(\ADD_/c[196] ) );
  XOR \ADD_/FAINST[195].FA_/U4  ( .A(\ADD_/FAINST[195].FA_/n1 ), .B(b[195]), 
        .Z(c[195]) );
  AND \ADD_/FAINST[195].FA_/U3  ( .A(\ADD_/FAINST[195].FA_/n1 ), .B(
        \ADD_/FAINST[195].FA_/n2 ), .Z(\ADD_/FAINST[195].FA_/n3 ) );
  XOR \ADD_/FAINST[195].FA_/U2  ( .A(b[195]), .B(\ADD_/c[195] ), .Z(
        \ADD_/FAINST[195].FA_/n2 ) );
  XOR \ADD_/FAINST[195].FA_/U1  ( .A(a[195]), .B(\ADD_/c[195] ), .Z(
        \ADD_/FAINST[195].FA_/n1 ) );
  XOR \ADD_/FAINST[194].FA_/U5  ( .A(\ADD_/FAINST[194].FA_/n3 ), .B(
        \ADD_/c[194] ), .Z(\ADD_/c[195] ) );
  XOR \ADD_/FAINST[194].FA_/U4  ( .A(\ADD_/FAINST[194].FA_/n1 ), .B(b[194]), 
        .Z(c[194]) );
  AND \ADD_/FAINST[194].FA_/U3  ( .A(\ADD_/FAINST[194].FA_/n1 ), .B(
        \ADD_/FAINST[194].FA_/n2 ), .Z(\ADD_/FAINST[194].FA_/n3 ) );
  XOR \ADD_/FAINST[194].FA_/U2  ( .A(b[194]), .B(\ADD_/c[194] ), .Z(
        \ADD_/FAINST[194].FA_/n2 ) );
  XOR \ADD_/FAINST[194].FA_/U1  ( .A(a[194]), .B(\ADD_/c[194] ), .Z(
        \ADD_/FAINST[194].FA_/n1 ) );
  XOR \ADD_/FAINST[193].FA_/U5  ( .A(\ADD_/FAINST[193].FA_/n3 ), .B(
        \ADD_/c[193] ), .Z(\ADD_/c[194] ) );
  XOR \ADD_/FAINST[193].FA_/U4  ( .A(\ADD_/FAINST[193].FA_/n1 ), .B(b[193]), 
        .Z(c[193]) );
  AND \ADD_/FAINST[193].FA_/U3  ( .A(\ADD_/FAINST[193].FA_/n1 ), .B(
        \ADD_/FAINST[193].FA_/n2 ), .Z(\ADD_/FAINST[193].FA_/n3 ) );
  XOR \ADD_/FAINST[193].FA_/U2  ( .A(b[193]), .B(\ADD_/c[193] ), .Z(
        \ADD_/FAINST[193].FA_/n2 ) );
  XOR \ADD_/FAINST[193].FA_/U1  ( .A(a[193]), .B(\ADD_/c[193] ), .Z(
        \ADD_/FAINST[193].FA_/n1 ) );
  XOR \ADD_/FAINST[192].FA_/U5  ( .A(\ADD_/FAINST[192].FA_/n3 ), .B(
        \ADD_/c[192] ), .Z(\ADD_/c[193] ) );
  XOR \ADD_/FAINST[192].FA_/U4  ( .A(\ADD_/FAINST[192].FA_/n1 ), .B(b[192]), 
        .Z(c[192]) );
  AND \ADD_/FAINST[192].FA_/U3  ( .A(\ADD_/FAINST[192].FA_/n1 ), .B(
        \ADD_/FAINST[192].FA_/n2 ), .Z(\ADD_/FAINST[192].FA_/n3 ) );
  XOR \ADD_/FAINST[192].FA_/U2  ( .A(b[192]), .B(\ADD_/c[192] ), .Z(
        \ADD_/FAINST[192].FA_/n2 ) );
  XOR \ADD_/FAINST[192].FA_/U1  ( .A(a[192]), .B(\ADD_/c[192] ), .Z(
        \ADD_/FAINST[192].FA_/n1 ) );
  XOR \ADD_/FAINST[191].FA_/U5  ( .A(\ADD_/FAINST[191].FA_/n3 ), .B(
        \ADD_/c[191] ), .Z(\ADD_/c[192] ) );
  XOR \ADD_/FAINST[191].FA_/U4  ( .A(\ADD_/FAINST[191].FA_/n1 ), .B(b[191]), 
        .Z(c[191]) );
  AND \ADD_/FAINST[191].FA_/U3  ( .A(\ADD_/FAINST[191].FA_/n1 ), .B(
        \ADD_/FAINST[191].FA_/n2 ), .Z(\ADD_/FAINST[191].FA_/n3 ) );
  XOR \ADD_/FAINST[191].FA_/U2  ( .A(b[191]), .B(\ADD_/c[191] ), .Z(
        \ADD_/FAINST[191].FA_/n2 ) );
  XOR \ADD_/FAINST[191].FA_/U1  ( .A(a[191]), .B(\ADD_/c[191] ), .Z(
        \ADD_/FAINST[191].FA_/n1 ) );
  XOR \ADD_/FAINST[190].FA_/U5  ( .A(\ADD_/FAINST[190].FA_/n3 ), .B(
        \ADD_/c[190] ), .Z(\ADD_/c[191] ) );
  XOR \ADD_/FAINST[190].FA_/U4  ( .A(\ADD_/FAINST[190].FA_/n1 ), .B(b[190]), 
        .Z(c[190]) );
  AND \ADD_/FAINST[190].FA_/U3  ( .A(\ADD_/FAINST[190].FA_/n1 ), .B(
        \ADD_/FAINST[190].FA_/n2 ), .Z(\ADD_/FAINST[190].FA_/n3 ) );
  XOR \ADD_/FAINST[190].FA_/U2  ( .A(b[190]), .B(\ADD_/c[190] ), .Z(
        \ADD_/FAINST[190].FA_/n2 ) );
  XOR \ADD_/FAINST[190].FA_/U1  ( .A(a[190]), .B(\ADD_/c[190] ), .Z(
        \ADD_/FAINST[190].FA_/n1 ) );
  XOR \ADD_/FAINST[189].FA_/U5  ( .A(\ADD_/FAINST[189].FA_/n3 ), .B(
        \ADD_/c[189] ), .Z(\ADD_/c[190] ) );
  XOR \ADD_/FAINST[189].FA_/U4  ( .A(\ADD_/FAINST[189].FA_/n1 ), .B(b[189]), 
        .Z(c[189]) );
  AND \ADD_/FAINST[189].FA_/U3  ( .A(\ADD_/FAINST[189].FA_/n1 ), .B(
        \ADD_/FAINST[189].FA_/n2 ), .Z(\ADD_/FAINST[189].FA_/n3 ) );
  XOR \ADD_/FAINST[189].FA_/U2  ( .A(b[189]), .B(\ADD_/c[189] ), .Z(
        \ADD_/FAINST[189].FA_/n2 ) );
  XOR \ADD_/FAINST[189].FA_/U1  ( .A(a[189]), .B(\ADD_/c[189] ), .Z(
        \ADD_/FAINST[189].FA_/n1 ) );
  XOR \ADD_/FAINST[188].FA_/U5  ( .A(\ADD_/FAINST[188].FA_/n3 ), .B(
        \ADD_/c[188] ), .Z(\ADD_/c[189] ) );
  XOR \ADD_/FAINST[188].FA_/U4  ( .A(\ADD_/FAINST[188].FA_/n1 ), .B(b[188]), 
        .Z(c[188]) );
  AND \ADD_/FAINST[188].FA_/U3  ( .A(\ADD_/FAINST[188].FA_/n1 ), .B(
        \ADD_/FAINST[188].FA_/n2 ), .Z(\ADD_/FAINST[188].FA_/n3 ) );
  XOR \ADD_/FAINST[188].FA_/U2  ( .A(b[188]), .B(\ADD_/c[188] ), .Z(
        \ADD_/FAINST[188].FA_/n2 ) );
  XOR \ADD_/FAINST[188].FA_/U1  ( .A(a[188]), .B(\ADD_/c[188] ), .Z(
        \ADD_/FAINST[188].FA_/n1 ) );
  XOR \ADD_/FAINST[187].FA_/U5  ( .A(\ADD_/FAINST[187].FA_/n3 ), .B(
        \ADD_/c[187] ), .Z(\ADD_/c[188] ) );
  XOR \ADD_/FAINST[187].FA_/U4  ( .A(\ADD_/FAINST[187].FA_/n1 ), .B(b[187]), 
        .Z(c[187]) );
  AND \ADD_/FAINST[187].FA_/U3  ( .A(\ADD_/FAINST[187].FA_/n1 ), .B(
        \ADD_/FAINST[187].FA_/n2 ), .Z(\ADD_/FAINST[187].FA_/n3 ) );
  XOR \ADD_/FAINST[187].FA_/U2  ( .A(b[187]), .B(\ADD_/c[187] ), .Z(
        \ADD_/FAINST[187].FA_/n2 ) );
  XOR \ADD_/FAINST[187].FA_/U1  ( .A(a[187]), .B(\ADD_/c[187] ), .Z(
        \ADD_/FAINST[187].FA_/n1 ) );
  XOR \ADD_/FAINST[186].FA_/U5  ( .A(\ADD_/FAINST[186].FA_/n3 ), .B(
        \ADD_/c[186] ), .Z(\ADD_/c[187] ) );
  XOR \ADD_/FAINST[186].FA_/U4  ( .A(\ADD_/FAINST[186].FA_/n1 ), .B(b[186]), 
        .Z(c[186]) );
  AND \ADD_/FAINST[186].FA_/U3  ( .A(\ADD_/FAINST[186].FA_/n1 ), .B(
        \ADD_/FAINST[186].FA_/n2 ), .Z(\ADD_/FAINST[186].FA_/n3 ) );
  XOR \ADD_/FAINST[186].FA_/U2  ( .A(b[186]), .B(\ADD_/c[186] ), .Z(
        \ADD_/FAINST[186].FA_/n2 ) );
  XOR \ADD_/FAINST[186].FA_/U1  ( .A(a[186]), .B(\ADD_/c[186] ), .Z(
        \ADD_/FAINST[186].FA_/n1 ) );
  XOR \ADD_/FAINST[185].FA_/U5  ( .A(\ADD_/FAINST[185].FA_/n3 ), .B(
        \ADD_/c[185] ), .Z(\ADD_/c[186] ) );
  XOR \ADD_/FAINST[185].FA_/U4  ( .A(\ADD_/FAINST[185].FA_/n1 ), .B(b[185]), 
        .Z(c[185]) );
  AND \ADD_/FAINST[185].FA_/U3  ( .A(\ADD_/FAINST[185].FA_/n1 ), .B(
        \ADD_/FAINST[185].FA_/n2 ), .Z(\ADD_/FAINST[185].FA_/n3 ) );
  XOR \ADD_/FAINST[185].FA_/U2  ( .A(b[185]), .B(\ADD_/c[185] ), .Z(
        \ADD_/FAINST[185].FA_/n2 ) );
  XOR \ADD_/FAINST[185].FA_/U1  ( .A(a[185]), .B(\ADD_/c[185] ), .Z(
        \ADD_/FAINST[185].FA_/n1 ) );
  XOR \ADD_/FAINST[184].FA_/U5  ( .A(\ADD_/FAINST[184].FA_/n3 ), .B(
        \ADD_/c[184] ), .Z(\ADD_/c[185] ) );
  XOR \ADD_/FAINST[184].FA_/U4  ( .A(\ADD_/FAINST[184].FA_/n1 ), .B(b[184]), 
        .Z(c[184]) );
  AND \ADD_/FAINST[184].FA_/U3  ( .A(\ADD_/FAINST[184].FA_/n1 ), .B(
        \ADD_/FAINST[184].FA_/n2 ), .Z(\ADD_/FAINST[184].FA_/n3 ) );
  XOR \ADD_/FAINST[184].FA_/U2  ( .A(b[184]), .B(\ADD_/c[184] ), .Z(
        \ADD_/FAINST[184].FA_/n2 ) );
  XOR \ADD_/FAINST[184].FA_/U1  ( .A(a[184]), .B(\ADD_/c[184] ), .Z(
        \ADD_/FAINST[184].FA_/n1 ) );
  XOR \ADD_/FAINST[183].FA_/U5  ( .A(\ADD_/FAINST[183].FA_/n3 ), .B(
        \ADD_/c[183] ), .Z(\ADD_/c[184] ) );
  XOR \ADD_/FAINST[183].FA_/U4  ( .A(\ADD_/FAINST[183].FA_/n1 ), .B(b[183]), 
        .Z(c[183]) );
  AND \ADD_/FAINST[183].FA_/U3  ( .A(\ADD_/FAINST[183].FA_/n1 ), .B(
        \ADD_/FAINST[183].FA_/n2 ), .Z(\ADD_/FAINST[183].FA_/n3 ) );
  XOR \ADD_/FAINST[183].FA_/U2  ( .A(b[183]), .B(\ADD_/c[183] ), .Z(
        \ADD_/FAINST[183].FA_/n2 ) );
  XOR \ADD_/FAINST[183].FA_/U1  ( .A(a[183]), .B(\ADD_/c[183] ), .Z(
        \ADD_/FAINST[183].FA_/n1 ) );
  XOR \ADD_/FAINST[182].FA_/U5  ( .A(\ADD_/FAINST[182].FA_/n3 ), .B(
        \ADD_/c[182] ), .Z(\ADD_/c[183] ) );
  XOR \ADD_/FAINST[182].FA_/U4  ( .A(\ADD_/FAINST[182].FA_/n1 ), .B(b[182]), 
        .Z(c[182]) );
  AND \ADD_/FAINST[182].FA_/U3  ( .A(\ADD_/FAINST[182].FA_/n1 ), .B(
        \ADD_/FAINST[182].FA_/n2 ), .Z(\ADD_/FAINST[182].FA_/n3 ) );
  XOR \ADD_/FAINST[182].FA_/U2  ( .A(b[182]), .B(\ADD_/c[182] ), .Z(
        \ADD_/FAINST[182].FA_/n2 ) );
  XOR \ADD_/FAINST[182].FA_/U1  ( .A(a[182]), .B(\ADD_/c[182] ), .Z(
        \ADD_/FAINST[182].FA_/n1 ) );
  XOR \ADD_/FAINST[181].FA_/U5  ( .A(\ADD_/FAINST[181].FA_/n3 ), .B(
        \ADD_/c[181] ), .Z(\ADD_/c[182] ) );
  XOR \ADD_/FAINST[181].FA_/U4  ( .A(\ADD_/FAINST[181].FA_/n1 ), .B(b[181]), 
        .Z(c[181]) );
  AND \ADD_/FAINST[181].FA_/U3  ( .A(\ADD_/FAINST[181].FA_/n1 ), .B(
        \ADD_/FAINST[181].FA_/n2 ), .Z(\ADD_/FAINST[181].FA_/n3 ) );
  XOR \ADD_/FAINST[181].FA_/U2  ( .A(b[181]), .B(\ADD_/c[181] ), .Z(
        \ADD_/FAINST[181].FA_/n2 ) );
  XOR \ADD_/FAINST[181].FA_/U1  ( .A(a[181]), .B(\ADD_/c[181] ), .Z(
        \ADD_/FAINST[181].FA_/n1 ) );
  XOR \ADD_/FAINST[180].FA_/U5  ( .A(\ADD_/FAINST[180].FA_/n3 ), .B(
        \ADD_/c[180] ), .Z(\ADD_/c[181] ) );
  XOR \ADD_/FAINST[180].FA_/U4  ( .A(\ADD_/FAINST[180].FA_/n1 ), .B(b[180]), 
        .Z(c[180]) );
  AND \ADD_/FAINST[180].FA_/U3  ( .A(\ADD_/FAINST[180].FA_/n1 ), .B(
        \ADD_/FAINST[180].FA_/n2 ), .Z(\ADD_/FAINST[180].FA_/n3 ) );
  XOR \ADD_/FAINST[180].FA_/U2  ( .A(b[180]), .B(\ADD_/c[180] ), .Z(
        \ADD_/FAINST[180].FA_/n2 ) );
  XOR \ADD_/FAINST[180].FA_/U1  ( .A(a[180]), .B(\ADD_/c[180] ), .Z(
        \ADD_/FAINST[180].FA_/n1 ) );
  XOR \ADD_/FAINST[179].FA_/U5  ( .A(\ADD_/FAINST[179].FA_/n3 ), .B(
        \ADD_/c[179] ), .Z(\ADD_/c[180] ) );
  XOR \ADD_/FAINST[179].FA_/U4  ( .A(\ADD_/FAINST[179].FA_/n1 ), .B(b[179]), 
        .Z(c[179]) );
  AND \ADD_/FAINST[179].FA_/U3  ( .A(\ADD_/FAINST[179].FA_/n1 ), .B(
        \ADD_/FAINST[179].FA_/n2 ), .Z(\ADD_/FAINST[179].FA_/n3 ) );
  XOR \ADD_/FAINST[179].FA_/U2  ( .A(b[179]), .B(\ADD_/c[179] ), .Z(
        \ADD_/FAINST[179].FA_/n2 ) );
  XOR \ADD_/FAINST[179].FA_/U1  ( .A(a[179]), .B(\ADD_/c[179] ), .Z(
        \ADD_/FAINST[179].FA_/n1 ) );
  XOR \ADD_/FAINST[178].FA_/U5  ( .A(\ADD_/FAINST[178].FA_/n3 ), .B(
        \ADD_/c[178] ), .Z(\ADD_/c[179] ) );
  XOR \ADD_/FAINST[178].FA_/U4  ( .A(\ADD_/FAINST[178].FA_/n1 ), .B(b[178]), 
        .Z(c[178]) );
  AND \ADD_/FAINST[178].FA_/U3  ( .A(\ADD_/FAINST[178].FA_/n1 ), .B(
        \ADD_/FAINST[178].FA_/n2 ), .Z(\ADD_/FAINST[178].FA_/n3 ) );
  XOR \ADD_/FAINST[178].FA_/U2  ( .A(b[178]), .B(\ADD_/c[178] ), .Z(
        \ADD_/FAINST[178].FA_/n2 ) );
  XOR \ADD_/FAINST[178].FA_/U1  ( .A(a[178]), .B(\ADD_/c[178] ), .Z(
        \ADD_/FAINST[178].FA_/n1 ) );
  XOR \ADD_/FAINST[177].FA_/U5  ( .A(\ADD_/FAINST[177].FA_/n3 ), .B(
        \ADD_/c[177] ), .Z(\ADD_/c[178] ) );
  XOR \ADD_/FAINST[177].FA_/U4  ( .A(\ADD_/FAINST[177].FA_/n1 ), .B(b[177]), 
        .Z(c[177]) );
  AND \ADD_/FAINST[177].FA_/U3  ( .A(\ADD_/FAINST[177].FA_/n1 ), .B(
        \ADD_/FAINST[177].FA_/n2 ), .Z(\ADD_/FAINST[177].FA_/n3 ) );
  XOR \ADD_/FAINST[177].FA_/U2  ( .A(b[177]), .B(\ADD_/c[177] ), .Z(
        \ADD_/FAINST[177].FA_/n2 ) );
  XOR \ADD_/FAINST[177].FA_/U1  ( .A(a[177]), .B(\ADD_/c[177] ), .Z(
        \ADD_/FAINST[177].FA_/n1 ) );
  XOR \ADD_/FAINST[176].FA_/U5  ( .A(\ADD_/FAINST[176].FA_/n3 ), .B(
        \ADD_/c[176] ), .Z(\ADD_/c[177] ) );
  XOR \ADD_/FAINST[176].FA_/U4  ( .A(\ADD_/FAINST[176].FA_/n1 ), .B(b[176]), 
        .Z(c[176]) );
  AND \ADD_/FAINST[176].FA_/U3  ( .A(\ADD_/FAINST[176].FA_/n1 ), .B(
        \ADD_/FAINST[176].FA_/n2 ), .Z(\ADD_/FAINST[176].FA_/n3 ) );
  XOR \ADD_/FAINST[176].FA_/U2  ( .A(b[176]), .B(\ADD_/c[176] ), .Z(
        \ADD_/FAINST[176].FA_/n2 ) );
  XOR \ADD_/FAINST[176].FA_/U1  ( .A(a[176]), .B(\ADD_/c[176] ), .Z(
        \ADD_/FAINST[176].FA_/n1 ) );
  XOR \ADD_/FAINST[175].FA_/U5  ( .A(\ADD_/FAINST[175].FA_/n3 ), .B(
        \ADD_/c[175] ), .Z(\ADD_/c[176] ) );
  XOR \ADD_/FAINST[175].FA_/U4  ( .A(\ADD_/FAINST[175].FA_/n1 ), .B(b[175]), 
        .Z(c[175]) );
  AND \ADD_/FAINST[175].FA_/U3  ( .A(\ADD_/FAINST[175].FA_/n1 ), .B(
        \ADD_/FAINST[175].FA_/n2 ), .Z(\ADD_/FAINST[175].FA_/n3 ) );
  XOR \ADD_/FAINST[175].FA_/U2  ( .A(b[175]), .B(\ADD_/c[175] ), .Z(
        \ADD_/FAINST[175].FA_/n2 ) );
  XOR \ADD_/FAINST[175].FA_/U1  ( .A(a[175]), .B(\ADD_/c[175] ), .Z(
        \ADD_/FAINST[175].FA_/n1 ) );
  XOR \ADD_/FAINST[174].FA_/U5  ( .A(\ADD_/FAINST[174].FA_/n3 ), .B(
        \ADD_/c[174] ), .Z(\ADD_/c[175] ) );
  XOR \ADD_/FAINST[174].FA_/U4  ( .A(\ADD_/FAINST[174].FA_/n1 ), .B(b[174]), 
        .Z(c[174]) );
  AND \ADD_/FAINST[174].FA_/U3  ( .A(\ADD_/FAINST[174].FA_/n1 ), .B(
        \ADD_/FAINST[174].FA_/n2 ), .Z(\ADD_/FAINST[174].FA_/n3 ) );
  XOR \ADD_/FAINST[174].FA_/U2  ( .A(b[174]), .B(\ADD_/c[174] ), .Z(
        \ADD_/FAINST[174].FA_/n2 ) );
  XOR \ADD_/FAINST[174].FA_/U1  ( .A(a[174]), .B(\ADD_/c[174] ), .Z(
        \ADD_/FAINST[174].FA_/n1 ) );
  XOR \ADD_/FAINST[173].FA_/U5  ( .A(\ADD_/FAINST[173].FA_/n3 ), .B(
        \ADD_/c[173] ), .Z(\ADD_/c[174] ) );
  XOR \ADD_/FAINST[173].FA_/U4  ( .A(\ADD_/FAINST[173].FA_/n1 ), .B(b[173]), 
        .Z(c[173]) );
  AND \ADD_/FAINST[173].FA_/U3  ( .A(\ADD_/FAINST[173].FA_/n1 ), .B(
        \ADD_/FAINST[173].FA_/n2 ), .Z(\ADD_/FAINST[173].FA_/n3 ) );
  XOR \ADD_/FAINST[173].FA_/U2  ( .A(b[173]), .B(\ADD_/c[173] ), .Z(
        \ADD_/FAINST[173].FA_/n2 ) );
  XOR \ADD_/FAINST[173].FA_/U1  ( .A(a[173]), .B(\ADD_/c[173] ), .Z(
        \ADD_/FAINST[173].FA_/n1 ) );
  XOR \ADD_/FAINST[172].FA_/U5  ( .A(\ADD_/FAINST[172].FA_/n3 ), .B(
        \ADD_/c[172] ), .Z(\ADD_/c[173] ) );
  XOR \ADD_/FAINST[172].FA_/U4  ( .A(\ADD_/FAINST[172].FA_/n1 ), .B(b[172]), 
        .Z(c[172]) );
  AND \ADD_/FAINST[172].FA_/U3  ( .A(\ADD_/FAINST[172].FA_/n1 ), .B(
        \ADD_/FAINST[172].FA_/n2 ), .Z(\ADD_/FAINST[172].FA_/n3 ) );
  XOR \ADD_/FAINST[172].FA_/U2  ( .A(b[172]), .B(\ADD_/c[172] ), .Z(
        \ADD_/FAINST[172].FA_/n2 ) );
  XOR \ADD_/FAINST[172].FA_/U1  ( .A(a[172]), .B(\ADD_/c[172] ), .Z(
        \ADD_/FAINST[172].FA_/n1 ) );
  XOR \ADD_/FAINST[171].FA_/U5  ( .A(\ADD_/FAINST[171].FA_/n3 ), .B(
        \ADD_/c[171] ), .Z(\ADD_/c[172] ) );
  XOR \ADD_/FAINST[171].FA_/U4  ( .A(\ADD_/FAINST[171].FA_/n1 ), .B(b[171]), 
        .Z(c[171]) );
  AND \ADD_/FAINST[171].FA_/U3  ( .A(\ADD_/FAINST[171].FA_/n1 ), .B(
        \ADD_/FAINST[171].FA_/n2 ), .Z(\ADD_/FAINST[171].FA_/n3 ) );
  XOR \ADD_/FAINST[171].FA_/U2  ( .A(b[171]), .B(\ADD_/c[171] ), .Z(
        \ADD_/FAINST[171].FA_/n2 ) );
  XOR \ADD_/FAINST[171].FA_/U1  ( .A(a[171]), .B(\ADD_/c[171] ), .Z(
        \ADD_/FAINST[171].FA_/n1 ) );
  XOR \ADD_/FAINST[170].FA_/U5  ( .A(\ADD_/FAINST[170].FA_/n3 ), .B(
        \ADD_/c[170] ), .Z(\ADD_/c[171] ) );
  XOR \ADD_/FAINST[170].FA_/U4  ( .A(\ADD_/FAINST[170].FA_/n1 ), .B(b[170]), 
        .Z(c[170]) );
  AND \ADD_/FAINST[170].FA_/U3  ( .A(\ADD_/FAINST[170].FA_/n1 ), .B(
        \ADD_/FAINST[170].FA_/n2 ), .Z(\ADD_/FAINST[170].FA_/n3 ) );
  XOR \ADD_/FAINST[170].FA_/U2  ( .A(b[170]), .B(\ADD_/c[170] ), .Z(
        \ADD_/FAINST[170].FA_/n2 ) );
  XOR \ADD_/FAINST[170].FA_/U1  ( .A(a[170]), .B(\ADD_/c[170] ), .Z(
        \ADD_/FAINST[170].FA_/n1 ) );
  XOR \ADD_/FAINST[169].FA_/U5  ( .A(\ADD_/FAINST[169].FA_/n3 ), .B(
        \ADD_/c[169] ), .Z(\ADD_/c[170] ) );
  XOR \ADD_/FAINST[169].FA_/U4  ( .A(\ADD_/FAINST[169].FA_/n1 ), .B(b[169]), 
        .Z(c[169]) );
  AND \ADD_/FAINST[169].FA_/U3  ( .A(\ADD_/FAINST[169].FA_/n1 ), .B(
        \ADD_/FAINST[169].FA_/n2 ), .Z(\ADD_/FAINST[169].FA_/n3 ) );
  XOR \ADD_/FAINST[169].FA_/U2  ( .A(b[169]), .B(\ADD_/c[169] ), .Z(
        \ADD_/FAINST[169].FA_/n2 ) );
  XOR \ADD_/FAINST[169].FA_/U1  ( .A(a[169]), .B(\ADD_/c[169] ), .Z(
        \ADD_/FAINST[169].FA_/n1 ) );
  XOR \ADD_/FAINST[168].FA_/U5  ( .A(\ADD_/FAINST[168].FA_/n3 ), .B(
        \ADD_/c[168] ), .Z(\ADD_/c[169] ) );
  XOR \ADD_/FAINST[168].FA_/U4  ( .A(\ADD_/FAINST[168].FA_/n1 ), .B(b[168]), 
        .Z(c[168]) );
  AND \ADD_/FAINST[168].FA_/U3  ( .A(\ADD_/FAINST[168].FA_/n1 ), .B(
        \ADD_/FAINST[168].FA_/n2 ), .Z(\ADD_/FAINST[168].FA_/n3 ) );
  XOR \ADD_/FAINST[168].FA_/U2  ( .A(b[168]), .B(\ADD_/c[168] ), .Z(
        \ADD_/FAINST[168].FA_/n2 ) );
  XOR \ADD_/FAINST[168].FA_/U1  ( .A(a[168]), .B(\ADD_/c[168] ), .Z(
        \ADD_/FAINST[168].FA_/n1 ) );
  XOR \ADD_/FAINST[167].FA_/U5  ( .A(\ADD_/FAINST[167].FA_/n3 ), .B(
        \ADD_/c[167] ), .Z(\ADD_/c[168] ) );
  XOR \ADD_/FAINST[167].FA_/U4  ( .A(\ADD_/FAINST[167].FA_/n1 ), .B(b[167]), 
        .Z(c[167]) );
  AND \ADD_/FAINST[167].FA_/U3  ( .A(\ADD_/FAINST[167].FA_/n1 ), .B(
        \ADD_/FAINST[167].FA_/n2 ), .Z(\ADD_/FAINST[167].FA_/n3 ) );
  XOR \ADD_/FAINST[167].FA_/U2  ( .A(b[167]), .B(\ADD_/c[167] ), .Z(
        \ADD_/FAINST[167].FA_/n2 ) );
  XOR \ADD_/FAINST[167].FA_/U1  ( .A(a[167]), .B(\ADD_/c[167] ), .Z(
        \ADD_/FAINST[167].FA_/n1 ) );
  XOR \ADD_/FAINST[166].FA_/U5  ( .A(\ADD_/FAINST[166].FA_/n3 ), .B(
        \ADD_/c[166] ), .Z(\ADD_/c[167] ) );
  XOR \ADD_/FAINST[166].FA_/U4  ( .A(\ADD_/FAINST[166].FA_/n1 ), .B(b[166]), 
        .Z(c[166]) );
  AND \ADD_/FAINST[166].FA_/U3  ( .A(\ADD_/FAINST[166].FA_/n1 ), .B(
        \ADD_/FAINST[166].FA_/n2 ), .Z(\ADD_/FAINST[166].FA_/n3 ) );
  XOR \ADD_/FAINST[166].FA_/U2  ( .A(b[166]), .B(\ADD_/c[166] ), .Z(
        \ADD_/FAINST[166].FA_/n2 ) );
  XOR \ADD_/FAINST[166].FA_/U1  ( .A(a[166]), .B(\ADD_/c[166] ), .Z(
        \ADD_/FAINST[166].FA_/n1 ) );
  XOR \ADD_/FAINST[165].FA_/U5  ( .A(\ADD_/FAINST[165].FA_/n3 ), .B(
        \ADD_/c[165] ), .Z(\ADD_/c[166] ) );
  XOR \ADD_/FAINST[165].FA_/U4  ( .A(\ADD_/FAINST[165].FA_/n1 ), .B(b[165]), 
        .Z(c[165]) );
  AND \ADD_/FAINST[165].FA_/U3  ( .A(\ADD_/FAINST[165].FA_/n1 ), .B(
        \ADD_/FAINST[165].FA_/n2 ), .Z(\ADD_/FAINST[165].FA_/n3 ) );
  XOR \ADD_/FAINST[165].FA_/U2  ( .A(b[165]), .B(\ADD_/c[165] ), .Z(
        \ADD_/FAINST[165].FA_/n2 ) );
  XOR \ADD_/FAINST[165].FA_/U1  ( .A(a[165]), .B(\ADD_/c[165] ), .Z(
        \ADD_/FAINST[165].FA_/n1 ) );
  XOR \ADD_/FAINST[164].FA_/U5  ( .A(\ADD_/FAINST[164].FA_/n3 ), .B(
        \ADD_/c[164] ), .Z(\ADD_/c[165] ) );
  XOR \ADD_/FAINST[164].FA_/U4  ( .A(\ADD_/FAINST[164].FA_/n1 ), .B(b[164]), 
        .Z(c[164]) );
  AND \ADD_/FAINST[164].FA_/U3  ( .A(\ADD_/FAINST[164].FA_/n1 ), .B(
        \ADD_/FAINST[164].FA_/n2 ), .Z(\ADD_/FAINST[164].FA_/n3 ) );
  XOR \ADD_/FAINST[164].FA_/U2  ( .A(b[164]), .B(\ADD_/c[164] ), .Z(
        \ADD_/FAINST[164].FA_/n2 ) );
  XOR \ADD_/FAINST[164].FA_/U1  ( .A(a[164]), .B(\ADD_/c[164] ), .Z(
        \ADD_/FAINST[164].FA_/n1 ) );
  XOR \ADD_/FAINST[163].FA_/U5  ( .A(\ADD_/FAINST[163].FA_/n3 ), .B(
        \ADD_/c[163] ), .Z(\ADD_/c[164] ) );
  XOR \ADD_/FAINST[163].FA_/U4  ( .A(\ADD_/FAINST[163].FA_/n1 ), .B(b[163]), 
        .Z(c[163]) );
  AND \ADD_/FAINST[163].FA_/U3  ( .A(\ADD_/FAINST[163].FA_/n1 ), .B(
        \ADD_/FAINST[163].FA_/n2 ), .Z(\ADD_/FAINST[163].FA_/n3 ) );
  XOR \ADD_/FAINST[163].FA_/U2  ( .A(b[163]), .B(\ADD_/c[163] ), .Z(
        \ADD_/FAINST[163].FA_/n2 ) );
  XOR \ADD_/FAINST[163].FA_/U1  ( .A(a[163]), .B(\ADD_/c[163] ), .Z(
        \ADD_/FAINST[163].FA_/n1 ) );
  XOR \ADD_/FAINST[162].FA_/U5  ( .A(\ADD_/FAINST[162].FA_/n3 ), .B(
        \ADD_/c[162] ), .Z(\ADD_/c[163] ) );
  XOR \ADD_/FAINST[162].FA_/U4  ( .A(\ADD_/FAINST[162].FA_/n1 ), .B(b[162]), 
        .Z(c[162]) );
  AND \ADD_/FAINST[162].FA_/U3  ( .A(\ADD_/FAINST[162].FA_/n1 ), .B(
        \ADD_/FAINST[162].FA_/n2 ), .Z(\ADD_/FAINST[162].FA_/n3 ) );
  XOR \ADD_/FAINST[162].FA_/U2  ( .A(b[162]), .B(\ADD_/c[162] ), .Z(
        \ADD_/FAINST[162].FA_/n2 ) );
  XOR \ADD_/FAINST[162].FA_/U1  ( .A(a[162]), .B(\ADD_/c[162] ), .Z(
        \ADD_/FAINST[162].FA_/n1 ) );
  XOR \ADD_/FAINST[161].FA_/U5  ( .A(\ADD_/FAINST[161].FA_/n3 ), .B(
        \ADD_/c[161] ), .Z(\ADD_/c[162] ) );
  XOR \ADD_/FAINST[161].FA_/U4  ( .A(\ADD_/FAINST[161].FA_/n1 ), .B(b[161]), 
        .Z(c[161]) );
  AND \ADD_/FAINST[161].FA_/U3  ( .A(\ADD_/FAINST[161].FA_/n1 ), .B(
        \ADD_/FAINST[161].FA_/n2 ), .Z(\ADD_/FAINST[161].FA_/n3 ) );
  XOR \ADD_/FAINST[161].FA_/U2  ( .A(b[161]), .B(\ADD_/c[161] ), .Z(
        \ADD_/FAINST[161].FA_/n2 ) );
  XOR \ADD_/FAINST[161].FA_/U1  ( .A(a[161]), .B(\ADD_/c[161] ), .Z(
        \ADD_/FAINST[161].FA_/n1 ) );
  XOR \ADD_/FAINST[160].FA_/U5  ( .A(\ADD_/FAINST[160].FA_/n3 ), .B(
        \ADD_/c[160] ), .Z(\ADD_/c[161] ) );
  XOR \ADD_/FAINST[160].FA_/U4  ( .A(\ADD_/FAINST[160].FA_/n1 ), .B(b[160]), 
        .Z(c[160]) );
  AND \ADD_/FAINST[160].FA_/U3  ( .A(\ADD_/FAINST[160].FA_/n1 ), .B(
        \ADD_/FAINST[160].FA_/n2 ), .Z(\ADD_/FAINST[160].FA_/n3 ) );
  XOR \ADD_/FAINST[160].FA_/U2  ( .A(b[160]), .B(\ADD_/c[160] ), .Z(
        \ADD_/FAINST[160].FA_/n2 ) );
  XOR \ADD_/FAINST[160].FA_/U1  ( .A(a[160]), .B(\ADD_/c[160] ), .Z(
        \ADD_/FAINST[160].FA_/n1 ) );
  XOR \ADD_/FAINST[159].FA_/U5  ( .A(\ADD_/FAINST[159].FA_/n3 ), .B(
        \ADD_/c[159] ), .Z(\ADD_/c[160] ) );
  XOR \ADD_/FAINST[159].FA_/U4  ( .A(\ADD_/FAINST[159].FA_/n1 ), .B(b[159]), 
        .Z(c[159]) );
  AND \ADD_/FAINST[159].FA_/U3  ( .A(\ADD_/FAINST[159].FA_/n1 ), .B(
        \ADD_/FAINST[159].FA_/n2 ), .Z(\ADD_/FAINST[159].FA_/n3 ) );
  XOR \ADD_/FAINST[159].FA_/U2  ( .A(b[159]), .B(\ADD_/c[159] ), .Z(
        \ADD_/FAINST[159].FA_/n2 ) );
  XOR \ADD_/FAINST[159].FA_/U1  ( .A(a[159]), .B(\ADD_/c[159] ), .Z(
        \ADD_/FAINST[159].FA_/n1 ) );
  XOR \ADD_/FAINST[158].FA_/U5  ( .A(\ADD_/FAINST[158].FA_/n3 ), .B(
        \ADD_/c[158] ), .Z(\ADD_/c[159] ) );
  XOR \ADD_/FAINST[158].FA_/U4  ( .A(\ADD_/FAINST[158].FA_/n1 ), .B(b[158]), 
        .Z(c[158]) );
  AND \ADD_/FAINST[158].FA_/U3  ( .A(\ADD_/FAINST[158].FA_/n1 ), .B(
        \ADD_/FAINST[158].FA_/n2 ), .Z(\ADD_/FAINST[158].FA_/n3 ) );
  XOR \ADD_/FAINST[158].FA_/U2  ( .A(b[158]), .B(\ADD_/c[158] ), .Z(
        \ADD_/FAINST[158].FA_/n2 ) );
  XOR \ADD_/FAINST[158].FA_/U1  ( .A(a[158]), .B(\ADD_/c[158] ), .Z(
        \ADD_/FAINST[158].FA_/n1 ) );
  XOR \ADD_/FAINST[157].FA_/U5  ( .A(\ADD_/FAINST[157].FA_/n3 ), .B(
        \ADD_/c[157] ), .Z(\ADD_/c[158] ) );
  XOR \ADD_/FAINST[157].FA_/U4  ( .A(\ADD_/FAINST[157].FA_/n1 ), .B(b[157]), 
        .Z(c[157]) );
  AND \ADD_/FAINST[157].FA_/U3  ( .A(\ADD_/FAINST[157].FA_/n1 ), .B(
        \ADD_/FAINST[157].FA_/n2 ), .Z(\ADD_/FAINST[157].FA_/n3 ) );
  XOR \ADD_/FAINST[157].FA_/U2  ( .A(b[157]), .B(\ADD_/c[157] ), .Z(
        \ADD_/FAINST[157].FA_/n2 ) );
  XOR \ADD_/FAINST[157].FA_/U1  ( .A(a[157]), .B(\ADD_/c[157] ), .Z(
        \ADD_/FAINST[157].FA_/n1 ) );
  XOR \ADD_/FAINST[156].FA_/U5  ( .A(\ADD_/FAINST[156].FA_/n3 ), .B(
        \ADD_/c[156] ), .Z(\ADD_/c[157] ) );
  XOR \ADD_/FAINST[156].FA_/U4  ( .A(\ADD_/FAINST[156].FA_/n1 ), .B(b[156]), 
        .Z(c[156]) );
  AND \ADD_/FAINST[156].FA_/U3  ( .A(\ADD_/FAINST[156].FA_/n1 ), .B(
        \ADD_/FAINST[156].FA_/n2 ), .Z(\ADD_/FAINST[156].FA_/n3 ) );
  XOR \ADD_/FAINST[156].FA_/U2  ( .A(b[156]), .B(\ADD_/c[156] ), .Z(
        \ADD_/FAINST[156].FA_/n2 ) );
  XOR \ADD_/FAINST[156].FA_/U1  ( .A(a[156]), .B(\ADD_/c[156] ), .Z(
        \ADD_/FAINST[156].FA_/n1 ) );
  XOR \ADD_/FAINST[155].FA_/U5  ( .A(\ADD_/FAINST[155].FA_/n3 ), .B(
        \ADD_/c[155] ), .Z(\ADD_/c[156] ) );
  XOR \ADD_/FAINST[155].FA_/U4  ( .A(\ADD_/FAINST[155].FA_/n1 ), .B(b[155]), 
        .Z(c[155]) );
  AND \ADD_/FAINST[155].FA_/U3  ( .A(\ADD_/FAINST[155].FA_/n1 ), .B(
        \ADD_/FAINST[155].FA_/n2 ), .Z(\ADD_/FAINST[155].FA_/n3 ) );
  XOR \ADD_/FAINST[155].FA_/U2  ( .A(b[155]), .B(\ADD_/c[155] ), .Z(
        \ADD_/FAINST[155].FA_/n2 ) );
  XOR \ADD_/FAINST[155].FA_/U1  ( .A(a[155]), .B(\ADD_/c[155] ), .Z(
        \ADD_/FAINST[155].FA_/n1 ) );
  XOR \ADD_/FAINST[154].FA_/U5  ( .A(\ADD_/FAINST[154].FA_/n3 ), .B(
        \ADD_/c[154] ), .Z(\ADD_/c[155] ) );
  XOR \ADD_/FAINST[154].FA_/U4  ( .A(\ADD_/FAINST[154].FA_/n1 ), .B(b[154]), 
        .Z(c[154]) );
  AND \ADD_/FAINST[154].FA_/U3  ( .A(\ADD_/FAINST[154].FA_/n1 ), .B(
        \ADD_/FAINST[154].FA_/n2 ), .Z(\ADD_/FAINST[154].FA_/n3 ) );
  XOR \ADD_/FAINST[154].FA_/U2  ( .A(b[154]), .B(\ADD_/c[154] ), .Z(
        \ADD_/FAINST[154].FA_/n2 ) );
  XOR \ADD_/FAINST[154].FA_/U1  ( .A(a[154]), .B(\ADD_/c[154] ), .Z(
        \ADD_/FAINST[154].FA_/n1 ) );
  XOR \ADD_/FAINST[153].FA_/U5  ( .A(\ADD_/FAINST[153].FA_/n3 ), .B(
        \ADD_/c[153] ), .Z(\ADD_/c[154] ) );
  XOR \ADD_/FAINST[153].FA_/U4  ( .A(\ADD_/FAINST[153].FA_/n1 ), .B(b[153]), 
        .Z(c[153]) );
  AND \ADD_/FAINST[153].FA_/U3  ( .A(\ADD_/FAINST[153].FA_/n1 ), .B(
        \ADD_/FAINST[153].FA_/n2 ), .Z(\ADD_/FAINST[153].FA_/n3 ) );
  XOR \ADD_/FAINST[153].FA_/U2  ( .A(b[153]), .B(\ADD_/c[153] ), .Z(
        \ADD_/FAINST[153].FA_/n2 ) );
  XOR \ADD_/FAINST[153].FA_/U1  ( .A(a[153]), .B(\ADD_/c[153] ), .Z(
        \ADD_/FAINST[153].FA_/n1 ) );
  XOR \ADD_/FAINST[152].FA_/U5  ( .A(\ADD_/FAINST[152].FA_/n3 ), .B(
        \ADD_/c[152] ), .Z(\ADD_/c[153] ) );
  XOR \ADD_/FAINST[152].FA_/U4  ( .A(\ADD_/FAINST[152].FA_/n1 ), .B(b[152]), 
        .Z(c[152]) );
  AND \ADD_/FAINST[152].FA_/U3  ( .A(\ADD_/FAINST[152].FA_/n1 ), .B(
        \ADD_/FAINST[152].FA_/n2 ), .Z(\ADD_/FAINST[152].FA_/n3 ) );
  XOR \ADD_/FAINST[152].FA_/U2  ( .A(b[152]), .B(\ADD_/c[152] ), .Z(
        \ADD_/FAINST[152].FA_/n2 ) );
  XOR \ADD_/FAINST[152].FA_/U1  ( .A(a[152]), .B(\ADD_/c[152] ), .Z(
        \ADD_/FAINST[152].FA_/n1 ) );
  XOR \ADD_/FAINST[151].FA_/U5  ( .A(\ADD_/FAINST[151].FA_/n3 ), .B(
        \ADD_/c[151] ), .Z(\ADD_/c[152] ) );
  XOR \ADD_/FAINST[151].FA_/U4  ( .A(\ADD_/FAINST[151].FA_/n1 ), .B(b[151]), 
        .Z(c[151]) );
  AND \ADD_/FAINST[151].FA_/U3  ( .A(\ADD_/FAINST[151].FA_/n1 ), .B(
        \ADD_/FAINST[151].FA_/n2 ), .Z(\ADD_/FAINST[151].FA_/n3 ) );
  XOR \ADD_/FAINST[151].FA_/U2  ( .A(b[151]), .B(\ADD_/c[151] ), .Z(
        \ADD_/FAINST[151].FA_/n2 ) );
  XOR \ADD_/FAINST[151].FA_/U1  ( .A(a[151]), .B(\ADD_/c[151] ), .Z(
        \ADD_/FAINST[151].FA_/n1 ) );
  XOR \ADD_/FAINST[150].FA_/U5  ( .A(\ADD_/FAINST[150].FA_/n3 ), .B(
        \ADD_/c[150] ), .Z(\ADD_/c[151] ) );
  XOR \ADD_/FAINST[150].FA_/U4  ( .A(\ADD_/FAINST[150].FA_/n1 ), .B(b[150]), 
        .Z(c[150]) );
  AND \ADD_/FAINST[150].FA_/U3  ( .A(\ADD_/FAINST[150].FA_/n1 ), .B(
        \ADD_/FAINST[150].FA_/n2 ), .Z(\ADD_/FAINST[150].FA_/n3 ) );
  XOR \ADD_/FAINST[150].FA_/U2  ( .A(b[150]), .B(\ADD_/c[150] ), .Z(
        \ADD_/FAINST[150].FA_/n2 ) );
  XOR \ADD_/FAINST[150].FA_/U1  ( .A(a[150]), .B(\ADD_/c[150] ), .Z(
        \ADD_/FAINST[150].FA_/n1 ) );
  XOR \ADD_/FAINST[149].FA_/U5  ( .A(\ADD_/FAINST[149].FA_/n3 ), .B(
        \ADD_/c[149] ), .Z(\ADD_/c[150] ) );
  XOR \ADD_/FAINST[149].FA_/U4  ( .A(\ADD_/FAINST[149].FA_/n1 ), .B(b[149]), 
        .Z(c[149]) );
  AND \ADD_/FAINST[149].FA_/U3  ( .A(\ADD_/FAINST[149].FA_/n1 ), .B(
        \ADD_/FAINST[149].FA_/n2 ), .Z(\ADD_/FAINST[149].FA_/n3 ) );
  XOR \ADD_/FAINST[149].FA_/U2  ( .A(b[149]), .B(\ADD_/c[149] ), .Z(
        \ADD_/FAINST[149].FA_/n2 ) );
  XOR \ADD_/FAINST[149].FA_/U1  ( .A(a[149]), .B(\ADD_/c[149] ), .Z(
        \ADD_/FAINST[149].FA_/n1 ) );
  XOR \ADD_/FAINST[148].FA_/U5  ( .A(\ADD_/FAINST[148].FA_/n3 ), .B(
        \ADD_/c[148] ), .Z(\ADD_/c[149] ) );
  XOR \ADD_/FAINST[148].FA_/U4  ( .A(\ADD_/FAINST[148].FA_/n1 ), .B(b[148]), 
        .Z(c[148]) );
  AND \ADD_/FAINST[148].FA_/U3  ( .A(\ADD_/FAINST[148].FA_/n1 ), .B(
        \ADD_/FAINST[148].FA_/n2 ), .Z(\ADD_/FAINST[148].FA_/n3 ) );
  XOR \ADD_/FAINST[148].FA_/U2  ( .A(b[148]), .B(\ADD_/c[148] ), .Z(
        \ADD_/FAINST[148].FA_/n2 ) );
  XOR \ADD_/FAINST[148].FA_/U1  ( .A(a[148]), .B(\ADD_/c[148] ), .Z(
        \ADD_/FAINST[148].FA_/n1 ) );
  XOR \ADD_/FAINST[147].FA_/U5  ( .A(\ADD_/FAINST[147].FA_/n3 ), .B(
        \ADD_/c[147] ), .Z(\ADD_/c[148] ) );
  XOR \ADD_/FAINST[147].FA_/U4  ( .A(\ADD_/FAINST[147].FA_/n1 ), .B(b[147]), 
        .Z(c[147]) );
  AND \ADD_/FAINST[147].FA_/U3  ( .A(\ADD_/FAINST[147].FA_/n1 ), .B(
        \ADD_/FAINST[147].FA_/n2 ), .Z(\ADD_/FAINST[147].FA_/n3 ) );
  XOR \ADD_/FAINST[147].FA_/U2  ( .A(b[147]), .B(\ADD_/c[147] ), .Z(
        \ADD_/FAINST[147].FA_/n2 ) );
  XOR \ADD_/FAINST[147].FA_/U1  ( .A(a[147]), .B(\ADD_/c[147] ), .Z(
        \ADD_/FAINST[147].FA_/n1 ) );
  XOR \ADD_/FAINST[146].FA_/U5  ( .A(\ADD_/FAINST[146].FA_/n3 ), .B(
        \ADD_/c[146] ), .Z(\ADD_/c[147] ) );
  XOR \ADD_/FAINST[146].FA_/U4  ( .A(\ADD_/FAINST[146].FA_/n1 ), .B(b[146]), 
        .Z(c[146]) );
  AND \ADD_/FAINST[146].FA_/U3  ( .A(\ADD_/FAINST[146].FA_/n1 ), .B(
        \ADD_/FAINST[146].FA_/n2 ), .Z(\ADD_/FAINST[146].FA_/n3 ) );
  XOR \ADD_/FAINST[146].FA_/U2  ( .A(b[146]), .B(\ADD_/c[146] ), .Z(
        \ADD_/FAINST[146].FA_/n2 ) );
  XOR \ADD_/FAINST[146].FA_/U1  ( .A(a[146]), .B(\ADD_/c[146] ), .Z(
        \ADD_/FAINST[146].FA_/n1 ) );
  XOR \ADD_/FAINST[145].FA_/U5  ( .A(\ADD_/FAINST[145].FA_/n3 ), .B(
        \ADD_/c[145] ), .Z(\ADD_/c[146] ) );
  XOR \ADD_/FAINST[145].FA_/U4  ( .A(\ADD_/FAINST[145].FA_/n1 ), .B(b[145]), 
        .Z(c[145]) );
  AND \ADD_/FAINST[145].FA_/U3  ( .A(\ADD_/FAINST[145].FA_/n1 ), .B(
        \ADD_/FAINST[145].FA_/n2 ), .Z(\ADD_/FAINST[145].FA_/n3 ) );
  XOR \ADD_/FAINST[145].FA_/U2  ( .A(b[145]), .B(\ADD_/c[145] ), .Z(
        \ADD_/FAINST[145].FA_/n2 ) );
  XOR \ADD_/FAINST[145].FA_/U1  ( .A(a[145]), .B(\ADD_/c[145] ), .Z(
        \ADD_/FAINST[145].FA_/n1 ) );
  XOR \ADD_/FAINST[144].FA_/U5  ( .A(\ADD_/FAINST[144].FA_/n3 ), .B(
        \ADD_/c[144] ), .Z(\ADD_/c[145] ) );
  XOR \ADD_/FAINST[144].FA_/U4  ( .A(\ADD_/FAINST[144].FA_/n1 ), .B(b[144]), 
        .Z(c[144]) );
  AND \ADD_/FAINST[144].FA_/U3  ( .A(\ADD_/FAINST[144].FA_/n1 ), .B(
        \ADD_/FAINST[144].FA_/n2 ), .Z(\ADD_/FAINST[144].FA_/n3 ) );
  XOR \ADD_/FAINST[144].FA_/U2  ( .A(b[144]), .B(\ADD_/c[144] ), .Z(
        \ADD_/FAINST[144].FA_/n2 ) );
  XOR \ADD_/FAINST[144].FA_/U1  ( .A(a[144]), .B(\ADD_/c[144] ), .Z(
        \ADD_/FAINST[144].FA_/n1 ) );
  XOR \ADD_/FAINST[143].FA_/U5  ( .A(\ADD_/FAINST[143].FA_/n3 ), .B(
        \ADD_/c[143] ), .Z(\ADD_/c[144] ) );
  XOR \ADD_/FAINST[143].FA_/U4  ( .A(\ADD_/FAINST[143].FA_/n1 ), .B(b[143]), 
        .Z(c[143]) );
  AND \ADD_/FAINST[143].FA_/U3  ( .A(\ADD_/FAINST[143].FA_/n1 ), .B(
        \ADD_/FAINST[143].FA_/n2 ), .Z(\ADD_/FAINST[143].FA_/n3 ) );
  XOR \ADD_/FAINST[143].FA_/U2  ( .A(b[143]), .B(\ADD_/c[143] ), .Z(
        \ADD_/FAINST[143].FA_/n2 ) );
  XOR \ADD_/FAINST[143].FA_/U1  ( .A(a[143]), .B(\ADD_/c[143] ), .Z(
        \ADD_/FAINST[143].FA_/n1 ) );
  XOR \ADD_/FAINST[142].FA_/U5  ( .A(\ADD_/FAINST[142].FA_/n3 ), .B(
        \ADD_/c[142] ), .Z(\ADD_/c[143] ) );
  XOR \ADD_/FAINST[142].FA_/U4  ( .A(\ADD_/FAINST[142].FA_/n1 ), .B(b[142]), 
        .Z(c[142]) );
  AND \ADD_/FAINST[142].FA_/U3  ( .A(\ADD_/FAINST[142].FA_/n1 ), .B(
        \ADD_/FAINST[142].FA_/n2 ), .Z(\ADD_/FAINST[142].FA_/n3 ) );
  XOR \ADD_/FAINST[142].FA_/U2  ( .A(b[142]), .B(\ADD_/c[142] ), .Z(
        \ADD_/FAINST[142].FA_/n2 ) );
  XOR \ADD_/FAINST[142].FA_/U1  ( .A(a[142]), .B(\ADD_/c[142] ), .Z(
        \ADD_/FAINST[142].FA_/n1 ) );
  XOR \ADD_/FAINST[141].FA_/U5  ( .A(\ADD_/FAINST[141].FA_/n3 ), .B(
        \ADD_/c[141] ), .Z(\ADD_/c[142] ) );
  XOR \ADD_/FAINST[141].FA_/U4  ( .A(\ADD_/FAINST[141].FA_/n1 ), .B(b[141]), 
        .Z(c[141]) );
  AND \ADD_/FAINST[141].FA_/U3  ( .A(\ADD_/FAINST[141].FA_/n1 ), .B(
        \ADD_/FAINST[141].FA_/n2 ), .Z(\ADD_/FAINST[141].FA_/n3 ) );
  XOR \ADD_/FAINST[141].FA_/U2  ( .A(b[141]), .B(\ADD_/c[141] ), .Z(
        \ADD_/FAINST[141].FA_/n2 ) );
  XOR \ADD_/FAINST[141].FA_/U1  ( .A(a[141]), .B(\ADD_/c[141] ), .Z(
        \ADD_/FAINST[141].FA_/n1 ) );
  XOR \ADD_/FAINST[140].FA_/U5  ( .A(\ADD_/FAINST[140].FA_/n3 ), .B(
        \ADD_/c[140] ), .Z(\ADD_/c[141] ) );
  XOR \ADD_/FAINST[140].FA_/U4  ( .A(\ADD_/FAINST[140].FA_/n1 ), .B(b[140]), 
        .Z(c[140]) );
  AND \ADD_/FAINST[140].FA_/U3  ( .A(\ADD_/FAINST[140].FA_/n1 ), .B(
        \ADD_/FAINST[140].FA_/n2 ), .Z(\ADD_/FAINST[140].FA_/n3 ) );
  XOR \ADD_/FAINST[140].FA_/U2  ( .A(b[140]), .B(\ADD_/c[140] ), .Z(
        \ADD_/FAINST[140].FA_/n2 ) );
  XOR \ADD_/FAINST[140].FA_/U1  ( .A(a[140]), .B(\ADD_/c[140] ), .Z(
        \ADD_/FAINST[140].FA_/n1 ) );
  XOR \ADD_/FAINST[139].FA_/U5  ( .A(\ADD_/FAINST[139].FA_/n3 ), .B(
        \ADD_/c[139] ), .Z(\ADD_/c[140] ) );
  XOR \ADD_/FAINST[139].FA_/U4  ( .A(\ADD_/FAINST[139].FA_/n1 ), .B(b[139]), 
        .Z(c[139]) );
  AND \ADD_/FAINST[139].FA_/U3  ( .A(\ADD_/FAINST[139].FA_/n1 ), .B(
        \ADD_/FAINST[139].FA_/n2 ), .Z(\ADD_/FAINST[139].FA_/n3 ) );
  XOR \ADD_/FAINST[139].FA_/U2  ( .A(b[139]), .B(\ADD_/c[139] ), .Z(
        \ADD_/FAINST[139].FA_/n2 ) );
  XOR \ADD_/FAINST[139].FA_/U1  ( .A(a[139]), .B(\ADD_/c[139] ), .Z(
        \ADD_/FAINST[139].FA_/n1 ) );
  XOR \ADD_/FAINST[138].FA_/U5  ( .A(\ADD_/FAINST[138].FA_/n3 ), .B(
        \ADD_/c[138] ), .Z(\ADD_/c[139] ) );
  XOR \ADD_/FAINST[138].FA_/U4  ( .A(\ADD_/FAINST[138].FA_/n1 ), .B(b[138]), 
        .Z(c[138]) );
  AND \ADD_/FAINST[138].FA_/U3  ( .A(\ADD_/FAINST[138].FA_/n1 ), .B(
        \ADD_/FAINST[138].FA_/n2 ), .Z(\ADD_/FAINST[138].FA_/n3 ) );
  XOR \ADD_/FAINST[138].FA_/U2  ( .A(b[138]), .B(\ADD_/c[138] ), .Z(
        \ADD_/FAINST[138].FA_/n2 ) );
  XOR \ADD_/FAINST[138].FA_/U1  ( .A(a[138]), .B(\ADD_/c[138] ), .Z(
        \ADD_/FAINST[138].FA_/n1 ) );
  XOR \ADD_/FAINST[137].FA_/U5  ( .A(\ADD_/FAINST[137].FA_/n3 ), .B(
        \ADD_/c[137] ), .Z(\ADD_/c[138] ) );
  XOR \ADD_/FAINST[137].FA_/U4  ( .A(\ADD_/FAINST[137].FA_/n1 ), .B(b[137]), 
        .Z(c[137]) );
  AND \ADD_/FAINST[137].FA_/U3  ( .A(\ADD_/FAINST[137].FA_/n1 ), .B(
        \ADD_/FAINST[137].FA_/n2 ), .Z(\ADD_/FAINST[137].FA_/n3 ) );
  XOR \ADD_/FAINST[137].FA_/U2  ( .A(b[137]), .B(\ADD_/c[137] ), .Z(
        \ADD_/FAINST[137].FA_/n2 ) );
  XOR \ADD_/FAINST[137].FA_/U1  ( .A(a[137]), .B(\ADD_/c[137] ), .Z(
        \ADD_/FAINST[137].FA_/n1 ) );
  XOR \ADD_/FAINST[136].FA_/U5  ( .A(\ADD_/FAINST[136].FA_/n3 ), .B(
        \ADD_/c[136] ), .Z(\ADD_/c[137] ) );
  XOR \ADD_/FAINST[136].FA_/U4  ( .A(\ADD_/FAINST[136].FA_/n1 ), .B(b[136]), 
        .Z(c[136]) );
  AND \ADD_/FAINST[136].FA_/U3  ( .A(\ADD_/FAINST[136].FA_/n1 ), .B(
        \ADD_/FAINST[136].FA_/n2 ), .Z(\ADD_/FAINST[136].FA_/n3 ) );
  XOR \ADD_/FAINST[136].FA_/U2  ( .A(b[136]), .B(\ADD_/c[136] ), .Z(
        \ADD_/FAINST[136].FA_/n2 ) );
  XOR \ADD_/FAINST[136].FA_/U1  ( .A(a[136]), .B(\ADD_/c[136] ), .Z(
        \ADD_/FAINST[136].FA_/n1 ) );
  XOR \ADD_/FAINST[135].FA_/U5  ( .A(\ADD_/FAINST[135].FA_/n3 ), .B(
        \ADD_/c[135] ), .Z(\ADD_/c[136] ) );
  XOR \ADD_/FAINST[135].FA_/U4  ( .A(\ADD_/FAINST[135].FA_/n1 ), .B(b[135]), 
        .Z(c[135]) );
  AND \ADD_/FAINST[135].FA_/U3  ( .A(\ADD_/FAINST[135].FA_/n1 ), .B(
        \ADD_/FAINST[135].FA_/n2 ), .Z(\ADD_/FAINST[135].FA_/n3 ) );
  XOR \ADD_/FAINST[135].FA_/U2  ( .A(b[135]), .B(\ADD_/c[135] ), .Z(
        \ADD_/FAINST[135].FA_/n2 ) );
  XOR \ADD_/FAINST[135].FA_/U1  ( .A(a[135]), .B(\ADD_/c[135] ), .Z(
        \ADD_/FAINST[135].FA_/n1 ) );
  XOR \ADD_/FAINST[134].FA_/U5  ( .A(\ADD_/FAINST[134].FA_/n3 ), .B(
        \ADD_/c[134] ), .Z(\ADD_/c[135] ) );
  XOR \ADD_/FAINST[134].FA_/U4  ( .A(\ADD_/FAINST[134].FA_/n1 ), .B(b[134]), 
        .Z(c[134]) );
  AND \ADD_/FAINST[134].FA_/U3  ( .A(\ADD_/FAINST[134].FA_/n1 ), .B(
        \ADD_/FAINST[134].FA_/n2 ), .Z(\ADD_/FAINST[134].FA_/n3 ) );
  XOR \ADD_/FAINST[134].FA_/U2  ( .A(b[134]), .B(\ADD_/c[134] ), .Z(
        \ADD_/FAINST[134].FA_/n2 ) );
  XOR \ADD_/FAINST[134].FA_/U1  ( .A(a[134]), .B(\ADD_/c[134] ), .Z(
        \ADD_/FAINST[134].FA_/n1 ) );
  XOR \ADD_/FAINST[133].FA_/U5  ( .A(\ADD_/FAINST[133].FA_/n3 ), .B(
        \ADD_/c[133] ), .Z(\ADD_/c[134] ) );
  XOR \ADD_/FAINST[133].FA_/U4  ( .A(\ADD_/FAINST[133].FA_/n1 ), .B(b[133]), 
        .Z(c[133]) );
  AND \ADD_/FAINST[133].FA_/U3  ( .A(\ADD_/FAINST[133].FA_/n1 ), .B(
        \ADD_/FAINST[133].FA_/n2 ), .Z(\ADD_/FAINST[133].FA_/n3 ) );
  XOR \ADD_/FAINST[133].FA_/U2  ( .A(b[133]), .B(\ADD_/c[133] ), .Z(
        \ADD_/FAINST[133].FA_/n2 ) );
  XOR \ADD_/FAINST[133].FA_/U1  ( .A(a[133]), .B(\ADD_/c[133] ), .Z(
        \ADD_/FAINST[133].FA_/n1 ) );
  XOR \ADD_/FAINST[132].FA_/U5  ( .A(\ADD_/FAINST[132].FA_/n3 ), .B(
        \ADD_/c[132] ), .Z(\ADD_/c[133] ) );
  XOR \ADD_/FAINST[132].FA_/U4  ( .A(\ADD_/FAINST[132].FA_/n1 ), .B(b[132]), 
        .Z(c[132]) );
  AND \ADD_/FAINST[132].FA_/U3  ( .A(\ADD_/FAINST[132].FA_/n1 ), .B(
        \ADD_/FAINST[132].FA_/n2 ), .Z(\ADD_/FAINST[132].FA_/n3 ) );
  XOR \ADD_/FAINST[132].FA_/U2  ( .A(b[132]), .B(\ADD_/c[132] ), .Z(
        \ADD_/FAINST[132].FA_/n2 ) );
  XOR \ADD_/FAINST[132].FA_/U1  ( .A(a[132]), .B(\ADD_/c[132] ), .Z(
        \ADD_/FAINST[132].FA_/n1 ) );
  XOR \ADD_/FAINST[131].FA_/U5  ( .A(\ADD_/FAINST[131].FA_/n3 ), .B(
        \ADD_/c[131] ), .Z(\ADD_/c[132] ) );
  XOR \ADD_/FAINST[131].FA_/U4  ( .A(\ADD_/FAINST[131].FA_/n1 ), .B(b[131]), 
        .Z(c[131]) );
  AND \ADD_/FAINST[131].FA_/U3  ( .A(\ADD_/FAINST[131].FA_/n1 ), .B(
        \ADD_/FAINST[131].FA_/n2 ), .Z(\ADD_/FAINST[131].FA_/n3 ) );
  XOR \ADD_/FAINST[131].FA_/U2  ( .A(b[131]), .B(\ADD_/c[131] ), .Z(
        \ADD_/FAINST[131].FA_/n2 ) );
  XOR \ADD_/FAINST[131].FA_/U1  ( .A(a[131]), .B(\ADD_/c[131] ), .Z(
        \ADD_/FAINST[131].FA_/n1 ) );
  XOR \ADD_/FAINST[130].FA_/U5  ( .A(\ADD_/FAINST[130].FA_/n3 ), .B(
        \ADD_/c[130] ), .Z(\ADD_/c[131] ) );
  XOR \ADD_/FAINST[130].FA_/U4  ( .A(\ADD_/FAINST[130].FA_/n1 ), .B(b[130]), 
        .Z(c[130]) );
  AND \ADD_/FAINST[130].FA_/U3  ( .A(\ADD_/FAINST[130].FA_/n1 ), .B(
        \ADD_/FAINST[130].FA_/n2 ), .Z(\ADD_/FAINST[130].FA_/n3 ) );
  XOR \ADD_/FAINST[130].FA_/U2  ( .A(b[130]), .B(\ADD_/c[130] ), .Z(
        \ADD_/FAINST[130].FA_/n2 ) );
  XOR \ADD_/FAINST[130].FA_/U1  ( .A(a[130]), .B(\ADD_/c[130] ), .Z(
        \ADD_/FAINST[130].FA_/n1 ) );
  XOR \ADD_/FAINST[129].FA_/U5  ( .A(\ADD_/FAINST[129].FA_/n3 ), .B(
        \ADD_/c[129] ), .Z(\ADD_/c[130] ) );
  XOR \ADD_/FAINST[129].FA_/U4  ( .A(\ADD_/FAINST[129].FA_/n1 ), .B(b[129]), 
        .Z(c[129]) );
  AND \ADD_/FAINST[129].FA_/U3  ( .A(\ADD_/FAINST[129].FA_/n1 ), .B(
        \ADD_/FAINST[129].FA_/n2 ), .Z(\ADD_/FAINST[129].FA_/n3 ) );
  XOR \ADD_/FAINST[129].FA_/U2  ( .A(b[129]), .B(\ADD_/c[129] ), .Z(
        \ADD_/FAINST[129].FA_/n2 ) );
  XOR \ADD_/FAINST[129].FA_/U1  ( .A(a[129]), .B(\ADD_/c[129] ), .Z(
        \ADD_/FAINST[129].FA_/n1 ) );
  XOR \ADD_/FAINST[128].FA_/U5  ( .A(\ADD_/FAINST[128].FA_/n3 ), .B(
        \ADD_/c[128] ), .Z(\ADD_/c[129] ) );
  XOR \ADD_/FAINST[128].FA_/U4  ( .A(\ADD_/FAINST[128].FA_/n1 ), .B(b[128]), 
        .Z(c[128]) );
  AND \ADD_/FAINST[128].FA_/U3  ( .A(\ADD_/FAINST[128].FA_/n1 ), .B(
        \ADD_/FAINST[128].FA_/n2 ), .Z(\ADD_/FAINST[128].FA_/n3 ) );
  XOR \ADD_/FAINST[128].FA_/U2  ( .A(b[128]), .B(\ADD_/c[128] ), .Z(
        \ADD_/FAINST[128].FA_/n2 ) );
  XOR \ADD_/FAINST[128].FA_/U1  ( .A(a[128]), .B(\ADD_/c[128] ), .Z(
        \ADD_/FAINST[128].FA_/n1 ) );
  XOR \ADD_/FAINST[127].FA_/U5  ( .A(\ADD_/FAINST[127].FA_/n3 ), .B(
        \ADD_/c[127] ), .Z(\ADD_/c[128] ) );
  XOR \ADD_/FAINST[127].FA_/U4  ( .A(\ADD_/FAINST[127].FA_/n1 ), .B(b[127]), 
        .Z(c[127]) );
  AND \ADD_/FAINST[127].FA_/U3  ( .A(\ADD_/FAINST[127].FA_/n1 ), .B(
        \ADD_/FAINST[127].FA_/n2 ), .Z(\ADD_/FAINST[127].FA_/n3 ) );
  XOR \ADD_/FAINST[127].FA_/U2  ( .A(b[127]), .B(\ADD_/c[127] ), .Z(
        \ADD_/FAINST[127].FA_/n2 ) );
  XOR \ADD_/FAINST[127].FA_/U1  ( .A(a[127]), .B(\ADD_/c[127] ), .Z(
        \ADD_/FAINST[127].FA_/n1 ) );
  XOR \ADD_/FAINST[126].FA_/U5  ( .A(\ADD_/FAINST[126].FA_/n3 ), .B(
        \ADD_/c[126] ), .Z(\ADD_/c[127] ) );
  XOR \ADD_/FAINST[126].FA_/U4  ( .A(\ADD_/FAINST[126].FA_/n1 ), .B(b[126]), 
        .Z(c[126]) );
  AND \ADD_/FAINST[126].FA_/U3  ( .A(\ADD_/FAINST[126].FA_/n1 ), .B(
        \ADD_/FAINST[126].FA_/n2 ), .Z(\ADD_/FAINST[126].FA_/n3 ) );
  XOR \ADD_/FAINST[126].FA_/U2  ( .A(b[126]), .B(\ADD_/c[126] ), .Z(
        \ADD_/FAINST[126].FA_/n2 ) );
  XOR \ADD_/FAINST[126].FA_/U1  ( .A(a[126]), .B(\ADD_/c[126] ), .Z(
        \ADD_/FAINST[126].FA_/n1 ) );
  XOR \ADD_/FAINST[125].FA_/U5  ( .A(\ADD_/FAINST[125].FA_/n3 ), .B(
        \ADD_/c[125] ), .Z(\ADD_/c[126] ) );
  XOR \ADD_/FAINST[125].FA_/U4  ( .A(\ADD_/FAINST[125].FA_/n1 ), .B(b[125]), 
        .Z(c[125]) );
  AND \ADD_/FAINST[125].FA_/U3  ( .A(\ADD_/FAINST[125].FA_/n1 ), .B(
        \ADD_/FAINST[125].FA_/n2 ), .Z(\ADD_/FAINST[125].FA_/n3 ) );
  XOR \ADD_/FAINST[125].FA_/U2  ( .A(b[125]), .B(\ADD_/c[125] ), .Z(
        \ADD_/FAINST[125].FA_/n2 ) );
  XOR \ADD_/FAINST[125].FA_/U1  ( .A(a[125]), .B(\ADD_/c[125] ), .Z(
        \ADD_/FAINST[125].FA_/n1 ) );
  XOR \ADD_/FAINST[124].FA_/U5  ( .A(\ADD_/FAINST[124].FA_/n3 ), .B(
        \ADD_/c[124] ), .Z(\ADD_/c[125] ) );
  XOR \ADD_/FAINST[124].FA_/U4  ( .A(\ADD_/FAINST[124].FA_/n1 ), .B(b[124]), 
        .Z(c[124]) );
  AND \ADD_/FAINST[124].FA_/U3  ( .A(\ADD_/FAINST[124].FA_/n1 ), .B(
        \ADD_/FAINST[124].FA_/n2 ), .Z(\ADD_/FAINST[124].FA_/n3 ) );
  XOR \ADD_/FAINST[124].FA_/U2  ( .A(b[124]), .B(\ADD_/c[124] ), .Z(
        \ADD_/FAINST[124].FA_/n2 ) );
  XOR \ADD_/FAINST[124].FA_/U1  ( .A(a[124]), .B(\ADD_/c[124] ), .Z(
        \ADD_/FAINST[124].FA_/n1 ) );
  XOR \ADD_/FAINST[123].FA_/U5  ( .A(\ADD_/FAINST[123].FA_/n3 ), .B(
        \ADD_/c[123] ), .Z(\ADD_/c[124] ) );
  XOR \ADD_/FAINST[123].FA_/U4  ( .A(\ADD_/FAINST[123].FA_/n1 ), .B(b[123]), 
        .Z(c[123]) );
  AND \ADD_/FAINST[123].FA_/U3  ( .A(\ADD_/FAINST[123].FA_/n1 ), .B(
        \ADD_/FAINST[123].FA_/n2 ), .Z(\ADD_/FAINST[123].FA_/n3 ) );
  XOR \ADD_/FAINST[123].FA_/U2  ( .A(b[123]), .B(\ADD_/c[123] ), .Z(
        \ADD_/FAINST[123].FA_/n2 ) );
  XOR \ADD_/FAINST[123].FA_/U1  ( .A(a[123]), .B(\ADD_/c[123] ), .Z(
        \ADD_/FAINST[123].FA_/n1 ) );
  XOR \ADD_/FAINST[122].FA_/U5  ( .A(\ADD_/FAINST[122].FA_/n3 ), .B(
        \ADD_/c[122] ), .Z(\ADD_/c[123] ) );
  XOR \ADD_/FAINST[122].FA_/U4  ( .A(\ADD_/FAINST[122].FA_/n1 ), .B(b[122]), 
        .Z(c[122]) );
  AND \ADD_/FAINST[122].FA_/U3  ( .A(\ADD_/FAINST[122].FA_/n1 ), .B(
        \ADD_/FAINST[122].FA_/n2 ), .Z(\ADD_/FAINST[122].FA_/n3 ) );
  XOR \ADD_/FAINST[122].FA_/U2  ( .A(b[122]), .B(\ADD_/c[122] ), .Z(
        \ADD_/FAINST[122].FA_/n2 ) );
  XOR \ADD_/FAINST[122].FA_/U1  ( .A(a[122]), .B(\ADD_/c[122] ), .Z(
        \ADD_/FAINST[122].FA_/n1 ) );
  XOR \ADD_/FAINST[121].FA_/U5  ( .A(\ADD_/FAINST[121].FA_/n3 ), .B(
        \ADD_/c[121] ), .Z(\ADD_/c[122] ) );
  XOR \ADD_/FAINST[121].FA_/U4  ( .A(\ADD_/FAINST[121].FA_/n1 ), .B(b[121]), 
        .Z(c[121]) );
  AND \ADD_/FAINST[121].FA_/U3  ( .A(\ADD_/FAINST[121].FA_/n1 ), .B(
        \ADD_/FAINST[121].FA_/n2 ), .Z(\ADD_/FAINST[121].FA_/n3 ) );
  XOR \ADD_/FAINST[121].FA_/U2  ( .A(b[121]), .B(\ADD_/c[121] ), .Z(
        \ADD_/FAINST[121].FA_/n2 ) );
  XOR \ADD_/FAINST[121].FA_/U1  ( .A(a[121]), .B(\ADD_/c[121] ), .Z(
        \ADD_/FAINST[121].FA_/n1 ) );
  XOR \ADD_/FAINST[120].FA_/U5  ( .A(\ADD_/FAINST[120].FA_/n3 ), .B(
        \ADD_/c[120] ), .Z(\ADD_/c[121] ) );
  XOR \ADD_/FAINST[120].FA_/U4  ( .A(\ADD_/FAINST[120].FA_/n1 ), .B(b[120]), 
        .Z(c[120]) );
  AND \ADD_/FAINST[120].FA_/U3  ( .A(\ADD_/FAINST[120].FA_/n1 ), .B(
        \ADD_/FAINST[120].FA_/n2 ), .Z(\ADD_/FAINST[120].FA_/n3 ) );
  XOR \ADD_/FAINST[120].FA_/U2  ( .A(b[120]), .B(\ADD_/c[120] ), .Z(
        \ADD_/FAINST[120].FA_/n2 ) );
  XOR \ADD_/FAINST[120].FA_/U1  ( .A(a[120]), .B(\ADD_/c[120] ), .Z(
        \ADD_/FAINST[120].FA_/n1 ) );
  XOR \ADD_/FAINST[119].FA_/U5  ( .A(\ADD_/FAINST[119].FA_/n3 ), .B(
        \ADD_/c[119] ), .Z(\ADD_/c[120] ) );
  XOR \ADD_/FAINST[119].FA_/U4  ( .A(\ADD_/FAINST[119].FA_/n1 ), .B(b[119]), 
        .Z(c[119]) );
  AND \ADD_/FAINST[119].FA_/U3  ( .A(\ADD_/FAINST[119].FA_/n1 ), .B(
        \ADD_/FAINST[119].FA_/n2 ), .Z(\ADD_/FAINST[119].FA_/n3 ) );
  XOR \ADD_/FAINST[119].FA_/U2  ( .A(b[119]), .B(\ADD_/c[119] ), .Z(
        \ADD_/FAINST[119].FA_/n2 ) );
  XOR \ADD_/FAINST[119].FA_/U1  ( .A(a[119]), .B(\ADD_/c[119] ), .Z(
        \ADD_/FAINST[119].FA_/n1 ) );
  XOR \ADD_/FAINST[118].FA_/U5  ( .A(\ADD_/FAINST[118].FA_/n3 ), .B(
        \ADD_/c[118] ), .Z(\ADD_/c[119] ) );
  XOR \ADD_/FAINST[118].FA_/U4  ( .A(\ADD_/FAINST[118].FA_/n1 ), .B(b[118]), 
        .Z(c[118]) );
  AND \ADD_/FAINST[118].FA_/U3  ( .A(\ADD_/FAINST[118].FA_/n1 ), .B(
        \ADD_/FAINST[118].FA_/n2 ), .Z(\ADD_/FAINST[118].FA_/n3 ) );
  XOR \ADD_/FAINST[118].FA_/U2  ( .A(b[118]), .B(\ADD_/c[118] ), .Z(
        \ADD_/FAINST[118].FA_/n2 ) );
  XOR \ADD_/FAINST[118].FA_/U1  ( .A(a[118]), .B(\ADD_/c[118] ), .Z(
        \ADD_/FAINST[118].FA_/n1 ) );
  XOR \ADD_/FAINST[117].FA_/U5  ( .A(\ADD_/FAINST[117].FA_/n3 ), .B(
        \ADD_/c[117] ), .Z(\ADD_/c[118] ) );
  XOR \ADD_/FAINST[117].FA_/U4  ( .A(\ADD_/FAINST[117].FA_/n1 ), .B(b[117]), 
        .Z(c[117]) );
  AND \ADD_/FAINST[117].FA_/U3  ( .A(\ADD_/FAINST[117].FA_/n1 ), .B(
        \ADD_/FAINST[117].FA_/n2 ), .Z(\ADD_/FAINST[117].FA_/n3 ) );
  XOR \ADD_/FAINST[117].FA_/U2  ( .A(b[117]), .B(\ADD_/c[117] ), .Z(
        \ADD_/FAINST[117].FA_/n2 ) );
  XOR \ADD_/FAINST[117].FA_/U1  ( .A(a[117]), .B(\ADD_/c[117] ), .Z(
        \ADD_/FAINST[117].FA_/n1 ) );
  XOR \ADD_/FAINST[116].FA_/U5  ( .A(\ADD_/FAINST[116].FA_/n3 ), .B(
        \ADD_/c[116] ), .Z(\ADD_/c[117] ) );
  XOR \ADD_/FAINST[116].FA_/U4  ( .A(\ADD_/FAINST[116].FA_/n1 ), .B(b[116]), 
        .Z(c[116]) );
  AND \ADD_/FAINST[116].FA_/U3  ( .A(\ADD_/FAINST[116].FA_/n1 ), .B(
        \ADD_/FAINST[116].FA_/n2 ), .Z(\ADD_/FAINST[116].FA_/n3 ) );
  XOR \ADD_/FAINST[116].FA_/U2  ( .A(b[116]), .B(\ADD_/c[116] ), .Z(
        \ADD_/FAINST[116].FA_/n2 ) );
  XOR \ADD_/FAINST[116].FA_/U1  ( .A(a[116]), .B(\ADD_/c[116] ), .Z(
        \ADD_/FAINST[116].FA_/n1 ) );
  XOR \ADD_/FAINST[115].FA_/U5  ( .A(\ADD_/FAINST[115].FA_/n3 ), .B(
        \ADD_/c[115] ), .Z(\ADD_/c[116] ) );
  XOR \ADD_/FAINST[115].FA_/U4  ( .A(\ADD_/FAINST[115].FA_/n1 ), .B(b[115]), 
        .Z(c[115]) );
  AND \ADD_/FAINST[115].FA_/U3  ( .A(\ADD_/FAINST[115].FA_/n1 ), .B(
        \ADD_/FAINST[115].FA_/n2 ), .Z(\ADD_/FAINST[115].FA_/n3 ) );
  XOR \ADD_/FAINST[115].FA_/U2  ( .A(b[115]), .B(\ADD_/c[115] ), .Z(
        \ADD_/FAINST[115].FA_/n2 ) );
  XOR \ADD_/FAINST[115].FA_/U1  ( .A(a[115]), .B(\ADD_/c[115] ), .Z(
        \ADD_/FAINST[115].FA_/n1 ) );
  XOR \ADD_/FAINST[114].FA_/U5  ( .A(\ADD_/FAINST[114].FA_/n3 ), .B(
        \ADD_/c[114] ), .Z(\ADD_/c[115] ) );
  XOR \ADD_/FAINST[114].FA_/U4  ( .A(\ADD_/FAINST[114].FA_/n1 ), .B(b[114]), 
        .Z(c[114]) );
  AND \ADD_/FAINST[114].FA_/U3  ( .A(\ADD_/FAINST[114].FA_/n1 ), .B(
        \ADD_/FAINST[114].FA_/n2 ), .Z(\ADD_/FAINST[114].FA_/n3 ) );
  XOR \ADD_/FAINST[114].FA_/U2  ( .A(b[114]), .B(\ADD_/c[114] ), .Z(
        \ADD_/FAINST[114].FA_/n2 ) );
  XOR \ADD_/FAINST[114].FA_/U1  ( .A(a[114]), .B(\ADD_/c[114] ), .Z(
        \ADD_/FAINST[114].FA_/n1 ) );
  XOR \ADD_/FAINST[113].FA_/U5  ( .A(\ADD_/FAINST[113].FA_/n3 ), .B(
        \ADD_/c[113] ), .Z(\ADD_/c[114] ) );
  XOR \ADD_/FAINST[113].FA_/U4  ( .A(\ADD_/FAINST[113].FA_/n1 ), .B(b[113]), 
        .Z(c[113]) );
  AND \ADD_/FAINST[113].FA_/U3  ( .A(\ADD_/FAINST[113].FA_/n1 ), .B(
        \ADD_/FAINST[113].FA_/n2 ), .Z(\ADD_/FAINST[113].FA_/n3 ) );
  XOR \ADD_/FAINST[113].FA_/U2  ( .A(b[113]), .B(\ADD_/c[113] ), .Z(
        \ADD_/FAINST[113].FA_/n2 ) );
  XOR \ADD_/FAINST[113].FA_/U1  ( .A(a[113]), .B(\ADD_/c[113] ), .Z(
        \ADD_/FAINST[113].FA_/n1 ) );
  XOR \ADD_/FAINST[112].FA_/U5  ( .A(\ADD_/FAINST[112].FA_/n3 ), .B(
        \ADD_/c[112] ), .Z(\ADD_/c[113] ) );
  XOR \ADD_/FAINST[112].FA_/U4  ( .A(\ADD_/FAINST[112].FA_/n1 ), .B(b[112]), 
        .Z(c[112]) );
  AND \ADD_/FAINST[112].FA_/U3  ( .A(\ADD_/FAINST[112].FA_/n1 ), .B(
        \ADD_/FAINST[112].FA_/n2 ), .Z(\ADD_/FAINST[112].FA_/n3 ) );
  XOR \ADD_/FAINST[112].FA_/U2  ( .A(b[112]), .B(\ADD_/c[112] ), .Z(
        \ADD_/FAINST[112].FA_/n2 ) );
  XOR \ADD_/FAINST[112].FA_/U1  ( .A(a[112]), .B(\ADD_/c[112] ), .Z(
        \ADD_/FAINST[112].FA_/n1 ) );
  XOR \ADD_/FAINST[111].FA_/U5  ( .A(\ADD_/FAINST[111].FA_/n3 ), .B(
        \ADD_/c[111] ), .Z(\ADD_/c[112] ) );
  XOR \ADD_/FAINST[111].FA_/U4  ( .A(\ADD_/FAINST[111].FA_/n1 ), .B(b[111]), 
        .Z(c[111]) );
  AND \ADD_/FAINST[111].FA_/U3  ( .A(\ADD_/FAINST[111].FA_/n1 ), .B(
        \ADD_/FAINST[111].FA_/n2 ), .Z(\ADD_/FAINST[111].FA_/n3 ) );
  XOR \ADD_/FAINST[111].FA_/U2  ( .A(b[111]), .B(\ADD_/c[111] ), .Z(
        \ADD_/FAINST[111].FA_/n2 ) );
  XOR \ADD_/FAINST[111].FA_/U1  ( .A(a[111]), .B(\ADD_/c[111] ), .Z(
        \ADD_/FAINST[111].FA_/n1 ) );
  XOR \ADD_/FAINST[110].FA_/U5  ( .A(\ADD_/FAINST[110].FA_/n3 ), .B(
        \ADD_/c[110] ), .Z(\ADD_/c[111] ) );
  XOR \ADD_/FAINST[110].FA_/U4  ( .A(\ADD_/FAINST[110].FA_/n1 ), .B(b[110]), 
        .Z(c[110]) );
  AND \ADD_/FAINST[110].FA_/U3  ( .A(\ADD_/FAINST[110].FA_/n1 ), .B(
        \ADD_/FAINST[110].FA_/n2 ), .Z(\ADD_/FAINST[110].FA_/n3 ) );
  XOR \ADD_/FAINST[110].FA_/U2  ( .A(b[110]), .B(\ADD_/c[110] ), .Z(
        \ADD_/FAINST[110].FA_/n2 ) );
  XOR \ADD_/FAINST[110].FA_/U1  ( .A(a[110]), .B(\ADD_/c[110] ), .Z(
        \ADD_/FAINST[110].FA_/n1 ) );
  XOR \ADD_/FAINST[109].FA_/U5  ( .A(\ADD_/FAINST[109].FA_/n3 ), .B(
        \ADD_/c[109] ), .Z(\ADD_/c[110] ) );
  XOR \ADD_/FAINST[109].FA_/U4  ( .A(\ADD_/FAINST[109].FA_/n1 ), .B(b[109]), 
        .Z(c[109]) );
  AND \ADD_/FAINST[109].FA_/U3  ( .A(\ADD_/FAINST[109].FA_/n1 ), .B(
        \ADD_/FAINST[109].FA_/n2 ), .Z(\ADD_/FAINST[109].FA_/n3 ) );
  XOR \ADD_/FAINST[109].FA_/U2  ( .A(b[109]), .B(\ADD_/c[109] ), .Z(
        \ADD_/FAINST[109].FA_/n2 ) );
  XOR \ADD_/FAINST[109].FA_/U1  ( .A(a[109]), .B(\ADD_/c[109] ), .Z(
        \ADD_/FAINST[109].FA_/n1 ) );
  XOR \ADD_/FAINST[108].FA_/U5  ( .A(\ADD_/FAINST[108].FA_/n3 ), .B(
        \ADD_/c[108] ), .Z(\ADD_/c[109] ) );
  XOR \ADD_/FAINST[108].FA_/U4  ( .A(\ADD_/FAINST[108].FA_/n1 ), .B(b[108]), 
        .Z(c[108]) );
  AND \ADD_/FAINST[108].FA_/U3  ( .A(\ADD_/FAINST[108].FA_/n1 ), .B(
        \ADD_/FAINST[108].FA_/n2 ), .Z(\ADD_/FAINST[108].FA_/n3 ) );
  XOR \ADD_/FAINST[108].FA_/U2  ( .A(b[108]), .B(\ADD_/c[108] ), .Z(
        \ADD_/FAINST[108].FA_/n2 ) );
  XOR \ADD_/FAINST[108].FA_/U1  ( .A(a[108]), .B(\ADD_/c[108] ), .Z(
        \ADD_/FAINST[108].FA_/n1 ) );
  XOR \ADD_/FAINST[107].FA_/U5  ( .A(\ADD_/FAINST[107].FA_/n3 ), .B(
        \ADD_/c[107] ), .Z(\ADD_/c[108] ) );
  XOR \ADD_/FAINST[107].FA_/U4  ( .A(\ADD_/FAINST[107].FA_/n1 ), .B(b[107]), 
        .Z(c[107]) );
  AND \ADD_/FAINST[107].FA_/U3  ( .A(\ADD_/FAINST[107].FA_/n1 ), .B(
        \ADD_/FAINST[107].FA_/n2 ), .Z(\ADD_/FAINST[107].FA_/n3 ) );
  XOR \ADD_/FAINST[107].FA_/U2  ( .A(b[107]), .B(\ADD_/c[107] ), .Z(
        \ADD_/FAINST[107].FA_/n2 ) );
  XOR \ADD_/FAINST[107].FA_/U1  ( .A(a[107]), .B(\ADD_/c[107] ), .Z(
        \ADD_/FAINST[107].FA_/n1 ) );
  XOR \ADD_/FAINST[106].FA_/U5  ( .A(\ADD_/FAINST[106].FA_/n3 ), .B(
        \ADD_/c[106] ), .Z(\ADD_/c[107] ) );
  XOR \ADD_/FAINST[106].FA_/U4  ( .A(\ADD_/FAINST[106].FA_/n1 ), .B(b[106]), 
        .Z(c[106]) );
  AND \ADD_/FAINST[106].FA_/U3  ( .A(\ADD_/FAINST[106].FA_/n1 ), .B(
        \ADD_/FAINST[106].FA_/n2 ), .Z(\ADD_/FAINST[106].FA_/n3 ) );
  XOR \ADD_/FAINST[106].FA_/U2  ( .A(b[106]), .B(\ADD_/c[106] ), .Z(
        \ADD_/FAINST[106].FA_/n2 ) );
  XOR \ADD_/FAINST[106].FA_/U1  ( .A(a[106]), .B(\ADD_/c[106] ), .Z(
        \ADD_/FAINST[106].FA_/n1 ) );
  XOR \ADD_/FAINST[105].FA_/U5  ( .A(\ADD_/FAINST[105].FA_/n3 ), .B(
        \ADD_/c[105] ), .Z(\ADD_/c[106] ) );
  XOR \ADD_/FAINST[105].FA_/U4  ( .A(\ADD_/FAINST[105].FA_/n1 ), .B(b[105]), 
        .Z(c[105]) );
  AND \ADD_/FAINST[105].FA_/U3  ( .A(\ADD_/FAINST[105].FA_/n1 ), .B(
        \ADD_/FAINST[105].FA_/n2 ), .Z(\ADD_/FAINST[105].FA_/n3 ) );
  XOR \ADD_/FAINST[105].FA_/U2  ( .A(b[105]), .B(\ADD_/c[105] ), .Z(
        \ADD_/FAINST[105].FA_/n2 ) );
  XOR \ADD_/FAINST[105].FA_/U1  ( .A(a[105]), .B(\ADD_/c[105] ), .Z(
        \ADD_/FAINST[105].FA_/n1 ) );
  XOR \ADD_/FAINST[104].FA_/U5  ( .A(\ADD_/FAINST[104].FA_/n3 ), .B(
        \ADD_/c[104] ), .Z(\ADD_/c[105] ) );
  XOR \ADD_/FAINST[104].FA_/U4  ( .A(\ADD_/FAINST[104].FA_/n1 ), .B(b[104]), 
        .Z(c[104]) );
  AND \ADD_/FAINST[104].FA_/U3  ( .A(\ADD_/FAINST[104].FA_/n1 ), .B(
        \ADD_/FAINST[104].FA_/n2 ), .Z(\ADD_/FAINST[104].FA_/n3 ) );
  XOR \ADD_/FAINST[104].FA_/U2  ( .A(b[104]), .B(\ADD_/c[104] ), .Z(
        \ADD_/FAINST[104].FA_/n2 ) );
  XOR \ADD_/FAINST[104].FA_/U1  ( .A(a[104]), .B(\ADD_/c[104] ), .Z(
        \ADD_/FAINST[104].FA_/n1 ) );
  XOR \ADD_/FAINST[103].FA_/U5  ( .A(\ADD_/FAINST[103].FA_/n3 ), .B(
        \ADD_/c[103] ), .Z(\ADD_/c[104] ) );
  XOR \ADD_/FAINST[103].FA_/U4  ( .A(\ADD_/FAINST[103].FA_/n1 ), .B(b[103]), 
        .Z(c[103]) );
  AND \ADD_/FAINST[103].FA_/U3  ( .A(\ADD_/FAINST[103].FA_/n1 ), .B(
        \ADD_/FAINST[103].FA_/n2 ), .Z(\ADD_/FAINST[103].FA_/n3 ) );
  XOR \ADD_/FAINST[103].FA_/U2  ( .A(b[103]), .B(\ADD_/c[103] ), .Z(
        \ADD_/FAINST[103].FA_/n2 ) );
  XOR \ADD_/FAINST[103].FA_/U1  ( .A(a[103]), .B(\ADD_/c[103] ), .Z(
        \ADD_/FAINST[103].FA_/n1 ) );
  XOR \ADD_/FAINST[102].FA_/U5  ( .A(\ADD_/FAINST[102].FA_/n3 ), .B(
        \ADD_/c[102] ), .Z(\ADD_/c[103] ) );
  XOR \ADD_/FAINST[102].FA_/U4  ( .A(\ADD_/FAINST[102].FA_/n1 ), .B(b[102]), 
        .Z(c[102]) );
  AND \ADD_/FAINST[102].FA_/U3  ( .A(\ADD_/FAINST[102].FA_/n1 ), .B(
        \ADD_/FAINST[102].FA_/n2 ), .Z(\ADD_/FAINST[102].FA_/n3 ) );
  XOR \ADD_/FAINST[102].FA_/U2  ( .A(b[102]), .B(\ADD_/c[102] ), .Z(
        \ADD_/FAINST[102].FA_/n2 ) );
  XOR \ADD_/FAINST[102].FA_/U1  ( .A(a[102]), .B(\ADD_/c[102] ), .Z(
        \ADD_/FAINST[102].FA_/n1 ) );
  XOR \ADD_/FAINST[101].FA_/U5  ( .A(\ADD_/FAINST[101].FA_/n3 ), .B(
        \ADD_/c[101] ), .Z(\ADD_/c[102] ) );
  XOR \ADD_/FAINST[101].FA_/U4  ( .A(\ADD_/FAINST[101].FA_/n1 ), .B(b[101]), 
        .Z(c[101]) );
  AND \ADD_/FAINST[101].FA_/U3  ( .A(\ADD_/FAINST[101].FA_/n1 ), .B(
        \ADD_/FAINST[101].FA_/n2 ), .Z(\ADD_/FAINST[101].FA_/n3 ) );
  XOR \ADD_/FAINST[101].FA_/U2  ( .A(b[101]), .B(\ADD_/c[101] ), .Z(
        \ADD_/FAINST[101].FA_/n2 ) );
  XOR \ADD_/FAINST[101].FA_/U1  ( .A(a[101]), .B(\ADD_/c[101] ), .Z(
        \ADD_/FAINST[101].FA_/n1 ) );
  XOR \ADD_/FAINST[100].FA_/U5  ( .A(\ADD_/FAINST[100].FA_/n3 ), .B(
        \ADD_/c[100] ), .Z(\ADD_/c[101] ) );
  XOR \ADD_/FAINST[100].FA_/U4  ( .A(\ADD_/FAINST[100].FA_/n1 ), .B(b[100]), 
        .Z(c[100]) );
  AND \ADD_/FAINST[100].FA_/U3  ( .A(\ADD_/FAINST[100].FA_/n1 ), .B(
        \ADD_/FAINST[100].FA_/n2 ), .Z(\ADD_/FAINST[100].FA_/n3 ) );
  XOR \ADD_/FAINST[100].FA_/U2  ( .A(b[100]), .B(\ADD_/c[100] ), .Z(
        \ADD_/FAINST[100].FA_/n2 ) );
  XOR \ADD_/FAINST[100].FA_/U1  ( .A(a[100]), .B(\ADD_/c[100] ), .Z(
        \ADD_/FAINST[100].FA_/n1 ) );
  XOR \ADD_/FAINST[99].FA_/U5  ( .A(\ADD_/FAINST[99].FA_/n3 ), .B(\ADD_/c[99] ), .Z(\ADD_/c[100] ) );
  XOR \ADD_/FAINST[99].FA_/U4  ( .A(\ADD_/FAINST[99].FA_/n1 ), .B(b[99]), .Z(
        c[99]) );
  AND \ADD_/FAINST[99].FA_/U3  ( .A(\ADD_/FAINST[99].FA_/n1 ), .B(
        \ADD_/FAINST[99].FA_/n2 ), .Z(\ADD_/FAINST[99].FA_/n3 ) );
  XOR \ADD_/FAINST[99].FA_/U2  ( .A(b[99]), .B(\ADD_/c[99] ), .Z(
        \ADD_/FAINST[99].FA_/n2 ) );
  XOR \ADD_/FAINST[99].FA_/U1  ( .A(a[99]), .B(\ADD_/c[99] ), .Z(
        \ADD_/FAINST[99].FA_/n1 ) );
  XOR \ADD_/FAINST[98].FA_/U5  ( .A(\ADD_/FAINST[98].FA_/n3 ), .B(\ADD_/c[98] ), .Z(\ADD_/c[99] ) );
  XOR \ADD_/FAINST[98].FA_/U4  ( .A(\ADD_/FAINST[98].FA_/n1 ), .B(b[98]), .Z(
        c[98]) );
  AND \ADD_/FAINST[98].FA_/U3  ( .A(\ADD_/FAINST[98].FA_/n1 ), .B(
        \ADD_/FAINST[98].FA_/n2 ), .Z(\ADD_/FAINST[98].FA_/n3 ) );
  XOR \ADD_/FAINST[98].FA_/U2  ( .A(b[98]), .B(\ADD_/c[98] ), .Z(
        \ADD_/FAINST[98].FA_/n2 ) );
  XOR \ADD_/FAINST[98].FA_/U1  ( .A(a[98]), .B(\ADD_/c[98] ), .Z(
        \ADD_/FAINST[98].FA_/n1 ) );
  XOR \ADD_/FAINST[97].FA_/U5  ( .A(\ADD_/FAINST[97].FA_/n3 ), .B(\ADD_/c[97] ), .Z(\ADD_/c[98] ) );
  XOR \ADD_/FAINST[97].FA_/U4  ( .A(\ADD_/FAINST[97].FA_/n1 ), .B(b[97]), .Z(
        c[97]) );
  AND \ADD_/FAINST[97].FA_/U3  ( .A(\ADD_/FAINST[97].FA_/n1 ), .B(
        \ADD_/FAINST[97].FA_/n2 ), .Z(\ADD_/FAINST[97].FA_/n3 ) );
  XOR \ADD_/FAINST[97].FA_/U2  ( .A(b[97]), .B(\ADD_/c[97] ), .Z(
        \ADD_/FAINST[97].FA_/n2 ) );
  XOR \ADD_/FAINST[97].FA_/U1  ( .A(a[97]), .B(\ADD_/c[97] ), .Z(
        \ADD_/FAINST[97].FA_/n1 ) );
  XOR \ADD_/FAINST[96].FA_/U5  ( .A(\ADD_/FAINST[96].FA_/n3 ), .B(\ADD_/c[96] ), .Z(\ADD_/c[97] ) );
  XOR \ADD_/FAINST[96].FA_/U4  ( .A(\ADD_/FAINST[96].FA_/n1 ), .B(b[96]), .Z(
        c[96]) );
  AND \ADD_/FAINST[96].FA_/U3  ( .A(\ADD_/FAINST[96].FA_/n1 ), .B(
        \ADD_/FAINST[96].FA_/n2 ), .Z(\ADD_/FAINST[96].FA_/n3 ) );
  XOR \ADD_/FAINST[96].FA_/U2  ( .A(b[96]), .B(\ADD_/c[96] ), .Z(
        \ADD_/FAINST[96].FA_/n2 ) );
  XOR \ADD_/FAINST[96].FA_/U1  ( .A(a[96]), .B(\ADD_/c[96] ), .Z(
        \ADD_/FAINST[96].FA_/n1 ) );
  XOR \ADD_/FAINST[95].FA_/U5  ( .A(\ADD_/FAINST[95].FA_/n3 ), .B(\ADD_/c[95] ), .Z(\ADD_/c[96] ) );
  XOR \ADD_/FAINST[95].FA_/U4  ( .A(\ADD_/FAINST[95].FA_/n1 ), .B(b[95]), .Z(
        c[95]) );
  AND \ADD_/FAINST[95].FA_/U3  ( .A(\ADD_/FAINST[95].FA_/n1 ), .B(
        \ADD_/FAINST[95].FA_/n2 ), .Z(\ADD_/FAINST[95].FA_/n3 ) );
  XOR \ADD_/FAINST[95].FA_/U2  ( .A(b[95]), .B(\ADD_/c[95] ), .Z(
        \ADD_/FAINST[95].FA_/n2 ) );
  XOR \ADD_/FAINST[95].FA_/U1  ( .A(a[95]), .B(\ADD_/c[95] ), .Z(
        \ADD_/FAINST[95].FA_/n1 ) );
  XOR \ADD_/FAINST[94].FA_/U5  ( .A(\ADD_/FAINST[94].FA_/n3 ), .B(\ADD_/c[94] ), .Z(\ADD_/c[95] ) );
  XOR \ADD_/FAINST[94].FA_/U4  ( .A(\ADD_/FAINST[94].FA_/n1 ), .B(b[94]), .Z(
        c[94]) );
  AND \ADD_/FAINST[94].FA_/U3  ( .A(\ADD_/FAINST[94].FA_/n1 ), .B(
        \ADD_/FAINST[94].FA_/n2 ), .Z(\ADD_/FAINST[94].FA_/n3 ) );
  XOR \ADD_/FAINST[94].FA_/U2  ( .A(b[94]), .B(\ADD_/c[94] ), .Z(
        \ADD_/FAINST[94].FA_/n2 ) );
  XOR \ADD_/FAINST[94].FA_/U1  ( .A(a[94]), .B(\ADD_/c[94] ), .Z(
        \ADD_/FAINST[94].FA_/n1 ) );
  XOR \ADD_/FAINST[93].FA_/U5  ( .A(\ADD_/FAINST[93].FA_/n3 ), .B(\ADD_/c[93] ), .Z(\ADD_/c[94] ) );
  XOR \ADD_/FAINST[93].FA_/U4  ( .A(\ADD_/FAINST[93].FA_/n1 ), .B(b[93]), .Z(
        c[93]) );
  AND \ADD_/FAINST[93].FA_/U3  ( .A(\ADD_/FAINST[93].FA_/n1 ), .B(
        \ADD_/FAINST[93].FA_/n2 ), .Z(\ADD_/FAINST[93].FA_/n3 ) );
  XOR \ADD_/FAINST[93].FA_/U2  ( .A(b[93]), .B(\ADD_/c[93] ), .Z(
        \ADD_/FAINST[93].FA_/n2 ) );
  XOR \ADD_/FAINST[93].FA_/U1  ( .A(a[93]), .B(\ADD_/c[93] ), .Z(
        \ADD_/FAINST[93].FA_/n1 ) );
  XOR \ADD_/FAINST[92].FA_/U5  ( .A(\ADD_/FAINST[92].FA_/n3 ), .B(\ADD_/c[92] ), .Z(\ADD_/c[93] ) );
  XOR \ADD_/FAINST[92].FA_/U4  ( .A(\ADD_/FAINST[92].FA_/n1 ), .B(b[92]), .Z(
        c[92]) );
  AND \ADD_/FAINST[92].FA_/U3  ( .A(\ADD_/FAINST[92].FA_/n1 ), .B(
        \ADD_/FAINST[92].FA_/n2 ), .Z(\ADD_/FAINST[92].FA_/n3 ) );
  XOR \ADD_/FAINST[92].FA_/U2  ( .A(b[92]), .B(\ADD_/c[92] ), .Z(
        \ADD_/FAINST[92].FA_/n2 ) );
  XOR \ADD_/FAINST[92].FA_/U1  ( .A(a[92]), .B(\ADD_/c[92] ), .Z(
        \ADD_/FAINST[92].FA_/n1 ) );
  XOR \ADD_/FAINST[91].FA_/U5  ( .A(\ADD_/FAINST[91].FA_/n3 ), .B(\ADD_/c[91] ), .Z(\ADD_/c[92] ) );
  XOR \ADD_/FAINST[91].FA_/U4  ( .A(\ADD_/FAINST[91].FA_/n1 ), .B(b[91]), .Z(
        c[91]) );
  AND \ADD_/FAINST[91].FA_/U3  ( .A(\ADD_/FAINST[91].FA_/n1 ), .B(
        \ADD_/FAINST[91].FA_/n2 ), .Z(\ADD_/FAINST[91].FA_/n3 ) );
  XOR \ADD_/FAINST[91].FA_/U2  ( .A(b[91]), .B(\ADD_/c[91] ), .Z(
        \ADD_/FAINST[91].FA_/n2 ) );
  XOR \ADD_/FAINST[91].FA_/U1  ( .A(a[91]), .B(\ADD_/c[91] ), .Z(
        \ADD_/FAINST[91].FA_/n1 ) );
  XOR \ADD_/FAINST[90].FA_/U5  ( .A(\ADD_/FAINST[90].FA_/n3 ), .B(\ADD_/c[90] ), .Z(\ADD_/c[91] ) );
  XOR \ADD_/FAINST[90].FA_/U4  ( .A(\ADD_/FAINST[90].FA_/n1 ), .B(b[90]), .Z(
        c[90]) );
  AND \ADD_/FAINST[90].FA_/U3  ( .A(\ADD_/FAINST[90].FA_/n1 ), .B(
        \ADD_/FAINST[90].FA_/n2 ), .Z(\ADD_/FAINST[90].FA_/n3 ) );
  XOR \ADD_/FAINST[90].FA_/U2  ( .A(b[90]), .B(\ADD_/c[90] ), .Z(
        \ADD_/FAINST[90].FA_/n2 ) );
  XOR \ADD_/FAINST[90].FA_/U1  ( .A(a[90]), .B(\ADD_/c[90] ), .Z(
        \ADD_/FAINST[90].FA_/n1 ) );
  XOR \ADD_/FAINST[89].FA_/U5  ( .A(\ADD_/FAINST[89].FA_/n3 ), .B(\ADD_/c[89] ), .Z(\ADD_/c[90] ) );
  XOR \ADD_/FAINST[89].FA_/U4  ( .A(\ADD_/FAINST[89].FA_/n1 ), .B(b[89]), .Z(
        c[89]) );
  AND \ADD_/FAINST[89].FA_/U3  ( .A(\ADD_/FAINST[89].FA_/n1 ), .B(
        \ADD_/FAINST[89].FA_/n2 ), .Z(\ADD_/FAINST[89].FA_/n3 ) );
  XOR \ADD_/FAINST[89].FA_/U2  ( .A(b[89]), .B(\ADD_/c[89] ), .Z(
        \ADD_/FAINST[89].FA_/n2 ) );
  XOR \ADD_/FAINST[89].FA_/U1  ( .A(a[89]), .B(\ADD_/c[89] ), .Z(
        \ADD_/FAINST[89].FA_/n1 ) );
  XOR \ADD_/FAINST[88].FA_/U5  ( .A(\ADD_/FAINST[88].FA_/n3 ), .B(\ADD_/c[88] ), .Z(\ADD_/c[89] ) );
  XOR \ADD_/FAINST[88].FA_/U4  ( .A(\ADD_/FAINST[88].FA_/n1 ), .B(b[88]), .Z(
        c[88]) );
  AND \ADD_/FAINST[88].FA_/U3  ( .A(\ADD_/FAINST[88].FA_/n1 ), .B(
        \ADD_/FAINST[88].FA_/n2 ), .Z(\ADD_/FAINST[88].FA_/n3 ) );
  XOR \ADD_/FAINST[88].FA_/U2  ( .A(b[88]), .B(\ADD_/c[88] ), .Z(
        \ADD_/FAINST[88].FA_/n2 ) );
  XOR \ADD_/FAINST[88].FA_/U1  ( .A(a[88]), .B(\ADD_/c[88] ), .Z(
        \ADD_/FAINST[88].FA_/n1 ) );
  XOR \ADD_/FAINST[87].FA_/U5  ( .A(\ADD_/FAINST[87].FA_/n3 ), .B(\ADD_/c[87] ), .Z(\ADD_/c[88] ) );
  XOR \ADD_/FAINST[87].FA_/U4  ( .A(\ADD_/FAINST[87].FA_/n1 ), .B(b[87]), .Z(
        c[87]) );
  AND \ADD_/FAINST[87].FA_/U3  ( .A(\ADD_/FAINST[87].FA_/n1 ), .B(
        \ADD_/FAINST[87].FA_/n2 ), .Z(\ADD_/FAINST[87].FA_/n3 ) );
  XOR \ADD_/FAINST[87].FA_/U2  ( .A(b[87]), .B(\ADD_/c[87] ), .Z(
        \ADD_/FAINST[87].FA_/n2 ) );
  XOR \ADD_/FAINST[87].FA_/U1  ( .A(a[87]), .B(\ADD_/c[87] ), .Z(
        \ADD_/FAINST[87].FA_/n1 ) );
  XOR \ADD_/FAINST[86].FA_/U5  ( .A(\ADD_/FAINST[86].FA_/n3 ), .B(\ADD_/c[86] ), .Z(\ADD_/c[87] ) );
  XOR \ADD_/FAINST[86].FA_/U4  ( .A(\ADD_/FAINST[86].FA_/n1 ), .B(b[86]), .Z(
        c[86]) );
  AND \ADD_/FAINST[86].FA_/U3  ( .A(\ADD_/FAINST[86].FA_/n1 ), .B(
        \ADD_/FAINST[86].FA_/n2 ), .Z(\ADD_/FAINST[86].FA_/n3 ) );
  XOR \ADD_/FAINST[86].FA_/U2  ( .A(b[86]), .B(\ADD_/c[86] ), .Z(
        \ADD_/FAINST[86].FA_/n2 ) );
  XOR \ADD_/FAINST[86].FA_/U1  ( .A(a[86]), .B(\ADD_/c[86] ), .Z(
        \ADD_/FAINST[86].FA_/n1 ) );
  XOR \ADD_/FAINST[85].FA_/U5  ( .A(\ADD_/FAINST[85].FA_/n3 ), .B(\ADD_/c[85] ), .Z(\ADD_/c[86] ) );
  XOR \ADD_/FAINST[85].FA_/U4  ( .A(\ADD_/FAINST[85].FA_/n1 ), .B(b[85]), .Z(
        c[85]) );
  AND \ADD_/FAINST[85].FA_/U3  ( .A(\ADD_/FAINST[85].FA_/n1 ), .B(
        \ADD_/FAINST[85].FA_/n2 ), .Z(\ADD_/FAINST[85].FA_/n3 ) );
  XOR \ADD_/FAINST[85].FA_/U2  ( .A(b[85]), .B(\ADD_/c[85] ), .Z(
        \ADD_/FAINST[85].FA_/n2 ) );
  XOR \ADD_/FAINST[85].FA_/U1  ( .A(a[85]), .B(\ADD_/c[85] ), .Z(
        \ADD_/FAINST[85].FA_/n1 ) );
  XOR \ADD_/FAINST[84].FA_/U5  ( .A(\ADD_/FAINST[84].FA_/n3 ), .B(\ADD_/c[84] ), .Z(\ADD_/c[85] ) );
  XOR \ADD_/FAINST[84].FA_/U4  ( .A(\ADD_/FAINST[84].FA_/n1 ), .B(b[84]), .Z(
        c[84]) );
  AND \ADD_/FAINST[84].FA_/U3  ( .A(\ADD_/FAINST[84].FA_/n1 ), .B(
        \ADD_/FAINST[84].FA_/n2 ), .Z(\ADD_/FAINST[84].FA_/n3 ) );
  XOR \ADD_/FAINST[84].FA_/U2  ( .A(b[84]), .B(\ADD_/c[84] ), .Z(
        \ADD_/FAINST[84].FA_/n2 ) );
  XOR \ADD_/FAINST[84].FA_/U1  ( .A(a[84]), .B(\ADD_/c[84] ), .Z(
        \ADD_/FAINST[84].FA_/n1 ) );
  XOR \ADD_/FAINST[83].FA_/U5  ( .A(\ADD_/FAINST[83].FA_/n3 ), .B(\ADD_/c[83] ), .Z(\ADD_/c[84] ) );
  XOR \ADD_/FAINST[83].FA_/U4  ( .A(\ADD_/FAINST[83].FA_/n1 ), .B(b[83]), .Z(
        c[83]) );
  AND \ADD_/FAINST[83].FA_/U3  ( .A(\ADD_/FAINST[83].FA_/n1 ), .B(
        \ADD_/FAINST[83].FA_/n2 ), .Z(\ADD_/FAINST[83].FA_/n3 ) );
  XOR \ADD_/FAINST[83].FA_/U2  ( .A(b[83]), .B(\ADD_/c[83] ), .Z(
        \ADD_/FAINST[83].FA_/n2 ) );
  XOR \ADD_/FAINST[83].FA_/U1  ( .A(a[83]), .B(\ADD_/c[83] ), .Z(
        \ADD_/FAINST[83].FA_/n1 ) );
  XOR \ADD_/FAINST[82].FA_/U5  ( .A(\ADD_/FAINST[82].FA_/n3 ), .B(\ADD_/c[82] ), .Z(\ADD_/c[83] ) );
  XOR \ADD_/FAINST[82].FA_/U4  ( .A(\ADD_/FAINST[82].FA_/n1 ), .B(b[82]), .Z(
        c[82]) );
  AND \ADD_/FAINST[82].FA_/U3  ( .A(\ADD_/FAINST[82].FA_/n1 ), .B(
        \ADD_/FAINST[82].FA_/n2 ), .Z(\ADD_/FAINST[82].FA_/n3 ) );
  XOR \ADD_/FAINST[82].FA_/U2  ( .A(b[82]), .B(\ADD_/c[82] ), .Z(
        \ADD_/FAINST[82].FA_/n2 ) );
  XOR \ADD_/FAINST[82].FA_/U1  ( .A(a[82]), .B(\ADD_/c[82] ), .Z(
        \ADD_/FAINST[82].FA_/n1 ) );
  XOR \ADD_/FAINST[81].FA_/U5  ( .A(\ADD_/FAINST[81].FA_/n3 ), .B(\ADD_/c[81] ), .Z(\ADD_/c[82] ) );
  XOR \ADD_/FAINST[81].FA_/U4  ( .A(\ADD_/FAINST[81].FA_/n1 ), .B(b[81]), .Z(
        c[81]) );
  AND \ADD_/FAINST[81].FA_/U3  ( .A(\ADD_/FAINST[81].FA_/n1 ), .B(
        \ADD_/FAINST[81].FA_/n2 ), .Z(\ADD_/FAINST[81].FA_/n3 ) );
  XOR \ADD_/FAINST[81].FA_/U2  ( .A(b[81]), .B(\ADD_/c[81] ), .Z(
        \ADD_/FAINST[81].FA_/n2 ) );
  XOR \ADD_/FAINST[81].FA_/U1  ( .A(a[81]), .B(\ADD_/c[81] ), .Z(
        \ADD_/FAINST[81].FA_/n1 ) );
  XOR \ADD_/FAINST[80].FA_/U5  ( .A(\ADD_/FAINST[80].FA_/n3 ), .B(\ADD_/c[80] ), .Z(\ADD_/c[81] ) );
  XOR \ADD_/FAINST[80].FA_/U4  ( .A(\ADD_/FAINST[80].FA_/n1 ), .B(b[80]), .Z(
        c[80]) );
  AND \ADD_/FAINST[80].FA_/U3  ( .A(\ADD_/FAINST[80].FA_/n1 ), .B(
        \ADD_/FAINST[80].FA_/n2 ), .Z(\ADD_/FAINST[80].FA_/n3 ) );
  XOR \ADD_/FAINST[80].FA_/U2  ( .A(b[80]), .B(\ADD_/c[80] ), .Z(
        \ADD_/FAINST[80].FA_/n2 ) );
  XOR \ADD_/FAINST[80].FA_/U1  ( .A(a[80]), .B(\ADD_/c[80] ), .Z(
        \ADD_/FAINST[80].FA_/n1 ) );
  XOR \ADD_/FAINST[79].FA_/U5  ( .A(\ADD_/FAINST[79].FA_/n3 ), .B(\ADD_/c[79] ), .Z(\ADD_/c[80] ) );
  XOR \ADD_/FAINST[79].FA_/U4  ( .A(\ADD_/FAINST[79].FA_/n1 ), .B(b[79]), .Z(
        c[79]) );
  AND \ADD_/FAINST[79].FA_/U3  ( .A(\ADD_/FAINST[79].FA_/n1 ), .B(
        \ADD_/FAINST[79].FA_/n2 ), .Z(\ADD_/FAINST[79].FA_/n3 ) );
  XOR \ADD_/FAINST[79].FA_/U2  ( .A(b[79]), .B(\ADD_/c[79] ), .Z(
        \ADD_/FAINST[79].FA_/n2 ) );
  XOR \ADD_/FAINST[79].FA_/U1  ( .A(a[79]), .B(\ADD_/c[79] ), .Z(
        \ADD_/FAINST[79].FA_/n1 ) );
  XOR \ADD_/FAINST[78].FA_/U5  ( .A(\ADD_/FAINST[78].FA_/n3 ), .B(\ADD_/c[78] ), .Z(\ADD_/c[79] ) );
  XOR \ADD_/FAINST[78].FA_/U4  ( .A(\ADD_/FAINST[78].FA_/n1 ), .B(b[78]), .Z(
        c[78]) );
  AND \ADD_/FAINST[78].FA_/U3  ( .A(\ADD_/FAINST[78].FA_/n1 ), .B(
        \ADD_/FAINST[78].FA_/n2 ), .Z(\ADD_/FAINST[78].FA_/n3 ) );
  XOR \ADD_/FAINST[78].FA_/U2  ( .A(b[78]), .B(\ADD_/c[78] ), .Z(
        \ADD_/FAINST[78].FA_/n2 ) );
  XOR \ADD_/FAINST[78].FA_/U1  ( .A(a[78]), .B(\ADD_/c[78] ), .Z(
        \ADD_/FAINST[78].FA_/n1 ) );
  XOR \ADD_/FAINST[77].FA_/U5  ( .A(\ADD_/FAINST[77].FA_/n3 ), .B(\ADD_/c[77] ), .Z(\ADD_/c[78] ) );
  XOR \ADD_/FAINST[77].FA_/U4  ( .A(\ADD_/FAINST[77].FA_/n1 ), .B(b[77]), .Z(
        c[77]) );
  AND \ADD_/FAINST[77].FA_/U3  ( .A(\ADD_/FAINST[77].FA_/n1 ), .B(
        \ADD_/FAINST[77].FA_/n2 ), .Z(\ADD_/FAINST[77].FA_/n3 ) );
  XOR \ADD_/FAINST[77].FA_/U2  ( .A(b[77]), .B(\ADD_/c[77] ), .Z(
        \ADD_/FAINST[77].FA_/n2 ) );
  XOR \ADD_/FAINST[77].FA_/U1  ( .A(a[77]), .B(\ADD_/c[77] ), .Z(
        \ADD_/FAINST[77].FA_/n1 ) );
  XOR \ADD_/FAINST[76].FA_/U5  ( .A(\ADD_/FAINST[76].FA_/n3 ), .B(\ADD_/c[76] ), .Z(\ADD_/c[77] ) );
  XOR \ADD_/FAINST[76].FA_/U4  ( .A(\ADD_/FAINST[76].FA_/n1 ), .B(b[76]), .Z(
        c[76]) );
  AND \ADD_/FAINST[76].FA_/U3  ( .A(\ADD_/FAINST[76].FA_/n1 ), .B(
        \ADD_/FAINST[76].FA_/n2 ), .Z(\ADD_/FAINST[76].FA_/n3 ) );
  XOR \ADD_/FAINST[76].FA_/U2  ( .A(b[76]), .B(\ADD_/c[76] ), .Z(
        \ADD_/FAINST[76].FA_/n2 ) );
  XOR \ADD_/FAINST[76].FA_/U1  ( .A(a[76]), .B(\ADD_/c[76] ), .Z(
        \ADD_/FAINST[76].FA_/n1 ) );
  XOR \ADD_/FAINST[75].FA_/U5  ( .A(\ADD_/FAINST[75].FA_/n3 ), .B(\ADD_/c[75] ), .Z(\ADD_/c[76] ) );
  XOR \ADD_/FAINST[75].FA_/U4  ( .A(\ADD_/FAINST[75].FA_/n1 ), .B(b[75]), .Z(
        c[75]) );
  AND \ADD_/FAINST[75].FA_/U3  ( .A(\ADD_/FAINST[75].FA_/n1 ), .B(
        \ADD_/FAINST[75].FA_/n2 ), .Z(\ADD_/FAINST[75].FA_/n3 ) );
  XOR \ADD_/FAINST[75].FA_/U2  ( .A(b[75]), .B(\ADD_/c[75] ), .Z(
        \ADD_/FAINST[75].FA_/n2 ) );
  XOR \ADD_/FAINST[75].FA_/U1  ( .A(a[75]), .B(\ADD_/c[75] ), .Z(
        \ADD_/FAINST[75].FA_/n1 ) );
  XOR \ADD_/FAINST[74].FA_/U5  ( .A(\ADD_/FAINST[74].FA_/n3 ), .B(\ADD_/c[74] ), .Z(\ADD_/c[75] ) );
  XOR \ADD_/FAINST[74].FA_/U4  ( .A(\ADD_/FAINST[74].FA_/n1 ), .B(b[74]), .Z(
        c[74]) );
  AND \ADD_/FAINST[74].FA_/U3  ( .A(\ADD_/FAINST[74].FA_/n1 ), .B(
        \ADD_/FAINST[74].FA_/n2 ), .Z(\ADD_/FAINST[74].FA_/n3 ) );
  XOR \ADD_/FAINST[74].FA_/U2  ( .A(b[74]), .B(\ADD_/c[74] ), .Z(
        \ADD_/FAINST[74].FA_/n2 ) );
  XOR \ADD_/FAINST[74].FA_/U1  ( .A(a[74]), .B(\ADD_/c[74] ), .Z(
        \ADD_/FAINST[74].FA_/n1 ) );
  XOR \ADD_/FAINST[73].FA_/U5  ( .A(\ADD_/FAINST[73].FA_/n3 ), .B(\ADD_/c[73] ), .Z(\ADD_/c[74] ) );
  XOR \ADD_/FAINST[73].FA_/U4  ( .A(\ADD_/FAINST[73].FA_/n1 ), .B(b[73]), .Z(
        c[73]) );
  AND \ADD_/FAINST[73].FA_/U3  ( .A(\ADD_/FAINST[73].FA_/n1 ), .B(
        \ADD_/FAINST[73].FA_/n2 ), .Z(\ADD_/FAINST[73].FA_/n3 ) );
  XOR \ADD_/FAINST[73].FA_/U2  ( .A(b[73]), .B(\ADD_/c[73] ), .Z(
        \ADD_/FAINST[73].FA_/n2 ) );
  XOR \ADD_/FAINST[73].FA_/U1  ( .A(a[73]), .B(\ADD_/c[73] ), .Z(
        \ADD_/FAINST[73].FA_/n1 ) );
  XOR \ADD_/FAINST[72].FA_/U5  ( .A(\ADD_/FAINST[72].FA_/n3 ), .B(\ADD_/c[72] ), .Z(\ADD_/c[73] ) );
  XOR \ADD_/FAINST[72].FA_/U4  ( .A(\ADD_/FAINST[72].FA_/n1 ), .B(b[72]), .Z(
        c[72]) );
  AND \ADD_/FAINST[72].FA_/U3  ( .A(\ADD_/FAINST[72].FA_/n1 ), .B(
        \ADD_/FAINST[72].FA_/n2 ), .Z(\ADD_/FAINST[72].FA_/n3 ) );
  XOR \ADD_/FAINST[72].FA_/U2  ( .A(b[72]), .B(\ADD_/c[72] ), .Z(
        \ADD_/FAINST[72].FA_/n2 ) );
  XOR \ADD_/FAINST[72].FA_/U1  ( .A(a[72]), .B(\ADD_/c[72] ), .Z(
        \ADD_/FAINST[72].FA_/n1 ) );
  XOR \ADD_/FAINST[71].FA_/U5  ( .A(\ADD_/FAINST[71].FA_/n3 ), .B(\ADD_/c[71] ), .Z(\ADD_/c[72] ) );
  XOR \ADD_/FAINST[71].FA_/U4  ( .A(\ADD_/FAINST[71].FA_/n1 ), .B(b[71]), .Z(
        c[71]) );
  AND \ADD_/FAINST[71].FA_/U3  ( .A(\ADD_/FAINST[71].FA_/n1 ), .B(
        \ADD_/FAINST[71].FA_/n2 ), .Z(\ADD_/FAINST[71].FA_/n3 ) );
  XOR \ADD_/FAINST[71].FA_/U2  ( .A(b[71]), .B(\ADD_/c[71] ), .Z(
        \ADD_/FAINST[71].FA_/n2 ) );
  XOR \ADD_/FAINST[71].FA_/U1  ( .A(a[71]), .B(\ADD_/c[71] ), .Z(
        \ADD_/FAINST[71].FA_/n1 ) );
  XOR \ADD_/FAINST[70].FA_/U5  ( .A(\ADD_/FAINST[70].FA_/n3 ), .B(\ADD_/c[70] ), .Z(\ADD_/c[71] ) );
  XOR \ADD_/FAINST[70].FA_/U4  ( .A(\ADD_/FAINST[70].FA_/n1 ), .B(b[70]), .Z(
        c[70]) );
  AND \ADD_/FAINST[70].FA_/U3  ( .A(\ADD_/FAINST[70].FA_/n1 ), .B(
        \ADD_/FAINST[70].FA_/n2 ), .Z(\ADD_/FAINST[70].FA_/n3 ) );
  XOR \ADD_/FAINST[70].FA_/U2  ( .A(b[70]), .B(\ADD_/c[70] ), .Z(
        \ADD_/FAINST[70].FA_/n2 ) );
  XOR \ADD_/FAINST[70].FA_/U1  ( .A(a[70]), .B(\ADD_/c[70] ), .Z(
        \ADD_/FAINST[70].FA_/n1 ) );
  XOR \ADD_/FAINST[69].FA_/U5  ( .A(\ADD_/FAINST[69].FA_/n3 ), .B(\ADD_/c[69] ), .Z(\ADD_/c[70] ) );
  XOR \ADD_/FAINST[69].FA_/U4  ( .A(\ADD_/FAINST[69].FA_/n1 ), .B(b[69]), .Z(
        c[69]) );
  AND \ADD_/FAINST[69].FA_/U3  ( .A(\ADD_/FAINST[69].FA_/n1 ), .B(
        \ADD_/FAINST[69].FA_/n2 ), .Z(\ADD_/FAINST[69].FA_/n3 ) );
  XOR \ADD_/FAINST[69].FA_/U2  ( .A(b[69]), .B(\ADD_/c[69] ), .Z(
        \ADD_/FAINST[69].FA_/n2 ) );
  XOR \ADD_/FAINST[69].FA_/U1  ( .A(a[69]), .B(\ADD_/c[69] ), .Z(
        \ADD_/FAINST[69].FA_/n1 ) );
  XOR \ADD_/FAINST[68].FA_/U5  ( .A(\ADD_/FAINST[68].FA_/n3 ), .B(\ADD_/c[68] ), .Z(\ADD_/c[69] ) );
  XOR \ADD_/FAINST[68].FA_/U4  ( .A(\ADD_/FAINST[68].FA_/n1 ), .B(b[68]), .Z(
        c[68]) );
  AND \ADD_/FAINST[68].FA_/U3  ( .A(\ADD_/FAINST[68].FA_/n1 ), .B(
        \ADD_/FAINST[68].FA_/n2 ), .Z(\ADD_/FAINST[68].FA_/n3 ) );
  XOR \ADD_/FAINST[68].FA_/U2  ( .A(b[68]), .B(\ADD_/c[68] ), .Z(
        \ADD_/FAINST[68].FA_/n2 ) );
  XOR \ADD_/FAINST[68].FA_/U1  ( .A(a[68]), .B(\ADD_/c[68] ), .Z(
        \ADD_/FAINST[68].FA_/n1 ) );
  XOR \ADD_/FAINST[67].FA_/U5  ( .A(\ADD_/FAINST[67].FA_/n3 ), .B(\ADD_/c[67] ), .Z(\ADD_/c[68] ) );
  XOR \ADD_/FAINST[67].FA_/U4  ( .A(\ADD_/FAINST[67].FA_/n1 ), .B(b[67]), .Z(
        c[67]) );
  AND \ADD_/FAINST[67].FA_/U3  ( .A(\ADD_/FAINST[67].FA_/n1 ), .B(
        \ADD_/FAINST[67].FA_/n2 ), .Z(\ADD_/FAINST[67].FA_/n3 ) );
  XOR \ADD_/FAINST[67].FA_/U2  ( .A(b[67]), .B(\ADD_/c[67] ), .Z(
        \ADD_/FAINST[67].FA_/n2 ) );
  XOR \ADD_/FAINST[67].FA_/U1  ( .A(a[67]), .B(\ADD_/c[67] ), .Z(
        \ADD_/FAINST[67].FA_/n1 ) );
  XOR \ADD_/FAINST[66].FA_/U5  ( .A(\ADD_/FAINST[66].FA_/n3 ), .B(\ADD_/c[66] ), .Z(\ADD_/c[67] ) );
  XOR \ADD_/FAINST[66].FA_/U4  ( .A(\ADD_/FAINST[66].FA_/n1 ), .B(b[66]), .Z(
        c[66]) );
  AND \ADD_/FAINST[66].FA_/U3  ( .A(\ADD_/FAINST[66].FA_/n1 ), .B(
        \ADD_/FAINST[66].FA_/n2 ), .Z(\ADD_/FAINST[66].FA_/n3 ) );
  XOR \ADD_/FAINST[66].FA_/U2  ( .A(b[66]), .B(\ADD_/c[66] ), .Z(
        \ADD_/FAINST[66].FA_/n2 ) );
  XOR \ADD_/FAINST[66].FA_/U1  ( .A(a[66]), .B(\ADD_/c[66] ), .Z(
        \ADD_/FAINST[66].FA_/n1 ) );
  XOR \ADD_/FAINST[65].FA_/U5  ( .A(\ADD_/FAINST[65].FA_/n3 ), .B(\ADD_/c[65] ), .Z(\ADD_/c[66] ) );
  XOR \ADD_/FAINST[65].FA_/U4  ( .A(\ADD_/FAINST[65].FA_/n1 ), .B(b[65]), .Z(
        c[65]) );
  AND \ADD_/FAINST[65].FA_/U3  ( .A(\ADD_/FAINST[65].FA_/n1 ), .B(
        \ADD_/FAINST[65].FA_/n2 ), .Z(\ADD_/FAINST[65].FA_/n3 ) );
  XOR \ADD_/FAINST[65].FA_/U2  ( .A(b[65]), .B(\ADD_/c[65] ), .Z(
        \ADD_/FAINST[65].FA_/n2 ) );
  XOR \ADD_/FAINST[65].FA_/U1  ( .A(a[65]), .B(\ADD_/c[65] ), .Z(
        \ADD_/FAINST[65].FA_/n1 ) );
  XOR \ADD_/FAINST[64].FA_/U5  ( .A(\ADD_/FAINST[64].FA_/n3 ), .B(\ADD_/c[64] ), .Z(\ADD_/c[65] ) );
  XOR \ADD_/FAINST[64].FA_/U4  ( .A(\ADD_/FAINST[64].FA_/n1 ), .B(b[64]), .Z(
        c[64]) );
  AND \ADD_/FAINST[64].FA_/U3  ( .A(\ADD_/FAINST[64].FA_/n1 ), .B(
        \ADD_/FAINST[64].FA_/n2 ), .Z(\ADD_/FAINST[64].FA_/n3 ) );
  XOR \ADD_/FAINST[64].FA_/U2  ( .A(b[64]), .B(\ADD_/c[64] ), .Z(
        \ADD_/FAINST[64].FA_/n2 ) );
  XOR \ADD_/FAINST[64].FA_/U1  ( .A(a[64]), .B(\ADD_/c[64] ), .Z(
        \ADD_/FAINST[64].FA_/n1 ) );
  XOR \ADD_/FAINST[63].FA_/U5  ( .A(\ADD_/FAINST[63].FA_/n3 ), .B(\ADD_/c[63] ), .Z(\ADD_/c[64] ) );
  XOR \ADD_/FAINST[63].FA_/U4  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(b[63]), .Z(
        c[63]) );
  AND \ADD_/FAINST[63].FA_/U3  ( .A(\ADD_/FAINST[63].FA_/n1 ), .B(
        \ADD_/FAINST[63].FA_/n2 ), .Z(\ADD_/FAINST[63].FA_/n3 ) );
  XOR \ADD_/FAINST[63].FA_/U2  ( .A(b[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n2 ) );
  XOR \ADD_/FAINST[63].FA_/U1  ( .A(a[63]), .B(\ADD_/c[63] ), .Z(
        \ADD_/FAINST[63].FA_/n1 ) );
  XOR \ADD_/FAINST[62].FA_/U5  ( .A(\ADD_/FAINST[62].FA_/n3 ), .B(\ADD_/c[62] ), .Z(\ADD_/c[63] ) );
  XOR \ADD_/FAINST[62].FA_/U4  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(b[62]), .Z(
        c[62]) );
  AND \ADD_/FAINST[62].FA_/U3  ( .A(\ADD_/FAINST[62].FA_/n1 ), .B(
        \ADD_/FAINST[62].FA_/n2 ), .Z(\ADD_/FAINST[62].FA_/n3 ) );
  XOR \ADD_/FAINST[62].FA_/U2  ( .A(b[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n2 ) );
  XOR \ADD_/FAINST[62].FA_/U1  ( .A(a[62]), .B(\ADD_/c[62] ), .Z(
        \ADD_/FAINST[62].FA_/n1 ) );
  XOR \ADD_/FAINST[61].FA_/U5  ( .A(\ADD_/FAINST[61].FA_/n3 ), .B(\ADD_/c[61] ), .Z(\ADD_/c[62] ) );
  XOR \ADD_/FAINST[61].FA_/U4  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(b[61]), .Z(
        c[61]) );
  AND \ADD_/FAINST[61].FA_/U3  ( .A(\ADD_/FAINST[61].FA_/n1 ), .B(
        \ADD_/FAINST[61].FA_/n2 ), .Z(\ADD_/FAINST[61].FA_/n3 ) );
  XOR \ADD_/FAINST[61].FA_/U2  ( .A(b[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n2 ) );
  XOR \ADD_/FAINST[61].FA_/U1  ( .A(a[61]), .B(\ADD_/c[61] ), .Z(
        \ADD_/FAINST[61].FA_/n1 ) );
  XOR \ADD_/FAINST[60].FA_/U5  ( .A(\ADD_/FAINST[60].FA_/n3 ), .B(\ADD_/c[60] ), .Z(\ADD_/c[61] ) );
  XOR \ADD_/FAINST[60].FA_/U4  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(b[60]), .Z(
        c[60]) );
  AND \ADD_/FAINST[60].FA_/U3  ( .A(\ADD_/FAINST[60].FA_/n1 ), .B(
        \ADD_/FAINST[60].FA_/n2 ), .Z(\ADD_/FAINST[60].FA_/n3 ) );
  XOR \ADD_/FAINST[60].FA_/U2  ( .A(b[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n2 ) );
  XOR \ADD_/FAINST[60].FA_/U1  ( .A(a[60]), .B(\ADD_/c[60] ), .Z(
        \ADD_/FAINST[60].FA_/n1 ) );
  XOR \ADD_/FAINST[59].FA_/U5  ( .A(\ADD_/FAINST[59].FA_/n3 ), .B(\ADD_/c[59] ), .Z(\ADD_/c[60] ) );
  XOR \ADD_/FAINST[59].FA_/U4  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(b[59]), .Z(
        c[59]) );
  AND \ADD_/FAINST[59].FA_/U3  ( .A(\ADD_/FAINST[59].FA_/n1 ), .B(
        \ADD_/FAINST[59].FA_/n2 ), .Z(\ADD_/FAINST[59].FA_/n3 ) );
  XOR \ADD_/FAINST[59].FA_/U2  ( .A(b[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n2 ) );
  XOR \ADD_/FAINST[59].FA_/U1  ( .A(a[59]), .B(\ADD_/c[59] ), .Z(
        \ADD_/FAINST[59].FA_/n1 ) );
  XOR \ADD_/FAINST[58].FA_/U5  ( .A(\ADD_/FAINST[58].FA_/n3 ), .B(\ADD_/c[58] ), .Z(\ADD_/c[59] ) );
  XOR \ADD_/FAINST[58].FA_/U4  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(b[58]), .Z(
        c[58]) );
  AND \ADD_/FAINST[58].FA_/U3  ( .A(\ADD_/FAINST[58].FA_/n1 ), .B(
        \ADD_/FAINST[58].FA_/n2 ), .Z(\ADD_/FAINST[58].FA_/n3 ) );
  XOR \ADD_/FAINST[58].FA_/U2  ( .A(b[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n2 ) );
  XOR \ADD_/FAINST[58].FA_/U1  ( .A(a[58]), .B(\ADD_/c[58] ), .Z(
        \ADD_/FAINST[58].FA_/n1 ) );
  XOR \ADD_/FAINST[57].FA_/U5  ( .A(\ADD_/FAINST[57].FA_/n3 ), .B(\ADD_/c[57] ), .Z(\ADD_/c[58] ) );
  XOR \ADD_/FAINST[57].FA_/U4  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(b[57]), .Z(
        c[57]) );
  AND \ADD_/FAINST[57].FA_/U3  ( .A(\ADD_/FAINST[57].FA_/n1 ), .B(
        \ADD_/FAINST[57].FA_/n2 ), .Z(\ADD_/FAINST[57].FA_/n3 ) );
  XOR \ADD_/FAINST[57].FA_/U2  ( .A(b[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n2 ) );
  XOR \ADD_/FAINST[57].FA_/U1  ( .A(a[57]), .B(\ADD_/c[57] ), .Z(
        \ADD_/FAINST[57].FA_/n1 ) );
  XOR \ADD_/FAINST[56].FA_/U5  ( .A(\ADD_/FAINST[56].FA_/n3 ), .B(\ADD_/c[56] ), .Z(\ADD_/c[57] ) );
  XOR \ADD_/FAINST[56].FA_/U4  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(b[56]), .Z(
        c[56]) );
  AND \ADD_/FAINST[56].FA_/U3  ( .A(\ADD_/FAINST[56].FA_/n1 ), .B(
        \ADD_/FAINST[56].FA_/n2 ), .Z(\ADD_/FAINST[56].FA_/n3 ) );
  XOR \ADD_/FAINST[56].FA_/U2  ( .A(b[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n2 ) );
  XOR \ADD_/FAINST[56].FA_/U1  ( .A(a[56]), .B(\ADD_/c[56] ), .Z(
        \ADD_/FAINST[56].FA_/n1 ) );
  XOR \ADD_/FAINST[55].FA_/U5  ( .A(\ADD_/FAINST[55].FA_/n3 ), .B(\ADD_/c[55] ), .Z(\ADD_/c[56] ) );
  XOR \ADD_/FAINST[55].FA_/U4  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(b[55]), .Z(
        c[55]) );
  AND \ADD_/FAINST[55].FA_/U3  ( .A(\ADD_/FAINST[55].FA_/n1 ), .B(
        \ADD_/FAINST[55].FA_/n2 ), .Z(\ADD_/FAINST[55].FA_/n3 ) );
  XOR \ADD_/FAINST[55].FA_/U2  ( .A(b[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n2 ) );
  XOR \ADD_/FAINST[55].FA_/U1  ( .A(a[55]), .B(\ADD_/c[55] ), .Z(
        \ADD_/FAINST[55].FA_/n1 ) );
  XOR \ADD_/FAINST[54].FA_/U5  ( .A(\ADD_/FAINST[54].FA_/n3 ), .B(\ADD_/c[54] ), .Z(\ADD_/c[55] ) );
  XOR \ADD_/FAINST[54].FA_/U4  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(b[54]), .Z(
        c[54]) );
  AND \ADD_/FAINST[54].FA_/U3  ( .A(\ADD_/FAINST[54].FA_/n1 ), .B(
        \ADD_/FAINST[54].FA_/n2 ), .Z(\ADD_/FAINST[54].FA_/n3 ) );
  XOR \ADD_/FAINST[54].FA_/U2  ( .A(b[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n2 ) );
  XOR \ADD_/FAINST[54].FA_/U1  ( .A(a[54]), .B(\ADD_/c[54] ), .Z(
        \ADD_/FAINST[54].FA_/n1 ) );
  XOR \ADD_/FAINST[53].FA_/U5  ( .A(\ADD_/FAINST[53].FA_/n3 ), .B(\ADD_/c[53] ), .Z(\ADD_/c[54] ) );
  XOR \ADD_/FAINST[53].FA_/U4  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(b[53]), .Z(
        c[53]) );
  AND \ADD_/FAINST[53].FA_/U3  ( .A(\ADD_/FAINST[53].FA_/n1 ), .B(
        \ADD_/FAINST[53].FA_/n2 ), .Z(\ADD_/FAINST[53].FA_/n3 ) );
  XOR \ADD_/FAINST[53].FA_/U2  ( .A(b[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n2 ) );
  XOR \ADD_/FAINST[53].FA_/U1  ( .A(a[53]), .B(\ADD_/c[53] ), .Z(
        \ADD_/FAINST[53].FA_/n1 ) );
  XOR \ADD_/FAINST[52].FA_/U5  ( .A(\ADD_/FAINST[52].FA_/n3 ), .B(\ADD_/c[52] ), .Z(\ADD_/c[53] ) );
  XOR \ADD_/FAINST[52].FA_/U4  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(b[52]), .Z(
        c[52]) );
  AND \ADD_/FAINST[52].FA_/U3  ( .A(\ADD_/FAINST[52].FA_/n1 ), .B(
        \ADD_/FAINST[52].FA_/n2 ), .Z(\ADD_/FAINST[52].FA_/n3 ) );
  XOR \ADD_/FAINST[52].FA_/U2  ( .A(b[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n2 ) );
  XOR \ADD_/FAINST[52].FA_/U1  ( .A(a[52]), .B(\ADD_/c[52] ), .Z(
        \ADD_/FAINST[52].FA_/n1 ) );
  XOR \ADD_/FAINST[51].FA_/U5  ( .A(\ADD_/FAINST[51].FA_/n3 ), .B(\ADD_/c[51] ), .Z(\ADD_/c[52] ) );
  XOR \ADD_/FAINST[51].FA_/U4  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(b[51]), .Z(
        c[51]) );
  AND \ADD_/FAINST[51].FA_/U3  ( .A(\ADD_/FAINST[51].FA_/n1 ), .B(
        \ADD_/FAINST[51].FA_/n2 ), .Z(\ADD_/FAINST[51].FA_/n3 ) );
  XOR \ADD_/FAINST[51].FA_/U2  ( .A(b[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n2 ) );
  XOR \ADD_/FAINST[51].FA_/U1  ( .A(a[51]), .B(\ADD_/c[51] ), .Z(
        \ADD_/FAINST[51].FA_/n1 ) );
  XOR \ADD_/FAINST[50].FA_/U5  ( .A(\ADD_/FAINST[50].FA_/n3 ), .B(\ADD_/c[50] ), .Z(\ADD_/c[51] ) );
  XOR \ADD_/FAINST[50].FA_/U4  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(b[50]), .Z(
        c[50]) );
  AND \ADD_/FAINST[50].FA_/U3  ( .A(\ADD_/FAINST[50].FA_/n1 ), .B(
        \ADD_/FAINST[50].FA_/n2 ), .Z(\ADD_/FAINST[50].FA_/n3 ) );
  XOR \ADD_/FAINST[50].FA_/U2  ( .A(b[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n2 ) );
  XOR \ADD_/FAINST[50].FA_/U1  ( .A(a[50]), .B(\ADD_/c[50] ), .Z(
        \ADD_/FAINST[50].FA_/n1 ) );
  XOR \ADD_/FAINST[49].FA_/U5  ( .A(\ADD_/FAINST[49].FA_/n3 ), .B(\ADD_/c[49] ), .Z(\ADD_/c[50] ) );
  XOR \ADD_/FAINST[49].FA_/U4  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(b[49]), .Z(
        c[49]) );
  AND \ADD_/FAINST[49].FA_/U3  ( .A(\ADD_/FAINST[49].FA_/n1 ), .B(
        \ADD_/FAINST[49].FA_/n2 ), .Z(\ADD_/FAINST[49].FA_/n3 ) );
  XOR \ADD_/FAINST[49].FA_/U2  ( .A(b[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n2 ) );
  XOR \ADD_/FAINST[49].FA_/U1  ( .A(a[49]), .B(\ADD_/c[49] ), .Z(
        \ADD_/FAINST[49].FA_/n1 ) );
  XOR \ADD_/FAINST[48].FA_/U5  ( .A(\ADD_/FAINST[48].FA_/n3 ), .B(\ADD_/c[48] ), .Z(\ADD_/c[49] ) );
  XOR \ADD_/FAINST[48].FA_/U4  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(b[48]), .Z(
        c[48]) );
  AND \ADD_/FAINST[48].FA_/U3  ( .A(\ADD_/FAINST[48].FA_/n1 ), .B(
        \ADD_/FAINST[48].FA_/n2 ), .Z(\ADD_/FAINST[48].FA_/n3 ) );
  XOR \ADD_/FAINST[48].FA_/U2  ( .A(b[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n2 ) );
  XOR \ADD_/FAINST[48].FA_/U1  ( .A(a[48]), .B(\ADD_/c[48] ), .Z(
        \ADD_/FAINST[48].FA_/n1 ) );
  XOR \ADD_/FAINST[47].FA_/U5  ( .A(\ADD_/FAINST[47].FA_/n3 ), .B(\ADD_/c[47] ), .Z(\ADD_/c[48] ) );
  XOR \ADD_/FAINST[47].FA_/U4  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(b[47]), .Z(
        c[47]) );
  AND \ADD_/FAINST[47].FA_/U3  ( .A(\ADD_/FAINST[47].FA_/n1 ), .B(
        \ADD_/FAINST[47].FA_/n2 ), .Z(\ADD_/FAINST[47].FA_/n3 ) );
  XOR \ADD_/FAINST[47].FA_/U2  ( .A(b[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n2 ) );
  XOR \ADD_/FAINST[47].FA_/U1  ( .A(a[47]), .B(\ADD_/c[47] ), .Z(
        \ADD_/FAINST[47].FA_/n1 ) );
  XOR \ADD_/FAINST[46].FA_/U5  ( .A(\ADD_/FAINST[46].FA_/n3 ), .B(\ADD_/c[46] ), .Z(\ADD_/c[47] ) );
  XOR \ADD_/FAINST[46].FA_/U4  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(b[46]), .Z(
        c[46]) );
  AND \ADD_/FAINST[46].FA_/U3  ( .A(\ADD_/FAINST[46].FA_/n1 ), .B(
        \ADD_/FAINST[46].FA_/n2 ), .Z(\ADD_/FAINST[46].FA_/n3 ) );
  XOR \ADD_/FAINST[46].FA_/U2  ( .A(b[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n2 ) );
  XOR \ADD_/FAINST[46].FA_/U1  ( .A(a[46]), .B(\ADD_/c[46] ), .Z(
        \ADD_/FAINST[46].FA_/n1 ) );
  XOR \ADD_/FAINST[45].FA_/U5  ( .A(\ADD_/FAINST[45].FA_/n3 ), .B(\ADD_/c[45] ), .Z(\ADD_/c[46] ) );
  XOR \ADD_/FAINST[45].FA_/U4  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(b[45]), .Z(
        c[45]) );
  AND \ADD_/FAINST[45].FA_/U3  ( .A(\ADD_/FAINST[45].FA_/n1 ), .B(
        \ADD_/FAINST[45].FA_/n2 ), .Z(\ADD_/FAINST[45].FA_/n3 ) );
  XOR \ADD_/FAINST[45].FA_/U2  ( .A(b[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n2 ) );
  XOR \ADD_/FAINST[45].FA_/U1  ( .A(a[45]), .B(\ADD_/c[45] ), .Z(
        \ADD_/FAINST[45].FA_/n1 ) );
  XOR \ADD_/FAINST[44].FA_/U5  ( .A(\ADD_/FAINST[44].FA_/n3 ), .B(\ADD_/c[44] ), .Z(\ADD_/c[45] ) );
  XOR \ADD_/FAINST[44].FA_/U4  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(b[44]), .Z(
        c[44]) );
  AND \ADD_/FAINST[44].FA_/U3  ( .A(\ADD_/FAINST[44].FA_/n1 ), .B(
        \ADD_/FAINST[44].FA_/n2 ), .Z(\ADD_/FAINST[44].FA_/n3 ) );
  XOR \ADD_/FAINST[44].FA_/U2  ( .A(b[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n2 ) );
  XOR \ADD_/FAINST[44].FA_/U1  ( .A(a[44]), .B(\ADD_/c[44] ), .Z(
        \ADD_/FAINST[44].FA_/n1 ) );
  XOR \ADD_/FAINST[43].FA_/U5  ( .A(\ADD_/FAINST[43].FA_/n3 ), .B(\ADD_/c[43] ), .Z(\ADD_/c[44] ) );
  XOR \ADD_/FAINST[43].FA_/U4  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(b[43]), .Z(
        c[43]) );
  AND \ADD_/FAINST[43].FA_/U3  ( .A(\ADD_/FAINST[43].FA_/n1 ), .B(
        \ADD_/FAINST[43].FA_/n2 ), .Z(\ADD_/FAINST[43].FA_/n3 ) );
  XOR \ADD_/FAINST[43].FA_/U2  ( .A(b[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n2 ) );
  XOR \ADD_/FAINST[43].FA_/U1  ( .A(a[43]), .B(\ADD_/c[43] ), .Z(
        \ADD_/FAINST[43].FA_/n1 ) );
  XOR \ADD_/FAINST[42].FA_/U5  ( .A(\ADD_/FAINST[42].FA_/n3 ), .B(\ADD_/c[42] ), .Z(\ADD_/c[43] ) );
  XOR \ADD_/FAINST[42].FA_/U4  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(b[42]), .Z(
        c[42]) );
  AND \ADD_/FAINST[42].FA_/U3  ( .A(\ADD_/FAINST[42].FA_/n1 ), .B(
        \ADD_/FAINST[42].FA_/n2 ), .Z(\ADD_/FAINST[42].FA_/n3 ) );
  XOR \ADD_/FAINST[42].FA_/U2  ( .A(b[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n2 ) );
  XOR \ADD_/FAINST[42].FA_/U1  ( .A(a[42]), .B(\ADD_/c[42] ), .Z(
        \ADD_/FAINST[42].FA_/n1 ) );
  XOR \ADD_/FAINST[41].FA_/U5  ( .A(\ADD_/FAINST[41].FA_/n3 ), .B(\ADD_/c[41] ), .Z(\ADD_/c[42] ) );
  XOR \ADD_/FAINST[41].FA_/U4  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(b[41]), .Z(
        c[41]) );
  AND \ADD_/FAINST[41].FA_/U3  ( .A(\ADD_/FAINST[41].FA_/n1 ), .B(
        \ADD_/FAINST[41].FA_/n2 ), .Z(\ADD_/FAINST[41].FA_/n3 ) );
  XOR \ADD_/FAINST[41].FA_/U2  ( .A(b[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n2 ) );
  XOR \ADD_/FAINST[41].FA_/U1  ( .A(a[41]), .B(\ADD_/c[41] ), .Z(
        \ADD_/FAINST[41].FA_/n1 ) );
  XOR \ADD_/FAINST[40].FA_/U5  ( .A(\ADD_/FAINST[40].FA_/n3 ), .B(\ADD_/c[40] ), .Z(\ADD_/c[41] ) );
  XOR \ADD_/FAINST[40].FA_/U4  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(b[40]), .Z(
        c[40]) );
  AND \ADD_/FAINST[40].FA_/U3  ( .A(\ADD_/FAINST[40].FA_/n1 ), .B(
        \ADD_/FAINST[40].FA_/n2 ), .Z(\ADD_/FAINST[40].FA_/n3 ) );
  XOR \ADD_/FAINST[40].FA_/U2  ( .A(b[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n2 ) );
  XOR \ADD_/FAINST[40].FA_/U1  ( .A(a[40]), .B(\ADD_/c[40] ), .Z(
        \ADD_/FAINST[40].FA_/n1 ) );
  XOR \ADD_/FAINST[39].FA_/U5  ( .A(\ADD_/FAINST[39].FA_/n3 ), .B(\ADD_/c[39] ), .Z(\ADD_/c[40] ) );
  XOR \ADD_/FAINST[39].FA_/U4  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(b[39]), .Z(
        c[39]) );
  AND \ADD_/FAINST[39].FA_/U3  ( .A(\ADD_/FAINST[39].FA_/n1 ), .B(
        \ADD_/FAINST[39].FA_/n2 ), .Z(\ADD_/FAINST[39].FA_/n3 ) );
  XOR \ADD_/FAINST[39].FA_/U2  ( .A(b[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n2 ) );
  XOR \ADD_/FAINST[39].FA_/U1  ( .A(a[39]), .B(\ADD_/c[39] ), .Z(
        \ADD_/FAINST[39].FA_/n1 ) );
  XOR \ADD_/FAINST[38].FA_/U5  ( .A(\ADD_/FAINST[38].FA_/n3 ), .B(\ADD_/c[38] ), .Z(\ADD_/c[39] ) );
  XOR \ADD_/FAINST[38].FA_/U4  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(b[38]), .Z(
        c[38]) );
  AND \ADD_/FAINST[38].FA_/U3  ( .A(\ADD_/FAINST[38].FA_/n1 ), .B(
        \ADD_/FAINST[38].FA_/n2 ), .Z(\ADD_/FAINST[38].FA_/n3 ) );
  XOR \ADD_/FAINST[38].FA_/U2  ( .A(b[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n2 ) );
  XOR \ADD_/FAINST[38].FA_/U1  ( .A(a[38]), .B(\ADD_/c[38] ), .Z(
        \ADD_/FAINST[38].FA_/n1 ) );
  XOR \ADD_/FAINST[37].FA_/U5  ( .A(\ADD_/FAINST[37].FA_/n3 ), .B(\ADD_/c[37] ), .Z(\ADD_/c[38] ) );
  XOR \ADD_/FAINST[37].FA_/U4  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(b[37]), .Z(
        c[37]) );
  AND \ADD_/FAINST[37].FA_/U3  ( .A(\ADD_/FAINST[37].FA_/n1 ), .B(
        \ADD_/FAINST[37].FA_/n2 ), .Z(\ADD_/FAINST[37].FA_/n3 ) );
  XOR \ADD_/FAINST[37].FA_/U2  ( .A(b[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n2 ) );
  XOR \ADD_/FAINST[37].FA_/U1  ( .A(a[37]), .B(\ADD_/c[37] ), .Z(
        \ADD_/FAINST[37].FA_/n1 ) );
  XOR \ADD_/FAINST[36].FA_/U5  ( .A(\ADD_/FAINST[36].FA_/n3 ), .B(\ADD_/c[36] ), .Z(\ADD_/c[37] ) );
  XOR \ADD_/FAINST[36].FA_/U4  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(b[36]), .Z(
        c[36]) );
  AND \ADD_/FAINST[36].FA_/U3  ( .A(\ADD_/FAINST[36].FA_/n1 ), .B(
        \ADD_/FAINST[36].FA_/n2 ), .Z(\ADD_/FAINST[36].FA_/n3 ) );
  XOR \ADD_/FAINST[36].FA_/U2  ( .A(b[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n2 ) );
  XOR \ADD_/FAINST[36].FA_/U1  ( .A(a[36]), .B(\ADD_/c[36] ), .Z(
        \ADD_/FAINST[36].FA_/n1 ) );
  XOR \ADD_/FAINST[35].FA_/U5  ( .A(\ADD_/FAINST[35].FA_/n3 ), .B(\ADD_/c[35] ), .Z(\ADD_/c[36] ) );
  XOR \ADD_/FAINST[35].FA_/U4  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(b[35]), .Z(
        c[35]) );
  AND \ADD_/FAINST[35].FA_/U3  ( .A(\ADD_/FAINST[35].FA_/n1 ), .B(
        \ADD_/FAINST[35].FA_/n2 ), .Z(\ADD_/FAINST[35].FA_/n3 ) );
  XOR \ADD_/FAINST[35].FA_/U2  ( .A(b[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n2 ) );
  XOR \ADD_/FAINST[35].FA_/U1  ( .A(a[35]), .B(\ADD_/c[35] ), .Z(
        \ADD_/FAINST[35].FA_/n1 ) );
  XOR \ADD_/FAINST[34].FA_/U5  ( .A(\ADD_/FAINST[34].FA_/n3 ), .B(\ADD_/c[34] ), .Z(\ADD_/c[35] ) );
  XOR \ADD_/FAINST[34].FA_/U4  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(b[34]), .Z(
        c[34]) );
  AND \ADD_/FAINST[34].FA_/U3  ( .A(\ADD_/FAINST[34].FA_/n1 ), .B(
        \ADD_/FAINST[34].FA_/n2 ), .Z(\ADD_/FAINST[34].FA_/n3 ) );
  XOR \ADD_/FAINST[34].FA_/U2  ( .A(b[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n2 ) );
  XOR \ADD_/FAINST[34].FA_/U1  ( .A(a[34]), .B(\ADD_/c[34] ), .Z(
        \ADD_/FAINST[34].FA_/n1 ) );
  XOR \ADD_/FAINST[33].FA_/U5  ( .A(\ADD_/FAINST[33].FA_/n3 ), .B(\ADD_/c[33] ), .Z(\ADD_/c[34] ) );
  XOR \ADD_/FAINST[33].FA_/U4  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(b[33]), .Z(
        c[33]) );
  AND \ADD_/FAINST[33].FA_/U3  ( .A(\ADD_/FAINST[33].FA_/n1 ), .B(
        \ADD_/FAINST[33].FA_/n2 ), .Z(\ADD_/FAINST[33].FA_/n3 ) );
  XOR \ADD_/FAINST[33].FA_/U2  ( .A(b[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n2 ) );
  XOR \ADD_/FAINST[33].FA_/U1  ( .A(a[33]), .B(\ADD_/c[33] ), .Z(
        \ADD_/FAINST[33].FA_/n1 ) );
  XOR \ADD_/FAINST[32].FA_/U5  ( .A(\ADD_/FAINST[32].FA_/n3 ), .B(\ADD_/c[32] ), .Z(\ADD_/c[33] ) );
  XOR \ADD_/FAINST[32].FA_/U4  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(b[32]), .Z(
        c[32]) );
  AND \ADD_/FAINST[32].FA_/U3  ( .A(\ADD_/FAINST[32].FA_/n1 ), .B(
        \ADD_/FAINST[32].FA_/n2 ), .Z(\ADD_/FAINST[32].FA_/n3 ) );
  XOR \ADD_/FAINST[32].FA_/U2  ( .A(b[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n2 ) );
  XOR \ADD_/FAINST[32].FA_/U1  ( .A(a[32]), .B(\ADD_/c[32] ), .Z(
        \ADD_/FAINST[32].FA_/n1 ) );
  XOR \ADD_/FAINST[31].FA_/U5  ( .A(\ADD_/FAINST[31].FA_/n3 ), .B(\ADD_/c[31] ), .Z(\ADD_/c[32] ) );
  XOR \ADD_/FAINST[31].FA_/U4  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(b[31]), .Z(
        c[31]) );
  AND \ADD_/FAINST[31].FA_/U3  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(
        \ADD_/FAINST[31].FA_/n2 ), .Z(\ADD_/FAINST[31].FA_/n3 ) );
  XOR \ADD_/FAINST[31].FA_/U2  ( .A(b[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n2 ) );
  XOR \ADD_/FAINST[31].FA_/U1  ( .A(a[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n1 ) );
  XOR \ADD_/FAINST[30].FA_/U5  ( .A(\ADD_/FAINST[30].FA_/n3 ), .B(\ADD_/c[30] ), .Z(\ADD_/c[31] ) );
  XOR \ADD_/FAINST[30].FA_/U4  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(b[30]), .Z(
        c[30]) );
  AND \ADD_/FAINST[30].FA_/U3  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(
        \ADD_/FAINST[30].FA_/n2 ), .Z(\ADD_/FAINST[30].FA_/n3 ) );
  XOR \ADD_/FAINST[30].FA_/U2  ( .A(b[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n2 ) );
  XOR \ADD_/FAINST[30].FA_/U1  ( .A(a[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n1 ) );
  XOR \ADD_/FAINST[29].FA_/U5  ( .A(\ADD_/FAINST[29].FA_/n3 ), .B(\ADD_/c[29] ), .Z(\ADD_/c[30] ) );
  XOR \ADD_/FAINST[29].FA_/U4  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(b[29]), .Z(
        c[29]) );
  AND \ADD_/FAINST[29].FA_/U3  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(
        \ADD_/FAINST[29].FA_/n2 ), .Z(\ADD_/FAINST[29].FA_/n3 ) );
  XOR \ADD_/FAINST[29].FA_/U2  ( .A(b[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n2 ) );
  XOR \ADD_/FAINST[29].FA_/U1  ( .A(a[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n1 ) );
  XOR \ADD_/FAINST[28].FA_/U5  ( .A(\ADD_/FAINST[28].FA_/n3 ), .B(\ADD_/c[28] ), .Z(\ADD_/c[29] ) );
  XOR \ADD_/FAINST[28].FA_/U4  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(b[28]), .Z(
        c[28]) );
  AND \ADD_/FAINST[28].FA_/U3  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(
        \ADD_/FAINST[28].FA_/n2 ), .Z(\ADD_/FAINST[28].FA_/n3 ) );
  XOR \ADD_/FAINST[28].FA_/U2  ( .A(b[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n2 ) );
  XOR \ADD_/FAINST[28].FA_/U1  ( .A(a[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n1 ) );
  XOR \ADD_/FAINST[27].FA_/U5  ( .A(\ADD_/FAINST[27].FA_/n3 ), .B(\ADD_/c[27] ), .Z(\ADD_/c[28] ) );
  XOR \ADD_/FAINST[27].FA_/U4  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(b[27]), .Z(
        c[27]) );
  AND \ADD_/FAINST[27].FA_/U3  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(
        \ADD_/FAINST[27].FA_/n2 ), .Z(\ADD_/FAINST[27].FA_/n3 ) );
  XOR \ADD_/FAINST[27].FA_/U2  ( .A(b[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n2 ) );
  XOR \ADD_/FAINST[27].FA_/U1  ( .A(a[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n1 ) );
  XOR \ADD_/FAINST[26].FA_/U5  ( .A(\ADD_/FAINST[26].FA_/n3 ), .B(\ADD_/c[26] ), .Z(\ADD_/c[27] ) );
  XOR \ADD_/FAINST[26].FA_/U4  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(b[26]), .Z(
        c[26]) );
  AND \ADD_/FAINST[26].FA_/U3  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(
        \ADD_/FAINST[26].FA_/n2 ), .Z(\ADD_/FAINST[26].FA_/n3 ) );
  XOR \ADD_/FAINST[26].FA_/U2  ( .A(b[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n2 ) );
  XOR \ADD_/FAINST[26].FA_/U1  ( .A(a[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n1 ) );
  XOR \ADD_/FAINST[25].FA_/U5  ( .A(\ADD_/FAINST[25].FA_/n3 ), .B(\ADD_/c[25] ), .Z(\ADD_/c[26] ) );
  XOR \ADD_/FAINST[25].FA_/U4  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(b[25]), .Z(
        c[25]) );
  AND \ADD_/FAINST[25].FA_/U3  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(
        \ADD_/FAINST[25].FA_/n2 ), .Z(\ADD_/FAINST[25].FA_/n3 ) );
  XOR \ADD_/FAINST[25].FA_/U2  ( .A(b[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n2 ) );
  XOR \ADD_/FAINST[25].FA_/U1  ( .A(a[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n1 ) );
  XOR \ADD_/FAINST[24].FA_/U5  ( .A(\ADD_/FAINST[24].FA_/n3 ), .B(\ADD_/c[24] ), .Z(\ADD_/c[25] ) );
  XOR \ADD_/FAINST[24].FA_/U4  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(b[24]), .Z(
        c[24]) );
  AND \ADD_/FAINST[24].FA_/U3  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(
        \ADD_/FAINST[24].FA_/n2 ), .Z(\ADD_/FAINST[24].FA_/n3 ) );
  XOR \ADD_/FAINST[24].FA_/U2  ( .A(b[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n2 ) );
  XOR \ADD_/FAINST[24].FA_/U1  ( .A(a[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n1 ) );
  XOR \ADD_/FAINST[23].FA_/U5  ( .A(\ADD_/FAINST[23].FA_/n3 ), .B(\ADD_/c[23] ), .Z(\ADD_/c[24] ) );
  XOR \ADD_/FAINST[23].FA_/U4  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(b[23]), .Z(
        c[23]) );
  AND \ADD_/FAINST[23].FA_/U3  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(
        \ADD_/FAINST[23].FA_/n2 ), .Z(\ADD_/FAINST[23].FA_/n3 ) );
  XOR \ADD_/FAINST[23].FA_/U2  ( .A(b[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n2 ) );
  XOR \ADD_/FAINST[23].FA_/U1  ( .A(a[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n1 ) );
  XOR \ADD_/FAINST[22].FA_/U5  ( .A(\ADD_/FAINST[22].FA_/n3 ), .B(\ADD_/c[22] ), .Z(\ADD_/c[23] ) );
  XOR \ADD_/FAINST[22].FA_/U4  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(b[22]), .Z(
        c[22]) );
  AND \ADD_/FAINST[22].FA_/U3  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(
        \ADD_/FAINST[22].FA_/n2 ), .Z(\ADD_/FAINST[22].FA_/n3 ) );
  XOR \ADD_/FAINST[22].FA_/U2  ( .A(b[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n2 ) );
  XOR \ADD_/FAINST[22].FA_/U1  ( .A(a[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n1 ) );
  XOR \ADD_/FAINST[21].FA_/U5  ( .A(\ADD_/FAINST[21].FA_/n3 ), .B(\ADD_/c[21] ), .Z(\ADD_/c[22] ) );
  XOR \ADD_/FAINST[21].FA_/U4  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(b[21]), .Z(
        c[21]) );
  AND \ADD_/FAINST[21].FA_/U3  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(
        \ADD_/FAINST[21].FA_/n2 ), .Z(\ADD_/FAINST[21].FA_/n3 ) );
  XOR \ADD_/FAINST[21].FA_/U2  ( .A(b[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n2 ) );
  XOR \ADD_/FAINST[21].FA_/U1  ( .A(a[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n1 ) );
  XOR \ADD_/FAINST[20].FA_/U5  ( .A(\ADD_/FAINST[20].FA_/n3 ), .B(\ADD_/c[20] ), .Z(\ADD_/c[21] ) );
  XOR \ADD_/FAINST[20].FA_/U4  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(b[20]), .Z(
        c[20]) );
  AND \ADD_/FAINST[20].FA_/U3  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(
        \ADD_/FAINST[20].FA_/n2 ), .Z(\ADD_/FAINST[20].FA_/n3 ) );
  XOR \ADD_/FAINST[20].FA_/U2  ( .A(b[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n2 ) );
  XOR \ADD_/FAINST[20].FA_/U1  ( .A(a[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n1 ) );
  XOR \ADD_/FAINST[19].FA_/U5  ( .A(\ADD_/FAINST[19].FA_/n3 ), .B(\ADD_/c[19] ), .Z(\ADD_/c[20] ) );
  XOR \ADD_/FAINST[19].FA_/U4  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(b[19]), .Z(
        c[19]) );
  AND \ADD_/FAINST[19].FA_/U3  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(
        \ADD_/FAINST[19].FA_/n2 ), .Z(\ADD_/FAINST[19].FA_/n3 ) );
  XOR \ADD_/FAINST[19].FA_/U2  ( .A(b[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n2 ) );
  XOR \ADD_/FAINST[19].FA_/U1  ( .A(a[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n1 ) );
  XOR \ADD_/FAINST[18].FA_/U5  ( .A(\ADD_/FAINST[18].FA_/n3 ), .B(\ADD_/c[18] ), .Z(\ADD_/c[19] ) );
  XOR \ADD_/FAINST[18].FA_/U4  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(b[18]), .Z(
        c[18]) );
  AND \ADD_/FAINST[18].FA_/U3  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(
        \ADD_/FAINST[18].FA_/n2 ), .Z(\ADD_/FAINST[18].FA_/n3 ) );
  XOR \ADD_/FAINST[18].FA_/U2  ( .A(b[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n2 ) );
  XOR \ADD_/FAINST[18].FA_/U1  ( .A(a[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n1 ) );
  XOR \ADD_/FAINST[17].FA_/U5  ( .A(\ADD_/FAINST[17].FA_/n3 ), .B(\ADD_/c[17] ), .Z(\ADD_/c[18] ) );
  XOR \ADD_/FAINST[17].FA_/U4  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(b[17]), .Z(
        c[17]) );
  AND \ADD_/FAINST[17].FA_/U3  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(
        \ADD_/FAINST[17].FA_/n2 ), .Z(\ADD_/FAINST[17].FA_/n3 ) );
  XOR \ADD_/FAINST[17].FA_/U2  ( .A(b[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n2 ) );
  XOR \ADD_/FAINST[17].FA_/U1  ( .A(a[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n1 ) );
  XOR \ADD_/FAINST[16].FA_/U5  ( .A(\ADD_/FAINST[16].FA_/n3 ), .B(\ADD_/c[16] ), .Z(\ADD_/c[17] ) );
  XOR \ADD_/FAINST[16].FA_/U4  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(b[16]), .Z(
        c[16]) );
  AND \ADD_/FAINST[16].FA_/U3  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(
        \ADD_/FAINST[16].FA_/n2 ), .Z(\ADD_/FAINST[16].FA_/n3 ) );
  XOR \ADD_/FAINST[16].FA_/U2  ( .A(b[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n2 ) );
  XOR \ADD_/FAINST[16].FA_/U1  ( .A(a[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n1 ) );
  XOR \ADD_/FAINST[15].FA_/U5  ( .A(\ADD_/FAINST[15].FA_/n3 ), .B(\ADD_/c[15] ), .Z(\ADD_/c[16] ) );
  XOR \ADD_/FAINST[15].FA_/U4  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(b[15]), .Z(
        c[15]) );
  AND \ADD_/FAINST[15].FA_/U3  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(
        \ADD_/FAINST[15].FA_/n2 ), .Z(\ADD_/FAINST[15].FA_/n3 ) );
  XOR \ADD_/FAINST[15].FA_/U2  ( .A(b[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n2 ) );
  XOR \ADD_/FAINST[15].FA_/U1  ( .A(a[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n1 ) );
  XOR \ADD_/FAINST[14].FA_/U5  ( .A(\ADD_/FAINST[14].FA_/n3 ), .B(\ADD_/c[14] ), .Z(\ADD_/c[15] ) );
  XOR \ADD_/FAINST[14].FA_/U4  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(b[14]), .Z(
        c[14]) );
  AND \ADD_/FAINST[14].FA_/U3  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(
        \ADD_/FAINST[14].FA_/n2 ), .Z(\ADD_/FAINST[14].FA_/n3 ) );
  XOR \ADD_/FAINST[14].FA_/U2  ( .A(b[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n2 ) );
  XOR \ADD_/FAINST[14].FA_/U1  ( .A(a[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n1 ) );
  XOR \ADD_/FAINST[13].FA_/U5  ( .A(\ADD_/FAINST[13].FA_/n3 ), .B(\ADD_/c[13] ), .Z(\ADD_/c[14] ) );
  XOR \ADD_/FAINST[13].FA_/U4  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(b[13]), .Z(
        c[13]) );
  AND \ADD_/FAINST[13].FA_/U3  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(
        \ADD_/FAINST[13].FA_/n2 ), .Z(\ADD_/FAINST[13].FA_/n3 ) );
  XOR \ADD_/FAINST[13].FA_/U2  ( .A(b[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n2 ) );
  XOR \ADD_/FAINST[13].FA_/U1  ( .A(a[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n1 ) );
  XOR \ADD_/FAINST[12].FA_/U5  ( .A(\ADD_/FAINST[12].FA_/n3 ), .B(\ADD_/c[12] ), .Z(\ADD_/c[13] ) );
  XOR \ADD_/FAINST[12].FA_/U4  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(b[12]), .Z(
        c[12]) );
  AND \ADD_/FAINST[12].FA_/U3  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(
        \ADD_/FAINST[12].FA_/n2 ), .Z(\ADD_/FAINST[12].FA_/n3 ) );
  XOR \ADD_/FAINST[12].FA_/U2  ( .A(b[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n2 ) );
  XOR \ADD_/FAINST[12].FA_/U1  ( .A(a[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n1 ) );
  XOR \ADD_/FAINST[11].FA_/U5  ( .A(\ADD_/FAINST[11].FA_/n3 ), .B(\ADD_/c[11] ), .Z(\ADD_/c[12] ) );
  XOR \ADD_/FAINST[11].FA_/U4  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(b[11]), .Z(
        c[11]) );
  AND \ADD_/FAINST[11].FA_/U3  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(
        \ADD_/FAINST[11].FA_/n2 ), .Z(\ADD_/FAINST[11].FA_/n3 ) );
  XOR \ADD_/FAINST[11].FA_/U2  ( .A(b[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n2 ) );
  XOR \ADD_/FAINST[11].FA_/U1  ( .A(a[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n1 ) );
  XOR \ADD_/FAINST[10].FA_/U5  ( .A(\ADD_/FAINST[10].FA_/n3 ), .B(\ADD_/c[10] ), .Z(\ADD_/c[11] ) );
  XOR \ADD_/FAINST[10].FA_/U4  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(b[10]), .Z(
        c[10]) );
  AND \ADD_/FAINST[10].FA_/U3  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(
        \ADD_/FAINST[10].FA_/n2 ), .Z(\ADD_/FAINST[10].FA_/n3 ) );
  XOR \ADD_/FAINST[10].FA_/U2  ( .A(b[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n2 ) );
  XOR \ADD_/FAINST[10].FA_/U1  ( .A(a[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n1 ) );
  XOR \ADD_/FAINST[9].FA_/U5  ( .A(\ADD_/FAINST[9].FA_/n3 ), .B(\ADD_/c[9] ), 
        .Z(\ADD_/c[10] ) );
  XOR \ADD_/FAINST[9].FA_/U4  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(b[9]), .Z(c[9]) );
  AND \ADD_/FAINST[9].FA_/U3  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(
        \ADD_/FAINST[9].FA_/n2 ), .Z(\ADD_/FAINST[9].FA_/n3 ) );
  XOR \ADD_/FAINST[9].FA_/U2  ( .A(b[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n2 ) );
  XOR \ADD_/FAINST[9].FA_/U1  ( .A(a[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n1 ) );
  XOR \ADD_/FAINST[8].FA_/U5  ( .A(\ADD_/FAINST[8].FA_/n3 ), .B(\ADD_/c[8] ), 
        .Z(\ADD_/c[9] ) );
  XOR \ADD_/FAINST[8].FA_/U4  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(b[8]), .Z(c[8]) );
  AND \ADD_/FAINST[8].FA_/U3  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(
        \ADD_/FAINST[8].FA_/n2 ), .Z(\ADD_/FAINST[8].FA_/n3 ) );
  XOR \ADD_/FAINST[8].FA_/U2  ( .A(b[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n2 ) );
  XOR \ADD_/FAINST[8].FA_/U1  ( .A(a[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n1 ) );
  XOR \ADD_/FAINST[7].FA_/U5  ( .A(\ADD_/FAINST[7].FA_/n3 ), .B(\ADD_/c[7] ), 
        .Z(\ADD_/c[8] ) );
  XOR \ADD_/FAINST[7].FA_/U4  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(b[7]), .Z(c[7]) );
  AND \ADD_/FAINST[7].FA_/U3  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(
        \ADD_/FAINST[7].FA_/n2 ), .Z(\ADD_/FAINST[7].FA_/n3 ) );
  XOR \ADD_/FAINST[7].FA_/U2  ( .A(b[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n2 ) );
  XOR \ADD_/FAINST[7].FA_/U1  ( .A(a[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n1 ) );
  XOR \ADD_/FAINST[6].FA_/U5  ( .A(\ADD_/FAINST[6].FA_/n3 ), .B(\ADD_/c[6] ), 
        .Z(\ADD_/c[7] ) );
  XOR \ADD_/FAINST[6].FA_/U4  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(b[6]), .Z(c[6]) );
  AND \ADD_/FAINST[6].FA_/U3  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(
        \ADD_/FAINST[6].FA_/n2 ), .Z(\ADD_/FAINST[6].FA_/n3 ) );
  XOR \ADD_/FAINST[6].FA_/U2  ( .A(b[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n2 ) );
  XOR \ADD_/FAINST[6].FA_/U1  ( .A(a[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n1 ) );
  XOR \ADD_/FAINST[5].FA_/U5  ( .A(\ADD_/FAINST[5].FA_/n3 ), .B(\ADD_/c[5] ), 
        .Z(\ADD_/c[6] ) );
  XOR \ADD_/FAINST[5].FA_/U4  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(b[5]), .Z(c[5]) );
  AND \ADD_/FAINST[5].FA_/U3  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(
        \ADD_/FAINST[5].FA_/n2 ), .Z(\ADD_/FAINST[5].FA_/n3 ) );
  XOR \ADD_/FAINST[5].FA_/U2  ( .A(b[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n2 ) );
  XOR \ADD_/FAINST[5].FA_/U1  ( .A(a[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n1 ) );
  XOR \ADD_/FAINST[4].FA_/U5  ( .A(\ADD_/FAINST[4].FA_/n3 ), .B(\ADD_/c[4] ), 
        .Z(\ADD_/c[5] ) );
  XOR \ADD_/FAINST[4].FA_/U4  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(b[4]), .Z(c[4]) );
  AND \ADD_/FAINST[4].FA_/U3  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(
        \ADD_/FAINST[4].FA_/n2 ), .Z(\ADD_/FAINST[4].FA_/n3 ) );
  XOR \ADD_/FAINST[4].FA_/U2  ( .A(b[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n2 ) );
  XOR \ADD_/FAINST[4].FA_/U1  ( .A(a[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n1 ) );
  XOR \ADD_/FAINST[3].FA_/U5  ( .A(\ADD_/FAINST[3].FA_/n3 ), .B(\ADD_/c[3] ), 
        .Z(\ADD_/c[4] ) );
  XOR \ADD_/FAINST[3].FA_/U4  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(b[3]), .Z(c[3]) );
  AND \ADD_/FAINST[3].FA_/U3  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(
        \ADD_/FAINST[3].FA_/n2 ), .Z(\ADD_/FAINST[3].FA_/n3 ) );
  XOR \ADD_/FAINST[3].FA_/U2  ( .A(b[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n2 ) );
  XOR \ADD_/FAINST[3].FA_/U1  ( .A(a[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n1 ) );
  XOR \ADD_/FAINST[2].FA_/U5  ( .A(\ADD_/FAINST[2].FA_/n3 ), .B(\ADD_/c[2] ), 
        .Z(\ADD_/c[3] ) );
  XOR \ADD_/FAINST[2].FA_/U4  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(b[2]), .Z(c[2]) );
  AND \ADD_/FAINST[2].FA_/U3  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(
        \ADD_/FAINST[2].FA_/n2 ), .Z(\ADD_/FAINST[2].FA_/n3 ) );
  XOR \ADD_/FAINST[2].FA_/U2  ( .A(b[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n2 ) );
  XOR \ADD_/FAINST[2].FA_/U1  ( .A(a[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n1 ) );
  XOR \ADD_/FAINST[1].FA_/U5  ( .A(\ADD_/FAINST[1].FA_/n3 ), .B(\ADD_/c[1] ), 
        .Z(\ADD_/c[2] ) );
  XOR \ADD_/FAINST[1].FA_/U4  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(b[1]), .Z(c[1]) );
  AND \ADD_/FAINST[1].FA_/U3  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(
        \ADD_/FAINST[1].FA_/n2 ), .Z(\ADD_/FAINST[1].FA_/n3 ) );
  XOR \ADD_/FAINST[1].FA_/U2  ( .A(b[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n2 ) );
  XOR \ADD_/FAINST[1].FA_/U1  ( .A(a[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n1 ) );
endmodule

