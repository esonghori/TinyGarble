
module modmult_N256_CC512 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;


endmodule


module modexp_2N_NN_N256_CC262144 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203;
  wire   [511:0] start_in;
  wire   [511:0] start_reg;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] x;
  wire   [255:0] y;

  modmult_N256_CC512 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .Q(
        start_reg[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .Q(
        start_reg[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .Q(
        start_reg[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .Q(
        start_reg[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .Q(
        start_reg[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .Q(
        start_reg[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .Q(
        start_reg[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .Q(
        start_reg[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .Q(
        start_reg[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .Q(
        start_reg[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .Q(
        start_reg[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .Q(
        start_reg[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .Q(
        start_reg[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .Q(
        start_reg[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .Q(
        start_reg[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .Q(
        start_reg[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .Q(
        start_reg[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .Q(
        start_reg[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .Q(
        start_reg[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .Q(
        start_reg[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .Q(
        start_reg[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .Q(
        start_reg[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .Q(
        start_reg[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .Q(
        start_reg[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .Q(
        start_reg[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .Q(
        start_reg[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .Q(
        start_reg[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .Q(
        start_reg[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .Q(
        start_reg[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .Q(
        start_reg[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .Q(
        start_reg[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .Q(
        start_reg[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .Q(
        start_reg[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .Q(
        start_reg[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .Q(
        start_reg[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .Q(
        start_reg[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .Q(
        start_reg[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .Q(
        start_reg[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .Q(
        start_reg[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .Q(
        start_reg[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .Q(
        start_reg[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .Q(
        start_reg[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .Q(
        start_reg[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .Q(
        start_reg[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .Q(
        start_reg[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .Q(
        start_reg[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .Q(
        start_reg[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .Q(
        start_reg[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .Q(
        start_reg[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .Q(
        start_reg[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .Q(
        start_reg[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .Q(
        start_reg[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .Q(
        start_reg[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .Q(
        start_reg[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .Q(
        start_reg[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .Q(
        start_reg[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .Q(
        start_reg[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .Q(
        start_reg[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .Q(
        start_reg[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .Q(
        start_reg[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .Q(
        start_reg[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .Q(
        start_reg[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .Q(
        start_reg[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .Q(
        start_reg[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .Q(
        start_reg[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .Q(
        start_reg[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .Q(
        start_reg[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .Q(
        start_reg[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .Q(
        start_reg[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .Q(
        start_reg[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .Q(
        start_reg[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .Q(
        start_reg[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .Q(
        start_reg[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .Q(
        start_reg[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .Q(
        start_reg[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .Q(
        start_reg[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .Q(
        start_reg[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .Q(
        start_reg[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .Q(
        start_reg[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .Q(
        start_reg[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .Q(
        start_reg[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .Q(
        start_reg[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .Q(
        start_reg[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .Q(
        start_reg[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .Q(
        start_reg[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .Q(
        start_reg[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .Q(
        start_reg[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .Q(
        start_reg[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .Q(
        start_reg[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .Q(
        start_reg[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .Q(
        start_reg[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .Q(
        start_reg[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .Q(
        start_reg[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .Q(
        start_reg[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .Q(
        start_reg[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .Q(
        start_reg[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .Q(
        start_reg[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .Q(
        start_reg[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .Q(
        start_reg[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .Q(
        start_reg[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .Q(
        start_reg[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .Q(
        start_reg[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .Q(
        start_reg[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .Q(
        start_reg[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .Q(
        start_reg[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .Q(
        start_reg[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .Q(
        start_reg[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .Q(
        start_reg[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .Q(
        start_reg[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .Q(
        start_reg[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .Q(
        start_reg[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .Q(
        start_reg[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .Q(
        start_reg[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .Q(
        start_reg[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .Q(
        start_reg[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .Q(
        start_reg[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .Q(
        start_reg[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .Q(
        start_reg[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .Q(
        start_reg[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .Q(
        start_reg[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .Q(
        start_reg[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .Q(
        start_reg[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .Q(
        start_reg[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .Q(
        start_reg[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .Q(
        start_reg[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .Q(
        start_reg[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .Q(
        start_reg[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .Q(
        start_reg[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .Q(
        start_reg[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .Q(
        start_reg[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .Q(
        start_reg[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .Q(
        start_reg[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .Q(
        start_reg[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .Q(
        start_reg[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .Q(
        start_reg[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .Q(
        start_reg[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .Q(
        start_reg[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .Q(
        start_reg[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .Q(
        start_reg[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .Q(
        start_reg[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .Q(
        start_reg[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .Q(
        start_reg[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .Q(
        start_reg[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .Q(
        start_reg[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .Q(
        start_reg[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .Q(
        start_reg[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .Q(
        start_reg[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .Q(
        start_reg[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .Q(
        start_reg[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .Q(
        start_reg[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .Q(
        start_reg[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .Q(
        start_reg[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .Q(
        start_reg[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .Q(
        start_reg[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .Q(
        start_reg[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .Q(
        start_reg[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .Q(
        start_reg[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .Q(
        start_reg[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .Q(
        start_reg[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .Q(
        start_reg[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .Q(
        start_reg[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .Q(
        start_reg[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .Q(
        start_reg[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .Q(
        start_reg[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .Q(
        start_reg[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .Q(
        start_reg[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .Q(
        start_reg[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .Q(
        start_reg[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .Q(
        start_reg[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .Q(
        start_reg[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .Q(
        start_reg[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .Q(
        start_reg[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .Q(
        start_reg[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .Q(
        start_reg[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .Q(
        start_reg[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .Q(
        start_reg[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .Q(
        start_reg[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .Q(
        start_reg[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .Q(
        start_reg[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .Q(
        start_reg[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .Q(
        start_reg[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .Q(
        start_reg[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .Q(
        start_reg[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .Q(
        start_reg[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .Q(
        start_reg[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .Q(
        start_reg[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .Q(
        start_reg[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .Q(
        start_reg[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .Q(
        start_reg[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .Q(
        start_reg[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .Q(
        start_reg[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .Q(
        start_reg[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .Q(
        start_reg[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .Q(
        start_reg[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .Q(
        start_reg[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .Q(
        start_reg[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .Q(
        start_reg[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .Q(
        start_reg[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .Q(
        start_reg[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .Q(
        start_reg[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .Q(
        start_reg[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .Q(
        start_reg[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .Q(
        start_reg[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .Q(
        start_reg[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .Q(
        start_reg[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .Q(
        start_reg[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .Q(
        start_reg[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .Q(
        start_reg[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .Q(
        start_reg[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .Q(
        start_reg[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .Q(
        start_reg[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .Q(
        start_reg[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .Q(
        start_reg[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .Q(
        start_reg[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .Q(
        start_reg[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .Q(
        start_reg[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .Q(
        start_reg[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .Q(
        start_reg[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .Q(
        start_reg[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .Q(
        start_reg[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .Q(
        start_reg[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .Q(
        start_reg[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .Q(
        start_reg[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .Q(
        start_reg[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .Q(
        start_reg[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .Q(
        start_reg[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .Q(
        start_reg[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .Q(
        start_reg[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .Q(
        start_reg[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .Q(
        start_reg[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .Q(
        start_reg[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .Q(
        start_reg[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .Q(
        start_reg[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .Q(
        start_reg[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .Q(
        start_reg[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .Q(
        start_reg[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .Q(
        start_reg[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .Q(
        start_reg[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .Q(
        start_reg[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .Q(
        start_reg[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .Q(
        start_reg[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .Q(
        start_reg[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .Q(
        start_reg[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .Q(
        start_reg[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .Q(
        start_reg[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .Q(
        start_reg[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .Q(
        start_reg[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .Q(
        start_reg[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .Q(
        start_reg[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .Q(
        start_reg[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .Q(
        start_reg[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .Q(
        start_reg[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .Q(
        start_reg[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .Q(
        start_reg[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .Q(
        start_reg[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .Q(
        start_reg[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .Q(
        start_reg[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .Q(
        start_reg[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .Q(
        start_reg[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .Q(
        start_reg[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .Q(
        start_reg[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .Q(
        start_reg[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .Q(
        start_reg[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .Q(
        start_reg[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .Q(
        start_reg[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .Q(
        start_reg[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .Q(
        start_reg[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .Q(
        start_reg[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .Q(
        start_reg[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .Q(
        start_reg[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .Q(
        start_reg[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .Q(
        start_reg[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .Q(
        start_reg[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .Q(
        start_reg[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .Q(
        start_reg[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .Q(
        start_reg[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .Q(
        start_reg[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .Q(
        start_reg[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .Q(
        start_reg[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .Q(
        start_reg[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .Q(
        start_reg[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .Q(
        start_reg[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .Q(
        start_reg[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .Q(
        start_reg[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .Q(
        start_reg[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .Q(
        start_reg[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .Q(
        start_reg[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .Q(
        start_reg[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .Q(
        start_reg[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .Q(
        start_reg[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .Q(
        start_reg[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .Q(
        start_reg[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .Q(
        start_reg[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .Q(
        start_reg[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .Q(
        start_reg[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .Q(
        start_reg[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .Q(
        start_reg[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .Q(
        start_reg[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .Q(
        start_reg[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .Q(
        start_reg[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .Q(
        start_reg[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .Q(
        start_reg[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .Q(
        start_reg[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .Q(
        start_reg[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .Q(
        start_reg[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .Q(
        start_reg[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .Q(
        start_reg[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .Q(
        start_reg[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .Q(
        start_reg[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .Q(
        start_reg[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .Q(
        start_reg[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .Q(
        start_reg[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .Q(
        start_reg[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .Q(
        start_reg[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .Q(
        start_reg[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .Q(
        start_reg[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .Q(
        start_reg[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .Q(
        start_reg[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .Q(
        start_reg[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .Q(
        start_reg[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .Q(
        start_reg[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .Q(
        start_reg[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .Q(
        start_reg[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .Q(
        start_reg[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .Q(
        start_reg[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .Q(
        start_reg[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .Q(
        start_reg[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .Q(
        start_reg[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .Q(
        start_reg[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .Q(
        start_reg[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .Q(
        start_reg[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .Q(
        start_reg[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .Q(
        start_reg[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .Q(
        start_reg[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .Q(
        start_reg[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .Q(
        start_reg[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .Q(
        start_reg[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .Q(
        start_reg[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .Q(
        start_reg[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .Q(
        start_reg[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .Q(
        start_reg[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .Q(
        start_reg[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .Q(
        start_reg[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .Q(
        start_reg[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .Q(
        start_reg[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .Q(
        start_reg[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .Q(
        start_reg[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .Q(
        start_reg[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .Q(
        start_reg[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .Q(
        start_reg[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .Q(
        start_reg[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .Q(
        start_reg[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .Q(
        start_reg[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .Q(
        start_reg[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .Q(
        start_reg[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .Q(
        start_reg[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .Q(
        start_reg[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .Q(
        start_reg[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .Q(
        start_reg[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .Q(
        start_reg[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .Q(
        start_reg[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .Q(
        start_reg[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .Q(
        start_reg[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .Q(
        start_reg[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .Q(
        start_reg[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .Q(
        start_reg[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .Q(
        start_reg[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .Q(
        start_reg[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .Q(
        start_reg[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .Q(
        start_reg[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .Q(
        start_reg[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .Q(
        start_reg[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .Q(
        start_reg[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .Q(
        start_reg[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .Q(
        start_reg[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .Q(
        start_reg[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .Q(
        start_reg[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .Q(
        start_reg[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .Q(
        start_reg[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .Q(
        start_reg[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .Q(
        start_reg[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .Q(
        start_reg[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .Q(
        start_reg[511]) );
  DFF mul_pow_reg ( .D(n3859), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n3858), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n3857), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n3856), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n3855), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n3854), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n3853), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n3852), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n3851), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n3850), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n3849), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n3848), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n3847), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n3846), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n3845), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n3844), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n3843), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n3842), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n3841), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n3840), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n3839), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n3838), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n3837), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n3836), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n3835), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n3834), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n3833), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n3832), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n3831), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n3830), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n3829), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n3828), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n3827), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n3826), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n3825), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n3824), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n3823), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n3822), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n3821), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n3820), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n3819), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n3818), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n3817), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n3816), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n3815), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n3814), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n3813), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n3812), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n3811), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n3810), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n3809), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n3808), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n3807), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n3806), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n3805), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n3804), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n3803), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n3802), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n3801), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n3800), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n3799), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n3798), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n3797), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n3796), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n3795), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n3794), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n3793), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n3792), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n3791), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n3790), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n3789), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n3788), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n3787), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n3786), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n3785), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n3784), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n3783), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n3782), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n3781), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n3780), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n3779), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n3778), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n3777), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n3776), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n3775), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n3774), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n3773), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n3772), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n3771), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n3770), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n3769), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n3768), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n3767), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n3766), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n3765), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n3764), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n3763), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n3762), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n3761), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n3760), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n3759), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n3758), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n3757), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n3756), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n3755), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n3754), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n3753), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n3752), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n3751), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n3750), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n3749), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n3748), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n3747), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n3746), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n3745), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n3744), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n3743), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n3742), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n3741), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n3740), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n3739), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n3738), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n3737), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n3736), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n3735), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n3734), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n3733), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n3732), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n3731), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n3730), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n3729), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n3728), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n3727), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n3726), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n3725), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n3724), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n3723), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n3722), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n3721), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n3720), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n3719), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n3718), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n3717), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n3716), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n3715), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n3714), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n3713), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n3712), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n3711), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n3710), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n3709), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n3708), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n3707), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n3706), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n3705), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n3704), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n3703), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n3702), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n3701), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n3700), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n3699), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n3698), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n3697), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n3696), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n3695), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n3694), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n3693), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n3692), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n3691), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n3690), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n3689), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n3688), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n3687), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n3686), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n3685), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n3684), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n3683), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n3682), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n3681), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n3680), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n3679), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n3678), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n3677), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n3676), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n3675), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n3674), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n3673), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n3672), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n3671), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n3670), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n3669), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n3668), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n3667), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n3666), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n3665), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n3664), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n3663), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n3662), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n3661), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n3660), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n3659), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n3658), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n3657), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n3656), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n3655), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n3654), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n3653), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n3652), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n3651), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n3650), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n3649), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n3648), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n3647), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n3646), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n3645), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n3644), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n3643), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n3642), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n3641), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n3640), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n3639), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n3638), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n3637), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n3636), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n3635), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n3634), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n3633), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n3632), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n3631), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n3630), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n3629), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n3628), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n3627), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n3626), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n3625), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n3624), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n3623), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n3622), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n3621), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n3620), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n3619), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n3618), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n3617), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n3616), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n3615), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n3614), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n3613), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n3612), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n3611), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n3610), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n3609), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n3608), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n3607), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n3606), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n3605), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n3604), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n3603), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF first_one_reg ( .D(n3346), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n3601), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n3600), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n3599), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n3598), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n3597), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n3596), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n3595), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n3594), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n3593), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n3592), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n3591), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n3590), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n3589), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n3588), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n3587), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n3586), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n3585), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n3584), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n3583), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n3582), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n3581), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n3580), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n3579), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n3578), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n3577), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n3576), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n3575), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n3574), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n3573), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n3572), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n3571), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n3570), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n3569), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n3568), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n3567), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n3566), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n3565), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n3564), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n3563), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n3562), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n3561), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n3560), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n3559), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n3558), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n3557), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n3556), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n3555), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n3554), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n3553), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n3552), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n3551), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n3550), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n3549), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n3548), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n3547), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n3546), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n3545), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n3544), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n3543), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n3542), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n3541), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n3540), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n3539), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n3538), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n3537), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n3536), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n3535), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n3534), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n3533), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n3532), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n3531), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n3530), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n3529), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n3528), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n3527), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n3526), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n3525), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n3524), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n3523), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n3522), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n3521), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n3520), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n3519), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n3518), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n3517), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n3516), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n3515), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n3514), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n3513), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n3512), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n3511), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n3510), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n3509), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n3508), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n3507), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n3506), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n3505), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n3504), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n3503), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n3502), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n3501), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n3500), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n3499), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n3498), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n3497), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n3496), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n3495), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n3494), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n3493), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n3492), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n3491), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n3490), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n3489), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n3488), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n3487), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n3486), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n3485), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n3484), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n3483), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n3482), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n3481), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n3480), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n3479), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n3478), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n3477), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n3476), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n3475), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n3474), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n3473), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n3472), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n3471), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n3470), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n3469), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n3468), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n3467), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n3466), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n3465), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n3464), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n3463), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n3462), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n3461), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n3460), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n3459), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n3458), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n3457), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n3456), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n3455), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n3454), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n3453), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n3452), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n3451), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n3450), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n3449), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n3448), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n3447), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n3446), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n3445), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n3444), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n3443), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n3442), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n3441), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n3440), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n3439), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n3438), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n3437), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n3436), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n3435), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n3434), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n3433), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n3432), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n3431), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n3430), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n3429), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n3428), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n3427), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n3426), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n3425), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n3424), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n3423), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n3422), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n3421), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n3420), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n3419), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n3418), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n3417), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n3416), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n3415), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n3414), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n3413), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n3412), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n3411), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n3410), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n3409), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n3408), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n3407), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n3406), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n3405), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n3404), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n3403), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n3402), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n3401), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n3400), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n3399), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n3398), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n3397), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n3396), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n3395), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n3394), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n3393), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n3392), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n3391), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n3390), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n3389), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n3388), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n3387), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n3386), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n3385), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n3384), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n3383), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n3382), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n3381), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n3380), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n3379), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n3378), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n3377), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n3376), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n3375), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n3374), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n3373), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n3372), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n3371), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n3370), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n3369), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n3368), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n3367), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n3366), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n3365), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n3364), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n3363), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n3362), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n3361), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n3360), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n3359), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n3358), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n3357), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n3356), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n3355), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n3354), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n3353), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n3352), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n3351), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n3350), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n3349), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n3348), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n3347), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n3602), .CLK(clk), .RST(rst), .Q(creg[255]) );
  NAND U5142 ( .A(n3860), .B(n3861), .Z(y[9]) );
  NAND U5143 ( .A(n3862), .B(m[9]), .Z(n3861) );
  NAND U5144 ( .A(n3863), .B(creg[9]), .Z(n3860) );
  NAND U5145 ( .A(n3864), .B(n3865), .Z(y[99]) );
  NAND U5146 ( .A(n3862), .B(m[99]), .Z(n3865) );
  NAND U5147 ( .A(n3863), .B(creg[99]), .Z(n3864) );
  NAND U5148 ( .A(n3866), .B(n3867), .Z(y[98]) );
  NAND U5149 ( .A(n3862), .B(m[98]), .Z(n3867) );
  NAND U5150 ( .A(n3863), .B(creg[98]), .Z(n3866) );
  NAND U5151 ( .A(n3868), .B(n3869), .Z(y[97]) );
  NAND U5152 ( .A(n3862), .B(m[97]), .Z(n3869) );
  NAND U5153 ( .A(n3863), .B(creg[97]), .Z(n3868) );
  NAND U5154 ( .A(n3870), .B(n3871), .Z(y[96]) );
  NAND U5155 ( .A(n3862), .B(m[96]), .Z(n3871) );
  NAND U5156 ( .A(n3863), .B(creg[96]), .Z(n3870) );
  NAND U5157 ( .A(n3872), .B(n3873), .Z(y[95]) );
  NAND U5158 ( .A(n3862), .B(m[95]), .Z(n3873) );
  NAND U5159 ( .A(n3863), .B(creg[95]), .Z(n3872) );
  NAND U5160 ( .A(n3874), .B(n3875), .Z(y[94]) );
  NAND U5161 ( .A(n3862), .B(m[94]), .Z(n3875) );
  NAND U5162 ( .A(n3863), .B(creg[94]), .Z(n3874) );
  NAND U5163 ( .A(n3876), .B(n3877), .Z(y[93]) );
  NAND U5164 ( .A(n3862), .B(m[93]), .Z(n3877) );
  NAND U5165 ( .A(n3863), .B(creg[93]), .Z(n3876) );
  NAND U5166 ( .A(n3878), .B(n3879), .Z(y[92]) );
  NAND U5167 ( .A(n3862), .B(m[92]), .Z(n3879) );
  NAND U5168 ( .A(n3863), .B(creg[92]), .Z(n3878) );
  NAND U5169 ( .A(n3880), .B(n3881), .Z(y[91]) );
  NAND U5170 ( .A(n3862), .B(m[91]), .Z(n3881) );
  NAND U5171 ( .A(n3863), .B(creg[91]), .Z(n3880) );
  NAND U5172 ( .A(n3882), .B(n3883), .Z(y[90]) );
  NAND U5173 ( .A(n3862), .B(m[90]), .Z(n3883) );
  NAND U5174 ( .A(n3863), .B(creg[90]), .Z(n3882) );
  NAND U5175 ( .A(n3884), .B(n3885), .Z(y[8]) );
  NAND U5176 ( .A(n3862), .B(m[8]), .Z(n3885) );
  NAND U5177 ( .A(n3863), .B(creg[8]), .Z(n3884) );
  NAND U5178 ( .A(n3886), .B(n3887), .Z(y[89]) );
  NAND U5179 ( .A(n3862), .B(m[89]), .Z(n3887) );
  NAND U5180 ( .A(n3863), .B(creg[89]), .Z(n3886) );
  NAND U5181 ( .A(n3888), .B(n3889), .Z(y[88]) );
  NAND U5182 ( .A(n3862), .B(m[88]), .Z(n3889) );
  NAND U5183 ( .A(n3863), .B(creg[88]), .Z(n3888) );
  NAND U5184 ( .A(n3890), .B(n3891), .Z(y[87]) );
  NAND U5185 ( .A(n3862), .B(m[87]), .Z(n3891) );
  NAND U5186 ( .A(n3863), .B(creg[87]), .Z(n3890) );
  NAND U5187 ( .A(n3892), .B(n3893), .Z(y[86]) );
  NAND U5188 ( .A(n3862), .B(m[86]), .Z(n3893) );
  NAND U5189 ( .A(n3863), .B(creg[86]), .Z(n3892) );
  NAND U5190 ( .A(n3894), .B(n3895), .Z(y[85]) );
  NAND U5191 ( .A(n3862), .B(m[85]), .Z(n3895) );
  NAND U5192 ( .A(n3863), .B(creg[85]), .Z(n3894) );
  NAND U5193 ( .A(n3896), .B(n3897), .Z(y[84]) );
  NAND U5194 ( .A(n3862), .B(m[84]), .Z(n3897) );
  NAND U5195 ( .A(n3863), .B(creg[84]), .Z(n3896) );
  NAND U5196 ( .A(n3898), .B(n3899), .Z(y[83]) );
  NAND U5197 ( .A(n3862), .B(m[83]), .Z(n3899) );
  NAND U5198 ( .A(n3863), .B(creg[83]), .Z(n3898) );
  NAND U5199 ( .A(n3900), .B(n3901), .Z(y[82]) );
  NAND U5200 ( .A(n3862), .B(m[82]), .Z(n3901) );
  NAND U5201 ( .A(n3863), .B(creg[82]), .Z(n3900) );
  NAND U5202 ( .A(n3902), .B(n3903), .Z(y[81]) );
  NAND U5203 ( .A(n3862), .B(m[81]), .Z(n3903) );
  NAND U5204 ( .A(n3863), .B(creg[81]), .Z(n3902) );
  NAND U5205 ( .A(n3904), .B(n3905), .Z(y[80]) );
  NAND U5206 ( .A(n3862), .B(m[80]), .Z(n3905) );
  NAND U5207 ( .A(n3863), .B(creg[80]), .Z(n3904) );
  NAND U5208 ( .A(n3906), .B(n3907), .Z(y[7]) );
  NAND U5209 ( .A(n3862), .B(m[7]), .Z(n3907) );
  NAND U5210 ( .A(n3863), .B(creg[7]), .Z(n3906) );
  NAND U5211 ( .A(n3908), .B(n3909), .Z(y[79]) );
  NAND U5212 ( .A(n3862), .B(m[79]), .Z(n3909) );
  NAND U5213 ( .A(n3863), .B(creg[79]), .Z(n3908) );
  NAND U5214 ( .A(n3910), .B(n3911), .Z(y[78]) );
  NAND U5215 ( .A(n3862), .B(m[78]), .Z(n3911) );
  NAND U5216 ( .A(n3863), .B(creg[78]), .Z(n3910) );
  NAND U5217 ( .A(n3912), .B(n3913), .Z(y[77]) );
  NAND U5218 ( .A(n3862), .B(m[77]), .Z(n3913) );
  NAND U5219 ( .A(n3863), .B(creg[77]), .Z(n3912) );
  NAND U5220 ( .A(n3914), .B(n3915), .Z(y[76]) );
  NAND U5221 ( .A(n3862), .B(m[76]), .Z(n3915) );
  NAND U5222 ( .A(n3863), .B(creg[76]), .Z(n3914) );
  NAND U5223 ( .A(n3916), .B(n3917), .Z(y[75]) );
  NAND U5224 ( .A(n3862), .B(m[75]), .Z(n3917) );
  NAND U5225 ( .A(n3863), .B(creg[75]), .Z(n3916) );
  NAND U5226 ( .A(n3918), .B(n3919), .Z(y[74]) );
  NAND U5227 ( .A(n3862), .B(m[74]), .Z(n3919) );
  NAND U5228 ( .A(n3863), .B(creg[74]), .Z(n3918) );
  NAND U5229 ( .A(n3920), .B(n3921), .Z(y[73]) );
  NAND U5230 ( .A(n3862), .B(m[73]), .Z(n3921) );
  NAND U5231 ( .A(n3863), .B(creg[73]), .Z(n3920) );
  NAND U5232 ( .A(n3922), .B(n3923), .Z(y[72]) );
  NAND U5233 ( .A(n3862), .B(m[72]), .Z(n3923) );
  NAND U5234 ( .A(n3863), .B(creg[72]), .Z(n3922) );
  NAND U5235 ( .A(n3924), .B(n3925), .Z(y[71]) );
  NAND U5236 ( .A(n3862), .B(m[71]), .Z(n3925) );
  NAND U5237 ( .A(n3863), .B(creg[71]), .Z(n3924) );
  NAND U5238 ( .A(n3926), .B(n3927), .Z(y[70]) );
  NAND U5239 ( .A(n3862), .B(m[70]), .Z(n3927) );
  NAND U5240 ( .A(n3863), .B(creg[70]), .Z(n3926) );
  NAND U5241 ( .A(n3928), .B(n3929), .Z(y[6]) );
  NAND U5242 ( .A(n3862), .B(m[6]), .Z(n3929) );
  NAND U5243 ( .A(n3863), .B(creg[6]), .Z(n3928) );
  NAND U5244 ( .A(n3930), .B(n3931), .Z(y[69]) );
  NAND U5245 ( .A(n3862), .B(m[69]), .Z(n3931) );
  NAND U5246 ( .A(n3863), .B(creg[69]), .Z(n3930) );
  NAND U5247 ( .A(n3932), .B(n3933), .Z(y[68]) );
  NAND U5248 ( .A(n3862), .B(m[68]), .Z(n3933) );
  NAND U5249 ( .A(n3863), .B(creg[68]), .Z(n3932) );
  NAND U5250 ( .A(n3934), .B(n3935), .Z(y[67]) );
  NAND U5251 ( .A(n3862), .B(m[67]), .Z(n3935) );
  NAND U5252 ( .A(n3863), .B(creg[67]), .Z(n3934) );
  NAND U5253 ( .A(n3936), .B(n3937), .Z(y[66]) );
  NAND U5254 ( .A(n3862), .B(m[66]), .Z(n3937) );
  NAND U5255 ( .A(n3863), .B(creg[66]), .Z(n3936) );
  NAND U5256 ( .A(n3938), .B(n3939), .Z(y[65]) );
  NAND U5257 ( .A(n3862), .B(m[65]), .Z(n3939) );
  NAND U5258 ( .A(n3863), .B(creg[65]), .Z(n3938) );
  NAND U5259 ( .A(n3940), .B(n3941), .Z(y[64]) );
  NAND U5260 ( .A(n3862), .B(m[64]), .Z(n3941) );
  NAND U5261 ( .A(n3863), .B(creg[64]), .Z(n3940) );
  NAND U5262 ( .A(n3942), .B(n3943), .Z(y[63]) );
  NAND U5263 ( .A(n3862), .B(m[63]), .Z(n3943) );
  NAND U5264 ( .A(n3863), .B(creg[63]), .Z(n3942) );
  NAND U5265 ( .A(n3944), .B(n3945), .Z(y[62]) );
  NAND U5266 ( .A(n3862), .B(m[62]), .Z(n3945) );
  NAND U5267 ( .A(n3863), .B(creg[62]), .Z(n3944) );
  NAND U5268 ( .A(n3946), .B(n3947), .Z(y[61]) );
  NAND U5269 ( .A(n3862), .B(m[61]), .Z(n3947) );
  NAND U5270 ( .A(n3863), .B(creg[61]), .Z(n3946) );
  NAND U5271 ( .A(n3948), .B(n3949), .Z(y[60]) );
  NAND U5272 ( .A(n3862), .B(m[60]), .Z(n3949) );
  NAND U5273 ( .A(n3863), .B(creg[60]), .Z(n3948) );
  NAND U5274 ( .A(n3950), .B(n3951), .Z(y[5]) );
  NAND U5275 ( .A(n3862), .B(m[5]), .Z(n3951) );
  NAND U5276 ( .A(n3863), .B(creg[5]), .Z(n3950) );
  NAND U5277 ( .A(n3952), .B(n3953), .Z(y[59]) );
  NAND U5278 ( .A(n3862), .B(m[59]), .Z(n3953) );
  NAND U5279 ( .A(n3863), .B(creg[59]), .Z(n3952) );
  NAND U5280 ( .A(n3954), .B(n3955), .Z(y[58]) );
  NAND U5281 ( .A(n3862), .B(m[58]), .Z(n3955) );
  NAND U5282 ( .A(n3863), .B(creg[58]), .Z(n3954) );
  NAND U5283 ( .A(n3956), .B(n3957), .Z(y[57]) );
  NAND U5284 ( .A(n3862), .B(m[57]), .Z(n3957) );
  NAND U5285 ( .A(n3863), .B(creg[57]), .Z(n3956) );
  NAND U5286 ( .A(n3958), .B(n3959), .Z(y[56]) );
  NAND U5287 ( .A(n3862), .B(m[56]), .Z(n3959) );
  NAND U5288 ( .A(n3863), .B(creg[56]), .Z(n3958) );
  NAND U5289 ( .A(n3960), .B(n3961), .Z(y[55]) );
  NAND U5290 ( .A(n3862), .B(m[55]), .Z(n3961) );
  NAND U5291 ( .A(n3863), .B(creg[55]), .Z(n3960) );
  NAND U5292 ( .A(n3962), .B(n3963), .Z(y[54]) );
  NAND U5293 ( .A(n3862), .B(m[54]), .Z(n3963) );
  NAND U5294 ( .A(n3863), .B(creg[54]), .Z(n3962) );
  NAND U5295 ( .A(n3964), .B(n3965), .Z(y[53]) );
  NAND U5296 ( .A(n3862), .B(m[53]), .Z(n3965) );
  NAND U5297 ( .A(n3863), .B(creg[53]), .Z(n3964) );
  NAND U5298 ( .A(n3966), .B(n3967), .Z(y[52]) );
  NAND U5299 ( .A(n3862), .B(m[52]), .Z(n3967) );
  NAND U5300 ( .A(n3863), .B(creg[52]), .Z(n3966) );
  NAND U5301 ( .A(n3968), .B(n3969), .Z(y[51]) );
  NAND U5302 ( .A(n3862), .B(m[51]), .Z(n3969) );
  NAND U5303 ( .A(n3863), .B(creg[51]), .Z(n3968) );
  NAND U5304 ( .A(n3970), .B(n3971), .Z(y[50]) );
  NAND U5305 ( .A(n3862), .B(m[50]), .Z(n3971) );
  NAND U5306 ( .A(n3863), .B(creg[50]), .Z(n3970) );
  NAND U5307 ( .A(n3972), .B(n3973), .Z(y[4]) );
  NAND U5308 ( .A(n3862), .B(m[4]), .Z(n3973) );
  NAND U5309 ( .A(n3863), .B(creg[4]), .Z(n3972) );
  NAND U5310 ( .A(n3974), .B(n3975), .Z(y[49]) );
  NAND U5311 ( .A(n3862), .B(m[49]), .Z(n3975) );
  NAND U5312 ( .A(n3863), .B(creg[49]), .Z(n3974) );
  NAND U5313 ( .A(n3976), .B(n3977), .Z(y[48]) );
  NAND U5314 ( .A(n3862), .B(m[48]), .Z(n3977) );
  NAND U5315 ( .A(n3863), .B(creg[48]), .Z(n3976) );
  NAND U5316 ( .A(n3978), .B(n3979), .Z(y[47]) );
  NAND U5317 ( .A(n3862), .B(m[47]), .Z(n3979) );
  NAND U5318 ( .A(n3863), .B(creg[47]), .Z(n3978) );
  NAND U5319 ( .A(n3980), .B(n3981), .Z(y[46]) );
  NAND U5320 ( .A(n3862), .B(m[46]), .Z(n3981) );
  NAND U5321 ( .A(n3863), .B(creg[46]), .Z(n3980) );
  NAND U5322 ( .A(n3982), .B(n3983), .Z(y[45]) );
  NAND U5323 ( .A(n3862), .B(m[45]), .Z(n3983) );
  NAND U5324 ( .A(n3863), .B(creg[45]), .Z(n3982) );
  NAND U5325 ( .A(n3984), .B(n3985), .Z(y[44]) );
  NAND U5326 ( .A(n3862), .B(m[44]), .Z(n3985) );
  NAND U5327 ( .A(n3863), .B(creg[44]), .Z(n3984) );
  NAND U5328 ( .A(n3986), .B(n3987), .Z(y[43]) );
  NAND U5329 ( .A(n3862), .B(m[43]), .Z(n3987) );
  NAND U5330 ( .A(n3863), .B(creg[43]), .Z(n3986) );
  NAND U5331 ( .A(n3988), .B(n3989), .Z(y[42]) );
  NAND U5332 ( .A(n3862), .B(m[42]), .Z(n3989) );
  NAND U5333 ( .A(n3863), .B(creg[42]), .Z(n3988) );
  NAND U5334 ( .A(n3990), .B(n3991), .Z(y[41]) );
  NAND U5335 ( .A(n3862), .B(m[41]), .Z(n3991) );
  NAND U5336 ( .A(n3863), .B(creg[41]), .Z(n3990) );
  NAND U5337 ( .A(n3992), .B(n3993), .Z(y[40]) );
  NAND U5338 ( .A(n3862), .B(m[40]), .Z(n3993) );
  NAND U5339 ( .A(n3863), .B(creg[40]), .Z(n3992) );
  NAND U5340 ( .A(n3994), .B(n3995), .Z(y[3]) );
  NAND U5341 ( .A(n3862), .B(m[3]), .Z(n3995) );
  NAND U5342 ( .A(n3863), .B(creg[3]), .Z(n3994) );
  NAND U5343 ( .A(n3996), .B(n3997), .Z(y[39]) );
  NAND U5344 ( .A(n3862), .B(m[39]), .Z(n3997) );
  NAND U5345 ( .A(n3863), .B(creg[39]), .Z(n3996) );
  NAND U5346 ( .A(n3998), .B(n3999), .Z(y[38]) );
  NAND U5347 ( .A(n3862), .B(m[38]), .Z(n3999) );
  NAND U5348 ( .A(n3863), .B(creg[38]), .Z(n3998) );
  NAND U5349 ( .A(n4000), .B(n4001), .Z(y[37]) );
  NAND U5350 ( .A(n3862), .B(m[37]), .Z(n4001) );
  NAND U5351 ( .A(n3863), .B(creg[37]), .Z(n4000) );
  NAND U5352 ( .A(n4002), .B(n4003), .Z(y[36]) );
  NAND U5353 ( .A(n3862), .B(m[36]), .Z(n4003) );
  NAND U5354 ( .A(n3863), .B(creg[36]), .Z(n4002) );
  NAND U5355 ( .A(n4004), .B(n4005), .Z(y[35]) );
  NAND U5356 ( .A(n3862), .B(m[35]), .Z(n4005) );
  NAND U5357 ( .A(n3863), .B(creg[35]), .Z(n4004) );
  NAND U5358 ( .A(n4006), .B(n4007), .Z(y[34]) );
  NAND U5359 ( .A(n3862), .B(m[34]), .Z(n4007) );
  NAND U5360 ( .A(n3863), .B(creg[34]), .Z(n4006) );
  NAND U5361 ( .A(n4008), .B(n4009), .Z(y[33]) );
  NAND U5362 ( .A(n3862), .B(m[33]), .Z(n4009) );
  NAND U5363 ( .A(n3863), .B(creg[33]), .Z(n4008) );
  NAND U5364 ( .A(n4010), .B(n4011), .Z(y[32]) );
  NAND U5365 ( .A(n3862), .B(m[32]), .Z(n4011) );
  NAND U5366 ( .A(n3863), .B(creg[32]), .Z(n4010) );
  NAND U5367 ( .A(n4012), .B(n4013), .Z(y[31]) );
  NAND U5368 ( .A(n3862), .B(m[31]), .Z(n4013) );
  NAND U5369 ( .A(n3863), .B(creg[31]), .Z(n4012) );
  NAND U5370 ( .A(n4014), .B(n4015), .Z(y[30]) );
  NAND U5371 ( .A(n3862), .B(m[30]), .Z(n4015) );
  NAND U5372 ( .A(n3863), .B(creg[30]), .Z(n4014) );
  NAND U5373 ( .A(n4016), .B(n4017), .Z(y[2]) );
  NAND U5374 ( .A(n3862), .B(m[2]), .Z(n4017) );
  NAND U5375 ( .A(n3863), .B(creg[2]), .Z(n4016) );
  NAND U5376 ( .A(n4018), .B(n4019), .Z(y[29]) );
  NAND U5377 ( .A(n3862), .B(m[29]), .Z(n4019) );
  NAND U5378 ( .A(n3863), .B(creg[29]), .Z(n4018) );
  NAND U5379 ( .A(n4020), .B(n4021), .Z(y[28]) );
  NAND U5380 ( .A(n3862), .B(m[28]), .Z(n4021) );
  NAND U5381 ( .A(n3863), .B(creg[28]), .Z(n4020) );
  NAND U5382 ( .A(n4022), .B(n4023), .Z(y[27]) );
  NAND U5383 ( .A(n3862), .B(m[27]), .Z(n4023) );
  NAND U5384 ( .A(n3863), .B(creg[27]), .Z(n4022) );
  NAND U5385 ( .A(n4024), .B(n4025), .Z(y[26]) );
  NAND U5386 ( .A(n3862), .B(m[26]), .Z(n4025) );
  NAND U5387 ( .A(n3863), .B(creg[26]), .Z(n4024) );
  NAND U5388 ( .A(n4026), .B(n4027), .Z(y[25]) );
  NAND U5389 ( .A(n3862), .B(m[25]), .Z(n4027) );
  NAND U5390 ( .A(n3863), .B(creg[25]), .Z(n4026) );
  NAND U5391 ( .A(n4028), .B(n4029), .Z(y[255]) );
  NAND U5392 ( .A(n3862), .B(m[255]), .Z(n4029) );
  NAND U5393 ( .A(n3863), .B(creg[255]), .Z(n4028) );
  NAND U5394 ( .A(n4030), .B(n4031), .Z(y[254]) );
  NAND U5395 ( .A(n3862), .B(m[254]), .Z(n4031) );
  NAND U5396 ( .A(n3863), .B(creg[254]), .Z(n4030) );
  NAND U5397 ( .A(n4032), .B(n4033), .Z(y[253]) );
  NAND U5398 ( .A(n3862), .B(m[253]), .Z(n4033) );
  NAND U5399 ( .A(n3863), .B(creg[253]), .Z(n4032) );
  NAND U5400 ( .A(n4034), .B(n4035), .Z(y[252]) );
  NAND U5401 ( .A(n3862), .B(m[252]), .Z(n4035) );
  NAND U5402 ( .A(n3863), .B(creg[252]), .Z(n4034) );
  NAND U5403 ( .A(n4036), .B(n4037), .Z(y[251]) );
  NAND U5404 ( .A(n3862), .B(m[251]), .Z(n4037) );
  NAND U5405 ( .A(n3863), .B(creg[251]), .Z(n4036) );
  NAND U5406 ( .A(n4038), .B(n4039), .Z(y[250]) );
  NAND U5407 ( .A(n3862), .B(m[250]), .Z(n4039) );
  NAND U5408 ( .A(n3863), .B(creg[250]), .Z(n4038) );
  NAND U5409 ( .A(n4040), .B(n4041), .Z(y[24]) );
  NAND U5410 ( .A(n3862), .B(m[24]), .Z(n4041) );
  NAND U5411 ( .A(n3863), .B(creg[24]), .Z(n4040) );
  NAND U5412 ( .A(n4042), .B(n4043), .Z(y[249]) );
  NAND U5413 ( .A(n3862), .B(m[249]), .Z(n4043) );
  NAND U5414 ( .A(n3863), .B(creg[249]), .Z(n4042) );
  NAND U5415 ( .A(n4044), .B(n4045), .Z(y[248]) );
  NAND U5416 ( .A(n3862), .B(m[248]), .Z(n4045) );
  NAND U5417 ( .A(n3863), .B(creg[248]), .Z(n4044) );
  NAND U5418 ( .A(n4046), .B(n4047), .Z(y[247]) );
  NAND U5419 ( .A(n3862), .B(m[247]), .Z(n4047) );
  NAND U5420 ( .A(n3863), .B(creg[247]), .Z(n4046) );
  NAND U5421 ( .A(n4048), .B(n4049), .Z(y[246]) );
  NAND U5422 ( .A(n3862), .B(m[246]), .Z(n4049) );
  NAND U5423 ( .A(n3863), .B(creg[246]), .Z(n4048) );
  NAND U5424 ( .A(n4050), .B(n4051), .Z(y[245]) );
  NAND U5425 ( .A(n3862), .B(m[245]), .Z(n4051) );
  NAND U5426 ( .A(n3863), .B(creg[245]), .Z(n4050) );
  NAND U5427 ( .A(n4052), .B(n4053), .Z(y[244]) );
  NAND U5428 ( .A(n3862), .B(m[244]), .Z(n4053) );
  NAND U5429 ( .A(n3863), .B(creg[244]), .Z(n4052) );
  NAND U5430 ( .A(n4054), .B(n4055), .Z(y[243]) );
  NAND U5431 ( .A(n3862), .B(m[243]), .Z(n4055) );
  NAND U5432 ( .A(n3863), .B(creg[243]), .Z(n4054) );
  NAND U5433 ( .A(n4056), .B(n4057), .Z(y[242]) );
  NAND U5434 ( .A(n3862), .B(m[242]), .Z(n4057) );
  NAND U5435 ( .A(n3863), .B(creg[242]), .Z(n4056) );
  NAND U5436 ( .A(n4058), .B(n4059), .Z(y[241]) );
  NAND U5437 ( .A(n3862), .B(m[241]), .Z(n4059) );
  NAND U5438 ( .A(n3863), .B(creg[241]), .Z(n4058) );
  NAND U5439 ( .A(n4060), .B(n4061), .Z(y[240]) );
  NAND U5440 ( .A(n3862), .B(m[240]), .Z(n4061) );
  NAND U5441 ( .A(n3863), .B(creg[240]), .Z(n4060) );
  NAND U5442 ( .A(n4062), .B(n4063), .Z(y[23]) );
  NAND U5443 ( .A(n3862), .B(m[23]), .Z(n4063) );
  NAND U5444 ( .A(n3863), .B(creg[23]), .Z(n4062) );
  NAND U5445 ( .A(n4064), .B(n4065), .Z(y[239]) );
  NAND U5446 ( .A(n3862), .B(m[239]), .Z(n4065) );
  NAND U5447 ( .A(n3863), .B(creg[239]), .Z(n4064) );
  NAND U5448 ( .A(n4066), .B(n4067), .Z(y[238]) );
  NAND U5449 ( .A(n3862), .B(m[238]), .Z(n4067) );
  NAND U5450 ( .A(n3863), .B(creg[238]), .Z(n4066) );
  NAND U5451 ( .A(n4068), .B(n4069), .Z(y[237]) );
  NAND U5452 ( .A(n3862), .B(m[237]), .Z(n4069) );
  NAND U5453 ( .A(n3863), .B(creg[237]), .Z(n4068) );
  NAND U5454 ( .A(n4070), .B(n4071), .Z(y[236]) );
  NAND U5455 ( .A(n3862), .B(m[236]), .Z(n4071) );
  NAND U5456 ( .A(n3863), .B(creg[236]), .Z(n4070) );
  NAND U5457 ( .A(n4072), .B(n4073), .Z(y[235]) );
  NAND U5458 ( .A(n3862), .B(m[235]), .Z(n4073) );
  NAND U5459 ( .A(n3863), .B(creg[235]), .Z(n4072) );
  NAND U5460 ( .A(n4074), .B(n4075), .Z(y[234]) );
  NAND U5461 ( .A(n3862), .B(m[234]), .Z(n4075) );
  NAND U5462 ( .A(n3863), .B(creg[234]), .Z(n4074) );
  NAND U5463 ( .A(n4076), .B(n4077), .Z(y[233]) );
  NAND U5464 ( .A(n3862), .B(m[233]), .Z(n4077) );
  NAND U5465 ( .A(n3863), .B(creg[233]), .Z(n4076) );
  NAND U5466 ( .A(n4078), .B(n4079), .Z(y[232]) );
  NAND U5467 ( .A(n3862), .B(m[232]), .Z(n4079) );
  NAND U5468 ( .A(n3863), .B(creg[232]), .Z(n4078) );
  NAND U5469 ( .A(n4080), .B(n4081), .Z(y[231]) );
  NAND U5470 ( .A(n3862), .B(m[231]), .Z(n4081) );
  NAND U5471 ( .A(n3863), .B(creg[231]), .Z(n4080) );
  NAND U5472 ( .A(n4082), .B(n4083), .Z(y[230]) );
  NAND U5473 ( .A(n3862), .B(m[230]), .Z(n4083) );
  NAND U5474 ( .A(n3863), .B(creg[230]), .Z(n4082) );
  NAND U5475 ( .A(n4084), .B(n4085), .Z(y[22]) );
  NAND U5476 ( .A(n3862), .B(m[22]), .Z(n4085) );
  NAND U5477 ( .A(n3863), .B(creg[22]), .Z(n4084) );
  NAND U5478 ( .A(n4086), .B(n4087), .Z(y[229]) );
  NAND U5479 ( .A(n3862), .B(m[229]), .Z(n4087) );
  NAND U5480 ( .A(n3863), .B(creg[229]), .Z(n4086) );
  NAND U5481 ( .A(n4088), .B(n4089), .Z(y[228]) );
  NAND U5482 ( .A(n3862), .B(m[228]), .Z(n4089) );
  NAND U5483 ( .A(n3863), .B(creg[228]), .Z(n4088) );
  NAND U5484 ( .A(n4090), .B(n4091), .Z(y[227]) );
  NAND U5485 ( .A(n3862), .B(m[227]), .Z(n4091) );
  NAND U5486 ( .A(n3863), .B(creg[227]), .Z(n4090) );
  NAND U5487 ( .A(n4092), .B(n4093), .Z(y[226]) );
  NAND U5488 ( .A(n3862), .B(m[226]), .Z(n4093) );
  NAND U5489 ( .A(n3863), .B(creg[226]), .Z(n4092) );
  NAND U5490 ( .A(n4094), .B(n4095), .Z(y[225]) );
  NAND U5491 ( .A(n3862), .B(m[225]), .Z(n4095) );
  NAND U5492 ( .A(n3863), .B(creg[225]), .Z(n4094) );
  NAND U5493 ( .A(n4096), .B(n4097), .Z(y[224]) );
  NAND U5494 ( .A(n3862), .B(m[224]), .Z(n4097) );
  NAND U5495 ( .A(n3863), .B(creg[224]), .Z(n4096) );
  NAND U5496 ( .A(n4098), .B(n4099), .Z(y[223]) );
  NAND U5497 ( .A(n3862), .B(m[223]), .Z(n4099) );
  NAND U5498 ( .A(n3863), .B(creg[223]), .Z(n4098) );
  NAND U5499 ( .A(n4100), .B(n4101), .Z(y[222]) );
  NAND U5500 ( .A(n3862), .B(m[222]), .Z(n4101) );
  NAND U5501 ( .A(n3863), .B(creg[222]), .Z(n4100) );
  NAND U5502 ( .A(n4102), .B(n4103), .Z(y[221]) );
  NAND U5503 ( .A(n3862), .B(m[221]), .Z(n4103) );
  NAND U5504 ( .A(n3863), .B(creg[221]), .Z(n4102) );
  NAND U5505 ( .A(n4104), .B(n4105), .Z(y[220]) );
  NAND U5506 ( .A(n3862), .B(m[220]), .Z(n4105) );
  NAND U5507 ( .A(n3863), .B(creg[220]), .Z(n4104) );
  NAND U5508 ( .A(n4106), .B(n4107), .Z(y[21]) );
  NAND U5509 ( .A(n3862), .B(m[21]), .Z(n4107) );
  NAND U5510 ( .A(n3863), .B(creg[21]), .Z(n4106) );
  NAND U5511 ( .A(n4108), .B(n4109), .Z(y[219]) );
  NAND U5512 ( .A(n3862), .B(m[219]), .Z(n4109) );
  NAND U5513 ( .A(n3863), .B(creg[219]), .Z(n4108) );
  NAND U5514 ( .A(n4110), .B(n4111), .Z(y[218]) );
  NAND U5515 ( .A(n3862), .B(m[218]), .Z(n4111) );
  NAND U5516 ( .A(n3863), .B(creg[218]), .Z(n4110) );
  NAND U5517 ( .A(n4112), .B(n4113), .Z(y[217]) );
  NAND U5518 ( .A(n3862), .B(m[217]), .Z(n4113) );
  NAND U5519 ( .A(n3863), .B(creg[217]), .Z(n4112) );
  NAND U5520 ( .A(n4114), .B(n4115), .Z(y[216]) );
  NAND U5521 ( .A(n3862), .B(m[216]), .Z(n4115) );
  NAND U5522 ( .A(n3863), .B(creg[216]), .Z(n4114) );
  NAND U5523 ( .A(n4116), .B(n4117), .Z(y[215]) );
  NAND U5524 ( .A(n3862), .B(m[215]), .Z(n4117) );
  NAND U5525 ( .A(n3863), .B(creg[215]), .Z(n4116) );
  NAND U5526 ( .A(n4118), .B(n4119), .Z(y[214]) );
  NAND U5527 ( .A(n3862), .B(m[214]), .Z(n4119) );
  NAND U5528 ( .A(n3863), .B(creg[214]), .Z(n4118) );
  NAND U5529 ( .A(n4120), .B(n4121), .Z(y[213]) );
  NAND U5530 ( .A(n3862), .B(m[213]), .Z(n4121) );
  NAND U5531 ( .A(n3863), .B(creg[213]), .Z(n4120) );
  NAND U5532 ( .A(n4122), .B(n4123), .Z(y[212]) );
  NAND U5533 ( .A(n3862), .B(m[212]), .Z(n4123) );
  NAND U5534 ( .A(n3863), .B(creg[212]), .Z(n4122) );
  NAND U5535 ( .A(n4124), .B(n4125), .Z(y[211]) );
  NAND U5536 ( .A(n3862), .B(m[211]), .Z(n4125) );
  NAND U5537 ( .A(n3863), .B(creg[211]), .Z(n4124) );
  NAND U5538 ( .A(n4126), .B(n4127), .Z(y[210]) );
  NAND U5539 ( .A(n3862), .B(m[210]), .Z(n4127) );
  NAND U5540 ( .A(n3863), .B(creg[210]), .Z(n4126) );
  NAND U5541 ( .A(n4128), .B(n4129), .Z(y[20]) );
  NAND U5542 ( .A(n3862), .B(m[20]), .Z(n4129) );
  NAND U5543 ( .A(n3863), .B(creg[20]), .Z(n4128) );
  NAND U5544 ( .A(n4130), .B(n4131), .Z(y[209]) );
  NAND U5545 ( .A(n3862), .B(m[209]), .Z(n4131) );
  NAND U5546 ( .A(n3863), .B(creg[209]), .Z(n4130) );
  NAND U5547 ( .A(n4132), .B(n4133), .Z(y[208]) );
  NAND U5548 ( .A(n3862), .B(m[208]), .Z(n4133) );
  NAND U5549 ( .A(n3863), .B(creg[208]), .Z(n4132) );
  NAND U5550 ( .A(n4134), .B(n4135), .Z(y[207]) );
  NAND U5551 ( .A(n3862), .B(m[207]), .Z(n4135) );
  NAND U5552 ( .A(n3863), .B(creg[207]), .Z(n4134) );
  NAND U5553 ( .A(n4136), .B(n4137), .Z(y[206]) );
  NAND U5554 ( .A(n3862), .B(m[206]), .Z(n4137) );
  NAND U5555 ( .A(n3863), .B(creg[206]), .Z(n4136) );
  NAND U5556 ( .A(n4138), .B(n4139), .Z(y[205]) );
  NAND U5557 ( .A(n3862), .B(m[205]), .Z(n4139) );
  NAND U5558 ( .A(n3863), .B(creg[205]), .Z(n4138) );
  NAND U5559 ( .A(n4140), .B(n4141), .Z(y[204]) );
  NAND U5560 ( .A(n3862), .B(m[204]), .Z(n4141) );
  NAND U5561 ( .A(n3863), .B(creg[204]), .Z(n4140) );
  NAND U5562 ( .A(n4142), .B(n4143), .Z(y[203]) );
  NAND U5563 ( .A(n3862), .B(m[203]), .Z(n4143) );
  NAND U5564 ( .A(n3863), .B(creg[203]), .Z(n4142) );
  NAND U5565 ( .A(n4144), .B(n4145), .Z(y[202]) );
  NAND U5566 ( .A(n3862), .B(m[202]), .Z(n4145) );
  NAND U5567 ( .A(n3863), .B(creg[202]), .Z(n4144) );
  NAND U5568 ( .A(n4146), .B(n4147), .Z(y[201]) );
  NAND U5569 ( .A(n3862), .B(m[201]), .Z(n4147) );
  NAND U5570 ( .A(n3863), .B(creg[201]), .Z(n4146) );
  NAND U5571 ( .A(n4148), .B(n4149), .Z(y[200]) );
  NAND U5572 ( .A(n3862), .B(m[200]), .Z(n4149) );
  NAND U5573 ( .A(n3863), .B(creg[200]), .Z(n4148) );
  NAND U5574 ( .A(n4150), .B(n4151), .Z(y[1]) );
  NAND U5575 ( .A(n3862), .B(m[1]), .Z(n4151) );
  NAND U5576 ( .A(n3863), .B(creg[1]), .Z(n4150) );
  NAND U5577 ( .A(n4152), .B(n4153), .Z(y[19]) );
  NAND U5578 ( .A(n3862), .B(m[19]), .Z(n4153) );
  NAND U5579 ( .A(n3863), .B(creg[19]), .Z(n4152) );
  NAND U5580 ( .A(n4154), .B(n4155), .Z(y[199]) );
  NAND U5581 ( .A(n3862), .B(m[199]), .Z(n4155) );
  NAND U5582 ( .A(n3863), .B(creg[199]), .Z(n4154) );
  NAND U5583 ( .A(n4156), .B(n4157), .Z(y[198]) );
  NAND U5584 ( .A(n3862), .B(m[198]), .Z(n4157) );
  NAND U5585 ( .A(n3863), .B(creg[198]), .Z(n4156) );
  NAND U5586 ( .A(n4158), .B(n4159), .Z(y[197]) );
  NAND U5587 ( .A(n3862), .B(m[197]), .Z(n4159) );
  NAND U5588 ( .A(n3863), .B(creg[197]), .Z(n4158) );
  NAND U5589 ( .A(n4160), .B(n4161), .Z(y[196]) );
  NAND U5590 ( .A(n3862), .B(m[196]), .Z(n4161) );
  NAND U5591 ( .A(n3863), .B(creg[196]), .Z(n4160) );
  NAND U5592 ( .A(n4162), .B(n4163), .Z(y[195]) );
  NAND U5593 ( .A(n3862), .B(m[195]), .Z(n4163) );
  NAND U5594 ( .A(n3863), .B(creg[195]), .Z(n4162) );
  NAND U5595 ( .A(n4164), .B(n4165), .Z(y[194]) );
  NAND U5596 ( .A(n3862), .B(m[194]), .Z(n4165) );
  NAND U5597 ( .A(n3863), .B(creg[194]), .Z(n4164) );
  NAND U5598 ( .A(n4166), .B(n4167), .Z(y[193]) );
  NAND U5599 ( .A(n3862), .B(m[193]), .Z(n4167) );
  NAND U5600 ( .A(n3863), .B(creg[193]), .Z(n4166) );
  NAND U5601 ( .A(n4168), .B(n4169), .Z(y[192]) );
  NAND U5602 ( .A(n3862), .B(m[192]), .Z(n4169) );
  NAND U5603 ( .A(n3863), .B(creg[192]), .Z(n4168) );
  NAND U5604 ( .A(n4170), .B(n4171), .Z(y[191]) );
  NAND U5605 ( .A(n3862), .B(m[191]), .Z(n4171) );
  NAND U5606 ( .A(n3863), .B(creg[191]), .Z(n4170) );
  NAND U5607 ( .A(n4172), .B(n4173), .Z(y[190]) );
  NAND U5608 ( .A(n3862), .B(m[190]), .Z(n4173) );
  NAND U5609 ( .A(n3863), .B(creg[190]), .Z(n4172) );
  NAND U5610 ( .A(n4174), .B(n4175), .Z(y[18]) );
  NAND U5611 ( .A(n3862), .B(m[18]), .Z(n4175) );
  NAND U5612 ( .A(n3863), .B(creg[18]), .Z(n4174) );
  NAND U5613 ( .A(n4176), .B(n4177), .Z(y[189]) );
  NAND U5614 ( .A(n3862), .B(m[189]), .Z(n4177) );
  NAND U5615 ( .A(n3863), .B(creg[189]), .Z(n4176) );
  NAND U5616 ( .A(n4178), .B(n4179), .Z(y[188]) );
  NAND U5617 ( .A(n3862), .B(m[188]), .Z(n4179) );
  NAND U5618 ( .A(n3863), .B(creg[188]), .Z(n4178) );
  NAND U5619 ( .A(n4180), .B(n4181), .Z(y[187]) );
  NAND U5620 ( .A(n3862), .B(m[187]), .Z(n4181) );
  NAND U5621 ( .A(n3863), .B(creg[187]), .Z(n4180) );
  NAND U5622 ( .A(n4182), .B(n4183), .Z(y[186]) );
  NAND U5623 ( .A(n3862), .B(m[186]), .Z(n4183) );
  NAND U5624 ( .A(n3863), .B(creg[186]), .Z(n4182) );
  NAND U5625 ( .A(n4184), .B(n4185), .Z(y[185]) );
  NAND U5626 ( .A(n3862), .B(m[185]), .Z(n4185) );
  NAND U5627 ( .A(n3863), .B(creg[185]), .Z(n4184) );
  NAND U5628 ( .A(n4186), .B(n4187), .Z(y[184]) );
  NAND U5629 ( .A(n3862), .B(m[184]), .Z(n4187) );
  NAND U5630 ( .A(n3863), .B(creg[184]), .Z(n4186) );
  NAND U5631 ( .A(n4188), .B(n4189), .Z(y[183]) );
  NAND U5632 ( .A(n3862), .B(m[183]), .Z(n4189) );
  NAND U5633 ( .A(n3863), .B(creg[183]), .Z(n4188) );
  NAND U5634 ( .A(n4190), .B(n4191), .Z(y[182]) );
  NAND U5635 ( .A(n3862), .B(m[182]), .Z(n4191) );
  NAND U5636 ( .A(n3863), .B(creg[182]), .Z(n4190) );
  NAND U5637 ( .A(n4192), .B(n4193), .Z(y[181]) );
  NAND U5638 ( .A(n3862), .B(m[181]), .Z(n4193) );
  NAND U5639 ( .A(n3863), .B(creg[181]), .Z(n4192) );
  NAND U5640 ( .A(n4194), .B(n4195), .Z(y[180]) );
  NAND U5641 ( .A(n3862), .B(m[180]), .Z(n4195) );
  NAND U5642 ( .A(n3863), .B(creg[180]), .Z(n4194) );
  NAND U5643 ( .A(n4196), .B(n4197), .Z(y[17]) );
  NAND U5644 ( .A(n3862), .B(m[17]), .Z(n4197) );
  NAND U5645 ( .A(n3863), .B(creg[17]), .Z(n4196) );
  NAND U5646 ( .A(n4198), .B(n4199), .Z(y[179]) );
  NAND U5647 ( .A(n3862), .B(m[179]), .Z(n4199) );
  NAND U5648 ( .A(n3863), .B(creg[179]), .Z(n4198) );
  NAND U5649 ( .A(n4200), .B(n4201), .Z(y[178]) );
  NAND U5650 ( .A(n3862), .B(m[178]), .Z(n4201) );
  NAND U5651 ( .A(n3863), .B(creg[178]), .Z(n4200) );
  NAND U5652 ( .A(n4202), .B(n4203), .Z(y[177]) );
  NAND U5653 ( .A(n3862), .B(m[177]), .Z(n4203) );
  NAND U5654 ( .A(n3863), .B(creg[177]), .Z(n4202) );
  NAND U5655 ( .A(n4204), .B(n4205), .Z(y[176]) );
  NAND U5656 ( .A(n3862), .B(m[176]), .Z(n4205) );
  NAND U5657 ( .A(n3863), .B(creg[176]), .Z(n4204) );
  NAND U5658 ( .A(n4206), .B(n4207), .Z(y[175]) );
  NAND U5659 ( .A(n3862), .B(m[175]), .Z(n4207) );
  NAND U5660 ( .A(n3863), .B(creg[175]), .Z(n4206) );
  NAND U5661 ( .A(n4208), .B(n4209), .Z(y[174]) );
  NAND U5662 ( .A(n3862), .B(m[174]), .Z(n4209) );
  NAND U5663 ( .A(n3863), .B(creg[174]), .Z(n4208) );
  NAND U5664 ( .A(n4210), .B(n4211), .Z(y[173]) );
  NAND U5665 ( .A(n3862), .B(m[173]), .Z(n4211) );
  NAND U5666 ( .A(n3863), .B(creg[173]), .Z(n4210) );
  NAND U5667 ( .A(n4212), .B(n4213), .Z(y[172]) );
  NAND U5668 ( .A(n3862), .B(m[172]), .Z(n4213) );
  NAND U5669 ( .A(n3863), .B(creg[172]), .Z(n4212) );
  NAND U5670 ( .A(n4214), .B(n4215), .Z(y[171]) );
  NAND U5671 ( .A(n3862), .B(m[171]), .Z(n4215) );
  NAND U5672 ( .A(n3863), .B(creg[171]), .Z(n4214) );
  NAND U5673 ( .A(n4216), .B(n4217), .Z(y[170]) );
  NAND U5674 ( .A(n3862), .B(m[170]), .Z(n4217) );
  NAND U5675 ( .A(n3863), .B(creg[170]), .Z(n4216) );
  NAND U5676 ( .A(n4218), .B(n4219), .Z(y[16]) );
  NAND U5677 ( .A(n3862), .B(m[16]), .Z(n4219) );
  NAND U5678 ( .A(n3863), .B(creg[16]), .Z(n4218) );
  NAND U5679 ( .A(n4220), .B(n4221), .Z(y[169]) );
  NAND U5680 ( .A(n3862), .B(m[169]), .Z(n4221) );
  NAND U5681 ( .A(n3863), .B(creg[169]), .Z(n4220) );
  NAND U5682 ( .A(n4222), .B(n4223), .Z(y[168]) );
  NAND U5683 ( .A(n3862), .B(m[168]), .Z(n4223) );
  NAND U5684 ( .A(n3863), .B(creg[168]), .Z(n4222) );
  NAND U5685 ( .A(n4224), .B(n4225), .Z(y[167]) );
  NAND U5686 ( .A(n3862), .B(m[167]), .Z(n4225) );
  NAND U5687 ( .A(n3863), .B(creg[167]), .Z(n4224) );
  NAND U5688 ( .A(n4226), .B(n4227), .Z(y[166]) );
  NAND U5689 ( .A(n3862), .B(m[166]), .Z(n4227) );
  NAND U5690 ( .A(n3863), .B(creg[166]), .Z(n4226) );
  NAND U5691 ( .A(n4228), .B(n4229), .Z(y[165]) );
  NAND U5692 ( .A(n3862), .B(m[165]), .Z(n4229) );
  NAND U5693 ( .A(n3863), .B(creg[165]), .Z(n4228) );
  NAND U5694 ( .A(n4230), .B(n4231), .Z(y[164]) );
  NAND U5695 ( .A(n3862), .B(m[164]), .Z(n4231) );
  NAND U5696 ( .A(n3863), .B(creg[164]), .Z(n4230) );
  NAND U5697 ( .A(n4232), .B(n4233), .Z(y[163]) );
  NAND U5698 ( .A(n3862), .B(m[163]), .Z(n4233) );
  NAND U5699 ( .A(n3863), .B(creg[163]), .Z(n4232) );
  NAND U5700 ( .A(n4234), .B(n4235), .Z(y[162]) );
  NAND U5701 ( .A(n3862), .B(m[162]), .Z(n4235) );
  NAND U5702 ( .A(n3863), .B(creg[162]), .Z(n4234) );
  NAND U5703 ( .A(n4236), .B(n4237), .Z(y[161]) );
  NAND U5704 ( .A(n3862), .B(m[161]), .Z(n4237) );
  NAND U5705 ( .A(n3863), .B(creg[161]), .Z(n4236) );
  NAND U5706 ( .A(n4238), .B(n4239), .Z(y[160]) );
  NAND U5707 ( .A(n3862), .B(m[160]), .Z(n4239) );
  NAND U5708 ( .A(n3863), .B(creg[160]), .Z(n4238) );
  NAND U5709 ( .A(n4240), .B(n4241), .Z(y[15]) );
  NAND U5710 ( .A(n3862), .B(m[15]), .Z(n4241) );
  NAND U5711 ( .A(n3863), .B(creg[15]), .Z(n4240) );
  NAND U5712 ( .A(n4242), .B(n4243), .Z(y[159]) );
  NAND U5713 ( .A(n3862), .B(m[159]), .Z(n4243) );
  NAND U5714 ( .A(n3863), .B(creg[159]), .Z(n4242) );
  NAND U5715 ( .A(n4244), .B(n4245), .Z(y[158]) );
  NAND U5716 ( .A(n3862), .B(m[158]), .Z(n4245) );
  NAND U5717 ( .A(n3863), .B(creg[158]), .Z(n4244) );
  NAND U5718 ( .A(n4246), .B(n4247), .Z(y[157]) );
  NAND U5719 ( .A(n3862), .B(m[157]), .Z(n4247) );
  NAND U5720 ( .A(n3863), .B(creg[157]), .Z(n4246) );
  NAND U5721 ( .A(n4248), .B(n4249), .Z(y[156]) );
  NAND U5722 ( .A(n3862), .B(m[156]), .Z(n4249) );
  NAND U5723 ( .A(n3863), .B(creg[156]), .Z(n4248) );
  NAND U5724 ( .A(n4250), .B(n4251), .Z(y[155]) );
  NAND U5725 ( .A(n3862), .B(m[155]), .Z(n4251) );
  NAND U5726 ( .A(n3863), .B(creg[155]), .Z(n4250) );
  NAND U5727 ( .A(n4252), .B(n4253), .Z(y[154]) );
  NAND U5728 ( .A(n3862), .B(m[154]), .Z(n4253) );
  NAND U5729 ( .A(n3863), .B(creg[154]), .Z(n4252) );
  NAND U5730 ( .A(n4254), .B(n4255), .Z(y[153]) );
  NAND U5731 ( .A(n3862), .B(m[153]), .Z(n4255) );
  NAND U5732 ( .A(n3863), .B(creg[153]), .Z(n4254) );
  NAND U5733 ( .A(n4256), .B(n4257), .Z(y[152]) );
  NAND U5734 ( .A(n3862), .B(m[152]), .Z(n4257) );
  NAND U5735 ( .A(n3863), .B(creg[152]), .Z(n4256) );
  NAND U5736 ( .A(n4258), .B(n4259), .Z(y[151]) );
  NAND U5737 ( .A(n3862), .B(m[151]), .Z(n4259) );
  NAND U5738 ( .A(n3863), .B(creg[151]), .Z(n4258) );
  NAND U5739 ( .A(n4260), .B(n4261), .Z(y[150]) );
  NAND U5740 ( .A(n3862), .B(m[150]), .Z(n4261) );
  NAND U5741 ( .A(n3863), .B(creg[150]), .Z(n4260) );
  NAND U5742 ( .A(n4262), .B(n4263), .Z(y[14]) );
  NAND U5743 ( .A(n3862), .B(m[14]), .Z(n4263) );
  NAND U5744 ( .A(n3863), .B(creg[14]), .Z(n4262) );
  NAND U5745 ( .A(n4264), .B(n4265), .Z(y[149]) );
  NAND U5746 ( .A(n3862), .B(m[149]), .Z(n4265) );
  NAND U5747 ( .A(n3863), .B(creg[149]), .Z(n4264) );
  NAND U5748 ( .A(n4266), .B(n4267), .Z(y[148]) );
  NAND U5749 ( .A(n3862), .B(m[148]), .Z(n4267) );
  NAND U5750 ( .A(n3863), .B(creg[148]), .Z(n4266) );
  NAND U5751 ( .A(n4268), .B(n4269), .Z(y[147]) );
  NAND U5752 ( .A(n3862), .B(m[147]), .Z(n4269) );
  NAND U5753 ( .A(n3863), .B(creg[147]), .Z(n4268) );
  NAND U5754 ( .A(n4270), .B(n4271), .Z(y[146]) );
  NAND U5755 ( .A(n3862), .B(m[146]), .Z(n4271) );
  NAND U5756 ( .A(n3863), .B(creg[146]), .Z(n4270) );
  NAND U5757 ( .A(n4272), .B(n4273), .Z(y[145]) );
  NAND U5758 ( .A(n3862), .B(m[145]), .Z(n4273) );
  NAND U5759 ( .A(n3863), .B(creg[145]), .Z(n4272) );
  NAND U5760 ( .A(n4274), .B(n4275), .Z(y[144]) );
  NAND U5761 ( .A(n3862), .B(m[144]), .Z(n4275) );
  NAND U5762 ( .A(n3863), .B(creg[144]), .Z(n4274) );
  NAND U5763 ( .A(n4276), .B(n4277), .Z(y[143]) );
  NAND U5764 ( .A(n3862), .B(m[143]), .Z(n4277) );
  NAND U5765 ( .A(n3863), .B(creg[143]), .Z(n4276) );
  NAND U5766 ( .A(n4278), .B(n4279), .Z(y[142]) );
  NAND U5767 ( .A(n3862), .B(m[142]), .Z(n4279) );
  NAND U5768 ( .A(n3863), .B(creg[142]), .Z(n4278) );
  NAND U5769 ( .A(n4280), .B(n4281), .Z(y[141]) );
  NAND U5770 ( .A(n3862), .B(m[141]), .Z(n4281) );
  NAND U5771 ( .A(n3863), .B(creg[141]), .Z(n4280) );
  NAND U5772 ( .A(n4282), .B(n4283), .Z(y[140]) );
  NAND U5773 ( .A(n3862), .B(m[140]), .Z(n4283) );
  NAND U5774 ( .A(n3863), .B(creg[140]), .Z(n4282) );
  NAND U5775 ( .A(n4284), .B(n4285), .Z(y[13]) );
  NAND U5776 ( .A(n3862), .B(m[13]), .Z(n4285) );
  NAND U5777 ( .A(n3863), .B(creg[13]), .Z(n4284) );
  NAND U5778 ( .A(n4286), .B(n4287), .Z(y[139]) );
  NAND U5779 ( .A(n3862), .B(m[139]), .Z(n4287) );
  NAND U5780 ( .A(n3863), .B(creg[139]), .Z(n4286) );
  NAND U5781 ( .A(n4288), .B(n4289), .Z(y[138]) );
  NAND U5782 ( .A(n3862), .B(m[138]), .Z(n4289) );
  NAND U5783 ( .A(n3863), .B(creg[138]), .Z(n4288) );
  NAND U5784 ( .A(n4290), .B(n4291), .Z(y[137]) );
  NAND U5785 ( .A(n3862), .B(m[137]), .Z(n4291) );
  NAND U5786 ( .A(n3863), .B(creg[137]), .Z(n4290) );
  NAND U5787 ( .A(n4292), .B(n4293), .Z(y[136]) );
  NAND U5788 ( .A(n3862), .B(m[136]), .Z(n4293) );
  NAND U5789 ( .A(n3863), .B(creg[136]), .Z(n4292) );
  NAND U5790 ( .A(n4294), .B(n4295), .Z(y[135]) );
  NAND U5791 ( .A(n3862), .B(m[135]), .Z(n4295) );
  NAND U5792 ( .A(n3863), .B(creg[135]), .Z(n4294) );
  NAND U5793 ( .A(n4296), .B(n4297), .Z(y[134]) );
  NAND U5794 ( .A(n3862), .B(m[134]), .Z(n4297) );
  NAND U5795 ( .A(n3863), .B(creg[134]), .Z(n4296) );
  NAND U5796 ( .A(n4298), .B(n4299), .Z(y[133]) );
  NAND U5797 ( .A(n3862), .B(m[133]), .Z(n4299) );
  NAND U5798 ( .A(n3863), .B(creg[133]), .Z(n4298) );
  NAND U5799 ( .A(n4300), .B(n4301), .Z(y[132]) );
  NAND U5800 ( .A(n3862), .B(m[132]), .Z(n4301) );
  NAND U5801 ( .A(n3863), .B(creg[132]), .Z(n4300) );
  NAND U5802 ( .A(n4302), .B(n4303), .Z(y[131]) );
  NAND U5803 ( .A(n3862), .B(m[131]), .Z(n4303) );
  NAND U5804 ( .A(n3863), .B(creg[131]), .Z(n4302) );
  NAND U5805 ( .A(n4304), .B(n4305), .Z(y[130]) );
  NAND U5806 ( .A(n3862), .B(m[130]), .Z(n4305) );
  NAND U5807 ( .A(n3863), .B(creg[130]), .Z(n4304) );
  NAND U5808 ( .A(n4306), .B(n4307), .Z(y[12]) );
  NAND U5809 ( .A(n3862), .B(m[12]), .Z(n4307) );
  NAND U5810 ( .A(n3863), .B(creg[12]), .Z(n4306) );
  NAND U5811 ( .A(n4308), .B(n4309), .Z(y[129]) );
  NAND U5812 ( .A(n3862), .B(m[129]), .Z(n4309) );
  NAND U5813 ( .A(n3863), .B(creg[129]), .Z(n4308) );
  NAND U5814 ( .A(n4310), .B(n4311), .Z(y[128]) );
  NAND U5815 ( .A(n3862), .B(m[128]), .Z(n4311) );
  NAND U5816 ( .A(n3863), .B(creg[128]), .Z(n4310) );
  NAND U5817 ( .A(n4312), .B(n4313), .Z(y[127]) );
  NAND U5818 ( .A(n3862), .B(m[127]), .Z(n4313) );
  NAND U5819 ( .A(n3863), .B(creg[127]), .Z(n4312) );
  NAND U5820 ( .A(n4314), .B(n4315), .Z(y[126]) );
  NAND U5821 ( .A(n3862), .B(m[126]), .Z(n4315) );
  NAND U5822 ( .A(n3863), .B(creg[126]), .Z(n4314) );
  NAND U5823 ( .A(n4316), .B(n4317), .Z(y[125]) );
  NAND U5824 ( .A(n3862), .B(m[125]), .Z(n4317) );
  NAND U5825 ( .A(n3863), .B(creg[125]), .Z(n4316) );
  NAND U5826 ( .A(n4318), .B(n4319), .Z(y[124]) );
  NAND U5827 ( .A(n3862), .B(m[124]), .Z(n4319) );
  NAND U5828 ( .A(n3863), .B(creg[124]), .Z(n4318) );
  NAND U5829 ( .A(n4320), .B(n4321), .Z(y[123]) );
  NAND U5830 ( .A(n3862), .B(m[123]), .Z(n4321) );
  NAND U5831 ( .A(n3863), .B(creg[123]), .Z(n4320) );
  NAND U5832 ( .A(n4322), .B(n4323), .Z(y[122]) );
  NAND U5833 ( .A(n3862), .B(m[122]), .Z(n4323) );
  NAND U5834 ( .A(n3863), .B(creg[122]), .Z(n4322) );
  NAND U5835 ( .A(n4324), .B(n4325), .Z(y[121]) );
  NAND U5836 ( .A(n3862), .B(m[121]), .Z(n4325) );
  NAND U5837 ( .A(n3863), .B(creg[121]), .Z(n4324) );
  NAND U5838 ( .A(n4326), .B(n4327), .Z(y[120]) );
  NAND U5839 ( .A(n3862), .B(m[120]), .Z(n4327) );
  NAND U5840 ( .A(n3863), .B(creg[120]), .Z(n4326) );
  NAND U5841 ( .A(n4328), .B(n4329), .Z(y[11]) );
  NAND U5842 ( .A(n3862), .B(m[11]), .Z(n4329) );
  NAND U5843 ( .A(n3863), .B(creg[11]), .Z(n4328) );
  NAND U5844 ( .A(n4330), .B(n4331), .Z(y[119]) );
  NAND U5845 ( .A(n3862), .B(m[119]), .Z(n4331) );
  NAND U5846 ( .A(n3863), .B(creg[119]), .Z(n4330) );
  NAND U5847 ( .A(n4332), .B(n4333), .Z(y[118]) );
  NAND U5848 ( .A(n3862), .B(m[118]), .Z(n4333) );
  NAND U5849 ( .A(n3863), .B(creg[118]), .Z(n4332) );
  NAND U5850 ( .A(n4334), .B(n4335), .Z(y[117]) );
  NAND U5851 ( .A(n3862), .B(m[117]), .Z(n4335) );
  NAND U5852 ( .A(n3863), .B(creg[117]), .Z(n4334) );
  NAND U5853 ( .A(n4336), .B(n4337), .Z(y[116]) );
  NAND U5854 ( .A(n3862), .B(m[116]), .Z(n4337) );
  NAND U5855 ( .A(n3863), .B(creg[116]), .Z(n4336) );
  NAND U5856 ( .A(n4338), .B(n4339), .Z(y[115]) );
  NAND U5857 ( .A(n3862), .B(m[115]), .Z(n4339) );
  NAND U5858 ( .A(n3863), .B(creg[115]), .Z(n4338) );
  NAND U5859 ( .A(n4340), .B(n4341), .Z(y[114]) );
  NAND U5860 ( .A(n3862), .B(m[114]), .Z(n4341) );
  NAND U5861 ( .A(n3863), .B(creg[114]), .Z(n4340) );
  NAND U5862 ( .A(n4342), .B(n4343), .Z(y[113]) );
  NAND U5863 ( .A(n3862), .B(m[113]), .Z(n4343) );
  NAND U5864 ( .A(n3863), .B(creg[113]), .Z(n4342) );
  NAND U5865 ( .A(n4344), .B(n4345), .Z(y[112]) );
  NAND U5866 ( .A(n3862), .B(m[112]), .Z(n4345) );
  NAND U5867 ( .A(n3863), .B(creg[112]), .Z(n4344) );
  NAND U5868 ( .A(n4346), .B(n4347), .Z(y[111]) );
  NAND U5869 ( .A(n3862), .B(m[111]), .Z(n4347) );
  NAND U5870 ( .A(n3863), .B(creg[111]), .Z(n4346) );
  NAND U5871 ( .A(n4348), .B(n4349), .Z(y[110]) );
  NAND U5872 ( .A(n3862), .B(m[110]), .Z(n4349) );
  NAND U5873 ( .A(n3863), .B(creg[110]), .Z(n4348) );
  NAND U5874 ( .A(n4350), .B(n4351), .Z(y[10]) );
  NAND U5875 ( .A(n3862), .B(m[10]), .Z(n4351) );
  NAND U5876 ( .A(n3863), .B(creg[10]), .Z(n4350) );
  NAND U5877 ( .A(n4352), .B(n4353), .Z(y[109]) );
  NAND U5878 ( .A(n3862), .B(m[109]), .Z(n4353) );
  NAND U5879 ( .A(n3863), .B(creg[109]), .Z(n4352) );
  NAND U5880 ( .A(n4354), .B(n4355), .Z(y[108]) );
  NAND U5881 ( .A(n3862), .B(m[108]), .Z(n4355) );
  NAND U5882 ( .A(n3863), .B(creg[108]), .Z(n4354) );
  NAND U5883 ( .A(n4356), .B(n4357), .Z(y[107]) );
  NAND U5884 ( .A(n3862), .B(m[107]), .Z(n4357) );
  NAND U5885 ( .A(n3863), .B(creg[107]), .Z(n4356) );
  NAND U5886 ( .A(n4358), .B(n4359), .Z(y[106]) );
  NAND U5887 ( .A(n3862), .B(m[106]), .Z(n4359) );
  NAND U5888 ( .A(n3863), .B(creg[106]), .Z(n4358) );
  NAND U5889 ( .A(n4360), .B(n4361), .Z(y[105]) );
  NAND U5890 ( .A(n3862), .B(m[105]), .Z(n4361) );
  NAND U5891 ( .A(n3863), .B(creg[105]), .Z(n4360) );
  NAND U5892 ( .A(n4362), .B(n4363), .Z(y[104]) );
  NAND U5893 ( .A(n3862), .B(m[104]), .Z(n4363) );
  NAND U5894 ( .A(n3863), .B(creg[104]), .Z(n4362) );
  NAND U5895 ( .A(n4364), .B(n4365), .Z(y[103]) );
  NAND U5896 ( .A(n3862), .B(m[103]), .Z(n4365) );
  NAND U5897 ( .A(n3863), .B(creg[103]), .Z(n4364) );
  NAND U5898 ( .A(n4366), .B(n4367), .Z(y[102]) );
  NAND U5899 ( .A(n3862), .B(m[102]), .Z(n4367) );
  NAND U5900 ( .A(n3863), .B(creg[102]), .Z(n4366) );
  NAND U5901 ( .A(n4368), .B(n4369), .Z(y[101]) );
  NAND U5902 ( .A(n3862), .B(m[101]), .Z(n4369) );
  NAND U5903 ( .A(n3863), .B(creg[101]), .Z(n4368) );
  NAND U5904 ( .A(n4370), .B(n4371), .Z(y[100]) );
  NAND U5905 ( .A(n3862), .B(m[100]), .Z(n4371) );
  NAND U5906 ( .A(n3863), .B(creg[100]), .Z(n4370) );
  NAND U5907 ( .A(n4372), .B(n4373), .Z(y[0]) );
  NAND U5908 ( .A(n3862), .B(m[0]), .Z(n4373) );
  NAND U5909 ( .A(n3863), .B(creg[0]), .Z(n4372) );
  NAND U5910 ( .A(n4374), .B(n4375), .Z(x[9]) );
  NAND U5911 ( .A(creg[9]), .B(init), .Z(n4374) );
  NAND U5912 ( .A(n4376), .B(n4377), .Z(x[99]) );
  NAND U5913 ( .A(creg[99]), .B(init), .Z(n4376) );
  NAND U5914 ( .A(n4378), .B(n4379), .Z(x[98]) );
  NAND U5915 ( .A(creg[98]), .B(init), .Z(n4378) );
  NAND U5916 ( .A(n4380), .B(n4381), .Z(x[97]) );
  NAND U5917 ( .A(creg[97]), .B(init), .Z(n4380) );
  NAND U5918 ( .A(n4382), .B(n4383), .Z(x[96]) );
  NAND U5919 ( .A(creg[96]), .B(init), .Z(n4382) );
  NAND U5920 ( .A(n4384), .B(n4385), .Z(x[95]) );
  NAND U5921 ( .A(creg[95]), .B(init), .Z(n4384) );
  NAND U5922 ( .A(n4386), .B(n4387), .Z(x[94]) );
  NAND U5923 ( .A(creg[94]), .B(init), .Z(n4386) );
  NAND U5924 ( .A(n4388), .B(n4389), .Z(x[93]) );
  NAND U5925 ( .A(creg[93]), .B(init), .Z(n4388) );
  NAND U5926 ( .A(n4390), .B(n4391), .Z(x[92]) );
  NAND U5927 ( .A(creg[92]), .B(init), .Z(n4390) );
  NAND U5928 ( .A(n4392), .B(n4393), .Z(x[91]) );
  NAND U5929 ( .A(creg[91]), .B(init), .Z(n4392) );
  NAND U5930 ( .A(n4394), .B(n4395), .Z(x[90]) );
  NAND U5931 ( .A(creg[90]), .B(init), .Z(n4394) );
  NAND U5932 ( .A(n4396), .B(n4397), .Z(x[8]) );
  NAND U5933 ( .A(creg[8]), .B(init), .Z(n4396) );
  NAND U5934 ( .A(n4398), .B(n4399), .Z(x[89]) );
  NAND U5935 ( .A(creg[89]), .B(init), .Z(n4398) );
  NAND U5936 ( .A(n4400), .B(n4401), .Z(x[88]) );
  NAND U5937 ( .A(creg[88]), .B(init), .Z(n4400) );
  NAND U5938 ( .A(n4402), .B(n4403), .Z(x[87]) );
  NAND U5939 ( .A(creg[87]), .B(init), .Z(n4402) );
  NAND U5940 ( .A(n4404), .B(n4405), .Z(x[86]) );
  NAND U5941 ( .A(creg[86]), .B(init), .Z(n4404) );
  NAND U5942 ( .A(n4406), .B(n4407), .Z(x[85]) );
  NAND U5943 ( .A(creg[85]), .B(init), .Z(n4406) );
  NAND U5944 ( .A(n4408), .B(n4409), .Z(x[84]) );
  NAND U5945 ( .A(creg[84]), .B(init), .Z(n4408) );
  NAND U5946 ( .A(n4410), .B(n4411), .Z(x[83]) );
  NAND U5947 ( .A(creg[83]), .B(init), .Z(n4410) );
  NAND U5948 ( .A(n4412), .B(n4413), .Z(x[82]) );
  NAND U5949 ( .A(creg[82]), .B(init), .Z(n4412) );
  NAND U5950 ( .A(n4414), .B(n4415), .Z(x[81]) );
  NAND U5951 ( .A(creg[81]), .B(init), .Z(n4414) );
  NAND U5952 ( .A(n4416), .B(n4417), .Z(x[80]) );
  NAND U5953 ( .A(creg[80]), .B(init), .Z(n4416) );
  NAND U5954 ( .A(n4418), .B(n4419), .Z(x[7]) );
  NAND U5955 ( .A(creg[7]), .B(init), .Z(n4418) );
  NAND U5956 ( .A(n4420), .B(n4421), .Z(x[79]) );
  NAND U5957 ( .A(creg[79]), .B(init), .Z(n4420) );
  NAND U5958 ( .A(n4422), .B(n4423), .Z(x[78]) );
  NAND U5959 ( .A(creg[78]), .B(init), .Z(n4422) );
  NAND U5960 ( .A(n4424), .B(n4425), .Z(x[77]) );
  NAND U5961 ( .A(creg[77]), .B(init), .Z(n4424) );
  NAND U5962 ( .A(n4426), .B(n4427), .Z(x[76]) );
  NAND U5963 ( .A(creg[76]), .B(init), .Z(n4426) );
  NAND U5964 ( .A(n4428), .B(n4429), .Z(x[75]) );
  NAND U5965 ( .A(creg[75]), .B(init), .Z(n4428) );
  NAND U5966 ( .A(n4430), .B(n4431), .Z(x[74]) );
  NAND U5967 ( .A(creg[74]), .B(init), .Z(n4430) );
  NAND U5968 ( .A(n4432), .B(n4433), .Z(x[73]) );
  NAND U5969 ( .A(creg[73]), .B(init), .Z(n4432) );
  NAND U5970 ( .A(n4434), .B(n4435), .Z(x[72]) );
  NAND U5971 ( .A(creg[72]), .B(init), .Z(n4434) );
  NAND U5972 ( .A(n4436), .B(n4437), .Z(x[71]) );
  NAND U5973 ( .A(creg[71]), .B(init), .Z(n4436) );
  NAND U5974 ( .A(n4438), .B(n4439), .Z(x[70]) );
  NAND U5975 ( .A(creg[70]), .B(init), .Z(n4438) );
  NAND U5976 ( .A(n4440), .B(n4441), .Z(x[6]) );
  NAND U5977 ( .A(creg[6]), .B(init), .Z(n4440) );
  NAND U5978 ( .A(n4442), .B(n4443), .Z(x[69]) );
  NAND U5979 ( .A(creg[69]), .B(init), .Z(n4442) );
  NAND U5980 ( .A(n4444), .B(n4445), .Z(x[68]) );
  NAND U5981 ( .A(creg[68]), .B(init), .Z(n4444) );
  NAND U5982 ( .A(n4446), .B(n4447), .Z(x[67]) );
  NAND U5983 ( .A(creg[67]), .B(init), .Z(n4446) );
  NAND U5984 ( .A(n4448), .B(n4449), .Z(x[66]) );
  NAND U5985 ( .A(creg[66]), .B(init), .Z(n4448) );
  NAND U5986 ( .A(n4450), .B(n4451), .Z(x[65]) );
  NAND U5987 ( .A(creg[65]), .B(init), .Z(n4450) );
  NAND U5988 ( .A(n4452), .B(n4453), .Z(x[64]) );
  NAND U5989 ( .A(creg[64]), .B(init), .Z(n4452) );
  NAND U5990 ( .A(n4454), .B(n4455), .Z(x[63]) );
  NAND U5991 ( .A(creg[63]), .B(init), .Z(n4454) );
  NAND U5992 ( .A(n4456), .B(n4457), .Z(x[62]) );
  NAND U5993 ( .A(creg[62]), .B(init), .Z(n4456) );
  NAND U5994 ( .A(n4458), .B(n4459), .Z(x[61]) );
  NAND U5995 ( .A(creg[61]), .B(init), .Z(n4458) );
  NAND U5996 ( .A(n4460), .B(n4461), .Z(x[60]) );
  NAND U5997 ( .A(creg[60]), .B(init), .Z(n4460) );
  NAND U5998 ( .A(n4462), .B(n4463), .Z(x[5]) );
  NAND U5999 ( .A(creg[5]), .B(init), .Z(n4462) );
  NAND U6000 ( .A(n4464), .B(n4465), .Z(x[59]) );
  NAND U6001 ( .A(creg[59]), .B(init), .Z(n4464) );
  NAND U6002 ( .A(n4466), .B(n4467), .Z(x[58]) );
  NAND U6003 ( .A(creg[58]), .B(init), .Z(n4466) );
  NAND U6004 ( .A(n4468), .B(n4469), .Z(x[57]) );
  NAND U6005 ( .A(creg[57]), .B(init), .Z(n4468) );
  NAND U6006 ( .A(n4470), .B(n4471), .Z(x[56]) );
  NAND U6007 ( .A(creg[56]), .B(init), .Z(n4470) );
  NAND U6008 ( .A(n4472), .B(n4473), .Z(x[55]) );
  NAND U6009 ( .A(creg[55]), .B(init), .Z(n4472) );
  NAND U6010 ( .A(n4474), .B(n4475), .Z(x[54]) );
  NAND U6011 ( .A(creg[54]), .B(init), .Z(n4474) );
  NAND U6012 ( .A(n4476), .B(n4477), .Z(x[53]) );
  NAND U6013 ( .A(creg[53]), .B(init), .Z(n4476) );
  NAND U6014 ( .A(n4478), .B(n4479), .Z(x[52]) );
  NAND U6015 ( .A(creg[52]), .B(init), .Z(n4478) );
  NAND U6016 ( .A(n4480), .B(n4481), .Z(x[51]) );
  NAND U6017 ( .A(creg[51]), .B(init), .Z(n4480) );
  NAND U6018 ( .A(n4482), .B(n4483), .Z(x[50]) );
  NAND U6019 ( .A(creg[50]), .B(init), .Z(n4482) );
  NAND U6020 ( .A(n4484), .B(n4485), .Z(x[4]) );
  NAND U6021 ( .A(creg[4]), .B(init), .Z(n4484) );
  NAND U6022 ( .A(n4486), .B(n4487), .Z(x[49]) );
  NAND U6023 ( .A(creg[49]), .B(init), .Z(n4486) );
  NAND U6024 ( .A(n4488), .B(n4489), .Z(x[48]) );
  NAND U6025 ( .A(creg[48]), .B(init), .Z(n4488) );
  NAND U6026 ( .A(n4490), .B(n4491), .Z(x[47]) );
  NAND U6027 ( .A(creg[47]), .B(init), .Z(n4490) );
  NAND U6028 ( .A(n4492), .B(n4493), .Z(x[46]) );
  NAND U6029 ( .A(creg[46]), .B(init), .Z(n4492) );
  NAND U6030 ( .A(n4494), .B(n4495), .Z(x[45]) );
  NAND U6031 ( .A(creg[45]), .B(init), .Z(n4494) );
  NAND U6032 ( .A(n4496), .B(n4497), .Z(x[44]) );
  NAND U6033 ( .A(creg[44]), .B(init), .Z(n4496) );
  NAND U6034 ( .A(n4498), .B(n4499), .Z(x[43]) );
  NAND U6035 ( .A(creg[43]), .B(init), .Z(n4498) );
  NAND U6036 ( .A(n4500), .B(n4501), .Z(x[42]) );
  NAND U6037 ( .A(creg[42]), .B(init), .Z(n4500) );
  NAND U6038 ( .A(n4502), .B(n4503), .Z(x[41]) );
  NAND U6039 ( .A(creg[41]), .B(init), .Z(n4502) );
  NAND U6040 ( .A(n4504), .B(n4505), .Z(x[40]) );
  NAND U6041 ( .A(creg[40]), .B(init), .Z(n4504) );
  NAND U6042 ( .A(n4506), .B(n4507), .Z(x[3]) );
  NAND U6043 ( .A(creg[3]), .B(init), .Z(n4506) );
  NAND U6044 ( .A(n4508), .B(n4509), .Z(x[39]) );
  NAND U6045 ( .A(creg[39]), .B(init), .Z(n4508) );
  NAND U6046 ( .A(n4510), .B(n4511), .Z(x[38]) );
  NAND U6047 ( .A(creg[38]), .B(init), .Z(n4510) );
  NAND U6048 ( .A(n4512), .B(n4513), .Z(x[37]) );
  NAND U6049 ( .A(creg[37]), .B(init), .Z(n4512) );
  NAND U6050 ( .A(n4514), .B(n4515), .Z(x[36]) );
  NAND U6051 ( .A(creg[36]), .B(init), .Z(n4514) );
  NAND U6052 ( .A(n4516), .B(n4517), .Z(x[35]) );
  NAND U6053 ( .A(creg[35]), .B(init), .Z(n4516) );
  NAND U6054 ( .A(n4518), .B(n4519), .Z(x[34]) );
  NAND U6055 ( .A(creg[34]), .B(init), .Z(n4518) );
  NAND U6056 ( .A(n4520), .B(n4521), .Z(x[33]) );
  NAND U6057 ( .A(creg[33]), .B(init), .Z(n4520) );
  NAND U6058 ( .A(n4522), .B(n4523), .Z(x[32]) );
  NAND U6059 ( .A(creg[32]), .B(init), .Z(n4522) );
  NAND U6060 ( .A(n4524), .B(n4525), .Z(x[31]) );
  NAND U6061 ( .A(creg[31]), .B(init), .Z(n4524) );
  NAND U6062 ( .A(n4526), .B(n4527), .Z(x[30]) );
  NAND U6063 ( .A(creg[30]), .B(init), .Z(n4526) );
  NAND U6064 ( .A(n4528), .B(n4529), .Z(x[2]) );
  NAND U6065 ( .A(creg[2]), .B(init), .Z(n4528) );
  NAND U6066 ( .A(n4530), .B(n4531), .Z(x[29]) );
  NAND U6067 ( .A(creg[29]), .B(init), .Z(n4530) );
  NAND U6068 ( .A(n4532), .B(n4533), .Z(x[28]) );
  NAND U6069 ( .A(creg[28]), .B(init), .Z(n4532) );
  NAND U6070 ( .A(n4534), .B(n4535), .Z(x[27]) );
  NAND U6071 ( .A(creg[27]), .B(init), .Z(n4534) );
  NAND U6072 ( .A(n4536), .B(n4537), .Z(x[26]) );
  NAND U6073 ( .A(creg[26]), .B(init), .Z(n4536) );
  NAND U6074 ( .A(n4538), .B(n4539), .Z(x[25]) );
  NAND U6075 ( .A(creg[25]), .B(init), .Z(n4538) );
  NAND U6076 ( .A(n4540), .B(n4541), .Z(x[255]) );
  NAND U6077 ( .A(creg[255]), .B(init), .Z(n4540) );
  NAND U6078 ( .A(n4542), .B(n4543), .Z(x[254]) );
  NAND U6079 ( .A(creg[254]), .B(init), .Z(n4542) );
  NAND U6080 ( .A(n4544), .B(n4545), .Z(x[253]) );
  NAND U6081 ( .A(creg[253]), .B(init), .Z(n4544) );
  NAND U6082 ( .A(n4546), .B(n4547), .Z(x[252]) );
  NAND U6083 ( .A(creg[252]), .B(init), .Z(n4546) );
  NAND U6084 ( .A(n4548), .B(n4549), .Z(x[251]) );
  NAND U6085 ( .A(creg[251]), .B(init), .Z(n4548) );
  NAND U6086 ( .A(n4550), .B(n4551), .Z(x[250]) );
  NAND U6087 ( .A(creg[250]), .B(init), .Z(n4550) );
  NAND U6088 ( .A(n4552), .B(n4553), .Z(x[24]) );
  NAND U6089 ( .A(creg[24]), .B(init), .Z(n4552) );
  NAND U6090 ( .A(n4554), .B(n4555), .Z(x[249]) );
  NAND U6091 ( .A(creg[249]), .B(init), .Z(n4554) );
  NAND U6092 ( .A(n4556), .B(n4557), .Z(x[248]) );
  NAND U6093 ( .A(creg[248]), .B(init), .Z(n4556) );
  NAND U6094 ( .A(n4558), .B(n4559), .Z(x[247]) );
  NAND U6095 ( .A(creg[247]), .B(init), .Z(n4558) );
  NAND U6096 ( .A(n4560), .B(n4561), .Z(x[246]) );
  NAND U6097 ( .A(creg[246]), .B(init), .Z(n4560) );
  NAND U6098 ( .A(n4562), .B(n4563), .Z(x[245]) );
  NAND U6099 ( .A(creg[245]), .B(init), .Z(n4562) );
  NAND U6100 ( .A(n4564), .B(n4565), .Z(x[244]) );
  NAND U6101 ( .A(creg[244]), .B(init), .Z(n4564) );
  NAND U6102 ( .A(n4566), .B(n4567), .Z(x[243]) );
  NAND U6103 ( .A(creg[243]), .B(init), .Z(n4566) );
  NAND U6104 ( .A(n4568), .B(n4569), .Z(x[242]) );
  NAND U6105 ( .A(creg[242]), .B(init), .Z(n4568) );
  NAND U6106 ( .A(n4570), .B(n4571), .Z(x[241]) );
  NAND U6107 ( .A(creg[241]), .B(init), .Z(n4570) );
  NAND U6108 ( .A(n4572), .B(n4573), .Z(x[240]) );
  NAND U6109 ( .A(creg[240]), .B(init), .Z(n4572) );
  NAND U6110 ( .A(n4574), .B(n4575), .Z(x[23]) );
  NAND U6111 ( .A(creg[23]), .B(init), .Z(n4574) );
  NAND U6112 ( .A(n4576), .B(n4577), .Z(x[239]) );
  NAND U6113 ( .A(creg[239]), .B(init), .Z(n4576) );
  NAND U6114 ( .A(n4578), .B(n4579), .Z(x[238]) );
  NAND U6115 ( .A(creg[238]), .B(init), .Z(n4578) );
  NAND U6116 ( .A(n4580), .B(n4581), .Z(x[237]) );
  NAND U6117 ( .A(creg[237]), .B(init), .Z(n4580) );
  NAND U6118 ( .A(n4582), .B(n4583), .Z(x[236]) );
  NAND U6119 ( .A(creg[236]), .B(init), .Z(n4582) );
  NAND U6120 ( .A(n4584), .B(n4585), .Z(x[235]) );
  NAND U6121 ( .A(creg[235]), .B(init), .Z(n4584) );
  NAND U6122 ( .A(n4586), .B(n4587), .Z(x[234]) );
  NAND U6123 ( .A(creg[234]), .B(init), .Z(n4586) );
  NAND U6124 ( .A(n4588), .B(n4589), .Z(x[233]) );
  NAND U6125 ( .A(creg[233]), .B(init), .Z(n4588) );
  NAND U6126 ( .A(n4590), .B(n4591), .Z(x[232]) );
  NAND U6127 ( .A(creg[232]), .B(init), .Z(n4590) );
  NAND U6128 ( .A(n4592), .B(n4593), .Z(x[231]) );
  NAND U6129 ( .A(creg[231]), .B(init), .Z(n4592) );
  NAND U6130 ( .A(n4594), .B(n4595), .Z(x[230]) );
  NAND U6131 ( .A(creg[230]), .B(init), .Z(n4594) );
  NAND U6132 ( .A(n4596), .B(n4597), .Z(x[22]) );
  NAND U6133 ( .A(creg[22]), .B(init), .Z(n4596) );
  NAND U6134 ( .A(n4598), .B(n4599), .Z(x[229]) );
  NAND U6135 ( .A(creg[229]), .B(init), .Z(n4598) );
  NAND U6136 ( .A(n4600), .B(n4601), .Z(x[228]) );
  NAND U6137 ( .A(creg[228]), .B(init), .Z(n4600) );
  NAND U6138 ( .A(n4602), .B(n4603), .Z(x[227]) );
  NAND U6139 ( .A(creg[227]), .B(init), .Z(n4602) );
  NAND U6140 ( .A(n4604), .B(n4605), .Z(x[226]) );
  NAND U6141 ( .A(creg[226]), .B(init), .Z(n4604) );
  NAND U6142 ( .A(n4606), .B(n4607), .Z(x[225]) );
  NAND U6143 ( .A(creg[225]), .B(init), .Z(n4606) );
  NAND U6144 ( .A(n4608), .B(n4609), .Z(x[224]) );
  NAND U6145 ( .A(creg[224]), .B(init), .Z(n4608) );
  NAND U6146 ( .A(n4610), .B(n4611), .Z(x[223]) );
  NAND U6147 ( .A(creg[223]), .B(init), .Z(n4610) );
  NAND U6148 ( .A(n4612), .B(n4613), .Z(x[222]) );
  NAND U6149 ( .A(creg[222]), .B(init), .Z(n4612) );
  NAND U6150 ( .A(n4614), .B(n4615), .Z(x[221]) );
  NAND U6151 ( .A(creg[221]), .B(init), .Z(n4614) );
  NAND U6152 ( .A(n4616), .B(n4617), .Z(x[220]) );
  NAND U6153 ( .A(creg[220]), .B(init), .Z(n4616) );
  NAND U6154 ( .A(n4618), .B(n4619), .Z(x[21]) );
  NAND U6155 ( .A(creg[21]), .B(init), .Z(n4618) );
  NAND U6156 ( .A(n4620), .B(n4621), .Z(x[219]) );
  NAND U6157 ( .A(creg[219]), .B(init), .Z(n4620) );
  NAND U6158 ( .A(n4622), .B(n4623), .Z(x[218]) );
  NAND U6159 ( .A(creg[218]), .B(init), .Z(n4622) );
  NAND U6160 ( .A(n4624), .B(n4625), .Z(x[217]) );
  NAND U6161 ( .A(creg[217]), .B(init), .Z(n4624) );
  NAND U6162 ( .A(n4626), .B(n4627), .Z(x[216]) );
  NAND U6163 ( .A(creg[216]), .B(init), .Z(n4626) );
  NAND U6164 ( .A(n4628), .B(n4629), .Z(x[215]) );
  NAND U6165 ( .A(creg[215]), .B(init), .Z(n4628) );
  NAND U6166 ( .A(n4630), .B(n4631), .Z(x[214]) );
  NAND U6167 ( .A(creg[214]), .B(init), .Z(n4630) );
  NAND U6168 ( .A(n4632), .B(n4633), .Z(x[213]) );
  NAND U6169 ( .A(creg[213]), .B(init), .Z(n4632) );
  NAND U6170 ( .A(n4634), .B(n4635), .Z(x[212]) );
  NAND U6171 ( .A(creg[212]), .B(init), .Z(n4634) );
  NAND U6172 ( .A(n4636), .B(n4637), .Z(x[211]) );
  NAND U6173 ( .A(creg[211]), .B(init), .Z(n4636) );
  NAND U6174 ( .A(n4638), .B(n4639), .Z(x[210]) );
  NAND U6175 ( .A(creg[210]), .B(init), .Z(n4638) );
  NAND U6176 ( .A(n4640), .B(n4641), .Z(x[20]) );
  NAND U6177 ( .A(creg[20]), .B(init), .Z(n4640) );
  NAND U6178 ( .A(n4642), .B(n4643), .Z(x[209]) );
  NAND U6179 ( .A(creg[209]), .B(init), .Z(n4642) );
  NAND U6180 ( .A(n4644), .B(n4645), .Z(x[208]) );
  NAND U6181 ( .A(creg[208]), .B(init), .Z(n4644) );
  NAND U6182 ( .A(n4646), .B(n4647), .Z(x[207]) );
  NAND U6183 ( .A(creg[207]), .B(init), .Z(n4646) );
  NAND U6184 ( .A(n4648), .B(n4649), .Z(x[206]) );
  NAND U6185 ( .A(creg[206]), .B(init), .Z(n4648) );
  NAND U6186 ( .A(n4650), .B(n4651), .Z(x[205]) );
  NAND U6187 ( .A(creg[205]), .B(init), .Z(n4650) );
  NAND U6188 ( .A(n4652), .B(n4653), .Z(x[204]) );
  NAND U6189 ( .A(creg[204]), .B(init), .Z(n4652) );
  NAND U6190 ( .A(n4654), .B(n4655), .Z(x[203]) );
  NAND U6191 ( .A(creg[203]), .B(init), .Z(n4654) );
  NAND U6192 ( .A(n4656), .B(n4657), .Z(x[202]) );
  NAND U6193 ( .A(creg[202]), .B(init), .Z(n4656) );
  NAND U6194 ( .A(n4658), .B(n4659), .Z(x[201]) );
  NAND U6195 ( .A(creg[201]), .B(init), .Z(n4658) );
  NAND U6196 ( .A(n4660), .B(n4661), .Z(x[200]) );
  NAND U6197 ( .A(creg[200]), .B(init), .Z(n4660) );
  NAND U6198 ( .A(n4662), .B(n4663), .Z(x[1]) );
  NAND U6199 ( .A(creg[1]), .B(init), .Z(n4662) );
  NAND U6200 ( .A(n4664), .B(n4665), .Z(x[19]) );
  NAND U6201 ( .A(creg[19]), .B(init), .Z(n4664) );
  NAND U6202 ( .A(n4666), .B(n4667), .Z(x[199]) );
  NAND U6203 ( .A(creg[199]), .B(init), .Z(n4666) );
  NAND U6204 ( .A(n4668), .B(n4669), .Z(x[198]) );
  NAND U6205 ( .A(creg[198]), .B(init), .Z(n4668) );
  NAND U6206 ( .A(n4670), .B(n4671), .Z(x[197]) );
  NAND U6207 ( .A(creg[197]), .B(init), .Z(n4670) );
  NAND U6208 ( .A(n4672), .B(n4673), .Z(x[196]) );
  NAND U6209 ( .A(creg[196]), .B(init), .Z(n4672) );
  NAND U6210 ( .A(n4674), .B(n4675), .Z(x[195]) );
  NAND U6211 ( .A(creg[195]), .B(init), .Z(n4674) );
  NAND U6212 ( .A(n4676), .B(n4677), .Z(x[194]) );
  NAND U6213 ( .A(creg[194]), .B(init), .Z(n4676) );
  NAND U6214 ( .A(n4678), .B(n4679), .Z(x[193]) );
  NAND U6215 ( .A(creg[193]), .B(init), .Z(n4678) );
  NAND U6216 ( .A(n4680), .B(n4681), .Z(x[192]) );
  NAND U6217 ( .A(creg[192]), .B(init), .Z(n4680) );
  NAND U6218 ( .A(n4682), .B(n4683), .Z(x[191]) );
  NAND U6219 ( .A(creg[191]), .B(init), .Z(n4682) );
  NAND U6220 ( .A(n4684), .B(n4685), .Z(x[190]) );
  NAND U6221 ( .A(creg[190]), .B(init), .Z(n4684) );
  NAND U6222 ( .A(n4686), .B(n4687), .Z(x[18]) );
  NAND U6223 ( .A(creg[18]), .B(init), .Z(n4686) );
  NAND U6224 ( .A(n4688), .B(n4689), .Z(x[189]) );
  NAND U6225 ( .A(creg[189]), .B(init), .Z(n4688) );
  NAND U6226 ( .A(n4690), .B(n4691), .Z(x[188]) );
  NAND U6227 ( .A(creg[188]), .B(init), .Z(n4690) );
  NAND U6228 ( .A(n4692), .B(n4693), .Z(x[187]) );
  NAND U6229 ( .A(creg[187]), .B(init), .Z(n4692) );
  NAND U6230 ( .A(n4694), .B(n4695), .Z(x[186]) );
  NAND U6231 ( .A(creg[186]), .B(init), .Z(n4694) );
  NAND U6232 ( .A(n4696), .B(n4697), .Z(x[185]) );
  NAND U6233 ( .A(creg[185]), .B(init), .Z(n4696) );
  NAND U6234 ( .A(n4698), .B(n4699), .Z(x[184]) );
  NAND U6235 ( .A(creg[184]), .B(init), .Z(n4698) );
  NAND U6236 ( .A(n4700), .B(n4701), .Z(x[183]) );
  NAND U6237 ( .A(creg[183]), .B(init), .Z(n4700) );
  NAND U6238 ( .A(n4702), .B(n4703), .Z(x[182]) );
  NAND U6239 ( .A(creg[182]), .B(init), .Z(n4702) );
  NAND U6240 ( .A(n4704), .B(n4705), .Z(x[181]) );
  NAND U6241 ( .A(creg[181]), .B(init), .Z(n4704) );
  NAND U6242 ( .A(n4706), .B(n4707), .Z(x[180]) );
  NAND U6243 ( .A(creg[180]), .B(init), .Z(n4706) );
  NAND U6244 ( .A(n4708), .B(n4709), .Z(x[17]) );
  NAND U6245 ( .A(creg[17]), .B(init), .Z(n4708) );
  NAND U6246 ( .A(n4710), .B(n4711), .Z(x[179]) );
  NAND U6247 ( .A(creg[179]), .B(init), .Z(n4710) );
  NAND U6248 ( .A(n4712), .B(n4713), .Z(x[178]) );
  NAND U6249 ( .A(creg[178]), .B(init), .Z(n4712) );
  NAND U6250 ( .A(n4714), .B(n4715), .Z(x[177]) );
  NAND U6251 ( .A(creg[177]), .B(init), .Z(n4714) );
  NAND U6252 ( .A(n4716), .B(n4717), .Z(x[176]) );
  NAND U6253 ( .A(creg[176]), .B(init), .Z(n4716) );
  NAND U6254 ( .A(n4718), .B(n4719), .Z(x[175]) );
  NAND U6255 ( .A(creg[175]), .B(init), .Z(n4718) );
  NAND U6256 ( .A(n4720), .B(n4721), .Z(x[174]) );
  NAND U6257 ( .A(creg[174]), .B(init), .Z(n4720) );
  NAND U6258 ( .A(n4722), .B(n4723), .Z(x[173]) );
  NAND U6259 ( .A(creg[173]), .B(init), .Z(n4722) );
  NAND U6260 ( .A(n4724), .B(n4725), .Z(x[172]) );
  NAND U6261 ( .A(creg[172]), .B(init), .Z(n4724) );
  NAND U6262 ( .A(n4726), .B(n4727), .Z(x[171]) );
  NAND U6263 ( .A(creg[171]), .B(init), .Z(n4726) );
  NAND U6264 ( .A(n4728), .B(n4729), .Z(x[170]) );
  NAND U6265 ( .A(creg[170]), .B(init), .Z(n4728) );
  NAND U6266 ( .A(n4730), .B(n4731), .Z(x[16]) );
  NAND U6267 ( .A(creg[16]), .B(init), .Z(n4730) );
  NAND U6268 ( .A(n4732), .B(n4733), .Z(x[169]) );
  NAND U6269 ( .A(creg[169]), .B(init), .Z(n4732) );
  NAND U6270 ( .A(n4734), .B(n4735), .Z(x[168]) );
  NAND U6271 ( .A(creg[168]), .B(init), .Z(n4734) );
  NAND U6272 ( .A(n4736), .B(n4737), .Z(x[167]) );
  NAND U6273 ( .A(creg[167]), .B(init), .Z(n4736) );
  NAND U6274 ( .A(n4738), .B(n4739), .Z(x[166]) );
  NAND U6275 ( .A(creg[166]), .B(init), .Z(n4738) );
  NAND U6276 ( .A(n4740), .B(n4741), .Z(x[165]) );
  NAND U6277 ( .A(creg[165]), .B(init), .Z(n4740) );
  NAND U6278 ( .A(n4742), .B(n4743), .Z(x[164]) );
  NAND U6279 ( .A(creg[164]), .B(init), .Z(n4742) );
  NAND U6280 ( .A(n4744), .B(n4745), .Z(x[163]) );
  NAND U6281 ( .A(creg[163]), .B(init), .Z(n4744) );
  NAND U6282 ( .A(n4746), .B(n4747), .Z(x[162]) );
  NAND U6283 ( .A(creg[162]), .B(init), .Z(n4746) );
  NAND U6284 ( .A(n4748), .B(n4749), .Z(x[161]) );
  NAND U6285 ( .A(creg[161]), .B(init), .Z(n4748) );
  NAND U6286 ( .A(n4750), .B(n4751), .Z(x[160]) );
  NAND U6287 ( .A(creg[160]), .B(init), .Z(n4750) );
  NAND U6288 ( .A(n4752), .B(n4753), .Z(x[15]) );
  NAND U6289 ( .A(creg[15]), .B(init), .Z(n4752) );
  NAND U6290 ( .A(n4754), .B(n4755), .Z(x[159]) );
  NAND U6291 ( .A(creg[159]), .B(init), .Z(n4754) );
  NAND U6292 ( .A(n4756), .B(n4757), .Z(x[158]) );
  NAND U6293 ( .A(creg[158]), .B(init), .Z(n4756) );
  NAND U6294 ( .A(n4758), .B(n4759), .Z(x[157]) );
  NAND U6295 ( .A(creg[157]), .B(init), .Z(n4758) );
  NAND U6296 ( .A(n4760), .B(n4761), .Z(x[156]) );
  NAND U6297 ( .A(creg[156]), .B(init), .Z(n4760) );
  NAND U6298 ( .A(n4762), .B(n4763), .Z(x[155]) );
  NAND U6299 ( .A(creg[155]), .B(init), .Z(n4762) );
  NAND U6300 ( .A(n4764), .B(n4765), .Z(x[154]) );
  NAND U6301 ( .A(creg[154]), .B(init), .Z(n4764) );
  NAND U6302 ( .A(n4766), .B(n4767), .Z(x[153]) );
  NAND U6303 ( .A(creg[153]), .B(init), .Z(n4766) );
  NAND U6304 ( .A(n4768), .B(n4769), .Z(x[152]) );
  NAND U6305 ( .A(creg[152]), .B(init), .Z(n4768) );
  NAND U6306 ( .A(n4770), .B(n4771), .Z(x[151]) );
  NAND U6307 ( .A(creg[151]), .B(init), .Z(n4770) );
  NAND U6308 ( .A(n4772), .B(n4773), .Z(x[150]) );
  NAND U6309 ( .A(creg[150]), .B(init), .Z(n4772) );
  NAND U6310 ( .A(n4774), .B(n4775), .Z(x[14]) );
  NAND U6311 ( .A(creg[14]), .B(init), .Z(n4774) );
  NAND U6312 ( .A(n4776), .B(n4777), .Z(x[149]) );
  NAND U6313 ( .A(creg[149]), .B(init), .Z(n4776) );
  NAND U6314 ( .A(n4778), .B(n4779), .Z(x[148]) );
  NAND U6315 ( .A(creg[148]), .B(init), .Z(n4778) );
  NAND U6316 ( .A(n4780), .B(n4781), .Z(x[147]) );
  NAND U6317 ( .A(creg[147]), .B(init), .Z(n4780) );
  NAND U6318 ( .A(n4782), .B(n4783), .Z(x[146]) );
  NAND U6319 ( .A(creg[146]), .B(init), .Z(n4782) );
  NAND U6320 ( .A(n4784), .B(n4785), .Z(x[145]) );
  NAND U6321 ( .A(creg[145]), .B(init), .Z(n4784) );
  NAND U6322 ( .A(n4786), .B(n4787), .Z(x[144]) );
  NAND U6323 ( .A(creg[144]), .B(init), .Z(n4786) );
  NAND U6324 ( .A(n4788), .B(n4789), .Z(x[143]) );
  NAND U6325 ( .A(creg[143]), .B(init), .Z(n4788) );
  NAND U6326 ( .A(n4790), .B(n4791), .Z(x[142]) );
  NAND U6327 ( .A(creg[142]), .B(init), .Z(n4790) );
  NAND U6328 ( .A(n4792), .B(n4793), .Z(x[141]) );
  NAND U6329 ( .A(creg[141]), .B(init), .Z(n4792) );
  NAND U6330 ( .A(n4794), .B(n4795), .Z(x[140]) );
  NAND U6331 ( .A(creg[140]), .B(init), .Z(n4794) );
  NAND U6332 ( .A(n4796), .B(n4797), .Z(x[13]) );
  NAND U6333 ( .A(creg[13]), .B(init), .Z(n4796) );
  NAND U6334 ( .A(n4798), .B(n4799), .Z(x[139]) );
  NAND U6335 ( .A(creg[139]), .B(init), .Z(n4798) );
  NAND U6336 ( .A(n4800), .B(n4801), .Z(x[138]) );
  NAND U6337 ( .A(creg[138]), .B(init), .Z(n4800) );
  NAND U6338 ( .A(n4802), .B(n4803), .Z(x[137]) );
  NAND U6339 ( .A(creg[137]), .B(init), .Z(n4802) );
  NAND U6340 ( .A(n4804), .B(n4805), .Z(x[136]) );
  NAND U6341 ( .A(creg[136]), .B(init), .Z(n4804) );
  NAND U6342 ( .A(n4806), .B(n4807), .Z(x[135]) );
  NAND U6343 ( .A(creg[135]), .B(init), .Z(n4806) );
  NAND U6344 ( .A(n4808), .B(n4809), .Z(x[134]) );
  NAND U6345 ( .A(creg[134]), .B(init), .Z(n4808) );
  NAND U6346 ( .A(n4810), .B(n4811), .Z(x[133]) );
  NAND U6347 ( .A(creg[133]), .B(init), .Z(n4810) );
  NAND U6348 ( .A(n4812), .B(n4813), .Z(x[132]) );
  NAND U6349 ( .A(creg[132]), .B(init), .Z(n4812) );
  NAND U6350 ( .A(n4814), .B(n4815), .Z(x[131]) );
  NAND U6351 ( .A(creg[131]), .B(init), .Z(n4814) );
  NAND U6352 ( .A(n4816), .B(n4817), .Z(x[130]) );
  NAND U6353 ( .A(creg[130]), .B(init), .Z(n4816) );
  NAND U6354 ( .A(n4818), .B(n4819), .Z(x[12]) );
  NAND U6355 ( .A(creg[12]), .B(init), .Z(n4818) );
  NAND U6356 ( .A(n4820), .B(n4821), .Z(x[129]) );
  NAND U6357 ( .A(creg[129]), .B(init), .Z(n4820) );
  NAND U6358 ( .A(n4822), .B(n4823), .Z(x[128]) );
  NAND U6359 ( .A(creg[128]), .B(init), .Z(n4822) );
  NAND U6360 ( .A(n4824), .B(n4825), .Z(x[127]) );
  NAND U6361 ( .A(creg[127]), .B(init), .Z(n4824) );
  NAND U6362 ( .A(n4826), .B(n4827), .Z(x[126]) );
  NAND U6363 ( .A(creg[126]), .B(init), .Z(n4826) );
  NAND U6364 ( .A(n4828), .B(n4829), .Z(x[125]) );
  NAND U6365 ( .A(creg[125]), .B(init), .Z(n4828) );
  NAND U6366 ( .A(n4830), .B(n4831), .Z(x[124]) );
  NAND U6367 ( .A(creg[124]), .B(init), .Z(n4830) );
  NAND U6368 ( .A(n4832), .B(n4833), .Z(x[123]) );
  NAND U6369 ( .A(creg[123]), .B(init), .Z(n4832) );
  NAND U6370 ( .A(n4834), .B(n4835), .Z(x[122]) );
  NAND U6371 ( .A(creg[122]), .B(init), .Z(n4834) );
  NAND U6372 ( .A(n4836), .B(n4837), .Z(x[121]) );
  NAND U6373 ( .A(creg[121]), .B(init), .Z(n4836) );
  NAND U6374 ( .A(n4838), .B(n4839), .Z(x[120]) );
  NAND U6375 ( .A(creg[120]), .B(init), .Z(n4838) );
  NAND U6376 ( .A(n4840), .B(n4841), .Z(x[11]) );
  NAND U6377 ( .A(creg[11]), .B(init), .Z(n4840) );
  NAND U6378 ( .A(n4842), .B(n4843), .Z(x[119]) );
  NAND U6379 ( .A(creg[119]), .B(init), .Z(n4842) );
  NAND U6380 ( .A(n4844), .B(n4845), .Z(x[118]) );
  NAND U6381 ( .A(creg[118]), .B(init), .Z(n4844) );
  NAND U6382 ( .A(n4846), .B(n4847), .Z(x[117]) );
  NAND U6383 ( .A(creg[117]), .B(init), .Z(n4846) );
  NAND U6384 ( .A(n4848), .B(n4849), .Z(x[116]) );
  NAND U6385 ( .A(creg[116]), .B(init), .Z(n4848) );
  NAND U6386 ( .A(n4850), .B(n4851), .Z(x[115]) );
  NAND U6387 ( .A(creg[115]), .B(init), .Z(n4850) );
  NAND U6388 ( .A(n4852), .B(n4853), .Z(x[114]) );
  NAND U6389 ( .A(creg[114]), .B(init), .Z(n4852) );
  NAND U6390 ( .A(n4854), .B(n4855), .Z(x[113]) );
  NAND U6391 ( .A(creg[113]), .B(init), .Z(n4854) );
  NAND U6392 ( .A(n4856), .B(n4857), .Z(x[112]) );
  NAND U6393 ( .A(creg[112]), .B(init), .Z(n4856) );
  NAND U6394 ( .A(n4858), .B(n4859), .Z(x[111]) );
  NAND U6395 ( .A(creg[111]), .B(init), .Z(n4858) );
  NAND U6396 ( .A(n4860), .B(n4861), .Z(x[110]) );
  NAND U6397 ( .A(creg[110]), .B(init), .Z(n4860) );
  NAND U6398 ( .A(n4862), .B(n4863), .Z(x[10]) );
  NAND U6399 ( .A(creg[10]), .B(init), .Z(n4862) );
  NAND U6400 ( .A(n4864), .B(n4865), .Z(x[109]) );
  NAND U6401 ( .A(creg[109]), .B(init), .Z(n4864) );
  NAND U6402 ( .A(n4866), .B(n4867), .Z(x[108]) );
  NAND U6403 ( .A(creg[108]), .B(init), .Z(n4866) );
  NAND U6404 ( .A(n4868), .B(n4869), .Z(x[107]) );
  NAND U6405 ( .A(creg[107]), .B(init), .Z(n4868) );
  NAND U6406 ( .A(n4870), .B(n4871), .Z(x[106]) );
  NAND U6407 ( .A(creg[106]), .B(init), .Z(n4870) );
  NAND U6408 ( .A(n4872), .B(n4873), .Z(x[105]) );
  NAND U6409 ( .A(creg[105]), .B(init), .Z(n4872) );
  NAND U6410 ( .A(n4874), .B(n4875), .Z(x[104]) );
  NAND U6411 ( .A(creg[104]), .B(init), .Z(n4874) );
  NAND U6412 ( .A(n4876), .B(n4877), .Z(x[103]) );
  NAND U6413 ( .A(creg[103]), .B(init), .Z(n4876) );
  NAND U6414 ( .A(n4878), .B(n4879), .Z(x[102]) );
  NAND U6415 ( .A(creg[102]), .B(init), .Z(n4878) );
  NAND U6416 ( .A(n4880), .B(n4881), .Z(x[101]) );
  NAND U6417 ( .A(creg[101]), .B(init), .Z(n4880) );
  NAND U6418 ( .A(n4882), .B(n4883), .Z(x[100]) );
  NAND U6419 ( .A(creg[100]), .B(init), .Z(n4882) );
  NAND U6420 ( .A(n4884), .B(n4885), .Z(x[0]) );
  NAND U6421 ( .A(creg[0]), .B(init), .Z(n4884) );
  AND U6422 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  AND U6423 ( .A(start_reg[99]), .B(init), .Z(start_in[99]) );
  AND U6424 ( .A(start_reg[98]), .B(init), .Z(start_in[98]) );
  AND U6425 ( .A(start_reg[97]), .B(init), .Z(start_in[97]) );
  AND U6426 ( .A(start_reg[96]), .B(init), .Z(start_in[96]) );
  AND U6427 ( .A(start_reg[95]), .B(init), .Z(start_in[95]) );
  AND U6428 ( .A(start_reg[94]), .B(init), .Z(start_in[94]) );
  AND U6429 ( .A(start_reg[93]), .B(init), .Z(start_in[93]) );
  AND U6430 ( .A(start_reg[92]), .B(init), .Z(start_in[92]) );
  AND U6431 ( .A(start_reg[91]), .B(init), .Z(start_in[91]) );
  AND U6432 ( .A(start_reg[90]), .B(init), .Z(start_in[90]) );
  AND U6433 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U6434 ( .A(start_reg[89]), .B(init), .Z(start_in[89]) );
  AND U6435 ( .A(start_reg[88]), .B(init), .Z(start_in[88]) );
  AND U6436 ( .A(start_reg[87]), .B(init), .Z(start_in[87]) );
  AND U6437 ( .A(start_reg[86]), .B(init), .Z(start_in[86]) );
  AND U6438 ( .A(start_reg[85]), .B(init), .Z(start_in[85]) );
  AND U6439 ( .A(start_reg[84]), .B(init), .Z(start_in[84]) );
  AND U6440 ( .A(start_reg[83]), .B(init), .Z(start_in[83]) );
  AND U6441 ( .A(start_reg[82]), .B(init), .Z(start_in[82]) );
  AND U6442 ( .A(start_reg[81]), .B(init), .Z(start_in[81]) );
  AND U6443 ( .A(start_reg[80]), .B(init), .Z(start_in[80]) );
  AND U6444 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U6445 ( .A(start_reg[79]), .B(init), .Z(start_in[79]) );
  AND U6446 ( .A(start_reg[78]), .B(init), .Z(start_in[78]) );
  AND U6447 ( .A(start_reg[77]), .B(init), .Z(start_in[77]) );
  AND U6448 ( .A(start_reg[76]), .B(init), .Z(start_in[76]) );
  AND U6449 ( .A(start_reg[75]), .B(init), .Z(start_in[75]) );
  AND U6450 ( .A(start_reg[74]), .B(init), .Z(start_in[74]) );
  AND U6451 ( .A(start_reg[73]), .B(init), .Z(start_in[73]) );
  AND U6452 ( .A(start_reg[72]), .B(init), .Z(start_in[72]) );
  AND U6453 ( .A(start_reg[71]), .B(init), .Z(start_in[71]) );
  AND U6454 ( .A(start_reg[70]), .B(init), .Z(start_in[70]) );
  AND U6455 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U6456 ( .A(start_reg[69]), .B(init), .Z(start_in[69]) );
  AND U6457 ( .A(start_reg[68]), .B(init), .Z(start_in[68]) );
  AND U6458 ( .A(start_reg[67]), .B(init), .Z(start_in[67]) );
  AND U6459 ( .A(start_reg[66]), .B(init), .Z(start_in[66]) );
  AND U6460 ( .A(start_reg[65]), .B(init), .Z(start_in[65]) );
  AND U6461 ( .A(start_reg[64]), .B(init), .Z(start_in[64]) );
  AND U6462 ( .A(start_reg[63]), .B(init), .Z(start_in[63]) );
  AND U6463 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U6464 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U6465 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U6466 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U6467 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U6468 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U6469 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U6470 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U6471 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U6472 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U6473 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U6474 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U6475 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U6476 ( .A(start_reg[510]), .B(init), .Z(start_in[510]) );
  AND U6477 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U6478 ( .A(start_reg[509]), .B(init), .Z(start_in[509]) );
  AND U6479 ( .A(start_reg[508]), .B(init), .Z(start_in[508]) );
  AND U6480 ( .A(start_reg[507]), .B(init), .Z(start_in[507]) );
  AND U6481 ( .A(start_reg[506]), .B(init), .Z(start_in[506]) );
  AND U6482 ( .A(start_reg[505]), .B(init), .Z(start_in[505]) );
  AND U6483 ( .A(start_reg[504]), .B(init), .Z(start_in[504]) );
  AND U6484 ( .A(start_reg[503]), .B(init), .Z(start_in[503]) );
  AND U6485 ( .A(start_reg[502]), .B(init), .Z(start_in[502]) );
  AND U6486 ( .A(start_reg[501]), .B(init), .Z(start_in[501]) );
  AND U6487 ( .A(start_reg[500]), .B(init), .Z(start_in[500]) );
  AND U6488 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U6489 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U6490 ( .A(start_reg[499]), .B(init), .Z(start_in[499]) );
  AND U6491 ( .A(start_reg[498]), .B(init), .Z(start_in[498]) );
  AND U6492 ( .A(start_reg[497]), .B(init), .Z(start_in[497]) );
  AND U6493 ( .A(start_reg[496]), .B(init), .Z(start_in[496]) );
  AND U6494 ( .A(start_reg[495]), .B(init), .Z(start_in[495]) );
  AND U6495 ( .A(start_reg[494]), .B(init), .Z(start_in[494]) );
  AND U6496 ( .A(start_reg[493]), .B(init), .Z(start_in[493]) );
  AND U6497 ( .A(start_reg[492]), .B(init), .Z(start_in[492]) );
  AND U6498 ( .A(start_reg[491]), .B(init), .Z(start_in[491]) );
  AND U6499 ( .A(start_reg[490]), .B(init), .Z(start_in[490]) );
  AND U6500 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U6501 ( .A(start_reg[489]), .B(init), .Z(start_in[489]) );
  AND U6502 ( .A(start_reg[488]), .B(init), .Z(start_in[488]) );
  AND U6503 ( .A(start_reg[487]), .B(init), .Z(start_in[487]) );
  AND U6504 ( .A(start_reg[486]), .B(init), .Z(start_in[486]) );
  AND U6505 ( .A(start_reg[485]), .B(init), .Z(start_in[485]) );
  AND U6506 ( .A(start_reg[484]), .B(init), .Z(start_in[484]) );
  AND U6507 ( .A(start_reg[483]), .B(init), .Z(start_in[483]) );
  AND U6508 ( .A(start_reg[482]), .B(init), .Z(start_in[482]) );
  AND U6509 ( .A(start_reg[481]), .B(init), .Z(start_in[481]) );
  AND U6510 ( .A(start_reg[480]), .B(init), .Z(start_in[480]) );
  AND U6511 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U6512 ( .A(start_reg[479]), .B(init), .Z(start_in[479]) );
  AND U6513 ( .A(start_reg[478]), .B(init), .Z(start_in[478]) );
  AND U6514 ( .A(start_reg[477]), .B(init), .Z(start_in[477]) );
  AND U6515 ( .A(start_reg[476]), .B(init), .Z(start_in[476]) );
  AND U6516 ( .A(start_reg[475]), .B(init), .Z(start_in[475]) );
  AND U6517 ( .A(start_reg[474]), .B(init), .Z(start_in[474]) );
  AND U6518 ( .A(start_reg[473]), .B(init), .Z(start_in[473]) );
  AND U6519 ( .A(start_reg[472]), .B(init), .Z(start_in[472]) );
  AND U6520 ( .A(start_reg[471]), .B(init), .Z(start_in[471]) );
  AND U6521 ( .A(start_reg[470]), .B(init), .Z(start_in[470]) );
  AND U6522 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U6523 ( .A(start_reg[469]), .B(init), .Z(start_in[469]) );
  AND U6524 ( .A(start_reg[468]), .B(init), .Z(start_in[468]) );
  AND U6525 ( .A(start_reg[467]), .B(init), .Z(start_in[467]) );
  AND U6526 ( .A(start_reg[466]), .B(init), .Z(start_in[466]) );
  AND U6527 ( .A(start_reg[465]), .B(init), .Z(start_in[465]) );
  AND U6528 ( .A(start_reg[464]), .B(init), .Z(start_in[464]) );
  AND U6529 ( .A(start_reg[463]), .B(init), .Z(start_in[463]) );
  AND U6530 ( .A(start_reg[462]), .B(init), .Z(start_in[462]) );
  AND U6531 ( .A(start_reg[461]), .B(init), .Z(start_in[461]) );
  AND U6532 ( .A(start_reg[460]), .B(init), .Z(start_in[460]) );
  AND U6533 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U6534 ( .A(start_reg[459]), .B(init), .Z(start_in[459]) );
  AND U6535 ( .A(start_reg[458]), .B(init), .Z(start_in[458]) );
  AND U6536 ( .A(start_reg[457]), .B(init), .Z(start_in[457]) );
  AND U6537 ( .A(start_reg[456]), .B(init), .Z(start_in[456]) );
  AND U6538 ( .A(start_reg[455]), .B(init), .Z(start_in[455]) );
  AND U6539 ( .A(start_reg[454]), .B(init), .Z(start_in[454]) );
  AND U6540 ( .A(start_reg[453]), .B(init), .Z(start_in[453]) );
  AND U6541 ( .A(start_reg[452]), .B(init), .Z(start_in[452]) );
  AND U6542 ( .A(start_reg[451]), .B(init), .Z(start_in[451]) );
  AND U6543 ( .A(start_reg[450]), .B(init), .Z(start_in[450]) );
  AND U6544 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U6545 ( .A(start_reg[449]), .B(init), .Z(start_in[449]) );
  AND U6546 ( .A(start_reg[448]), .B(init), .Z(start_in[448]) );
  AND U6547 ( .A(start_reg[447]), .B(init), .Z(start_in[447]) );
  AND U6548 ( .A(start_reg[446]), .B(init), .Z(start_in[446]) );
  AND U6549 ( .A(start_reg[445]), .B(init), .Z(start_in[445]) );
  AND U6550 ( .A(start_reg[444]), .B(init), .Z(start_in[444]) );
  AND U6551 ( .A(start_reg[443]), .B(init), .Z(start_in[443]) );
  AND U6552 ( .A(start_reg[442]), .B(init), .Z(start_in[442]) );
  AND U6553 ( .A(start_reg[441]), .B(init), .Z(start_in[441]) );
  AND U6554 ( .A(start_reg[440]), .B(init), .Z(start_in[440]) );
  AND U6555 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U6556 ( .A(start_reg[439]), .B(init), .Z(start_in[439]) );
  AND U6557 ( .A(start_reg[438]), .B(init), .Z(start_in[438]) );
  AND U6558 ( .A(start_reg[437]), .B(init), .Z(start_in[437]) );
  AND U6559 ( .A(start_reg[436]), .B(init), .Z(start_in[436]) );
  AND U6560 ( .A(start_reg[435]), .B(init), .Z(start_in[435]) );
  AND U6561 ( .A(start_reg[434]), .B(init), .Z(start_in[434]) );
  AND U6562 ( .A(start_reg[433]), .B(init), .Z(start_in[433]) );
  AND U6563 ( .A(start_reg[432]), .B(init), .Z(start_in[432]) );
  AND U6564 ( .A(start_reg[431]), .B(init), .Z(start_in[431]) );
  AND U6565 ( .A(start_reg[430]), .B(init), .Z(start_in[430]) );
  AND U6566 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U6567 ( .A(start_reg[429]), .B(init), .Z(start_in[429]) );
  AND U6568 ( .A(start_reg[428]), .B(init), .Z(start_in[428]) );
  AND U6569 ( .A(start_reg[427]), .B(init), .Z(start_in[427]) );
  AND U6570 ( .A(start_reg[426]), .B(init), .Z(start_in[426]) );
  AND U6571 ( .A(start_reg[425]), .B(init), .Z(start_in[425]) );
  AND U6572 ( .A(start_reg[424]), .B(init), .Z(start_in[424]) );
  AND U6573 ( .A(start_reg[423]), .B(init), .Z(start_in[423]) );
  AND U6574 ( .A(start_reg[422]), .B(init), .Z(start_in[422]) );
  AND U6575 ( .A(start_reg[421]), .B(init), .Z(start_in[421]) );
  AND U6576 ( .A(start_reg[420]), .B(init), .Z(start_in[420]) );
  AND U6577 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U6578 ( .A(start_reg[419]), .B(init), .Z(start_in[419]) );
  AND U6579 ( .A(start_reg[418]), .B(init), .Z(start_in[418]) );
  AND U6580 ( .A(start_reg[417]), .B(init), .Z(start_in[417]) );
  AND U6581 ( .A(start_reg[416]), .B(init), .Z(start_in[416]) );
  AND U6582 ( .A(start_reg[415]), .B(init), .Z(start_in[415]) );
  AND U6583 ( .A(start_reg[414]), .B(init), .Z(start_in[414]) );
  AND U6584 ( .A(start_reg[413]), .B(init), .Z(start_in[413]) );
  AND U6585 ( .A(start_reg[412]), .B(init), .Z(start_in[412]) );
  AND U6586 ( .A(start_reg[411]), .B(init), .Z(start_in[411]) );
  AND U6587 ( .A(start_reg[410]), .B(init), .Z(start_in[410]) );
  AND U6588 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U6589 ( .A(start_reg[409]), .B(init), .Z(start_in[409]) );
  AND U6590 ( .A(start_reg[408]), .B(init), .Z(start_in[408]) );
  AND U6591 ( .A(start_reg[407]), .B(init), .Z(start_in[407]) );
  AND U6592 ( .A(start_reg[406]), .B(init), .Z(start_in[406]) );
  AND U6593 ( .A(start_reg[405]), .B(init), .Z(start_in[405]) );
  AND U6594 ( .A(start_reg[404]), .B(init), .Z(start_in[404]) );
  AND U6595 ( .A(start_reg[403]), .B(init), .Z(start_in[403]) );
  AND U6596 ( .A(start_reg[402]), .B(init), .Z(start_in[402]) );
  AND U6597 ( .A(start_reg[401]), .B(init), .Z(start_in[401]) );
  AND U6598 ( .A(start_reg[400]), .B(init), .Z(start_in[400]) );
  AND U6599 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U6600 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U6601 ( .A(start_reg[399]), .B(init), .Z(start_in[399]) );
  AND U6602 ( .A(start_reg[398]), .B(init), .Z(start_in[398]) );
  AND U6603 ( .A(start_reg[397]), .B(init), .Z(start_in[397]) );
  AND U6604 ( .A(start_reg[396]), .B(init), .Z(start_in[396]) );
  AND U6605 ( .A(start_reg[395]), .B(init), .Z(start_in[395]) );
  AND U6606 ( .A(start_reg[394]), .B(init), .Z(start_in[394]) );
  AND U6607 ( .A(start_reg[393]), .B(init), .Z(start_in[393]) );
  AND U6608 ( .A(start_reg[392]), .B(init), .Z(start_in[392]) );
  AND U6609 ( .A(start_reg[391]), .B(init), .Z(start_in[391]) );
  AND U6610 ( .A(start_reg[390]), .B(init), .Z(start_in[390]) );
  AND U6611 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U6612 ( .A(start_reg[389]), .B(init), .Z(start_in[389]) );
  AND U6613 ( .A(start_reg[388]), .B(init), .Z(start_in[388]) );
  AND U6614 ( .A(start_reg[387]), .B(init), .Z(start_in[387]) );
  AND U6615 ( .A(start_reg[386]), .B(init), .Z(start_in[386]) );
  AND U6616 ( .A(start_reg[385]), .B(init), .Z(start_in[385]) );
  AND U6617 ( .A(start_reg[384]), .B(init), .Z(start_in[384]) );
  AND U6618 ( .A(start_reg[383]), .B(init), .Z(start_in[383]) );
  AND U6619 ( .A(start_reg[382]), .B(init), .Z(start_in[382]) );
  AND U6620 ( .A(start_reg[381]), .B(init), .Z(start_in[381]) );
  AND U6621 ( .A(start_reg[380]), .B(init), .Z(start_in[380]) );
  AND U6622 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U6623 ( .A(start_reg[379]), .B(init), .Z(start_in[379]) );
  AND U6624 ( .A(start_reg[378]), .B(init), .Z(start_in[378]) );
  AND U6625 ( .A(start_reg[377]), .B(init), .Z(start_in[377]) );
  AND U6626 ( .A(start_reg[376]), .B(init), .Z(start_in[376]) );
  AND U6627 ( .A(start_reg[375]), .B(init), .Z(start_in[375]) );
  AND U6628 ( .A(start_reg[374]), .B(init), .Z(start_in[374]) );
  AND U6629 ( .A(start_reg[373]), .B(init), .Z(start_in[373]) );
  AND U6630 ( .A(start_reg[372]), .B(init), .Z(start_in[372]) );
  AND U6631 ( .A(start_reg[371]), .B(init), .Z(start_in[371]) );
  AND U6632 ( .A(start_reg[370]), .B(init), .Z(start_in[370]) );
  AND U6633 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U6634 ( .A(start_reg[369]), .B(init), .Z(start_in[369]) );
  AND U6635 ( .A(start_reg[368]), .B(init), .Z(start_in[368]) );
  AND U6636 ( .A(start_reg[367]), .B(init), .Z(start_in[367]) );
  AND U6637 ( .A(start_reg[366]), .B(init), .Z(start_in[366]) );
  AND U6638 ( .A(start_reg[365]), .B(init), .Z(start_in[365]) );
  AND U6639 ( .A(start_reg[364]), .B(init), .Z(start_in[364]) );
  AND U6640 ( .A(start_reg[363]), .B(init), .Z(start_in[363]) );
  AND U6641 ( .A(start_reg[362]), .B(init), .Z(start_in[362]) );
  AND U6642 ( .A(start_reg[361]), .B(init), .Z(start_in[361]) );
  AND U6643 ( .A(start_reg[360]), .B(init), .Z(start_in[360]) );
  AND U6644 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U6645 ( .A(start_reg[359]), .B(init), .Z(start_in[359]) );
  AND U6646 ( .A(start_reg[358]), .B(init), .Z(start_in[358]) );
  AND U6647 ( .A(start_reg[357]), .B(init), .Z(start_in[357]) );
  AND U6648 ( .A(start_reg[356]), .B(init), .Z(start_in[356]) );
  AND U6649 ( .A(start_reg[355]), .B(init), .Z(start_in[355]) );
  AND U6650 ( .A(start_reg[354]), .B(init), .Z(start_in[354]) );
  AND U6651 ( .A(start_reg[353]), .B(init), .Z(start_in[353]) );
  AND U6652 ( .A(start_reg[352]), .B(init), .Z(start_in[352]) );
  AND U6653 ( .A(start_reg[351]), .B(init), .Z(start_in[351]) );
  AND U6654 ( .A(start_reg[350]), .B(init), .Z(start_in[350]) );
  AND U6655 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U6656 ( .A(start_reg[349]), .B(init), .Z(start_in[349]) );
  AND U6657 ( .A(start_reg[348]), .B(init), .Z(start_in[348]) );
  AND U6658 ( .A(start_reg[347]), .B(init), .Z(start_in[347]) );
  AND U6659 ( .A(start_reg[346]), .B(init), .Z(start_in[346]) );
  AND U6660 ( .A(start_reg[345]), .B(init), .Z(start_in[345]) );
  AND U6661 ( .A(start_reg[344]), .B(init), .Z(start_in[344]) );
  AND U6662 ( .A(start_reg[343]), .B(init), .Z(start_in[343]) );
  AND U6663 ( .A(start_reg[342]), .B(init), .Z(start_in[342]) );
  AND U6664 ( .A(start_reg[341]), .B(init), .Z(start_in[341]) );
  AND U6665 ( .A(start_reg[340]), .B(init), .Z(start_in[340]) );
  AND U6666 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U6667 ( .A(start_reg[339]), .B(init), .Z(start_in[339]) );
  AND U6668 ( .A(start_reg[338]), .B(init), .Z(start_in[338]) );
  AND U6669 ( .A(start_reg[337]), .B(init), .Z(start_in[337]) );
  AND U6670 ( .A(start_reg[336]), .B(init), .Z(start_in[336]) );
  AND U6671 ( .A(start_reg[335]), .B(init), .Z(start_in[335]) );
  AND U6672 ( .A(start_reg[334]), .B(init), .Z(start_in[334]) );
  AND U6673 ( .A(start_reg[333]), .B(init), .Z(start_in[333]) );
  AND U6674 ( .A(start_reg[332]), .B(init), .Z(start_in[332]) );
  AND U6675 ( .A(start_reg[331]), .B(init), .Z(start_in[331]) );
  AND U6676 ( .A(start_reg[330]), .B(init), .Z(start_in[330]) );
  AND U6677 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U6678 ( .A(start_reg[329]), .B(init), .Z(start_in[329]) );
  AND U6679 ( .A(start_reg[328]), .B(init), .Z(start_in[328]) );
  AND U6680 ( .A(start_reg[327]), .B(init), .Z(start_in[327]) );
  AND U6681 ( .A(start_reg[326]), .B(init), .Z(start_in[326]) );
  AND U6682 ( .A(start_reg[325]), .B(init), .Z(start_in[325]) );
  AND U6683 ( .A(start_reg[324]), .B(init), .Z(start_in[324]) );
  AND U6684 ( .A(start_reg[323]), .B(init), .Z(start_in[323]) );
  AND U6685 ( .A(start_reg[322]), .B(init), .Z(start_in[322]) );
  AND U6686 ( .A(start_reg[321]), .B(init), .Z(start_in[321]) );
  AND U6687 ( .A(start_reg[320]), .B(init), .Z(start_in[320]) );
  AND U6688 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U6689 ( .A(start_reg[319]), .B(init), .Z(start_in[319]) );
  AND U6690 ( .A(start_reg[318]), .B(init), .Z(start_in[318]) );
  AND U6691 ( .A(start_reg[317]), .B(init), .Z(start_in[317]) );
  AND U6692 ( .A(start_reg[316]), .B(init), .Z(start_in[316]) );
  AND U6693 ( .A(start_reg[315]), .B(init), .Z(start_in[315]) );
  AND U6694 ( .A(start_reg[314]), .B(init), .Z(start_in[314]) );
  AND U6695 ( .A(start_reg[313]), .B(init), .Z(start_in[313]) );
  AND U6696 ( .A(start_reg[312]), .B(init), .Z(start_in[312]) );
  AND U6697 ( .A(start_reg[311]), .B(init), .Z(start_in[311]) );
  AND U6698 ( .A(start_reg[310]), .B(init), .Z(start_in[310]) );
  AND U6699 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U6700 ( .A(start_reg[309]), .B(init), .Z(start_in[309]) );
  AND U6701 ( .A(start_reg[308]), .B(init), .Z(start_in[308]) );
  AND U6702 ( .A(start_reg[307]), .B(init), .Z(start_in[307]) );
  AND U6703 ( .A(start_reg[306]), .B(init), .Z(start_in[306]) );
  AND U6704 ( .A(start_reg[305]), .B(init), .Z(start_in[305]) );
  AND U6705 ( .A(start_reg[304]), .B(init), .Z(start_in[304]) );
  AND U6706 ( .A(start_reg[303]), .B(init), .Z(start_in[303]) );
  AND U6707 ( .A(start_reg[302]), .B(init), .Z(start_in[302]) );
  AND U6708 ( .A(start_reg[301]), .B(init), .Z(start_in[301]) );
  AND U6709 ( .A(start_reg[300]), .B(init), .Z(start_in[300]) );
  AND U6710 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U6711 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U6712 ( .A(start_reg[299]), .B(init), .Z(start_in[299]) );
  AND U6713 ( .A(start_reg[298]), .B(init), .Z(start_in[298]) );
  AND U6714 ( .A(start_reg[297]), .B(init), .Z(start_in[297]) );
  AND U6715 ( .A(start_reg[296]), .B(init), .Z(start_in[296]) );
  AND U6716 ( .A(start_reg[295]), .B(init), .Z(start_in[295]) );
  AND U6717 ( .A(start_reg[294]), .B(init), .Z(start_in[294]) );
  AND U6718 ( .A(start_reg[293]), .B(init), .Z(start_in[293]) );
  AND U6719 ( .A(start_reg[292]), .B(init), .Z(start_in[292]) );
  AND U6720 ( .A(start_reg[291]), .B(init), .Z(start_in[291]) );
  AND U6721 ( .A(start_reg[290]), .B(init), .Z(start_in[290]) );
  AND U6722 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U6723 ( .A(start_reg[289]), .B(init), .Z(start_in[289]) );
  AND U6724 ( .A(start_reg[288]), .B(init), .Z(start_in[288]) );
  AND U6725 ( .A(start_reg[287]), .B(init), .Z(start_in[287]) );
  AND U6726 ( .A(start_reg[286]), .B(init), .Z(start_in[286]) );
  AND U6727 ( .A(start_reg[285]), .B(init), .Z(start_in[285]) );
  AND U6728 ( .A(start_reg[284]), .B(init), .Z(start_in[284]) );
  AND U6729 ( .A(start_reg[283]), .B(init), .Z(start_in[283]) );
  AND U6730 ( .A(start_reg[282]), .B(init), .Z(start_in[282]) );
  AND U6731 ( .A(start_reg[281]), .B(init), .Z(start_in[281]) );
  AND U6732 ( .A(start_reg[280]), .B(init), .Z(start_in[280]) );
  AND U6733 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U6734 ( .A(start_reg[279]), .B(init), .Z(start_in[279]) );
  AND U6735 ( .A(start_reg[278]), .B(init), .Z(start_in[278]) );
  AND U6736 ( .A(start_reg[277]), .B(init), .Z(start_in[277]) );
  AND U6737 ( .A(start_reg[276]), .B(init), .Z(start_in[276]) );
  AND U6738 ( .A(start_reg[275]), .B(init), .Z(start_in[275]) );
  AND U6739 ( .A(start_reg[274]), .B(init), .Z(start_in[274]) );
  AND U6740 ( .A(start_reg[273]), .B(init), .Z(start_in[273]) );
  AND U6741 ( .A(start_reg[272]), .B(init), .Z(start_in[272]) );
  AND U6742 ( .A(start_reg[271]), .B(init), .Z(start_in[271]) );
  AND U6743 ( .A(start_reg[270]), .B(init), .Z(start_in[270]) );
  AND U6744 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U6745 ( .A(start_reg[269]), .B(init), .Z(start_in[269]) );
  AND U6746 ( .A(start_reg[268]), .B(init), .Z(start_in[268]) );
  AND U6747 ( .A(start_reg[267]), .B(init), .Z(start_in[267]) );
  AND U6748 ( .A(start_reg[266]), .B(init), .Z(start_in[266]) );
  AND U6749 ( .A(start_reg[265]), .B(init), .Z(start_in[265]) );
  AND U6750 ( .A(start_reg[264]), .B(init), .Z(start_in[264]) );
  AND U6751 ( .A(start_reg[263]), .B(init), .Z(start_in[263]) );
  AND U6752 ( .A(start_reg[262]), .B(init), .Z(start_in[262]) );
  AND U6753 ( .A(start_reg[261]), .B(init), .Z(start_in[261]) );
  AND U6754 ( .A(start_reg[260]), .B(init), .Z(start_in[260]) );
  AND U6755 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U6756 ( .A(start_reg[259]), .B(init), .Z(start_in[259]) );
  AND U6757 ( .A(start_reg[258]), .B(init), .Z(start_in[258]) );
  AND U6758 ( .A(start_reg[257]), .B(init), .Z(start_in[257]) );
  AND U6759 ( .A(start_reg[256]), .B(init), .Z(start_in[256]) );
  AND U6760 ( .A(start_reg[255]), .B(init), .Z(start_in[255]) );
  AND U6761 ( .A(start_reg[254]), .B(init), .Z(start_in[254]) );
  AND U6762 ( .A(start_reg[253]), .B(init), .Z(start_in[253]) );
  AND U6763 ( .A(start_reg[252]), .B(init), .Z(start_in[252]) );
  AND U6764 ( .A(start_reg[251]), .B(init), .Z(start_in[251]) );
  AND U6765 ( .A(start_reg[250]), .B(init), .Z(start_in[250]) );
  AND U6766 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U6767 ( .A(start_reg[249]), .B(init), .Z(start_in[249]) );
  AND U6768 ( .A(start_reg[248]), .B(init), .Z(start_in[248]) );
  AND U6769 ( .A(start_reg[247]), .B(init), .Z(start_in[247]) );
  AND U6770 ( .A(start_reg[246]), .B(init), .Z(start_in[246]) );
  AND U6771 ( .A(start_reg[245]), .B(init), .Z(start_in[245]) );
  AND U6772 ( .A(start_reg[244]), .B(init), .Z(start_in[244]) );
  AND U6773 ( .A(start_reg[243]), .B(init), .Z(start_in[243]) );
  AND U6774 ( .A(start_reg[242]), .B(init), .Z(start_in[242]) );
  AND U6775 ( .A(start_reg[241]), .B(init), .Z(start_in[241]) );
  AND U6776 ( .A(start_reg[240]), .B(init), .Z(start_in[240]) );
  AND U6777 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U6778 ( .A(start_reg[239]), .B(init), .Z(start_in[239]) );
  AND U6779 ( .A(start_reg[238]), .B(init), .Z(start_in[238]) );
  AND U6780 ( .A(start_reg[237]), .B(init), .Z(start_in[237]) );
  AND U6781 ( .A(start_reg[236]), .B(init), .Z(start_in[236]) );
  AND U6782 ( .A(start_reg[235]), .B(init), .Z(start_in[235]) );
  AND U6783 ( .A(start_reg[234]), .B(init), .Z(start_in[234]) );
  AND U6784 ( .A(start_reg[233]), .B(init), .Z(start_in[233]) );
  AND U6785 ( .A(start_reg[232]), .B(init), .Z(start_in[232]) );
  AND U6786 ( .A(start_reg[231]), .B(init), .Z(start_in[231]) );
  AND U6787 ( .A(start_reg[230]), .B(init), .Z(start_in[230]) );
  AND U6788 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U6789 ( .A(start_reg[229]), .B(init), .Z(start_in[229]) );
  AND U6790 ( .A(start_reg[228]), .B(init), .Z(start_in[228]) );
  AND U6791 ( .A(start_reg[227]), .B(init), .Z(start_in[227]) );
  AND U6792 ( .A(start_reg[226]), .B(init), .Z(start_in[226]) );
  AND U6793 ( .A(start_reg[225]), .B(init), .Z(start_in[225]) );
  AND U6794 ( .A(start_reg[224]), .B(init), .Z(start_in[224]) );
  AND U6795 ( .A(start_reg[223]), .B(init), .Z(start_in[223]) );
  AND U6796 ( .A(start_reg[222]), .B(init), .Z(start_in[222]) );
  AND U6797 ( .A(start_reg[221]), .B(init), .Z(start_in[221]) );
  AND U6798 ( .A(start_reg[220]), .B(init), .Z(start_in[220]) );
  AND U6799 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U6800 ( .A(start_reg[219]), .B(init), .Z(start_in[219]) );
  AND U6801 ( .A(start_reg[218]), .B(init), .Z(start_in[218]) );
  AND U6802 ( .A(start_reg[217]), .B(init), .Z(start_in[217]) );
  AND U6803 ( .A(start_reg[216]), .B(init), .Z(start_in[216]) );
  AND U6804 ( .A(start_reg[215]), .B(init), .Z(start_in[215]) );
  AND U6805 ( .A(start_reg[214]), .B(init), .Z(start_in[214]) );
  AND U6806 ( .A(start_reg[213]), .B(init), .Z(start_in[213]) );
  AND U6807 ( .A(start_reg[212]), .B(init), .Z(start_in[212]) );
  AND U6808 ( .A(start_reg[211]), .B(init), .Z(start_in[211]) );
  AND U6809 ( .A(start_reg[210]), .B(init), .Z(start_in[210]) );
  AND U6810 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U6811 ( .A(start_reg[209]), .B(init), .Z(start_in[209]) );
  AND U6812 ( .A(start_reg[208]), .B(init), .Z(start_in[208]) );
  AND U6813 ( .A(start_reg[207]), .B(init), .Z(start_in[207]) );
  AND U6814 ( .A(start_reg[206]), .B(init), .Z(start_in[206]) );
  AND U6815 ( .A(start_reg[205]), .B(init), .Z(start_in[205]) );
  AND U6816 ( .A(start_reg[204]), .B(init), .Z(start_in[204]) );
  AND U6817 ( .A(start_reg[203]), .B(init), .Z(start_in[203]) );
  AND U6818 ( .A(start_reg[202]), .B(init), .Z(start_in[202]) );
  AND U6819 ( .A(start_reg[201]), .B(init), .Z(start_in[201]) );
  AND U6820 ( .A(start_reg[200]), .B(init), .Z(start_in[200]) );
  AND U6821 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U6822 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U6823 ( .A(start_reg[199]), .B(init), .Z(start_in[199]) );
  AND U6824 ( .A(start_reg[198]), .B(init), .Z(start_in[198]) );
  AND U6825 ( .A(start_reg[197]), .B(init), .Z(start_in[197]) );
  AND U6826 ( .A(start_reg[196]), .B(init), .Z(start_in[196]) );
  AND U6827 ( .A(start_reg[195]), .B(init), .Z(start_in[195]) );
  AND U6828 ( .A(start_reg[194]), .B(init), .Z(start_in[194]) );
  AND U6829 ( .A(start_reg[193]), .B(init), .Z(start_in[193]) );
  AND U6830 ( .A(start_reg[192]), .B(init), .Z(start_in[192]) );
  AND U6831 ( .A(start_reg[191]), .B(init), .Z(start_in[191]) );
  AND U6832 ( .A(start_reg[190]), .B(init), .Z(start_in[190]) );
  AND U6833 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U6834 ( .A(start_reg[189]), .B(init), .Z(start_in[189]) );
  AND U6835 ( .A(start_reg[188]), .B(init), .Z(start_in[188]) );
  AND U6836 ( .A(start_reg[187]), .B(init), .Z(start_in[187]) );
  AND U6837 ( .A(start_reg[186]), .B(init), .Z(start_in[186]) );
  AND U6838 ( .A(start_reg[185]), .B(init), .Z(start_in[185]) );
  AND U6839 ( .A(start_reg[184]), .B(init), .Z(start_in[184]) );
  AND U6840 ( .A(start_reg[183]), .B(init), .Z(start_in[183]) );
  AND U6841 ( .A(start_reg[182]), .B(init), .Z(start_in[182]) );
  AND U6842 ( .A(start_reg[181]), .B(init), .Z(start_in[181]) );
  AND U6843 ( .A(start_reg[180]), .B(init), .Z(start_in[180]) );
  AND U6844 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U6845 ( .A(start_reg[179]), .B(init), .Z(start_in[179]) );
  AND U6846 ( .A(start_reg[178]), .B(init), .Z(start_in[178]) );
  AND U6847 ( .A(start_reg[177]), .B(init), .Z(start_in[177]) );
  AND U6848 ( .A(start_reg[176]), .B(init), .Z(start_in[176]) );
  AND U6849 ( .A(start_reg[175]), .B(init), .Z(start_in[175]) );
  AND U6850 ( .A(start_reg[174]), .B(init), .Z(start_in[174]) );
  AND U6851 ( .A(start_reg[173]), .B(init), .Z(start_in[173]) );
  AND U6852 ( .A(start_reg[172]), .B(init), .Z(start_in[172]) );
  AND U6853 ( .A(start_reg[171]), .B(init), .Z(start_in[171]) );
  AND U6854 ( .A(start_reg[170]), .B(init), .Z(start_in[170]) );
  AND U6855 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U6856 ( .A(start_reg[169]), .B(init), .Z(start_in[169]) );
  AND U6857 ( .A(start_reg[168]), .B(init), .Z(start_in[168]) );
  AND U6858 ( .A(start_reg[167]), .B(init), .Z(start_in[167]) );
  AND U6859 ( .A(start_reg[166]), .B(init), .Z(start_in[166]) );
  AND U6860 ( .A(start_reg[165]), .B(init), .Z(start_in[165]) );
  AND U6861 ( .A(start_reg[164]), .B(init), .Z(start_in[164]) );
  AND U6862 ( .A(start_reg[163]), .B(init), .Z(start_in[163]) );
  AND U6863 ( .A(start_reg[162]), .B(init), .Z(start_in[162]) );
  AND U6864 ( .A(start_reg[161]), .B(init), .Z(start_in[161]) );
  AND U6865 ( .A(start_reg[160]), .B(init), .Z(start_in[160]) );
  AND U6866 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U6867 ( .A(start_reg[159]), .B(init), .Z(start_in[159]) );
  AND U6868 ( .A(start_reg[158]), .B(init), .Z(start_in[158]) );
  AND U6869 ( .A(start_reg[157]), .B(init), .Z(start_in[157]) );
  AND U6870 ( .A(start_reg[156]), .B(init), .Z(start_in[156]) );
  AND U6871 ( .A(start_reg[155]), .B(init), .Z(start_in[155]) );
  AND U6872 ( .A(start_reg[154]), .B(init), .Z(start_in[154]) );
  AND U6873 ( .A(start_reg[153]), .B(init), .Z(start_in[153]) );
  AND U6874 ( .A(start_reg[152]), .B(init), .Z(start_in[152]) );
  AND U6875 ( .A(start_reg[151]), .B(init), .Z(start_in[151]) );
  AND U6876 ( .A(start_reg[150]), .B(init), .Z(start_in[150]) );
  AND U6877 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U6878 ( .A(start_reg[149]), .B(init), .Z(start_in[149]) );
  AND U6879 ( .A(start_reg[148]), .B(init), .Z(start_in[148]) );
  AND U6880 ( .A(start_reg[147]), .B(init), .Z(start_in[147]) );
  AND U6881 ( .A(start_reg[146]), .B(init), .Z(start_in[146]) );
  AND U6882 ( .A(start_reg[145]), .B(init), .Z(start_in[145]) );
  AND U6883 ( .A(start_reg[144]), .B(init), .Z(start_in[144]) );
  AND U6884 ( .A(start_reg[143]), .B(init), .Z(start_in[143]) );
  AND U6885 ( .A(start_reg[142]), .B(init), .Z(start_in[142]) );
  AND U6886 ( .A(start_reg[141]), .B(init), .Z(start_in[141]) );
  AND U6887 ( .A(start_reg[140]), .B(init), .Z(start_in[140]) );
  AND U6888 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U6889 ( .A(start_reg[139]), .B(init), .Z(start_in[139]) );
  AND U6890 ( .A(start_reg[138]), .B(init), .Z(start_in[138]) );
  AND U6891 ( .A(start_reg[137]), .B(init), .Z(start_in[137]) );
  AND U6892 ( .A(start_reg[136]), .B(init), .Z(start_in[136]) );
  AND U6893 ( .A(start_reg[135]), .B(init), .Z(start_in[135]) );
  AND U6894 ( .A(start_reg[134]), .B(init), .Z(start_in[134]) );
  AND U6895 ( .A(start_reg[133]), .B(init), .Z(start_in[133]) );
  AND U6896 ( .A(start_reg[132]), .B(init), .Z(start_in[132]) );
  AND U6897 ( .A(start_reg[131]), .B(init), .Z(start_in[131]) );
  AND U6898 ( .A(start_reg[130]), .B(init), .Z(start_in[130]) );
  AND U6899 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U6900 ( .A(start_reg[129]), .B(init), .Z(start_in[129]) );
  AND U6901 ( .A(start_reg[128]), .B(init), .Z(start_in[128]) );
  AND U6902 ( .A(start_reg[127]), .B(init), .Z(start_in[127]) );
  AND U6903 ( .A(start_reg[126]), .B(init), .Z(start_in[126]) );
  AND U6904 ( .A(start_reg[125]), .B(init), .Z(start_in[125]) );
  AND U6905 ( .A(start_reg[124]), .B(init), .Z(start_in[124]) );
  AND U6906 ( .A(start_reg[123]), .B(init), .Z(start_in[123]) );
  AND U6907 ( .A(start_reg[122]), .B(init), .Z(start_in[122]) );
  AND U6908 ( .A(start_reg[121]), .B(init), .Z(start_in[121]) );
  AND U6909 ( .A(start_reg[120]), .B(init), .Z(start_in[120]) );
  AND U6910 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U6911 ( .A(start_reg[119]), .B(init), .Z(start_in[119]) );
  AND U6912 ( .A(start_reg[118]), .B(init), .Z(start_in[118]) );
  AND U6913 ( .A(start_reg[117]), .B(init), .Z(start_in[117]) );
  AND U6914 ( .A(start_reg[116]), .B(init), .Z(start_in[116]) );
  AND U6915 ( .A(start_reg[115]), .B(init), .Z(start_in[115]) );
  AND U6916 ( .A(start_reg[114]), .B(init), .Z(start_in[114]) );
  AND U6917 ( .A(start_reg[113]), .B(init), .Z(start_in[113]) );
  AND U6918 ( .A(start_reg[112]), .B(init), .Z(start_in[112]) );
  AND U6919 ( .A(start_reg[111]), .B(init), .Z(start_in[111]) );
  AND U6920 ( .A(start_reg[110]), .B(init), .Z(start_in[110]) );
  AND U6921 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  AND U6922 ( .A(start_reg[109]), .B(init), .Z(start_in[109]) );
  AND U6923 ( .A(start_reg[108]), .B(init), .Z(start_in[108]) );
  AND U6924 ( .A(start_reg[107]), .B(init), .Z(start_in[107]) );
  AND U6925 ( .A(start_reg[106]), .B(init), .Z(start_in[106]) );
  AND U6926 ( .A(start_reg[105]), .B(init), .Z(start_in[105]) );
  AND U6927 ( .A(start_reg[104]), .B(init), .Z(start_in[104]) );
  AND U6928 ( .A(start_reg[103]), .B(init), .Z(start_in[103]) );
  AND U6929 ( .A(start_reg[102]), .B(init), .Z(start_in[102]) );
  AND U6930 ( .A(start_reg[101]), .B(init), .Z(start_in[101]) );
  AND U6931 ( .A(start_reg[100]), .B(init), .Z(start_in[100]) );
  NANDN U6932 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  NAND U6933 ( .A(n4886), .B(n4887), .Z(n3859) );
  NAND U6934 ( .A(n3863), .B(start_reg[511]), .Z(n4887) );
  IV U6935 ( .A(n3862), .Z(n3863) );
  NANDN U6936 ( .A(start_in[511]), .B(mul_pow), .Z(n4886) );
  NAND U6937 ( .A(n4888), .B(n4889), .Z(n3858) );
  NANDN U6938 ( .A(n4890), .B(ereg[0]), .Z(n4889) );
  NANDN U6939 ( .A(init), .B(e[0]), .Z(n4888) );
  NAND U6940 ( .A(n4891), .B(n4892), .Z(n3857) );
  NANDN U6941 ( .A(init), .B(e[1]), .Z(n4892) );
  AND U6942 ( .A(n4893), .B(n4894), .Z(n4891) );
  NAND U6943 ( .A(n4895), .B(ereg[0]), .Z(n4894) );
  NANDN U6944 ( .A(n4890), .B(ereg[1]), .Z(n4893) );
  NAND U6945 ( .A(n4896), .B(n4897), .Z(n3856) );
  NANDN U6946 ( .A(init), .B(e[2]), .Z(n4897) );
  AND U6947 ( .A(n4898), .B(n4899), .Z(n4896) );
  NAND U6948 ( .A(ereg[1]), .B(n4895), .Z(n4899) );
  NANDN U6949 ( .A(n4890), .B(ereg[2]), .Z(n4898) );
  NAND U6950 ( .A(n4900), .B(n4901), .Z(n3855) );
  NANDN U6951 ( .A(init), .B(e[3]), .Z(n4901) );
  AND U6952 ( .A(n4902), .B(n4903), .Z(n4900) );
  NAND U6953 ( .A(ereg[2]), .B(n4895), .Z(n4903) );
  NANDN U6954 ( .A(n4890), .B(ereg[3]), .Z(n4902) );
  NAND U6955 ( .A(n4904), .B(n4905), .Z(n3854) );
  NANDN U6956 ( .A(init), .B(e[4]), .Z(n4905) );
  AND U6957 ( .A(n4906), .B(n4907), .Z(n4904) );
  NAND U6958 ( .A(ereg[3]), .B(n4895), .Z(n4907) );
  NANDN U6959 ( .A(n4890), .B(ereg[4]), .Z(n4906) );
  NAND U6960 ( .A(n4908), .B(n4909), .Z(n3853) );
  NANDN U6961 ( .A(init), .B(e[5]), .Z(n4909) );
  AND U6962 ( .A(n4910), .B(n4911), .Z(n4908) );
  NAND U6963 ( .A(ereg[4]), .B(n4895), .Z(n4911) );
  NANDN U6964 ( .A(n4890), .B(ereg[5]), .Z(n4910) );
  NAND U6965 ( .A(n4912), .B(n4913), .Z(n3852) );
  NANDN U6966 ( .A(init), .B(e[6]), .Z(n4913) );
  AND U6967 ( .A(n4914), .B(n4915), .Z(n4912) );
  NAND U6968 ( .A(ereg[5]), .B(n4895), .Z(n4915) );
  NANDN U6969 ( .A(n4890), .B(ereg[6]), .Z(n4914) );
  NAND U6970 ( .A(n4916), .B(n4917), .Z(n3851) );
  NANDN U6971 ( .A(init), .B(e[7]), .Z(n4917) );
  AND U6972 ( .A(n4918), .B(n4919), .Z(n4916) );
  NAND U6973 ( .A(ereg[6]), .B(n4895), .Z(n4919) );
  NANDN U6974 ( .A(n4890), .B(ereg[7]), .Z(n4918) );
  NAND U6975 ( .A(n4920), .B(n4921), .Z(n3850) );
  NANDN U6976 ( .A(init), .B(e[8]), .Z(n4921) );
  AND U6977 ( .A(n4922), .B(n4923), .Z(n4920) );
  NAND U6978 ( .A(ereg[7]), .B(n4895), .Z(n4923) );
  NANDN U6979 ( .A(n4890), .B(ereg[8]), .Z(n4922) );
  NAND U6980 ( .A(n4924), .B(n4925), .Z(n3849) );
  NANDN U6981 ( .A(init), .B(e[9]), .Z(n4925) );
  AND U6982 ( .A(n4926), .B(n4927), .Z(n4924) );
  NAND U6983 ( .A(ereg[8]), .B(n4895), .Z(n4927) );
  NANDN U6984 ( .A(n4890), .B(ereg[9]), .Z(n4926) );
  NAND U6985 ( .A(n4928), .B(n4929), .Z(n3848) );
  NANDN U6986 ( .A(init), .B(e[10]), .Z(n4929) );
  AND U6987 ( .A(n4930), .B(n4931), .Z(n4928) );
  NAND U6988 ( .A(ereg[9]), .B(n4895), .Z(n4931) );
  NANDN U6989 ( .A(n4890), .B(ereg[10]), .Z(n4930) );
  NAND U6990 ( .A(n4932), .B(n4933), .Z(n3847) );
  NANDN U6991 ( .A(init), .B(e[11]), .Z(n4933) );
  AND U6992 ( .A(n4934), .B(n4935), .Z(n4932) );
  NAND U6993 ( .A(ereg[10]), .B(n4895), .Z(n4935) );
  NANDN U6994 ( .A(n4890), .B(ereg[11]), .Z(n4934) );
  NAND U6995 ( .A(n4936), .B(n4937), .Z(n3846) );
  NANDN U6996 ( .A(init), .B(e[12]), .Z(n4937) );
  AND U6997 ( .A(n4938), .B(n4939), .Z(n4936) );
  NAND U6998 ( .A(ereg[11]), .B(n4895), .Z(n4939) );
  NANDN U6999 ( .A(n4890), .B(ereg[12]), .Z(n4938) );
  NAND U7000 ( .A(n4940), .B(n4941), .Z(n3845) );
  NANDN U7001 ( .A(init), .B(e[13]), .Z(n4941) );
  AND U7002 ( .A(n4942), .B(n4943), .Z(n4940) );
  NAND U7003 ( .A(ereg[12]), .B(n4895), .Z(n4943) );
  NANDN U7004 ( .A(n4890), .B(ereg[13]), .Z(n4942) );
  NAND U7005 ( .A(n4944), .B(n4945), .Z(n3844) );
  NANDN U7006 ( .A(init), .B(e[14]), .Z(n4945) );
  AND U7007 ( .A(n4946), .B(n4947), .Z(n4944) );
  NAND U7008 ( .A(ereg[13]), .B(n4895), .Z(n4947) );
  NANDN U7009 ( .A(n4890), .B(ereg[14]), .Z(n4946) );
  NAND U7010 ( .A(n4948), .B(n4949), .Z(n3843) );
  NANDN U7011 ( .A(init), .B(e[15]), .Z(n4949) );
  AND U7012 ( .A(n4950), .B(n4951), .Z(n4948) );
  NAND U7013 ( .A(ereg[14]), .B(n4895), .Z(n4951) );
  NANDN U7014 ( .A(n4890), .B(ereg[15]), .Z(n4950) );
  NAND U7015 ( .A(n4952), .B(n4953), .Z(n3842) );
  NANDN U7016 ( .A(init), .B(e[16]), .Z(n4953) );
  AND U7017 ( .A(n4954), .B(n4955), .Z(n4952) );
  NAND U7018 ( .A(ereg[15]), .B(n4895), .Z(n4955) );
  NANDN U7019 ( .A(n4890), .B(ereg[16]), .Z(n4954) );
  NAND U7020 ( .A(n4956), .B(n4957), .Z(n3841) );
  NANDN U7021 ( .A(init), .B(e[17]), .Z(n4957) );
  AND U7022 ( .A(n4958), .B(n4959), .Z(n4956) );
  NAND U7023 ( .A(ereg[16]), .B(n4895), .Z(n4959) );
  NANDN U7024 ( .A(n4890), .B(ereg[17]), .Z(n4958) );
  NAND U7025 ( .A(n4960), .B(n4961), .Z(n3840) );
  NANDN U7026 ( .A(init), .B(e[18]), .Z(n4961) );
  AND U7027 ( .A(n4962), .B(n4963), .Z(n4960) );
  NAND U7028 ( .A(ereg[17]), .B(n4895), .Z(n4963) );
  NANDN U7029 ( .A(n4890), .B(ereg[18]), .Z(n4962) );
  NAND U7030 ( .A(n4964), .B(n4965), .Z(n3839) );
  NANDN U7031 ( .A(init), .B(e[19]), .Z(n4965) );
  AND U7032 ( .A(n4966), .B(n4967), .Z(n4964) );
  NAND U7033 ( .A(ereg[18]), .B(n4895), .Z(n4967) );
  NANDN U7034 ( .A(n4890), .B(ereg[19]), .Z(n4966) );
  NAND U7035 ( .A(n4968), .B(n4969), .Z(n3838) );
  NANDN U7036 ( .A(init), .B(e[20]), .Z(n4969) );
  AND U7037 ( .A(n4970), .B(n4971), .Z(n4968) );
  NAND U7038 ( .A(ereg[19]), .B(n4895), .Z(n4971) );
  NANDN U7039 ( .A(n4890), .B(ereg[20]), .Z(n4970) );
  NAND U7040 ( .A(n4972), .B(n4973), .Z(n3837) );
  NANDN U7041 ( .A(init), .B(e[21]), .Z(n4973) );
  AND U7042 ( .A(n4974), .B(n4975), .Z(n4972) );
  NAND U7043 ( .A(ereg[20]), .B(n4895), .Z(n4975) );
  NANDN U7044 ( .A(n4890), .B(ereg[21]), .Z(n4974) );
  NAND U7045 ( .A(n4976), .B(n4977), .Z(n3836) );
  NANDN U7046 ( .A(init), .B(e[22]), .Z(n4977) );
  AND U7047 ( .A(n4978), .B(n4979), .Z(n4976) );
  NAND U7048 ( .A(ereg[21]), .B(n4895), .Z(n4979) );
  NANDN U7049 ( .A(n4890), .B(ereg[22]), .Z(n4978) );
  NAND U7050 ( .A(n4980), .B(n4981), .Z(n3835) );
  NANDN U7051 ( .A(init), .B(e[23]), .Z(n4981) );
  AND U7052 ( .A(n4982), .B(n4983), .Z(n4980) );
  NAND U7053 ( .A(ereg[22]), .B(n4895), .Z(n4983) );
  NANDN U7054 ( .A(n4890), .B(ereg[23]), .Z(n4982) );
  NAND U7055 ( .A(n4984), .B(n4985), .Z(n3834) );
  NANDN U7056 ( .A(init), .B(e[24]), .Z(n4985) );
  AND U7057 ( .A(n4986), .B(n4987), .Z(n4984) );
  NAND U7058 ( .A(ereg[23]), .B(n4895), .Z(n4987) );
  NANDN U7059 ( .A(n4890), .B(ereg[24]), .Z(n4986) );
  NAND U7060 ( .A(n4988), .B(n4989), .Z(n3833) );
  NANDN U7061 ( .A(init), .B(e[25]), .Z(n4989) );
  AND U7062 ( .A(n4990), .B(n4991), .Z(n4988) );
  NAND U7063 ( .A(ereg[24]), .B(n4895), .Z(n4991) );
  NANDN U7064 ( .A(n4890), .B(ereg[25]), .Z(n4990) );
  NAND U7065 ( .A(n4992), .B(n4993), .Z(n3832) );
  NANDN U7066 ( .A(init), .B(e[26]), .Z(n4993) );
  AND U7067 ( .A(n4994), .B(n4995), .Z(n4992) );
  NAND U7068 ( .A(ereg[25]), .B(n4895), .Z(n4995) );
  NANDN U7069 ( .A(n4890), .B(ereg[26]), .Z(n4994) );
  NAND U7070 ( .A(n4996), .B(n4997), .Z(n3831) );
  NANDN U7071 ( .A(init), .B(e[27]), .Z(n4997) );
  AND U7072 ( .A(n4998), .B(n4999), .Z(n4996) );
  NAND U7073 ( .A(ereg[26]), .B(n4895), .Z(n4999) );
  NANDN U7074 ( .A(n4890), .B(ereg[27]), .Z(n4998) );
  NAND U7075 ( .A(n5000), .B(n5001), .Z(n3830) );
  NANDN U7076 ( .A(init), .B(e[28]), .Z(n5001) );
  AND U7077 ( .A(n5002), .B(n5003), .Z(n5000) );
  NAND U7078 ( .A(ereg[27]), .B(n4895), .Z(n5003) );
  NANDN U7079 ( .A(n4890), .B(ereg[28]), .Z(n5002) );
  NAND U7080 ( .A(n5004), .B(n5005), .Z(n3829) );
  NANDN U7081 ( .A(init), .B(e[29]), .Z(n5005) );
  AND U7082 ( .A(n5006), .B(n5007), .Z(n5004) );
  NAND U7083 ( .A(ereg[28]), .B(n4895), .Z(n5007) );
  NANDN U7084 ( .A(n4890), .B(ereg[29]), .Z(n5006) );
  NAND U7085 ( .A(n5008), .B(n5009), .Z(n3828) );
  NANDN U7086 ( .A(init), .B(e[30]), .Z(n5009) );
  AND U7087 ( .A(n5010), .B(n5011), .Z(n5008) );
  NAND U7088 ( .A(ereg[29]), .B(n4895), .Z(n5011) );
  NANDN U7089 ( .A(n4890), .B(ereg[30]), .Z(n5010) );
  NAND U7090 ( .A(n5012), .B(n5013), .Z(n3827) );
  NANDN U7091 ( .A(init), .B(e[31]), .Z(n5013) );
  AND U7092 ( .A(n5014), .B(n5015), .Z(n5012) );
  NAND U7093 ( .A(ereg[30]), .B(n4895), .Z(n5015) );
  NANDN U7094 ( .A(n4890), .B(ereg[31]), .Z(n5014) );
  NAND U7095 ( .A(n5016), .B(n5017), .Z(n3826) );
  NANDN U7096 ( .A(init), .B(e[32]), .Z(n5017) );
  AND U7097 ( .A(n5018), .B(n5019), .Z(n5016) );
  NAND U7098 ( .A(ereg[31]), .B(n4895), .Z(n5019) );
  NANDN U7099 ( .A(n4890), .B(ereg[32]), .Z(n5018) );
  NAND U7100 ( .A(n5020), .B(n5021), .Z(n3825) );
  NANDN U7101 ( .A(init), .B(e[33]), .Z(n5021) );
  AND U7102 ( .A(n5022), .B(n5023), .Z(n5020) );
  NAND U7103 ( .A(ereg[32]), .B(n4895), .Z(n5023) );
  NANDN U7104 ( .A(n4890), .B(ereg[33]), .Z(n5022) );
  NAND U7105 ( .A(n5024), .B(n5025), .Z(n3824) );
  NANDN U7106 ( .A(init), .B(e[34]), .Z(n5025) );
  AND U7107 ( .A(n5026), .B(n5027), .Z(n5024) );
  NAND U7108 ( .A(ereg[33]), .B(n4895), .Z(n5027) );
  NANDN U7109 ( .A(n4890), .B(ereg[34]), .Z(n5026) );
  NAND U7110 ( .A(n5028), .B(n5029), .Z(n3823) );
  NANDN U7111 ( .A(init), .B(e[35]), .Z(n5029) );
  AND U7112 ( .A(n5030), .B(n5031), .Z(n5028) );
  NAND U7113 ( .A(ereg[34]), .B(n4895), .Z(n5031) );
  NANDN U7114 ( .A(n4890), .B(ereg[35]), .Z(n5030) );
  NAND U7115 ( .A(n5032), .B(n5033), .Z(n3822) );
  NANDN U7116 ( .A(init), .B(e[36]), .Z(n5033) );
  AND U7117 ( .A(n5034), .B(n5035), .Z(n5032) );
  NAND U7118 ( .A(ereg[35]), .B(n4895), .Z(n5035) );
  NANDN U7119 ( .A(n4890), .B(ereg[36]), .Z(n5034) );
  NAND U7120 ( .A(n5036), .B(n5037), .Z(n3821) );
  NANDN U7121 ( .A(init), .B(e[37]), .Z(n5037) );
  AND U7122 ( .A(n5038), .B(n5039), .Z(n5036) );
  NAND U7123 ( .A(ereg[36]), .B(n4895), .Z(n5039) );
  NANDN U7124 ( .A(n4890), .B(ereg[37]), .Z(n5038) );
  NAND U7125 ( .A(n5040), .B(n5041), .Z(n3820) );
  NANDN U7126 ( .A(init), .B(e[38]), .Z(n5041) );
  AND U7127 ( .A(n5042), .B(n5043), .Z(n5040) );
  NAND U7128 ( .A(ereg[37]), .B(n4895), .Z(n5043) );
  NANDN U7129 ( .A(n4890), .B(ereg[38]), .Z(n5042) );
  NAND U7130 ( .A(n5044), .B(n5045), .Z(n3819) );
  NANDN U7131 ( .A(init), .B(e[39]), .Z(n5045) );
  AND U7132 ( .A(n5046), .B(n5047), .Z(n5044) );
  NAND U7133 ( .A(ereg[38]), .B(n4895), .Z(n5047) );
  NANDN U7134 ( .A(n4890), .B(ereg[39]), .Z(n5046) );
  NAND U7135 ( .A(n5048), .B(n5049), .Z(n3818) );
  NANDN U7136 ( .A(init), .B(e[40]), .Z(n5049) );
  AND U7137 ( .A(n5050), .B(n5051), .Z(n5048) );
  NAND U7138 ( .A(ereg[39]), .B(n4895), .Z(n5051) );
  NANDN U7139 ( .A(n4890), .B(ereg[40]), .Z(n5050) );
  NAND U7140 ( .A(n5052), .B(n5053), .Z(n3817) );
  NANDN U7141 ( .A(init), .B(e[41]), .Z(n5053) );
  AND U7142 ( .A(n5054), .B(n5055), .Z(n5052) );
  NAND U7143 ( .A(ereg[40]), .B(n4895), .Z(n5055) );
  NANDN U7144 ( .A(n4890), .B(ereg[41]), .Z(n5054) );
  NAND U7145 ( .A(n5056), .B(n5057), .Z(n3816) );
  NANDN U7146 ( .A(init), .B(e[42]), .Z(n5057) );
  AND U7147 ( .A(n5058), .B(n5059), .Z(n5056) );
  NAND U7148 ( .A(ereg[41]), .B(n4895), .Z(n5059) );
  NANDN U7149 ( .A(n4890), .B(ereg[42]), .Z(n5058) );
  NAND U7150 ( .A(n5060), .B(n5061), .Z(n3815) );
  NANDN U7151 ( .A(init), .B(e[43]), .Z(n5061) );
  AND U7152 ( .A(n5062), .B(n5063), .Z(n5060) );
  NAND U7153 ( .A(ereg[42]), .B(n4895), .Z(n5063) );
  NANDN U7154 ( .A(n4890), .B(ereg[43]), .Z(n5062) );
  NAND U7155 ( .A(n5064), .B(n5065), .Z(n3814) );
  NANDN U7156 ( .A(init), .B(e[44]), .Z(n5065) );
  AND U7157 ( .A(n5066), .B(n5067), .Z(n5064) );
  NAND U7158 ( .A(ereg[43]), .B(n4895), .Z(n5067) );
  NANDN U7159 ( .A(n4890), .B(ereg[44]), .Z(n5066) );
  NAND U7160 ( .A(n5068), .B(n5069), .Z(n3813) );
  NANDN U7161 ( .A(init), .B(e[45]), .Z(n5069) );
  AND U7162 ( .A(n5070), .B(n5071), .Z(n5068) );
  NAND U7163 ( .A(ereg[44]), .B(n4895), .Z(n5071) );
  NANDN U7164 ( .A(n4890), .B(ereg[45]), .Z(n5070) );
  NAND U7165 ( .A(n5072), .B(n5073), .Z(n3812) );
  NANDN U7166 ( .A(init), .B(e[46]), .Z(n5073) );
  AND U7167 ( .A(n5074), .B(n5075), .Z(n5072) );
  NAND U7168 ( .A(ereg[45]), .B(n4895), .Z(n5075) );
  NANDN U7169 ( .A(n4890), .B(ereg[46]), .Z(n5074) );
  NAND U7170 ( .A(n5076), .B(n5077), .Z(n3811) );
  NANDN U7171 ( .A(init), .B(e[47]), .Z(n5077) );
  AND U7172 ( .A(n5078), .B(n5079), .Z(n5076) );
  NAND U7173 ( .A(ereg[46]), .B(n4895), .Z(n5079) );
  NANDN U7174 ( .A(n4890), .B(ereg[47]), .Z(n5078) );
  NAND U7175 ( .A(n5080), .B(n5081), .Z(n3810) );
  NANDN U7176 ( .A(init), .B(e[48]), .Z(n5081) );
  AND U7177 ( .A(n5082), .B(n5083), .Z(n5080) );
  NAND U7178 ( .A(ereg[47]), .B(n4895), .Z(n5083) );
  NANDN U7179 ( .A(n4890), .B(ereg[48]), .Z(n5082) );
  NAND U7180 ( .A(n5084), .B(n5085), .Z(n3809) );
  NANDN U7181 ( .A(init), .B(e[49]), .Z(n5085) );
  AND U7182 ( .A(n5086), .B(n5087), .Z(n5084) );
  NAND U7183 ( .A(ereg[48]), .B(n4895), .Z(n5087) );
  NANDN U7184 ( .A(n4890), .B(ereg[49]), .Z(n5086) );
  NAND U7185 ( .A(n5088), .B(n5089), .Z(n3808) );
  NANDN U7186 ( .A(init), .B(e[50]), .Z(n5089) );
  AND U7187 ( .A(n5090), .B(n5091), .Z(n5088) );
  NAND U7188 ( .A(ereg[49]), .B(n4895), .Z(n5091) );
  NANDN U7189 ( .A(n4890), .B(ereg[50]), .Z(n5090) );
  NAND U7190 ( .A(n5092), .B(n5093), .Z(n3807) );
  NANDN U7191 ( .A(init), .B(e[51]), .Z(n5093) );
  AND U7192 ( .A(n5094), .B(n5095), .Z(n5092) );
  NAND U7193 ( .A(ereg[50]), .B(n4895), .Z(n5095) );
  NANDN U7194 ( .A(n4890), .B(ereg[51]), .Z(n5094) );
  NAND U7195 ( .A(n5096), .B(n5097), .Z(n3806) );
  NANDN U7196 ( .A(init), .B(e[52]), .Z(n5097) );
  AND U7197 ( .A(n5098), .B(n5099), .Z(n5096) );
  NAND U7198 ( .A(ereg[51]), .B(n4895), .Z(n5099) );
  NANDN U7199 ( .A(n4890), .B(ereg[52]), .Z(n5098) );
  NAND U7200 ( .A(n5100), .B(n5101), .Z(n3805) );
  NANDN U7201 ( .A(init), .B(e[53]), .Z(n5101) );
  AND U7202 ( .A(n5102), .B(n5103), .Z(n5100) );
  NAND U7203 ( .A(ereg[52]), .B(n4895), .Z(n5103) );
  NANDN U7204 ( .A(n4890), .B(ereg[53]), .Z(n5102) );
  NAND U7205 ( .A(n5104), .B(n5105), .Z(n3804) );
  NANDN U7206 ( .A(init), .B(e[54]), .Z(n5105) );
  AND U7207 ( .A(n5106), .B(n5107), .Z(n5104) );
  NAND U7208 ( .A(ereg[53]), .B(n4895), .Z(n5107) );
  NANDN U7209 ( .A(n4890), .B(ereg[54]), .Z(n5106) );
  NAND U7210 ( .A(n5108), .B(n5109), .Z(n3803) );
  NANDN U7211 ( .A(init), .B(e[55]), .Z(n5109) );
  AND U7212 ( .A(n5110), .B(n5111), .Z(n5108) );
  NAND U7213 ( .A(ereg[54]), .B(n4895), .Z(n5111) );
  NANDN U7214 ( .A(n4890), .B(ereg[55]), .Z(n5110) );
  NAND U7215 ( .A(n5112), .B(n5113), .Z(n3802) );
  NANDN U7216 ( .A(init), .B(e[56]), .Z(n5113) );
  AND U7217 ( .A(n5114), .B(n5115), .Z(n5112) );
  NAND U7218 ( .A(ereg[55]), .B(n4895), .Z(n5115) );
  NANDN U7219 ( .A(n4890), .B(ereg[56]), .Z(n5114) );
  NAND U7220 ( .A(n5116), .B(n5117), .Z(n3801) );
  NANDN U7221 ( .A(init), .B(e[57]), .Z(n5117) );
  AND U7222 ( .A(n5118), .B(n5119), .Z(n5116) );
  NAND U7223 ( .A(ereg[56]), .B(n4895), .Z(n5119) );
  NANDN U7224 ( .A(n4890), .B(ereg[57]), .Z(n5118) );
  NAND U7225 ( .A(n5120), .B(n5121), .Z(n3800) );
  NANDN U7226 ( .A(init), .B(e[58]), .Z(n5121) );
  AND U7227 ( .A(n5122), .B(n5123), .Z(n5120) );
  NAND U7228 ( .A(ereg[57]), .B(n4895), .Z(n5123) );
  NANDN U7229 ( .A(n4890), .B(ereg[58]), .Z(n5122) );
  NAND U7230 ( .A(n5124), .B(n5125), .Z(n3799) );
  NANDN U7231 ( .A(init), .B(e[59]), .Z(n5125) );
  AND U7232 ( .A(n5126), .B(n5127), .Z(n5124) );
  NAND U7233 ( .A(ereg[58]), .B(n4895), .Z(n5127) );
  NANDN U7234 ( .A(n4890), .B(ereg[59]), .Z(n5126) );
  NAND U7235 ( .A(n5128), .B(n5129), .Z(n3798) );
  NANDN U7236 ( .A(init), .B(e[60]), .Z(n5129) );
  AND U7237 ( .A(n5130), .B(n5131), .Z(n5128) );
  NAND U7238 ( .A(ereg[59]), .B(n4895), .Z(n5131) );
  NANDN U7239 ( .A(n4890), .B(ereg[60]), .Z(n5130) );
  NAND U7240 ( .A(n5132), .B(n5133), .Z(n3797) );
  NANDN U7241 ( .A(init), .B(e[61]), .Z(n5133) );
  AND U7242 ( .A(n5134), .B(n5135), .Z(n5132) );
  NAND U7243 ( .A(ereg[60]), .B(n4895), .Z(n5135) );
  NANDN U7244 ( .A(n4890), .B(ereg[61]), .Z(n5134) );
  NAND U7245 ( .A(n5136), .B(n5137), .Z(n3796) );
  NANDN U7246 ( .A(init), .B(e[62]), .Z(n5137) );
  AND U7247 ( .A(n5138), .B(n5139), .Z(n5136) );
  NAND U7248 ( .A(ereg[61]), .B(n4895), .Z(n5139) );
  NANDN U7249 ( .A(n4890), .B(ereg[62]), .Z(n5138) );
  NAND U7250 ( .A(n5140), .B(n5141), .Z(n3795) );
  NANDN U7251 ( .A(init), .B(e[63]), .Z(n5141) );
  AND U7252 ( .A(n5142), .B(n5143), .Z(n5140) );
  NAND U7253 ( .A(ereg[62]), .B(n4895), .Z(n5143) );
  NANDN U7254 ( .A(n4890), .B(ereg[63]), .Z(n5142) );
  NAND U7255 ( .A(n5144), .B(n5145), .Z(n3794) );
  NANDN U7256 ( .A(init), .B(e[64]), .Z(n5145) );
  AND U7257 ( .A(n5146), .B(n5147), .Z(n5144) );
  NAND U7258 ( .A(ereg[63]), .B(n4895), .Z(n5147) );
  NANDN U7259 ( .A(n4890), .B(ereg[64]), .Z(n5146) );
  NAND U7260 ( .A(n5148), .B(n5149), .Z(n3793) );
  NANDN U7261 ( .A(init), .B(e[65]), .Z(n5149) );
  AND U7262 ( .A(n5150), .B(n5151), .Z(n5148) );
  NAND U7263 ( .A(ereg[64]), .B(n4895), .Z(n5151) );
  NANDN U7264 ( .A(n4890), .B(ereg[65]), .Z(n5150) );
  NAND U7265 ( .A(n5152), .B(n5153), .Z(n3792) );
  NANDN U7266 ( .A(init), .B(e[66]), .Z(n5153) );
  AND U7267 ( .A(n5154), .B(n5155), .Z(n5152) );
  NAND U7268 ( .A(ereg[65]), .B(n4895), .Z(n5155) );
  NANDN U7269 ( .A(n4890), .B(ereg[66]), .Z(n5154) );
  NAND U7270 ( .A(n5156), .B(n5157), .Z(n3791) );
  NANDN U7271 ( .A(init), .B(e[67]), .Z(n5157) );
  AND U7272 ( .A(n5158), .B(n5159), .Z(n5156) );
  NAND U7273 ( .A(ereg[66]), .B(n4895), .Z(n5159) );
  NANDN U7274 ( .A(n4890), .B(ereg[67]), .Z(n5158) );
  NAND U7275 ( .A(n5160), .B(n5161), .Z(n3790) );
  NANDN U7276 ( .A(init), .B(e[68]), .Z(n5161) );
  AND U7277 ( .A(n5162), .B(n5163), .Z(n5160) );
  NAND U7278 ( .A(ereg[67]), .B(n4895), .Z(n5163) );
  NANDN U7279 ( .A(n4890), .B(ereg[68]), .Z(n5162) );
  NAND U7280 ( .A(n5164), .B(n5165), .Z(n3789) );
  NANDN U7281 ( .A(init), .B(e[69]), .Z(n5165) );
  AND U7282 ( .A(n5166), .B(n5167), .Z(n5164) );
  NAND U7283 ( .A(ereg[68]), .B(n4895), .Z(n5167) );
  NANDN U7284 ( .A(n4890), .B(ereg[69]), .Z(n5166) );
  NAND U7285 ( .A(n5168), .B(n5169), .Z(n3788) );
  NANDN U7286 ( .A(init), .B(e[70]), .Z(n5169) );
  AND U7287 ( .A(n5170), .B(n5171), .Z(n5168) );
  NAND U7288 ( .A(ereg[69]), .B(n4895), .Z(n5171) );
  NANDN U7289 ( .A(n4890), .B(ereg[70]), .Z(n5170) );
  NAND U7290 ( .A(n5172), .B(n5173), .Z(n3787) );
  NANDN U7291 ( .A(init), .B(e[71]), .Z(n5173) );
  AND U7292 ( .A(n5174), .B(n5175), .Z(n5172) );
  NAND U7293 ( .A(ereg[70]), .B(n4895), .Z(n5175) );
  NANDN U7294 ( .A(n4890), .B(ereg[71]), .Z(n5174) );
  NAND U7295 ( .A(n5176), .B(n5177), .Z(n3786) );
  NANDN U7296 ( .A(init), .B(e[72]), .Z(n5177) );
  AND U7297 ( .A(n5178), .B(n5179), .Z(n5176) );
  NAND U7298 ( .A(ereg[71]), .B(n4895), .Z(n5179) );
  NANDN U7299 ( .A(n4890), .B(ereg[72]), .Z(n5178) );
  NAND U7300 ( .A(n5180), .B(n5181), .Z(n3785) );
  NANDN U7301 ( .A(init), .B(e[73]), .Z(n5181) );
  AND U7302 ( .A(n5182), .B(n5183), .Z(n5180) );
  NAND U7303 ( .A(ereg[72]), .B(n4895), .Z(n5183) );
  NANDN U7304 ( .A(n4890), .B(ereg[73]), .Z(n5182) );
  NAND U7305 ( .A(n5184), .B(n5185), .Z(n3784) );
  NANDN U7306 ( .A(init), .B(e[74]), .Z(n5185) );
  AND U7307 ( .A(n5186), .B(n5187), .Z(n5184) );
  NAND U7308 ( .A(ereg[73]), .B(n4895), .Z(n5187) );
  NANDN U7309 ( .A(n4890), .B(ereg[74]), .Z(n5186) );
  NAND U7310 ( .A(n5188), .B(n5189), .Z(n3783) );
  NANDN U7311 ( .A(init), .B(e[75]), .Z(n5189) );
  AND U7312 ( .A(n5190), .B(n5191), .Z(n5188) );
  NAND U7313 ( .A(ereg[74]), .B(n4895), .Z(n5191) );
  NANDN U7314 ( .A(n4890), .B(ereg[75]), .Z(n5190) );
  NAND U7315 ( .A(n5192), .B(n5193), .Z(n3782) );
  NANDN U7316 ( .A(init), .B(e[76]), .Z(n5193) );
  AND U7317 ( .A(n5194), .B(n5195), .Z(n5192) );
  NAND U7318 ( .A(ereg[75]), .B(n4895), .Z(n5195) );
  NANDN U7319 ( .A(n4890), .B(ereg[76]), .Z(n5194) );
  NAND U7320 ( .A(n5196), .B(n5197), .Z(n3781) );
  NANDN U7321 ( .A(init), .B(e[77]), .Z(n5197) );
  AND U7322 ( .A(n5198), .B(n5199), .Z(n5196) );
  NAND U7323 ( .A(ereg[76]), .B(n4895), .Z(n5199) );
  NANDN U7324 ( .A(n4890), .B(ereg[77]), .Z(n5198) );
  NAND U7325 ( .A(n5200), .B(n5201), .Z(n3780) );
  NANDN U7326 ( .A(init), .B(e[78]), .Z(n5201) );
  AND U7327 ( .A(n5202), .B(n5203), .Z(n5200) );
  NAND U7328 ( .A(ereg[77]), .B(n4895), .Z(n5203) );
  NANDN U7329 ( .A(n4890), .B(ereg[78]), .Z(n5202) );
  NAND U7330 ( .A(n5204), .B(n5205), .Z(n3779) );
  NANDN U7331 ( .A(init), .B(e[79]), .Z(n5205) );
  AND U7332 ( .A(n5206), .B(n5207), .Z(n5204) );
  NAND U7333 ( .A(ereg[78]), .B(n4895), .Z(n5207) );
  NANDN U7334 ( .A(n4890), .B(ereg[79]), .Z(n5206) );
  NAND U7335 ( .A(n5208), .B(n5209), .Z(n3778) );
  NANDN U7336 ( .A(init), .B(e[80]), .Z(n5209) );
  AND U7337 ( .A(n5210), .B(n5211), .Z(n5208) );
  NAND U7338 ( .A(ereg[79]), .B(n4895), .Z(n5211) );
  NANDN U7339 ( .A(n4890), .B(ereg[80]), .Z(n5210) );
  NAND U7340 ( .A(n5212), .B(n5213), .Z(n3777) );
  NANDN U7341 ( .A(init), .B(e[81]), .Z(n5213) );
  AND U7342 ( .A(n5214), .B(n5215), .Z(n5212) );
  NAND U7343 ( .A(ereg[80]), .B(n4895), .Z(n5215) );
  NANDN U7344 ( .A(n4890), .B(ereg[81]), .Z(n5214) );
  NAND U7345 ( .A(n5216), .B(n5217), .Z(n3776) );
  NANDN U7346 ( .A(init), .B(e[82]), .Z(n5217) );
  AND U7347 ( .A(n5218), .B(n5219), .Z(n5216) );
  NAND U7348 ( .A(ereg[81]), .B(n4895), .Z(n5219) );
  NANDN U7349 ( .A(n4890), .B(ereg[82]), .Z(n5218) );
  NAND U7350 ( .A(n5220), .B(n5221), .Z(n3775) );
  NANDN U7351 ( .A(init), .B(e[83]), .Z(n5221) );
  AND U7352 ( .A(n5222), .B(n5223), .Z(n5220) );
  NAND U7353 ( .A(ereg[82]), .B(n4895), .Z(n5223) );
  NANDN U7354 ( .A(n4890), .B(ereg[83]), .Z(n5222) );
  NAND U7355 ( .A(n5224), .B(n5225), .Z(n3774) );
  NANDN U7356 ( .A(init), .B(e[84]), .Z(n5225) );
  AND U7357 ( .A(n5226), .B(n5227), .Z(n5224) );
  NAND U7358 ( .A(ereg[83]), .B(n4895), .Z(n5227) );
  NANDN U7359 ( .A(n4890), .B(ereg[84]), .Z(n5226) );
  NAND U7360 ( .A(n5228), .B(n5229), .Z(n3773) );
  NANDN U7361 ( .A(init), .B(e[85]), .Z(n5229) );
  AND U7362 ( .A(n5230), .B(n5231), .Z(n5228) );
  NAND U7363 ( .A(ereg[84]), .B(n4895), .Z(n5231) );
  NANDN U7364 ( .A(n4890), .B(ereg[85]), .Z(n5230) );
  NAND U7365 ( .A(n5232), .B(n5233), .Z(n3772) );
  NANDN U7366 ( .A(init), .B(e[86]), .Z(n5233) );
  AND U7367 ( .A(n5234), .B(n5235), .Z(n5232) );
  NAND U7368 ( .A(ereg[85]), .B(n4895), .Z(n5235) );
  NANDN U7369 ( .A(n4890), .B(ereg[86]), .Z(n5234) );
  NAND U7370 ( .A(n5236), .B(n5237), .Z(n3771) );
  NANDN U7371 ( .A(init), .B(e[87]), .Z(n5237) );
  AND U7372 ( .A(n5238), .B(n5239), .Z(n5236) );
  NAND U7373 ( .A(ereg[86]), .B(n4895), .Z(n5239) );
  NANDN U7374 ( .A(n4890), .B(ereg[87]), .Z(n5238) );
  NAND U7375 ( .A(n5240), .B(n5241), .Z(n3770) );
  NANDN U7376 ( .A(init), .B(e[88]), .Z(n5241) );
  AND U7377 ( .A(n5242), .B(n5243), .Z(n5240) );
  NAND U7378 ( .A(ereg[87]), .B(n4895), .Z(n5243) );
  NANDN U7379 ( .A(n4890), .B(ereg[88]), .Z(n5242) );
  NAND U7380 ( .A(n5244), .B(n5245), .Z(n3769) );
  NANDN U7381 ( .A(init), .B(e[89]), .Z(n5245) );
  AND U7382 ( .A(n5246), .B(n5247), .Z(n5244) );
  NAND U7383 ( .A(ereg[88]), .B(n4895), .Z(n5247) );
  NANDN U7384 ( .A(n4890), .B(ereg[89]), .Z(n5246) );
  NAND U7385 ( .A(n5248), .B(n5249), .Z(n3768) );
  NANDN U7386 ( .A(init), .B(e[90]), .Z(n5249) );
  AND U7387 ( .A(n5250), .B(n5251), .Z(n5248) );
  NAND U7388 ( .A(ereg[89]), .B(n4895), .Z(n5251) );
  NANDN U7389 ( .A(n4890), .B(ereg[90]), .Z(n5250) );
  NAND U7390 ( .A(n5252), .B(n5253), .Z(n3767) );
  NANDN U7391 ( .A(init), .B(e[91]), .Z(n5253) );
  AND U7392 ( .A(n5254), .B(n5255), .Z(n5252) );
  NAND U7393 ( .A(ereg[90]), .B(n4895), .Z(n5255) );
  NANDN U7394 ( .A(n4890), .B(ereg[91]), .Z(n5254) );
  NAND U7395 ( .A(n5256), .B(n5257), .Z(n3766) );
  NANDN U7396 ( .A(init), .B(e[92]), .Z(n5257) );
  AND U7397 ( .A(n5258), .B(n5259), .Z(n5256) );
  NAND U7398 ( .A(ereg[91]), .B(n4895), .Z(n5259) );
  NANDN U7399 ( .A(n4890), .B(ereg[92]), .Z(n5258) );
  NAND U7400 ( .A(n5260), .B(n5261), .Z(n3765) );
  NANDN U7401 ( .A(init), .B(e[93]), .Z(n5261) );
  AND U7402 ( .A(n5262), .B(n5263), .Z(n5260) );
  NAND U7403 ( .A(ereg[92]), .B(n4895), .Z(n5263) );
  NANDN U7404 ( .A(n4890), .B(ereg[93]), .Z(n5262) );
  NAND U7405 ( .A(n5264), .B(n5265), .Z(n3764) );
  NANDN U7406 ( .A(init), .B(e[94]), .Z(n5265) );
  AND U7407 ( .A(n5266), .B(n5267), .Z(n5264) );
  NAND U7408 ( .A(ereg[93]), .B(n4895), .Z(n5267) );
  NANDN U7409 ( .A(n4890), .B(ereg[94]), .Z(n5266) );
  NAND U7410 ( .A(n5268), .B(n5269), .Z(n3763) );
  NANDN U7411 ( .A(init), .B(e[95]), .Z(n5269) );
  AND U7412 ( .A(n5270), .B(n5271), .Z(n5268) );
  NAND U7413 ( .A(ereg[94]), .B(n4895), .Z(n5271) );
  NANDN U7414 ( .A(n4890), .B(ereg[95]), .Z(n5270) );
  NAND U7415 ( .A(n5272), .B(n5273), .Z(n3762) );
  NANDN U7416 ( .A(init), .B(e[96]), .Z(n5273) );
  AND U7417 ( .A(n5274), .B(n5275), .Z(n5272) );
  NAND U7418 ( .A(ereg[95]), .B(n4895), .Z(n5275) );
  NANDN U7419 ( .A(n4890), .B(ereg[96]), .Z(n5274) );
  NAND U7420 ( .A(n5276), .B(n5277), .Z(n3761) );
  NANDN U7421 ( .A(init), .B(e[97]), .Z(n5277) );
  AND U7422 ( .A(n5278), .B(n5279), .Z(n5276) );
  NAND U7423 ( .A(ereg[96]), .B(n4895), .Z(n5279) );
  NANDN U7424 ( .A(n4890), .B(ereg[97]), .Z(n5278) );
  NAND U7425 ( .A(n5280), .B(n5281), .Z(n3760) );
  NANDN U7426 ( .A(init), .B(e[98]), .Z(n5281) );
  AND U7427 ( .A(n5282), .B(n5283), .Z(n5280) );
  NAND U7428 ( .A(ereg[97]), .B(n4895), .Z(n5283) );
  NANDN U7429 ( .A(n4890), .B(ereg[98]), .Z(n5282) );
  NAND U7430 ( .A(n5284), .B(n5285), .Z(n3759) );
  NANDN U7431 ( .A(init), .B(e[99]), .Z(n5285) );
  AND U7432 ( .A(n5286), .B(n5287), .Z(n5284) );
  NAND U7433 ( .A(ereg[98]), .B(n4895), .Z(n5287) );
  NANDN U7434 ( .A(n4890), .B(ereg[99]), .Z(n5286) );
  NAND U7435 ( .A(n5288), .B(n5289), .Z(n3758) );
  NANDN U7436 ( .A(init), .B(e[100]), .Z(n5289) );
  AND U7437 ( .A(n5290), .B(n5291), .Z(n5288) );
  NAND U7438 ( .A(ereg[99]), .B(n4895), .Z(n5291) );
  NANDN U7439 ( .A(n4890), .B(ereg[100]), .Z(n5290) );
  NAND U7440 ( .A(n5292), .B(n5293), .Z(n3757) );
  NANDN U7441 ( .A(init), .B(e[101]), .Z(n5293) );
  AND U7442 ( .A(n5294), .B(n5295), .Z(n5292) );
  NAND U7443 ( .A(ereg[100]), .B(n4895), .Z(n5295) );
  NANDN U7444 ( .A(n4890), .B(ereg[101]), .Z(n5294) );
  NAND U7445 ( .A(n5296), .B(n5297), .Z(n3756) );
  NANDN U7446 ( .A(init), .B(e[102]), .Z(n5297) );
  AND U7447 ( .A(n5298), .B(n5299), .Z(n5296) );
  NAND U7448 ( .A(ereg[101]), .B(n4895), .Z(n5299) );
  NANDN U7449 ( .A(n4890), .B(ereg[102]), .Z(n5298) );
  NAND U7450 ( .A(n5300), .B(n5301), .Z(n3755) );
  NANDN U7451 ( .A(init), .B(e[103]), .Z(n5301) );
  AND U7452 ( .A(n5302), .B(n5303), .Z(n5300) );
  NAND U7453 ( .A(ereg[102]), .B(n4895), .Z(n5303) );
  NANDN U7454 ( .A(n4890), .B(ereg[103]), .Z(n5302) );
  NAND U7455 ( .A(n5304), .B(n5305), .Z(n3754) );
  NANDN U7456 ( .A(init), .B(e[104]), .Z(n5305) );
  AND U7457 ( .A(n5306), .B(n5307), .Z(n5304) );
  NAND U7458 ( .A(ereg[103]), .B(n4895), .Z(n5307) );
  NANDN U7459 ( .A(n4890), .B(ereg[104]), .Z(n5306) );
  NAND U7460 ( .A(n5308), .B(n5309), .Z(n3753) );
  NANDN U7461 ( .A(init), .B(e[105]), .Z(n5309) );
  AND U7462 ( .A(n5310), .B(n5311), .Z(n5308) );
  NAND U7463 ( .A(ereg[104]), .B(n4895), .Z(n5311) );
  NANDN U7464 ( .A(n4890), .B(ereg[105]), .Z(n5310) );
  NAND U7465 ( .A(n5312), .B(n5313), .Z(n3752) );
  NANDN U7466 ( .A(init), .B(e[106]), .Z(n5313) );
  AND U7467 ( .A(n5314), .B(n5315), .Z(n5312) );
  NAND U7468 ( .A(ereg[105]), .B(n4895), .Z(n5315) );
  NANDN U7469 ( .A(n4890), .B(ereg[106]), .Z(n5314) );
  NAND U7470 ( .A(n5316), .B(n5317), .Z(n3751) );
  NANDN U7471 ( .A(init), .B(e[107]), .Z(n5317) );
  AND U7472 ( .A(n5318), .B(n5319), .Z(n5316) );
  NAND U7473 ( .A(ereg[106]), .B(n4895), .Z(n5319) );
  NANDN U7474 ( .A(n4890), .B(ereg[107]), .Z(n5318) );
  NAND U7475 ( .A(n5320), .B(n5321), .Z(n3750) );
  NANDN U7476 ( .A(init), .B(e[108]), .Z(n5321) );
  AND U7477 ( .A(n5322), .B(n5323), .Z(n5320) );
  NAND U7478 ( .A(ereg[107]), .B(n4895), .Z(n5323) );
  NANDN U7479 ( .A(n4890), .B(ereg[108]), .Z(n5322) );
  NAND U7480 ( .A(n5324), .B(n5325), .Z(n3749) );
  NANDN U7481 ( .A(init), .B(e[109]), .Z(n5325) );
  AND U7482 ( .A(n5326), .B(n5327), .Z(n5324) );
  NAND U7483 ( .A(ereg[108]), .B(n4895), .Z(n5327) );
  NANDN U7484 ( .A(n4890), .B(ereg[109]), .Z(n5326) );
  NAND U7485 ( .A(n5328), .B(n5329), .Z(n3748) );
  NANDN U7486 ( .A(init), .B(e[110]), .Z(n5329) );
  AND U7487 ( .A(n5330), .B(n5331), .Z(n5328) );
  NAND U7488 ( .A(ereg[109]), .B(n4895), .Z(n5331) );
  NANDN U7489 ( .A(n4890), .B(ereg[110]), .Z(n5330) );
  NAND U7490 ( .A(n5332), .B(n5333), .Z(n3747) );
  NANDN U7491 ( .A(init), .B(e[111]), .Z(n5333) );
  AND U7492 ( .A(n5334), .B(n5335), .Z(n5332) );
  NAND U7493 ( .A(ereg[110]), .B(n4895), .Z(n5335) );
  NANDN U7494 ( .A(n4890), .B(ereg[111]), .Z(n5334) );
  NAND U7495 ( .A(n5336), .B(n5337), .Z(n3746) );
  NANDN U7496 ( .A(init), .B(e[112]), .Z(n5337) );
  AND U7497 ( .A(n5338), .B(n5339), .Z(n5336) );
  NAND U7498 ( .A(ereg[111]), .B(n4895), .Z(n5339) );
  NANDN U7499 ( .A(n4890), .B(ereg[112]), .Z(n5338) );
  NAND U7500 ( .A(n5340), .B(n5341), .Z(n3745) );
  NANDN U7501 ( .A(init), .B(e[113]), .Z(n5341) );
  AND U7502 ( .A(n5342), .B(n5343), .Z(n5340) );
  NAND U7503 ( .A(ereg[112]), .B(n4895), .Z(n5343) );
  NANDN U7504 ( .A(n4890), .B(ereg[113]), .Z(n5342) );
  NAND U7505 ( .A(n5344), .B(n5345), .Z(n3744) );
  NANDN U7506 ( .A(init), .B(e[114]), .Z(n5345) );
  AND U7507 ( .A(n5346), .B(n5347), .Z(n5344) );
  NAND U7508 ( .A(ereg[113]), .B(n4895), .Z(n5347) );
  NANDN U7509 ( .A(n4890), .B(ereg[114]), .Z(n5346) );
  NAND U7510 ( .A(n5348), .B(n5349), .Z(n3743) );
  NANDN U7511 ( .A(init), .B(e[115]), .Z(n5349) );
  AND U7512 ( .A(n5350), .B(n5351), .Z(n5348) );
  NAND U7513 ( .A(ereg[114]), .B(n4895), .Z(n5351) );
  NANDN U7514 ( .A(n4890), .B(ereg[115]), .Z(n5350) );
  NAND U7515 ( .A(n5352), .B(n5353), .Z(n3742) );
  NANDN U7516 ( .A(init), .B(e[116]), .Z(n5353) );
  AND U7517 ( .A(n5354), .B(n5355), .Z(n5352) );
  NAND U7518 ( .A(ereg[115]), .B(n4895), .Z(n5355) );
  NANDN U7519 ( .A(n4890), .B(ereg[116]), .Z(n5354) );
  NAND U7520 ( .A(n5356), .B(n5357), .Z(n3741) );
  NANDN U7521 ( .A(init), .B(e[117]), .Z(n5357) );
  AND U7522 ( .A(n5358), .B(n5359), .Z(n5356) );
  NAND U7523 ( .A(ereg[116]), .B(n4895), .Z(n5359) );
  NANDN U7524 ( .A(n4890), .B(ereg[117]), .Z(n5358) );
  NAND U7525 ( .A(n5360), .B(n5361), .Z(n3740) );
  NANDN U7526 ( .A(init), .B(e[118]), .Z(n5361) );
  AND U7527 ( .A(n5362), .B(n5363), .Z(n5360) );
  NAND U7528 ( .A(ereg[117]), .B(n4895), .Z(n5363) );
  NANDN U7529 ( .A(n4890), .B(ereg[118]), .Z(n5362) );
  NAND U7530 ( .A(n5364), .B(n5365), .Z(n3739) );
  NANDN U7531 ( .A(init), .B(e[119]), .Z(n5365) );
  AND U7532 ( .A(n5366), .B(n5367), .Z(n5364) );
  NAND U7533 ( .A(ereg[118]), .B(n4895), .Z(n5367) );
  NANDN U7534 ( .A(n4890), .B(ereg[119]), .Z(n5366) );
  NAND U7535 ( .A(n5368), .B(n5369), .Z(n3738) );
  NANDN U7536 ( .A(init), .B(e[120]), .Z(n5369) );
  AND U7537 ( .A(n5370), .B(n5371), .Z(n5368) );
  NAND U7538 ( .A(ereg[119]), .B(n4895), .Z(n5371) );
  NANDN U7539 ( .A(n4890), .B(ereg[120]), .Z(n5370) );
  NAND U7540 ( .A(n5372), .B(n5373), .Z(n3737) );
  NANDN U7541 ( .A(init), .B(e[121]), .Z(n5373) );
  AND U7542 ( .A(n5374), .B(n5375), .Z(n5372) );
  NAND U7543 ( .A(ereg[120]), .B(n4895), .Z(n5375) );
  NANDN U7544 ( .A(n4890), .B(ereg[121]), .Z(n5374) );
  NAND U7545 ( .A(n5376), .B(n5377), .Z(n3736) );
  NANDN U7546 ( .A(init), .B(e[122]), .Z(n5377) );
  AND U7547 ( .A(n5378), .B(n5379), .Z(n5376) );
  NAND U7548 ( .A(ereg[121]), .B(n4895), .Z(n5379) );
  NANDN U7549 ( .A(n4890), .B(ereg[122]), .Z(n5378) );
  NAND U7550 ( .A(n5380), .B(n5381), .Z(n3735) );
  NANDN U7551 ( .A(init), .B(e[123]), .Z(n5381) );
  AND U7552 ( .A(n5382), .B(n5383), .Z(n5380) );
  NAND U7553 ( .A(ereg[122]), .B(n4895), .Z(n5383) );
  NANDN U7554 ( .A(n4890), .B(ereg[123]), .Z(n5382) );
  NAND U7555 ( .A(n5384), .B(n5385), .Z(n3734) );
  NANDN U7556 ( .A(init), .B(e[124]), .Z(n5385) );
  AND U7557 ( .A(n5386), .B(n5387), .Z(n5384) );
  NAND U7558 ( .A(ereg[123]), .B(n4895), .Z(n5387) );
  NANDN U7559 ( .A(n4890), .B(ereg[124]), .Z(n5386) );
  NAND U7560 ( .A(n5388), .B(n5389), .Z(n3733) );
  NANDN U7561 ( .A(init), .B(e[125]), .Z(n5389) );
  AND U7562 ( .A(n5390), .B(n5391), .Z(n5388) );
  NAND U7563 ( .A(ereg[124]), .B(n4895), .Z(n5391) );
  NANDN U7564 ( .A(n4890), .B(ereg[125]), .Z(n5390) );
  NAND U7565 ( .A(n5392), .B(n5393), .Z(n3732) );
  NANDN U7566 ( .A(init), .B(e[126]), .Z(n5393) );
  AND U7567 ( .A(n5394), .B(n5395), .Z(n5392) );
  NAND U7568 ( .A(ereg[125]), .B(n4895), .Z(n5395) );
  NANDN U7569 ( .A(n4890), .B(ereg[126]), .Z(n5394) );
  NAND U7570 ( .A(n5396), .B(n5397), .Z(n3731) );
  NANDN U7571 ( .A(init), .B(e[127]), .Z(n5397) );
  AND U7572 ( .A(n5398), .B(n5399), .Z(n5396) );
  NAND U7573 ( .A(ereg[126]), .B(n4895), .Z(n5399) );
  NANDN U7574 ( .A(n4890), .B(ereg[127]), .Z(n5398) );
  NAND U7575 ( .A(n5400), .B(n5401), .Z(n3730) );
  NANDN U7576 ( .A(init), .B(e[128]), .Z(n5401) );
  AND U7577 ( .A(n5402), .B(n5403), .Z(n5400) );
  NAND U7578 ( .A(ereg[127]), .B(n4895), .Z(n5403) );
  NANDN U7579 ( .A(n4890), .B(ereg[128]), .Z(n5402) );
  NAND U7580 ( .A(n5404), .B(n5405), .Z(n3729) );
  NANDN U7581 ( .A(init), .B(e[129]), .Z(n5405) );
  AND U7582 ( .A(n5406), .B(n5407), .Z(n5404) );
  NAND U7583 ( .A(ereg[128]), .B(n4895), .Z(n5407) );
  NANDN U7584 ( .A(n4890), .B(ereg[129]), .Z(n5406) );
  NAND U7585 ( .A(n5408), .B(n5409), .Z(n3728) );
  NANDN U7586 ( .A(init), .B(e[130]), .Z(n5409) );
  AND U7587 ( .A(n5410), .B(n5411), .Z(n5408) );
  NAND U7588 ( .A(ereg[129]), .B(n4895), .Z(n5411) );
  NANDN U7589 ( .A(n4890), .B(ereg[130]), .Z(n5410) );
  NAND U7590 ( .A(n5412), .B(n5413), .Z(n3727) );
  NANDN U7591 ( .A(init), .B(e[131]), .Z(n5413) );
  AND U7592 ( .A(n5414), .B(n5415), .Z(n5412) );
  NAND U7593 ( .A(ereg[130]), .B(n4895), .Z(n5415) );
  NANDN U7594 ( .A(n4890), .B(ereg[131]), .Z(n5414) );
  NAND U7595 ( .A(n5416), .B(n5417), .Z(n3726) );
  NANDN U7596 ( .A(init), .B(e[132]), .Z(n5417) );
  AND U7597 ( .A(n5418), .B(n5419), .Z(n5416) );
  NAND U7598 ( .A(ereg[131]), .B(n4895), .Z(n5419) );
  NANDN U7599 ( .A(n4890), .B(ereg[132]), .Z(n5418) );
  NAND U7600 ( .A(n5420), .B(n5421), .Z(n3725) );
  NANDN U7601 ( .A(init), .B(e[133]), .Z(n5421) );
  AND U7602 ( .A(n5422), .B(n5423), .Z(n5420) );
  NAND U7603 ( .A(ereg[132]), .B(n4895), .Z(n5423) );
  NANDN U7604 ( .A(n4890), .B(ereg[133]), .Z(n5422) );
  NAND U7605 ( .A(n5424), .B(n5425), .Z(n3724) );
  NANDN U7606 ( .A(init), .B(e[134]), .Z(n5425) );
  AND U7607 ( .A(n5426), .B(n5427), .Z(n5424) );
  NAND U7608 ( .A(ereg[133]), .B(n4895), .Z(n5427) );
  NANDN U7609 ( .A(n4890), .B(ereg[134]), .Z(n5426) );
  NAND U7610 ( .A(n5428), .B(n5429), .Z(n3723) );
  NANDN U7611 ( .A(init), .B(e[135]), .Z(n5429) );
  AND U7612 ( .A(n5430), .B(n5431), .Z(n5428) );
  NAND U7613 ( .A(ereg[134]), .B(n4895), .Z(n5431) );
  NANDN U7614 ( .A(n4890), .B(ereg[135]), .Z(n5430) );
  NAND U7615 ( .A(n5432), .B(n5433), .Z(n3722) );
  NANDN U7616 ( .A(init), .B(e[136]), .Z(n5433) );
  AND U7617 ( .A(n5434), .B(n5435), .Z(n5432) );
  NAND U7618 ( .A(ereg[135]), .B(n4895), .Z(n5435) );
  NANDN U7619 ( .A(n4890), .B(ereg[136]), .Z(n5434) );
  NAND U7620 ( .A(n5436), .B(n5437), .Z(n3721) );
  NANDN U7621 ( .A(init), .B(e[137]), .Z(n5437) );
  AND U7622 ( .A(n5438), .B(n5439), .Z(n5436) );
  NAND U7623 ( .A(ereg[136]), .B(n4895), .Z(n5439) );
  NANDN U7624 ( .A(n4890), .B(ereg[137]), .Z(n5438) );
  NAND U7625 ( .A(n5440), .B(n5441), .Z(n3720) );
  NANDN U7626 ( .A(init), .B(e[138]), .Z(n5441) );
  AND U7627 ( .A(n5442), .B(n5443), .Z(n5440) );
  NAND U7628 ( .A(ereg[137]), .B(n4895), .Z(n5443) );
  NANDN U7629 ( .A(n4890), .B(ereg[138]), .Z(n5442) );
  NAND U7630 ( .A(n5444), .B(n5445), .Z(n3719) );
  NANDN U7631 ( .A(init), .B(e[139]), .Z(n5445) );
  AND U7632 ( .A(n5446), .B(n5447), .Z(n5444) );
  NAND U7633 ( .A(ereg[138]), .B(n4895), .Z(n5447) );
  NANDN U7634 ( .A(n4890), .B(ereg[139]), .Z(n5446) );
  NAND U7635 ( .A(n5448), .B(n5449), .Z(n3718) );
  NANDN U7636 ( .A(init), .B(e[140]), .Z(n5449) );
  AND U7637 ( .A(n5450), .B(n5451), .Z(n5448) );
  NAND U7638 ( .A(ereg[139]), .B(n4895), .Z(n5451) );
  NANDN U7639 ( .A(n4890), .B(ereg[140]), .Z(n5450) );
  NAND U7640 ( .A(n5452), .B(n5453), .Z(n3717) );
  NANDN U7641 ( .A(init), .B(e[141]), .Z(n5453) );
  AND U7642 ( .A(n5454), .B(n5455), .Z(n5452) );
  NAND U7643 ( .A(ereg[140]), .B(n4895), .Z(n5455) );
  NANDN U7644 ( .A(n4890), .B(ereg[141]), .Z(n5454) );
  NAND U7645 ( .A(n5456), .B(n5457), .Z(n3716) );
  NANDN U7646 ( .A(init), .B(e[142]), .Z(n5457) );
  AND U7647 ( .A(n5458), .B(n5459), .Z(n5456) );
  NAND U7648 ( .A(ereg[141]), .B(n4895), .Z(n5459) );
  NANDN U7649 ( .A(n4890), .B(ereg[142]), .Z(n5458) );
  NAND U7650 ( .A(n5460), .B(n5461), .Z(n3715) );
  NANDN U7651 ( .A(init), .B(e[143]), .Z(n5461) );
  AND U7652 ( .A(n5462), .B(n5463), .Z(n5460) );
  NAND U7653 ( .A(ereg[142]), .B(n4895), .Z(n5463) );
  NANDN U7654 ( .A(n4890), .B(ereg[143]), .Z(n5462) );
  NAND U7655 ( .A(n5464), .B(n5465), .Z(n3714) );
  NANDN U7656 ( .A(init), .B(e[144]), .Z(n5465) );
  AND U7657 ( .A(n5466), .B(n5467), .Z(n5464) );
  NAND U7658 ( .A(ereg[143]), .B(n4895), .Z(n5467) );
  NANDN U7659 ( .A(n4890), .B(ereg[144]), .Z(n5466) );
  NAND U7660 ( .A(n5468), .B(n5469), .Z(n3713) );
  NANDN U7661 ( .A(init), .B(e[145]), .Z(n5469) );
  AND U7662 ( .A(n5470), .B(n5471), .Z(n5468) );
  NAND U7663 ( .A(ereg[144]), .B(n4895), .Z(n5471) );
  NANDN U7664 ( .A(n4890), .B(ereg[145]), .Z(n5470) );
  NAND U7665 ( .A(n5472), .B(n5473), .Z(n3712) );
  NANDN U7666 ( .A(init), .B(e[146]), .Z(n5473) );
  AND U7667 ( .A(n5474), .B(n5475), .Z(n5472) );
  NAND U7668 ( .A(ereg[145]), .B(n4895), .Z(n5475) );
  NANDN U7669 ( .A(n4890), .B(ereg[146]), .Z(n5474) );
  NAND U7670 ( .A(n5476), .B(n5477), .Z(n3711) );
  NANDN U7671 ( .A(init), .B(e[147]), .Z(n5477) );
  AND U7672 ( .A(n5478), .B(n5479), .Z(n5476) );
  NAND U7673 ( .A(ereg[146]), .B(n4895), .Z(n5479) );
  NANDN U7674 ( .A(n4890), .B(ereg[147]), .Z(n5478) );
  NAND U7675 ( .A(n5480), .B(n5481), .Z(n3710) );
  NANDN U7676 ( .A(init), .B(e[148]), .Z(n5481) );
  AND U7677 ( .A(n5482), .B(n5483), .Z(n5480) );
  NAND U7678 ( .A(ereg[147]), .B(n4895), .Z(n5483) );
  NANDN U7679 ( .A(n4890), .B(ereg[148]), .Z(n5482) );
  NAND U7680 ( .A(n5484), .B(n5485), .Z(n3709) );
  NANDN U7681 ( .A(init), .B(e[149]), .Z(n5485) );
  AND U7682 ( .A(n5486), .B(n5487), .Z(n5484) );
  NAND U7683 ( .A(ereg[148]), .B(n4895), .Z(n5487) );
  NANDN U7684 ( .A(n4890), .B(ereg[149]), .Z(n5486) );
  NAND U7685 ( .A(n5488), .B(n5489), .Z(n3708) );
  NANDN U7686 ( .A(init), .B(e[150]), .Z(n5489) );
  AND U7687 ( .A(n5490), .B(n5491), .Z(n5488) );
  NAND U7688 ( .A(ereg[149]), .B(n4895), .Z(n5491) );
  NANDN U7689 ( .A(n4890), .B(ereg[150]), .Z(n5490) );
  NAND U7690 ( .A(n5492), .B(n5493), .Z(n3707) );
  NANDN U7691 ( .A(init), .B(e[151]), .Z(n5493) );
  AND U7692 ( .A(n5494), .B(n5495), .Z(n5492) );
  NAND U7693 ( .A(ereg[150]), .B(n4895), .Z(n5495) );
  NANDN U7694 ( .A(n4890), .B(ereg[151]), .Z(n5494) );
  NAND U7695 ( .A(n5496), .B(n5497), .Z(n3706) );
  NANDN U7696 ( .A(init), .B(e[152]), .Z(n5497) );
  AND U7697 ( .A(n5498), .B(n5499), .Z(n5496) );
  NAND U7698 ( .A(ereg[151]), .B(n4895), .Z(n5499) );
  NANDN U7699 ( .A(n4890), .B(ereg[152]), .Z(n5498) );
  NAND U7700 ( .A(n5500), .B(n5501), .Z(n3705) );
  NANDN U7701 ( .A(init), .B(e[153]), .Z(n5501) );
  AND U7702 ( .A(n5502), .B(n5503), .Z(n5500) );
  NAND U7703 ( .A(ereg[152]), .B(n4895), .Z(n5503) );
  NANDN U7704 ( .A(n4890), .B(ereg[153]), .Z(n5502) );
  NAND U7705 ( .A(n5504), .B(n5505), .Z(n3704) );
  NANDN U7706 ( .A(init), .B(e[154]), .Z(n5505) );
  AND U7707 ( .A(n5506), .B(n5507), .Z(n5504) );
  NAND U7708 ( .A(ereg[153]), .B(n4895), .Z(n5507) );
  NANDN U7709 ( .A(n4890), .B(ereg[154]), .Z(n5506) );
  NAND U7710 ( .A(n5508), .B(n5509), .Z(n3703) );
  NANDN U7711 ( .A(init), .B(e[155]), .Z(n5509) );
  AND U7712 ( .A(n5510), .B(n5511), .Z(n5508) );
  NAND U7713 ( .A(ereg[154]), .B(n4895), .Z(n5511) );
  NANDN U7714 ( .A(n4890), .B(ereg[155]), .Z(n5510) );
  NAND U7715 ( .A(n5512), .B(n5513), .Z(n3702) );
  NANDN U7716 ( .A(init), .B(e[156]), .Z(n5513) );
  AND U7717 ( .A(n5514), .B(n5515), .Z(n5512) );
  NAND U7718 ( .A(ereg[155]), .B(n4895), .Z(n5515) );
  NANDN U7719 ( .A(n4890), .B(ereg[156]), .Z(n5514) );
  NAND U7720 ( .A(n5516), .B(n5517), .Z(n3701) );
  NANDN U7721 ( .A(init), .B(e[157]), .Z(n5517) );
  AND U7722 ( .A(n5518), .B(n5519), .Z(n5516) );
  NAND U7723 ( .A(ereg[156]), .B(n4895), .Z(n5519) );
  NANDN U7724 ( .A(n4890), .B(ereg[157]), .Z(n5518) );
  NAND U7725 ( .A(n5520), .B(n5521), .Z(n3700) );
  NANDN U7726 ( .A(init), .B(e[158]), .Z(n5521) );
  AND U7727 ( .A(n5522), .B(n5523), .Z(n5520) );
  NAND U7728 ( .A(ereg[157]), .B(n4895), .Z(n5523) );
  NANDN U7729 ( .A(n4890), .B(ereg[158]), .Z(n5522) );
  NAND U7730 ( .A(n5524), .B(n5525), .Z(n3699) );
  NANDN U7731 ( .A(init), .B(e[159]), .Z(n5525) );
  AND U7732 ( .A(n5526), .B(n5527), .Z(n5524) );
  NAND U7733 ( .A(ereg[158]), .B(n4895), .Z(n5527) );
  NANDN U7734 ( .A(n4890), .B(ereg[159]), .Z(n5526) );
  NAND U7735 ( .A(n5528), .B(n5529), .Z(n3698) );
  NANDN U7736 ( .A(init), .B(e[160]), .Z(n5529) );
  AND U7737 ( .A(n5530), .B(n5531), .Z(n5528) );
  NAND U7738 ( .A(ereg[159]), .B(n4895), .Z(n5531) );
  NANDN U7739 ( .A(n4890), .B(ereg[160]), .Z(n5530) );
  NAND U7740 ( .A(n5532), .B(n5533), .Z(n3697) );
  NANDN U7741 ( .A(init), .B(e[161]), .Z(n5533) );
  AND U7742 ( .A(n5534), .B(n5535), .Z(n5532) );
  NAND U7743 ( .A(ereg[160]), .B(n4895), .Z(n5535) );
  NANDN U7744 ( .A(n4890), .B(ereg[161]), .Z(n5534) );
  NAND U7745 ( .A(n5536), .B(n5537), .Z(n3696) );
  NANDN U7746 ( .A(init), .B(e[162]), .Z(n5537) );
  AND U7747 ( .A(n5538), .B(n5539), .Z(n5536) );
  NAND U7748 ( .A(ereg[161]), .B(n4895), .Z(n5539) );
  NANDN U7749 ( .A(n4890), .B(ereg[162]), .Z(n5538) );
  NAND U7750 ( .A(n5540), .B(n5541), .Z(n3695) );
  NANDN U7751 ( .A(init), .B(e[163]), .Z(n5541) );
  AND U7752 ( .A(n5542), .B(n5543), .Z(n5540) );
  NAND U7753 ( .A(ereg[162]), .B(n4895), .Z(n5543) );
  NANDN U7754 ( .A(n4890), .B(ereg[163]), .Z(n5542) );
  NAND U7755 ( .A(n5544), .B(n5545), .Z(n3694) );
  NANDN U7756 ( .A(init), .B(e[164]), .Z(n5545) );
  AND U7757 ( .A(n5546), .B(n5547), .Z(n5544) );
  NAND U7758 ( .A(ereg[163]), .B(n4895), .Z(n5547) );
  NANDN U7759 ( .A(n4890), .B(ereg[164]), .Z(n5546) );
  NAND U7760 ( .A(n5548), .B(n5549), .Z(n3693) );
  NANDN U7761 ( .A(init), .B(e[165]), .Z(n5549) );
  AND U7762 ( .A(n5550), .B(n5551), .Z(n5548) );
  NAND U7763 ( .A(ereg[164]), .B(n4895), .Z(n5551) );
  NANDN U7764 ( .A(n4890), .B(ereg[165]), .Z(n5550) );
  NAND U7765 ( .A(n5552), .B(n5553), .Z(n3692) );
  NANDN U7766 ( .A(init), .B(e[166]), .Z(n5553) );
  AND U7767 ( .A(n5554), .B(n5555), .Z(n5552) );
  NAND U7768 ( .A(ereg[165]), .B(n4895), .Z(n5555) );
  NANDN U7769 ( .A(n4890), .B(ereg[166]), .Z(n5554) );
  NAND U7770 ( .A(n5556), .B(n5557), .Z(n3691) );
  NANDN U7771 ( .A(init), .B(e[167]), .Z(n5557) );
  AND U7772 ( .A(n5558), .B(n5559), .Z(n5556) );
  NAND U7773 ( .A(ereg[166]), .B(n4895), .Z(n5559) );
  NANDN U7774 ( .A(n4890), .B(ereg[167]), .Z(n5558) );
  NAND U7775 ( .A(n5560), .B(n5561), .Z(n3690) );
  NANDN U7776 ( .A(init), .B(e[168]), .Z(n5561) );
  AND U7777 ( .A(n5562), .B(n5563), .Z(n5560) );
  NAND U7778 ( .A(ereg[167]), .B(n4895), .Z(n5563) );
  NANDN U7779 ( .A(n4890), .B(ereg[168]), .Z(n5562) );
  NAND U7780 ( .A(n5564), .B(n5565), .Z(n3689) );
  NANDN U7781 ( .A(init), .B(e[169]), .Z(n5565) );
  AND U7782 ( .A(n5566), .B(n5567), .Z(n5564) );
  NAND U7783 ( .A(ereg[168]), .B(n4895), .Z(n5567) );
  NANDN U7784 ( .A(n4890), .B(ereg[169]), .Z(n5566) );
  NAND U7785 ( .A(n5568), .B(n5569), .Z(n3688) );
  NANDN U7786 ( .A(init), .B(e[170]), .Z(n5569) );
  AND U7787 ( .A(n5570), .B(n5571), .Z(n5568) );
  NAND U7788 ( .A(ereg[169]), .B(n4895), .Z(n5571) );
  NANDN U7789 ( .A(n4890), .B(ereg[170]), .Z(n5570) );
  NAND U7790 ( .A(n5572), .B(n5573), .Z(n3687) );
  NANDN U7791 ( .A(init), .B(e[171]), .Z(n5573) );
  AND U7792 ( .A(n5574), .B(n5575), .Z(n5572) );
  NAND U7793 ( .A(ereg[170]), .B(n4895), .Z(n5575) );
  NANDN U7794 ( .A(n4890), .B(ereg[171]), .Z(n5574) );
  NAND U7795 ( .A(n5576), .B(n5577), .Z(n3686) );
  NANDN U7796 ( .A(init), .B(e[172]), .Z(n5577) );
  AND U7797 ( .A(n5578), .B(n5579), .Z(n5576) );
  NAND U7798 ( .A(ereg[171]), .B(n4895), .Z(n5579) );
  NANDN U7799 ( .A(n4890), .B(ereg[172]), .Z(n5578) );
  NAND U7800 ( .A(n5580), .B(n5581), .Z(n3685) );
  NANDN U7801 ( .A(init), .B(e[173]), .Z(n5581) );
  AND U7802 ( .A(n5582), .B(n5583), .Z(n5580) );
  NAND U7803 ( .A(ereg[172]), .B(n4895), .Z(n5583) );
  NANDN U7804 ( .A(n4890), .B(ereg[173]), .Z(n5582) );
  NAND U7805 ( .A(n5584), .B(n5585), .Z(n3684) );
  NANDN U7806 ( .A(init), .B(e[174]), .Z(n5585) );
  AND U7807 ( .A(n5586), .B(n5587), .Z(n5584) );
  NAND U7808 ( .A(ereg[173]), .B(n4895), .Z(n5587) );
  NANDN U7809 ( .A(n4890), .B(ereg[174]), .Z(n5586) );
  NAND U7810 ( .A(n5588), .B(n5589), .Z(n3683) );
  NANDN U7811 ( .A(init), .B(e[175]), .Z(n5589) );
  AND U7812 ( .A(n5590), .B(n5591), .Z(n5588) );
  NAND U7813 ( .A(ereg[174]), .B(n4895), .Z(n5591) );
  NANDN U7814 ( .A(n4890), .B(ereg[175]), .Z(n5590) );
  NAND U7815 ( .A(n5592), .B(n5593), .Z(n3682) );
  NANDN U7816 ( .A(init), .B(e[176]), .Z(n5593) );
  AND U7817 ( .A(n5594), .B(n5595), .Z(n5592) );
  NAND U7818 ( .A(ereg[175]), .B(n4895), .Z(n5595) );
  NANDN U7819 ( .A(n4890), .B(ereg[176]), .Z(n5594) );
  NAND U7820 ( .A(n5596), .B(n5597), .Z(n3681) );
  NANDN U7821 ( .A(init), .B(e[177]), .Z(n5597) );
  AND U7822 ( .A(n5598), .B(n5599), .Z(n5596) );
  NAND U7823 ( .A(ereg[176]), .B(n4895), .Z(n5599) );
  NANDN U7824 ( .A(n4890), .B(ereg[177]), .Z(n5598) );
  NAND U7825 ( .A(n5600), .B(n5601), .Z(n3680) );
  NANDN U7826 ( .A(init), .B(e[178]), .Z(n5601) );
  AND U7827 ( .A(n5602), .B(n5603), .Z(n5600) );
  NAND U7828 ( .A(ereg[177]), .B(n4895), .Z(n5603) );
  NANDN U7829 ( .A(n4890), .B(ereg[178]), .Z(n5602) );
  NAND U7830 ( .A(n5604), .B(n5605), .Z(n3679) );
  NANDN U7831 ( .A(init), .B(e[179]), .Z(n5605) );
  AND U7832 ( .A(n5606), .B(n5607), .Z(n5604) );
  NAND U7833 ( .A(ereg[178]), .B(n4895), .Z(n5607) );
  NANDN U7834 ( .A(n4890), .B(ereg[179]), .Z(n5606) );
  NAND U7835 ( .A(n5608), .B(n5609), .Z(n3678) );
  NANDN U7836 ( .A(init), .B(e[180]), .Z(n5609) );
  AND U7837 ( .A(n5610), .B(n5611), .Z(n5608) );
  NAND U7838 ( .A(ereg[179]), .B(n4895), .Z(n5611) );
  NANDN U7839 ( .A(n4890), .B(ereg[180]), .Z(n5610) );
  NAND U7840 ( .A(n5612), .B(n5613), .Z(n3677) );
  NANDN U7841 ( .A(init), .B(e[181]), .Z(n5613) );
  AND U7842 ( .A(n5614), .B(n5615), .Z(n5612) );
  NAND U7843 ( .A(ereg[180]), .B(n4895), .Z(n5615) );
  NANDN U7844 ( .A(n4890), .B(ereg[181]), .Z(n5614) );
  NAND U7845 ( .A(n5616), .B(n5617), .Z(n3676) );
  NANDN U7846 ( .A(init), .B(e[182]), .Z(n5617) );
  AND U7847 ( .A(n5618), .B(n5619), .Z(n5616) );
  NAND U7848 ( .A(ereg[181]), .B(n4895), .Z(n5619) );
  NANDN U7849 ( .A(n4890), .B(ereg[182]), .Z(n5618) );
  NAND U7850 ( .A(n5620), .B(n5621), .Z(n3675) );
  NANDN U7851 ( .A(init), .B(e[183]), .Z(n5621) );
  AND U7852 ( .A(n5622), .B(n5623), .Z(n5620) );
  NAND U7853 ( .A(ereg[182]), .B(n4895), .Z(n5623) );
  NANDN U7854 ( .A(n4890), .B(ereg[183]), .Z(n5622) );
  NAND U7855 ( .A(n5624), .B(n5625), .Z(n3674) );
  NANDN U7856 ( .A(init), .B(e[184]), .Z(n5625) );
  AND U7857 ( .A(n5626), .B(n5627), .Z(n5624) );
  NAND U7858 ( .A(ereg[183]), .B(n4895), .Z(n5627) );
  NANDN U7859 ( .A(n4890), .B(ereg[184]), .Z(n5626) );
  NAND U7860 ( .A(n5628), .B(n5629), .Z(n3673) );
  NANDN U7861 ( .A(init), .B(e[185]), .Z(n5629) );
  AND U7862 ( .A(n5630), .B(n5631), .Z(n5628) );
  NAND U7863 ( .A(ereg[184]), .B(n4895), .Z(n5631) );
  NANDN U7864 ( .A(n4890), .B(ereg[185]), .Z(n5630) );
  NAND U7865 ( .A(n5632), .B(n5633), .Z(n3672) );
  NANDN U7866 ( .A(init), .B(e[186]), .Z(n5633) );
  AND U7867 ( .A(n5634), .B(n5635), .Z(n5632) );
  NAND U7868 ( .A(ereg[185]), .B(n4895), .Z(n5635) );
  NANDN U7869 ( .A(n4890), .B(ereg[186]), .Z(n5634) );
  NAND U7870 ( .A(n5636), .B(n5637), .Z(n3671) );
  NANDN U7871 ( .A(init), .B(e[187]), .Z(n5637) );
  AND U7872 ( .A(n5638), .B(n5639), .Z(n5636) );
  NAND U7873 ( .A(ereg[186]), .B(n4895), .Z(n5639) );
  NANDN U7874 ( .A(n4890), .B(ereg[187]), .Z(n5638) );
  NAND U7875 ( .A(n5640), .B(n5641), .Z(n3670) );
  NANDN U7876 ( .A(init), .B(e[188]), .Z(n5641) );
  AND U7877 ( .A(n5642), .B(n5643), .Z(n5640) );
  NAND U7878 ( .A(ereg[187]), .B(n4895), .Z(n5643) );
  NANDN U7879 ( .A(n4890), .B(ereg[188]), .Z(n5642) );
  NAND U7880 ( .A(n5644), .B(n5645), .Z(n3669) );
  NANDN U7881 ( .A(init), .B(e[189]), .Z(n5645) );
  AND U7882 ( .A(n5646), .B(n5647), .Z(n5644) );
  NAND U7883 ( .A(ereg[188]), .B(n4895), .Z(n5647) );
  NANDN U7884 ( .A(n4890), .B(ereg[189]), .Z(n5646) );
  NAND U7885 ( .A(n5648), .B(n5649), .Z(n3668) );
  NANDN U7886 ( .A(init), .B(e[190]), .Z(n5649) );
  AND U7887 ( .A(n5650), .B(n5651), .Z(n5648) );
  NAND U7888 ( .A(ereg[189]), .B(n4895), .Z(n5651) );
  NANDN U7889 ( .A(n4890), .B(ereg[190]), .Z(n5650) );
  NAND U7890 ( .A(n5652), .B(n5653), .Z(n3667) );
  NANDN U7891 ( .A(init), .B(e[191]), .Z(n5653) );
  AND U7892 ( .A(n5654), .B(n5655), .Z(n5652) );
  NAND U7893 ( .A(ereg[190]), .B(n4895), .Z(n5655) );
  NANDN U7894 ( .A(n4890), .B(ereg[191]), .Z(n5654) );
  NAND U7895 ( .A(n5656), .B(n5657), .Z(n3666) );
  NANDN U7896 ( .A(init), .B(e[192]), .Z(n5657) );
  AND U7897 ( .A(n5658), .B(n5659), .Z(n5656) );
  NAND U7898 ( .A(ereg[191]), .B(n4895), .Z(n5659) );
  NANDN U7899 ( .A(n4890), .B(ereg[192]), .Z(n5658) );
  NAND U7900 ( .A(n5660), .B(n5661), .Z(n3665) );
  NANDN U7901 ( .A(init), .B(e[193]), .Z(n5661) );
  AND U7902 ( .A(n5662), .B(n5663), .Z(n5660) );
  NAND U7903 ( .A(ereg[192]), .B(n4895), .Z(n5663) );
  NANDN U7904 ( .A(n4890), .B(ereg[193]), .Z(n5662) );
  NAND U7905 ( .A(n5664), .B(n5665), .Z(n3664) );
  NANDN U7906 ( .A(init), .B(e[194]), .Z(n5665) );
  AND U7907 ( .A(n5666), .B(n5667), .Z(n5664) );
  NAND U7908 ( .A(ereg[193]), .B(n4895), .Z(n5667) );
  NANDN U7909 ( .A(n4890), .B(ereg[194]), .Z(n5666) );
  NAND U7910 ( .A(n5668), .B(n5669), .Z(n3663) );
  NANDN U7911 ( .A(init), .B(e[195]), .Z(n5669) );
  AND U7912 ( .A(n5670), .B(n5671), .Z(n5668) );
  NAND U7913 ( .A(ereg[194]), .B(n4895), .Z(n5671) );
  NANDN U7914 ( .A(n4890), .B(ereg[195]), .Z(n5670) );
  NAND U7915 ( .A(n5672), .B(n5673), .Z(n3662) );
  NANDN U7916 ( .A(init), .B(e[196]), .Z(n5673) );
  AND U7917 ( .A(n5674), .B(n5675), .Z(n5672) );
  NAND U7918 ( .A(ereg[195]), .B(n4895), .Z(n5675) );
  NANDN U7919 ( .A(n4890), .B(ereg[196]), .Z(n5674) );
  NAND U7920 ( .A(n5676), .B(n5677), .Z(n3661) );
  NANDN U7921 ( .A(init), .B(e[197]), .Z(n5677) );
  AND U7922 ( .A(n5678), .B(n5679), .Z(n5676) );
  NAND U7923 ( .A(ereg[196]), .B(n4895), .Z(n5679) );
  NANDN U7924 ( .A(n4890), .B(ereg[197]), .Z(n5678) );
  NAND U7925 ( .A(n5680), .B(n5681), .Z(n3660) );
  NANDN U7926 ( .A(init), .B(e[198]), .Z(n5681) );
  AND U7927 ( .A(n5682), .B(n5683), .Z(n5680) );
  NAND U7928 ( .A(ereg[197]), .B(n4895), .Z(n5683) );
  NANDN U7929 ( .A(n4890), .B(ereg[198]), .Z(n5682) );
  NAND U7930 ( .A(n5684), .B(n5685), .Z(n3659) );
  NANDN U7931 ( .A(init), .B(e[199]), .Z(n5685) );
  AND U7932 ( .A(n5686), .B(n5687), .Z(n5684) );
  NAND U7933 ( .A(ereg[198]), .B(n4895), .Z(n5687) );
  NANDN U7934 ( .A(n4890), .B(ereg[199]), .Z(n5686) );
  NAND U7935 ( .A(n5688), .B(n5689), .Z(n3658) );
  NANDN U7936 ( .A(init), .B(e[200]), .Z(n5689) );
  AND U7937 ( .A(n5690), .B(n5691), .Z(n5688) );
  NAND U7938 ( .A(ereg[199]), .B(n4895), .Z(n5691) );
  NANDN U7939 ( .A(n4890), .B(ereg[200]), .Z(n5690) );
  NAND U7940 ( .A(n5692), .B(n5693), .Z(n3657) );
  NANDN U7941 ( .A(init), .B(e[201]), .Z(n5693) );
  AND U7942 ( .A(n5694), .B(n5695), .Z(n5692) );
  NAND U7943 ( .A(ereg[200]), .B(n4895), .Z(n5695) );
  NANDN U7944 ( .A(n4890), .B(ereg[201]), .Z(n5694) );
  NAND U7945 ( .A(n5696), .B(n5697), .Z(n3656) );
  NANDN U7946 ( .A(init), .B(e[202]), .Z(n5697) );
  AND U7947 ( .A(n5698), .B(n5699), .Z(n5696) );
  NAND U7948 ( .A(ereg[201]), .B(n4895), .Z(n5699) );
  NANDN U7949 ( .A(n4890), .B(ereg[202]), .Z(n5698) );
  NAND U7950 ( .A(n5700), .B(n5701), .Z(n3655) );
  NANDN U7951 ( .A(init), .B(e[203]), .Z(n5701) );
  AND U7952 ( .A(n5702), .B(n5703), .Z(n5700) );
  NAND U7953 ( .A(ereg[202]), .B(n4895), .Z(n5703) );
  NANDN U7954 ( .A(n4890), .B(ereg[203]), .Z(n5702) );
  NAND U7955 ( .A(n5704), .B(n5705), .Z(n3654) );
  NANDN U7956 ( .A(init), .B(e[204]), .Z(n5705) );
  AND U7957 ( .A(n5706), .B(n5707), .Z(n5704) );
  NAND U7958 ( .A(ereg[203]), .B(n4895), .Z(n5707) );
  NANDN U7959 ( .A(n4890), .B(ereg[204]), .Z(n5706) );
  NAND U7960 ( .A(n5708), .B(n5709), .Z(n3653) );
  NANDN U7961 ( .A(init), .B(e[205]), .Z(n5709) );
  AND U7962 ( .A(n5710), .B(n5711), .Z(n5708) );
  NAND U7963 ( .A(ereg[204]), .B(n4895), .Z(n5711) );
  NANDN U7964 ( .A(n4890), .B(ereg[205]), .Z(n5710) );
  NAND U7965 ( .A(n5712), .B(n5713), .Z(n3652) );
  NANDN U7966 ( .A(init), .B(e[206]), .Z(n5713) );
  AND U7967 ( .A(n5714), .B(n5715), .Z(n5712) );
  NAND U7968 ( .A(ereg[205]), .B(n4895), .Z(n5715) );
  NANDN U7969 ( .A(n4890), .B(ereg[206]), .Z(n5714) );
  NAND U7970 ( .A(n5716), .B(n5717), .Z(n3651) );
  NANDN U7971 ( .A(init), .B(e[207]), .Z(n5717) );
  AND U7972 ( .A(n5718), .B(n5719), .Z(n5716) );
  NAND U7973 ( .A(ereg[206]), .B(n4895), .Z(n5719) );
  NANDN U7974 ( .A(n4890), .B(ereg[207]), .Z(n5718) );
  NAND U7975 ( .A(n5720), .B(n5721), .Z(n3650) );
  NANDN U7976 ( .A(init), .B(e[208]), .Z(n5721) );
  AND U7977 ( .A(n5722), .B(n5723), .Z(n5720) );
  NAND U7978 ( .A(ereg[207]), .B(n4895), .Z(n5723) );
  NANDN U7979 ( .A(n4890), .B(ereg[208]), .Z(n5722) );
  NAND U7980 ( .A(n5724), .B(n5725), .Z(n3649) );
  NANDN U7981 ( .A(init), .B(e[209]), .Z(n5725) );
  AND U7982 ( .A(n5726), .B(n5727), .Z(n5724) );
  NAND U7983 ( .A(ereg[208]), .B(n4895), .Z(n5727) );
  NANDN U7984 ( .A(n4890), .B(ereg[209]), .Z(n5726) );
  NAND U7985 ( .A(n5728), .B(n5729), .Z(n3648) );
  NANDN U7986 ( .A(init), .B(e[210]), .Z(n5729) );
  AND U7987 ( .A(n5730), .B(n5731), .Z(n5728) );
  NAND U7988 ( .A(ereg[209]), .B(n4895), .Z(n5731) );
  NANDN U7989 ( .A(n4890), .B(ereg[210]), .Z(n5730) );
  NAND U7990 ( .A(n5732), .B(n5733), .Z(n3647) );
  NANDN U7991 ( .A(init), .B(e[211]), .Z(n5733) );
  AND U7992 ( .A(n5734), .B(n5735), .Z(n5732) );
  NAND U7993 ( .A(ereg[210]), .B(n4895), .Z(n5735) );
  NANDN U7994 ( .A(n4890), .B(ereg[211]), .Z(n5734) );
  NAND U7995 ( .A(n5736), .B(n5737), .Z(n3646) );
  NANDN U7996 ( .A(init), .B(e[212]), .Z(n5737) );
  AND U7997 ( .A(n5738), .B(n5739), .Z(n5736) );
  NAND U7998 ( .A(ereg[211]), .B(n4895), .Z(n5739) );
  NANDN U7999 ( .A(n4890), .B(ereg[212]), .Z(n5738) );
  NAND U8000 ( .A(n5740), .B(n5741), .Z(n3645) );
  NANDN U8001 ( .A(init), .B(e[213]), .Z(n5741) );
  AND U8002 ( .A(n5742), .B(n5743), .Z(n5740) );
  NAND U8003 ( .A(ereg[212]), .B(n4895), .Z(n5743) );
  NANDN U8004 ( .A(n4890), .B(ereg[213]), .Z(n5742) );
  NAND U8005 ( .A(n5744), .B(n5745), .Z(n3644) );
  NANDN U8006 ( .A(init), .B(e[214]), .Z(n5745) );
  AND U8007 ( .A(n5746), .B(n5747), .Z(n5744) );
  NAND U8008 ( .A(ereg[213]), .B(n4895), .Z(n5747) );
  NANDN U8009 ( .A(n4890), .B(ereg[214]), .Z(n5746) );
  NAND U8010 ( .A(n5748), .B(n5749), .Z(n3643) );
  NANDN U8011 ( .A(init), .B(e[215]), .Z(n5749) );
  AND U8012 ( .A(n5750), .B(n5751), .Z(n5748) );
  NAND U8013 ( .A(ereg[214]), .B(n4895), .Z(n5751) );
  NANDN U8014 ( .A(n4890), .B(ereg[215]), .Z(n5750) );
  NAND U8015 ( .A(n5752), .B(n5753), .Z(n3642) );
  NANDN U8016 ( .A(init), .B(e[216]), .Z(n5753) );
  AND U8017 ( .A(n5754), .B(n5755), .Z(n5752) );
  NAND U8018 ( .A(ereg[215]), .B(n4895), .Z(n5755) );
  NANDN U8019 ( .A(n4890), .B(ereg[216]), .Z(n5754) );
  NAND U8020 ( .A(n5756), .B(n5757), .Z(n3641) );
  NANDN U8021 ( .A(init), .B(e[217]), .Z(n5757) );
  AND U8022 ( .A(n5758), .B(n5759), .Z(n5756) );
  NAND U8023 ( .A(ereg[216]), .B(n4895), .Z(n5759) );
  NANDN U8024 ( .A(n4890), .B(ereg[217]), .Z(n5758) );
  NAND U8025 ( .A(n5760), .B(n5761), .Z(n3640) );
  NANDN U8026 ( .A(init), .B(e[218]), .Z(n5761) );
  AND U8027 ( .A(n5762), .B(n5763), .Z(n5760) );
  NAND U8028 ( .A(ereg[217]), .B(n4895), .Z(n5763) );
  NANDN U8029 ( .A(n4890), .B(ereg[218]), .Z(n5762) );
  NAND U8030 ( .A(n5764), .B(n5765), .Z(n3639) );
  NANDN U8031 ( .A(init), .B(e[219]), .Z(n5765) );
  AND U8032 ( .A(n5766), .B(n5767), .Z(n5764) );
  NAND U8033 ( .A(ereg[218]), .B(n4895), .Z(n5767) );
  NANDN U8034 ( .A(n4890), .B(ereg[219]), .Z(n5766) );
  NAND U8035 ( .A(n5768), .B(n5769), .Z(n3638) );
  NANDN U8036 ( .A(init), .B(e[220]), .Z(n5769) );
  AND U8037 ( .A(n5770), .B(n5771), .Z(n5768) );
  NAND U8038 ( .A(ereg[219]), .B(n4895), .Z(n5771) );
  NANDN U8039 ( .A(n4890), .B(ereg[220]), .Z(n5770) );
  NAND U8040 ( .A(n5772), .B(n5773), .Z(n3637) );
  NANDN U8041 ( .A(init), .B(e[221]), .Z(n5773) );
  AND U8042 ( .A(n5774), .B(n5775), .Z(n5772) );
  NAND U8043 ( .A(ereg[220]), .B(n4895), .Z(n5775) );
  NANDN U8044 ( .A(n4890), .B(ereg[221]), .Z(n5774) );
  NAND U8045 ( .A(n5776), .B(n5777), .Z(n3636) );
  NANDN U8046 ( .A(init), .B(e[222]), .Z(n5777) );
  AND U8047 ( .A(n5778), .B(n5779), .Z(n5776) );
  NAND U8048 ( .A(ereg[221]), .B(n4895), .Z(n5779) );
  NANDN U8049 ( .A(n4890), .B(ereg[222]), .Z(n5778) );
  NAND U8050 ( .A(n5780), .B(n5781), .Z(n3635) );
  NANDN U8051 ( .A(init), .B(e[223]), .Z(n5781) );
  AND U8052 ( .A(n5782), .B(n5783), .Z(n5780) );
  NAND U8053 ( .A(ereg[222]), .B(n4895), .Z(n5783) );
  NANDN U8054 ( .A(n4890), .B(ereg[223]), .Z(n5782) );
  NAND U8055 ( .A(n5784), .B(n5785), .Z(n3634) );
  NANDN U8056 ( .A(init), .B(e[224]), .Z(n5785) );
  AND U8057 ( .A(n5786), .B(n5787), .Z(n5784) );
  NAND U8058 ( .A(ereg[223]), .B(n4895), .Z(n5787) );
  NANDN U8059 ( .A(n4890), .B(ereg[224]), .Z(n5786) );
  NAND U8060 ( .A(n5788), .B(n5789), .Z(n3633) );
  NANDN U8061 ( .A(init), .B(e[225]), .Z(n5789) );
  AND U8062 ( .A(n5790), .B(n5791), .Z(n5788) );
  NAND U8063 ( .A(ereg[224]), .B(n4895), .Z(n5791) );
  NANDN U8064 ( .A(n4890), .B(ereg[225]), .Z(n5790) );
  NAND U8065 ( .A(n5792), .B(n5793), .Z(n3632) );
  NANDN U8066 ( .A(init), .B(e[226]), .Z(n5793) );
  AND U8067 ( .A(n5794), .B(n5795), .Z(n5792) );
  NAND U8068 ( .A(ereg[225]), .B(n4895), .Z(n5795) );
  NANDN U8069 ( .A(n4890), .B(ereg[226]), .Z(n5794) );
  NAND U8070 ( .A(n5796), .B(n5797), .Z(n3631) );
  NANDN U8071 ( .A(init), .B(e[227]), .Z(n5797) );
  AND U8072 ( .A(n5798), .B(n5799), .Z(n5796) );
  NAND U8073 ( .A(ereg[226]), .B(n4895), .Z(n5799) );
  NANDN U8074 ( .A(n4890), .B(ereg[227]), .Z(n5798) );
  NAND U8075 ( .A(n5800), .B(n5801), .Z(n3630) );
  NANDN U8076 ( .A(init), .B(e[228]), .Z(n5801) );
  AND U8077 ( .A(n5802), .B(n5803), .Z(n5800) );
  NAND U8078 ( .A(ereg[227]), .B(n4895), .Z(n5803) );
  NANDN U8079 ( .A(n4890), .B(ereg[228]), .Z(n5802) );
  NAND U8080 ( .A(n5804), .B(n5805), .Z(n3629) );
  NANDN U8081 ( .A(init), .B(e[229]), .Z(n5805) );
  AND U8082 ( .A(n5806), .B(n5807), .Z(n5804) );
  NAND U8083 ( .A(ereg[228]), .B(n4895), .Z(n5807) );
  NANDN U8084 ( .A(n4890), .B(ereg[229]), .Z(n5806) );
  NAND U8085 ( .A(n5808), .B(n5809), .Z(n3628) );
  NANDN U8086 ( .A(init), .B(e[230]), .Z(n5809) );
  AND U8087 ( .A(n5810), .B(n5811), .Z(n5808) );
  NAND U8088 ( .A(ereg[229]), .B(n4895), .Z(n5811) );
  NANDN U8089 ( .A(n4890), .B(ereg[230]), .Z(n5810) );
  NAND U8090 ( .A(n5812), .B(n5813), .Z(n3627) );
  NANDN U8091 ( .A(init), .B(e[231]), .Z(n5813) );
  AND U8092 ( .A(n5814), .B(n5815), .Z(n5812) );
  NAND U8093 ( .A(ereg[230]), .B(n4895), .Z(n5815) );
  NANDN U8094 ( .A(n4890), .B(ereg[231]), .Z(n5814) );
  NAND U8095 ( .A(n5816), .B(n5817), .Z(n3626) );
  NANDN U8096 ( .A(init), .B(e[232]), .Z(n5817) );
  AND U8097 ( .A(n5818), .B(n5819), .Z(n5816) );
  NAND U8098 ( .A(ereg[231]), .B(n4895), .Z(n5819) );
  NANDN U8099 ( .A(n4890), .B(ereg[232]), .Z(n5818) );
  NAND U8100 ( .A(n5820), .B(n5821), .Z(n3625) );
  NANDN U8101 ( .A(init), .B(e[233]), .Z(n5821) );
  AND U8102 ( .A(n5822), .B(n5823), .Z(n5820) );
  NAND U8103 ( .A(ereg[232]), .B(n4895), .Z(n5823) );
  NANDN U8104 ( .A(n4890), .B(ereg[233]), .Z(n5822) );
  NAND U8105 ( .A(n5824), .B(n5825), .Z(n3624) );
  NANDN U8106 ( .A(init), .B(e[234]), .Z(n5825) );
  AND U8107 ( .A(n5826), .B(n5827), .Z(n5824) );
  NAND U8108 ( .A(ereg[233]), .B(n4895), .Z(n5827) );
  NANDN U8109 ( .A(n4890), .B(ereg[234]), .Z(n5826) );
  NAND U8110 ( .A(n5828), .B(n5829), .Z(n3623) );
  NANDN U8111 ( .A(init), .B(e[235]), .Z(n5829) );
  AND U8112 ( .A(n5830), .B(n5831), .Z(n5828) );
  NAND U8113 ( .A(ereg[234]), .B(n4895), .Z(n5831) );
  NANDN U8114 ( .A(n4890), .B(ereg[235]), .Z(n5830) );
  NAND U8115 ( .A(n5832), .B(n5833), .Z(n3622) );
  NANDN U8116 ( .A(init), .B(e[236]), .Z(n5833) );
  AND U8117 ( .A(n5834), .B(n5835), .Z(n5832) );
  NAND U8118 ( .A(ereg[235]), .B(n4895), .Z(n5835) );
  NANDN U8119 ( .A(n4890), .B(ereg[236]), .Z(n5834) );
  NAND U8120 ( .A(n5836), .B(n5837), .Z(n3621) );
  NANDN U8121 ( .A(init), .B(e[237]), .Z(n5837) );
  AND U8122 ( .A(n5838), .B(n5839), .Z(n5836) );
  NAND U8123 ( .A(ereg[236]), .B(n4895), .Z(n5839) );
  NANDN U8124 ( .A(n4890), .B(ereg[237]), .Z(n5838) );
  NAND U8125 ( .A(n5840), .B(n5841), .Z(n3620) );
  NANDN U8126 ( .A(init), .B(e[238]), .Z(n5841) );
  AND U8127 ( .A(n5842), .B(n5843), .Z(n5840) );
  NAND U8128 ( .A(ereg[237]), .B(n4895), .Z(n5843) );
  NANDN U8129 ( .A(n4890), .B(ereg[238]), .Z(n5842) );
  NAND U8130 ( .A(n5844), .B(n5845), .Z(n3619) );
  NANDN U8131 ( .A(init), .B(e[239]), .Z(n5845) );
  AND U8132 ( .A(n5846), .B(n5847), .Z(n5844) );
  NAND U8133 ( .A(ereg[238]), .B(n4895), .Z(n5847) );
  NANDN U8134 ( .A(n4890), .B(ereg[239]), .Z(n5846) );
  NAND U8135 ( .A(n5848), .B(n5849), .Z(n3618) );
  NANDN U8136 ( .A(init), .B(e[240]), .Z(n5849) );
  AND U8137 ( .A(n5850), .B(n5851), .Z(n5848) );
  NAND U8138 ( .A(ereg[239]), .B(n4895), .Z(n5851) );
  NANDN U8139 ( .A(n4890), .B(ereg[240]), .Z(n5850) );
  NAND U8140 ( .A(n5852), .B(n5853), .Z(n3617) );
  NANDN U8141 ( .A(init), .B(e[241]), .Z(n5853) );
  AND U8142 ( .A(n5854), .B(n5855), .Z(n5852) );
  NAND U8143 ( .A(ereg[240]), .B(n4895), .Z(n5855) );
  NANDN U8144 ( .A(n4890), .B(ereg[241]), .Z(n5854) );
  NAND U8145 ( .A(n5856), .B(n5857), .Z(n3616) );
  NANDN U8146 ( .A(init), .B(e[242]), .Z(n5857) );
  AND U8147 ( .A(n5858), .B(n5859), .Z(n5856) );
  NAND U8148 ( .A(ereg[241]), .B(n4895), .Z(n5859) );
  NANDN U8149 ( .A(n4890), .B(ereg[242]), .Z(n5858) );
  NAND U8150 ( .A(n5860), .B(n5861), .Z(n3615) );
  NANDN U8151 ( .A(init), .B(e[243]), .Z(n5861) );
  AND U8152 ( .A(n5862), .B(n5863), .Z(n5860) );
  NAND U8153 ( .A(ereg[242]), .B(n4895), .Z(n5863) );
  NANDN U8154 ( .A(n4890), .B(ereg[243]), .Z(n5862) );
  NAND U8155 ( .A(n5864), .B(n5865), .Z(n3614) );
  NANDN U8156 ( .A(init), .B(e[244]), .Z(n5865) );
  AND U8157 ( .A(n5866), .B(n5867), .Z(n5864) );
  NAND U8158 ( .A(ereg[243]), .B(n4895), .Z(n5867) );
  NANDN U8159 ( .A(n4890), .B(ereg[244]), .Z(n5866) );
  NAND U8160 ( .A(n5868), .B(n5869), .Z(n3613) );
  NANDN U8161 ( .A(init), .B(e[245]), .Z(n5869) );
  AND U8162 ( .A(n5870), .B(n5871), .Z(n5868) );
  NAND U8163 ( .A(ereg[244]), .B(n4895), .Z(n5871) );
  NANDN U8164 ( .A(n4890), .B(ereg[245]), .Z(n5870) );
  NAND U8165 ( .A(n5872), .B(n5873), .Z(n3612) );
  NANDN U8166 ( .A(init), .B(e[246]), .Z(n5873) );
  AND U8167 ( .A(n5874), .B(n5875), .Z(n5872) );
  NAND U8168 ( .A(ereg[245]), .B(n4895), .Z(n5875) );
  NANDN U8169 ( .A(n4890), .B(ereg[246]), .Z(n5874) );
  NAND U8170 ( .A(n5876), .B(n5877), .Z(n3611) );
  NANDN U8171 ( .A(init), .B(e[247]), .Z(n5877) );
  AND U8172 ( .A(n5878), .B(n5879), .Z(n5876) );
  NAND U8173 ( .A(ereg[246]), .B(n4895), .Z(n5879) );
  NANDN U8174 ( .A(n4890), .B(ereg[247]), .Z(n5878) );
  NAND U8175 ( .A(n5880), .B(n5881), .Z(n3610) );
  NANDN U8176 ( .A(init), .B(e[248]), .Z(n5881) );
  AND U8177 ( .A(n5882), .B(n5883), .Z(n5880) );
  NAND U8178 ( .A(ereg[247]), .B(n4895), .Z(n5883) );
  NANDN U8179 ( .A(n4890), .B(ereg[248]), .Z(n5882) );
  NAND U8180 ( .A(n5884), .B(n5885), .Z(n3609) );
  NANDN U8181 ( .A(init), .B(e[249]), .Z(n5885) );
  AND U8182 ( .A(n5886), .B(n5887), .Z(n5884) );
  NAND U8183 ( .A(ereg[248]), .B(n4895), .Z(n5887) );
  NANDN U8184 ( .A(n4890), .B(ereg[249]), .Z(n5886) );
  NAND U8185 ( .A(n5888), .B(n5889), .Z(n3608) );
  NANDN U8186 ( .A(init), .B(e[250]), .Z(n5889) );
  AND U8187 ( .A(n5890), .B(n5891), .Z(n5888) );
  NAND U8188 ( .A(ereg[249]), .B(n4895), .Z(n5891) );
  NANDN U8189 ( .A(n4890), .B(ereg[250]), .Z(n5890) );
  NAND U8190 ( .A(n5892), .B(n5893), .Z(n3607) );
  NANDN U8191 ( .A(init), .B(e[251]), .Z(n5893) );
  AND U8192 ( .A(n5894), .B(n5895), .Z(n5892) );
  NAND U8193 ( .A(ereg[250]), .B(n4895), .Z(n5895) );
  NANDN U8194 ( .A(n4890), .B(ereg[251]), .Z(n5894) );
  NAND U8195 ( .A(n5896), .B(n5897), .Z(n3606) );
  NANDN U8196 ( .A(init), .B(e[252]), .Z(n5897) );
  AND U8197 ( .A(n5898), .B(n5899), .Z(n5896) );
  NAND U8198 ( .A(ereg[251]), .B(n4895), .Z(n5899) );
  NANDN U8199 ( .A(n4890), .B(ereg[252]), .Z(n5898) );
  NAND U8200 ( .A(n5900), .B(n5901), .Z(n3605) );
  NANDN U8201 ( .A(init), .B(e[253]), .Z(n5901) );
  AND U8202 ( .A(n5902), .B(n5903), .Z(n5900) );
  NAND U8203 ( .A(ereg[252]), .B(n4895), .Z(n5903) );
  NANDN U8204 ( .A(n4890), .B(ereg[253]), .Z(n5902) );
  NAND U8205 ( .A(n5904), .B(n5905), .Z(n3604) );
  NANDN U8206 ( .A(init), .B(e[254]), .Z(n5905) );
  AND U8207 ( .A(n5906), .B(n5907), .Z(n5904) );
  NAND U8208 ( .A(ereg[253]), .B(n4895), .Z(n5907) );
  NANDN U8209 ( .A(n4890), .B(ereg[254]), .Z(n5906) );
  NAND U8210 ( .A(n5908), .B(n5909), .Z(n3603) );
  NANDN U8211 ( .A(init), .B(e[255]), .Z(n5909) );
  AND U8212 ( .A(n5910), .B(n5911), .Z(n5908) );
  NAND U8213 ( .A(ereg[254]), .B(n4895), .Z(n5911) );
  AND U8214 ( .A(n4890), .B(start_in[511]), .Z(n4895) );
  NANDN U8215 ( .A(n4890), .B(ereg[255]), .Z(n5910) );
  AND U8216 ( .A(n5912), .B(n3862), .Z(n4890) );
  NANDN U8217 ( .A(mul_pow), .B(init), .Z(n3862) );
  NANDN U8218 ( .A(start_reg[511]), .B(init), .Z(n5912) );
  NAND U8219 ( .A(n5913), .B(n4541), .Z(n3602) );
  NANDN U8220 ( .A(init), .B(m[255]), .Z(n4541) );
  AND U8221 ( .A(n5914), .B(n5915), .Z(n5913) );
  NAND U8222 ( .A(o[255]), .B(n5916), .Z(n5915) );
  NANDN U8223 ( .A(n5917), .B(creg[255]), .Z(n5914) );
  NAND U8224 ( .A(n5918), .B(n4885), .Z(n3601) );
  NANDN U8225 ( .A(init), .B(m[0]), .Z(n4885) );
  AND U8226 ( .A(n5919), .B(n5920), .Z(n5918) );
  NAND U8227 ( .A(o[0]), .B(n5916), .Z(n5920) );
  NANDN U8228 ( .A(n5917), .B(creg[0]), .Z(n5919) );
  NAND U8229 ( .A(n5921), .B(n4663), .Z(n3600) );
  NANDN U8230 ( .A(init), .B(m[1]), .Z(n4663) );
  AND U8231 ( .A(n5922), .B(n5923), .Z(n5921) );
  NAND U8232 ( .A(o[1]), .B(n5916), .Z(n5923) );
  NANDN U8233 ( .A(n5917), .B(creg[1]), .Z(n5922) );
  NAND U8234 ( .A(n5924), .B(n4529), .Z(n3599) );
  NANDN U8235 ( .A(init), .B(m[2]), .Z(n4529) );
  AND U8236 ( .A(n5925), .B(n5926), .Z(n5924) );
  NAND U8237 ( .A(o[2]), .B(n5916), .Z(n5926) );
  NANDN U8238 ( .A(n5917), .B(creg[2]), .Z(n5925) );
  NAND U8239 ( .A(n5927), .B(n4507), .Z(n3598) );
  NANDN U8240 ( .A(init), .B(m[3]), .Z(n4507) );
  AND U8241 ( .A(n5928), .B(n5929), .Z(n5927) );
  NAND U8242 ( .A(o[3]), .B(n5916), .Z(n5929) );
  NANDN U8243 ( .A(n5917), .B(creg[3]), .Z(n5928) );
  NAND U8244 ( .A(n5930), .B(n4485), .Z(n3597) );
  NANDN U8245 ( .A(init), .B(m[4]), .Z(n4485) );
  AND U8246 ( .A(n5931), .B(n5932), .Z(n5930) );
  NAND U8247 ( .A(o[4]), .B(n5916), .Z(n5932) );
  NANDN U8248 ( .A(n5917), .B(creg[4]), .Z(n5931) );
  NAND U8249 ( .A(n5933), .B(n4463), .Z(n3596) );
  NANDN U8250 ( .A(init), .B(m[5]), .Z(n4463) );
  AND U8251 ( .A(n5934), .B(n5935), .Z(n5933) );
  NAND U8252 ( .A(o[5]), .B(n5916), .Z(n5935) );
  NANDN U8253 ( .A(n5917), .B(creg[5]), .Z(n5934) );
  NAND U8254 ( .A(n5936), .B(n4441), .Z(n3595) );
  NANDN U8255 ( .A(init), .B(m[6]), .Z(n4441) );
  AND U8256 ( .A(n5937), .B(n5938), .Z(n5936) );
  NAND U8257 ( .A(o[6]), .B(n5916), .Z(n5938) );
  NANDN U8258 ( .A(n5917), .B(creg[6]), .Z(n5937) );
  NAND U8259 ( .A(n5939), .B(n4419), .Z(n3594) );
  NANDN U8260 ( .A(init), .B(m[7]), .Z(n4419) );
  AND U8261 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U8262 ( .A(o[7]), .B(n5916), .Z(n5941) );
  NANDN U8263 ( .A(n5917), .B(creg[7]), .Z(n5940) );
  NAND U8264 ( .A(n5942), .B(n4397), .Z(n3593) );
  NANDN U8265 ( .A(init), .B(m[8]), .Z(n4397) );
  AND U8266 ( .A(n5943), .B(n5944), .Z(n5942) );
  NAND U8267 ( .A(o[8]), .B(n5916), .Z(n5944) );
  NANDN U8268 ( .A(n5917), .B(creg[8]), .Z(n5943) );
  NAND U8269 ( .A(n5945), .B(n4375), .Z(n3592) );
  NANDN U8270 ( .A(init), .B(m[9]), .Z(n4375) );
  AND U8271 ( .A(n5946), .B(n5947), .Z(n5945) );
  NAND U8272 ( .A(o[9]), .B(n5916), .Z(n5947) );
  NANDN U8273 ( .A(n5917), .B(creg[9]), .Z(n5946) );
  NAND U8274 ( .A(n5948), .B(n4863), .Z(n3591) );
  NANDN U8275 ( .A(init), .B(m[10]), .Z(n4863) );
  AND U8276 ( .A(n5949), .B(n5950), .Z(n5948) );
  NAND U8277 ( .A(o[10]), .B(n5916), .Z(n5950) );
  NANDN U8278 ( .A(n5917), .B(creg[10]), .Z(n5949) );
  NAND U8279 ( .A(n5951), .B(n4841), .Z(n3590) );
  NANDN U8280 ( .A(init), .B(m[11]), .Z(n4841) );
  AND U8281 ( .A(n5952), .B(n5953), .Z(n5951) );
  NAND U8282 ( .A(o[11]), .B(n5916), .Z(n5953) );
  NANDN U8283 ( .A(n5917), .B(creg[11]), .Z(n5952) );
  NAND U8284 ( .A(n5954), .B(n4819), .Z(n3589) );
  NANDN U8285 ( .A(init), .B(m[12]), .Z(n4819) );
  AND U8286 ( .A(n5955), .B(n5956), .Z(n5954) );
  NAND U8287 ( .A(o[12]), .B(n5916), .Z(n5956) );
  NANDN U8288 ( .A(n5917), .B(creg[12]), .Z(n5955) );
  NAND U8289 ( .A(n5957), .B(n4797), .Z(n3588) );
  NANDN U8290 ( .A(init), .B(m[13]), .Z(n4797) );
  AND U8291 ( .A(n5958), .B(n5959), .Z(n5957) );
  NAND U8292 ( .A(o[13]), .B(n5916), .Z(n5959) );
  NANDN U8293 ( .A(n5917), .B(creg[13]), .Z(n5958) );
  NAND U8294 ( .A(n5960), .B(n4775), .Z(n3587) );
  NANDN U8295 ( .A(init), .B(m[14]), .Z(n4775) );
  AND U8296 ( .A(n5961), .B(n5962), .Z(n5960) );
  NAND U8297 ( .A(o[14]), .B(n5916), .Z(n5962) );
  NANDN U8298 ( .A(n5917), .B(creg[14]), .Z(n5961) );
  NAND U8299 ( .A(n5963), .B(n4753), .Z(n3586) );
  NANDN U8300 ( .A(init), .B(m[15]), .Z(n4753) );
  AND U8301 ( .A(n5964), .B(n5965), .Z(n5963) );
  NAND U8302 ( .A(o[15]), .B(n5916), .Z(n5965) );
  NANDN U8303 ( .A(n5917), .B(creg[15]), .Z(n5964) );
  NAND U8304 ( .A(n5966), .B(n4731), .Z(n3585) );
  NANDN U8305 ( .A(init), .B(m[16]), .Z(n4731) );
  AND U8306 ( .A(n5967), .B(n5968), .Z(n5966) );
  NAND U8307 ( .A(o[16]), .B(n5916), .Z(n5968) );
  NANDN U8308 ( .A(n5917), .B(creg[16]), .Z(n5967) );
  NAND U8309 ( .A(n5969), .B(n4709), .Z(n3584) );
  NANDN U8310 ( .A(init), .B(m[17]), .Z(n4709) );
  AND U8311 ( .A(n5970), .B(n5971), .Z(n5969) );
  NAND U8312 ( .A(o[17]), .B(n5916), .Z(n5971) );
  NANDN U8313 ( .A(n5917), .B(creg[17]), .Z(n5970) );
  NAND U8314 ( .A(n5972), .B(n4687), .Z(n3583) );
  NANDN U8315 ( .A(init), .B(m[18]), .Z(n4687) );
  AND U8316 ( .A(n5973), .B(n5974), .Z(n5972) );
  NAND U8317 ( .A(o[18]), .B(n5916), .Z(n5974) );
  NANDN U8318 ( .A(n5917), .B(creg[18]), .Z(n5973) );
  NAND U8319 ( .A(n5975), .B(n4665), .Z(n3582) );
  NANDN U8320 ( .A(init), .B(m[19]), .Z(n4665) );
  AND U8321 ( .A(n5976), .B(n5977), .Z(n5975) );
  NAND U8322 ( .A(o[19]), .B(n5916), .Z(n5977) );
  NANDN U8323 ( .A(n5917), .B(creg[19]), .Z(n5976) );
  NAND U8324 ( .A(n5978), .B(n4641), .Z(n3581) );
  NANDN U8325 ( .A(init), .B(m[20]), .Z(n4641) );
  AND U8326 ( .A(n5979), .B(n5980), .Z(n5978) );
  NAND U8327 ( .A(o[20]), .B(n5916), .Z(n5980) );
  NANDN U8328 ( .A(n5917), .B(creg[20]), .Z(n5979) );
  NAND U8329 ( .A(n5981), .B(n4619), .Z(n3580) );
  NANDN U8330 ( .A(init), .B(m[21]), .Z(n4619) );
  AND U8331 ( .A(n5982), .B(n5983), .Z(n5981) );
  NAND U8332 ( .A(o[21]), .B(n5916), .Z(n5983) );
  NANDN U8333 ( .A(n5917), .B(creg[21]), .Z(n5982) );
  NAND U8334 ( .A(n5984), .B(n4597), .Z(n3579) );
  NANDN U8335 ( .A(init), .B(m[22]), .Z(n4597) );
  AND U8336 ( .A(n5985), .B(n5986), .Z(n5984) );
  NAND U8337 ( .A(o[22]), .B(n5916), .Z(n5986) );
  NANDN U8338 ( .A(n5917), .B(creg[22]), .Z(n5985) );
  NAND U8339 ( .A(n5987), .B(n4575), .Z(n3578) );
  NANDN U8340 ( .A(init), .B(m[23]), .Z(n4575) );
  AND U8341 ( .A(n5988), .B(n5989), .Z(n5987) );
  NAND U8342 ( .A(o[23]), .B(n5916), .Z(n5989) );
  NANDN U8343 ( .A(n5917), .B(creg[23]), .Z(n5988) );
  NAND U8344 ( .A(n5990), .B(n4553), .Z(n3577) );
  NANDN U8345 ( .A(init), .B(m[24]), .Z(n4553) );
  AND U8346 ( .A(n5991), .B(n5992), .Z(n5990) );
  NAND U8347 ( .A(o[24]), .B(n5916), .Z(n5992) );
  NANDN U8348 ( .A(n5917), .B(creg[24]), .Z(n5991) );
  NAND U8349 ( .A(n5993), .B(n4539), .Z(n3576) );
  NANDN U8350 ( .A(init), .B(m[25]), .Z(n4539) );
  AND U8351 ( .A(n5994), .B(n5995), .Z(n5993) );
  NAND U8352 ( .A(o[25]), .B(n5916), .Z(n5995) );
  NANDN U8353 ( .A(n5917), .B(creg[25]), .Z(n5994) );
  NAND U8354 ( .A(n5996), .B(n4537), .Z(n3575) );
  NANDN U8355 ( .A(init), .B(m[26]), .Z(n4537) );
  AND U8356 ( .A(n5997), .B(n5998), .Z(n5996) );
  NAND U8357 ( .A(o[26]), .B(n5916), .Z(n5998) );
  NANDN U8358 ( .A(n5917), .B(creg[26]), .Z(n5997) );
  NAND U8359 ( .A(n5999), .B(n4535), .Z(n3574) );
  NANDN U8360 ( .A(init), .B(m[27]), .Z(n4535) );
  AND U8361 ( .A(n6000), .B(n6001), .Z(n5999) );
  NAND U8362 ( .A(o[27]), .B(n5916), .Z(n6001) );
  NANDN U8363 ( .A(n5917), .B(creg[27]), .Z(n6000) );
  NAND U8364 ( .A(n6002), .B(n4533), .Z(n3573) );
  NANDN U8365 ( .A(init), .B(m[28]), .Z(n4533) );
  AND U8366 ( .A(n6003), .B(n6004), .Z(n6002) );
  NAND U8367 ( .A(o[28]), .B(n5916), .Z(n6004) );
  NANDN U8368 ( .A(n5917), .B(creg[28]), .Z(n6003) );
  NAND U8369 ( .A(n6005), .B(n4531), .Z(n3572) );
  NANDN U8370 ( .A(init), .B(m[29]), .Z(n4531) );
  AND U8371 ( .A(n6006), .B(n6007), .Z(n6005) );
  NAND U8372 ( .A(o[29]), .B(n5916), .Z(n6007) );
  NANDN U8373 ( .A(n5917), .B(creg[29]), .Z(n6006) );
  NAND U8374 ( .A(n6008), .B(n4527), .Z(n3571) );
  NANDN U8375 ( .A(init), .B(m[30]), .Z(n4527) );
  AND U8376 ( .A(n6009), .B(n6010), .Z(n6008) );
  NAND U8377 ( .A(o[30]), .B(n5916), .Z(n6010) );
  NANDN U8378 ( .A(n5917), .B(creg[30]), .Z(n6009) );
  NAND U8379 ( .A(n6011), .B(n4525), .Z(n3570) );
  NANDN U8380 ( .A(init), .B(m[31]), .Z(n4525) );
  AND U8381 ( .A(n6012), .B(n6013), .Z(n6011) );
  NAND U8382 ( .A(o[31]), .B(n5916), .Z(n6013) );
  NANDN U8383 ( .A(n5917), .B(creg[31]), .Z(n6012) );
  NAND U8384 ( .A(n6014), .B(n4523), .Z(n3569) );
  NANDN U8385 ( .A(init), .B(m[32]), .Z(n4523) );
  AND U8386 ( .A(n6015), .B(n6016), .Z(n6014) );
  NAND U8387 ( .A(o[32]), .B(n5916), .Z(n6016) );
  NANDN U8388 ( .A(n5917), .B(creg[32]), .Z(n6015) );
  NAND U8389 ( .A(n6017), .B(n4521), .Z(n3568) );
  NANDN U8390 ( .A(init), .B(m[33]), .Z(n4521) );
  AND U8391 ( .A(n6018), .B(n6019), .Z(n6017) );
  NAND U8392 ( .A(o[33]), .B(n5916), .Z(n6019) );
  NANDN U8393 ( .A(n5917), .B(creg[33]), .Z(n6018) );
  NAND U8394 ( .A(n6020), .B(n4519), .Z(n3567) );
  NANDN U8395 ( .A(init), .B(m[34]), .Z(n4519) );
  AND U8396 ( .A(n6021), .B(n6022), .Z(n6020) );
  NAND U8397 ( .A(o[34]), .B(n5916), .Z(n6022) );
  NANDN U8398 ( .A(n5917), .B(creg[34]), .Z(n6021) );
  NAND U8399 ( .A(n6023), .B(n4517), .Z(n3566) );
  NANDN U8400 ( .A(init), .B(m[35]), .Z(n4517) );
  AND U8401 ( .A(n6024), .B(n6025), .Z(n6023) );
  NAND U8402 ( .A(o[35]), .B(n5916), .Z(n6025) );
  NANDN U8403 ( .A(n5917), .B(creg[35]), .Z(n6024) );
  NAND U8404 ( .A(n6026), .B(n4515), .Z(n3565) );
  NANDN U8405 ( .A(init), .B(m[36]), .Z(n4515) );
  AND U8406 ( .A(n6027), .B(n6028), .Z(n6026) );
  NAND U8407 ( .A(o[36]), .B(n5916), .Z(n6028) );
  NANDN U8408 ( .A(n5917), .B(creg[36]), .Z(n6027) );
  NAND U8409 ( .A(n6029), .B(n4513), .Z(n3564) );
  NANDN U8410 ( .A(init), .B(m[37]), .Z(n4513) );
  AND U8411 ( .A(n6030), .B(n6031), .Z(n6029) );
  NAND U8412 ( .A(o[37]), .B(n5916), .Z(n6031) );
  NANDN U8413 ( .A(n5917), .B(creg[37]), .Z(n6030) );
  NAND U8414 ( .A(n6032), .B(n4511), .Z(n3563) );
  NANDN U8415 ( .A(init), .B(m[38]), .Z(n4511) );
  AND U8416 ( .A(n6033), .B(n6034), .Z(n6032) );
  NAND U8417 ( .A(o[38]), .B(n5916), .Z(n6034) );
  NANDN U8418 ( .A(n5917), .B(creg[38]), .Z(n6033) );
  NAND U8419 ( .A(n6035), .B(n4509), .Z(n3562) );
  NANDN U8420 ( .A(init), .B(m[39]), .Z(n4509) );
  AND U8421 ( .A(n6036), .B(n6037), .Z(n6035) );
  NAND U8422 ( .A(o[39]), .B(n5916), .Z(n6037) );
  NANDN U8423 ( .A(n5917), .B(creg[39]), .Z(n6036) );
  NAND U8424 ( .A(n6038), .B(n4505), .Z(n3561) );
  NANDN U8425 ( .A(init), .B(m[40]), .Z(n4505) );
  AND U8426 ( .A(n6039), .B(n6040), .Z(n6038) );
  NAND U8427 ( .A(o[40]), .B(n5916), .Z(n6040) );
  NANDN U8428 ( .A(n5917), .B(creg[40]), .Z(n6039) );
  NAND U8429 ( .A(n6041), .B(n4503), .Z(n3560) );
  NANDN U8430 ( .A(init), .B(m[41]), .Z(n4503) );
  AND U8431 ( .A(n6042), .B(n6043), .Z(n6041) );
  NAND U8432 ( .A(o[41]), .B(n5916), .Z(n6043) );
  NANDN U8433 ( .A(n5917), .B(creg[41]), .Z(n6042) );
  NAND U8434 ( .A(n6044), .B(n4501), .Z(n3559) );
  NANDN U8435 ( .A(init), .B(m[42]), .Z(n4501) );
  AND U8436 ( .A(n6045), .B(n6046), .Z(n6044) );
  NAND U8437 ( .A(o[42]), .B(n5916), .Z(n6046) );
  NANDN U8438 ( .A(n5917), .B(creg[42]), .Z(n6045) );
  NAND U8439 ( .A(n6047), .B(n4499), .Z(n3558) );
  NANDN U8440 ( .A(init), .B(m[43]), .Z(n4499) );
  AND U8441 ( .A(n6048), .B(n6049), .Z(n6047) );
  NAND U8442 ( .A(o[43]), .B(n5916), .Z(n6049) );
  NANDN U8443 ( .A(n5917), .B(creg[43]), .Z(n6048) );
  NAND U8444 ( .A(n6050), .B(n4497), .Z(n3557) );
  NANDN U8445 ( .A(init), .B(m[44]), .Z(n4497) );
  AND U8446 ( .A(n6051), .B(n6052), .Z(n6050) );
  NAND U8447 ( .A(o[44]), .B(n5916), .Z(n6052) );
  NANDN U8448 ( .A(n5917), .B(creg[44]), .Z(n6051) );
  NAND U8449 ( .A(n6053), .B(n4495), .Z(n3556) );
  NANDN U8450 ( .A(init), .B(m[45]), .Z(n4495) );
  AND U8451 ( .A(n6054), .B(n6055), .Z(n6053) );
  NAND U8452 ( .A(o[45]), .B(n5916), .Z(n6055) );
  NANDN U8453 ( .A(n5917), .B(creg[45]), .Z(n6054) );
  NAND U8454 ( .A(n6056), .B(n4493), .Z(n3555) );
  NANDN U8455 ( .A(init), .B(m[46]), .Z(n4493) );
  AND U8456 ( .A(n6057), .B(n6058), .Z(n6056) );
  NAND U8457 ( .A(o[46]), .B(n5916), .Z(n6058) );
  NANDN U8458 ( .A(n5917), .B(creg[46]), .Z(n6057) );
  NAND U8459 ( .A(n6059), .B(n4491), .Z(n3554) );
  NANDN U8460 ( .A(init), .B(m[47]), .Z(n4491) );
  AND U8461 ( .A(n6060), .B(n6061), .Z(n6059) );
  NAND U8462 ( .A(o[47]), .B(n5916), .Z(n6061) );
  NANDN U8463 ( .A(n5917), .B(creg[47]), .Z(n6060) );
  NAND U8464 ( .A(n6062), .B(n4489), .Z(n3553) );
  NANDN U8465 ( .A(init), .B(m[48]), .Z(n4489) );
  AND U8466 ( .A(n6063), .B(n6064), .Z(n6062) );
  NAND U8467 ( .A(o[48]), .B(n5916), .Z(n6064) );
  NANDN U8468 ( .A(n5917), .B(creg[48]), .Z(n6063) );
  NAND U8469 ( .A(n6065), .B(n4487), .Z(n3552) );
  NANDN U8470 ( .A(init), .B(m[49]), .Z(n4487) );
  AND U8471 ( .A(n6066), .B(n6067), .Z(n6065) );
  NAND U8472 ( .A(o[49]), .B(n5916), .Z(n6067) );
  NANDN U8473 ( .A(n5917), .B(creg[49]), .Z(n6066) );
  NAND U8474 ( .A(n6068), .B(n4483), .Z(n3551) );
  NANDN U8475 ( .A(init), .B(m[50]), .Z(n4483) );
  AND U8476 ( .A(n6069), .B(n6070), .Z(n6068) );
  NAND U8477 ( .A(o[50]), .B(n5916), .Z(n6070) );
  NANDN U8478 ( .A(n5917), .B(creg[50]), .Z(n6069) );
  NAND U8479 ( .A(n6071), .B(n4481), .Z(n3550) );
  NANDN U8480 ( .A(init), .B(m[51]), .Z(n4481) );
  AND U8481 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U8482 ( .A(o[51]), .B(n5916), .Z(n6073) );
  NANDN U8483 ( .A(n5917), .B(creg[51]), .Z(n6072) );
  NAND U8484 ( .A(n6074), .B(n4479), .Z(n3549) );
  NANDN U8485 ( .A(init), .B(m[52]), .Z(n4479) );
  AND U8486 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U8487 ( .A(o[52]), .B(n5916), .Z(n6076) );
  NANDN U8488 ( .A(n5917), .B(creg[52]), .Z(n6075) );
  NAND U8489 ( .A(n6077), .B(n4477), .Z(n3548) );
  NANDN U8490 ( .A(init), .B(m[53]), .Z(n4477) );
  AND U8491 ( .A(n6078), .B(n6079), .Z(n6077) );
  NAND U8492 ( .A(o[53]), .B(n5916), .Z(n6079) );
  NANDN U8493 ( .A(n5917), .B(creg[53]), .Z(n6078) );
  NAND U8494 ( .A(n6080), .B(n4475), .Z(n3547) );
  NANDN U8495 ( .A(init), .B(m[54]), .Z(n4475) );
  AND U8496 ( .A(n6081), .B(n6082), .Z(n6080) );
  NAND U8497 ( .A(o[54]), .B(n5916), .Z(n6082) );
  NANDN U8498 ( .A(n5917), .B(creg[54]), .Z(n6081) );
  NAND U8499 ( .A(n6083), .B(n4473), .Z(n3546) );
  NANDN U8500 ( .A(init), .B(m[55]), .Z(n4473) );
  AND U8501 ( .A(n6084), .B(n6085), .Z(n6083) );
  NAND U8502 ( .A(o[55]), .B(n5916), .Z(n6085) );
  NANDN U8503 ( .A(n5917), .B(creg[55]), .Z(n6084) );
  NAND U8504 ( .A(n6086), .B(n4471), .Z(n3545) );
  NANDN U8505 ( .A(init), .B(m[56]), .Z(n4471) );
  AND U8506 ( .A(n6087), .B(n6088), .Z(n6086) );
  NAND U8507 ( .A(o[56]), .B(n5916), .Z(n6088) );
  NANDN U8508 ( .A(n5917), .B(creg[56]), .Z(n6087) );
  NAND U8509 ( .A(n6089), .B(n4469), .Z(n3544) );
  NANDN U8510 ( .A(init), .B(m[57]), .Z(n4469) );
  AND U8511 ( .A(n6090), .B(n6091), .Z(n6089) );
  NAND U8512 ( .A(o[57]), .B(n5916), .Z(n6091) );
  NANDN U8513 ( .A(n5917), .B(creg[57]), .Z(n6090) );
  NAND U8514 ( .A(n6092), .B(n4467), .Z(n3543) );
  NANDN U8515 ( .A(init), .B(m[58]), .Z(n4467) );
  AND U8516 ( .A(n6093), .B(n6094), .Z(n6092) );
  NAND U8517 ( .A(o[58]), .B(n5916), .Z(n6094) );
  NANDN U8518 ( .A(n5917), .B(creg[58]), .Z(n6093) );
  NAND U8519 ( .A(n6095), .B(n4465), .Z(n3542) );
  NANDN U8520 ( .A(init), .B(m[59]), .Z(n4465) );
  AND U8521 ( .A(n6096), .B(n6097), .Z(n6095) );
  NAND U8522 ( .A(o[59]), .B(n5916), .Z(n6097) );
  NANDN U8523 ( .A(n5917), .B(creg[59]), .Z(n6096) );
  NAND U8524 ( .A(n6098), .B(n4461), .Z(n3541) );
  NANDN U8525 ( .A(init), .B(m[60]), .Z(n4461) );
  AND U8526 ( .A(n6099), .B(n6100), .Z(n6098) );
  NAND U8527 ( .A(o[60]), .B(n5916), .Z(n6100) );
  NANDN U8528 ( .A(n5917), .B(creg[60]), .Z(n6099) );
  NAND U8529 ( .A(n6101), .B(n4459), .Z(n3540) );
  NANDN U8530 ( .A(init), .B(m[61]), .Z(n4459) );
  AND U8531 ( .A(n6102), .B(n6103), .Z(n6101) );
  NAND U8532 ( .A(o[61]), .B(n5916), .Z(n6103) );
  NANDN U8533 ( .A(n5917), .B(creg[61]), .Z(n6102) );
  NAND U8534 ( .A(n6104), .B(n4457), .Z(n3539) );
  NANDN U8535 ( .A(init), .B(m[62]), .Z(n4457) );
  AND U8536 ( .A(n6105), .B(n6106), .Z(n6104) );
  NAND U8537 ( .A(o[62]), .B(n5916), .Z(n6106) );
  NANDN U8538 ( .A(n5917), .B(creg[62]), .Z(n6105) );
  NAND U8539 ( .A(n6107), .B(n4455), .Z(n3538) );
  NANDN U8540 ( .A(init), .B(m[63]), .Z(n4455) );
  AND U8541 ( .A(n6108), .B(n6109), .Z(n6107) );
  NAND U8542 ( .A(o[63]), .B(n5916), .Z(n6109) );
  NANDN U8543 ( .A(n5917), .B(creg[63]), .Z(n6108) );
  NAND U8544 ( .A(n6110), .B(n4453), .Z(n3537) );
  NANDN U8545 ( .A(init), .B(m[64]), .Z(n4453) );
  AND U8546 ( .A(n6111), .B(n6112), .Z(n6110) );
  NAND U8547 ( .A(o[64]), .B(n5916), .Z(n6112) );
  NANDN U8548 ( .A(n5917), .B(creg[64]), .Z(n6111) );
  NAND U8549 ( .A(n6113), .B(n4451), .Z(n3536) );
  NANDN U8550 ( .A(init), .B(m[65]), .Z(n4451) );
  AND U8551 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U8552 ( .A(o[65]), .B(n5916), .Z(n6115) );
  NANDN U8553 ( .A(n5917), .B(creg[65]), .Z(n6114) );
  NAND U8554 ( .A(n6116), .B(n4449), .Z(n3535) );
  NANDN U8555 ( .A(init), .B(m[66]), .Z(n4449) );
  AND U8556 ( .A(n6117), .B(n6118), .Z(n6116) );
  NAND U8557 ( .A(o[66]), .B(n5916), .Z(n6118) );
  NANDN U8558 ( .A(n5917), .B(creg[66]), .Z(n6117) );
  NAND U8559 ( .A(n6119), .B(n4447), .Z(n3534) );
  NANDN U8560 ( .A(init), .B(m[67]), .Z(n4447) );
  AND U8561 ( .A(n6120), .B(n6121), .Z(n6119) );
  NAND U8562 ( .A(o[67]), .B(n5916), .Z(n6121) );
  NANDN U8563 ( .A(n5917), .B(creg[67]), .Z(n6120) );
  NAND U8564 ( .A(n6122), .B(n4445), .Z(n3533) );
  NANDN U8565 ( .A(init), .B(m[68]), .Z(n4445) );
  AND U8566 ( .A(n6123), .B(n6124), .Z(n6122) );
  NAND U8567 ( .A(o[68]), .B(n5916), .Z(n6124) );
  NANDN U8568 ( .A(n5917), .B(creg[68]), .Z(n6123) );
  NAND U8569 ( .A(n6125), .B(n4443), .Z(n3532) );
  NANDN U8570 ( .A(init), .B(m[69]), .Z(n4443) );
  AND U8571 ( .A(n6126), .B(n6127), .Z(n6125) );
  NAND U8572 ( .A(o[69]), .B(n5916), .Z(n6127) );
  NANDN U8573 ( .A(n5917), .B(creg[69]), .Z(n6126) );
  NAND U8574 ( .A(n6128), .B(n4439), .Z(n3531) );
  NANDN U8575 ( .A(init), .B(m[70]), .Z(n4439) );
  AND U8576 ( .A(n6129), .B(n6130), .Z(n6128) );
  NAND U8577 ( .A(o[70]), .B(n5916), .Z(n6130) );
  NANDN U8578 ( .A(n5917), .B(creg[70]), .Z(n6129) );
  NAND U8579 ( .A(n6131), .B(n4437), .Z(n3530) );
  NANDN U8580 ( .A(init), .B(m[71]), .Z(n4437) );
  AND U8581 ( .A(n6132), .B(n6133), .Z(n6131) );
  NAND U8582 ( .A(o[71]), .B(n5916), .Z(n6133) );
  NANDN U8583 ( .A(n5917), .B(creg[71]), .Z(n6132) );
  NAND U8584 ( .A(n6134), .B(n4435), .Z(n3529) );
  NANDN U8585 ( .A(init), .B(m[72]), .Z(n4435) );
  AND U8586 ( .A(n6135), .B(n6136), .Z(n6134) );
  NAND U8587 ( .A(o[72]), .B(n5916), .Z(n6136) );
  NANDN U8588 ( .A(n5917), .B(creg[72]), .Z(n6135) );
  NAND U8589 ( .A(n6137), .B(n4433), .Z(n3528) );
  NANDN U8590 ( .A(init), .B(m[73]), .Z(n4433) );
  AND U8591 ( .A(n6138), .B(n6139), .Z(n6137) );
  NAND U8592 ( .A(o[73]), .B(n5916), .Z(n6139) );
  NANDN U8593 ( .A(n5917), .B(creg[73]), .Z(n6138) );
  NAND U8594 ( .A(n6140), .B(n4431), .Z(n3527) );
  NANDN U8595 ( .A(init), .B(m[74]), .Z(n4431) );
  AND U8596 ( .A(n6141), .B(n6142), .Z(n6140) );
  NAND U8597 ( .A(o[74]), .B(n5916), .Z(n6142) );
  NANDN U8598 ( .A(n5917), .B(creg[74]), .Z(n6141) );
  NAND U8599 ( .A(n6143), .B(n4429), .Z(n3526) );
  NANDN U8600 ( .A(init), .B(m[75]), .Z(n4429) );
  AND U8601 ( .A(n6144), .B(n6145), .Z(n6143) );
  NAND U8602 ( .A(o[75]), .B(n5916), .Z(n6145) );
  NANDN U8603 ( .A(n5917), .B(creg[75]), .Z(n6144) );
  NAND U8604 ( .A(n6146), .B(n4427), .Z(n3525) );
  NANDN U8605 ( .A(init), .B(m[76]), .Z(n4427) );
  AND U8606 ( .A(n6147), .B(n6148), .Z(n6146) );
  NAND U8607 ( .A(o[76]), .B(n5916), .Z(n6148) );
  NANDN U8608 ( .A(n5917), .B(creg[76]), .Z(n6147) );
  NAND U8609 ( .A(n6149), .B(n4425), .Z(n3524) );
  NANDN U8610 ( .A(init), .B(m[77]), .Z(n4425) );
  AND U8611 ( .A(n6150), .B(n6151), .Z(n6149) );
  NAND U8612 ( .A(o[77]), .B(n5916), .Z(n6151) );
  NANDN U8613 ( .A(n5917), .B(creg[77]), .Z(n6150) );
  NAND U8614 ( .A(n6152), .B(n4423), .Z(n3523) );
  NANDN U8615 ( .A(init), .B(m[78]), .Z(n4423) );
  AND U8616 ( .A(n6153), .B(n6154), .Z(n6152) );
  NAND U8617 ( .A(o[78]), .B(n5916), .Z(n6154) );
  NANDN U8618 ( .A(n5917), .B(creg[78]), .Z(n6153) );
  NAND U8619 ( .A(n6155), .B(n4421), .Z(n3522) );
  NANDN U8620 ( .A(init), .B(m[79]), .Z(n4421) );
  AND U8621 ( .A(n6156), .B(n6157), .Z(n6155) );
  NAND U8622 ( .A(o[79]), .B(n5916), .Z(n6157) );
  NANDN U8623 ( .A(n5917), .B(creg[79]), .Z(n6156) );
  NAND U8624 ( .A(n6158), .B(n4417), .Z(n3521) );
  NANDN U8625 ( .A(init), .B(m[80]), .Z(n4417) );
  AND U8626 ( .A(n6159), .B(n6160), .Z(n6158) );
  NAND U8627 ( .A(o[80]), .B(n5916), .Z(n6160) );
  NANDN U8628 ( .A(n5917), .B(creg[80]), .Z(n6159) );
  NAND U8629 ( .A(n6161), .B(n4415), .Z(n3520) );
  NANDN U8630 ( .A(init), .B(m[81]), .Z(n4415) );
  AND U8631 ( .A(n6162), .B(n6163), .Z(n6161) );
  NAND U8632 ( .A(o[81]), .B(n5916), .Z(n6163) );
  NANDN U8633 ( .A(n5917), .B(creg[81]), .Z(n6162) );
  NAND U8634 ( .A(n6164), .B(n4413), .Z(n3519) );
  NANDN U8635 ( .A(init), .B(m[82]), .Z(n4413) );
  AND U8636 ( .A(n6165), .B(n6166), .Z(n6164) );
  NAND U8637 ( .A(o[82]), .B(n5916), .Z(n6166) );
  NANDN U8638 ( .A(n5917), .B(creg[82]), .Z(n6165) );
  NAND U8639 ( .A(n6167), .B(n4411), .Z(n3518) );
  NANDN U8640 ( .A(init), .B(m[83]), .Z(n4411) );
  AND U8641 ( .A(n6168), .B(n6169), .Z(n6167) );
  NAND U8642 ( .A(o[83]), .B(n5916), .Z(n6169) );
  NANDN U8643 ( .A(n5917), .B(creg[83]), .Z(n6168) );
  NAND U8644 ( .A(n6170), .B(n4409), .Z(n3517) );
  NANDN U8645 ( .A(init), .B(m[84]), .Z(n4409) );
  AND U8646 ( .A(n6171), .B(n6172), .Z(n6170) );
  NAND U8647 ( .A(o[84]), .B(n5916), .Z(n6172) );
  NANDN U8648 ( .A(n5917), .B(creg[84]), .Z(n6171) );
  NAND U8649 ( .A(n6173), .B(n4407), .Z(n3516) );
  NANDN U8650 ( .A(init), .B(m[85]), .Z(n4407) );
  AND U8651 ( .A(n6174), .B(n6175), .Z(n6173) );
  NAND U8652 ( .A(o[85]), .B(n5916), .Z(n6175) );
  NANDN U8653 ( .A(n5917), .B(creg[85]), .Z(n6174) );
  NAND U8654 ( .A(n6176), .B(n4405), .Z(n3515) );
  NANDN U8655 ( .A(init), .B(m[86]), .Z(n4405) );
  AND U8656 ( .A(n6177), .B(n6178), .Z(n6176) );
  NAND U8657 ( .A(o[86]), .B(n5916), .Z(n6178) );
  NANDN U8658 ( .A(n5917), .B(creg[86]), .Z(n6177) );
  NAND U8659 ( .A(n6179), .B(n4403), .Z(n3514) );
  NANDN U8660 ( .A(init), .B(m[87]), .Z(n4403) );
  AND U8661 ( .A(n6180), .B(n6181), .Z(n6179) );
  NAND U8662 ( .A(o[87]), .B(n5916), .Z(n6181) );
  NANDN U8663 ( .A(n5917), .B(creg[87]), .Z(n6180) );
  NAND U8664 ( .A(n6182), .B(n4401), .Z(n3513) );
  NANDN U8665 ( .A(init), .B(m[88]), .Z(n4401) );
  AND U8666 ( .A(n6183), .B(n6184), .Z(n6182) );
  NAND U8667 ( .A(o[88]), .B(n5916), .Z(n6184) );
  NANDN U8668 ( .A(n5917), .B(creg[88]), .Z(n6183) );
  NAND U8669 ( .A(n6185), .B(n4399), .Z(n3512) );
  NANDN U8670 ( .A(init), .B(m[89]), .Z(n4399) );
  AND U8671 ( .A(n6186), .B(n6187), .Z(n6185) );
  NAND U8672 ( .A(o[89]), .B(n5916), .Z(n6187) );
  NANDN U8673 ( .A(n5917), .B(creg[89]), .Z(n6186) );
  NAND U8674 ( .A(n6188), .B(n4395), .Z(n3511) );
  NANDN U8675 ( .A(init), .B(m[90]), .Z(n4395) );
  AND U8676 ( .A(n6189), .B(n6190), .Z(n6188) );
  NAND U8677 ( .A(o[90]), .B(n5916), .Z(n6190) );
  NANDN U8678 ( .A(n5917), .B(creg[90]), .Z(n6189) );
  NAND U8679 ( .A(n6191), .B(n4393), .Z(n3510) );
  NANDN U8680 ( .A(init), .B(m[91]), .Z(n4393) );
  AND U8681 ( .A(n6192), .B(n6193), .Z(n6191) );
  NAND U8682 ( .A(o[91]), .B(n5916), .Z(n6193) );
  NANDN U8683 ( .A(n5917), .B(creg[91]), .Z(n6192) );
  NAND U8684 ( .A(n6194), .B(n4391), .Z(n3509) );
  NANDN U8685 ( .A(init), .B(m[92]), .Z(n4391) );
  AND U8686 ( .A(n6195), .B(n6196), .Z(n6194) );
  NAND U8687 ( .A(o[92]), .B(n5916), .Z(n6196) );
  NANDN U8688 ( .A(n5917), .B(creg[92]), .Z(n6195) );
  NAND U8689 ( .A(n6197), .B(n4389), .Z(n3508) );
  NANDN U8690 ( .A(init), .B(m[93]), .Z(n4389) );
  AND U8691 ( .A(n6198), .B(n6199), .Z(n6197) );
  NAND U8692 ( .A(o[93]), .B(n5916), .Z(n6199) );
  NANDN U8693 ( .A(n5917), .B(creg[93]), .Z(n6198) );
  NAND U8694 ( .A(n6200), .B(n4387), .Z(n3507) );
  NANDN U8695 ( .A(init), .B(m[94]), .Z(n4387) );
  AND U8696 ( .A(n6201), .B(n6202), .Z(n6200) );
  NAND U8697 ( .A(o[94]), .B(n5916), .Z(n6202) );
  NANDN U8698 ( .A(n5917), .B(creg[94]), .Z(n6201) );
  NAND U8699 ( .A(n6203), .B(n4385), .Z(n3506) );
  NANDN U8700 ( .A(init), .B(m[95]), .Z(n4385) );
  AND U8701 ( .A(n6204), .B(n6205), .Z(n6203) );
  NAND U8702 ( .A(o[95]), .B(n5916), .Z(n6205) );
  NANDN U8703 ( .A(n5917), .B(creg[95]), .Z(n6204) );
  NAND U8704 ( .A(n6206), .B(n4383), .Z(n3505) );
  NANDN U8705 ( .A(init), .B(m[96]), .Z(n4383) );
  AND U8706 ( .A(n6207), .B(n6208), .Z(n6206) );
  NAND U8707 ( .A(o[96]), .B(n5916), .Z(n6208) );
  NANDN U8708 ( .A(n5917), .B(creg[96]), .Z(n6207) );
  NAND U8709 ( .A(n6209), .B(n4381), .Z(n3504) );
  NANDN U8710 ( .A(init), .B(m[97]), .Z(n4381) );
  AND U8711 ( .A(n6210), .B(n6211), .Z(n6209) );
  NAND U8712 ( .A(o[97]), .B(n5916), .Z(n6211) );
  NANDN U8713 ( .A(n5917), .B(creg[97]), .Z(n6210) );
  NAND U8714 ( .A(n6212), .B(n4379), .Z(n3503) );
  NANDN U8715 ( .A(init), .B(m[98]), .Z(n4379) );
  AND U8716 ( .A(n6213), .B(n6214), .Z(n6212) );
  NAND U8717 ( .A(o[98]), .B(n5916), .Z(n6214) );
  NANDN U8718 ( .A(n5917), .B(creg[98]), .Z(n6213) );
  NAND U8719 ( .A(n6215), .B(n4377), .Z(n3502) );
  NANDN U8720 ( .A(init), .B(m[99]), .Z(n4377) );
  AND U8721 ( .A(n6216), .B(n6217), .Z(n6215) );
  NAND U8722 ( .A(o[99]), .B(n5916), .Z(n6217) );
  NANDN U8723 ( .A(n5917), .B(creg[99]), .Z(n6216) );
  NAND U8724 ( .A(n6218), .B(n4883), .Z(n3501) );
  NANDN U8725 ( .A(init), .B(m[100]), .Z(n4883) );
  AND U8726 ( .A(n6219), .B(n6220), .Z(n6218) );
  NAND U8727 ( .A(o[100]), .B(n5916), .Z(n6220) );
  NANDN U8728 ( .A(n5917), .B(creg[100]), .Z(n6219) );
  NAND U8729 ( .A(n6221), .B(n4881), .Z(n3500) );
  NANDN U8730 ( .A(init), .B(m[101]), .Z(n4881) );
  AND U8731 ( .A(n6222), .B(n6223), .Z(n6221) );
  NAND U8732 ( .A(o[101]), .B(n5916), .Z(n6223) );
  NANDN U8733 ( .A(n5917), .B(creg[101]), .Z(n6222) );
  NAND U8734 ( .A(n6224), .B(n4879), .Z(n3499) );
  NANDN U8735 ( .A(init), .B(m[102]), .Z(n4879) );
  AND U8736 ( .A(n6225), .B(n6226), .Z(n6224) );
  NAND U8737 ( .A(o[102]), .B(n5916), .Z(n6226) );
  NANDN U8738 ( .A(n5917), .B(creg[102]), .Z(n6225) );
  NAND U8739 ( .A(n6227), .B(n4877), .Z(n3498) );
  NANDN U8740 ( .A(init), .B(m[103]), .Z(n4877) );
  AND U8741 ( .A(n6228), .B(n6229), .Z(n6227) );
  NAND U8742 ( .A(o[103]), .B(n5916), .Z(n6229) );
  NANDN U8743 ( .A(n5917), .B(creg[103]), .Z(n6228) );
  NAND U8744 ( .A(n6230), .B(n4875), .Z(n3497) );
  NANDN U8745 ( .A(init), .B(m[104]), .Z(n4875) );
  AND U8746 ( .A(n6231), .B(n6232), .Z(n6230) );
  NAND U8747 ( .A(o[104]), .B(n5916), .Z(n6232) );
  NANDN U8748 ( .A(n5917), .B(creg[104]), .Z(n6231) );
  NAND U8749 ( .A(n6233), .B(n4873), .Z(n3496) );
  NANDN U8750 ( .A(init), .B(m[105]), .Z(n4873) );
  AND U8751 ( .A(n6234), .B(n6235), .Z(n6233) );
  NAND U8752 ( .A(o[105]), .B(n5916), .Z(n6235) );
  NANDN U8753 ( .A(n5917), .B(creg[105]), .Z(n6234) );
  NAND U8754 ( .A(n6236), .B(n4871), .Z(n3495) );
  NANDN U8755 ( .A(init), .B(m[106]), .Z(n4871) );
  AND U8756 ( .A(n6237), .B(n6238), .Z(n6236) );
  NAND U8757 ( .A(o[106]), .B(n5916), .Z(n6238) );
  NANDN U8758 ( .A(n5917), .B(creg[106]), .Z(n6237) );
  NAND U8759 ( .A(n6239), .B(n4869), .Z(n3494) );
  NANDN U8760 ( .A(init), .B(m[107]), .Z(n4869) );
  AND U8761 ( .A(n6240), .B(n6241), .Z(n6239) );
  NAND U8762 ( .A(o[107]), .B(n5916), .Z(n6241) );
  NANDN U8763 ( .A(n5917), .B(creg[107]), .Z(n6240) );
  NAND U8764 ( .A(n6242), .B(n4867), .Z(n3493) );
  NANDN U8765 ( .A(init), .B(m[108]), .Z(n4867) );
  AND U8766 ( .A(n6243), .B(n6244), .Z(n6242) );
  NAND U8767 ( .A(o[108]), .B(n5916), .Z(n6244) );
  NANDN U8768 ( .A(n5917), .B(creg[108]), .Z(n6243) );
  NAND U8769 ( .A(n6245), .B(n4865), .Z(n3492) );
  NANDN U8770 ( .A(init), .B(m[109]), .Z(n4865) );
  AND U8771 ( .A(n6246), .B(n6247), .Z(n6245) );
  NAND U8772 ( .A(o[109]), .B(n5916), .Z(n6247) );
  NANDN U8773 ( .A(n5917), .B(creg[109]), .Z(n6246) );
  NAND U8774 ( .A(n6248), .B(n4861), .Z(n3491) );
  NANDN U8775 ( .A(init), .B(m[110]), .Z(n4861) );
  AND U8776 ( .A(n6249), .B(n6250), .Z(n6248) );
  NAND U8777 ( .A(o[110]), .B(n5916), .Z(n6250) );
  NANDN U8778 ( .A(n5917), .B(creg[110]), .Z(n6249) );
  NAND U8779 ( .A(n6251), .B(n4859), .Z(n3490) );
  NANDN U8780 ( .A(init), .B(m[111]), .Z(n4859) );
  AND U8781 ( .A(n6252), .B(n6253), .Z(n6251) );
  NAND U8782 ( .A(o[111]), .B(n5916), .Z(n6253) );
  NANDN U8783 ( .A(n5917), .B(creg[111]), .Z(n6252) );
  NAND U8784 ( .A(n6254), .B(n4857), .Z(n3489) );
  NANDN U8785 ( .A(init), .B(m[112]), .Z(n4857) );
  AND U8786 ( .A(n6255), .B(n6256), .Z(n6254) );
  NAND U8787 ( .A(o[112]), .B(n5916), .Z(n6256) );
  NANDN U8788 ( .A(n5917), .B(creg[112]), .Z(n6255) );
  NAND U8789 ( .A(n6257), .B(n4855), .Z(n3488) );
  NANDN U8790 ( .A(init), .B(m[113]), .Z(n4855) );
  AND U8791 ( .A(n6258), .B(n6259), .Z(n6257) );
  NAND U8792 ( .A(o[113]), .B(n5916), .Z(n6259) );
  NANDN U8793 ( .A(n5917), .B(creg[113]), .Z(n6258) );
  NAND U8794 ( .A(n6260), .B(n4853), .Z(n3487) );
  NANDN U8795 ( .A(init), .B(m[114]), .Z(n4853) );
  AND U8796 ( .A(n6261), .B(n6262), .Z(n6260) );
  NAND U8797 ( .A(o[114]), .B(n5916), .Z(n6262) );
  NANDN U8798 ( .A(n5917), .B(creg[114]), .Z(n6261) );
  NAND U8799 ( .A(n6263), .B(n4851), .Z(n3486) );
  NANDN U8800 ( .A(init), .B(m[115]), .Z(n4851) );
  AND U8801 ( .A(n6264), .B(n6265), .Z(n6263) );
  NAND U8802 ( .A(o[115]), .B(n5916), .Z(n6265) );
  NANDN U8803 ( .A(n5917), .B(creg[115]), .Z(n6264) );
  NAND U8804 ( .A(n6266), .B(n4849), .Z(n3485) );
  NANDN U8805 ( .A(init), .B(m[116]), .Z(n4849) );
  AND U8806 ( .A(n6267), .B(n6268), .Z(n6266) );
  NAND U8807 ( .A(o[116]), .B(n5916), .Z(n6268) );
  NANDN U8808 ( .A(n5917), .B(creg[116]), .Z(n6267) );
  NAND U8809 ( .A(n6269), .B(n4847), .Z(n3484) );
  NANDN U8810 ( .A(init), .B(m[117]), .Z(n4847) );
  AND U8811 ( .A(n6270), .B(n6271), .Z(n6269) );
  NAND U8812 ( .A(o[117]), .B(n5916), .Z(n6271) );
  NANDN U8813 ( .A(n5917), .B(creg[117]), .Z(n6270) );
  NAND U8814 ( .A(n6272), .B(n4845), .Z(n3483) );
  NANDN U8815 ( .A(init), .B(m[118]), .Z(n4845) );
  AND U8816 ( .A(n6273), .B(n6274), .Z(n6272) );
  NAND U8817 ( .A(o[118]), .B(n5916), .Z(n6274) );
  NANDN U8818 ( .A(n5917), .B(creg[118]), .Z(n6273) );
  NAND U8819 ( .A(n6275), .B(n4843), .Z(n3482) );
  NANDN U8820 ( .A(init), .B(m[119]), .Z(n4843) );
  AND U8821 ( .A(n6276), .B(n6277), .Z(n6275) );
  NAND U8822 ( .A(o[119]), .B(n5916), .Z(n6277) );
  NANDN U8823 ( .A(n5917), .B(creg[119]), .Z(n6276) );
  NAND U8824 ( .A(n6278), .B(n4839), .Z(n3481) );
  NANDN U8825 ( .A(init), .B(m[120]), .Z(n4839) );
  AND U8826 ( .A(n6279), .B(n6280), .Z(n6278) );
  NAND U8827 ( .A(o[120]), .B(n5916), .Z(n6280) );
  NANDN U8828 ( .A(n5917), .B(creg[120]), .Z(n6279) );
  NAND U8829 ( .A(n6281), .B(n4837), .Z(n3480) );
  NANDN U8830 ( .A(init), .B(m[121]), .Z(n4837) );
  AND U8831 ( .A(n6282), .B(n6283), .Z(n6281) );
  NAND U8832 ( .A(o[121]), .B(n5916), .Z(n6283) );
  NANDN U8833 ( .A(n5917), .B(creg[121]), .Z(n6282) );
  NAND U8834 ( .A(n6284), .B(n4835), .Z(n3479) );
  NANDN U8835 ( .A(init), .B(m[122]), .Z(n4835) );
  AND U8836 ( .A(n6285), .B(n6286), .Z(n6284) );
  NAND U8837 ( .A(o[122]), .B(n5916), .Z(n6286) );
  NANDN U8838 ( .A(n5917), .B(creg[122]), .Z(n6285) );
  NAND U8839 ( .A(n6287), .B(n4833), .Z(n3478) );
  NANDN U8840 ( .A(init), .B(m[123]), .Z(n4833) );
  AND U8841 ( .A(n6288), .B(n6289), .Z(n6287) );
  NAND U8842 ( .A(o[123]), .B(n5916), .Z(n6289) );
  NANDN U8843 ( .A(n5917), .B(creg[123]), .Z(n6288) );
  NAND U8844 ( .A(n6290), .B(n4831), .Z(n3477) );
  NANDN U8845 ( .A(init), .B(m[124]), .Z(n4831) );
  AND U8846 ( .A(n6291), .B(n6292), .Z(n6290) );
  NAND U8847 ( .A(o[124]), .B(n5916), .Z(n6292) );
  NANDN U8848 ( .A(n5917), .B(creg[124]), .Z(n6291) );
  NAND U8849 ( .A(n6293), .B(n4829), .Z(n3476) );
  NANDN U8850 ( .A(init), .B(m[125]), .Z(n4829) );
  AND U8851 ( .A(n6294), .B(n6295), .Z(n6293) );
  NAND U8852 ( .A(o[125]), .B(n5916), .Z(n6295) );
  NANDN U8853 ( .A(n5917), .B(creg[125]), .Z(n6294) );
  NAND U8854 ( .A(n6296), .B(n4827), .Z(n3475) );
  NANDN U8855 ( .A(init), .B(m[126]), .Z(n4827) );
  AND U8856 ( .A(n6297), .B(n6298), .Z(n6296) );
  NAND U8857 ( .A(o[126]), .B(n5916), .Z(n6298) );
  NANDN U8858 ( .A(n5917), .B(creg[126]), .Z(n6297) );
  NAND U8859 ( .A(n6299), .B(n4825), .Z(n3474) );
  NANDN U8860 ( .A(init), .B(m[127]), .Z(n4825) );
  AND U8861 ( .A(n6300), .B(n6301), .Z(n6299) );
  NAND U8862 ( .A(o[127]), .B(n5916), .Z(n6301) );
  NANDN U8863 ( .A(n5917), .B(creg[127]), .Z(n6300) );
  NAND U8864 ( .A(n6302), .B(n4823), .Z(n3473) );
  NANDN U8865 ( .A(init), .B(m[128]), .Z(n4823) );
  AND U8866 ( .A(n6303), .B(n6304), .Z(n6302) );
  NAND U8867 ( .A(o[128]), .B(n5916), .Z(n6304) );
  NANDN U8868 ( .A(n5917), .B(creg[128]), .Z(n6303) );
  NAND U8869 ( .A(n6305), .B(n4821), .Z(n3472) );
  NANDN U8870 ( .A(init), .B(m[129]), .Z(n4821) );
  AND U8871 ( .A(n6306), .B(n6307), .Z(n6305) );
  NAND U8872 ( .A(o[129]), .B(n5916), .Z(n6307) );
  NANDN U8873 ( .A(n5917), .B(creg[129]), .Z(n6306) );
  NAND U8874 ( .A(n6308), .B(n4817), .Z(n3471) );
  NANDN U8875 ( .A(init), .B(m[130]), .Z(n4817) );
  AND U8876 ( .A(n6309), .B(n6310), .Z(n6308) );
  NAND U8877 ( .A(o[130]), .B(n5916), .Z(n6310) );
  NANDN U8878 ( .A(n5917), .B(creg[130]), .Z(n6309) );
  NAND U8879 ( .A(n6311), .B(n4815), .Z(n3470) );
  NANDN U8880 ( .A(init), .B(m[131]), .Z(n4815) );
  AND U8881 ( .A(n6312), .B(n6313), .Z(n6311) );
  NAND U8882 ( .A(o[131]), .B(n5916), .Z(n6313) );
  NANDN U8883 ( .A(n5917), .B(creg[131]), .Z(n6312) );
  NAND U8884 ( .A(n6314), .B(n4813), .Z(n3469) );
  NANDN U8885 ( .A(init), .B(m[132]), .Z(n4813) );
  AND U8886 ( .A(n6315), .B(n6316), .Z(n6314) );
  NAND U8887 ( .A(o[132]), .B(n5916), .Z(n6316) );
  NANDN U8888 ( .A(n5917), .B(creg[132]), .Z(n6315) );
  NAND U8889 ( .A(n6317), .B(n4811), .Z(n3468) );
  NANDN U8890 ( .A(init), .B(m[133]), .Z(n4811) );
  AND U8891 ( .A(n6318), .B(n6319), .Z(n6317) );
  NAND U8892 ( .A(o[133]), .B(n5916), .Z(n6319) );
  NANDN U8893 ( .A(n5917), .B(creg[133]), .Z(n6318) );
  NAND U8894 ( .A(n6320), .B(n4809), .Z(n3467) );
  NANDN U8895 ( .A(init), .B(m[134]), .Z(n4809) );
  AND U8896 ( .A(n6321), .B(n6322), .Z(n6320) );
  NAND U8897 ( .A(o[134]), .B(n5916), .Z(n6322) );
  NANDN U8898 ( .A(n5917), .B(creg[134]), .Z(n6321) );
  NAND U8899 ( .A(n6323), .B(n4807), .Z(n3466) );
  NANDN U8900 ( .A(init), .B(m[135]), .Z(n4807) );
  AND U8901 ( .A(n6324), .B(n6325), .Z(n6323) );
  NAND U8902 ( .A(o[135]), .B(n5916), .Z(n6325) );
  NANDN U8903 ( .A(n5917), .B(creg[135]), .Z(n6324) );
  NAND U8904 ( .A(n6326), .B(n4805), .Z(n3465) );
  NANDN U8905 ( .A(init), .B(m[136]), .Z(n4805) );
  AND U8906 ( .A(n6327), .B(n6328), .Z(n6326) );
  NAND U8907 ( .A(o[136]), .B(n5916), .Z(n6328) );
  NANDN U8908 ( .A(n5917), .B(creg[136]), .Z(n6327) );
  NAND U8909 ( .A(n6329), .B(n4803), .Z(n3464) );
  NANDN U8910 ( .A(init), .B(m[137]), .Z(n4803) );
  AND U8911 ( .A(n6330), .B(n6331), .Z(n6329) );
  NAND U8912 ( .A(o[137]), .B(n5916), .Z(n6331) );
  NANDN U8913 ( .A(n5917), .B(creg[137]), .Z(n6330) );
  NAND U8914 ( .A(n6332), .B(n4801), .Z(n3463) );
  NANDN U8915 ( .A(init), .B(m[138]), .Z(n4801) );
  AND U8916 ( .A(n6333), .B(n6334), .Z(n6332) );
  NAND U8917 ( .A(o[138]), .B(n5916), .Z(n6334) );
  NANDN U8918 ( .A(n5917), .B(creg[138]), .Z(n6333) );
  NAND U8919 ( .A(n6335), .B(n4799), .Z(n3462) );
  NANDN U8920 ( .A(init), .B(m[139]), .Z(n4799) );
  AND U8921 ( .A(n6336), .B(n6337), .Z(n6335) );
  NAND U8922 ( .A(o[139]), .B(n5916), .Z(n6337) );
  NANDN U8923 ( .A(n5917), .B(creg[139]), .Z(n6336) );
  NAND U8924 ( .A(n6338), .B(n4795), .Z(n3461) );
  NANDN U8925 ( .A(init), .B(m[140]), .Z(n4795) );
  AND U8926 ( .A(n6339), .B(n6340), .Z(n6338) );
  NAND U8927 ( .A(o[140]), .B(n5916), .Z(n6340) );
  NANDN U8928 ( .A(n5917), .B(creg[140]), .Z(n6339) );
  NAND U8929 ( .A(n6341), .B(n4793), .Z(n3460) );
  NANDN U8930 ( .A(init), .B(m[141]), .Z(n4793) );
  AND U8931 ( .A(n6342), .B(n6343), .Z(n6341) );
  NAND U8932 ( .A(o[141]), .B(n5916), .Z(n6343) );
  NANDN U8933 ( .A(n5917), .B(creg[141]), .Z(n6342) );
  NAND U8934 ( .A(n6344), .B(n4791), .Z(n3459) );
  NANDN U8935 ( .A(init), .B(m[142]), .Z(n4791) );
  AND U8936 ( .A(n6345), .B(n6346), .Z(n6344) );
  NAND U8937 ( .A(o[142]), .B(n5916), .Z(n6346) );
  NANDN U8938 ( .A(n5917), .B(creg[142]), .Z(n6345) );
  NAND U8939 ( .A(n6347), .B(n4789), .Z(n3458) );
  NANDN U8940 ( .A(init), .B(m[143]), .Z(n4789) );
  AND U8941 ( .A(n6348), .B(n6349), .Z(n6347) );
  NAND U8942 ( .A(o[143]), .B(n5916), .Z(n6349) );
  NANDN U8943 ( .A(n5917), .B(creg[143]), .Z(n6348) );
  NAND U8944 ( .A(n6350), .B(n4787), .Z(n3457) );
  NANDN U8945 ( .A(init), .B(m[144]), .Z(n4787) );
  AND U8946 ( .A(n6351), .B(n6352), .Z(n6350) );
  NAND U8947 ( .A(o[144]), .B(n5916), .Z(n6352) );
  NANDN U8948 ( .A(n5917), .B(creg[144]), .Z(n6351) );
  NAND U8949 ( .A(n6353), .B(n4785), .Z(n3456) );
  NANDN U8950 ( .A(init), .B(m[145]), .Z(n4785) );
  AND U8951 ( .A(n6354), .B(n6355), .Z(n6353) );
  NAND U8952 ( .A(o[145]), .B(n5916), .Z(n6355) );
  NANDN U8953 ( .A(n5917), .B(creg[145]), .Z(n6354) );
  NAND U8954 ( .A(n6356), .B(n4783), .Z(n3455) );
  NANDN U8955 ( .A(init), .B(m[146]), .Z(n4783) );
  AND U8956 ( .A(n6357), .B(n6358), .Z(n6356) );
  NAND U8957 ( .A(o[146]), .B(n5916), .Z(n6358) );
  NANDN U8958 ( .A(n5917), .B(creg[146]), .Z(n6357) );
  NAND U8959 ( .A(n6359), .B(n4781), .Z(n3454) );
  NANDN U8960 ( .A(init), .B(m[147]), .Z(n4781) );
  AND U8961 ( .A(n6360), .B(n6361), .Z(n6359) );
  NAND U8962 ( .A(o[147]), .B(n5916), .Z(n6361) );
  NANDN U8963 ( .A(n5917), .B(creg[147]), .Z(n6360) );
  NAND U8964 ( .A(n6362), .B(n4779), .Z(n3453) );
  NANDN U8965 ( .A(init), .B(m[148]), .Z(n4779) );
  AND U8966 ( .A(n6363), .B(n6364), .Z(n6362) );
  NAND U8967 ( .A(o[148]), .B(n5916), .Z(n6364) );
  NANDN U8968 ( .A(n5917), .B(creg[148]), .Z(n6363) );
  NAND U8969 ( .A(n6365), .B(n4777), .Z(n3452) );
  NANDN U8970 ( .A(init), .B(m[149]), .Z(n4777) );
  AND U8971 ( .A(n6366), .B(n6367), .Z(n6365) );
  NAND U8972 ( .A(o[149]), .B(n5916), .Z(n6367) );
  NANDN U8973 ( .A(n5917), .B(creg[149]), .Z(n6366) );
  NAND U8974 ( .A(n6368), .B(n4773), .Z(n3451) );
  NANDN U8975 ( .A(init), .B(m[150]), .Z(n4773) );
  AND U8976 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U8977 ( .A(o[150]), .B(n5916), .Z(n6370) );
  NANDN U8978 ( .A(n5917), .B(creg[150]), .Z(n6369) );
  NAND U8979 ( .A(n6371), .B(n4771), .Z(n3450) );
  NANDN U8980 ( .A(init), .B(m[151]), .Z(n4771) );
  AND U8981 ( .A(n6372), .B(n6373), .Z(n6371) );
  NAND U8982 ( .A(o[151]), .B(n5916), .Z(n6373) );
  NANDN U8983 ( .A(n5917), .B(creg[151]), .Z(n6372) );
  NAND U8984 ( .A(n6374), .B(n4769), .Z(n3449) );
  NANDN U8985 ( .A(init), .B(m[152]), .Z(n4769) );
  AND U8986 ( .A(n6375), .B(n6376), .Z(n6374) );
  NAND U8987 ( .A(o[152]), .B(n5916), .Z(n6376) );
  NANDN U8988 ( .A(n5917), .B(creg[152]), .Z(n6375) );
  NAND U8989 ( .A(n6377), .B(n4767), .Z(n3448) );
  NANDN U8990 ( .A(init), .B(m[153]), .Z(n4767) );
  AND U8991 ( .A(n6378), .B(n6379), .Z(n6377) );
  NAND U8992 ( .A(o[153]), .B(n5916), .Z(n6379) );
  NANDN U8993 ( .A(n5917), .B(creg[153]), .Z(n6378) );
  NAND U8994 ( .A(n6380), .B(n4765), .Z(n3447) );
  NANDN U8995 ( .A(init), .B(m[154]), .Z(n4765) );
  AND U8996 ( .A(n6381), .B(n6382), .Z(n6380) );
  NAND U8997 ( .A(o[154]), .B(n5916), .Z(n6382) );
  NANDN U8998 ( .A(n5917), .B(creg[154]), .Z(n6381) );
  NAND U8999 ( .A(n6383), .B(n4763), .Z(n3446) );
  NANDN U9000 ( .A(init), .B(m[155]), .Z(n4763) );
  AND U9001 ( .A(n6384), .B(n6385), .Z(n6383) );
  NAND U9002 ( .A(o[155]), .B(n5916), .Z(n6385) );
  NANDN U9003 ( .A(n5917), .B(creg[155]), .Z(n6384) );
  NAND U9004 ( .A(n6386), .B(n4761), .Z(n3445) );
  NANDN U9005 ( .A(init), .B(m[156]), .Z(n4761) );
  AND U9006 ( .A(n6387), .B(n6388), .Z(n6386) );
  NAND U9007 ( .A(o[156]), .B(n5916), .Z(n6388) );
  NANDN U9008 ( .A(n5917), .B(creg[156]), .Z(n6387) );
  NAND U9009 ( .A(n6389), .B(n4759), .Z(n3444) );
  NANDN U9010 ( .A(init), .B(m[157]), .Z(n4759) );
  AND U9011 ( .A(n6390), .B(n6391), .Z(n6389) );
  NAND U9012 ( .A(o[157]), .B(n5916), .Z(n6391) );
  NANDN U9013 ( .A(n5917), .B(creg[157]), .Z(n6390) );
  NAND U9014 ( .A(n6392), .B(n4757), .Z(n3443) );
  NANDN U9015 ( .A(init), .B(m[158]), .Z(n4757) );
  AND U9016 ( .A(n6393), .B(n6394), .Z(n6392) );
  NAND U9017 ( .A(o[158]), .B(n5916), .Z(n6394) );
  NANDN U9018 ( .A(n5917), .B(creg[158]), .Z(n6393) );
  NAND U9019 ( .A(n6395), .B(n4755), .Z(n3442) );
  NANDN U9020 ( .A(init), .B(m[159]), .Z(n4755) );
  AND U9021 ( .A(n6396), .B(n6397), .Z(n6395) );
  NAND U9022 ( .A(o[159]), .B(n5916), .Z(n6397) );
  NANDN U9023 ( .A(n5917), .B(creg[159]), .Z(n6396) );
  NAND U9024 ( .A(n6398), .B(n4751), .Z(n3441) );
  NANDN U9025 ( .A(init), .B(m[160]), .Z(n4751) );
  AND U9026 ( .A(n6399), .B(n6400), .Z(n6398) );
  NAND U9027 ( .A(o[160]), .B(n5916), .Z(n6400) );
  NANDN U9028 ( .A(n5917), .B(creg[160]), .Z(n6399) );
  NAND U9029 ( .A(n6401), .B(n4749), .Z(n3440) );
  NANDN U9030 ( .A(init), .B(m[161]), .Z(n4749) );
  AND U9031 ( .A(n6402), .B(n6403), .Z(n6401) );
  NAND U9032 ( .A(o[161]), .B(n5916), .Z(n6403) );
  NANDN U9033 ( .A(n5917), .B(creg[161]), .Z(n6402) );
  NAND U9034 ( .A(n6404), .B(n4747), .Z(n3439) );
  NANDN U9035 ( .A(init), .B(m[162]), .Z(n4747) );
  AND U9036 ( .A(n6405), .B(n6406), .Z(n6404) );
  NAND U9037 ( .A(o[162]), .B(n5916), .Z(n6406) );
  NANDN U9038 ( .A(n5917), .B(creg[162]), .Z(n6405) );
  NAND U9039 ( .A(n6407), .B(n4745), .Z(n3438) );
  NANDN U9040 ( .A(init), .B(m[163]), .Z(n4745) );
  AND U9041 ( .A(n6408), .B(n6409), .Z(n6407) );
  NAND U9042 ( .A(o[163]), .B(n5916), .Z(n6409) );
  NANDN U9043 ( .A(n5917), .B(creg[163]), .Z(n6408) );
  NAND U9044 ( .A(n6410), .B(n4743), .Z(n3437) );
  NANDN U9045 ( .A(init), .B(m[164]), .Z(n4743) );
  AND U9046 ( .A(n6411), .B(n6412), .Z(n6410) );
  NAND U9047 ( .A(o[164]), .B(n5916), .Z(n6412) );
  NANDN U9048 ( .A(n5917), .B(creg[164]), .Z(n6411) );
  NAND U9049 ( .A(n6413), .B(n4741), .Z(n3436) );
  NANDN U9050 ( .A(init), .B(m[165]), .Z(n4741) );
  AND U9051 ( .A(n6414), .B(n6415), .Z(n6413) );
  NAND U9052 ( .A(o[165]), .B(n5916), .Z(n6415) );
  NANDN U9053 ( .A(n5917), .B(creg[165]), .Z(n6414) );
  NAND U9054 ( .A(n6416), .B(n4739), .Z(n3435) );
  NANDN U9055 ( .A(init), .B(m[166]), .Z(n4739) );
  AND U9056 ( .A(n6417), .B(n6418), .Z(n6416) );
  NAND U9057 ( .A(o[166]), .B(n5916), .Z(n6418) );
  NANDN U9058 ( .A(n5917), .B(creg[166]), .Z(n6417) );
  NAND U9059 ( .A(n6419), .B(n4737), .Z(n3434) );
  NANDN U9060 ( .A(init), .B(m[167]), .Z(n4737) );
  AND U9061 ( .A(n6420), .B(n6421), .Z(n6419) );
  NAND U9062 ( .A(o[167]), .B(n5916), .Z(n6421) );
  NANDN U9063 ( .A(n5917), .B(creg[167]), .Z(n6420) );
  NAND U9064 ( .A(n6422), .B(n4735), .Z(n3433) );
  NANDN U9065 ( .A(init), .B(m[168]), .Z(n4735) );
  AND U9066 ( .A(n6423), .B(n6424), .Z(n6422) );
  NAND U9067 ( .A(o[168]), .B(n5916), .Z(n6424) );
  NANDN U9068 ( .A(n5917), .B(creg[168]), .Z(n6423) );
  NAND U9069 ( .A(n6425), .B(n4733), .Z(n3432) );
  NANDN U9070 ( .A(init), .B(m[169]), .Z(n4733) );
  AND U9071 ( .A(n6426), .B(n6427), .Z(n6425) );
  NAND U9072 ( .A(o[169]), .B(n5916), .Z(n6427) );
  NANDN U9073 ( .A(n5917), .B(creg[169]), .Z(n6426) );
  NAND U9074 ( .A(n6428), .B(n4729), .Z(n3431) );
  NANDN U9075 ( .A(init), .B(m[170]), .Z(n4729) );
  AND U9076 ( .A(n6429), .B(n6430), .Z(n6428) );
  NAND U9077 ( .A(o[170]), .B(n5916), .Z(n6430) );
  NANDN U9078 ( .A(n5917), .B(creg[170]), .Z(n6429) );
  NAND U9079 ( .A(n6431), .B(n4727), .Z(n3430) );
  NANDN U9080 ( .A(init), .B(m[171]), .Z(n4727) );
  AND U9081 ( .A(n6432), .B(n6433), .Z(n6431) );
  NAND U9082 ( .A(o[171]), .B(n5916), .Z(n6433) );
  NANDN U9083 ( .A(n5917), .B(creg[171]), .Z(n6432) );
  NAND U9084 ( .A(n6434), .B(n4725), .Z(n3429) );
  NANDN U9085 ( .A(init), .B(m[172]), .Z(n4725) );
  AND U9086 ( .A(n6435), .B(n6436), .Z(n6434) );
  NAND U9087 ( .A(o[172]), .B(n5916), .Z(n6436) );
  NANDN U9088 ( .A(n5917), .B(creg[172]), .Z(n6435) );
  NAND U9089 ( .A(n6437), .B(n4723), .Z(n3428) );
  NANDN U9090 ( .A(init), .B(m[173]), .Z(n4723) );
  AND U9091 ( .A(n6438), .B(n6439), .Z(n6437) );
  NAND U9092 ( .A(o[173]), .B(n5916), .Z(n6439) );
  NANDN U9093 ( .A(n5917), .B(creg[173]), .Z(n6438) );
  NAND U9094 ( .A(n6440), .B(n4721), .Z(n3427) );
  NANDN U9095 ( .A(init), .B(m[174]), .Z(n4721) );
  AND U9096 ( .A(n6441), .B(n6442), .Z(n6440) );
  NAND U9097 ( .A(o[174]), .B(n5916), .Z(n6442) );
  NANDN U9098 ( .A(n5917), .B(creg[174]), .Z(n6441) );
  NAND U9099 ( .A(n6443), .B(n4719), .Z(n3426) );
  NANDN U9100 ( .A(init), .B(m[175]), .Z(n4719) );
  AND U9101 ( .A(n6444), .B(n6445), .Z(n6443) );
  NAND U9102 ( .A(o[175]), .B(n5916), .Z(n6445) );
  NANDN U9103 ( .A(n5917), .B(creg[175]), .Z(n6444) );
  NAND U9104 ( .A(n6446), .B(n4717), .Z(n3425) );
  NANDN U9105 ( .A(init), .B(m[176]), .Z(n4717) );
  AND U9106 ( .A(n6447), .B(n6448), .Z(n6446) );
  NAND U9107 ( .A(o[176]), .B(n5916), .Z(n6448) );
  NANDN U9108 ( .A(n5917), .B(creg[176]), .Z(n6447) );
  NAND U9109 ( .A(n6449), .B(n4715), .Z(n3424) );
  NANDN U9110 ( .A(init), .B(m[177]), .Z(n4715) );
  AND U9111 ( .A(n6450), .B(n6451), .Z(n6449) );
  NAND U9112 ( .A(o[177]), .B(n5916), .Z(n6451) );
  NANDN U9113 ( .A(n5917), .B(creg[177]), .Z(n6450) );
  NAND U9114 ( .A(n6452), .B(n4713), .Z(n3423) );
  NANDN U9115 ( .A(init), .B(m[178]), .Z(n4713) );
  AND U9116 ( .A(n6453), .B(n6454), .Z(n6452) );
  NAND U9117 ( .A(o[178]), .B(n5916), .Z(n6454) );
  NANDN U9118 ( .A(n5917), .B(creg[178]), .Z(n6453) );
  NAND U9119 ( .A(n6455), .B(n4711), .Z(n3422) );
  NANDN U9120 ( .A(init), .B(m[179]), .Z(n4711) );
  AND U9121 ( .A(n6456), .B(n6457), .Z(n6455) );
  NAND U9122 ( .A(o[179]), .B(n5916), .Z(n6457) );
  NANDN U9123 ( .A(n5917), .B(creg[179]), .Z(n6456) );
  NAND U9124 ( .A(n6458), .B(n4707), .Z(n3421) );
  NANDN U9125 ( .A(init), .B(m[180]), .Z(n4707) );
  AND U9126 ( .A(n6459), .B(n6460), .Z(n6458) );
  NAND U9127 ( .A(o[180]), .B(n5916), .Z(n6460) );
  NANDN U9128 ( .A(n5917), .B(creg[180]), .Z(n6459) );
  NAND U9129 ( .A(n6461), .B(n4705), .Z(n3420) );
  NANDN U9130 ( .A(init), .B(m[181]), .Z(n4705) );
  AND U9131 ( .A(n6462), .B(n6463), .Z(n6461) );
  NAND U9132 ( .A(o[181]), .B(n5916), .Z(n6463) );
  NANDN U9133 ( .A(n5917), .B(creg[181]), .Z(n6462) );
  NAND U9134 ( .A(n6464), .B(n4703), .Z(n3419) );
  NANDN U9135 ( .A(init), .B(m[182]), .Z(n4703) );
  AND U9136 ( .A(n6465), .B(n6466), .Z(n6464) );
  NAND U9137 ( .A(o[182]), .B(n5916), .Z(n6466) );
  NANDN U9138 ( .A(n5917), .B(creg[182]), .Z(n6465) );
  NAND U9139 ( .A(n6467), .B(n4701), .Z(n3418) );
  NANDN U9140 ( .A(init), .B(m[183]), .Z(n4701) );
  AND U9141 ( .A(n6468), .B(n6469), .Z(n6467) );
  NAND U9142 ( .A(o[183]), .B(n5916), .Z(n6469) );
  NANDN U9143 ( .A(n5917), .B(creg[183]), .Z(n6468) );
  NAND U9144 ( .A(n6470), .B(n4699), .Z(n3417) );
  NANDN U9145 ( .A(init), .B(m[184]), .Z(n4699) );
  AND U9146 ( .A(n6471), .B(n6472), .Z(n6470) );
  NAND U9147 ( .A(o[184]), .B(n5916), .Z(n6472) );
  NANDN U9148 ( .A(n5917), .B(creg[184]), .Z(n6471) );
  NAND U9149 ( .A(n6473), .B(n4697), .Z(n3416) );
  NANDN U9150 ( .A(init), .B(m[185]), .Z(n4697) );
  AND U9151 ( .A(n6474), .B(n6475), .Z(n6473) );
  NAND U9152 ( .A(o[185]), .B(n5916), .Z(n6475) );
  NANDN U9153 ( .A(n5917), .B(creg[185]), .Z(n6474) );
  NAND U9154 ( .A(n6476), .B(n4695), .Z(n3415) );
  NANDN U9155 ( .A(init), .B(m[186]), .Z(n4695) );
  AND U9156 ( .A(n6477), .B(n6478), .Z(n6476) );
  NAND U9157 ( .A(o[186]), .B(n5916), .Z(n6478) );
  NANDN U9158 ( .A(n5917), .B(creg[186]), .Z(n6477) );
  NAND U9159 ( .A(n6479), .B(n4693), .Z(n3414) );
  NANDN U9160 ( .A(init), .B(m[187]), .Z(n4693) );
  AND U9161 ( .A(n6480), .B(n6481), .Z(n6479) );
  NAND U9162 ( .A(o[187]), .B(n5916), .Z(n6481) );
  NANDN U9163 ( .A(n5917), .B(creg[187]), .Z(n6480) );
  NAND U9164 ( .A(n6482), .B(n4691), .Z(n3413) );
  NANDN U9165 ( .A(init), .B(m[188]), .Z(n4691) );
  AND U9166 ( .A(n6483), .B(n6484), .Z(n6482) );
  NAND U9167 ( .A(o[188]), .B(n5916), .Z(n6484) );
  NANDN U9168 ( .A(n5917), .B(creg[188]), .Z(n6483) );
  NAND U9169 ( .A(n6485), .B(n4689), .Z(n3412) );
  NANDN U9170 ( .A(init), .B(m[189]), .Z(n4689) );
  AND U9171 ( .A(n6486), .B(n6487), .Z(n6485) );
  NAND U9172 ( .A(o[189]), .B(n5916), .Z(n6487) );
  NANDN U9173 ( .A(n5917), .B(creg[189]), .Z(n6486) );
  NAND U9174 ( .A(n6488), .B(n4685), .Z(n3411) );
  NANDN U9175 ( .A(init), .B(m[190]), .Z(n4685) );
  AND U9176 ( .A(n6489), .B(n6490), .Z(n6488) );
  NAND U9177 ( .A(o[190]), .B(n5916), .Z(n6490) );
  NANDN U9178 ( .A(n5917), .B(creg[190]), .Z(n6489) );
  NAND U9179 ( .A(n6491), .B(n4683), .Z(n3410) );
  NANDN U9180 ( .A(init), .B(m[191]), .Z(n4683) );
  AND U9181 ( .A(n6492), .B(n6493), .Z(n6491) );
  NAND U9182 ( .A(o[191]), .B(n5916), .Z(n6493) );
  NANDN U9183 ( .A(n5917), .B(creg[191]), .Z(n6492) );
  NAND U9184 ( .A(n6494), .B(n4681), .Z(n3409) );
  NANDN U9185 ( .A(init), .B(m[192]), .Z(n4681) );
  AND U9186 ( .A(n6495), .B(n6496), .Z(n6494) );
  NAND U9187 ( .A(o[192]), .B(n5916), .Z(n6496) );
  NANDN U9188 ( .A(n5917), .B(creg[192]), .Z(n6495) );
  NAND U9189 ( .A(n6497), .B(n4679), .Z(n3408) );
  NANDN U9190 ( .A(init), .B(m[193]), .Z(n4679) );
  AND U9191 ( .A(n6498), .B(n6499), .Z(n6497) );
  NAND U9192 ( .A(o[193]), .B(n5916), .Z(n6499) );
  NANDN U9193 ( .A(n5917), .B(creg[193]), .Z(n6498) );
  NAND U9194 ( .A(n6500), .B(n4677), .Z(n3407) );
  NANDN U9195 ( .A(init), .B(m[194]), .Z(n4677) );
  AND U9196 ( .A(n6501), .B(n6502), .Z(n6500) );
  NAND U9197 ( .A(o[194]), .B(n5916), .Z(n6502) );
  NANDN U9198 ( .A(n5917), .B(creg[194]), .Z(n6501) );
  NAND U9199 ( .A(n6503), .B(n4675), .Z(n3406) );
  NANDN U9200 ( .A(init), .B(m[195]), .Z(n4675) );
  AND U9201 ( .A(n6504), .B(n6505), .Z(n6503) );
  NAND U9202 ( .A(o[195]), .B(n5916), .Z(n6505) );
  NANDN U9203 ( .A(n5917), .B(creg[195]), .Z(n6504) );
  NAND U9204 ( .A(n6506), .B(n4673), .Z(n3405) );
  NANDN U9205 ( .A(init), .B(m[196]), .Z(n4673) );
  AND U9206 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U9207 ( .A(o[196]), .B(n5916), .Z(n6508) );
  NANDN U9208 ( .A(n5917), .B(creg[196]), .Z(n6507) );
  NAND U9209 ( .A(n6509), .B(n4671), .Z(n3404) );
  NANDN U9210 ( .A(init), .B(m[197]), .Z(n4671) );
  AND U9211 ( .A(n6510), .B(n6511), .Z(n6509) );
  NAND U9212 ( .A(o[197]), .B(n5916), .Z(n6511) );
  NANDN U9213 ( .A(n5917), .B(creg[197]), .Z(n6510) );
  NAND U9214 ( .A(n6512), .B(n4669), .Z(n3403) );
  NANDN U9215 ( .A(init), .B(m[198]), .Z(n4669) );
  AND U9216 ( .A(n6513), .B(n6514), .Z(n6512) );
  NAND U9217 ( .A(o[198]), .B(n5916), .Z(n6514) );
  NANDN U9218 ( .A(n5917), .B(creg[198]), .Z(n6513) );
  NAND U9219 ( .A(n6515), .B(n4667), .Z(n3402) );
  NANDN U9220 ( .A(init), .B(m[199]), .Z(n4667) );
  AND U9221 ( .A(n6516), .B(n6517), .Z(n6515) );
  NAND U9222 ( .A(o[199]), .B(n5916), .Z(n6517) );
  NANDN U9223 ( .A(n5917), .B(creg[199]), .Z(n6516) );
  NAND U9224 ( .A(n6518), .B(n4661), .Z(n3401) );
  NANDN U9225 ( .A(init), .B(m[200]), .Z(n4661) );
  AND U9226 ( .A(n6519), .B(n6520), .Z(n6518) );
  NAND U9227 ( .A(o[200]), .B(n5916), .Z(n6520) );
  NANDN U9228 ( .A(n5917), .B(creg[200]), .Z(n6519) );
  NAND U9229 ( .A(n6521), .B(n4659), .Z(n3400) );
  NANDN U9230 ( .A(init), .B(m[201]), .Z(n4659) );
  AND U9231 ( .A(n6522), .B(n6523), .Z(n6521) );
  NAND U9232 ( .A(o[201]), .B(n5916), .Z(n6523) );
  NANDN U9233 ( .A(n5917), .B(creg[201]), .Z(n6522) );
  NAND U9234 ( .A(n6524), .B(n4657), .Z(n3399) );
  NANDN U9235 ( .A(init), .B(m[202]), .Z(n4657) );
  AND U9236 ( .A(n6525), .B(n6526), .Z(n6524) );
  NAND U9237 ( .A(o[202]), .B(n5916), .Z(n6526) );
  NANDN U9238 ( .A(n5917), .B(creg[202]), .Z(n6525) );
  NAND U9239 ( .A(n6527), .B(n4655), .Z(n3398) );
  NANDN U9240 ( .A(init), .B(m[203]), .Z(n4655) );
  AND U9241 ( .A(n6528), .B(n6529), .Z(n6527) );
  NAND U9242 ( .A(o[203]), .B(n5916), .Z(n6529) );
  NANDN U9243 ( .A(n5917), .B(creg[203]), .Z(n6528) );
  NAND U9244 ( .A(n6530), .B(n4653), .Z(n3397) );
  NANDN U9245 ( .A(init), .B(m[204]), .Z(n4653) );
  AND U9246 ( .A(n6531), .B(n6532), .Z(n6530) );
  NAND U9247 ( .A(o[204]), .B(n5916), .Z(n6532) );
  NANDN U9248 ( .A(n5917), .B(creg[204]), .Z(n6531) );
  NAND U9249 ( .A(n6533), .B(n4651), .Z(n3396) );
  NANDN U9250 ( .A(init), .B(m[205]), .Z(n4651) );
  AND U9251 ( .A(n6534), .B(n6535), .Z(n6533) );
  NAND U9252 ( .A(o[205]), .B(n5916), .Z(n6535) );
  NANDN U9253 ( .A(n5917), .B(creg[205]), .Z(n6534) );
  NAND U9254 ( .A(n6536), .B(n4649), .Z(n3395) );
  NANDN U9255 ( .A(init), .B(m[206]), .Z(n4649) );
  AND U9256 ( .A(n6537), .B(n6538), .Z(n6536) );
  NAND U9257 ( .A(o[206]), .B(n5916), .Z(n6538) );
  NANDN U9258 ( .A(n5917), .B(creg[206]), .Z(n6537) );
  NAND U9259 ( .A(n6539), .B(n4647), .Z(n3394) );
  NANDN U9260 ( .A(init), .B(m[207]), .Z(n4647) );
  AND U9261 ( .A(n6540), .B(n6541), .Z(n6539) );
  NAND U9262 ( .A(o[207]), .B(n5916), .Z(n6541) );
  NANDN U9263 ( .A(n5917), .B(creg[207]), .Z(n6540) );
  NAND U9264 ( .A(n6542), .B(n4645), .Z(n3393) );
  NANDN U9265 ( .A(init), .B(m[208]), .Z(n4645) );
  AND U9266 ( .A(n6543), .B(n6544), .Z(n6542) );
  NAND U9267 ( .A(o[208]), .B(n5916), .Z(n6544) );
  NANDN U9268 ( .A(n5917), .B(creg[208]), .Z(n6543) );
  NAND U9269 ( .A(n6545), .B(n4643), .Z(n3392) );
  NANDN U9270 ( .A(init), .B(m[209]), .Z(n4643) );
  AND U9271 ( .A(n6546), .B(n6547), .Z(n6545) );
  NAND U9272 ( .A(o[209]), .B(n5916), .Z(n6547) );
  NANDN U9273 ( .A(n5917), .B(creg[209]), .Z(n6546) );
  NAND U9274 ( .A(n6548), .B(n4639), .Z(n3391) );
  NANDN U9275 ( .A(init), .B(m[210]), .Z(n4639) );
  AND U9276 ( .A(n6549), .B(n6550), .Z(n6548) );
  NAND U9277 ( .A(o[210]), .B(n5916), .Z(n6550) );
  NANDN U9278 ( .A(n5917), .B(creg[210]), .Z(n6549) );
  NAND U9279 ( .A(n6551), .B(n4637), .Z(n3390) );
  NANDN U9280 ( .A(init), .B(m[211]), .Z(n4637) );
  AND U9281 ( .A(n6552), .B(n6553), .Z(n6551) );
  NAND U9282 ( .A(o[211]), .B(n5916), .Z(n6553) );
  NANDN U9283 ( .A(n5917), .B(creg[211]), .Z(n6552) );
  NAND U9284 ( .A(n6554), .B(n4635), .Z(n3389) );
  NANDN U9285 ( .A(init), .B(m[212]), .Z(n4635) );
  AND U9286 ( .A(n6555), .B(n6556), .Z(n6554) );
  NAND U9287 ( .A(o[212]), .B(n5916), .Z(n6556) );
  NANDN U9288 ( .A(n5917), .B(creg[212]), .Z(n6555) );
  NAND U9289 ( .A(n6557), .B(n4633), .Z(n3388) );
  NANDN U9290 ( .A(init), .B(m[213]), .Z(n4633) );
  AND U9291 ( .A(n6558), .B(n6559), .Z(n6557) );
  NAND U9292 ( .A(o[213]), .B(n5916), .Z(n6559) );
  NANDN U9293 ( .A(n5917), .B(creg[213]), .Z(n6558) );
  NAND U9294 ( .A(n6560), .B(n4631), .Z(n3387) );
  NANDN U9295 ( .A(init), .B(m[214]), .Z(n4631) );
  AND U9296 ( .A(n6561), .B(n6562), .Z(n6560) );
  NAND U9297 ( .A(o[214]), .B(n5916), .Z(n6562) );
  NANDN U9298 ( .A(n5917), .B(creg[214]), .Z(n6561) );
  NAND U9299 ( .A(n6563), .B(n4629), .Z(n3386) );
  NANDN U9300 ( .A(init), .B(m[215]), .Z(n4629) );
  AND U9301 ( .A(n6564), .B(n6565), .Z(n6563) );
  NAND U9302 ( .A(o[215]), .B(n5916), .Z(n6565) );
  NANDN U9303 ( .A(n5917), .B(creg[215]), .Z(n6564) );
  NAND U9304 ( .A(n6566), .B(n4627), .Z(n3385) );
  NANDN U9305 ( .A(init), .B(m[216]), .Z(n4627) );
  AND U9306 ( .A(n6567), .B(n6568), .Z(n6566) );
  NAND U9307 ( .A(o[216]), .B(n5916), .Z(n6568) );
  NANDN U9308 ( .A(n5917), .B(creg[216]), .Z(n6567) );
  NAND U9309 ( .A(n6569), .B(n4625), .Z(n3384) );
  NANDN U9310 ( .A(init), .B(m[217]), .Z(n4625) );
  AND U9311 ( .A(n6570), .B(n6571), .Z(n6569) );
  NAND U9312 ( .A(o[217]), .B(n5916), .Z(n6571) );
  NANDN U9313 ( .A(n5917), .B(creg[217]), .Z(n6570) );
  NAND U9314 ( .A(n6572), .B(n4623), .Z(n3383) );
  NANDN U9315 ( .A(init), .B(m[218]), .Z(n4623) );
  AND U9316 ( .A(n6573), .B(n6574), .Z(n6572) );
  NAND U9317 ( .A(o[218]), .B(n5916), .Z(n6574) );
  NANDN U9318 ( .A(n5917), .B(creg[218]), .Z(n6573) );
  NAND U9319 ( .A(n6575), .B(n4621), .Z(n3382) );
  NANDN U9320 ( .A(init), .B(m[219]), .Z(n4621) );
  AND U9321 ( .A(n6576), .B(n6577), .Z(n6575) );
  NAND U9322 ( .A(o[219]), .B(n5916), .Z(n6577) );
  NANDN U9323 ( .A(n5917), .B(creg[219]), .Z(n6576) );
  NAND U9324 ( .A(n6578), .B(n4617), .Z(n3381) );
  NANDN U9325 ( .A(init), .B(m[220]), .Z(n4617) );
  AND U9326 ( .A(n6579), .B(n6580), .Z(n6578) );
  NAND U9327 ( .A(o[220]), .B(n5916), .Z(n6580) );
  NANDN U9328 ( .A(n5917), .B(creg[220]), .Z(n6579) );
  NAND U9329 ( .A(n6581), .B(n4615), .Z(n3380) );
  NANDN U9330 ( .A(init), .B(m[221]), .Z(n4615) );
  AND U9331 ( .A(n6582), .B(n6583), .Z(n6581) );
  NAND U9332 ( .A(o[221]), .B(n5916), .Z(n6583) );
  NANDN U9333 ( .A(n5917), .B(creg[221]), .Z(n6582) );
  NAND U9334 ( .A(n6584), .B(n4613), .Z(n3379) );
  NANDN U9335 ( .A(init), .B(m[222]), .Z(n4613) );
  AND U9336 ( .A(n6585), .B(n6586), .Z(n6584) );
  NAND U9337 ( .A(o[222]), .B(n5916), .Z(n6586) );
  NANDN U9338 ( .A(n5917), .B(creg[222]), .Z(n6585) );
  NAND U9339 ( .A(n6587), .B(n4611), .Z(n3378) );
  NANDN U9340 ( .A(init), .B(m[223]), .Z(n4611) );
  AND U9341 ( .A(n6588), .B(n6589), .Z(n6587) );
  NAND U9342 ( .A(o[223]), .B(n5916), .Z(n6589) );
  NANDN U9343 ( .A(n5917), .B(creg[223]), .Z(n6588) );
  NAND U9344 ( .A(n6590), .B(n4609), .Z(n3377) );
  NANDN U9345 ( .A(init), .B(m[224]), .Z(n4609) );
  AND U9346 ( .A(n6591), .B(n6592), .Z(n6590) );
  NAND U9347 ( .A(o[224]), .B(n5916), .Z(n6592) );
  NANDN U9348 ( .A(n5917), .B(creg[224]), .Z(n6591) );
  NAND U9349 ( .A(n6593), .B(n4607), .Z(n3376) );
  NANDN U9350 ( .A(init), .B(m[225]), .Z(n4607) );
  AND U9351 ( .A(n6594), .B(n6595), .Z(n6593) );
  NAND U9352 ( .A(o[225]), .B(n5916), .Z(n6595) );
  NANDN U9353 ( .A(n5917), .B(creg[225]), .Z(n6594) );
  NAND U9354 ( .A(n6596), .B(n4605), .Z(n3375) );
  NANDN U9355 ( .A(init), .B(m[226]), .Z(n4605) );
  AND U9356 ( .A(n6597), .B(n6598), .Z(n6596) );
  NAND U9357 ( .A(o[226]), .B(n5916), .Z(n6598) );
  NANDN U9358 ( .A(n5917), .B(creg[226]), .Z(n6597) );
  NAND U9359 ( .A(n6599), .B(n4603), .Z(n3374) );
  NANDN U9360 ( .A(init), .B(m[227]), .Z(n4603) );
  AND U9361 ( .A(n6600), .B(n6601), .Z(n6599) );
  NAND U9362 ( .A(o[227]), .B(n5916), .Z(n6601) );
  NANDN U9363 ( .A(n5917), .B(creg[227]), .Z(n6600) );
  NAND U9364 ( .A(n6602), .B(n4601), .Z(n3373) );
  NANDN U9365 ( .A(init), .B(m[228]), .Z(n4601) );
  AND U9366 ( .A(n6603), .B(n6604), .Z(n6602) );
  NAND U9367 ( .A(o[228]), .B(n5916), .Z(n6604) );
  NANDN U9368 ( .A(n5917), .B(creg[228]), .Z(n6603) );
  NAND U9369 ( .A(n6605), .B(n4599), .Z(n3372) );
  NANDN U9370 ( .A(init), .B(m[229]), .Z(n4599) );
  AND U9371 ( .A(n6606), .B(n6607), .Z(n6605) );
  NAND U9372 ( .A(o[229]), .B(n5916), .Z(n6607) );
  NANDN U9373 ( .A(n5917), .B(creg[229]), .Z(n6606) );
  NAND U9374 ( .A(n6608), .B(n4595), .Z(n3371) );
  NANDN U9375 ( .A(init), .B(m[230]), .Z(n4595) );
  AND U9376 ( .A(n6609), .B(n6610), .Z(n6608) );
  NAND U9377 ( .A(o[230]), .B(n5916), .Z(n6610) );
  NANDN U9378 ( .A(n5917), .B(creg[230]), .Z(n6609) );
  NAND U9379 ( .A(n6611), .B(n4593), .Z(n3370) );
  NANDN U9380 ( .A(init), .B(m[231]), .Z(n4593) );
  AND U9381 ( .A(n6612), .B(n6613), .Z(n6611) );
  NAND U9382 ( .A(o[231]), .B(n5916), .Z(n6613) );
  NANDN U9383 ( .A(n5917), .B(creg[231]), .Z(n6612) );
  NAND U9384 ( .A(n6614), .B(n4591), .Z(n3369) );
  NANDN U9385 ( .A(init), .B(m[232]), .Z(n4591) );
  AND U9386 ( .A(n6615), .B(n6616), .Z(n6614) );
  NAND U9387 ( .A(o[232]), .B(n5916), .Z(n6616) );
  NANDN U9388 ( .A(n5917), .B(creg[232]), .Z(n6615) );
  NAND U9389 ( .A(n6617), .B(n4589), .Z(n3368) );
  NANDN U9390 ( .A(init), .B(m[233]), .Z(n4589) );
  AND U9391 ( .A(n6618), .B(n6619), .Z(n6617) );
  NAND U9392 ( .A(o[233]), .B(n5916), .Z(n6619) );
  NANDN U9393 ( .A(n5917), .B(creg[233]), .Z(n6618) );
  NAND U9394 ( .A(n6620), .B(n4587), .Z(n3367) );
  NANDN U9395 ( .A(init), .B(m[234]), .Z(n4587) );
  AND U9396 ( .A(n6621), .B(n6622), .Z(n6620) );
  NAND U9397 ( .A(o[234]), .B(n5916), .Z(n6622) );
  NANDN U9398 ( .A(n5917), .B(creg[234]), .Z(n6621) );
  NAND U9399 ( .A(n6623), .B(n4585), .Z(n3366) );
  NANDN U9400 ( .A(init), .B(m[235]), .Z(n4585) );
  AND U9401 ( .A(n6624), .B(n6625), .Z(n6623) );
  NAND U9402 ( .A(o[235]), .B(n5916), .Z(n6625) );
  NANDN U9403 ( .A(n5917), .B(creg[235]), .Z(n6624) );
  NAND U9404 ( .A(n6626), .B(n4583), .Z(n3365) );
  NANDN U9405 ( .A(init), .B(m[236]), .Z(n4583) );
  AND U9406 ( .A(n6627), .B(n6628), .Z(n6626) );
  NAND U9407 ( .A(o[236]), .B(n5916), .Z(n6628) );
  NANDN U9408 ( .A(n5917), .B(creg[236]), .Z(n6627) );
  NAND U9409 ( .A(n6629), .B(n4581), .Z(n3364) );
  NANDN U9410 ( .A(init), .B(m[237]), .Z(n4581) );
  AND U9411 ( .A(n6630), .B(n6631), .Z(n6629) );
  NAND U9412 ( .A(o[237]), .B(n5916), .Z(n6631) );
  NANDN U9413 ( .A(n5917), .B(creg[237]), .Z(n6630) );
  NAND U9414 ( .A(n6632), .B(n4579), .Z(n3363) );
  NANDN U9415 ( .A(init), .B(m[238]), .Z(n4579) );
  AND U9416 ( .A(n6633), .B(n6634), .Z(n6632) );
  NAND U9417 ( .A(o[238]), .B(n5916), .Z(n6634) );
  NANDN U9418 ( .A(n5917), .B(creg[238]), .Z(n6633) );
  NAND U9419 ( .A(n6635), .B(n4577), .Z(n3362) );
  NANDN U9420 ( .A(init), .B(m[239]), .Z(n4577) );
  AND U9421 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U9422 ( .A(o[239]), .B(n5916), .Z(n6637) );
  NANDN U9423 ( .A(n5917), .B(creg[239]), .Z(n6636) );
  NAND U9424 ( .A(n6638), .B(n4573), .Z(n3361) );
  NANDN U9425 ( .A(init), .B(m[240]), .Z(n4573) );
  AND U9426 ( .A(n6639), .B(n6640), .Z(n6638) );
  NAND U9427 ( .A(o[240]), .B(n5916), .Z(n6640) );
  NANDN U9428 ( .A(n5917), .B(creg[240]), .Z(n6639) );
  NAND U9429 ( .A(n6641), .B(n4571), .Z(n3360) );
  NANDN U9430 ( .A(init), .B(m[241]), .Z(n4571) );
  AND U9431 ( .A(n6642), .B(n6643), .Z(n6641) );
  NAND U9432 ( .A(o[241]), .B(n5916), .Z(n6643) );
  NANDN U9433 ( .A(n5917), .B(creg[241]), .Z(n6642) );
  NAND U9434 ( .A(n6644), .B(n4569), .Z(n3359) );
  NANDN U9435 ( .A(init), .B(m[242]), .Z(n4569) );
  AND U9436 ( .A(n6645), .B(n6646), .Z(n6644) );
  NAND U9437 ( .A(o[242]), .B(n5916), .Z(n6646) );
  NANDN U9438 ( .A(n5917), .B(creg[242]), .Z(n6645) );
  NAND U9439 ( .A(n6647), .B(n4567), .Z(n3358) );
  NANDN U9440 ( .A(init), .B(m[243]), .Z(n4567) );
  AND U9441 ( .A(n6648), .B(n6649), .Z(n6647) );
  NAND U9442 ( .A(o[243]), .B(n5916), .Z(n6649) );
  NANDN U9443 ( .A(n5917), .B(creg[243]), .Z(n6648) );
  NAND U9444 ( .A(n6650), .B(n4565), .Z(n3357) );
  NANDN U9445 ( .A(init), .B(m[244]), .Z(n4565) );
  AND U9446 ( .A(n6651), .B(n6652), .Z(n6650) );
  NAND U9447 ( .A(o[244]), .B(n5916), .Z(n6652) );
  NANDN U9448 ( .A(n5917), .B(creg[244]), .Z(n6651) );
  NAND U9449 ( .A(n6653), .B(n4563), .Z(n3356) );
  NANDN U9450 ( .A(init), .B(m[245]), .Z(n4563) );
  AND U9451 ( .A(n6654), .B(n6655), .Z(n6653) );
  NAND U9452 ( .A(o[245]), .B(n5916), .Z(n6655) );
  NANDN U9453 ( .A(n5917), .B(creg[245]), .Z(n6654) );
  NAND U9454 ( .A(n6656), .B(n4561), .Z(n3355) );
  NANDN U9455 ( .A(init), .B(m[246]), .Z(n4561) );
  AND U9456 ( .A(n6657), .B(n6658), .Z(n6656) );
  NAND U9457 ( .A(o[246]), .B(n5916), .Z(n6658) );
  NANDN U9458 ( .A(n5917), .B(creg[246]), .Z(n6657) );
  NAND U9459 ( .A(n6659), .B(n4559), .Z(n3354) );
  NANDN U9460 ( .A(init), .B(m[247]), .Z(n4559) );
  AND U9461 ( .A(n6660), .B(n6661), .Z(n6659) );
  NAND U9462 ( .A(o[247]), .B(n5916), .Z(n6661) );
  NANDN U9463 ( .A(n5917), .B(creg[247]), .Z(n6660) );
  NAND U9464 ( .A(n6662), .B(n4557), .Z(n3353) );
  NANDN U9465 ( .A(init), .B(m[248]), .Z(n4557) );
  AND U9466 ( .A(n6663), .B(n6664), .Z(n6662) );
  NAND U9467 ( .A(o[248]), .B(n5916), .Z(n6664) );
  NANDN U9468 ( .A(n5917), .B(creg[248]), .Z(n6663) );
  NAND U9469 ( .A(n6665), .B(n4555), .Z(n3352) );
  NANDN U9470 ( .A(init), .B(m[249]), .Z(n4555) );
  AND U9471 ( .A(n6666), .B(n6667), .Z(n6665) );
  NAND U9472 ( .A(o[249]), .B(n5916), .Z(n6667) );
  NANDN U9473 ( .A(n5917), .B(creg[249]), .Z(n6666) );
  NAND U9474 ( .A(n6668), .B(n4551), .Z(n3351) );
  NANDN U9475 ( .A(init), .B(m[250]), .Z(n4551) );
  AND U9476 ( .A(n6669), .B(n6670), .Z(n6668) );
  NAND U9477 ( .A(o[250]), .B(n5916), .Z(n6670) );
  NANDN U9478 ( .A(n5917), .B(creg[250]), .Z(n6669) );
  NAND U9479 ( .A(n6671), .B(n4549), .Z(n3350) );
  NANDN U9480 ( .A(init), .B(m[251]), .Z(n4549) );
  AND U9481 ( .A(n6672), .B(n6673), .Z(n6671) );
  NAND U9482 ( .A(o[251]), .B(n5916), .Z(n6673) );
  NANDN U9483 ( .A(n5917), .B(creg[251]), .Z(n6672) );
  NAND U9484 ( .A(n6674), .B(n4547), .Z(n3349) );
  NANDN U9485 ( .A(init), .B(m[252]), .Z(n4547) );
  AND U9486 ( .A(n6675), .B(n6676), .Z(n6674) );
  NAND U9487 ( .A(o[252]), .B(n5916), .Z(n6676) );
  NANDN U9488 ( .A(n5917), .B(creg[252]), .Z(n6675) );
  NAND U9489 ( .A(n6677), .B(n4545), .Z(n3348) );
  NANDN U9490 ( .A(init), .B(m[253]), .Z(n4545) );
  AND U9491 ( .A(n6678), .B(n6679), .Z(n6677) );
  NAND U9492 ( .A(o[253]), .B(n5916), .Z(n6679) );
  NANDN U9493 ( .A(n5917), .B(creg[253]), .Z(n6678) );
  NAND U9494 ( .A(n6680), .B(n4543), .Z(n3347) );
  NANDN U9495 ( .A(init), .B(m[254]), .Z(n4543) );
  AND U9496 ( .A(n6681), .B(n6682), .Z(n6680) );
  NAND U9497 ( .A(o[254]), .B(n5916), .Z(n6682) );
  AND U9498 ( .A(start_in[511]), .B(n5917), .Z(n5916) );
  NANDN U9499 ( .A(n5917), .B(creg[254]), .Z(n6681) );
  NAND U9500 ( .A(init), .B(n6683), .Z(n5917) );
  NAND U9501 ( .A(first_one), .B(n6684), .Z(n6683) );
  AND U9502 ( .A(start_reg[511]), .B(n6685), .Z(n6684) );
  NAND U9503 ( .A(n6686), .B(mul_pow), .Z(n6685) );
  NANDN U9504 ( .A(first_one), .B(n6687), .Z(n3346) );
  NAND U9505 ( .A(n6688), .B(ereg[255]), .Z(n6687) );
  AND U9506 ( .A(start_in[511]), .B(mul_pow), .Z(n6688) );
  AND U9507 ( .A(start_reg[511]), .B(init), .Z(start_in[511]) );
  NAND U9508 ( .A(n6689), .B(n6690), .Z(c[9]) );
  NAND U9509 ( .A(n6691), .B(o[9]), .Z(n6690) );
  NAND U9510 ( .A(n6686), .B(creg[9]), .Z(n6689) );
  NAND U9511 ( .A(n6692), .B(n6693), .Z(c[99]) );
  NAND U9512 ( .A(n6691), .B(o[99]), .Z(n6693) );
  NAND U9513 ( .A(n6686), .B(creg[99]), .Z(n6692) );
  NAND U9514 ( .A(n6694), .B(n6695), .Z(c[98]) );
  NAND U9515 ( .A(n6691), .B(o[98]), .Z(n6695) );
  NAND U9516 ( .A(n6686), .B(creg[98]), .Z(n6694) );
  NAND U9517 ( .A(n6696), .B(n6697), .Z(c[97]) );
  NAND U9518 ( .A(n6691), .B(o[97]), .Z(n6697) );
  NAND U9519 ( .A(n6686), .B(creg[97]), .Z(n6696) );
  NAND U9520 ( .A(n6698), .B(n6699), .Z(c[96]) );
  NAND U9521 ( .A(n6691), .B(o[96]), .Z(n6699) );
  NAND U9522 ( .A(n6686), .B(creg[96]), .Z(n6698) );
  NAND U9523 ( .A(n6700), .B(n6701), .Z(c[95]) );
  NAND U9524 ( .A(n6691), .B(o[95]), .Z(n6701) );
  NAND U9525 ( .A(n6686), .B(creg[95]), .Z(n6700) );
  NAND U9526 ( .A(n6702), .B(n6703), .Z(c[94]) );
  NAND U9527 ( .A(n6691), .B(o[94]), .Z(n6703) );
  NAND U9528 ( .A(n6686), .B(creg[94]), .Z(n6702) );
  NAND U9529 ( .A(n6704), .B(n6705), .Z(c[93]) );
  NAND U9530 ( .A(n6691), .B(o[93]), .Z(n6705) );
  NAND U9531 ( .A(n6686), .B(creg[93]), .Z(n6704) );
  NAND U9532 ( .A(n6706), .B(n6707), .Z(c[92]) );
  NAND U9533 ( .A(n6691), .B(o[92]), .Z(n6707) );
  NAND U9534 ( .A(n6686), .B(creg[92]), .Z(n6706) );
  NAND U9535 ( .A(n6708), .B(n6709), .Z(c[91]) );
  NAND U9536 ( .A(n6691), .B(o[91]), .Z(n6709) );
  NAND U9537 ( .A(n6686), .B(creg[91]), .Z(n6708) );
  NAND U9538 ( .A(n6710), .B(n6711), .Z(c[90]) );
  NAND U9539 ( .A(n6691), .B(o[90]), .Z(n6711) );
  NAND U9540 ( .A(n6686), .B(creg[90]), .Z(n6710) );
  NAND U9541 ( .A(n6712), .B(n6713), .Z(c[8]) );
  NAND U9542 ( .A(n6691), .B(o[8]), .Z(n6713) );
  NAND U9543 ( .A(n6686), .B(creg[8]), .Z(n6712) );
  NAND U9544 ( .A(n6714), .B(n6715), .Z(c[89]) );
  NAND U9545 ( .A(n6691), .B(o[89]), .Z(n6715) );
  NAND U9546 ( .A(n6686), .B(creg[89]), .Z(n6714) );
  NAND U9547 ( .A(n6716), .B(n6717), .Z(c[88]) );
  NAND U9548 ( .A(n6691), .B(o[88]), .Z(n6717) );
  NAND U9549 ( .A(n6686), .B(creg[88]), .Z(n6716) );
  NAND U9550 ( .A(n6718), .B(n6719), .Z(c[87]) );
  NAND U9551 ( .A(n6691), .B(o[87]), .Z(n6719) );
  NAND U9552 ( .A(n6686), .B(creg[87]), .Z(n6718) );
  NAND U9553 ( .A(n6720), .B(n6721), .Z(c[86]) );
  NAND U9554 ( .A(n6691), .B(o[86]), .Z(n6721) );
  NAND U9555 ( .A(n6686), .B(creg[86]), .Z(n6720) );
  NAND U9556 ( .A(n6722), .B(n6723), .Z(c[85]) );
  NAND U9557 ( .A(n6691), .B(o[85]), .Z(n6723) );
  NAND U9558 ( .A(n6686), .B(creg[85]), .Z(n6722) );
  NAND U9559 ( .A(n6724), .B(n6725), .Z(c[84]) );
  NAND U9560 ( .A(n6691), .B(o[84]), .Z(n6725) );
  NAND U9561 ( .A(n6686), .B(creg[84]), .Z(n6724) );
  NAND U9562 ( .A(n6726), .B(n6727), .Z(c[83]) );
  NAND U9563 ( .A(n6691), .B(o[83]), .Z(n6727) );
  NAND U9564 ( .A(n6686), .B(creg[83]), .Z(n6726) );
  NAND U9565 ( .A(n6728), .B(n6729), .Z(c[82]) );
  NAND U9566 ( .A(n6691), .B(o[82]), .Z(n6729) );
  NAND U9567 ( .A(n6686), .B(creg[82]), .Z(n6728) );
  NAND U9568 ( .A(n6730), .B(n6731), .Z(c[81]) );
  NAND U9569 ( .A(n6691), .B(o[81]), .Z(n6731) );
  NAND U9570 ( .A(n6686), .B(creg[81]), .Z(n6730) );
  NAND U9571 ( .A(n6732), .B(n6733), .Z(c[80]) );
  NAND U9572 ( .A(n6691), .B(o[80]), .Z(n6733) );
  NAND U9573 ( .A(n6686), .B(creg[80]), .Z(n6732) );
  NAND U9574 ( .A(n6734), .B(n6735), .Z(c[7]) );
  NAND U9575 ( .A(n6691), .B(o[7]), .Z(n6735) );
  NAND U9576 ( .A(n6686), .B(creg[7]), .Z(n6734) );
  NAND U9577 ( .A(n6736), .B(n6737), .Z(c[79]) );
  NAND U9578 ( .A(n6691), .B(o[79]), .Z(n6737) );
  NAND U9579 ( .A(n6686), .B(creg[79]), .Z(n6736) );
  NAND U9580 ( .A(n6738), .B(n6739), .Z(c[78]) );
  NAND U9581 ( .A(n6691), .B(o[78]), .Z(n6739) );
  NAND U9582 ( .A(n6686), .B(creg[78]), .Z(n6738) );
  NAND U9583 ( .A(n6740), .B(n6741), .Z(c[77]) );
  NAND U9584 ( .A(n6691), .B(o[77]), .Z(n6741) );
  NAND U9585 ( .A(n6686), .B(creg[77]), .Z(n6740) );
  NAND U9586 ( .A(n6742), .B(n6743), .Z(c[76]) );
  NAND U9587 ( .A(n6691), .B(o[76]), .Z(n6743) );
  NAND U9588 ( .A(n6686), .B(creg[76]), .Z(n6742) );
  NAND U9589 ( .A(n6744), .B(n6745), .Z(c[75]) );
  NAND U9590 ( .A(n6691), .B(o[75]), .Z(n6745) );
  NAND U9591 ( .A(n6686), .B(creg[75]), .Z(n6744) );
  NAND U9592 ( .A(n6746), .B(n6747), .Z(c[74]) );
  NAND U9593 ( .A(n6691), .B(o[74]), .Z(n6747) );
  NAND U9594 ( .A(n6686), .B(creg[74]), .Z(n6746) );
  NAND U9595 ( .A(n6748), .B(n6749), .Z(c[73]) );
  NAND U9596 ( .A(n6691), .B(o[73]), .Z(n6749) );
  NAND U9597 ( .A(n6686), .B(creg[73]), .Z(n6748) );
  NAND U9598 ( .A(n6750), .B(n6751), .Z(c[72]) );
  NAND U9599 ( .A(n6691), .B(o[72]), .Z(n6751) );
  NAND U9600 ( .A(n6686), .B(creg[72]), .Z(n6750) );
  NAND U9601 ( .A(n6752), .B(n6753), .Z(c[71]) );
  NAND U9602 ( .A(n6691), .B(o[71]), .Z(n6753) );
  NAND U9603 ( .A(n6686), .B(creg[71]), .Z(n6752) );
  NAND U9604 ( .A(n6754), .B(n6755), .Z(c[70]) );
  NAND U9605 ( .A(n6691), .B(o[70]), .Z(n6755) );
  NAND U9606 ( .A(n6686), .B(creg[70]), .Z(n6754) );
  NAND U9607 ( .A(n6756), .B(n6757), .Z(c[6]) );
  NAND U9608 ( .A(n6691), .B(o[6]), .Z(n6757) );
  NAND U9609 ( .A(n6686), .B(creg[6]), .Z(n6756) );
  NAND U9610 ( .A(n6758), .B(n6759), .Z(c[69]) );
  NAND U9611 ( .A(n6691), .B(o[69]), .Z(n6759) );
  NAND U9612 ( .A(n6686), .B(creg[69]), .Z(n6758) );
  NAND U9613 ( .A(n6760), .B(n6761), .Z(c[68]) );
  NAND U9614 ( .A(n6691), .B(o[68]), .Z(n6761) );
  NAND U9615 ( .A(n6686), .B(creg[68]), .Z(n6760) );
  NAND U9616 ( .A(n6762), .B(n6763), .Z(c[67]) );
  NAND U9617 ( .A(n6691), .B(o[67]), .Z(n6763) );
  NAND U9618 ( .A(n6686), .B(creg[67]), .Z(n6762) );
  NAND U9619 ( .A(n6764), .B(n6765), .Z(c[66]) );
  NAND U9620 ( .A(n6691), .B(o[66]), .Z(n6765) );
  NAND U9621 ( .A(n6686), .B(creg[66]), .Z(n6764) );
  NAND U9622 ( .A(n6766), .B(n6767), .Z(c[65]) );
  NAND U9623 ( .A(n6691), .B(o[65]), .Z(n6767) );
  NAND U9624 ( .A(n6686), .B(creg[65]), .Z(n6766) );
  NAND U9625 ( .A(n6768), .B(n6769), .Z(c[64]) );
  NAND U9626 ( .A(n6691), .B(o[64]), .Z(n6769) );
  NAND U9627 ( .A(n6686), .B(creg[64]), .Z(n6768) );
  NAND U9628 ( .A(n6770), .B(n6771), .Z(c[63]) );
  NAND U9629 ( .A(n6691), .B(o[63]), .Z(n6771) );
  NAND U9630 ( .A(n6686), .B(creg[63]), .Z(n6770) );
  NAND U9631 ( .A(n6772), .B(n6773), .Z(c[62]) );
  NAND U9632 ( .A(n6691), .B(o[62]), .Z(n6773) );
  NAND U9633 ( .A(n6686), .B(creg[62]), .Z(n6772) );
  NAND U9634 ( .A(n6774), .B(n6775), .Z(c[61]) );
  NAND U9635 ( .A(n6691), .B(o[61]), .Z(n6775) );
  NAND U9636 ( .A(n6686), .B(creg[61]), .Z(n6774) );
  NAND U9637 ( .A(n6776), .B(n6777), .Z(c[60]) );
  NAND U9638 ( .A(n6691), .B(o[60]), .Z(n6777) );
  NAND U9639 ( .A(n6686), .B(creg[60]), .Z(n6776) );
  NAND U9640 ( .A(n6778), .B(n6779), .Z(c[5]) );
  NAND U9641 ( .A(n6691), .B(o[5]), .Z(n6779) );
  NAND U9642 ( .A(n6686), .B(creg[5]), .Z(n6778) );
  NAND U9643 ( .A(n6780), .B(n6781), .Z(c[59]) );
  NAND U9644 ( .A(n6691), .B(o[59]), .Z(n6781) );
  NAND U9645 ( .A(n6686), .B(creg[59]), .Z(n6780) );
  NAND U9646 ( .A(n6782), .B(n6783), .Z(c[58]) );
  NAND U9647 ( .A(n6691), .B(o[58]), .Z(n6783) );
  NAND U9648 ( .A(n6686), .B(creg[58]), .Z(n6782) );
  NAND U9649 ( .A(n6784), .B(n6785), .Z(c[57]) );
  NAND U9650 ( .A(n6691), .B(o[57]), .Z(n6785) );
  NAND U9651 ( .A(n6686), .B(creg[57]), .Z(n6784) );
  NAND U9652 ( .A(n6786), .B(n6787), .Z(c[56]) );
  NAND U9653 ( .A(n6691), .B(o[56]), .Z(n6787) );
  NAND U9654 ( .A(n6686), .B(creg[56]), .Z(n6786) );
  NAND U9655 ( .A(n6788), .B(n6789), .Z(c[55]) );
  NAND U9656 ( .A(n6691), .B(o[55]), .Z(n6789) );
  NAND U9657 ( .A(n6686), .B(creg[55]), .Z(n6788) );
  NAND U9658 ( .A(n6790), .B(n6791), .Z(c[54]) );
  NAND U9659 ( .A(n6691), .B(o[54]), .Z(n6791) );
  NAND U9660 ( .A(n6686), .B(creg[54]), .Z(n6790) );
  NAND U9661 ( .A(n6792), .B(n6793), .Z(c[53]) );
  NAND U9662 ( .A(n6691), .B(o[53]), .Z(n6793) );
  NAND U9663 ( .A(n6686), .B(creg[53]), .Z(n6792) );
  NAND U9664 ( .A(n6794), .B(n6795), .Z(c[52]) );
  NAND U9665 ( .A(n6691), .B(o[52]), .Z(n6795) );
  NAND U9666 ( .A(n6686), .B(creg[52]), .Z(n6794) );
  NAND U9667 ( .A(n6796), .B(n6797), .Z(c[51]) );
  NAND U9668 ( .A(n6691), .B(o[51]), .Z(n6797) );
  NAND U9669 ( .A(n6686), .B(creg[51]), .Z(n6796) );
  NAND U9670 ( .A(n6798), .B(n6799), .Z(c[50]) );
  NAND U9671 ( .A(n6691), .B(o[50]), .Z(n6799) );
  NAND U9672 ( .A(n6686), .B(creg[50]), .Z(n6798) );
  NAND U9673 ( .A(n6800), .B(n6801), .Z(c[4]) );
  NAND U9674 ( .A(n6691), .B(o[4]), .Z(n6801) );
  NAND U9675 ( .A(n6686), .B(creg[4]), .Z(n6800) );
  NAND U9676 ( .A(n6802), .B(n6803), .Z(c[49]) );
  NAND U9677 ( .A(n6691), .B(o[49]), .Z(n6803) );
  NAND U9678 ( .A(n6686), .B(creg[49]), .Z(n6802) );
  NAND U9679 ( .A(n6804), .B(n6805), .Z(c[48]) );
  NAND U9680 ( .A(n6691), .B(o[48]), .Z(n6805) );
  NAND U9681 ( .A(n6686), .B(creg[48]), .Z(n6804) );
  NAND U9682 ( .A(n6806), .B(n6807), .Z(c[47]) );
  NAND U9683 ( .A(n6691), .B(o[47]), .Z(n6807) );
  NAND U9684 ( .A(n6686), .B(creg[47]), .Z(n6806) );
  NAND U9685 ( .A(n6808), .B(n6809), .Z(c[46]) );
  NAND U9686 ( .A(n6691), .B(o[46]), .Z(n6809) );
  NAND U9687 ( .A(n6686), .B(creg[46]), .Z(n6808) );
  NAND U9688 ( .A(n6810), .B(n6811), .Z(c[45]) );
  NAND U9689 ( .A(n6691), .B(o[45]), .Z(n6811) );
  NAND U9690 ( .A(n6686), .B(creg[45]), .Z(n6810) );
  NAND U9691 ( .A(n6812), .B(n6813), .Z(c[44]) );
  NAND U9692 ( .A(n6691), .B(o[44]), .Z(n6813) );
  NAND U9693 ( .A(n6686), .B(creg[44]), .Z(n6812) );
  NAND U9694 ( .A(n6814), .B(n6815), .Z(c[43]) );
  NAND U9695 ( .A(n6691), .B(o[43]), .Z(n6815) );
  NAND U9696 ( .A(n6686), .B(creg[43]), .Z(n6814) );
  NAND U9697 ( .A(n6816), .B(n6817), .Z(c[42]) );
  NAND U9698 ( .A(n6691), .B(o[42]), .Z(n6817) );
  NAND U9699 ( .A(n6686), .B(creg[42]), .Z(n6816) );
  NAND U9700 ( .A(n6818), .B(n6819), .Z(c[41]) );
  NAND U9701 ( .A(n6691), .B(o[41]), .Z(n6819) );
  NAND U9702 ( .A(n6686), .B(creg[41]), .Z(n6818) );
  NAND U9703 ( .A(n6820), .B(n6821), .Z(c[40]) );
  NAND U9704 ( .A(n6691), .B(o[40]), .Z(n6821) );
  NAND U9705 ( .A(n6686), .B(creg[40]), .Z(n6820) );
  NAND U9706 ( .A(n6822), .B(n6823), .Z(c[3]) );
  NAND U9707 ( .A(n6691), .B(o[3]), .Z(n6823) );
  NAND U9708 ( .A(n6686), .B(creg[3]), .Z(n6822) );
  NAND U9709 ( .A(n6824), .B(n6825), .Z(c[39]) );
  NAND U9710 ( .A(n6691), .B(o[39]), .Z(n6825) );
  NAND U9711 ( .A(n6686), .B(creg[39]), .Z(n6824) );
  NAND U9712 ( .A(n6826), .B(n6827), .Z(c[38]) );
  NAND U9713 ( .A(n6691), .B(o[38]), .Z(n6827) );
  NAND U9714 ( .A(n6686), .B(creg[38]), .Z(n6826) );
  NAND U9715 ( .A(n6828), .B(n6829), .Z(c[37]) );
  NAND U9716 ( .A(n6691), .B(o[37]), .Z(n6829) );
  NAND U9717 ( .A(n6686), .B(creg[37]), .Z(n6828) );
  NAND U9718 ( .A(n6830), .B(n6831), .Z(c[36]) );
  NAND U9719 ( .A(n6691), .B(o[36]), .Z(n6831) );
  NAND U9720 ( .A(n6686), .B(creg[36]), .Z(n6830) );
  NAND U9721 ( .A(n6832), .B(n6833), .Z(c[35]) );
  NAND U9722 ( .A(n6691), .B(o[35]), .Z(n6833) );
  NAND U9723 ( .A(n6686), .B(creg[35]), .Z(n6832) );
  NAND U9724 ( .A(n6834), .B(n6835), .Z(c[34]) );
  NAND U9725 ( .A(n6691), .B(o[34]), .Z(n6835) );
  NAND U9726 ( .A(n6686), .B(creg[34]), .Z(n6834) );
  NAND U9727 ( .A(n6836), .B(n6837), .Z(c[33]) );
  NAND U9728 ( .A(n6691), .B(o[33]), .Z(n6837) );
  NAND U9729 ( .A(n6686), .B(creg[33]), .Z(n6836) );
  NAND U9730 ( .A(n6838), .B(n6839), .Z(c[32]) );
  NAND U9731 ( .A(n6691), .B(o[32]), .Z(n6839) );
  NAND U9732 ( .A(n6686), .B(creg[32]), .Z(n6838) );
  NAND U9733 ( .A(n6840), .B(n6841), .Z(c[31]) );
  NAND U9734 ( .A(n6691), .B(o[31]), .Z(n6841) );
  NAND U9735 ( .A(n6686), .B(creg[31]), .Z(n6840) );
  NAND U9736 ( .A(n6842), .B(n6843), .Z(c[30]) );
  NAND U9737 ( .A(n6691), .B(o[30]), .Z(n6843) );
  NAND U9738 ( .A(n6686), .B(creg[30]), .Z(n6842) );
  NAND U9739 ( .A(n6844), .B(n6845), .Z(c[2]) );
  NAND U9740 ( .A(n6691), .B(o[2]), .Z(n6845) );
  NAND U9741 ( .A(n6686), .B(creg[2]), .Z(n6844) );
  NAND U9742 ( .A(n6846), .B(n6847), .Z(c[29]) );
  NAND U9743 ( .A(n6691), .B(o[29]), .Z(n6847) );
  NAND U9744 ( .A(n6686), .B(creg[29]), .Z(n6846) );
  NAND U9745 ( .A(n6848), .B(n6849), .Z(c[28]) );
  NAND U9746 ( .A(n6691), .B(o[28]), .Z(n6849) );
  NAND U9747 ( .A(n6686), .B(creg[28]), .Z(n6848) );
  NAND U9748 ( .A(n6850), .B(n6851), .Z(c[27]) );
  NAND U9749 ( .A(n6691), .B(o[27]), .Z(n6851) );
  NAND U9750 ( .A(n6686), .B(creg[27]), .Z(n6850) );
  NAND U9751 ( .A(n6852), .B(n6853), .Z(c[26]) );
  NAND U9752 ( .A(n6691), .B(o[26]), .Z(n6853) );
  NAND U9753 ( .A(n6686), .B(creg[26]), .Z(n6852) );
  NAND U9754 ( .A(n6854), .B(n6855), .Z(c[25]) );
  NAND U9755 ( .A(n6691), .B(o[25]), .Z(n6855) );
  NAND U9756 ( .A(n6686), .B(creg[25]), .Z(n6854) );
  NAND U9757 ( .A(n6856), .B(n6857), .Z(c[255]) );
  NAND U9758 ( .A(n6691), .B(o[255]), .Z(n6857) );
  NAND U9759 ( .A(n6686), .B(creg[255]), .Z(n6856) );
  NAND U9760 ( .A(n6858), .B(n6859), .Z(c[254]) );
  NAND U9761 ( .A(n6691), .B(o[254]), .Z(n6859) );
  NAND U9762 ( .A(n6686), .B(creg[254]), .Z(n6858) );
  NAND U9763 ( .A(n6860), .B(n6861), .Z(c[253]) );
  NAND U9764 ( .A(n6691), .B(o[253]), .Z(n6861) );
  NAND U9765 ( .A(n6686), .B(creg[253]), .Z(n6860) );
  NAND U9766 ( .A(n6862), .B(n6863), .Z(c[252]) );
  NAND U9767 ( .A(n6691), .B(o[252]), .Z(n6863) );
  NAND U9768 ( .A(n6686), .B(creg[252]), .Z(n6862) );
  NAND U9769 ( .A(n6864), .B(n6865), .Z(c[251]) );
  NAND U9770 ( .A(n6691), .B(o[251]), .Z(n6865) );
  NAND U9771 ( .A(n6686), .B(creg[251]), .Z(n6864) );
  NAND U9772 ( .A(n6866), .B(n6867), .Z(c[250]) );
  NAND U9773 ( .A(n6691), .B(o[250]), .Z(n6867) );
  NAND U9774 ( .A(n6686), .B(creg[250]), .Z(n6866) );
  NAND U9775 ( .A(n6868), .B(n6869), .Z(c[24]) );
  NAND U9776 ( .A(n6691), .B(o[24]), .Z(n6869) );
  NAND U9777 ( .A(n6686), .B(creg[24]), .Z(n6868) );
  NAND U9778 ( .A(n6870), .B(n6871), .Z(c[249]) );
  NAND U9779 ( .A(n6691), .B(o[249]), .Z(n6871) );
  NAND U9780 ( .A(n6686), .B(creg[249]), .Z(n6870) );
  NAND U9781 ( .A(n6872), .B(n6873), .Z(c[248]) );
  NAND U9782 ( .A(n6691), .B(o[248]), .Z(n6873) );
  NAND U9783 ( .A(n6686), .B(creg[248]), .Z(n6872) );
  NAND U9784 ( .A(n6874), .B(n6875), .Z(c[247]) );
  NAND U9785 ( .A(n6691), .B(o[247]), .Z(n6875) );
  NAND U9786 ( .A(n6686), .B(creg[247]), .Z(n6874) );
  NAND U9787 ( .A(n6876), .B(n6877), .Z(c[246]) );
  NAND U9788 ( .A(n6691), .B(o[246]), .Z(n6877) );
  NAND U9789 ( .A(n6686), .B(creg[246]), .Z(n6876) );
  NAND U9790 ( .A(n6878), .B(n6879), .Z(c[245]) );
  NAND U9791 ( .A(n6691), .B(o[245]), .Z(n6879) );
  NAND U9792 ( .A(n6686), .B(creg[245]), .Z(n6878) );
  NAND U9793 ( .A(n6880), .B(n6881), .Z(c[244]) );
  NAND U9794 ( .A(n6691), .B(o[244]), .Z(n6881) );
  NAND U9795 ( .A(n6686), .B(creg[244]), .Z(n6880) );
  NAND U9796 ( .A(n6882), .B(n6883), .Z(c[243]) );
  NAND U9797 ( .A(n6691), .B(o[243]), .Z(n6883) );
  NAND U9798 ( .A(n6686), .B(creg[243]), .Z(n6882) );
  NAND U9799 ( .A(n6884), .B(n6885), .Z(c[242]) );
  NAND U9800 ( .A(n6691), .B(o[242]), .Z(n6885) );
  NAND U9801 ( .A(n6686), .B(creg[242]), .Z(n6884) );
  NAND U9802 ( .A(n6886), .B(n6887), .Z(c[241]) );
  NAND U9803 ( .A(n6691), .B(o[241]), .Z(n6887) );
  NAND U9804 ( .A(n6686), .B(creg[241]), .Z(n6886) );
  NAND U9805 ( .A(n6888), .B(n6889), .Z(c[240]) );
  NAND U9806 ( .A(n6691), .B(o[240]), .Z(n6889) );
  NAND U9807 ( .A(n6686), .B(creg[240]), .Z(n6888) );
  NAND U9808 ( .A(n6890), .B(n6891), .Z(c[23]) );
  NAND U9809 ( .A(n6691), .B(o[23]), .Z(n6891) );
  NAND U9810 ( .A(n6686), .B(creg[23]), .Z(n6890) );
  NAND U9811 ( .A(n6892), .B(n6893), .Z(c[239]) );
  NAND U9812 ( .A(n6691), .B(o[239]), .Z(n6893) );
  NAND U9813 ( .A(n6686), .B(creg[239]), .Z(n6892) );
  NAND U9814 ( .A(n6894), .B(n6895), .Z(c[238]) );
  NAND U9815 ( .A(n6691), .B(o[238]), .Z(n6895) );
  NAND U9816 ( .A(n6686), .B(creg[238]), .Z(n6894) );
  NAND U9817 ( .A(n6896), .B(n6897), .Z(c[237]) );
  NAND U9818 ( .A(n6691), .B(o[237]), .Z(n6897) );
  NAND U9819 ( .A(n6686), .B(creg[237]), .Z(n6896) );
  NAND U9820 ( .A(n6898), .B(n6899), .Z(c[236]) );
  NAND U9821 ( .A(n6691), .B(o[236]), .Z(n6899) );
  NAND U9822 ( .A(n6686), .B(creg[236]), .Z(n6898) );
  NAND U9823 ( .A(n6900), .B(n6901), .Z(c[235]) );
  NAND U9824 ( .A(n6691), .B(o[235]), .Z(n6901) );
  NAND U9825 ( .A(n6686), .B(creg[235]), .Z(n6900) );
  NAND U9826 ( .A(n6902), .B(n6903), .Z(c[234]) );
  NAND U9827 ( .A(n6691), .B(o[234]), .Z(n6903) );
  NAND U9828 ( .A(n6686), .B(creg[234]), .Z(n6902) );
  NAND U9829 ( .A(n6904), .B(n6905), .Z(c[233]) );
  NAND U9830 ( .A(n6691), .B(o[233]), .Z(n6905) );
  NAND U9831 ( .A(n6686), .B(creg[233]), .Z(n6904) );
  NAND U9832 ( .A(n6906), .B(n6907), .Z(c[232]) );
  NAND U9833 ( .A(n6691), .B(o[232]), .Z(n6907) );
  NAND U9834 ( .A(n6686), .B(creg[232]), .Z(n6906) );
  NAND U9835 ( .A(n6908), .B(n6909), .Z(c[231]) );
  NAND U9836 ( .A(n6691), .B(o[231]), .Z(n6909) );
  NAND U9837 ( .A(n6686), .B(creg[231]), .Z(n6908) );
  NAND U9838 ( .A(n6910), .B(n6911), .Z(c[230]) );
  NAND U9839 ( .A(n6691), .B(o[230]), .Z(n6911) );
  NAND U9840 ( .A(n6686), .B(creg[230]), .Z(n6910) );
  NAND U9841 ( .A(n6912), .B(n6913), .Z(c[22]) );
  NAND U9842 ( .A(n6691), .B(o[22]), .Z(n6913) );
  NAND U9843 ( .A(n6686), .B(creg[22]), .Z(n6912) );
  NAND U9844 ( .A(n6914), .B(n6915), .Z(c[229]) );
  NAND U9845 ( .A(n6691), .B(o[229]), .Z(n6915) );
  NAND U9846 ( .A(n6686), .B(creg[229]), .Z(n6914) );
  NAND U9847 ( .A(n6916), .B(n6917), .Z(c[228]) );
  NAND U9848 ( .A(n6691), .B(o[228]), .Z(n6917) );
  NAND U9849 ( .A(n6686), .B(creg[228]), .Z(n6916) );
  NAND U9850 ( .A(n6918), .B(n6919), .Z(c[227]) );
  NAND U9851 ( .A(n6691), .B(o[227]), .Z(n6919) );
  NAND U9852 ( .A(n6686), .B(creg[227]), .Z(n6918) );
  NAND U9853 ( .A(n6920), .B(n6921), .Z(c[226]) );
  NAND U9854 ( .A(n6691), .B(o[226]), .Z(n6921) );
  NAND U9855 ( .A(n6686), .B(creg[226]), .Z(n6920) );
  NAND U9856 ( .A(n6922), .B(n6923), .Z(c[225]) );
  NAND U9857 ( .A(n6691), .B(o[225]), .Z(n6923) );
  NAND U9858 ( .A(n6686), .B(creg[225]), .Z(n6922) );
  NAND U9859 ( .A(n6924), .B(n6925), .Z(c[224]) );
  NAND U9860 ( .A(n6691), .B(o[224]), .Z(n6925) );
  NAND U9861 ( .A(n6686), .B(creg[224]), .Z(n6924) );
  NAND U9862 ( .A(n6926), .B(n6927), .Z(c[223]) );
  NAND U9863 ( .A(n6691), .B(o[223]), .Z(n6927) );
  NAND U9864 ( .A(n6686), .B(creg[223]), .Z(n6926) );
  NAND U9865 ( .A(n6928), .B(n6929), .Z(c[222]) );
  NAND U9866 ( .A(n6691), .B(o[222]), .Z(n6929) );
  NAND U9867 ( .A(n6686), .B(creg[222]), .Z(n6928) );
  NAND U9868 ( .A(n6930), .B(n6931), .Z(c[221]) );
  NAND U9869 ( .A(n6691), .B(o[221]), .Z(n6931) );
  NAND U9870 ( .A(n6686), .B(creg[221]), .Z(n6930) );
  NAND U9871 ( .A(n6932), .B(n6933), .Z(c[220]) );
  NAND U9872 ( .A(n6691), .B(o[220]), .Z(n6933) );
  NAND U9873 ( .A(n6686), .B(creg[220]), .Z(n6932) );
  NAND U9874 ( .A(n6934), .B(n6935), .Z(c[21]) );
  NAND U9875 ( .A(n6691), .B(o[21]), .Z(n6935) );
  NAND U9876 ( .A(n6686), .B(creg[21]), .Z(n6934) );
  NAND U9877 ( .A(n6936), .B(n6937), .Z(c[219]) );
  NAND U9878 ( .A(n6691), .B(o[219]), .Z(n6937) );
  NAND U9879 ( .A(n6686), .B(creg[219]), .Z(n6936) );
  NAND U9880 ( .A(n6938), .B(n6939), .Z(c[218]) );
  NAND U9881 ( .A(n6691), .B(o[218]), .Z(n6939) );
  NAND U9882 ( .A(n6686), .B(creg[218]), .Z(n6938) );
  NAND U9883 ( .A(n6940), .B(n6941), .Z(c[217]) );
  NAND U9884 ( .A(n6691), .B(o[217]), .Z(n6941) );
  NAND U9885 ( .A(n6686), .B(creg[217]), .Z(n6940) );
  NAND U9886 ( .A(n6942), .B(n6943), .Z(c[216]) );
  NAND U9887 ( .A(n6691), .B(o[216]), .Z(n6943) );
  NAND U9888 ( .A(n6686), .B(creg[216]), .Z(n6942) );
  NAND U9889 ( .A(n6944), .B(n6945), .Z(c[215]) );
  NAND U9890 ( .A(n6691), .B(o[215]), .Z(n6945) );
  NAND U9891 ( .A(n6686), .B(creg[215]), .Z(n6944) );
  NAND U9892 ( .A(n6946), .B(n6947), .Z(c[214]) );
  NAND U9893 ( .A(n6691), .B(o[214]), .Z(n6947) );
  NAND U9894 ( .A(n6686), .B(creg[214]), .Z(n6946) );
  NAND U9895 ( .A(n6948), .B(n6949), .Z(c[213]) );
  NAND U9896 ( .A(n6691), .B(o[213]), .Z(n6949) );
  NAND U9897 ( .A(n6686), .B(creg[213]), .Z(n6948) );
  NAND U9898 ( .A(n6950), .B(n6951), .Z(c[212]) );
  NAND U9899 ( .A(n6691), .B(o[212]), .Z(n6951) );
  NAND U9900 ( .A(n6686), .B(creg[212]), .Z(n6950) );
  NAND U9901 ( .A(n6952), .B(n6953), .Z(c[211]) );
  NAND U9902 ( .A(n6691), .B(o[211]), .Z(n6953) );
  NAND U9903 ( .A(n6686), .B(creg[211]), .Z(n6952) );
  NAND U9904 ( .A(n6954), .B(n6955), .Z(c[210]) );
  NAND U9905 ( .A(n6691), .B(o[210]), .Z(n6955) );
  NAND U9906 ( .A(n6686), .B(creg[210]), .Z(n6954) );
  NAND U9907 ( .A(n6956), .B(n6957), .Z(c[20]) );
  NAND U9908 ( .A(n6691), .B(o[20]), .Z(n6957) );
  NAND U9909 ( .A(n6686), .B(creg[20]), .Z(n6956) );
  NAND U9910 ( .A(n6958), .B(n6959), .Z(c[209]) );
  NAND U9911 ( .A(n6691), .B(o[209]), .Z(n6959) );
  NAND U9912 ( .A(n6686), .B(creg[209]), .Z(n6958) );
  NAND U9913 ( .A(n6960), .B(n6961), .Z(c[208]) );
  NAND U9914 ( .A(n6691), .B(o[208]), .Z(n6961) );
  NAND U9915 ( .A(n6686), .B(creg[208]), .Z(n6960) );
  NAND U9916 ( .A(n6962), .B(n6963), .Z(c[207]) );
  NAND U9917 ( .A(n6691), .B(o[207]), .Z(n6963) );
  NAND U9918 ( .A(n6686), .B(creg[207]), .Z(n6962) );
  NAND U9919 ( .A(n6964), .B(n6965), .Z(c[206]) );
  NAND U9920 ( .A(n6691), .B(o[206]), .Z(n6965) );
  NAND U9921 ( .A(n6686), .B(creg[206]), .Z(n6964) );
  NAND U9922 ( .A(n6966), .B(n6967), .Z(c[205]) );
  NAND U9923 ( .A(n6691), .B(o[205]), .Z(n6967) );
  NAND U9924 ( .A(n6686), .B(creg[205]), .Z(n6966) );
  NAND U9925 ( .A(n6968), .B(n6969), .Z(c[204]) );
  NAND U9926 ( .A(n6691), .B(o[204]), .Z(n6969) );
  NAND U9927 ( .A(n6686), .B(creg[204]), .Z(n6968) );
  NAND U9928 ( .A(n6970), .B(n6971), .Z(c[203]) );
  NAND U9929 ( .A(n6691), .B(o[203]), .Z(n6971) );
  NAND U9930 ( .A(n6686), .B(creg[203]), .Z(n6970) );
  NAND U9931 ( .A(n6972), .B(n6973), .Z(c[202]) );
  NAND U9932 ( .A(n6691), .B(o[202]), .Z(n6973) );
  NAND U9933 ( .A(n6686), .B(creg[202]), .Z(n6972) );
  NAND U9934 ( .A(n6974), .B(n6975), .Z(c[201]) );
  NAND U9935 ( .A(n6691), .B(o[201]), .Z(n6975) );
  NAND U9936 ( .A(n6686), .B(creg[201]), .Z(n6974) );
  NAND U9937 ( .A(n6976), .B(n6977), .Z(c[200]) );
  NAND U9938 ( .A(n6691), .B(o[200]), .Z(n6977) );
  NAND U9939 ( .A(n6686), .B(creg[200]), .Z(n6976) );
  NAND U9940 ( .A(n6978), .B(n6979), .Z(c[1]) );
  NAND U9941 ( .A(n6691), .B(o[1]), .Z(n6979) );
  NAND U9942 ( .A(n6686), .B(creg[1]), .Z(n6978) );
  NAND U9943 ( .A(n6980), .B(n6981), .Z(c[19]) );
  NAND U9944 ( .A(n6691), .B(o[19]), .Z(n6981) );
  NAND U9945 ( .A(n6686), .B(creg[19]), .Z(n6980) );
  NAND U9946 ( .A(n6982), .B(n6983), .Z(c[199]) );
  NAND U9947 ( .A(n6691), .B(o[199]), .Z(n6983) );
  NAND U9948 ( .A(n6686), .B(creg[199]), .Z(n6982) );
  NAND U9949 ( .A(n6984), .B(n6985), .Z(c[198]) );
  NAND U9950 ( .A(n6691), .B(o[198]), .Z(n6985) );
  NAND U9951 ( .A(n6686), .B(creg[198]), .Z(n6984) );
  NAND U9952 ( .A(n6986), .B(n6987), .Z(c[197]) );
  NAND U9953 ( .A(n6691), .B(o[197]), .Z(n6987) );
  NAND U9954 ( .A(n6686), .B(creg[197]), .Z(n6986) );
  NAND U9955 ( .A(n6988), .B(n6989), .Z(c[196]) );
  NAND U9956 ( .A(n6691), .B(o[196]), .Z(n6989) );
  NAND U9957 ( .A(n6686), .B(creg[196]), .Z(n6988) );
  NAND U9958 ( .A(n6990), .B(n6991), .Z(c[195]) );
  NAND U9959 ( .A(n6691), .B(o[195]), .Z(n6991) );
  NAND U9960 ( .A(n6686), .B(creg[195]), .Z(n6990) );
  NAND U9961 ( .A(n6992), .B(n6993), .Z(c[194]) );
  NAND U9962 ( .A(n6691), .B(o[194]), .Z(n6993) );
  NAND U9963 ( .A(n6686), .B(creg[194]), .Z(n6992) );
  NAND U9964 ( .A(n6994), .B(n6995), .Z(c[193]) );
  NAND U9965 ( .A(n6691), .B(o[193]), .Z(n6995) );
  NAND U9966 ( .A(n6686), .B(creg[193]), .Z(n6994) );
  NAND U9967 ( .A(n6996), .B(n6997), .Z(c[192]) );
  NAND U9968 ( .A(n6691), .B(o[192]), .Z(n6997) );
  NAND U9969 ( .A(n6686), .B(creg[192]), .Z(n6996) );
  NAND U9970 ( .A(n6998), .B(n6999), .Z(c[191]) );
  NAND U9971 ( .A(n6691), .B(o[191]), .Z(n6999) );
  NAND U9972 ( .A(n6686), .B(creg[191]), .Z(n6998) );
  NAND U9973 ( .A(n7000), .B(n7001), .Z(c[190]) );
  NAND U9974 ( .A(n6691), .B(o[190]), .Z(n7001) );
  NAND U9975 ( .A(n6686), .B(creg[190]), .Z(n7000) );
  NAND U9976 ( .A(n7002), .B(n7003), .Z(c[18]) );
  NAND U9977 ( .A(n6691), .B(o[18]), .Z(n7003) );
  NAND U9978 ( .A(n6686), .B(creg[18]), .Z(n7002) );
  NAND U9979 ( .A(n7004), .B(n7005), .Z(c[189]) );
  NAND U9980 ( .A(n6691), .B(o[189]), .Z(n7005) );
  NAND U9981 ( .A(n6686), .B(creg[189]), .Z(n7004) );
  NAND U9982 ( .A(n7006), .B(n7007), .Z(c[188]) );
  NAND U9983 ( .A(n6691), .B(o[188]), .Z(n7007) );
  NAND U9984 ( .A(n6686), .B(creg[188]), .Z(n7006) );
  NAND U9985 ( .A(n7008), .B(n7009), .Z(c[187]) );
  NAND U9986 ( .A(n6691), .B(o[187]), .Z(n7009) );
  NAND U9987 ( .A(n6686), .B(creg[187]), .Z(n7008) );
  NAND U9988 ( .A(n7010), .B(n7011), .Z(c[186]) );
  NAND U9989 ( .A(n6691), .B(o[186]), .Z(n7011) );
  NAND U9990 ( .A(n6686), .B(creg[186]), .Z(n7010) );
  NAND U9991 ( .A(n7012), .B(n7013), .Z(c[185]) );
  NAND U9992 ( .A(n6691), .B(o[185]), .Z(n7013) );
  NAND U9993 ( .A(n6686), .B(creg[185]), .Z(n7012) );
  NAND U9994 ( .A(n7014), .B(n7015), .Z(c[184]) );
  NAND U9995 ( .A(n6691), .B(o[184]), .Z(n7015) );
  NAND U9996 ( .A(n6686), .B(creg[184]), .Z(n7014) );
  NAND U9997 ( .A(n7016), .B(n7017), .Z(c[183]) );
  NAND U9998 ( .A(n6691), .B(o[183]), .Z(n7017) );
  NAND U9999 ( .A(n6686), .B(creg[183]), .Z(n7016) );
  NAND U10000 ( .A(n7018), .B(n7019), .Z(c[182]) );
  NAND U10001 ( .A(n6691), .B(o[182]), .Z(n7019) );
  NAND U10002 ( .A(n6686), .B(creg[182]), .Z(n7018) );
  NAND U10003 ( .A(n7020), .B(n7021), .Z(c[181]) );
  NAND U10004 ( .A(n6691), .B(o[181]), .Z(n7021) );
  NAND U10005 ( .A(n6686), .B(creg[181]), .Z(n7020) );
  NAND U10006 ( .A(n7022), .B(n7023), .Z(c[180]) );
  NAND U10007 ( .A(n6691), .B(o[180]), .Z(n7023) );
  NAND U10008 ( .A(n6686), .B(creg[180]), .Z(n7022) );
  NAND U10009 ( .A(n7024), .B(n7025), .Z(c[17]) );
  NAND U10010 ( .A(n6691), .B(o[17]), .Z(n7025) );
  NAND U10011 ( .A(n6686), .B(creg[17]), .Z(n7024) );
  NAND U10012 ( .A(n7026), .B(n7027), .Z(c[179]) );
  NAND U10013 ( .A(n6691), .B(o[179]), .Z(n7027) );
  NAND U10014 ( .A(n6686), .B(creg[179]), .Z(n7026) );
  NAND U10015 ( .A(n7028), .B(n7029), .Z(c[178]) );
  NAND U10016 ( .A(n6691), .B(o[178]), .Z(n7029) );
  NAND U10017 ( .A(n6686), .B(creg[178]), .Z(n7028) );
  NAND U10018 ( .A(n7030), .B(n7031), .Z(c[177]) );
  NAND U10019 ( .A(n6691), .B(o[177]), .Z(n7031) );
  NAND U10020 ( .A(n6686), .B(creg[177]), .Z(n7030) );
  NAND U10021 ( .A(n7032), .B(n7033), .Z(c[176]) );
  NAND U10022 ( .A(n6691), .B(o[176]), .Z(n7033) );
  NAND U10023 ( .A(n6686), .B(creg[176]), .Z(n7032) );
  NAND U10024 ( .A(n7034), .B(n7035), .Z(c[175]) );
  NAND U10025 ( .A(n6691), .B(o[175]), .Z(n7035) );
  NAND U10026 ( .A(n6686), .B(creg[175]), .Z(n7034) );
  NAND U10027 ( .A(n7036), .B(n7037), .Z(c[174]) );
  NAND U10028 ( .A(n6691), .B(o[174]), .Z(n7037) );
  NAND U10029 ( .A(n6686), .B(creg[174]), .Z(n7036) );
  NAND U10030 ( .A(n7038), .B(n7039), .Z(c[173]) );
  NAND U10031 ( .A(n6691), .B(o[173]), .Z(n7039) );
  NAND U10032 ( .A(n6686), .B(creg[173]), .Z(n7038) );
  NAND U10033 ( .A(n7040), .B(n7041), .Z(c[172]) );
  NAND U10034 ( .A(n6691), .B(o[172]), .Z(n7041) );
  NAND U10035 ( .A(n6686), .B(creg[172]), .Z(n7040) );
  NAND U10036 ( .A(n7042), .B(n7043), .Z(c[171]) );
  NAND U10037 ( .A(n6691), .B(o[171]), .Z(n7043) );
  NAND U10038 ( .A(n6686), .B(creg[171]), .Z(n7042) );
  NAND U10039 ( .A(n7044), .B(n7045), .Z(c[170]) );
  NAND U10040 ( .A(n6691), .B(o[170]), .Z(n7045) );
  NAND U10041 ( .A(n6686), .B(creg[170]), .Z(n7044) );
  NAND U10042 ( .A(n7046), .B(n7047), .Z(c[16]) );
  NAND U10043 ( .A(n6691), .B(o[16]), .Z(n7047) );
  NAND U10044 ( .A(n6686), .B(creg[16]), .Z(n7046) );
  NAND U10045 ( .A(n7048), .B(n7049), .Z(c[169]) );
  NAND U10046 ( .A(n6691), .B(o[169]), .Z(n7049) );
  NAND U10047 ( .A(n6686), .B(creg[169]), .Z(n7048) );
  NAND U10048 ( .A(n7050), .B(n7051), .Z(c[168]) );
  NAND U10049 ( .A(n6691), .B(o[168]), .Z(n7051) );
  NAND U10050 ( .A(n6686), .B(creg[168]), .Z(n7050) );
  NAND U10051 ( .A(n7052), .B(n7053), .Z(c[167]) );
  NAND U10052 ( .A(n6691), .B(o[167]), .Z(n7053) );
  NAND U10053 ( .A(n6686), .B(creg[167]), .Z(n7052) );
  NAND U10054 ( .A(n7054), .B(n7055), .Z(c[166]) );
  NAND U10055 ( .A(n6691), .B(o[166]), .Z(n7055) );
  NAND U10056 ( .A(n6686), .B(creg[166]), .Z(n7054) );
  NAND U10057 ( .A(n7056), .B(n7057), .Z(c[165]) );
  NAND U10058 ( .A(n6691), .B(o[165]), .Z(n7057) );
  NAND U10059 ( .A(n6686), .B(creg[165]), .Z(n7056) );
  NAND U10060 ( .A(n7058), .B(n7059), .Z(c[164]) );
  NAND U10061 ( .A(n6691), .B(o[164]), .Z(n7059) );
  NAND U10062 ( .A(n6686), .B(creg[164]), .Z(n7058) );
  NAND U10063 ( .A(n7060), .B(n7061), .Z(c[163]) );
  NAND U10064 ( .A(n6691), .B(o[163]), .Z(n7061) );
  NAND U10065 ( .A(n6686), .B(creg[163]), .Z(n7060) );
  NAND U10066 ( .A(n7062), .B(n7063), .Z(c[162]) );
  NAND U10067 ( .A(n6691), .B(o[162]), .Z(n7063) );
  NAND U10068 ( .A(n6686), .B(creg[162]), .Z(n7062) );
  NAND U10069 ( .A(n7064), .B(n7065), .Z(c[161]) );
  NAND U10070 ( .A(n6691), .B(o[161]), .Z(n7065) );
  NAND U10071 ( .A(n6686), .B(creg[161]), .Z(n7064) );
  NAND U10072 ( .A(n7066), .B(n7067), .Z(c[160]) );
  NAND U10073 ( .A(n6691), .B(o[160]), .Z(n7067) );
  NAND U10074 ( .A(n6686), .B(creg[160]), .Z(n7066) );
  NAND U10075 ( .A(n7068), .B(n7069), .Z(c[15]) );
  NAND U10076 ( .A(n6691), .B(o[15]), .Z(n7069) );
  NAND U10077 ( .A(n6686), .B(creg[15]), .Z(n7068) );
  NAND U10078 ( .A(n7070), .B(n7071), .Z(c[159]) );
  NAND U10079 ( .A(n6691), .B(o[159]), .Z(n7071) );
  NAND U10080 ( .A(n6686), .B(creg[159]), .Z(n7070) );
  NAND U10081 ( .A(n7072), .B(n7073), .Z(c[158]) );
  NAND U10082 ( .A(n6691), .B(o[158]), .Z(n7073) );
  NAND U10083 ( .A(n6686), .B(creg[158]), .Z(n7072) );
  NAND U10084 ( .A(n7074), .B(n7075), .Z(c[157]) );
  NAND U10085 ( .A(n6691), .B(o[157]), .Z(n7075) );
  NAND U10086 ( .A(n6686), .B(creg[157]), .Z(n7074) );
  NAND U10087 ( .A(n7076), .B(n7077), .Z(c[156]) );
  NAND U10088 ( .A(n6691), .B(o[156]), .Z(n7077) );
  NAND U10089 ( .A(n6686), .B(creg[156]), .Z(n7076) );
  NAND U10090 ( .A(n7078), .B(n7079), .Z(c[155]) );
  NAND U10091 ( .A(n6691), .B(o[155]), .Z(n7079) );
  NAND U10092 ( .A(n6686), .B(creg[155]), .Z(n7078) );
  NAND U10093 ( .A(n7080), .B(n7081), .Z(c[154]) );
  NAND U10094 ( .A(n6691), .B(o[154]), .Z(n7081) );
  NAND U10095 ( .A(n6686), .B(creg[154]), .Z(n7080) );
  NAND U10096 ( .A(n7082), .B(n7083), .Z(c[153]) );
  NAND U10097 ( .A(n6691), .B(o[153]), .Z(n7083) );
  NAND U10098 ( .A(n6686), .B(creg[153]), .Z(n7082) );
  NAND U10099 ( .A(n7084), .B(n7085), .Z(c[152]) );
  NAND U10100 ( .A(n6691), .B(o[152]), .Z(n7085) );
  NAND U10101 ( .A(n6686), .B(creg[152]), .Z(n7084) );
  NAND U10102 ( .A(n7086), .B(n7087), .Z(c[151]) );
  NAND U10103 ( .A(n6691), .B(o[151]), .Z(n7087) );
  NAND U10104 ( .A(n6686), .B(creg[151]), .Z(n7086) );
  NAND U10105 ( .A(n7088), .B(n7089), .Z(c[150]) );
  NAND U10106 ( .A(n6691), .B(o[150]), .Z(n7089) );
  NAND U10107 ( .A(n6686), .B(creg[150]), .Z(n7088) );
  NAND U10108 ( .A(n7090), .B(n7091), .Z(c[14]) );
  NAND U10109 ( .A(n6691), .B(o[14]), .Z(n7091) );
  NAND U10110 ( .A(n6686), .B(creg[14]), .Z(n7090) );
  NAND U10111 ( .A(n7092), .B(n7093), .Z(c[149]) );
  NAND U10112 ( .A(n6691), .B(o[149]), .Z(n7093) );
  NAND U10113 ( .A(n6686), .B(creg[149]), .Z(n7092) );
  NAND U10114 ( .A(n7094), .B(n7095), .Z(c[148]) );
  NAND U10115 ( .A(n6691), .B(o[148]), .Z(n7095) );
  NAND U10116 ( .A(n6686), .B(creg[148]), .Z(n7094) );
  NAND U10117 ( .A(n7096), .B(n7097), .Z(c[147]) );
  NAND U10118 ( .A(n6691), .B(o[147]), .Z(n7097) );
  NAND U10119 ( .A(n6686), .B(creg[147]), .Z(n7096) );
  NAND U10120 ( .A(n7098), .B(n7099), .Z(c[146]) );
  NAND U10121 ( .A(n6691), .B(o[146]), .Z(n7099) );
  NAND U10122 ( .A(n6686), .B(creg[146]), .Z(n7098) );
  NAND U10123 ( .A(n7100), .B(n7101), .Z(c[145]) );
  NAND U10124 ( .A(n6691), .B(o[145]), .Z(n7101) );
  NAND U10125 ( .A(n6686), .B(creg[145]), .Z(n7100) );
  NAND U10126 ( .A(n7102), .B(n7103), .Z(c[144]) );
  NAND U10127 ( .A(n6691), .B(o[144]), .Z(n7103) );
  NAND U10128 ( .A(n6686), .B(creg[144]), .Z(n7102) );
  NAND U10129 ( .A(n7104), .B(n7105), .Z(c[143]) );
  NAND U10130 ( .A(n6691), .B(o[143]), .Z(n7105) );
  NAND U10131 ( .A(n6686), .B(creg[143]), .Z(n7104) );
  NAND U10132 ( .A(n7106), .B(n7107), .Z(c[142]) );
  NAND U10133 ( .A(n6691), .B(o[142]), .Z(n7107) );
  NAND U10134 ( .A(n6686), .B(creg[142]), .Z(n7106) );
  NAND U10135 ( .A(n7108), .B(n7109), .Z(c[141]) );
  NAND U10136 ( .A(n6691), .B(o[141]), .Z(n7109) );
  NAND U10137 ( .A(n6686), .B(creg[141]), .Z(n7108) );
  NAND U10138 ( .A(n7110), .B(n7111), .Z(c[140]) );
  NAND U10139 ( .A(n6691), .B(o[140]), .Z(n7111) );
  NAND U10140 ( .A(n6686), .B(creg[140]), .Z(n7110) );
  NAND U10141 ( .A(n7112), .B(n7113), .Z(c[13]) );
  NAND U10142 ( .A(n6691), .B(o[13]), .Z(n7113) );
  NAND U10143 ( .A(n6686), .B(creg[13]), .Z(n7112) );
  NAND U10144 ( .A(n7114), .B(n7115), .Z(c[139]) );
  NAND U10145 ( .A(n6691), .B(o[139]), .Z(n7115) );
  NAND U10146 ( .A(n6686), .B(creg[139]), .Z(n7114) );
  NAND U10147 ( .A(n7116), .B(n7117), .Z(c[138]) );
  NAND U10148 ( .A(n6691), .B(o[138]), .Z(n7117) );
  NAND U10149 ( .A(n6686), .B(creg[138]), .Z(n7116) );
  NAND U10150 ( .A(n7118), .B(n7119), .Z(c[137]) );
  NAND U10151 ( .A(n6691), .B(o[137]), .Z(n7119) );
  NAND U10152 ( .A(n6686), .B(creg[137]), .Z(n7118) );
  NAND U10153 ( .A(n7120), .B(n7121), .Z(c[136]) );
  NAND U10154 ( .A(n6691), .B(o[136]), .Z(n7121) );
  NAND U10155 ( .A(n6686), .B(creg[136]), .Z(n7120) );
  NAND U10156 ( .A(n7122), .B(n7123), .Z(c[135]) );
  NAND U10157 ( .A(n6691), .B(o[135]), .Z(n7123) );
  NAND U10158 ( .A(n6686), .B(creg[135]), .Z(n7122) );
  NAND U10159 ( .A(n7124), .B(n7125), .Z(c[134]) );
  NAND U10160 ( .A(n6691), .B(o[134]), .Z(n7125) );
  NAND U10161 ( .A(n6686), .B(creg[134]), .Z(n7124) );
  NAND U10162 ( .A(n7126), .B(n7127), .Z(c[133]) );
  NAND U10163 ( .A(n6691), .B(o[133]), .Z(n7127) );
  NAND U10164 ( .A(n6686), .B(creg[133]), .Z(n7126) );
  NAND U10165 ( .A(n7128), .B(n7129), .Z(c[132]) );
  NAND U10166 ( .A(n6691), .B(o[132]), .Z(n7129) );
  NAND U10167 ( .A(n6686), .B(creg[132]), .Z(n7128) );
  NAND U10168 ( .A(n7130), .B(n7131), .Z(c[131]) );
  NAND U10169 ( .A(n6691), .B(o[131]), .Z(n7131) );
  NAND U10170 ( .A(n6686), .B(creg[131]), .Z(n7130) );
  NAND U10171 ( .A(n7132), .B(n7133), .Z(c[130]) );
  NAND U10172 ( .A(n6691), .B(o[130]), .Z(n7133) );
  NAND U10173 ( .A(n6686), .B(creg[130]), .Z(n7132) );
  NAND U10174 ( .A(n7134), .B(n7135), .Z(c[12]) );
  NAND U10175 ( .A(n6691), .B(o[12]), .Z(n7135) );
  NAND U10176 ( .A(n6686), .B(creg[12]), .Z(n7134) );
  NAND U10177 ( .A(n7136), .B(n7137), .Z(c[129]) );
  NAND U10178 ( .A(n6691), .B(o[129]), .Z(n7137) );
  NAND U10179 ( .A(n6686), .B(creg[129]), .Z(n7136) );
  NAND U10180 ( .A(n7138), .B(n7139), .Z(c[128]) );
  NAND U10181 ( .A(n6691), .B(o[128]), .Z(n7139) );
  NAND U10182 ( .A(n6686), .B(creg[128]), .Z(n7138) );
  NAND U10183 ( .A(n7140), .B(n7141), .Z(c[127]) );
  NAND U10184 ( .A(n6691), .B(o[127]), .Z(n7141) );
  NAND U10185 ( .A(n6686), .B(creg[127]), .Z(n7140) );
  NAND U10186 ( .A(n7142), .B(n7143), .Z(c[126]) );
  NAND U10187 ( .A(n6691), .B(o[126]), .Z(n7143) );
  NAND U10188 ( .A(n6686), .B(creg[126]), .Z(n7142) );
  NAND U10189 ( .A(n7144), .B(n7145), .Z(c[125]) );
  NAND U10190 ( .A(n6691), .B(o[125]), .Z(n7145) );
  NAND U10191 ( .A(n6686), .B(creg[125]), .Z(n7144) );
  NAND U10192 ( .A(n7146), .B(n7147), .Z(c[124]) );
  NAND U10193 ( .A(n6691), .B(o[124]), .Z(n7147) );
  NAND U10194 ( .A(n6686), .B(creg[124]), .Z(n7146) );
  NAND U10195 ( .A(n7148), .B(n7149), .Z(c[123]) );
  NAND U10196 ( .A(n6691), .B(o[123]), .Z(n7149) );
  NAND U10197 ( .A(n6686), .B(creg[123]), .Z(n7148) );
  NAND U10198 ( .A(n7150), .B(n7151), .Z(c[122]) );
  NAND U10199 ( .A(n6691), .B(o[122]), .Z(n7151) );
  NAND U10200 ( .A(n6686), .B(creg[122]), .Z(n7150) );
  NAND U10201 ( .A(n7152), .B(n7153), .Z(c[121]) );
  NAND U10202 ( .A(n6691), .B(o[121]), .Z(n7153) );
  NAND U10203 ( .A(n6686), .B(creg[121]), .Z(n7152) );
  NAND U10204 ( .A(n7154), .B(n7155), .Z(c[120]) );
  NAND U10205 ( .A(n6691), .B(o[120]), .Z(n7155) );
  NAND U10206 ( .A(n6686), .B(creg[120]), .Z(n7154) );
  NAND U10207 ( .A(n7156), .B(n7157), .Z(c[11]) );
  NAND U10208 ( .A(n6691), .B(o[11]), .Z(n7157) );
  NAND U10209 ( .A(n6686), .B(creg[11]), .Z(n7156) );
  NAND U10210 ( .A(n7158), .B(n7159), .Z(c[119]) );
  NAND U10211 ( .A(n6691), .B(o[119]), .Z(n7159) );
  NAND U10212 ( .A(n6686), .B(creg[119]), .Z(n7158) );
  NAND U10213 ( .A(n7160), .B(n7161), .Z(c[118]) );
  NAND U10214 ( .A(n6691), .B(o[118]), .Z(n7161) );
  NAND U10215 ( .A(n6686), .B(creg[118]), .Z(n7160) );
  NAND U10216 ( .A(n7162), .B(n7163), .Z(c[117]) );
  NAND U10217 ( .A(n6691), .B(o[117]), .Z(n7163) );
  NAND U10218 ( .A(n6686), .B(creg[117]), .Z(n7162) );
  NAND U10219 ( .A(n7164), .B(n7165), .Z(c[116]) );
  NAND U10220 ( .A(n6691), .B(o[116]), .Z(n7165) );
  NAND U10221 ( .A(n6686), .B(creg[116]), .Z(n7164) );
  NAND U10222 ( .A(n7166), .B(n7167), .Z(c[115]) );
  NAND U10223 ( .A(n6691), .B(o[115]), .Z(n7167) );
  NAND U10224 ( .A(n6686), .B(creg[115]), .Z(n7166) );
  NAND U10225 ( .A(n7168), .B(n7169), .Z(c[114]) );
  NAND U10226 ( .A(n6691), .B(o[114]), .Z(n7169) );
  NAND U10227 ( .A(n6686), .B(creg[114]), .Z(n7168) );
  NAND U10228 ( .A(n7170), .B(n7171), .Z(c[113]) );
  NAND U10229 ( .A(n6691), .B(o[113]), .Z(n7171) );
  NAND U10230 ( .A(n6686), .B(creg[113]), .Z(n7170) );
  NAND U10231 ( .A(n7172), .B(n7173), .Z(c[112]) );
  NAND U10232 ( .A(n6691), .B(o[112]), .Z(n7173) );
  NAND U10233 ( .A(n6686), .B(creg[112]), .Z(n7172) );
  NAND U10234 ( .A(n7174), .B(n7175), .Z(c[111]) );
  NAND U10235 ( .A(n6691), .B(o[111]), .Z(n7175) );
  NAND U10236 ( .A(n6686), .B(creg[111]), .Z(n7174) );
  NAND U10237 ( .A(n7176), .B(n7177), .Z(c[110]) );
  NAND U10238 ( .A(n6691), .B(o[110]), .Z(n7177) );
  NAND U10239 ( .A(n6686), .B(creg[110]), .Z(n7176) );
  NAND U10240 ( .A(n7178), .B(n7179), .Z(c[10]) );
  NAND U10241 ( .A(n6691), .B(o[10]), .Z(n7179) );
  NAND U10242 ( .A(n6686), .B(creg[10]), .Z(n7178) );
  NAND U10243 ( .A(n7180), .B(n7181), .Z(c[109]) );
  NAND U10244 ( .A(n6691), .B(o[109]), .Z(n7181) );
  NAND U10245 ( .A(n6686), .B(creg[109]), .Z(n7180) );
  NAND U10246 ( .A(n7182), .B(n7183), .Z(c[108]) );
  NAND U10247 ( .A(n6691), .B(o[108]), .Z(n7183) );
  NAND U10248 ( .A(n6686), .B(creg[108]), .Z(n7182) );
  NAND U10249 ( .A(n7184), .B(n7185), .Z(c[107]) );
  NAND U10250 ( .A(n6691), .B(o[107]), .Z(n7185) );
  NAND U10251 ( .A(n6686), .B(creg[107]), .Z(n7184) );
  NAND U10252 ( .A(n7186), .B(n7187), .Z(c[106]) );
  NAND U10253 ( .A(n6691), .B(o[106]), .Z(n7187) );
  NAND U10254 ( .A(n6686), .B(creg[106]), .Z(n7186) );
  NAND U10255 ( .A(n7188), .B(n7189), .Z(c[105]) );
  NAND U10256 ( .A(n6691), .B(o[105]), .Z(n7189) );
  NAND U10257 ( .A(n6686), .B(creg[105]), .Z(n7188) );
  NAND U10258 ( .A(n7190), .B(n7191), .Z(c[104]) );
  NAND U10259 ( .A(n6691), .B(o[104]), .Z(n7191) );
  NAND U10260 ( .A(n6686), .B(creg[104]), .Z(n7190) );
  NAND U10261 ( .A(n7192), .B(n7193), .Z(c[103]) );
  NAND U10262 ( .A(n6691), .B(o[103]), .Z(n7193) );
  NAND U10263 ( .A(n6686), .B(creg[103]), .Z(n7192) );
  NAND U10264 ( .A(n7194), .B(n7195), .Z(c[102]) );
  NAND U10265 ( .A(n6691), .B(o[102]), .Z(n7195) );
  NAND U10266 ( .A(n6686), .B(creg[102]), .Z(n7194) );
  NAND U10267 ( .A(n7196), .B(n7197), .Z(c[101]) );
  NAND U10268 ( .A(n6691), .B(o[101]), .Z(n7197) );
  NAND U10269 ( .A(n6686), .B(creg[101]), .Z(n7196) );
  NAND U10270 ( .A(n7198), .B(n7199), .Z(c[100]) );
  NAND U10271 ( .A(n6691), .B(o[100]), .Z(n7199) );
  NAND U10272 ( .A(n6686), .B(creg[100]), .Z(n7198) );
  NAND U10273 ( .A(n7200), .B(n7201), .Z(c[0]) );
  NAND U10274 ( .A(n6691), .B(o[0]), .Z(n7201) );
  IV U10275 ( .A(n6686), .Z(n6691) );
  NAND U10276 ( .A(n6686), .B(creg[0]), .Z(n7200) );
  NAND U10277 ( .A(n7202), .B(n7203), .Z(n6686) );
  NANDN U10278 ( .A(ereg[255]), .B(init), .Z(n7203) );
  OR U10279 ( .A(init), .B(e[255]), .Z(n7202) );
endmodule

